module basic_2500_25000_3000_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_467,In_1853);
or U1 (N_1,In_1744,In_1567);
and U2 (N_2,In_293,In_528);
nor U3 (N_3,In_1757,In_897);
and U4 (N_4,In_885,In_937);
nand U5 (N_5,In_1242,In_1137);
nor U6 (N_6,In_1181,In_1706);
nor U7 (N_7,In_1462,In_2387);
nor U8 (N_8,In_874,In_33);
or U9 (N_9,In_1539,In_1285);
nand U10 (N_10,In_1495,In_1351);
or U11 (N_11,In_1445,In_1770);
or U12 (N_12,In_97,In_357);
nor U13 (N_13,In_1374,In_427);
or U14 (N_14,In_1936,In_2135);
and U15 (N_15,In_1662,In_568);
nand U16 (N_16,In_2144,In_1459);
nor U17 (N_17,In_1433,In_758);
xor U18 (N_18,In_1911,In_388);
or U19 (N_19,In_1334,In_798);
xnor U20 (N_20,In_2146,In_173);
or U21 (N_21,In_430,In_1829);
or U22 (N_22,In_285,In_1307);
nor U23 (N_23,In_449,In_2470);
nor U24 (N_24,In_690,In_527);
and U25 (N_25,In_1295,In_678);
nand U26 (N_26,In_2254,In_490);
and U27 (N_27,In_878,In_325);
and U28 (N_28,In_2370,In_1230);
nor U29 (N_29,In_434,In_753);
nor U30 (N_30,In_40,In_978);
and U31 (N_31,In_729,In_1812);
nor U32 (N_32,In_183,In_446);
or U33 (N_33,In_851,In_89);
nor U34 (N_34,In_26,In_86);
nand U35 (N_35,In_537,In_1768);
nor U36 (N_36,In_941,In_801);
nor U37 (N_37,In_942,In_719);
nor U38 (N_38,In_807,In_633);
or U39 (N_39,In_2420,In_2468);
and U40 (N_40,In_811,In_2352);
nor U41 (N_41,In_1160,In_473);
nand U42 (N_42,In_253,In_1650);
xor U43 (N_43,In_2444,In_1405);
nand U44 (N_44,In_628,In_927);
nand U45 (N_45,In_1298,In_1147);
or U46 (N_46,In_1475,In_1625);
xnor U47 (N_47,In_1983,In_2257);
xnor U48 (N_48,In_961,In_267);
nor U49 (N_49,In_737,In_644);
and U50 (N_50,In_862,In_2067);
nor U51 (N_51,In_2455,In_122);
or U52 (N_52,In_19,In_1751);
nand U53 (N_53,In_1600,In_1328);
or U54 (N_54,In_42,In_2175);
and U55 (N_55,In_1860,In_1225);
and U56 (N_56,In_364,In_513);
xor U57 (N_57,In_1886,In_1873);
nor U58 (N_58,In_2103,In_2161);
nand U59 (N_59,In_2162,In_971);
and U60 (N_60,In_2231,In_2125);
or U61 (N_61,In_257,In_410);
and U62 (N_62,In_1320,In_636);
xor U63 (N_63,In_53,In_1244);
nand U64 (N_64,In_1472,In_2339);
or U65 (N_65,In_1721,In_1330);
and U66 (N_66,In_1724,In_134);
and U67 (N_67,In_2378,In_1776);
or U68 (N_68,In_1595,In_128);
or U69 (N_69,In_2082,In_46);
xnor U70 (N_70,In_698,In_91);
nor U71 (N_71,In_853,In_2223);
or U72 (N_72,In_2026,In_457);
and U73 (N_73,In_544,In_6);
or U74 (N_74,In_279,In_308);
or U75 (N_75,In_1274,In_1091);
and U76 (N_76,In_1893,In_1458);
nand U77 (N_77,In_2188,In_1530);
nor U78 (N_78,In_431,In_1191);
and U79 (N_79,In_237,In_1669);
nand U80 (N_80,In_1962,In_451);
nor U81 (N_81,In_1894,In_664);
or U82 (N_82,In_1104,In_1037);
nand U83 (N_83,In_229,In_1221);
and U84 (N_84,In_588,In_893);
nand U85 (N_85,In_1825,In_779);
and U86 (N_86,In_1167,In_1766);
and U87 (N_87,In_1386,In_1813);
nor U88 (N_88,In_1837,In_931);
or U89 (N_89,In_2405,In_2268);
nor U90 (N_90,In_112,In_1193);
and U91 (N_91,In_101,In_368);
and U92 (N_92,In_2438,In_1066);
or U93 (N_93,In_718,In_1960);
or U94 (N_94,In_1814,In_954);
and U95 (N_95,In_1185,In_1196);
nand U96 (N_96,In_71,In_164);
nand U97 (N_97,In_1550,In_1942);
and U98 (N_98,In_830,In_1272);
xor U99 (N_99,In_1831,In_324);
nand U100 (N_100,In_1786,In_2007);
and U101 (N_101,In_2119,In_795);
or U102 (N_102,In_135,In_1856);
and U103 (N_103,In_1933,In_326);
nor U104 (N_104,In_1746,In_981);
xnor U105 (N_105,In_2051,In_1965);
nand U106 (N_106,In_875,In_1769);
nor U107 (N_107,In_1392,In_1881);
nor U108 (N_108,In_2399,In_738);
nor U109 (N_109,In_2418,In_2005);
or U110 (N_110,In_1521,In_13);
and U111 (N_111,In_2105,In_2467);
and U112 (N_112,In_1562,In_1705);
or U113 (N_113,In_369,In_881);
nor U114 (N_114,In_284,In_2475);
and U115 (N_115,In_1948,In_1996);
and U116 (N_116,In_1908,In_1799);
and U117 (N_117,In_2141,In_298);
nand U118 (N_118,In_2099,In_713);
or U119 (N_119,In_1127,In_1093);
and U120 (N_120,In_1577,In_2375);
or U121 (N_121,In_2240,In_1738);
or U122 (N_122,In_381,In_825);
nor U123 (N_123,In_2190,In_2404);
or U124 (N_124,In_1924,In_123);
nor U125 (N_125,In_2213,In_1250);
nor U126 (N_126,In_1531,In_1760);
nor U127 (N_127,In_270,In_549);
or U128 (N_128,In_374,In_76);
and U129 (N_129,In_1419,In_2344);
nand U130 (N_130,In_2351,In_469);
and U131 (N_131,In_1861,In_1581);
and U132 (N_132,In_367,In_294);
nand U133 (N_133,In_579,In_976);
or U134 (N_134,In_500,In_131);
nand U135 (N_135,In_1155,In_1323);
nor U136 (N_136,In_1062,In_1707);
and U137 (N_137,In_2272,In_965);
nor U138 (N_138,In_805,In_1821);
or U139 (N_139,In_2476,In_2073);
and U140 (N_140,In_2250,In_426);
and U141 (N_141,In_1771,In_319);
nand U142 (N_142,In_2021,In_555);
nand U143 (N_143,In_1199,In_697);
nor U144 (N_144,In_2490,In_596);
nand U145 (N_145,In_1851,In_1197);
and U146 (N_146,In_1439,In_432);
and U147 (N_147,In_2143,In_204);
nor U148 (N_148,In_423,In_231);
nand U149 (N_149,In_1465,In_2400);
nor U150 (N_150,In_619,In_439);
and U151 (N_151,In_1761,In_121);
and U152 (N_152,In_37,In_1736);
and U153 (N_153,In_493,In_1229);
nor U154 (N_154,In_919,In_1626);
or U155 (N_155,In_36,In_1442);
or U156 (N_156,In_1002,In_1341);
and U157 (N_157,In_2496,In_1251);
and U158 (N_158,In_625,In_580);
and U159 (N_159,In_967,In_1823);
nand U160 (N_160,In_720,In_924);
and U161 (N_161,In_2140,In_574);
and U162 (N_162,In_2466,In_1178);
and U163 (N_163,In_395,In_750);
nor U164 (N_164,In_309,In_1087);
and U165 (N_165,In_1725,In_2410);
nand U166 (N_166,In_95,In_571);
nor U167 (N_167,In_435,In_607);
or U168 (N_168,In_989,In_1780);
xnor U169 (N_169,In_1114,In_465);
nand U170 (N_170,In_440,In_2178);
xor U171 (N_171,In_1676,In_2227);
nand U172 (N_172,In_988,In_1533);
or U173 (N_173,In_2445,In_1299);
nor U174 (N_174,In_428,In_754);
or U175 (N_175,In_711,In_1362);
and U176 (N_176,In_206,In_70);
and U177 (N_177,In_1943,In_1143);
nor U178 (N_178,In_1205,In_1003);
or U179 (N_179,In_1171,In_559);
nand U180 (N_180,In_458,In_404);
nand U181 (N_181,In_262,In_2171);
nor U182 (N_182,In_1702,In_703);
nor U183 (N_183,In_1399,In_2156);
nand U184 (N_184,In_517,In_2331);
and U185 (N_185,In_2469,In_2300);
or U186 (N_186,In_1249,In_769);
nor U187 (N_187,In_84,In_39);
nor U188 (N_188,In_1556,In_460);
and U189 (N_189,In_721,In_2392);
xor U190 (N_190,In_1028,In_1947);
nor U191 (N_191,In_2487,In_2491);
and U192 (N_192,In_2301,In_1237);
nand U193 (N_193,In_2166,In_1578);
nor U194 (N_194,In_1258,In_987);
nor U195 (N_195,In_154,In_1068);
xor U196 (N_196,In_578,In_2186);
nand U197 (N_197,In_1228,In_340);
or U198 (N_198,In_2308,In_2441);
xor U199 (N_199,In_543,In_845);
and U200 (N_200,In_1880,In_2118);
nand U201 (N_201,In_2292,In_483);
and U202 (N_202,In_2435,In_934);
and U203 (N_203,In_2397,In_2337);
or U204 (N_204,In_85,In_417);
and U205 (N_205,In_2388,In_98);
and U206 (N_206,In_1170,In_1324);
nor U207 (N_207,In_641,In_125);
and U208 (N_208,In_2147,In_386);
nand U209 (N_209,In_2484,In_918);
nor U210 (N_210,In_225,In_1266);
nor U211 (N_211,In_1735,In_320);
or U212 (N_212,In_41,In_288);
nand U213 (N_213,In_2043,In_200);
or U214 (N_214,In_249,In_15);
nor U215 (N_215,In_2041,In_287);
or U216 (N_216,In_497,In_2310);
and U217 (N_217,In_1801,In_561);
nor U218 (N_218,In_870,In_1985);
nand U219 (N_219,In_1796,In_847);
nand U220 (N_220,In_511,In_539);
and U221 (N_221,In_1236,In_1046);
or U222 (N_222,In_1051,In_892);
and U223 (N_223,In_1265,In_389);
nor U224 (N_224,In_133,In_2480);
or U225 (N_225,In_2189,In_1546);
nor U226 (N_226,In_1708,In_1079);
nand U227 (N_227,In_2080,In_2235);
or U228 (N_228,In_531,In_1906);
nand U229 (N_229,In_169,In_1726);
nand U230 (N_230,In_2278,In_1429);
nand U231 (N_231,In_43,In_1292);
nor U232 (N_232,In_1899,In_906);
and U233 (N_233,In_24,In_733);
nand U234 (N_234,In_1594,In_1461);
nor U235 (N_235,In_969,In_1389);
or U236 (N_236,In_1819,In_624);
nand U237 (N_237,In_2002,In_2124);
and U238 (N_238,In_1692,In_215);
nor U239 (N_239,In_932,In_346);
or U240 (N_240,In_510,In_12);
and U241 (N_241,In_1917,In_1105);
and U242 (N_242,In_2004,In_952);
nor U243 (N_243,In_2208,In_2336);
nor U244 (N_244,In_673,In_1510);
nor U245 (N_245,In_2245,In_692);
nand U246 (N_246,In_1930,In_419);
nor U247 (N_247,In_182,In_1077);
and U248 (N_248,In_258,In_356);
nor U249 (N_249,In_1756,In_478);
nor U250 (N_250,In_2229,In_2053);
or U251 (N_251,In_1593,In_546);
or U252 (N_252,In_1050,In_1779);
or U253 (N_253,In_360,In_998);
nor U254 (N_254,In_2111,In_1226);
or U255 (N_255,In_1551,In_2039);
xnor U256 (N_256,In_1060,In_1280);
nand U257 (N_257,In_353,In_2032);
nor U258 (N_258,In_796,In_1407);
nor U259 (N_259,In_1503,In_1496);
nor U260 (N_260,In_727,In_2120);
or U261 (N_261,In_1762,In_663);
nor U262 (N_262,In_2133,In_1640);
or U263 (N_263,In_216,In_1219);
nor U264 (N_264,In_1246,In_382);
nand U265 (N_265,In_2389,In_522);
and U266 (N_266,In_659,In_2282);
xor U267 (N_267,In_1214,In_2411);
nand U268 (N_268,In_2197,In_1234);
and U269 (N_269,In_1076,In_1014);
or U270 (N_270,In_1264,In_1587);
nor U271 (N_271,In_1984,In_1279);
and U272 (N_272,In_212,In_75);
or U273 (N_273,In_1381,In_749);
nand U274 (N_274,In_1345,In_476);
and U275 (N_275,In_2325,In_463);
nand U276 (N_276,In_1333,In_2176);
and U277 (N_277,In_1281,In_72);
and U278 (N_278,In_2277,In_366);
or U279 (N_279,In_953,In_709);
and U280 (N_280,In_1806,In_226);
nor U281 (N_281,In_2371,In_2068);
nand U282 (N_282,In_1565,In_1869);
nand U283 (N_283,In_806,In_512);
nand U284 (N_284,In_1053,In_1968);
nor U285 (N_285,In_917,In_1652);
or U286 (N_286,In_1490,In_1332);
or U287 (N_287,In_2341,In_1103);
or U288 (N_288,In_722,In_1343);
and U289 (N_289,In_492,In_2035);
or U290 (N_290,In_150,In_2194);
or U291 (N_291,In_929,In_301);
nand U292 (N_292,In_371,In_790);
nand U293 (N_293,In_1891,In_909);
or U294 (N_294,In_841,In_1287);
nand U295 (N_295,In_1056,In_2107);
nor U296 (N_296,In_305,In_2377);
or U297 (N_297,In_1356,In_2233);
nor U298 (N_298,In_2309,In_1291);
nand U299 (N_299,In_1455,In_116);
xnor U300 (N_300,In_1576,In_2362);
nand U301 (N_301,In_1732,In_1142);
xnor U302 (N_302,In_418,In_1207);
nand U303 (N_303,In_387,In_627);
and U304 (N_304,In_1646,In_997);
nand U305 (N_305,In_425,In_278);
and U306 (N_306,In_2038,In_2131);
or U307 (N_307,In_1457,In_2409);
and U308 (N_308,In_1108,In_973);
nor U309 (N_309,In_1271,In_2137);
nor U310 (N_310,In_1019,In_1359);
or U311 (N_311,In_1741,In_877);
or U312 (N_312,In_1651,In_1540);
nand U313 (N_313,In_1492,In_1951);
nand U314 (N_314,In_1921,In_2092);
or U315 (N_315,In_349,In_281);
nand U316 (N_316,In_1635,In_1119);
nand U317 (N_317,In_323,In_534);
nand U318 (N_318,In_1470,In_264);
or U319 (N_319,In_705,In_694);
nor U320 (N_320,In_612,In_1634);
nand U321 (N_321,In_495,In_2184);
and U322 (N_322,In_773,In_2203);
and U323 (N_323,In_858,In_2323);
nand U324 (N_324,In_774,In_2207);
or U325 (N_325,In_1717,In_1730);
or U326 (N_326,In_900,In_563);
xor U327 (N_327,In_902,In_637);
and U328 (N_328,In_2173,In_2440);
or U329 (N_329,In_2001,In_1876);
and U330 (N_330,In_2328,In_2181);
and U331 (N_331,In_1179,In_876);
and U332 (N_332,In_746,In_1665);
nand U333 (N_333,In_259,In_1310);
nand U334 (N_334,In_2211,In_1448);
or U335 (N_335,In_2474,In_1052);
nor U336 (N_336,In_455,In_250);
nor U337 (N_337,In_2047,In_1585);
nor U338 (N_338,In_1004,In_1859);
or U339 (N_339,In_1146,In_1413);
nor U340 (N_340,In_1346,In_1690);
nand U341 (N_341,In_794,In_744);
nor U342 (N_342,In_1605,In_129);
or U343 (N_343,In_321,In_159);
or U344 (N_344,In_370,In_195);
or U345 (N_345,In_1945,In_90);
or U346 (N_346,In_1609,In_2210);
or U347 (N_347,In_1248,In_1628);
nor U348 (N_348,In_1339,In_1875);
nand U349 (N_349,In_2322,In_105);
or U350 (N_350,In_1570,In_1532);
or U351 (N_351,In_652,In_1139);
and U352 (N_352,In_2366,In_2094);
or U353 (N_353,In_1005,In_922);
or U354 (N_354,In_2183,In_1542);
nor U355 (N_355,In_1522,In_838);
xor U356 (N_356,In_2413,In_1866);
nand U357 (N_357,In_1558,In_1376);
nand U358 (N_358,In_1603,In_2066);
or U359 (N_359,In_1569,In_2030);
or U360 (N_360,In_274,In_1239);
xnor U361 (N_361,In_1745,In_951);
nand U362 (N_362,In_487,In_1306);
or U363 (N_363,In_1422,In_1807);
and U364 (N_364,In_824,In_634);
or U365 (N_365,In_1101,In_93);
or U366 (N_366,In_127,In_2429);
nor U367 (N_367,In_2084,In_2011);
nor U368 (N_368,In_148,In_843);
nand U369 (N_369,In_896,In_1506);
nor U370 (N_370,In_2369,In_1180);
nor U371 (N_371,In_1254,In_2456);
or U372 (N_372,In_2307,In_1607);
nor U373 (N_373,In_963,In_2372);
and U374 (N_374,In_728,In_1957);
and U375 (N_375,In_180,In_1024);
nand U376 (N_376,In_1820,In_861);
xor U377 (N_377,In_2033,In_1293);
or U378 (N_378,In_1253,In_1526);
nand U379 (N_379,In_584,In_2477);
nand U380 (N_380,In_1840,In_303);
and U381 (N_381,In_295,In_1703);
or U382 (N_382,In_178,In_448);
or U383 (N_383,In_1009,In_1846);
nand U384 (N_384,In_142,In_1549);
and U385 (N_385,In_974,In_1358);
and U386 (N_386,In_1063,In_479);
or U387 (N_387,In_1728,In_111);
and U388 (N_388,In_1141,In_251);
or U389 (N_389,In_1391,In_984);
nor U390 (N_390,In_1710,In_2158);
nor U391 (N_391,In_1308,In_409);
xor U392 (N_392,In_158,In_1660);
or U393 (N_393,In_810,In_403);
nand U394 (N_394,In_660,In_181);
or U395 (N_395,In_1203,In_2269);
or U396 (N_396,In_1102,In_1591);
nor U397 (N_397,In_940,In_100);
nand U398 (N_398,In_1109,In_1410);
nand U399 (N_399,In_545,In_868);
nor U400 (N_400,In_291,In_943);
nand U401 (N_401,In_2015,In_1126);
nor U402 (N_402,In_2354,In_1067);
nor U403 (N_403,In_1713,In_130);
nor U404 (N_404,In_1689,In_704);
nor U405 (N_405,In_863,In_1054);
xor U406 (N_406,In_422,In_1035);
nor U407 (N_407,In_1502,In_926);
and U408 (N_408,In_1504,In_1304);
nand U409 (N_409,In_1431,In_839);
nand U410 (N_410,In_187,In_23);
nor U411 (N_411,In_681,In_2110);
nor U412 (N_412,In_411,In_189);
and U413 (N_413,In_157,In_2017);
nor U414 (N_414,In_840,In_1666);
or U415 (N_415,In_1120,In_2303);
nor U416 (N_416,In_526,In_28);
nor U417 (N_417,In_1447,In_499);
nor U418 (N_418,In_2408,In_211);
nand U419 (N_419,In_92,In_759);
and U420 (N_420,In_2316,In_856);
nand U421 (N_421,In_2382,In_508);
nor U422 (N_422,In_1973,In_2020);
nor U423 (N_423,In_2312,In_1709);
nor U424 (N_424,In_307,In_1283);
nor U425 (N_425,In_1377,In_1497);
nand U426 (N_426,In_342,In_1424);
or U427 (N_427,In_1697,In_2174);
or U428 (N_428,In_1017,In_2010);
and U429 (N_429,In_2267,In_1566);
or U430 (N_430,In_1696,In_668);
nor U431 (N_431,In_156,In_760);
or U432 (N_432,In_67,In_1560);
nor U433 (N_433,In_1110,In_1029);
or U434 (N_434,In_1564,In_1427);
nand U435 (N_435,In_81,In_1773);
nand U436 (N_436,In_1694,In_2342);
and U437 (N_437,In_1255,In_2464);
or U438 (N_438,In_1064,In_1509);
or U439 (N_439,In_421,In_777);
and U440 (N_440,In_126,In_252);
nor U441 (N_441,In_530,In_640);
or U442 (N_442,In_1959,In_2070);
xnor U443 (N_443,In_152,In_1486);
and U444 (N_444,In_59,In_725);
nor U445 (N_445,In_2136,In_272);
and U446 (N_446,In_1493,In_2165);
nand U447 (N_447,In_762,In_1342);
or U448 (N_448,In_1241,In_666);
and U449 (N_449,In_827,In_1602);
nand U450 (N_450,In_199,In_907);
and U451 (N_451,In_322,In_363);
nor U452 (N_452,In_821,In_1897);
and U453 (N_453,In_1647,In_2494);
nand U454 (N_454,In_1300,In_2048);
nor U455 (N_455,In_2034,In_27);
and U456 (N_456,In_2473,In_350);
nor U457 (N_457,In_238,In_1286);
nand U458 (N_458,In_1030,In_2074);
or U459 (N_459,In_1739,In_866);
and U460 (N_460,In_1568,In_2044);
or U461 (N_461,In_1808,In_1775);
nand U462 (N_462,In_1387,In_2139);
nor U463 (N_463,In_593,In_1619);
or U464 (N_464,In_223,In_1123);
nand U465 (N_465,In_2391,In_1245);
nor U466 (N_466,In_1210,In_1044);
nand U467 (N_467,In_1150,In_2390);
or U468 (N_468,In_2234,In_1608);
and U469 (N_469,In_2416,In_2115);
and U470 (N_470,In_175,In_677);
nand U471 (N_471,In_1369,In_1798);
nand U472 (N_472,In_1670,In_819);
or U473 (N_473,In_1890,In_1072);
nor U474 (N_474,In_4,In_1731);
or U475 (N_475,In_831,In_1220);
nor U476 (N_476,In_2395,In_2152);
and U477 (N_477,In_1477,In_748);
nand U478 (N_478,In_514,In_1033);
or U479 (N_479,In_797,In_755);
or U480 (N_480,In_1976,In_64);
nand U481 (N_481,In_1797,In_2338);
nor U482 (N_482,In_1999,In_2142);
nor U483 (N_483,In_2355,In_602);
nor U484 (N_484,In_51,In_1481);
nor U485 (N_485,In_1482,In_1588);
or U486 (N_486,In_203,In_535);
and U487 (N_487,In_768,In_1294);
nand U488 (N_488,In_1073,In_1096);
nor U489 (N_489,In_502,In_2315);
or U490 (N_490,In_2014,In_609);
and U491 (N_491,In_1303,In_2381);
or U492 (N_492,In_1733,In_83);
nand U493 (N_493,In_1367,In_1130);
and U494 (N_494,In_1722,In_935);
or U495 (N_495,In_1879,In_1473);
nor U496 (N_496,In_2126,In_2205);
nor U497 (N_497,In_1518,In_2083);
nor U498 (N_498,In_977,In_1058);
nand U499 (N_499,In_726,In_1015);
and U500 (N_500,In_814,In_1681);
nand U501 (N_501,In_2195,In_1136);
nor U502 (N_502,In_1049,In_2081);
or U503 (N_503,In_207,In_2290);
xor U504 (N_504,In_1488,In_1355);
or U505 (N_505,In_1896,In_1528);
nand U506 (N_506,In_1070,In_699);
or U507 (N_507,In_466,In_194);
or U508 (N_508,In_1094,In_167);
nand U509 (N_509,In_489,In_2465);
or U510 (N_510,In_1997,In_1107);
nor U511 (N_511,In_2028,In_836);
nand U512 (N_512,In_1946,In_2122);
and U513 (N_513,In_611,In_1855);
nand U514 (N_514,In_1397,In_327);
nand U515 (N_515,In_1252,In_1041);
nand U516 (N_516,In_519,In_1464);
nor U517 (N_517,In_147,In_2275);
nand U518 (N_518,In_334,In_683);
nand U519 (N_519,In_114,In_747);
or U520 (N_520,In_415,In_1836);
nand U521 (N_521,In_35,In_2498);
and U522 (N_522,In_1699,In_5);
and U523 (N_523,In_424,In_2148);
nor U524 (N_524,In_889,In_151);
xnor U525 (N_525,In_1366,In_1641);
xor U526 (N_526,In_372,In_2478);
nand U527 (N_527,In_515,In_617);
nor U528 (N_528,In_1520,In_2423);
and U529 (N_529,In_1157,In_2398);
nand U530 (N_530,In_1128,In_1479);
nand U531 (N_531,In_701,In_1514);
or U532 (N_532,In_506,In_1315);
nand U533 (N_533,In_783,In_1277);
nand U534 (N_534,In_1729,In_280);
and U535 (N_535,In_2116,In_550);
or U536 (N_536,In_899,In_2252);
or U537 (N_537,In_1584,In_1038);
and U538 (N_538,In_2485,In_1572);
or U539 (N_539,In_2169,In_1231);
and U540 (N_540,In_104,In_1432);
and U541 (N_541,In_646,In_1852);
and U542 (N_542,In_260,In_1571);
or U543 (N_543,In_438,In_192);
or U544 (N_544,In_2072,In_828);
nand U545 (N_545,In_865,In_2360);
or U546 (N_546,In_864,In_2209);
nor U547 (N_547,In_2128,In_11);
and U548 (N_548,In_1348,In_276);
nand U549 (N_549,In_375,In_542);
or U550 (N_550,In_854,In_2076);
and U551 (N_551,In_1750,In_1671);
nand U552 (N_552,In_1329,In_1742);
or U553 (N_553,In_2164,In_2151);
or U554 (N_554,In_708,In_1451);
nand U555 (N_555,In_1867,In_1240);
nand U556 (N_556,In_2317,In_2220);
or U557 (N_557,In_1057,In_576);
nor U558 (N_558,In_66,In_1222);
nor U559 (N_559,In_220,In_1525);
xor U560 (N_560,In_775,In_2138);
xnor U561 (N_561,In_1878,In_557);
and U562 (N_562,In_1273,In_3);
nand U563 (N_563,In_339,In_1512);
nor U564 (N_564,In_995,In_1508);
nand U565 (N_565,In_338,In_236);
or U566 (N_566,In_1679,In_1289);
nand U567 (N_567,In_1026,In_261);
or U568 (N_568,In_21,In_964);
and U569 (N_569,In_1624,In_1400);
and U570 (N_570,In_911,In_1887);
nor U571 (N_571,In_143,In_645);
nand U572 (N_572,In_1988,In_1599);
nor U573 (N_573,In_1922,In_1805);
and U574 (N_574,In_184,In_1971);
and U575 (N_575,In_1085,In_908);
nand U576 (N_576,In_275,In_672);
or U577 (N_577,In_1791,In_494);
and U578 (N_578,In_503,In_842);
or U579 (N_579,In_1169,In_1900);
or U580 (N_580,In_2170,In_406);
nand U581 (N_581,In_29,In_1316);
or U582 (N_582,In_1187,In_1872);
nor U583 (N_583,In_1611,In_1858);
or U584 (N_584,In_329,In_1753);
nor U585 (N_585,In_1685,In_1688);
or U586 (N_586,In_1135,In_2318);
nor U587 (N_587,In_399,In_582);
nor U588 (N_588,In_1261,In_1554);
or U589 (N_589,In_119,In_2396);
nor U590 (N_590,In_1618,In_344);
nor U591 (N_591,In_2086,In_365);
or U592 (N_592,In_1275,In_994);
or U593 (N_593,In_1190,In_1672);
nand U594 (N_594,In_1450,In_2452);
nand U595 (N_595,In_740,In_2394);
and U596 (N_596,In_1408,In_916);
nand U597 (N_597,In_741,In_1124);
xor U598 (N_598,In_551,In_1006);
and U599 (N_599,In_1215,In_1916);
and U600 (N_600,In_402,In_1974);
nor U601 (N_601,In_1966,In_1443);
nand U602 (N_602,In_1013,In_883);
nand U603 (N_603,In_475,In_572);
or U604 (N_604,In_176,In_1826);
or U605 (N_605,In_68,In_2442);
and U606 (N_606,In_2199,In_1010);
nand U607 (N_607,In_2459,In_2281);
nand U608 (N_608,In_2291,In_2449);
and U609 (N_609,In_1284,In_1793);
and U610 (N_610,In_2299,In_731);
nor U611 (N_611,In_771,In_2261);
or U612 (N_612,In_1818,In_2499);
nor U613 (N_613,In_2129,In_1347);
nor U614 (N_614,In_2305,In_1574);
nor U615 (N_615,In_1772,In_1767);
and U616 (N_616,In_1684,In_1099);
and U617 (N_617,In_1537,In_700);
nand U618 (N_618,In_1370,In_1501);
nor U619 (N_619,In_992,In_848);
xnor U620 (N_620,In_1469,In_263);
or U621 (N_621,In_2095,In_1617);
and U622 (N_622,In_554,In_2090);
nand U623 (N_623,In_233,In_591);
or U624 (N_624,In_2238,In_390);
nand U625 (N_625,In_408,In_1478);
or U626 (N_626,In_1610,In_804);
or U627 (N_627,In_669,In_1269);
nor U628 (N_628,In_2472,In_716);
nand U629 (N_629,In_1941,In_1944);
nor U630 (N_630,In_1835,In_1373);
nor U631 (N_631,In_1716,In_283);
and U632 (N_632,In_910,In_394);
and U633 (N_633,In_1969,In_2289);
and U634 (N_634,In_986,In_1174);
or U635 (N_635,In_2471,In_635);
and U636 (N_636,In_1235,In_2012);
nor U637 (N_637,In_498,In_826);
nor U638 (N_638,In_2460,In_944);
or U639 (N_639,In_58,In_1082);
nand U640 (N_640,In_454,In_1485);
xor U641 (N_641,In_1583,In_1202);
or U642 (N_642,In_1888,In_1597);
and U643 (N_643,In_352,In_1877);
nand U644 (N_644,In_2177,In_1555);
nor U645 (N_645,In_1515,In_936);
nor U646 (N_646,In_377,In_960);
nor U647 (N_647,In_1327,In_416);
or U648 (N_648,In_396,In_647);
nand U649 (N_649,In_990,In_1);
or U650 (N_650,In_2433,In_400);
or U651 (N_651,In_1045,In_1350);
and U652 (N_652,In_452,In_879);
and U653 (N_653,In_1256,In_2180);
and U654 (N_654,In_1749,In_2349);
nand U655 (N_655,In_1952,In_1517);
nand U656 (N_656,In_536,In_570);
nand U657 (N_657,In_62,In_2160);
nand U658 (N_658,In_1711,In_1553);
nand U659 (N_659,In_197,In_315);
nor U660 (N_660,In_643,In_1950);
nor U661 (N_661,In_1257,In_1204);
or U662 (N_662,In_577,In_1993);
or U663 (N_663,In_662,In_52);
or U664 (N_664,In_241,In_2045);
nor U665 (N_665,In_1613,In_757);
xor U666 (N_666,In_480,In_1216);
or U667 (N_667,In_132,In_955);
or U668 (N_668,In_915,In_1121);
or U669 (N_669,In_1080,In_541);
xnor U670 (N_670,In_2258,In_1939);
nor U671 (N_671,In_1401,In_393);
nor U672 (N_672,In_74,In_631);
nand U673 (N_673,In_1718,In_1832);
and U674 (N_674,In_2000,In_778);
nor U675 (N_675,In_1027,In_149);
nand U676 (N_676,In_2285,In_653);
and U677 (N_677,In_2302,In_2350);
nand U678 (N_678,In_1403,In_2274);
xor U679 (N_679,In_2324,In_61);
nand U680 (N_680,In_950,In_484);
xor U681 (N_681,In_2191,In_174);
nand U682 (N_682,In_1040,In_706);
and U683 (N_683,In_1276,In_985);
nor U684 (N_684,In_2373,In_2424);
or U685 (N_685,In_1385,In_1787);
and U686 (N_686,In_115,In_1227);
nor U687 (N_687,In_835,In_2306);
nor U688 (N_688,In_1474,In_2376);
xnor U689 (N_689,In_2270,In_2439);
nand U690 (N_690,In_1484,In_504);
nor U691 (N_691,In_2481,In_696);
or U692 (N_692,In_336,In_560);
nor U693 (N_693,In_834,In_445);
nor U694 (N_694,In_2434,In_949);
nor U695 (N_695,In_2488,In_145);
or U696 (N_696,In_335,In_1932);
nand U697 (N_697,In_799,In_891);
nor U698 (N_698,In_957,In_347);
and U699 (N_699,In_714,In_1809);
nand U700 (N_700,In_2088,In_1441);
nand U701 (N_701,In_1357,In_1036);
and U702 (N_702,In_65,In_1654);
nor U703 (N_703,In_1949,In_2006);
and U704 (N_704,In_1200,In_1854);
nor U705 (N_705,In_2153,In_859);
or U706 (N_706,In_2271,In_1489);
or U707 (N_707,In_1217,In_829);
and U708 (N_708,In_1644,In_1663);
nor U709 (N_709,In_1209,In_2264);
and U710 (N_710,In_2486,In_345);
and U711 (N_711,In_595,In_1788);
nor U712 (N_712,In_1168,In_1326);
nor U713 (N_713,In_110,In_2430);
nand U714 (N_714,In_781,In_470);
and U715 (N_715,In_1926,In_1870);
nor U716 (N_716,In_243,In_2448);
nor U717 (N_717,In_49,In_1981);
nor U718 (N_718,In_1561,In_1092);
xnor U719 (N_719,In_193,In_109);
and U720 (N_720,In_2332,In_1129);
and U721 (N_721,In_2321,In_1601);
nand U722 (N_722,In_1631,In_1428);
or U723 (N_723,In_518,In_656);
nor U724 (N_724,In_1892,In_1606);
or U725 (N_725,In_605,In_1811);
or U726 (N_726,In_880,In_1259);
nand U727 (N_727,In_1331,In_832);
or U728 (N_728,In_975,In_1655);
or U729 (N_729,In_464,In_54);
nand U730 (N_730,In_2242,In_1804);
nand U731 (N_731,In_1075,In_2367);
and U732 (N_732,In_743,In_242);
nand U733 (N_733,In_311,In_1695);
nor U734 (N_734,In_752,In_1305);
and U735 (N_735,In_2348,In_2100);
and U736 (N_736,In_354,In_2123);
and U737 (N_737,In_1792,In_564);
and U738 (N_738,In_1789,In_2364);
nand U739 (N_739,In_1675,In_1012);
or U740 (N_740,In_2359,In_1632);
nand U741 (N_741,In_846,In_1164);
nor U742 (N_742,In_923,In_1838);
nor U743 (N_743,In_792,In_1083);
or U744 (N_744,In_1582,In_277);
or U745 (N_745,In_1186,In_2432);
nand U746 (N_746,In_1383,In_565);
nand U747 (N_747,In_1955,In_548);
and U748 (N_748,In_616,In_1415);
or U749 (N_749,In_1149,In_1848);
and U750 (N_750,In_1822,In_318);
or U751 (N_751,In_407,In_485);
and U752 (N_752,In_1008,In_1483);
or U753 (N_753,In_172,In_688);
and U754 (N_754,In_1314,In_1964);
and U755 (N_755,In_1777,In_676);
and U756 (N_756,In_1816,In_671);
or U757 (N_757,In_1198,In_1627);
nand U758 (N_758,In_1523,In_613);
nor U759 (N_759,In_1309,In_1545);
and U760 (N_760,In_2241,In_1925);
nand U761 (N_761,In_736,In_1884);
or U762 (N_762,In_1380,In_2427);
or U763 (N_763,In_2217,In_124);
and U764 (N_764,In_2365,In_1622);
nor U765 (N_765,In_1842,In_1991);
nand U766 (N_766,In_1755,In_933);
or U767 (N_767,In_1547,In_1025);
or U768 (N_768,In_437,In_2451);
and U769 (N_769,In_1325,In_2091);
or U770 (N_770,In_1638,In_234);
and U771 (N_771,In_1039,In_852);
nor U772 (N_772,In_1543,In_2057);
or U773 (N_773,In_615,In_1267);
and U774 (N_774,In_1363,In_1420);
nor U775 (N_775,In_1071,In_2079);
or U776 (N_776,In_343,In_785);
or U777 (N_777,In_928,In_255);
nor U778 (N_778,In_1586,In_108);
and U779 (N_779,In_1302,In_2216);
nor U780 (N_780,In_2172,In_1471);
or U781 (N_781,In_2255,In_1368);
or U782 (N_782,In_599,In_1460);
and U783 (N_783,In_2461,In_2069);
xor U784 (N_784,In_1857,In_1453);
and U785 (N_785,In_385,In_1794);
or U786 (N_786,In_1633,In_88);
or U787 (N_787,In_1156,In_1406);
or U788 (N_788,In_140,In_898);
nand U789 (N_789,In_2236,In_946);
nand U790 (N_790,In_2206,In_373);
nor U791 (N_791,In_1112,In_702);
and U792 (N_792,In_453,In_1938);
nor U793 (N_793,In_397,In_650);
or U794 (N_794,In_1183,In_1935);
nor U795 (N_795,In_639,In_618);
or U796 (N_796,In_8,In_1673);
nand U797 (N_797,In_265,In_2251);
and U798 (N_798,In_1290,In_592);
nand U799 (N_799,In_219,In_2109);
or U800 (N_800,In_1589,In_1616);
and U801 (N_801,In_2293,In_1648);
nor U802 (N_802,In_1604,In_1499);
and U803 (N_803,In_82,In_18);
nor U804 (N_804,In_632,In_1425);
or U805 (N_805,In_57,In_614);
or U806 (N_806,In_1620,In_2062);
or U807 (N_807,In_1151,In_1904);
or U808 (N_808,In_1700,In_217);
nand U809 (N_809,In_800,In_1579);
nor U810 (N_810,In_1923,In_1195);
nand U811 (N_811,In_903,In_482);
and U812 (N_812,In_815,In_2296);
nand U813 (N_813,In_106,In_1782);
and U814 (N_814,In_179,In_78);
and U815 (N_815,In_1165,In_1158);
nor U816 (N_816,In_2426,In_938);
nor U817 (N_817,In_2345,In_2393);
or U818 (N_818,In_1995,In_1452);
nand U819 (N_819,In_447,In_2042);
or U820 (N_820,In_2096,In_818);
nor U821 (N_821,In_405,In_1903);
nand U822 (N_822,In_351,In_1833);
nor U823 (N_823,In_675,In_25);
or U824 (N_824,In_1182,In_1153);
nor U825 (N_825,In_1642,In_1232);
nor U826 (N_826,In_1764,In_2428);
nand U827 (N_827,In_655,In_247);
or U828 (N_828,In_2121,In_1544);
and U829 (N_829,In_2482,In_930);
nor U830 (N_830,In_820,In_398);
and U831 (N_831,In_103,In_1352);
or U832 (N_832,In_501,In_2247);
and U833 (N_833,In_767,In_763);
nor U834 (N_834,In_1541,In_73);
nor U835 (N_835,In_674,In_1340);
nand U836 (N_836,In_2385,In_1727);
and U837 (N_837,In_505,In_1783);
and U838 (N_838,In_471,In_1580);
or U839 (N_839,In_523,In_297);
nor U840 (N_840,In_710,In_1111);
or U841 (N_841,In_2112,In_118);
nand U842 (N_842,In_0,In_837);
or U843 (N_843,In_230,In_136);
nor U844 (N_844,In_2061,In_2025);
or U845 (N_845,In_2117,In_533);
or U846 (N_846,In_60,In_2077);
and U847 (N_847,In_218,In_391);
or U848 (N_848,In_2029,In_31);
nand U849 (N_849,In_707,In_2202);
and U850 (N_850,In_520,In_1910);
and U851 (N_851,In_948,In_844);
or U852 (N_852,In_2108,In_1138);
nand U853 (N_853,In_2379,In_2446);
nor U854 (N_854,In_196,In_1667);
nand U855 (N_855,In_2243,In_273);
and U856 (N_856,In_1394,In_328);
or U857 (N_857,In_1335,In_120);
and U858 (N_858,In_1296,In_780);
nand U859 (N_859,In_925,In_442);
and U860 (N_860,In_629,In_1132);
or U861 (N_861,In_1018,In_654);
or U862 (N_862,In_855,In_300);
and U863 (N_863,In_2054,In_2221);
and U864 (N_864,In_1830,In_2497);
and U865 (N_865,In_2248,In_1687);
nand U866 (N_866,In_2023,In_687);
or U867 (N_867,In_914,In_1636);
or U868 (N_868,In_380,In_715);
nand U869 (N_869,In_2295,In_153);
or U870 (N_870,In_341,In_1061);
or U871 (N_871,In_1042,In_1865);
and U872 (N_872,In_2085,In_2330);
nor U873 (N_873,In_553,In_1774);
nor U874 (N_874,In_1172,In_1436);
or U875 (N_875,In_2215,In_80);
nor U876 (N_876,In_69,In_648);
xnor U877 (N_877,In_1683,In_1388);
or U878 (N_878,In_1423,In_1529);
or U879 (N_879,In_1714,In_1095);
or U880 (N_880,In_751,In_461);
nand U881 (N_881,In_1417,In_102);
and U882 (N_882,In_1524,In_982);
nor U883 (N_883,In_2193,In_1864);
and U884 (N_884,In_2022,In_312);
nand U885 (N_885,In_1630,In_962);
nand U886 (N_886,In_79,In_1972);
nor U887 (N_887,In_2056,In_2150);
nand U888 (N_888,In_1734,In_1089);
nand U889 (N_889,In_137,In_2078);
and U890 (N_890,In_459,In_2340);
or U891 (N_891,In_802,In_1778);
or U892 (N_892,In_966,In_1698);
nand U893 (N_893,In_1790,In_573);
and U894 (N_894,In_598,In_2168);
nand U895 (N_895,In_1763,In_496);
xor U896 (N_896,In_1177,In_1021);
and U897 (N_897,In_723,In_32);
and U898 (N_898,In_412,In_1319);
or U899 (N_899,In_1444,In_895);
nor U900 (N_900,In_793,In_2225);
and U901 (N_901,In_2287,In_1653);
and U902 (N_902,In_1844,In_850);
nor U903 (N_903,In_2,In_1847);
or U904 (N_904,In_16,In_547);
xnor U905 (N_905,In_1889,In_2263);
or U906 (N_906,In_833,In_2027);
or U907 (N_907,In_472,In_1312);
nand U908 (N_908,In_1527,In_524);
nor U909 (N_909,In_170,In_630);
or U910 (N_910,In_1321,In_286);
nand U911 (N_911,In_1435,In_441);
nor U912 (N_912,In_107,In_477);
nor U913 (N_913,In_516,In_2063);
nor U914 (N_914,In_788,In_1557);
nor U915 (N_915,In_1915,In_1592);
or U916 (N_916,In_1322,In_362);
nand U917 (N_917,In_486,In_638);
nor U918 (N_918,In_2232,In_7);
and U919 (N_919,In_56,In_739);
and U920 (N_920,In_146,In_956);
or U921 (N_921,In_1480,In_764);
nor U922 (N_922,In_1173,In_2273);
nor U923 (N_923,In_2230,In_1885);
and U924 (N_924,In_2256,In_1491);
nor U925 (N_925,In_1970,In_289);
nor U926 (N_926,In_1396,In_2008);
nor U927 (N_927,In_1288,In_1022);
nand U928 (N_928,In_585,In_2450);
or U929 (N_929,In_606,In_2326);
nand U930 (N_930,In_1883,In_474);
or U931 (N_931,In_1979,In_198);
and U932 (N_932,In_1839,In_857);
and U933 (N_933,In_1931,In_1133);
and U934 (N_934,In_1691,In_48);
nand U935 (N_935,In_2113,In_1901);
and U936 (N_936,In_2415,In_603);
nand U937 (N_937,In_620,In_113);
nand U938 (N_938,In_2368,In_2334);
or U939 (N_939,In_1426,In_1643);
nor U940 (N_940,In_1361,In_2458);
and U941 (N_941,In_2419,In_1118);
or U942 (N_942,In_2163,In_2358);
and U943 (N_943,In_208,In_1055);
and U944 (N_944,In_1353,In_468);
or U945 (N_945,In_1994,In_867);
or U946 (N_946,In_1260,In_525);
nand U947 (N_947,In_784,In_1411);
nand U948 (N_948,In_1000,In_886);
nor U949 (N_949,In_1134,In_665);
or U950 (N_950,In_913,In_809);
and U951 (N_951,In_959,In_1463);
and U952 (N_952,In_2253,In_1693);
nand U953 (N_953,In_1048,In_1098);
nor U954 (N_954,In_256,In_47);
or U955 (N_955,In_2196,In_246);
nor U956 (N_956,In_316,In_2288);
and U957 (N_957,In_299,In_1987);
nor U958 (N_958,In_2314,In_1047);
nand U959 (N_959,In_1031,In_433);
and U960 (N_960,In_972,In_2417);
and U961 (N_961,In_1536,In_2276);
nor U962 (N_962,In_1507,In_1430);
nand U963 (N_963,In_282,In_717);
nor U964 (N_964,In_1349,In_163);
or U965 (N_965,In_1224,In_689);
nand U966 (N_966,In_2187,In_968);
and U967 (N_967,In_1117,In_589);
or U968 (N_968,In_695,In_2425);
nand U969 (N_969,In_1871,In_2246);
nand U970 (N_970,In_1645,In_1747);
or U971 (N_971,In_1723,In_1704);
or U972 (N_972,In_205,In_1843);
or U973 (N_973,In_2298,In_191);
or U974 (N_974,In_787,In_2214);
and U975 (N_975,In_392,In_2453);
nor U976 (N_976,In_1152,In_1337);
and U977 (N_977,In_1548,In_444);
nor U978 (N_978,In_1466,In_2401);
nor U979 (N_979,In_443,In_601);
nor U980 (N_980,In_1317,In_224);
nor U981 (N_981,In_1032,In_1449);
nor U982 (N_982,In_2431,In_2104);
nand U983 (N_983,In_745,In_2106);
and U984 (N_984,In_1715,In_849);
or U985 (N_985,In_2283,In_1678);
or U986 (N_986,In_2266,In_420);
and U987 (N_987,In_770,In_2361);
and U988 (N_988,In_38,In_254);
nor U989 (N_989,In_1212,In_888);
or U990 (N_990,In_2049,In_567);
nand U991 (N_991,In_2130,In_188);
or U992 (N_992,In_887,In_14);
and U993 (N_993,In_1639,In_1113);
nand U994 (N_994,In_1680,In_1815);
nor U995 (N_995,In_921,In_1827);
nor U996 (N_996,In_1563,In_1122);
or U997 (N_997,In_144,In_558);
or U998 (N_998,In_904,In_413);
or U999 (N_999,In_304,In_1958);
or U1000 (N_1000,In_355,In_1086);
nor U1001 (N_1001,In_2265,In_594);
or U1002 (N_1002,In_912,In_1505);
nand U1003 (N_1003,In_1498,In_10);
and U1004 (N_1004,In_1023,In_1404);
or U1005 (N_1005,In_2249,In_1078);
or U1006 (N_1006,In_2159,In_2075);
and U1007 (N_1007,In_2055,In_1937);
and U1008 (N_1008,In_1011,In_776);
nor U1009 (N_1009,In_117,In_2402);
nor U1010 (N_1010,In_2237,In_138);
xnor U1011 (N_1011,In_1412,In_766);
nor U1012 (N_1012,In_2114,In_1573);
and U1013 (N_1013,In_456,In_2060);
nand U1014 (N_1014,In_348,In_450);
or U1015 (N_1015,In_871,In_45);
or U1016 (N_1016,In_901,In_96);
or U1017 (N_1017,In_22,In_1919);
and U1018 (N_1018,In_1849,In_761);
nand U1019 (N_1019,In_1596,In_2320);
nor U1020 (N_1020,In_575,In_562);
nand U1021 (N_1021,In_1233,In_1914);
or U1022 (N_1022,In_1297,In_1656);
nor U1023 (N_1023,In_999,In_2421);
nand U1024 (N_1024,In_1365,In_2437);
nor U1025 (N_1025,In_649,In_1552);
or U1026 (N_1026,In_532,In_2447);
nand U1027 (N_1027,In_1781,In_2003);
nor U1028 (N_1028,In_317,In_610);
and U1029 (N_1029,In_2226,In_685);
nand U1030 (N_1030,In_742,In_1162);
and U1031 (N_1031,In_1059,In_2462);
nor U1032 (N_1032,In_1262,In_2319);
or U1033 (N_1033,In_1395,In_1487);
nor U1034 (N_1034,In_2479,In_1034);
or U1035 (N_1035,In_1159,In_1834);
and U1036 (N_1036,In_658,In_1975);
and U1037 (N_1037,In_667,In_1682);
nor U1038 (N_1038,In_2155,In_813);
or U1039 (N_1039,In_1980,In_1081);
xnor U1040 (N_1040,In_1148,In_2495);
or U1041 (N_1041,In_1743,In_17);
or U1042 (N_1042,In_314,In_2097);
nor U1043 (N_1043,In_1318,In_735);
and U1044 (N_1044,In_1270,In_1375);
or U1045 (N_1045,In_2327,In_2013);
and U1046 (N_1046,In_873,In_1100);
or U1047 (N_1047,In_1795,In_2333);
or U1048 (N_1048,In_1629,In_2407);
or U1049 (N_1049,In_2384,In_724);
and U1050 (N_1050,In_1414,In_2101);
nor U1051 (N_1051,In_186,In_1494);
and U1052 (N_1052,In_2260,In_808);
and U1053 (N_1053,In_732,In_1393);
or U1054 (N_1054,In_1929,In_1863);
or U1055 (N_1055,In_2239,In_2483);
nor U1056 (N_1056,In_1097,In_803);
and U1057 (N_1057,In_590,In_1940);
or U1058 (N_1058,In_1175,In_1378);
or U1059 (N_1059,In_608,In_2037);
and U1060 (N_1060,In_1534,In_507);
nand U1061 (N_1061,In_1421,In_1372);
and U1062 (N_1062,In_313,In_581);
or U1063 (N_1063,In_1686,In_2157);
nand U1064 (N_1064,In_521,In_1278);
nand U1065 (N_1065,In_1398,In_1379);
or U1066 (N_1066,In_165,In_2093);
and U1067 (N_1067,In_30,In_1967);
nand U1068 (N_1068,In_248,In_1674);
and U1069 (N_1069,In_2065,In_583);
or U1070 (N_1070,In_1211,In_2098);
and U1071 (N_1071,In_2192,In_337);
and U1072 (N_1072,In_2212,In_214);
or U1073 (N_1073,In_812,In_1598);
xnor U1074 (N_1074,In_2386,In_166);
nor U1075 (N_1075,In_2329,In_869);
nor U1076 (N_1076,In_1759,In_201);
or U1077 (N_1077,In_209,In_1802);
and U1078 (N_1078,In_2064,In_2019);
nor U1079 (N_1079,In_141,In_734);
or U1080 (N_1080,In_1192,In_600);
nor U1081 (N_1081,In_2443,In_2304);
nand U1082 (N_1082,In_2313,In_2218);
or U1083 (N_1083,In_1208,In_1238);
nand U1084 (N_1084,In_556,In_2198);
and U1085 (N_1085,In_2071,In_1874);
nand U1086 (N_1086,In_569,In_1862);
nand U1087 (N_1087,In_266,In_980);
or U1088 (N_1088,In_604,In_1538);
nand U1089 (N_1089,In_2149,In_1088);
or U1090 (N_1090,In_1882,In_292);
nor U1091 (N_1091,In_2374,In_684);
and U1092 (N_1092,In_1737,In_383);
and U1093 (N_1093,In_623,In_2380);
nor U1094 (N_1094,In_1243,In_1785);
and U1095 (N_1095,In_1007,In_2036);
nand U1096 (N_1096,In_235,In_1637);
nand U1097 (N_1097,In_202,In_1115);
and U1098 (N_1098,In_1953,In_882);
and U1099 (N_1099,In_786,In_1069);
or U1100 (N_1100,In_94,In_2059);
or U1101 (N_1101,In_1268,In_2134);
or U1102 (N_1102,In_1409,In_2201);
nand U1103 (N_1103,In_2262,In_1928);
or U1104 (N_1104,In_1977,In_1247);
nand U1105 (N_1105,In_2052,In_63);
or U1106 (N_1106,In_872,In_358);
or U1107 (N_1107,In_1282,In_268);
and U1108 (N_1108,In_1661,In_1354);
and U1109 (N_1109,In_1963,In_991);
xor U1110 (N_1110,In_333,In_462);
and U1111 (N_1111,In_1074,In_1001);
nor U1112 (N_1112,In_1511,In_2335);
or U1113 (N_1113,In_1201,In_2259);
nand U1114 (N_1114,In_509,In_2294);
or U1115 (N_1115,In_1765,In_228);
nor U1116 (N_1116,In_376,In_621);
and U1117 (N_1117,In_2492,In_1658);
nor U1118 (N_1118,In_993,In_945);
nor U1119 (N_1119,In_1440,In_332);
or U1120 (N_1120,In_1194,In_622);
and U1121 (N_1121,In_2024,In_1438);
and U1122 (N_1122,In_970,In_1559);
or U1123 (N_1123,In_791,In_2058);
nor U1124 (N_1124,In_2406,In_765);
nand U1125 (N_1125,In_979,In_782);
and U1126 (N_1126,In_310,In_290);
and U1127 (N_1127,In_2412,In_1612);
nand U1128 (N_1128,In_1084,In_271);
and U1129 (N_1129,In_2403,In_2016);
nor U1130 (N_1130,In_691,In_1740);
nor U1131 (N_1131,In_2357,In_642);
xor U1132 (N_1132,In_651,In_884);
nor U1133 (N_1133,In_1800,In_429);
nor U1134 (N_1134,In_1263,In_587);
or U1135 (N_1135,In_680,In_1437);
nand U1136 (N_1136,In_1090,In_823);
nand U1137 (N_1137,In_1895,In_1913);
or U1138 (N_1138,In_1154,In_626);
nor U1139 (N_1139,In_9,In_1043);
nor U1140 (N_1140,In_1978,In_1817);
nor U1141 (N_1141,In_2089,In_682);
nor U1142 (N_1142,In_1575,In_2179);
nor U1143 (N_1143,In_240,In_414);
nor U1144 (N_1144,In_983,In_2031);
or U1145 (N_1145,In_1720,In_1918);
and U1146 (N_1146,In_1476,In_2383);
or U1147 (N_1147,In_2127,In_401);
and U1148 (N_1148,In_2145,In_1898);
and U1149 (N_1149,In_1927,In_1934);
or U1150 (N_1150,In_2244,In_1621);
xnor U1151 (N_1151,In_1615,In_1912);
xor U1152 (N_1152,In_160,In_239);
or U1153 (N_1153,In_436,In_1188);
and U1154 (N_1154,In_245,In_1752);
nand U1155 (N_1155,In_772,In_2222);
nor U1156 (N_1156,In_1384,In_1218);
nor U1157 (N_1157,In_2279,In_1954);
nand U1158 (N_1158,In_50,In_2414);
and U1159 (N_1159,In_2280,In_481);
nand U1160 (N_1160,In_1920,In_730);
and U1161 (N_1161,In_1850,In_1982);
nand U1162 (N_1162,In_1456,In_905);
nor U1163 (N_1163,In_1454,In_378);
and U1164 (N_1164,In_1364,In_2346);
nand U1165 (N_1165,In_232,In_1206);
and U1166 (N_1166,In_686,In_2050);
nand U1167 (N_1167,In_817,In_302);
or U1168 (N_1168,In_1535,In_379);
or U1169 (N_1169,In_996,In_2353);
or U1170 (N_1170,In_1467,In_1614);
nor U1171 (N_1171,In_1668,In_1907);
and U1172 (N_1172,In_2454,In_1500);
nor U1173 (N_1173,In_920,In_1868);
nor U1174 (N_1174,In_939,In_1418);
nor U1175 (N_1175,In_2200,In_1902);
or U1176 (N_1176,In_171,In_1140);
nand U1177 (N_1177,In_162,In_1590);
nor U1178 (N_1178,In_1519,In_1810);
nor U1179 (N_1179,In_99,In_529);
or U1180 (N_1180,In_1516,In_2457);
nor U1181 (N_1181,In_566,In_2009);
nor U1182 (N_1182,In_1905,In_1344);
xnor U1183 (N_1183,In_1845,In_1301);
and U1184 (N_1184,In_894,In_168);
nor U1185 (N_1185,In_1338,In_488);
nand U1186 (N_1186,In_2347,In_2204);
and U1187 (N_1187,In_2087,In_2154);
nand U1188 (N_1188,In_2422,In_1828);
or U1189 (N_1189,In_1986,In_185);
nor U1190 (N_1190,In_1144,In_1712);
and U1191 (N_1191,In_1719,In_2132);
or U1192 (N_1192,In_269,In_2046);
nand U1193 (N_1193,In_1166,In_210);
nor U1194 (N_1194,In_1382,In_1989);
or U1195 (N_1195,In_2343,In_55);
and U1196 (N_1196,In_2286,In_2284);
nand U1197 (N_1197,In_2185,In_491);
and U1198 (N_1198,In_1402,In_1961);
nor U1199 (N_1199,In_1623,In_1360);
nand U1200 (N_1200,In_1701,In_552);
and U1201 (N_1201,In_1116,In_213);
or U1202 (N_1202,In_1956,In_679);
nand U1203 (N_1203,In_1390,In_139);
nor U1204 (N_1204,In_1992,In_1664);
nand U1205 (N_1205,In_177,In_822);
nor U1206 (N_1206,In_947,In_1784);
and U1207 (N_1207,In_221,In_2493);
or U1208 (N_1208,In_661,In_1336);
nor U1209 (N_1209,In_190,In_2228);
nand U1210 (N_1210,In_1131,In_1677);
and U1211 (N_1211,In_2311,In_222);
nor U1212 (N_1212,In_1416,In_244);
nor U1213 (N_1213,In_1909,In_586);
or U1214 (N_1214,In_890,In_361);
and U1215 (N_1215,In_1065,In_1659);
or U1216 (N_1216,In_2018,In_384);
nor U1217 (N_1217,In_87,In_306);
and U1218 (N_1218,In_1998,In_1161);
nor U1219 (N_1219,In_1841,In_1754);
nand U1220 (N_1220,In_540,In_1803);
or U1221 (N_1221,In_958,In_1189);
or U1222 (N_1222,In_1213,In_1748);
and U1223 (N_1223,In_34,In_860);
nor U1224 (N_1224,In_2219,In_789);
and U1225 (N_1225,In_2182,In_1446);
and U1226 (N_1226,In_2436,In_161);
or U1227 (N_1227,In_1434,In_670);
nor U1228 (N_1228,In_1313,In_712);
xnor U1229 (N_1229,In_2356,In_77);
and U1230 (N_1230,In_2489,In_538);
or U1231 (N_1231,In_2463,In_1163);
nor U1232 (N_1232,In_44,In_2102);
or U1233 (N_1233,In_1758,In_1649);
nand U1234 (N_1234,In_2297,In_693);
and U1235 (N_1235,In_1125,In_1184);
or U1236 (N_1236,In_1371,In_1020);
nor U1237 (N_1237,In_1311,In_1223);
nor U1238 (N_1238,In_1468,In_296);
nor U1239 (N_1239,In_597,In_1145);
xor U1240 (N_1240,In_2040,In_330);
nand U1241 (N_1241,In_756,In_816);
nor U1242 (N_1242,In_20,In_331);
nor U1243 (N_1243,In_2167,In_1824);
and U1244 (N_1244,In_1657,In_1513);
or U1245 (N_1245,In_1106,In_657);
and U1246 (N_1246,In_1990,In_155);
and U1247 (N_1247,In_1016,In_359);
xnor U1248 (N_1248,In_2224,In_227);
or U1249 (N_1249,In_2363,In_1176);
nor U1250 (N_1250,In_2114,In_194);
and U1251 (N_1251,In_971,In_1921);
or U1252 (N_1252,In_2104,In_1396);
and U1253 (N_1253,In_1028,In_1382);
and U1254 (N_1254,In_1989,In_11);
nand U1255 (N_1255,In_2286,In_810);
and U1256 (N_1256,In_1414,In_1264);
and U1257 (N_1257,In_1839,In_432);
nor U1258 (N_1258,In_1794,In_1009);
and U1259 (N_1259,In_1733,In_1585);
nor U1260 (N_1260,In_1892,In_837);
nand U1261 (N_1261,In_505,In_724);
nor U1262 (N_1262,In_260,In_1931);
or U1263 (N_1263,In_692,In_2361);
nor U1264 (N_1264,In_22,In_1253);
nor U1265 (N_1265,In_2433,In_1068);
nor U1266 (N_1266,In_1470,In_1055);
nor U1267 (N_1267,In_1688,In_629);
and U1268 (N_1268,In_584,In_1692);
nor U1269 (N_1269,In_2271,In_1427);
or U1270 (N_1270,In_884,In_1587);
or U1271 (N_1271,In_387,In_1735);
nand U1272 (N_1272,In_335,In_1130);
and U1273 (N_1273,In_1531,In_592);
nor U1274 (N_1274,In_1504,In_227);
and U1275 (N_1275,In_396,In_2286);
nand U1276 (N_1276,In_58,In_996);
nand U1277 (N_1277,In_2224,In_1126);
and U1278 (N_1278,In_1061,In_1352);
and U1279 (N_1279,In_1385,In_138);
nand U1280 (N_1280,In_102,In_990);
and U1281 (N_1281,In_598,In_706);
and U1282 (N_1282,In_425,In_1856);
nand U1283 (N_1283,In_48,In_388);
nand U1284 (N_1284,In_2339,In_481);
nor U1285 (N_1285,In_1773,In_2421);
nor U1286 (N_1286,In_1542,In_1951);
and U1287 (N_1287,In_1151,In_1202);
and U1288 (N_1288,In_1405,In_1888);
and U1289 (N_1289,In_1403,In_1888);
or U1290 (N_1290,In_1606,In_222);
nand U1291 (N_1291,In_2082,In_811);
nor U1292 (N_1292,In_1079,In_2209);
nor U1293 (N_1293,In_2356,In_2086);
and U1294 (N_1294,In_2441,In_1922);
nor U1295 (N_1295,In_249,In_518);
nand U1296 (N_1296,In_703,In_1658);
nand U1297 (N_1297,In_1456,In_231);
nand U1298 (N_1298,In_298,In_225);
and U1299 (N_1299,In_2075,In_810);
and U1300 (N_1300,In_166,In_2329);
nor U1301 (N_1301,In_851,In_1596);
and U1302 (N_1302,In_2175,In_267);
nor U1303 (N_1303,In_1905,In_2106);
nand U1304 (N_1304,In_167,In_2248);
nand U1305 (N_1305,In_582,In_1742);
and U1306 (N_1306,In_1185,In_2037);
xor U1307 (N_1307,In_1631,In_660);
and U1308 (N_1308,In_250,In_1459);
nand U1309 (N_1309,In_257,In_14);
nand U1310 (N_1310,In_247,In_2227);
nor U1311 (N_1311,In_173,In_791);
nand U1312 (N_1312,In_2418,In_1415);
xnor U1313 (N_1313,In_1575,In_2428);
or U1314 (N_1314,In_1177,In_2018);
nor U1315 (N_1315,In_2378,In_2030);
xor U1316 (N_1316,In_541,In_1153);
or U1317 (N_1317,In_1980,In_2399);
or U1318 (N_1318,In_1480,In_2079);
xor U1319 (N_1319,In_230,In_1145);
or U1320 (N_1320,In_234,In_2164);
nor U1321 (N_1321,In_1708,In_1416);
nand U1322 (N_1322,In_901,In_998);
nor U1323 (N_1323,In_2076,In_95);
and U1324 (N_1324,In_1680,In_264);
or U1325 (N_1325,In_514,In_1260);
and U1326 (N_1326,In_2062,In_877);
or U1327 (N_1327,In_1489,In_1185);
or U1328 (N_1328,In_2169,In_861);
and U1329 (N_1329,In_1579,In_1043);
nand U1330 (N_1330,In_2240,In_1169);
nand U1331 (N_1331,In_9,In_184);
nor U1332 (N_1332,In_1983,In_1266);
nor U1333 (N_1333,In_889,In_1677);
or U1334 (N_1334,In_283,In_281);
nand U1335 (N_1335,In_435,In_2306);
and U1336 (N_1336,In_20,In_1812);
nor U1337 (N_1337,In_2405,In_1831);
nor U1338 (N_1338,In_2329,In_1238);
nand U1339 (N_1339,In_1133,In_720);
and U1340 (N_1340,In_27,In_1882);
or U1341 (N_1341,In_2196,In_1015);
nor U1342 (N_1342,In_759,In_478);
nor U1343 (N_1343,In_1834,In_1870);
or U1344 (N_1344,In_1327,In_689);
and U1345 (N_1345,In_1666,In_1890);
nor U1346 (N_1346,In_809,In_1485);
or U1347 (N_1347,In_1639,In_1215);
nand U1348 (N_1348,In_2054,In_2108);
nor U1349 (N_1349,In_561,In_2262);
xnor U1350 (N_1350,In_1047,In_1821);
nand U1351 (N_1351,In_1521,In_2143);
nor U1352 (N_1352,In_2464,In_1582);
nor U1353 (N_1353,In_705,In_833);
or U1354 (N_1354,In_274,In_342);
nor U1355 (N_1355,In_1473,In_726);
nand U1356 (N_1356,In_1149,In_1201);
nor U1357 (N_1357,In_72,In_806);
nand U1358 (N_1358,In_1619,In_1755);
nor U1359 (N_1359,In_1347,In_1198);
nor U1360 (N_1360,In_2241,In_1176);
or U1361 (N_1361,In_1372,In_2008);
nor U1362 (N_1362,In_478,In_1426);
nand U1363 (N_1363,In_1469,In_1345);
nand U1364 (N_1364,In_2004,In_2297);
or U1365 (N_1365,In_804,In_1147);
or U1366 (N_1366,In_2119,In_2009);
or U1367 (N_1367,In_2160,In_943);
or U1368 (N_1368,In_1637,In_2377);
and U1369 (N_1369,In_1402,In_2487);
nand U1370 (N_1370,In_937,In_2069);
or U1371 (N_1371,In_10,In_865);
nand U1372 (N_1372,In_1055,In_444);
nor U1373 (N_1373,In_495,In_207);
and U1374 (N_1374,In_1421,In_451);
nand U1375 (N_1375,In_834,In_1147);
nor U1376 (N_1376,In_611,In_2123);
nand U1377 (N_1377,In_460,In_411);
nor U1378 (N_1378,In_2366,In_1401);
nor U1379 (N_1379,In_2155,In_1989);
and U1380 (N_1380,In_275,In_125);
nand U1381 (N_1381,In_454,In_2107);
or U1382 (N_1382,In_435,In_916);
or U1383 (N_1383,In_788,In_1190);
nor U1384 (N_1384,In_2277,In_569);
and U1385 (N_1385,In_1279,In_467);
and U1386 (N_1386,In_2177,In_2000);
nor U1387 (N_1387,In_1972,In_2308);
nand U1388 (N_1388,In_1045,In_1318);
and U1389 (N_1389,In_620,In_2423);
nor U1390 (N_1390,In_1948,In_214);
nand U1391 (N_1391,In_1368,In_290);
or U1392 (N_1392,In_548,In_47);
or U1393 (N_1393,In_649,In_2411);
or U1394 (N_1394,In_51,In_1896);
nor U1395 (N_1395,In_1730,In_860);
nor U1396 (N_1396,In_1465,In_353);
and U1397 (N_1397,In_1184,In_176);
and U1398 (N_1398,In_1713,In_47);
and U1399 (N_1399,In_381,In_972);
and U1400 (N_1400,In_1696,In_1046);
nor U1401 (N_1401,In_1827,In_361);
nand U1402 (N_1402,In_189,In_746);
or U1403 (N_1403,In_1163,In_854);
nand U1404 (N_1404,In_1649,In_2427);
and U1405 (N_1405,In_854,In_1957);
nand U1406 (N_1406,In_979,In_2356);
and U1407 (N_1407,In_1740,In_137);
nor U1408 (N_1408,In_1129,In_2079);
nor U1409 (N_1409,In_117,In_1817);
and U1410 (N_1410,In_1418,In_946);
or U1411 (N_1411,In_802,In_1298);
and U1412 (N_1412,In_240,In_1427);
nor U1413 (N_1413,In_2235,In_401);
nor U1414 (N_1414,In_57,In_2163);
or U1415 (N_1415,In_1905,In_754);
and U1416 (N_1416,In_1132,In_1999);
nand U1417 (N_1417,In_126,In_619);
nand U1418 (N_1418,In_2035,In_1470);
and U1419 (N_1419,In_191,In_1983);
nor U1420 (N_1420,In_845,In_2443);
or U1421 (N_1421,In_1441,In_1467);
or U1422 (N_1422,In_2079,In_2235);
nand U1423 (N_1423,In_1817,In_860);
nor U1424 (N_1424,In_665,In_1750);
nand U1425 (N_1425,In_1813,In_16);
or U1426 (N_1426,In_2114,In_2254);
nand U1427 (N_1427,In_1228,In_95);
or U1428 (N_1428,In_1107,In_1200);
xor U1429 (N_1429,In_895,In_687);
and U1430 (N_1430,In_2448,In_443);
nand U1431 (N_1431,In_811,In_1186);
and U1432 (N_1432,In_955,In_1738);
and U1433 (N_1433,In_485,In_632);
nor U1434 (N_1434,In_1217,In_1893);
and U1435 (N_1435,In_836,In_1322);
nor U1436 (N_1436,In_72,In_580);
and U1437 (N_1437,In_1766,In_217);
or U1438 (N_1438,In_204,In_2208);
nand U1439 (N_1439,In_1371,In_1599);
and U1440 (N_1440,In_130,In_537);
and U1441 (N_1441,In_1656,In_1533);
nand U1442 (N_1442,In_2227,In_441);
or U1443 (N_1443,In_580,In_729);
and U1444 (N_1444,In_558,In_1328);
nor U1445 (N_1445,In_299,In_1681);
and U1446 (N_1446,In_2294,In_272);
nand U1447 (N_1447,In_257,In_560);
and U1448 (N_1448,In_1504,In_2174);
nor U1449 (N_1449,In_1188,In_426);
or U1450 (N_1450,In_1544,In_1667);
and U1451 (N_1451,In_777,In_632);
and U1452 (N_1452,In_745,In_2387);
and U1453 (N_1453,In_1666,In_2468);
nand U1454 (N_1454,In_236,In_1567);
nor U1455 (N_1455,In_1990,In_737);
nor U1456 (N_1456,In_2257,In_560);
nor U1457 (N_1457,In_54,In_2088);
nand U1458 (N_1458,In_1141,In_2264);
or U1459 (N_1459,In_1884,In_99);
or U1460 (N_1460,In_1823,In_970);
or U1461 (N_1461,In_1248,In_798);
nand U1462 (N_1462,In_2171,In_1516);
nor U1463 (N_1463,In_1980,In_1966);
nand U1464 (N_1464,In_2131,In_1421);
or U1465 (N_1465,In_332,In_772);
or U1466 (N_1466,In_1519,In_1382);
and U1467 (N_1467,In_352,In_874);
nand U1468 (N_1468,In_108,In_505);
nand U1469 (N_1469,In_429,In_1555);
nor U1470 (N_1470,In_1682,In_873);
and U1471 (N_1471,In_522,In_669);
nor U1472 (N_1472,In_889,In_806);
or U1473 (N_1473,In_1485,In_2201);
nor U1474 (N_1474,In_1496,In_731);
and U1475 (N_1475,In_1208,In_201);
nor U1476 (N_1476,In_572,In_2276);
nor U1477 (N_1477,In_2315,In_1252);
nor U1478 (N_1478,In_2287,In_514);
nor U1479 (N_1479,In_1905,In_2343);
and U1480 (N_1480,In_860,In_436);
nor U1481 (N_1481,In_44,In_490);
and U1482 (N_1482,In_2135,In_260);
and U1483 (N_1483,In_1326,In_1217);
nor U1484 (N_1484,In_20,In_779);
and U1485 (N_1485,In_1251,In_1049);
nand U1486 (N_1486,In_1349,In_405);
and U1487 (N_1487,In_1332,In_451);
and U1488 (N_1488,In_846,In_2014);
or U1489 (N_1489,In_2094,In_305);
nand U1490 (N_1490,In_1251,In_650);
nor U1491 (N_1491,In_2349,In_1659);
or U1492 (N_1492,In_196,In_517);
xnor U1493 (N_1493,In_1292,In_1671);
nor U1494 (N_1494,In_1694,In_1421);
nor U1495 (N_1495,In_1311,In_312);
or U1496 (N_1496,In_1510,In_2334);
nor U1497 (N_1497,In_2410,In_460);
or U1498 (N_1498,In_2442,In_722);
nand U1499 (N_1499,In_244,In_1850);
nor U1500 (N_1500,In_807,In_2479);
xnor U1501 (N_1501,In_865,In_453);
or U1502 (N_1502,In_1573,In_346);
or U1503 (N_1503,In_2281,In_328);
and U1504 (N_1504,In_1764,In_528);
or U1505 (N_1505,In_1943,In_2092);
or U1506 (N_1506,In_1651,In_2437);
or U1507 (N_1507,In_1558,In_2301);
or U1508 (N_1508,In_808,In_1029);
nor U1509 (N_1509,In_274,In_1323);
or U1510 (N_1510,In_2469,In_2005);
nand U1511 (N_1511,In_1806,In_682);
nor U1512 (N_1512,In_534,In_2174);
nand U1513 (N_1513,In_785,In_662);
or U1514 (N_1514,In_194,In_1451);
and U1515 (N_1515,In_52,In_2144);
nand U1516 (N_1516,In_280,In_1716);
nand U1517 (N_1517,In_1286,In_1399);
and U1518 (N_1518,In_157,In_1549);
and U1519 (N_1519,In_1711,In_186);
or U1520 (N_1520,In_651,In_1692);
or U1521 (N_1521,In_835,In_2046);
nor U1522 (N_1522,In_1845,In_2073);
or U1523 (N_1523,In_1919,In_1229);
or U1524 (N_1524,In_2336,In_571);
nor U1525 (N_1525,In_399,In_2276);
nor U1526 (N_1526,In_2148,In_1106);
or U1527 (N_1527,In_1867,In_47);
nand U1528 (N_1528,In_1434,In_2315);
nand U1529 (N_1529,In_1638,In_2140);
nor U1530 (N_1530,In_1931,In_1874);
nor U1531 (N_1531,In_1686,In_400);
or U1532 (N_1532,In_1837,In_1197);
and U1533 (N_1533,In_2276,In_1516);
or U1534 (N_1534,In_1143,In_1222);
or U1535 (N_1535,In_796,In_1638);
nand U1536 (N_1536,In_2068,In_436);
nand U1537 (N_1537,In_1233,In_366);
or U1538 (N_1538,In_1795,In_847);
and U1539 (N_1539,In_46,In_940);
nand U1540 (N_1540,In_861,In_1016);
nand U1541 (N_1541,In_774,In_518);
and U1542 (N_1542,In_730,In_1630);
nand U1543 (N_1543,In_1962,In_1098);
or U1544 (N_1544,In_206,In_598);
and U1545 (N_1545,In_2362,In_130);
or U1546 (N_1546,In_1797,In_727);
nor U1547 (N_1547,In_2484,In_1818);
and U1548 (N_1548,In_964,In_1142);
and U1549 (N_1549,In_200,In_9);
nor U1550 (N_1550,In_552,In_1198);
and U1551 (N_1551,In_682,In_1748);
or U1552 (N_1552,In_1411,In_764);
or U1553 (N_1553,In_1405,In_219);
nand U1554 (N_1554,In_1256,In_2422);
and U1555 (N_1555,In_2405,In_853);
or U1556 (N_1556,In_221,In_1080);
and U1557 (N_1557,In_1775,In_407);
nand U1558 (N_1558,In_1027,In_2454);
or U1559 (N_1559,In_211,In_565);
or U1560 (N_1560,In_2210,In_1944);
and U1561 (N_1561,In_1198,In_2386);
and U1562 (N_1562,In_885,In_289);
nand U1563 (N_1563,In_1052,In_1220);
xor U1564 (N_1564,In_1100,In_445);
and U1565 (N_1565,In_2425,In_628);
nand U1566 (N_1566,In_1526,In_2132);
or U1567 (N_1567,In_1278,In_558);
nand U1568 (N_1568,In_2088,In_1975);
nor U1569 (N_1569,In_2257,In_1936);
nor U1570 (N_1570,In_677,In_1733);
nand U1571 (N_1571,In_2161,In_1785);
xnor U1572 (N_1572,In_84,In_813);
nor U1573 (N_1573,In_548,In_1036);
or U1574 (N_1574,In_1873,In_1856);
or U1575 (N_1575,In_631,In_2217);
nor U1576 (N_1576,In_2018,In_2285);
or U1577 (N_1577,In_1544,In_2417);
nand U1578 (N_1578,In_1869,In_2432);
nand U1579 (N_1579,In_1860,In_1456);
and U1580 (N_1580,In_179,In_1391);
and U1581 (N_1581,In_263,In_2014);
nand U1582 (N_1582,In_4,In_787);
and U1583 (N_1583,In_414,In_1339);
or U1584 (N_1584,In_753,In_347);
and U1585 (N_1585,In_2328,In_269);
nand U1586 (N_1586,In_2139,In_1342);
or U1587 (N_1587,In_928,In_2432);
nand U1588 (N_1588,In_1076,In_1099);
or U1589 (N_1589,In_42,In_1358);
and U1590 (N_1590,In_2489,In_1980);
or U1591 (N_1591,In_2069,In_2351);
and U1592 (N_1592,In_226,In_1266);
nor U1593 (N_1593,In_1533,In_62);
nor U1594 (N_1594,In_1685,In_476);
or U1595 (N_1595,In_1925,In_2486);
nor U1596 (N_1596,In_1182,In_1777);
nand U1597 (N_1597,In_207,In_1896);
or U1598 (N_1598,In_111,In_840);
nand U1599 (N_1599,In_641,In_2151);
nor U1600 (N_1600,In_59,In_1280);
nand U1601 (N_1601,In_692,In_1733);
and U1602 (N_1602,In_2344,In_1314);
or U1603 (N_1603,In_1193,In_321);
nand U1604 (N_1604,In_81,In_946);
nor U1605 (N_1605,In_776,In_1766);
nand U1606 (N_1606,In_33,In_1646);
or U1607 (N_1607,In_2436,In_1677);
nand U1608 (N_1608,In_1977,In_1618);
nor U1609 (N_1609,In_2320,In_6);
and U1610 (N_1610,In_723,In_1204);
and U1611 (N_1611,In_562,In_2390);
nand U1612 (N_1612,In_716,In_789);
nor U1613 (N_1613,In_2492,In_586);
or U1614 (N_1614,In_1774,In_2305);
nand U1615 (N_1615,In_332,In_2170);
nor U1616 (N_1616,In_1468,In_777);
and U1617 (N_1617,In_1213,In_1526);
and U1618 (N_1618,In_1194,In_2493);
nor U1619 (N_1619,In_1433,In_984);
nand U1620 (N_1620,In_1337,In_34);
and U1621 (N_1621,In_697,In_1976);
nand U1622 (N_1622,In_408,In_2205);
and U1623 (N_1623,In_2168,In_847);
nand U1624 (N_1624,In_2004,In_2415);
and U1625 (N_1625,In_1066,In_1599);
nand U1626 (N_1626,In_1919,In_180);
nand U1627 (N_1627,In_714,In_559);
or U1628 (N_1628,In_479,In_1061);
nor U1629 (N_1629,In_487,In_1540);
and U1630 (N_1630,In_1112,In_1973);
nand U1631 (N_1631,In_988,In_1225);
nand U1632 (N_1632,In_1844,In_2017);
or U1633 (N_1633,In_2091,In_270);
or U1634 (N_1634,In_1371,In_672);
or U1635 (N_1635,In_814,In_15);
and U1636 (N_1636,In_305,In_322);
or U1637 (N_1637,In_1157,In_1465);
nand U1638 (N_1638,In_810,In_2393);
nand U1639 (N_1639,In_1013,In_1635);
or U1640 (N_1640,In_311,In_1272);
or U1641 (N_1641,In_1040,In_1509);
and U1642 (N_1642,In_199,In_1332);
nor U1643 (N_1643,In_2259,In_1789);
nand U1644 (N_1644,In_1122,In_1317);
nor U1645 (N_1645,In_1858,In_1519);
and U1646 (N_1646,In_597,In_2226);
nor U1647 (N_1647,In_2372,In_1209);
and U1648 (N_1648,In_2131,In_1633);
nand U1649 (N_1649,In_1287,In_137);
xor U1650 (N_1650,In_2017,In_926);
nand U1651 (N_1651,In_1793,In_2101);
nor U1652 (N_1652,In_2161,In_887);
nor U1653 (N_1653,In_1837,In_845);
or U1654 (N_1654,In_881,In_770);
nor U1655 (N_1655,In_732,In_957);
nor U1656 (N_1656,In_1334,In_408);
or U1657 (N_1657,In_1483,In_1129);
xnor U1658 (N_1658,In_687,In_1629);
nor U1659 (N_1659,In_2337,In_725);
nand U1660 (N_1660,In_2137,In_357);
and U1661 (N_1661,In_1470,In_319);
nor U1662 (N_1662,In_1289,In_77);
nor U1663 (N_1663,In_1963,In_1296);
nor U1664 (N_1664,In_1224,In_1249);
xor U1665 (N_1665,In_920,In_257);
nor U1666 (N_1666,In_522,In_1065);
and U1667 (N_1667,In_1920,In_590);
and U1668 (N_1668,In_2141,In_2294);
and U1669 (N_1669,In_871,In_696);
nor U1670 (N_1670,In_288,In_2376);
nand U1671 (N_1671,In_952,In_1386);
nor U1672 (N_1672,In_1481,In_2272);
nor U1673 (N_1673,In_1673,In_223);
nand U1674 (N_1674,In_2414,In_1997);
nand U1675 (N_1675,In_1028,In_214);
nor U1676 (N_1676,In_1164,In_154);
and U1677 (N_1677,In_2200,In_853);
nor U1678 (N_1678,In_727,In_374);
nand U1679 (N_1679,In_1872,In_1098);
nand U1680 (N_1680,In_704,In_572);
nor U1681 (N_1681,In_1387,In_1692);
xnor U1682 (N_1682,In_1097,In_1282);
nand U1683 (N_1683,In_2004,In_231);
xnor U1684 (N_1684,In_1578,In_393);
nand U1685 (N_1685,In_220,In_586);
and U1686 (N_1686,In_1360,In_1546);
nand U1687 (N_1687,In_1676,In_704);
nand U1688 (N_1688,In_10,In_1834);
nor U1689 (N_1689,In_146,In_1947);
or U1690 (N_1690,In_1742,In_568);
and U1691 (N_1691,In_837,In_702);
and U1692 (N_1692,In_1031,In_2318);
and U1693 (N_1693,In_917,In_1448);
and U1694 (N_1694,In_2127,In_2070);
or U1695 (N_1695,In_81,In_2278);
and U1696 (N_1696,In_776,In_563);
nand U1697 (N_1697,In_157,In_1032);
nand U1698 (N_1698,In_1512,In_734);
nand U1699 (N_1699,In_1652,In_1545);
or U1700 (N_1700,In_2126,In_472);
nor U1701 (N_1701,In_2456,In_46);
and U1702 (N_1702,In_1109,In_1062);
and U1703 (N_1703,In_1257,In_1934);
or U1704 (N_1704,In_250,In_2067);
and U1705 (N_1705,In_1844,In_1354);
or U1706 (N_1706,In_966,In_338);
nand U1707 (N_1707,In_391,In_326);
nand U1708 (N_1708,In_337,In_1711);
nor U1709 (N_1709,In_559,In_228);
and U1710 (N_1710,In_2365,In_945);
xnor U1711 (N_1711,In_738,In_341);
nand U1712 (N_1712,In_153,In_808);
nand U1713 (N_1713,In_1745,In_1125);
nor U1714 (N_1714,In_2127,In_1757);
nor U1715 (N_1715,In_1986,In_123);
nor U1716 (N_1716,In_520,In_1171);
nand U1717 (N_1717,In_1694,In_1494);
or U1718 (N_1718,In_62,In_51);
and U1719 (N_1719,In_641,In_721);
and U1720 (N_1720,In_2396,In_2470);
or U1721 (N_1721,In_1266,In_1198);
or U1722 (N_1722,In_367,In_167);
nor U1723 (N_1723,In_331,In_1135);
nor U1724 (N_1724,In_1679,In_501);
nor U1725 (N_1725,In_2176,In_703);
and U1726 (N_1726,In_2461,In_1392);
nor U1727 (N_1727,In_2036,In_1317);
nand U1728 (N_1728,In_736,In_1847);
and U1729 (N_1729,In_269,In_28);
and U1730 (N_1730,In_424,In_918);
nand U1731 (N_1731,In_2350,In_1918);
nor U1732 (N_1732,In_1534,In_721);
xor U1733 (N_1733,In_2203,In_1146);
nand U1734 (N_1734,In_996,In_2084);
nor U1735 (N_1735,In_1154,In_1590);
and U1736 (N_1736,In_2469,In_1124);
and U1737 (N_1737,In_1185,In_1625);
nor U1738 (N_1738,In_2151,In_788);
nor U1739 (N_1739,In_782,In_1231);
or U1740 (N_1740,In_1196,In_2379);
nor U1741 (N_1741,In_1320,In_2387);
and U1742 (N_1742,In_1653,In_960);
nand U1743 (N_1743,In_2006,In_2265);
nand U1744 (N_1744,In_2237,In_925);
nand U1745 (N_1745,In_653,In_404);
or U1746 (N_1746,In_2381,In_913);
nand U1747 (N_1747,In_1722,In_1794);
nand U1748 (N_1748,In_1251,In_2335);
nand U1749 (N_1749,In_2330,In_385);
and U1750 (N_1750,In_726,In_1328);
and U1751 (N_1751,In_994,In_915);
nand U1752 (N_1752,In_1320,In_1600);
nand U1753 (N_1753,In_2487,In_320);
nor U1754 (N_1754,In_141,In_589);
nand U1755 (N_1755,In_2488,In_2136);
nor U1756 (N_1756,In_2217,In_598);
nand U1757 (N_1757,In_423,In_2127);
or U1758 (N_1758,In_269,In_1420);
and U1759 (N_1759,In_1655,In_803);
and U1760 (N_1760,In_867,In_2075);
and U1761 (N_1761,In_912,In_1119);
nor U1762 (N_1762,In_2463,In_875);
or U1763 (N_1763,In_787,In_95);
nor U1764 (N_1764,In_1079,In_2256);
nor U1765 (N_1765,In_467,In_1115);
nand U1766 (N_1766,In_200,In_2281);
and U1767 (N_1767,In_1493,In_1508);
nor U1768 (N_1768,In_825,In_2047);
or U1769 (N_1769,In_16,In_2043);
nor U1770 (N_1770,In_61,In_482);
nor U1771 (N_1771,In_1361,In_1962);
and U1772 (N_1772,In_2240,In_2060);
nor U1773 (N_1773,In_1663,In_141);
nand U1774 (N_1774,In_2234,In_1800);
or U1775 (N_1775,In_1677,In_2086);
nand U1776 (N_1776,In_438,In_1015);
nand U1777 (N_1777,In_2320,In_719);
xor U1778 (N_1778,In_441,In_894);
or U1779 (N_1779,In_2434,In_328);
and U1780 (N_1780,In_2358,In_2329);
and U1781 (N_1781,In_1433,In_312);
and U1782 (N_1782,In_1558,In_2267);
and U1783 (N_1783,In_1693,In_558);
and U1784 (N_1784,In_1923,In_1996);
and U1785 (N_1785,In_644,In_37);
nor U1786 (N_1786,In_1156,In_2401);
or U1787 (N_1787,In_455,In_1957);
and U1788 (N_1788,In_57,In_994);
nand U1789 (N_1789,In_772,In_1749);
nor U1790 (N_1790,In_450,In_1657);
or U1791 (N_1791,In_1972,In_1069);
nor U1792 (N_1792,In_200,In_493);
nor U1793 (N_1793,In_1499,In_304);
nor U1794 (N_1794,In_797,In_1862);
nor U1795 (N_1795,In_1337,In_360);
nand U1796 (N_1796,In_1663,In_1671);
or U1797 (N_1797,In_39,In_1734);
or U1798 (N_1798,In_1655,In_1648);
nand U1799 (N_1799,In_1090,In_2190);
nand U1800 (N_1800,In_1121,In_1569);
or U1801 (N_1801,In_1794,In_1407);
nand U1802 (N_1802,In_1702,In_2095);
and U1803 (N_1803,In_1808,In_881);
nor U1804 (N_1804,In_1275,In_427);
and U1805 (N_1805,In_155,In_2010);
nand U1806 (N_1806,In_1906,In_900);
nor U1807 (N_1807,In_1187,In_586);
nand U1808 (N_1808,In_762,In_348);
or U1809 (N_1809,In_1699,In_1922);
or U1810 (N_1810,In_174,In_2212);
nand U1811 (N_1811,In_85,In_2255);
nand U1812 (N_1812,In_1985,In_1478);
nand U1813 (N_1813,In_2450,In_546);
nor U1814 (N_1814,In_850,In_1901);
and U1815 (N_1815,In_1572,In_846);
nand U1816 (N_1816,In_2459,In_756);
nor U1817 (N_1817,In_720,In_519);
and U1818 (N_1818,In_939,In_1980);
nor U1819 (N_1819,In_725,In_517);
nand U1820 (N_1820,In_418,In_26);
nor U1821 (N_1821,In_1875,In_1246);
nand U1822 (N_1822,In_720,In_453);
nor U1823 (N_1823,In_1908,In_323);
nand U1824 (N_1824,In_681,In_801);
nor U1825 (N_1825,In_2020,In_1032);
nor U1826 (N_1826,In_2210,In_705);
nor U1827 (N_1827,In_1134,In_1427);
xor U1828 (N_1828,In_1007,In_319);
nand U1829 (N_1829,In_680,In_1742);
or U1830 (N_1830,In_2295,In_1807);
xnor U1831 (N_1831,In_1842,In_1566);
or U1832 (N_1832,In_2230,In_352);
nand U1833 (N_1833,In_927,In_1801);
or U1834 (N_1834,In_1195,In_1109);
nor U1835 (N_1835,In_866,In_1096);
nor U1836 (N_1836,In_1283,In_879);
and U1837 (N_1837,In_1163,In_1505);
nor U1838 (N_1838,In_505,In_755);
or U1839 (N_1839,In_1508,In_2465);
and U1840 (N_1840,In_1636,In_390);
and U1841 (N_1841,In_0,In_62);
nand U1842 (N_1842,In_906,In_1209);
xor U1843 (N_1843,In_2309,In_2248);
nand U1844 (N_1844,In_1011,In_1560);
or U1845 (N_1845,In_519,In_2288);
nand U1846 (N_1846,In_268,In_2408);
or U1847 (N_1847,In_1938,In_2118);
nand U1848 (N_1848,In_1480,In_1451);
nor U1849 (N_1849,In_683,In_2106);
or U1850 (N_1850,In_1562,In_958);
and U1851 (N_1851,In_436,In_1421);
xor U1852 (N_1852,In_2251,In_1929);
and U1853 (N_1853,In_2400,In_578);
nor U1854 (N_1854,In_1183,In_958);
or U1855 (N_1855,In_1008,In_233);
nor U1856 (N_1856,In_648,In_68);
and U1857 (N_1857,In_1381,In_128);
and U1858 (N_1858,In_414,In_356);
nor U1859 (N_1859,In_1338,In_186);
and U1860 (N_1860,In_735,In_2031);
nor U1861 (N_1861,In_1606,In_577);
or U1862 (N_1862,In_685,In_415);
or U1863 (N_1863,In_2478,In_1039);
nor U1864 (N_1864,In_1454,In_1946);
or U1865 (N_1865,In_1613,In_252);
nand U1866 (N_1866,In_1514,In_1334);
and U1867 (N_1867,In_611,In_1349);
nor U1868 (N_1868,In_1573,In_1109);
nand U1869 (N_1869,In_1743,In_1600);
nor U1870 (N_1870,In_120,In_325);
nor U1871 (N_1871,In_2099,In_2213);
nor U1872 (N_1872,In_409,In_163);
nor U1873 (N_1873,In_792,In_1814);
nor U1874 (N_1874,In_503,In_1390);
xnor U1875 (N_1875,In_1476,In_479);
nand U1876 (N_1876,In_1261,In_1343);
nor U1877 (N_1877,In_1053,In_774);
nor U1878 (N_1878,In_539,In_1771);
nor U1879 (N_1879,In_1422,In_1504);
nor U1880 (N_1880,In_2200,In_1526);
and U1881 (N_1881,In_985,In_1878);
nand U1882 (N_1882,In_1213,In_871);
nand U1883 (N_1883,In_909,In_2258);
nand U1884 (N_1884,In_1704,In_1667);
nand U1885 (N_1885,In_1618,In_509);
nand U1886 (N_1886,In_2479,In_237);
or U1887 (N_1887,In_566,In_2203);
and U1888 (N_1888,In_2469,In_1241);
nand U1889 (N_1889,In_1365,In_666);
nor U1890 (N_1890,In_1669,In_341);
nand U1891 (N_1891,In_1669,In_1774);
or U1892 (N_1892,In_1113,In_434);
or U1893 (N_1893,In_876,In_1808);
and U1894 (N_1894,In_653,In_1869);
nor U1895 (N_1895,In_1119,In_1582);
nand U1896 (N_1896,In_2167,In_1105);
and U1897 (N_1897,In_427,In_84);
nor U1898 (N_1898,In_2369,In_990);
nor U1899 (N_1899,In_165,In_5);
nand U1900 (N_1900,In_2200,In_1028);
nor U1901 (N_1901,In_602,In_729);
nand U1902 (N_1902,In_395,In_73);
nor U1903 (N_1903,In_1127,In_310);
or U1904 (N_1904,In_1728,In_1852);
nor U1905 (N_1905,In_1009,In_572);
or U1906 (N_1906,In_1813,In_1794);
nand U1907 (N_1907,In_260,In_661);
nand U1908 (N_1908,In_552,In_885);
or U1909 (N_1909,In_132,In_1083);
and U1910 (N_1910,In_1018,In_1209);
nor U1911 (N_1911,In_164,In_397);
nand U1912 (N_1912,In_497,In_1598);
nand U1913 (N_1913,In_1529,In_798);
and U1914 (N_1914,In_263,In_1047);
and U1915 (N_1915,In_1216,In_222);
xnor U1916 (N_1916,In_1225,In_1487);
nand U1917 (N_1917,In_850,In_2208);
nor U1918 (N_1918,In_968,In_1848);
nand U1919 (N_1919,In_119,In_2297);
nand U1920 (N_1920,In_1780,In_925);
or U1921 (N_1921,In_305,In_1899);
or U1922 (N_1922,In_1981,In_93);
nand U1923 (N_1923,In_1365,In_655);
nand U1924 (N_1924,In_1813,In_2133);
xnor U1925 (N_1925,In_1839,In_1861);
nor U1926 (N_1926,In_1915,In_697);
and U1927 (N_1927,In_1813,In_258);
nor U1928 (N_1928,In_789,In_2261);
and U1929 (N_1929,In_638,In_1762);
nor U1930 (N_1930,In_400,In_2378);
or U1931 (N_1931,In_2319,In_600);
or U1932 (N_1932,In_1496,In_1256);
and U1933 (N_1933,In_2377,In_1182);
nor U1934 (N_1934,In_1804,In_1974);
nand U1935 (N_1935,In_954,In_2065);
or U1936 (N_1936,In_1735,In_568);
nor U1937 (N_1937,In_1993,In_2133);
or U1938 (N_1938,In_1371,In_2264);
nor U1939 (N_1939,In_899,In_783);
and U1940 (N_1940,In_1327,In_2394);
and U1941 (N_1941,In_1019,In_2452);
and U1942 (N_1942,In_2362,In_2345);
nor U1943 (N_1943,In_2276,In_2397);
or U1944 (N_1944,In_2160,In_1881);
nand U1945 (N_1945,In_1968,In_1062);
or U1946 (N_1946,In_1358,In_2362);
and U1947 (N_1947,In_252,In_1291);
nor U1948 (N_1948,In_846,In_1871);
nand U1949 (N_1949,In_978,In_59);
nand U1950 (N_1950,In_1430,In_1898);
or U1951 (N_1951,In_2305,In_1390);
or U1952 (N_1952,In_2088,In_205);
nand U1953 (N_1953,In_1184,In_2413);
or U1954 (N_1954,In_139,In_371);
and U1955 (N_1955,In_1560,In_1006);
nand U1956 (N_1956,In_1943,In_1243);
and U1957 (N_1957,In_103,In_1641);
or U1958 (N_1958,In_1720,In_1914);
or U1959 (N_1959,In_61,In_1757);
or U1960 (N_1960,In_1691,In_788);
nor U1961 (N_1961,In_2294,In_2148);
or U1962 (N_1962,In_789,In_928);
and U1963 (N_1963,In_2262,In_652);
nand U1964 (N_1964,In_127,In_1937);
or U1965 (N_1965,In_608,In_2295);
nand U1966 (N_1966,In_1741,In_2004);
or U1967 (N_1967,In_2160,In_399);
nand U1968 (N_1968,In_551,In_1870);
or U1969 (N_1969,In_2152,In_350);
xnor U1970 (N_1970,In_2306,In_212);
nor U1971 (N_1971,In_1670,In_334);
xnor U1972 (N_1972,In_222,In_1267);
nor U1973 (N_1973,In_939,In_192);
nor U1974 (N_1974,In_2300,In_756);
and U1975 (N_1975,In_1689,In_2365);
and U1976 (N_1976,In_2149,In_2462);
or U1977 (N_1977,In_406,In_1493);
or U1978 (N_1978,In_1697,In_2314);
and U1979 (N_1979,In_2147,In_2124);
xnor U1980 (N_1980,In_901,In_1318);
and U1981 (N_1981,In_292,In_47);
and U1982 (N_1982,In_359,In_483);
or U1983 (N_1983,In_2159,In_1384);
nor U1984 (N_1984,In_2008,In_408);
and U1985 (N_1985,In_2421,In_235);
nor U1986 (N_1986,In_2172,In_1185);
and U1987 (N_1987,In_774,In_1215);
nand U1988 (N_1988,In_955,In_1122);
nand U1989 (N_1989,In_456,In_900);
xnor U1990 (N_1990,In_946,In_674);
nor U1991 (N_1991,In_989,In_454);
nand U1992 (N_1992,In_1395,In_114);
or U1993 (N_1993,In_1697,In_1123);
or U1994 (N_1994,In_1949,In_476);
or U1995 (N_1995,In_1742,In_985);
xnor U1996 (N_1996,In_1881,In_1845);
and U1997 (N_1997,In_2349,In_1170);
nor U1998 (N_1998,In_154,In_2155);
nor U1999 (N_1999,In_1938,In_808);
nand U2000 (N_2000,In_1332,In_2024);
nand U2001 (N_2001,In_2291,In_1754);
and U2002 (N_2002,In_2314,In_2396);
nor U2003 (N_2003,In_931,In_2217);
xor U2004 (N_2004,In_1268,In_1625);
and U2005 (N_2005,In_1606,In_2381);
and U2006 (N_2006,In_1828,In_1694);
or U2007 (N_2007,In_2,In_2425);
and U2008 (N_2008,In_570,In_1892);
nand U2009 (N_2009,In_425,In_1186);
nand U2010 (N_2010,In_242,In_1266);
nor U2011 (N_2011,In_2002,In_2303);
nand U2012 (N_2012,In_1432,In_1896);
nand U2013 (N_2013,In_1466,In_1434);
or U2014 (N_2014,In_390,In_1362);
nand U2015 (N_2015,In_968,In_914);
and U2016 (N_2016,In_2078,In_1761);
or U2017 (N_2017,In_8,In_215);
or U2018 (N_2018,In_1968,In_654);
or U2019 (N_2019,In_284,In_167);
nor U2020 (N_2020,In_2027,In_2299);
and U2021 (N_2021,In_440,In_1072);
nor U2022 (N_2022,In_1856,In_2044);
nand U2023 (N_2023,In_430,In_2497);
and U2024 (N_2024,In_2156,In_2032);
nand U2025 (N_2025,In_1504,In_2475);
nand U2026 (N_2026,In_974,In_204);
nand U2027 (N_2027,In_71,In_876);
nor U2028 (N_2028,In_1413,In_617);
nor U2029 (N_2029,In_1470,In_759);
and U2030 (N_2030,In_332,In_459);
and U2031 (N_2031,In_89,In_319);
and U2032 (N_2032,In_60,In_827);
or U2033 (N_2033,In_1464,In_2072);
nor U2034 (N_2034,In_2312,In_2245);
nand U2035 (N_2035,In_226,In_427);
and U2036 (N_2036,In_1049,In_1925);
nor U2037 (N_2037,In_1155,In_800);
or U2038 (N_2038,In_968,In_2237);
and U2039 (N_2039,In_2469,In_1371);
and U2040 (N_2040,In_1624,In_112);
or U2041 (N_2041,In_455,In_2472);
and U2042 (N_2042,In_216,In_2499);
nand U2043 (N_2043,In_835,In_2116);
and U2044 (N_2044,In_1455,In_1982);
nand U2045 (N_2045,In_172,In_1967);
and U2046 (N_2046,In_904,In_654);
or U2047 (N_2047,In_817,In_63);
nand U2048 (N_2048,In_920,In_1059);
or U2049 (N_2049,In_1933,In_572);
or U2050 (N_2050,In_1805,In_672);
or U2051 (N_2051,In_1688,In_2468);
or U2052 (N_2052,In_2316,In_1881);
or U2053 (N_2053,In_2240,In_1501);
or U2054 (N_2054,In_1115,In_1420);
and U2055 (N_2055,In_2256,In_1836);
and U2056 (N_2056,In_2404,In_247);
or U2057 (N_2057,In_251,In_425);
and U2058 (N_2058,In_1216,In_2215);
or U2059 (N_2059,In_1482,In_1703);
nand U2060 (N_2060,In_192,In_1444);
nor U2061 (N_2061,In_2397,In_1220);
and U2062 (N_2062,In_2109,In_804);
xnor U2063 (N_2063,In_1820,In_1712);
or U2064 (N_2064,In_373,In_1626);
and U2065 (N_2065,In_2346,In_1160);
nor U2066 (N_2066,In_2130,In_1046);
or U2067 (N_2067,In_189,In_617);
and U2068 (N_2068,In_397,In_611);
nor U2069 (N_2069,In_1283,In_1442);
nor U2070 (N_2070,In_973,In_1997);
nand U2071 (N_2071,In_1763,In_87);
xor U2072 (N_2072,In_966,In_867);
or U2073 (N_2073,In_151,In_1333);
or U2074 (N_2074,In_112,In_1595);
nor U2075 (N_2075,In_768,In_2318);
nor U2076 (N_2076,In_924,In_369);
nor U2077 (N_2077,In_301,In_641);
or U2078 (N_2078,In_1741,In_1434);
and U2079 (N_2079,In_1809,In_2497);
and U2080 (N_2080,In_594,In_1699);
nor U2081 (N_2081,In_2098,In_1522);
nand U2082 (N_2082,In_1821,In_2255);
nor U2083 (N_2083,In_1890,In_796);
nand U2084 (N_2084,In_1696,In_1719);
and U2085 (N_2085,In_1872,In_101);
nand U2086 (N_2086,In_1728,In_2196);
nand U2087 (N_2087,In_865,In_755);
nand U2088 (N_2088,In_1240,In_2080);
or U2089 (N_2089,In_47,In_1055);
xnor U2090 (N_2090,In_487,In_334);
nor U2091 (N_2091,In_2070,In_1695);
and U2092 (N_2092,In_632,In_1722);
or U2093 (N_2093,In_2388,In_1496);
nand U2094 (N_2094,In_1274,In_246);
nor U2095 (N_2095,In_257,In_1224);
and U2096 (N_2096,In_2294,In_1362);
and U2097 (N_2097,In_938,In_929);
nand U2098 (N_2098,In_1477,In_1575);
and U2099 (N_2099,In_224,In_1600);
or U2100 (N_2100,In_520,In_913);
nand U2101 (N_2101,In_1097,In_529);
or U2102 (N_2102,In_2131,In_1167);
and U2103 (N_2103,In_207,In_1797);
nor U2104 (N_2104,In_2301,In_1017);
or U2105 (N_2105,In_791,In_1969);
nor U2106 (N_2106,In_2189,In_1070);
nand U2107 (N_2107,In_2257,In_1021);
and U2108 (N_2108,In_2055,In_1255);
nor U2109 (N_2109,In_2077,In_1757);
nand U2110 (N_2110,In_250,In_303);
or U2111 (N_2111,In_2207,In_2155);
or U2112 (N_2112,In_2230,In_174);
or U2113 (N_2113,In_1671,In_1423);
xor U2114 (N_2114,In_1293,In_528);
or U2115 (N_2115,In_567,In_853);
and U2116 (N_2116,In_1372,In_1309);
and U2117 (N_2117,In_2268,In_1324);
nor U2118 (N_2118,In_765,In_225);
nor U2119 (N_2119,In_468,In_2121);
or U2120 (N_2120,In_2457,In_555);
nand U2121 (N_2121,In_1523,In_1038);
xnor U2122 (N_2122,In_517,In_1879);
nor U2123 (N_2123,In_2206,In_1637);
nand U2124 (N_2124,In_1705,In_1689);
xnor U2125 (N_2125,In_1141,In_2020);
xor U2126 (N_2126,In_1896,In_1384);
nand U2127 (N_2127,In_126,In_132);
or U2128 (N_2128,In_238,In_2316);
nor U2129 (N_2129,In_2143,In_256);
and U2130 (N_2130,In_1636,In_727);
nand U2131 (N_2131,In_2096,In_309);
nand U2132 (N_2132,In_1726,In_2441);
and U2133 (N_2133,In_2016,In_1236);
and U2134 (N_2134,In_817,In_2210);
and U2135 (N_2135,In_53,In_113);
nand U2136 (N_2136,In_861,In_481);
or U2137 (N_2137,In_1916,In_798);
nor U2138 (N_2138,In_999,In_1666);
or U2139 (N_2139,In_743,In_2167);
or U2140 (N_2140,In_309,In_1711);
nand U2141 (N_2141,In_2303,In_14);
or U2142 (N_2142,In_984,In_838);
nand U2143 (N_2143,In_436,In_2009);
nor U2144 (N_2144,In_1766,In_2432);
and U2145 (N_2145,In_926,In_2200);
nor U2146 (N_2146,In_432,In_2154);
and U2147 (N_2147,In_1542,In_2249);
and U2148 (N_2148,In_412,In_2407);
or U2149 (N_2149,In_313,In_1807);
or U2150 (N_2150,In_681,In_607);
nand U2151 (N_2151,In_552,In_757);
nand U2152 (N_2152,In_2026,In_846);
or U2153 (N_2153,In_2460,In_2351);
and U2154 (N_2154,In_528,In_1924);
nand U2155 (N_2155,In_116,In_471);
and U2156 (N_2156,In_1132,In_523);
nor U2157 (N_2157,In_157,In_1896);
and U2158 (N_2158,In_1676,In_1419);
or U2159 (N_2159,In_219,In_438);
nor U2160 (N_2160,In_1571,In_837);
nand U2161 (N_2161,In_164,In_467);
and U2162 (N_2162,In_1311,In_1639);
and U2163 (N_2163,In_175,In_1232);
nor U2164 (N_2164,In_1969,In_389);
or U2165 (N_2165,In_1948,In_582);
or U2166 (N_2166,In_1731,In_488);
nand U2167 (N_2167,In_349,In_1219);
and U2168 (N_2168,In_588,In_957);
nand U2169 (N_2169,In_328,In_593);
and U2170 (N_2170,In_653,In_415);
or U2171 (N_2171,In_1497,In_2324);
nor U2172 (N_2172,In_1405,In_1445);
nand U2173 (N_2173,In_1298,In_2285);
and U2174 (N_2174,In_159,In_1612);
nand U2175 (N_2175,In_303,In_1299);
nand U2176 (N_2176,In_1866,In_2096);
or U2177 (N_2177,In_1144,In_1585);
nand U2178 (N_2178,In_2056,In_202);
or U2179 (N_2179,In_1962,In_2149);
nand U2180 (N_2180,In_36,In_2184);
nand U2181 (N_2181,In_2060,In_58);
and U2182 (N_2182,In_1442,In_1831);
nand U2183 (N_2183,In_1627,In_1474);
and U2184 (N_2184,In_749,In_1284);
or U2185 (N_2185,In_2269,In_1625);
nor U2186 (N_2186,In_2185,In_171);
nand U2187 (N_2187,In_1193,In_1752);
and U2188 (N_2188,In_2077,In_556);
and U2189 (N_2189,In_1982,In_2464);
nand U2190 (N_2190,In_1793,In_929);
nor U2191 (N_2191,In_2435,In_257);
nand U2192 (N_2192,In_1956,In_1836);
and U2193 (N_2193,In_382,In_1981);
or U2194 (N_2194,In_80,In_1274);
or U2195 (N_2195,In_701,In_1827);
and U2196 (N_2196,In_1989,In_2466);
nand U2197 (N_2197,In_1259,In_1360);
or U2198 (N_2198,In_1198,In_1322);
nor U2199 (N_2199,In_9,In_1411);
or U2200 (N_2200,In_1494,In_2267);
xor U2201 (N_2201,In_801,In_133);
or U2202 (N_2202,In_1727,In_1933);
nand U2203 (N_2203,In_1580,In_1839);
and U2204 (N_2204,In_2219,In_1618);
nand U2205 (N_2205,In_816,In_1794);
and U2206 (N_2206,In_111,In_1557);
xnor U2207 (N_2207,In_2175,In_917);
nand U2208 (N_2208,In_605,In_624);
nor U2209 (N_2209,In_472,In_1772);
or U2210 (N_2210,In_1572,In_1322);
or U2211 (N_2211,In_1161,In_1221);
nor U2212 (N_2212,In_2359,In_478);
nor U2213 (N_2213,In_2181,In_1447);
nand U2214 (N_2214,In_385,In_733);
and U2215 (N_2215,In_1730,In_547);
nand U2216 (N_2216,In_2462,In_1691);
nand U2217 (N_2217,In_186,In_189);
nor U2218 (N_2218,In_651,In_659);
nor U2219 (N_2219,In_1304,In_1026);
nand U2220 (N_2220,In_214,In_1186);
nor U2221 (N_2221,In_964,In_247);
or U2222 (N_2222,In_659,In_2333);
and U2223 (N_2223,In_286,In_2378);
xor U2224 (N_2224,In_2055,In_2122);
nand U2225 (N_2225,In_677,In_2079);
and U2226 (N_2226,In_2165,In_2452);
nor U2227 (N_2227,In_1007,In_844);
or U2228 (N_2228,In_1106,In_2232);
or U2229 (N_2229,In_1365,In_934);
nor U2230 (N_2230,In_1195,In_1304);
nor U2231 (N_2231,In_324,In_1275);
nand U2232 (N_2232,In_1991,In_2091);
or U2233 (N_2233,In_200,In_1812);
nand U2234 (N_2234,In_487,In_1144);
or U2235 (N_2235,In_148,In_1814);
and U2236 (N_2236,In_423,In_1861);
nand U2237 (N_2237,In_1065,In_993);
nor U2238 (N_2238,In_1984,In_569);
nand U2239 (N_2239,In_1612,In_1752);
nand U2240 (N_2240,In_1325,In_44);
nor U2241 (N_2241,In_1987,In_1366);
or U2242 (N_2242,In_1795,In_1716);
nor U2243 (N_2243,In_1659,In_2366);
nand U2244 (N_2244,In_1231,In_2098);
nor U2245 (N_2245,In_1797,In_1998);
nor U2246 (N_2246,In_446,In_2031);
or U2247 (N_2247,In_1070,In_1688);
and U2248 (N_2248,In_2364,In_1317);
or U2249 (N_2249,In_463,In_1279);
and U2250 (N_2250,In_1345,In_1207);
and U2251 (N_2251,In_790,In_1873);
xnor U2252 (N_2252,In_2468,In_951);
or U2253 (N_2253,In_1040,In_2185);
and U2254 (N_2254,In_2466,In_2411);
nor U2255 (N_2255,In_249,In_1596);
nand U2256 (N_2256,In_1453,In_752);
nor U2257 (N_2257,In_1218,In_876);
nor U2258 (N_2258,In_1910,In_249);
nand U2259 (N_2259,In_1830,In_942);
nand U2260 (N_2260,In_325,In_2229);
nor U2261 (N_2261,In_193,In_908);
or U2262 (N_2262,In_2464,In_307);
nand U2263 (N_2263,In_324,In_246);
or U2264 (N_2264,In_72,In_2008);
and U2265 (N_2265,In_755,In_273);
nor U2266 (N_2266,In_2111,In_1134);
nand U2267 (N_2267,In_1912,In_1255);
or U2268 (N_2268,In_2077,In_1933);
and U2269 (N_2269,In_1002,In_16);
nor U2270 (N_2270,In_274,In_1447);
nor U2271 (N_2271,In_2438,In_1434);
nor U2272 (N_2272,In_52,In_1596);
nand U2273 (N_2273,In_2153,In_2162);
or U2274 (N_2274,In_600,In_1142);
or U2275 (N_2275,In_768,In_2413);
nor U2276 (N_2276,In_1352,In_586);
or U2277 (N_2277,In_2334,In_1525);
nand U2278 (N_2278,In_195,In_2258);
nor U2279 (N_2279,In_2246,In_2373);
or U2280 (N_2280,In_1232,In_460);
and U2281 (N_2281,In_674,In_2007);
or U2282 (N_2282,In_2381,In_1323);
and U2283 (N_2283,In_1379,In_558);
or U2284 (N_2284,In_1970,In_1095);
or U2285 (N_2285,In_671,In_221);
or U2286 (N_2286,In_1973,In_483);
nand U2287 (N_2287,In_611,In_515);
nand U2288 (N_2288,In_1081,In_938);
nand U2289 (N_2289,In_2335,In_640);
nor U2290 (N_2290,In_1332,In_321);
nand U2291 (N_2291,In_1623,In_1388);
nand U2292 (N_2292,In_1442,In_1644);
and U2293 (N_2293,In_999,In_2067);
or U2294 (N_2294,In_1213,In_2106);
and U2295 (N_2295,In_2321,In_650);
or U2296 (N_2296,In_1796,In_185);
nand U2297 (N_2297,In_1344,In_787);
or U2298 (N_2298,In_1193,In_1613);
nor U2299 (N_2299,In_1160,In_1772);
nand U2300 (N_2300,In_1915,In_1484);
and U2301 (N_2301,In_932,In_1611);
and U2302 (N_2302,In_873,In_1611);
or U2303 (N_2303,In_1044,In_841);
and U2304 (N_2304,In_1261,In_878);
or U2305 (N_2305,In_1749,In_1742);
and U2306 (N_2306,In_84,In_1914);
or U2307 (N_2307,In_1852,In_1162);
nor U2308 (N_2308,In_1373,In_2089);
nor U2309 (N_2309,In_179,In_2199);
nand U2310 (N_2310,In_514,In_1474);
and U2311 (N_2311,In_670,In_1110);
nand U2312 (N_2312,In_133,In_1790);
nand U2313 (N_2313,In_1723,In_1194);
nor U2314 (N_2314,In_2228,In_1461);
and U2315 (N_2315,In_1337,In_1235);
nand U2316 (N_2316,In_204,In_2142);
nor U2317 (N_2317,In_1017,In_1096);
nand U2318 (N_2318,In_1864,In_811);
nand U2319 (N_2319,In_2017,In_607);
or U2320 (N_2320,In_1221,In_1114);
and U2321 (N_2321,In_2064,In_1606);
nand U2322 (N_2322,In_1695,In_301);
nor U2323 (N_2323,In_1299,In_669);
nor U2324 (N_2324,In_733,In_1587);
and U2325 (N_2325,In_1556,In_1080);
and U2326 (N_2326,In_659,In_530);
or U2327 (N_2327,In_1930,In_1063);
and U2328 (N_2328,In_162,In_1126);
and U2329 (N_2329,In_1568,In_1880);
and U2330 (N_2330,In_383,In_684);
and U2331 (N_2331,In_406,In_2445);
or U2332 (N_2332,In_1490,In_930);
and U2333 (N_2333,In_1454,In_2002);
or U2334 (N_2334,In_2261,In_34);
or U2335 (N_2335,In_980,In_283);
nor U2336 (N_2336,In_560,In_1248);
nor U2337 (N_2337,In_205,In_1083);
or U2338 (N_2338,In_1501,In_900);
or U2339 (N_2339,In_2471,In_560);
nand U2340 (N_2340,In_1872,In_1311);
and U2341 (N_2341,In_988,In_2341);
nor U2342 (N_2342,In_2023,In_1542);
or U2343 (N_2343,In_1773,In_1398);
and U2344 (N_2344,In_5,In_2298);
or U2345 (N_2345,In_654,In_397);
nand U2346 (N_2346,In_1256,In_693);
nand U2347 (N_2347,In_2454,In_994);
nand U2348 (N_2348,In_722,In_780);
nor U2349 (N_2349,In_1257,In_1644);
or U2350 (N_2350,In_995,In_2242);
and U2351 (N_2351,In_1387,In_2048);
and U2352 (N_2352,In_829,In_1087);
or U2353 (N_2353,In_1732,In_1920);
or U2354 (N_2354,In_1219,In_2195);
nor U2355 (N_2355,In_880,In_1507);
nand U2356 (N_2356,In_2439,In_729);
or U2357 (N_2357,In_250,In_219);
nand U2358 (N_2358,In_873,In_1974);
nor U2359 (N_2359,In_535,In_1106);
nor U2360 (N_2360,In_736,In_1607);
or U2361 (N_2361,In_1172,In_307);
and U2362 (N_2362,In_670,In_2418);
xor U2363 (N_2363,In_674,In_1836);
nand U2364 (N_2364,In_2296,In_1157);
nand U2365 (N_2365,In_1128,In_2356);
and U2366 (N_2366,In_407,In_470);
nand U2367 (N_2367,In_1002,In_1975);
or U2368 (N_2368,In_785,In_1929);
nand U2369 (N_2369,In_1445,In_665);
nor U2370 (N_2370,In_2273,In_1116);
nor U2371 (N_2371,In_2272,In_62);
nand U2372 (N_2372,In_2097,In_2482);
nand U2373 (N_2373,In_2434,In_1778);
or U2374 (N_2374,In_23,In_809);
and U2375 (N_2375,In_1370,In_596);
nor U2376 (N_2376,In_1467,In_2329);
and U2377 (N_2377,In_1207,In_2345);
and U2378 (N_2378,In_38,In_718);
nand U2379 (N_2379,In_834,In_2346);
nor U2380 (N_2380,In_2142,In_1667);
or U2381 (N_2381,In_11,In_706);
and U2382 (N_2382,In_2117,In_374);
nor U2383 (N_2383,In_652,In_2370);
and U2384 (N_2384,In_1820,In_597);
nand U2385 (N_2385,In_1682,In_1013);
nand U2386 (N_2386,In_1337,In_2318);
nor U2387 (N_2387,In_208,In_1591);
nand U2388 (N_2388,In_559,In_1602);
nand U2389 (N_2389,In_1748,In_1991);
nor U2390 (N_2390,In_193,In_88);
nor U2391 (N_2391,In_1474,In_831);
nor U2392 (N_2392,In_2403,In_1732);
nand U2393 (N_2393,In_1448,In_715);
and U2394 (N_2394,In_240,In_1233);
nand U2395 (N_2395,In_1483,In_1539);
nor U2396 (N_2396,In_2356,In_498);
or U2397 (N_2397,In_1689,In_1871);
and U2398 (N_2398,In_2227,In_547);
nand U2399 (N_2399,In_33,In_917);
or U2400 (N_2400,In_794,In_539);
and U2401 (N_2401,In_881,In_2239);
and U2402 (N_2402,In_1555,In_2297);
and U2403 (N_2403,In_829,In_765);
and U2404 (N_2404,In_1104,In_961);
and U2405 (N_2405,In_177,In_2146);
xor U2406 (N_2406,In_1841,In_1368);
and U2407 (N_2407,In_929,In_2381);
or U2408 (N_2408,In_1206,In_895);
nand U2409 (N_2409,In_1162,In_1921);
nand U2410 (N_2410,In_2112,In_2109);
nand U2411 (N_2411,In_2071,In_863);
and U2412 (N_2412,In_1716,In_449);
nor U2413 (N_2413,In_2354,In_353);
or U2414 (N_2414,In_869,In_1131);
or U2415 (N_2415,In_791,In_823);
nor U2416 (N_2416,In_2477,In_608);
nor U2417 (N_2417,In_1902,In_1845);
nand U2418 (N_2418,In_2079,In_1591);
and U2419 (N_2419,In_1252,In_2058);
nand U2420 (N_2420,In_1751,In_492);
nand U2421 (N_2421,In_180,In_2133);
and U2422 (N_2422,In_1947,In_2079);
nor U2423 (N_2423,In_2033,In_1981);
or U2424 (N_2424,In_1307,In_1170);
nor U2425 (N_2425,In_771,In_593);
and U2426 (N_2426,In_1643,In_275);
xnor U2427 (N_2427,In_1579,In_689);
and U2428 (N_2428,In_168,In_804);
nor U2429 (N_2429,In_1502,In_474);
nor U2430 (N_2430,In_2352,In_1036);
and U2431 (N_2431,In_1205,In_708);
nand U2432 (N_2432,In_970,In_124);
nor U2433 (N_2433,In_885,In_665);
or U2434 (N_2434,In_2460,In_91);
or U2435 (N_2435,In_210,In_2220);
or U2436 (N_2436,In_1961,In_1114);
nand U2437 (N_2437,In_2172,In_98);
and U2438 (N_2438,In_1975,In_560);
and U2439 (N_2439,In_1153,In_1318);
or U2440 (N_2440,In_116,In_1104);
nand U2441 (N_2441,In_257,In_1831);
and U2442 (N_2442,In_1054,In_2266);
and U2443 (N_2443,In_1240,In_1165);
nand U2444 (N_2444,In_968,In_190);
and U2445 (N_2445,In_1873,In_31);
and U2446 (N_2446,In_761,In_14);
and U2447 (N_2447,In_1294,In_1619);
nand U2448 (N_2448,In_1085,In_1302);
and U2449 (N_2449,In_1475,In_1427);
nor U2450 (N_2450,In_2409,In_2077);
xor U2451 (N_2451,In_617,In_2026);
nor U2452 (N_2452,In_596,In_1360);
nand U2453 (N_2453,In_1195,In_2322);
nor U2454 (N_2454,In_1231,In_1066);
or U2455 (N_2455,In_690,In_303);
nor U2456 (N_2456,In_1334,In_306);
and U2457 (N_2457,In_1505,In_896);
or U2458 (N_2458,In_462,In_985);
and U2459 (N_2459,In_750,In_2467);
nand U2460 (N_2460,In_1222,In_650);
and U2461 (N_2461,In_2447,In_111);
or U2462 (N_2462,In_1756,In_988);
nand U2463 (N_2463,In_1151,In_755);
or U2464 (N_2464,In_987,In_469);
nand U2465 (N_2465,In_676,In_349);
nor U2466 (N_2466,In_465,In_490);
nand U2467 (N_2467,In_1950,In_1666);
or U2468 (N_2468,In_519,In_1416);
nor U2469 (N_2469,In_512,In_1857);
nand U2470 (N_2470,In_842,In_211);
nand U2471 (N_2471,In_2048,In_41);
or U2472 (N_2472,In_654,In_214);
nor U2473 (N_2473,In_21,In_2039);
or U2474 (N_2474,In_850,In_705);
or U2475 (N_2475,In_1250,In_711);
and U2476 (N_2476,In_2496,In_287);
nand U2477 (N_2477,In_2006,In_104);
or U2478 (N_2478,In_1600,In_753);
nand U2479 (N_2479,In_72,In_1276);
nand U2480 (N_2480,In_2095,In_430);
nor U2481 (N_2481,In_1448,In_294);
or U2482 (N_2482,In_33,In_1552);
or U2483 (N_2483,In_1410,In_1915);
nor U2484 (N_2484,In_2166,In_739);
or U2485 (N_2485,In_2329,In_1317);
or U2486 (N_2486,In_2469,In_861);
and U2487 (N_2487,In_286,In_971);
nor U2488 (N_2488,In_121,In_1155);
or U2489 (N_2489,In_1931,In_8);
nand U2490 (N_2490,In_1375,In_78);
nor U2491 (N_2491,In_1466,In_899);
or U2492 (N_2492,In_1749,In_428);
and U2493 (N_2493,In_1384,In_1058);
and U2494 (N_2494,In_2024,In_563);
or U2495 (N_2495,In_872,In_2268);
nor U2496 (N_2496,In_236,In_1928);
nor U2497 (N_2497,In_1557,In_487);
or U2498 (N_2498,In_660,In_245);
or U2499 (N_2499,In_69,In_1618);
or U2500 (N_2500,In_1083,In_2281);
nand U2501 (N_2501,In_835,In_1850);
xor U2502 (N_2502,In_1117,In_1028);
xnor U2503 (N_2503,In_1960,In_2369);
and U2504 (N_2504,In_1091,In_919);
nand U2505 (N_2505,In_2060,In_1901);
nor U2506 (N_2506,In_1974,In_746);
nand U2507 (N_2507,In_1338,In_169);
nand U2508 (N_2508,In_2232,In_2252);
nand U2509 (N_2509,In_1507,In_1068);
or U2510 (N_2510,In_827,In_2306);
nand U2511 (N_2511,In_1426,In_1705);
nand U2512 (N_2512,In_2322,In_1087);
and U2513 (N_2513,In_264,In_2239);
nand U2514 (N_2514,In_201,In_194);
nand U2515 (N_2515,In_767,In_1719);
and U2516 (N_2516,In_1017,In_569);
or U2517 (N_2517,In_1759,In_226);
nor U2518 (N_2518,In_686,In_1755);
nand U2519 (N_2519,In_2474,In_838);
nor U2520 (N_2520,In_1948,In_739);
nor U2521 (N_2521,In_587,In_432);
nand U2522 (N_2522,In_679,In_1182);
and U2523 (N_2523,In_1564,In_533);
and U2524 (N_2524,In_901,In_324);
or U2525 (N_2525,In_2023,In_2407);
and U2526 (N_2526,In_1047,In_1023);
nor U2527 (N_2527,In_803,In_1059);
or U2528 (N_2528,In_853,In_2029);
or U2529 (N_2529,In_2190,In_282);
nand U2530 (N_2530,In_779,In_489);
nand U2531 (N_2531,In_2411,In_2210);
nor U2532 (N_2532,In_2170,In_1124);
nand U2533 (N_2533,In_548,In_2340);
nand U2534 (N_2534,In_168,In_1826);
nand U2535 (N_2535,In_1153,In_142);
nand U2536 (N_2536,In_170,In_2330);
nor U2537 (N_2537,In_1899,In_229);
and U2538 (N_2538,In_1185,In_2424);
and U2539 (N_2539,In_1485,In_2434);
or U2540 (N_2540,In_2379,In_99);
and U2541 (N_2541,In_2063,In_1389);
nor U2542 (N_2542,In_2351,In_97);
nand U2543 (N_2543,In_2242,In_1523);
and U2544 (N_2544,In_781,In_1786);
nand U2545 (N_2545,In_1872,In_456);
nand U2546 (N_2546,In_2417,In_1736);
nor U2547 (N_2547,In_1729,In_59);
nor U2548 (N_2548,In_1018,In_2335);
nor U2549 (N_2549,In_2028,In_1094);
and U2550 (N_2550,In_1464,In_1167);
nor U2551 (N_2551,In_1881,In_471);
or U2552 (N_2552,In_1396,In_1136);
and U2553 (N_2553,In_2291,In_1618);
nor U2554 (N_2554,In_202,In_2081);
or U2555 (N_2555,In_538,In_1973);
nor U2556 (N_2556,In_2379,In_2173);
xnor U2557 (N_2557,In_720,In_2360);
or U2558 (N_2558,In_640,In_886);
and U2559 (N_2559,In_1665,In_1976);
and U2560 (N_2560,In_1762,In_1183);
nor U2561 (N_2561,In_2270,In_47);
or U2562 (N_2562,In_148,In_1812);
and U2563 (N_2563,In_1111,In_280);
nor U2564 (N_2564,In_1548,In_776);
xor U2565 (N_2565,In_487,In_1633);
and U2566 (N_2566,In_1422,In_1208);
nor U2567 (N_2567,In_1029,In_1136);
or U2568 (N_2568,In_2162,In_1442);
or U2569 (N_2569,In_530,In_1508);
and U2570 (N_2570,In_2344,In_1164);
and U2571 (N_2571,In_790,In_6);
nand U2572 (N_2572,In_1645,In_445);
nor U2573 (N_2573,In_305,In_2448);
nand U2574 (N_2574,In_633,In_2303);
or U2575 (N_2575,In_857,In_2244);
nor U2576 (N_2576,In_1904,In_1573);
xnor U2577 (N_2577,In_1842,In_1683);
nand U2578 (N_2578,In_601,In_40);
nand U2579 (N_2579,In_2101,In_2433);
nand U2580 (N_2580,In_2187,In_514);
and U2581 (N_2581,In_1942,In_1250);
and U2582 (N_2582,In_1311,In_1936);
or U2583 (N_2583,In_1103,In_712);
nor U2584 (N_2584,In_1667,In_1101);
and U2585 (N_2585,In_1427,In_2347);
or U2586 (N_2586,In_2460,In_1852);
and U2587 (N_2587,In_184,In_1924);
nor U2588 (N_2588,In_2362,In_902);
and U2589 (N_2589,In_657,In_714);
nor U2590 (N_2590,In_871,In_1300);
nand U2591 (N_2591,In_688,In_853);
and U2592 (N_2592,In_1191,In_1024);
and U2593 (N_2593,In_1996,In_227);
nor U2594 (N_2594,In_1846,In_945);
and U2595 (N_2595,In_170,In_1528);
nor U2596 (N_2596,In_1563,In_1901);
and U2597 (N_2597,In_1881,In_1750);
and U2598 (N_2598,In_2131,In_1298);
nand U2599 (N_2599,In_1752,In_364);
nand U2600 (N_2600,In_2413,In_1950);
and U2601 (N_2601,In_2367,In_2076);
or U2602 (N_2602,In_13,In_1572);
xor U2603 (N_2603,In_335,In_1675);
and U2604 (N_2604,In_1878,In_853);
and U2605 (N_2605,In_586,In_1019);
or U2606 (N_2606,In_406,In_543);
or U2607 (N_2607,In_348,In_2355);
or U2608 (N_2608,In_2256,In_1708);
nand U2609 (N_2609,In_1868,In_1199);
and U2610 (N_2610,In_1964,In_2318);
xnor U2611 (N_2611,In_829,In_848);
nand U2612 (N_2612,In_2351,In_815);
or U2613 (N_2613,In_365,In_419);
and U2614 (N_2614,In_1144,In_2099);
nor U2615 (N_2615,In_452,In_818);
and U2616 (N_2616,In_379,In_687);
nor U2617 (N_2617,In_360,In_438);
nand U2618 (N_2618,In_877,In_1790);
nor U2619 (N_2619,In_500,In_2222);
nand U2620 (N_2620,In_1075,In_1017);
xor U2621 (N_2621,In_1710,In_693);
or U2622 (N_2622,In_1054,In_58);
and U2623 (N_2623,In_1412,In_917);
nor U2624 (N_2624,In_2017,In_1755);
nor U2625 (N_2625,In_2493,In_817);
or U2626 (N_2626,In_941,In_2273);
or U2627 (N_2627,In_2076,In_2282);
nor U2628 (N_2628,In_422,In_656);
and U2629 (N_2629,In_1895,In_2138);
or U2630 (N_2630,In_2189,In_912);
or U2631 (N_2631,In_1025,In_393);
nand U2632 (N_2632,In_405,In_97);
nor U2633 (N_2633,In_1486,In_2079);
and U2634 (N_2634,In_1243,In_2320);
nor U2635 (N_2635,In_1919,In_497);
xnor U2636 (N_2636,In_2390,In_783);
nor U2637 (N_2637,In_1369,In_2331);
or U2638 (N_2638,In_2183,In_113);
xnor U2639 (N_2639,In_1169,In_1475);
and U2640 (N_2640,In_339,In_2139);
nand U2641 (N_2641,In_16,In_554);
nor U2642 (N_2642,In_2071,In_177);
and U2643 (N_2643,In_326,In_1496);
nor U2644 (N_2644,In_777,In_912);
or U2645 (N_2645,In_1335,In_1063);
and U2646 (N_2646,In_1845,In_1330);
and U2647 (N_2647,In_763,In_1371);
nor U2648 (N_2648,In_1023,In_291);
and U2649 (N_2649,In_2126,In_343);
nor U2650 (N_2650,In_1178,In_2454);
or U2651 (N_2651,In_1332,In_2258);
nor U2652 (N_2652,In_2463,In_678);
nor U2653 (N_2653,In_578,In_1292);
xnor U2654 (N_2654,In_1637,In_1857);
nand U2655 (N_2655,In_2243,In_2178);
or U2656 (N_2656,In_1699,In_2163);
and U2657 (N_2657,In_1576,In_1902);
and U2658 (N_2658,In_770,In_3);
or U2659 (N_2659,In_1757,In_1662);
and U2660 (N_2660,In_415,In_1566);
nor U2661 (N_2661,In_278,In_581);
or U2662 (N_2662,In_878,In_2429);
or U2663 (N_2663,In_47,In_1129);
nor U2664 (N_2664,In_224,In_426);
or U2665 (N_2665,In_30,In_636);
nor U2666 (N_2666,In_934,In_1123);
and U2667 (N_2667,In_1281,In_457);
nor U2668 (N_2668,In_421,In_764);
or U2669 (N_2669,In_404,In_1938);
and U2670 (N_2670,In_1605,In_1939);
nor U2671 (N_2671,In_1195,In_2442);
or U2672 (N_2672,In_911,In_1504);
or U2673 (N_2673,In_537,In_2457);
or U2674 (N_2674,In_437,In_956);
and U2675 (N_2675,In_1762,In_1366);
or U2676 (N_2676,In_240,In_249);
nand U2677 (N_2677,In_2195,In_1242);
nand U2678 (N_2678,In_1394,In_1558);
nor U2679 (N_2679,In_2338,In_402);
and U2680 (N_2680,In_1899,In_1258);
and U2681 (N_2681,In_584,In_453);
or U2682 (N_2682,In_376,In_2483);
xor U2683 (N_2683,In_1649,In_1744);
or U2684 (N_2684,In_395,In_1262);
nor U2685 (N_2685,In_2412,In_2026);
nand U2686 (N_2686,In_2256,In_1129);
nor U2687 (N_2687,In_2210,In_860);
xor U2688 (N_2688,In_1220,In_1519);
or U2689 (N_2689,In_1597,In_2333);
and U2690 (N_2690,In_1793,In_2314);
and U2691 (N_2691,In_794,In_138);
or U2692 (N_2692,In_2220,In_1175);
xor U2693 (N_2693,In_588,In_411);
and U2694 (N_2694,In_1291,In_233);
and U2695 (N_2695,In_1579,In_1507);
and U2696 (N_2696,In_1649,In_970);
nand U2697 (N_2697,In_2127,In_2058);
or U2698 (N_2698,In_1972,In_603);
nand U2699 (N_2699,In_75,In_29);
or U2700 (N_2700,In_465,In_2451);
or U2701 (N_2701,In_1299,In_1106);
and U2702 (N_2702,In_218,In_2353);
nand U2703 (N_2703,In_1078,In_1207);
or U2704 (N_2704,In_2029,In_1036);
or U2705 (N_2705,In_827,In_1261);
nor U2706 (N_2706,In_867,In_4);
nor U2707 (N_2707,In_2340,In_1472);
nor U2708 (N_2708,In_2352,In_2413);
nand U2709 (N_2709,In_1454,In_2430);
nor U2710 (N_2710,In_2194,In_1946);
and U2711 (N_2711,In_2192,In_572);
nand U2712 (N_2712,In_1484,In_1761);
and U2713 (N_2713,In_2474,In_447);
or U2714 (N_2714,In_2178,In_1525);
nor U2715 (N_2715,In_2156,In_839);
nand U2716 (N_2716,In_2408,In_449);
xnor U2717 (N_2717,In_44,In_999);
and U2718 (N_2718,In_392,In_928);
or U2719 (N_2719,In_78,In_1729);
nor U2720 (N_2720,In_1928,In_331);
and U2721 (N_2721,In_1695,In_624);
nand U2722 (N_2722,In_210,In_1003);
and U2723 (N_2723,In_391,In_129);
nor U2724 (N_2724,In_257,In_2249);
and U2725 (N_2725,In_443,In_744);
xnor U2726 (N_2726,In_1957,In_193);
nor U2727 (N_2727,In_2164,In_1292);
or U2728 (N_2728,In_222,In_1073);
nor U2729 (N_2729,In_682,In_803);
nor U2730 (N_2730,In_1317,In_1506);
nand U2731 (N_2731,In_165,In_339);
and U2732 (N_2732,In_716,In_2069);
nand U2733 (N_2733,In_772,In_321);
and U2734 (N_2734,In_1770,In_128);
or U2735 (N_2735,In_1017,In_1227);
nand U2736 (N_2736,In_1801,In_1658);
nand U2737 (N_2737,In_757,In_1042);
and U2738 (N_2738,In_2279,In_1095);
or U2739 (N_2739,In_146,In_258);
nand U2740 (N_2740,In_2199,In_371);
nor U2741 (N_2741,In_384,In_1146);
nand U2742 (N_2742,In_382,In_1622);
and U2743 (N_2743,In_1854,In_809);
and U2744 (N_2744,In_714,In_1852);
nand U2745 (N_2745,In_1816,In_1548);
nand U2746 (N_2746,In_1659,In_1007);
nor U2747 (N_2747,In_724,In_2380);
or U2748 (N_2748,In_682,In_227);
xor U2749 (N_2749,In_1192,In_2329);
nand U2750 (N_2750,In_739,In_337);
and U2751 (N_2751,In_1504,In_499);
and U2752 (N_2752,In_1114,In_2077);
or U2753 (N_2753,In_813,In_1562);
or U2754 (N_2754,In_1247,In_305);
xnor U2755 (N_2755,In_1350,In_2481);
or U2756 (N_2756,In_1192,In_1419);
and U2757 (N_2757,In_1881,In_1991);
nand U2758 (N_2758,In_1711,In_1922);
or U2759 (N_2759,In_1362,In_2190);
and U2760 (N_2760,In_93,In_1904);
nor U2761 (N_2761,In_2382,In_95);
nor U2762 (N_2762,In_1830,In_2072);
and U2763 (N_2763,In_1540,In_358);
and U2764 (N_2764,In_643,In_707);
nand U2765 (N_2765,In_1556,In_75);
nand U2766 (N_2766,In_2130,In_13);
nand U2767 (N_2767,In_886,In_508);
nor U2768 (N_2768,In_2074,In_729);
or U2769 (N_2769,In_533,In_589);
nand U2770 (N_2770,In_2471,In_2380);
nand U2771 (N_2771,In_1060,In_706);
and U2772 (N_2772,In_2198,In_2108);
and U2773 (N_2773,In_585,In_376);
nor U2774 (N_2774,In_2071,In_1970);
nand U2775 (N_2775,In_2277,In_260);
nand U2776 (N_2776,In_1065,In_1402);
nand U2777 (N_2777,In_1928,In_15);
nand U2778 (N_2778,In_560,In_50);
and U2779 (N_2779,In_1818,In_1908);
nor U2780 (N_2780,In_386,In_619);
and U2781 (N_2781,In_1876,In_1488);
and U2782 (N_2782,In_1285,In_1582);
xnor U2783 (N_2783,In_98,In_1614);
and U2784 (N_2784,In_2068,In_1779);
and U2785 (N_2785,In_640,In_1439);
or U2786 (N_2786,In_221,In_75);
or U2787 (N_2787,In_511,In_2481);
nor U2788 (N_2788,In_1726,In_1437);
or U2789 (N_2789,In_2256,In_1161);
and U2790 (N_2790,In_933,In_321);
nor U2791 (N_2791,In_1091,In_1485);
and U2792 (N_2792,In_2392,In_935);
or U2793 (N_2793,In_2380,In_571);
xor U2794 (N_2794,In_1710,In_1504);
nor U2795 (N_2795,In_2298,In_25);
nor U2796 (N_2796,In_1646,In_1462);
nand U2797 (N_2797,In_542,In_1206);
and U2798 (N_2798,In_1172,In_227);
or U2799 (N_2799,In_1267,In_2144);
or U2800 (N_2800,In_1117,In_1491);
nor U2801 (N_2801,In_1337,In_1962);
nor U2802 (N_2802,In_2206,In_111);
nand U2803 (N_2803,In_1891,In_272);
nor U2804 (N_2804,In_2006,In_1084);
nor U2805 (N_2805,In_1384,In_1154);
or U2806 (N_2806,In_1573,In_100);
or U2807 (N_2807,In_2248,In_2280);
nand U2808 (N_2808,In_2411,In_587);
nand U2809 (N_2809,In_1232,In_2384);
nand U2810 (N_2810,In_812,In_65);
nand U2811 (N_2811,In_1755,In_694);
or U2812 (N_2812,In_1391,In_1431);
and U2813 (N_2813,In_88,In_315);
and U2814 (N_2814,In_389,In_2203);
nor U2815 (N_2815,In_1523,In_798);
nand U2816 (N_2816,In_563,In_2444);
nand U2817 (N_2817,In_1408,In_572);
nor U2818 (N_2818,In_94,In_2308);
nor U2819 (N_2819,In_2208,In_429);
or U2820 (N_2820,In_522,In_419);
nor U2821 (N_2821,In_694,In_1070);
or U2822 (N_2822,In_1576,In_1693);
and U2823 (N_2823,In_1625,In_324);
nor U2824 (N_2824,In_2336,In_2435);
or U2825 (N_2825,In_324,In_460);
nand U2826 (N_2826,In_2024,In_2425);
nand U2827 (N_2827,In_279,In_1253);
or U2828 (N_2828,In_2283,In_139);
nor U2829 (N_2829,In_987,In_1561);
or U2830 (N_2830,In_1467,In_1885);
and U2831 (N_2831,In_764,In_1884);
nor U2832 (N_2832,In_1800,In_2017);
nand U2833 (N_2833,In_1881,In_687);
nor U2834 (N_2834,In_1953,In_1285);
and U2835 (N_2835,In_1111,In_171);
and U2836 (N_2836,In_2291,In_1635);
nor U2837 (N_2837,In_1365,In_118);
or U2838 (N_2838,In_2025,In_2028);
nand U2839 (N_2839,In_1808,In_1508);
nand U2840 (N_2840,In_1659,In_1805);
nand U2841 (N_2841,In_2400,In_428);
xor U2842 (N_2842,In_1733,In_2382);
or U2843 (N_2843,In_1714,In_1893);
xnor U2844 (N_2844,In_496,In_1001);
nor U2845 (N_2845,In_757,In_1631);
or U2846 (N_2846,In_2290,In_560);
or U2847 (N_2847,In_870,In_511);
and U2848 (N_2848,In_480,In_690);
xor U2849 (N_2849,In_1467,In_1);
nor U2850 (N_2850,In_1397,In_823);
nor U2851 (N_2851,In_877,In_1613);
nor U2852 (N_2852,In_957,In_710);
and U2853 (N_2853,In_1566,In_564);
nor U2854 (N_2854,In_2353,In_2322);
xnor U2855 (N_2855,In_2342,In_1262);
or U2856 (N_2856,In_786,In_669);
or U2857 (N_2857,In_1952,In_395);
nor U2858 (N_2858,In_917,In_1695);
nand U2859 (N_2859,In_1956,In_75);
or U2860 (N_2860,In_1527,In_1079);
nand U2861 (N_2861,In_567,In_96);
nand U2862 (N_2862,In_543,In_202);
xnor U2863 (N_2863,In_863,In_994);
nand U2864 (N_2864,In_456,In_854);
nand U2865 (N_2865,In_1657,In_1745);
or U2866 (N_2866,In_1910,In_151);
or U2867 (N_2867,In_1812,In_485);
and U2868 (N_2868,In_1045,In_2451);
or U2869 (N_2869,In_578,In_2483);
or U2870 (N_2870,In_2230,In_1038);
and U2871 (N_2871,In_672,In_404);
and U2872 (N_2872,In_114,In_342);
and U2873 (N_2873,In_796,In_431);
nor U2874 (N_2874,In_1388,In_2252);
and U2875 (N_2875,In_1559,In_928);
or U2876 (N_2876,In_1720,In_1390);
nand U2877 (N_2877,In_2137,In_611);
or U2878 (N_2878,In_2270,In_924);
nand U2879 (N_2879,In_55,In_1203);
nor U2880 (N_2880,In_14,In_2132);
xor U2881 (N_2881,In_1835,In_897);
and U2882 (N_2882,In_1338,In_2180);
xnor U2883 (N_2883,In_1766,In_264);
nor U2884 (N_2884,In_1354,In_1655);
and U2885 (N_2885,In_1847,In_2279);
nor U2886 (N_2886,In_942,In_1456);
nand U2887 (N_2887,In_1179,In_153);
nor U2888 (N_2888,In_166,In_0);
nand U2889 (N_2889,In_1231,In_1155);
and U2890 (N_2890,In_1285,In_1179);
nor U2891 (N_2891,In_1477,In_1647);
nor U2892 (N_2892,In_1123,In_1840);
nand U2893 (N_2893,In_1027,In_1499);
or U2894 (N_2894,In_1088,In_2253);
nor U2895 (N_2895,In_648,In_27);
nand U2896 (N_2896,In_484,In_635);
nand U2897 (N_2897,In_2216,In_1090);
nor U2898 (N_2898,In_1901,In_1436);
nand U2899 (N_2899,In_1503,In_247);
nand U2900 (N_2900,In_1085,In_1478);
and U2901 (N_2901,In_741,In_1045);
or U2902 (N_2902,In_1929,In_2185);
nor U2903 (N_2903,In_1033,In_1253);
nor U2904 (N_2904,In_1491,In_1326);
or U2905 (N_2905,In_1178,In_60);
and U2906 (N_2906,In_1648,In_2121);
nand U2907 (N_2907,In_969,In_1475);
nand U2908 (N_2908,In_2108,In_351);
nor U2909 (N_2909,In_2150,In_7);
and U2910 (N_2910,In_1830,In_2229);
nand U2911 (N_2911,In_91,In_102);
nand U2912 (N_2912,In_228,In_1107);
nand U2913 (N_2913,In_132,In_450);
or U2914 (N_2914,In_1195,In_2098);
and U2915 (N_2915,In_186,In_880);
nand U2916 (N_2916,In_82,In_2358);
nor U2917 (N_2917,In_50,In_1129);
nor U2918 (N_2918,In_667,In_1203);
nand U2919 (N_2919,In_806,In_1154);
nand U2920 (N_2920,In_1498,In_1976);
and U2921 (N_2921,In_1957,In_981);
nand U2922 (N_2922,In_2039,In_567);
nor U2923 (N_2923,In_1987,In_439);
and U2924 (N_2924,In_245,In_103);
nand U2925 (N_2925,In_1623,In_1110);
or U2926 (N_2926,In_890,In_2315);
or U2927 (N_2927,In_441,In_1663);
xor U2928 (N_2928,In_965,In_838);
nand U2929 (N_2929,In_1537,In_2195);
nand U2930 (N_2930,In_1415,In_1184);
nand U2931 (N_2931,In_398,In_2308);
or U2932 (N_2932,In_1952,In_1577);
nor U2933 (N_2933,In_1957,In_2221);
or U2934 (N_2934,In_2169,In_2331);
or U2935 (N_2935,In_1318,In_444);
nor U2936 (N_2936,In_2240,In_786);
or U2937 (N_2937,In_2494,In_835);
nand U2938 (N_2938,In_295,In_2462);
nor U2939 (N_2939,In_1487,In_2049);
nor U2940 (N_2940,In_758,In_760);
and U2941 (N_2941,In_2474,In_1336);
and U2942 (N_2942,In_1614,In_1230);
and U2943 (N_2943,In_552,In_1230);
nand U2944 (N_2944,In_1798,In_1082);
nand U2945 (N_2945,In_1350,In_1771);
nand U2946 (N_2946,In_1973,In_648);
or U2947 (N_2947,In_1558,In_2023);
nor U2948 (N_2948,In_2091,In_1965);
nand U2949 (N_2949,In_1359,In_150);
nor U2950 (N_2950,In_1377,In_2082);
nand U2951 (N_2951,In_443,In_675);
nand U2952 (N_2952,In_481,In_1747);
nand U2953 (N_2953,In_1335,In_1429);
or U2954 (N_2954,In_588,In_882);
nand U2955 (N_2955,In_1079,In_131);
nor U2956 (N_2956,In_1920,In_1929);
nand U2957 (N_2957,In_1394,In_1303);
or U2958 (N_2958,In_1094,In_2386);
nand U2959 (N_2959,In_566,In_1626);
and U2960 (N_2960,In_1247,In_628);
or U2961 (N_2961,In_68,In_732);
and U2962 (N_2962,In_606,In_1706);
nand U2963 (N_2963,In_2004,In_211);
nand U2964 (N_2964,In_1338,In_1061);
or U2965 (N_2965,In_1703,In_1285);
nor U2966 (N_2966,In_413,In_1305);
or U2967 (N_2967,In_401,In_1544);
nor U2968 (N_2968,In_974,In_358);
or U2969 (N_2969,In_1805,In_922);
nor U2970 (N_2970,In_2191,In_996);
nor U2971 (N_2971,In_415,In_2054);
and U2972 (N_2972,In_95,In_1847);
nor U2973 (N_2973,In_324,In_199);
or U2974 (N_2974,In_544,In_20);
nand U2975 (N_2975,In_932,In_1539);
or U2976 (N_2976,In_359,In_1574);
nor U2977 (N_2977,In_452,In_235);
or U2978 (N_2978,In_981,In_1232);
nand U2979 (N_2979,In_1452,In_205);
or U2980 (N_2980,In_843,In_2040);
or U2981 (N_2981,In_2415,In_544);
and U2982 (N_2982,In_466,In_2349);
nand U2983 (N_2983,In_1592,In_316);
and U2984 (N_2984,In_2135,In_1912);
nand U2985 (N_2985,In_58,In_1531);
and U2986 (N_2986,In_481,In_1325);
nor U2987 (N_2987,In_1563,In_250);
and U2988 (N_2988,In_1294,In_1485);
xnor U2989 (N_2989,In_1934,In_1849);
nor U2990 (N_2990,In_1609,In_51);
and U2991 (N_2991,In_1593,In_2340);
nor U2992 (N_2992,In_1000,In_1264);
nor U2993 (N_2993,In_443,In_2118);
nand U2994 (N_2994,In_713,In_835);
nor U2995 (N_2995,In_177,In_2102);
or U2996 (N_2996,In_2363,In_87);
or U2997 (N_2997,In_974,In_540);
nand U2998 (N_2998,In_1979,In_2006);
and U2999 (N_2999,In_2491,In_2230);
nor U3000 (N_3000,In_1426,In_537);
and U3001 (N_3001,In_1701,In_246);
xor U3002 (N_3002,In_1136,In_974);
and U3003 (N_3003,In_365,In_1049);
or U3004 (N_3004,In_1477,In_1771);
or U3005 (N_3005,In_676,In_2456);
nand U3006 (N_3006,In_1196,In_1972);
or U3007 (N_3007,In_1769,In_615);
xor U3008 (N_3008,In_903,In_551);
nand U3009 (N_3009,In_1803,In_1020);
nor U3010 (N_3010,In_2424,In_771);
nand U3011 (N_3011,In_2447,In_1050);
xor U3012 (N_3012,In_2383,In_811);
nor U3013 (N_3013,In_1261,In_1910);
and U3014 (N_3014,In_1101,In_2407);
and U3015 (N_3015,In_1673,In_1191);
or U3016 (N_3016,In_2248,In_1872);
and U3017 (N_3017,In_2358,In_425);
nor U3018 (N_3018,In_1874,In_2077);
nand U3019 (N_3019,In_1769,In_1839);
nand U3020 (N_3020,In_64,In_1728);
and U3021 (N_3021,In_2054,In_533);
and U3022 (N_3022,In_2171,In_975);
or U3023 (N_3023,In_1523,In_1086);
or U3024 (N_3024,In_663,In_1681);
or U3025 (N_3025,In_1064,In_1806);
xor U3026 (N_3026,In_2049,In_884);
and U3027 (N_3027,In_85,In_1795);
or U3028 (N_3028,In_1717,In_688);
nor U3029 (N_3029,In_276,In_1888);
or U3030 (N_3030,In_1817,In_853);
nand U3031 (N_3031,In_2489,In_2404);
nand U3032 (N_3032,In_2497,In_2076);
nand U3033 (N_3033,In_263,In_1314);
or U3034 (N_3034,In_102,In_1942);
nand U3035 (N_3035,In_199,In_1047);
and U3036 (N_3036,In_2402,In_2147);
and U3037 (N_3037,In_1866,In_831);
or U3038 (N_3038,In_2429,In_196);
nand U3039 (N_3039,In_803,In_1199);
nand U3040 (N_3040,In_1626,In_174);
nand U3041 (N_3041,In_1364,In_2450);
or U3042 (N_3042,In_185,In_101);
and U3043 (N_3043,In_119,In_2209);
or U3044 (N_3044,In_796,In_1192);
or U3045 (N_3045,In_1994,In_2119);
nand U3046 (N_3046,In_2489,In_959);
and U3047 (N_3047,In_255,In_2051);
or U3048 (N_3048,In_1105,In_908);
and U3049 (N_3049,In_553,In_2243);
nand U3050 (N_3050,In_2054,In_1024);
and U3051 (N_3051,In_1560,In_1728);
and U3052 (N_3052,In_2303,In_707);
or U3053 (N_3053,In_1488,In_691);
nand U3054 (N_3054,In_2289,In_1143);
nand U3055 (N_3055,In_1917,In_1642);
nor U3056 (N_3056,In_1309,In_1878);
and U3057 (N_3057,In_804,In_2135);
and U3058 (N_3058,In_707,In_1083);
nor U3059 (N_3059,In_3,In_2444);
nand U3060 (N_3060,In_822,In_1433);
nand U3061 (N_3061,In_1029,In_1824);
and U3062 (N_3062,In_645,In_764);
nand U3063 (N_3063,In_773,In_1553);
nand U3064 (N_3064,In_601,In_1592);
and U3065 (N_3065,In_282,In_1900);
or U3066 (N_3066,In_2339,In_2109);
nor U3067 (N_3067,In_195,In_1337);
and U3068 (N_3068,In_196,In_293);
or U3069 (N_3069,In_2087,In_1356);
or U3070 (N_3070,In_757,In_2383);
nor U3071 (N_3071,In_1143,In_420);
nor U3072 (N_3072,In_794,In_2135);
nand U3073 (N_3073,In_1394,In_611);
nor U3074 (N_3074,In_1011,In_932);
nor U3075 (N_3075,In_1831,In_1645);
and U3076 (N_3076,In_1594,In_1886);
xor U3077 (N_3077,In_1143,In_1887);
and U3078 (N_3078,In_1292,In_25);
or U3079 (N_3079,In_439,In_336);
nand U3080 (N_3080,In_0,In_1688);
nor U3081 (N_3081,In_1074,In_333);
nand U3082 (N_3082,In_859,In_1461);
nor U3083 (N_3083,In_929,In_1756);
nor U3084 (N_3084,In_1863,In_372);
xor U3085 (N_3085,In_1625,In_149);
or U3086 (N_3086,In_910,In_201);
nand U3087 (N_3087,In_969,In_2219);
and U3088 (N_3088,In_2355,In_1610);
and U3089 (N_3089,In_784,In_197);
nor U3090 (N_3090,In_770,In_2358);
xor U3091 (N_3091,In_1638,In_1623);
or U3092 (N_3092,In_901,In_1745);
and U3093 (N_3093,In_2037,In_786);
and U3094 (N_3094,In_140,In_1633);
nor U3095 (N_3095,In_902,In_2171);
nor U3096 (N_3096,In_303,In_1738);
nand U3097 (N_3097,In_860,In_1178);
and U3098 (N_3098,In_333,In_135);
and U3099 (N_3099,In_1542,In_211);
and U3100 (N_3100,In_2464,In_2360);
nor U3101 (N_3101,In_455,In_320);
or U3102 (N_3102,In_602,In_1571);
or U3103 (N_3103,In_2335,In_1640);
and U3104 (N_3104,In_2305,In_1919);
nor U3105 (N_3105,In_2421,In_506);
nand U3106 (N_3106,In_1364,In_422);
or U3107 (N_3107,In_2369,In_1574);
and U3108 (N_3108,In_508,In_2301);
or U3109 (N_3109,In_1295,In_1556);
nor U3110 (N_3110,In_1602,In_2109);
nand U3111 (N_3111,In_2417,In_1813);
nand U3112 (N_3112,In_1969,In_1407);
nand U3113 (N_3113,In_348,In_2065);
and U3114 (N_3114,In_800,In_2465);
nand U3115 (N_3115,In_2456,In_2173);
and U3116 (N_3116,In_2464,In_1355);
nand U3117 (N_3117,In_445,In_306);
and U3118 (N_3118,In_132,In_1142);
nand U3119 (N_3119,In_1626,In_667);
or U3120 (N_3120,In_2428,In_591);
nor U3121 (N_3121,In_513,In_1973);
or U3122 (N_3122,In_809,In_2354);
and U3123 (N_3123,In_1979,In_882);
xor U3124 (N_3124,In_998,In_726);
and U3125 (N_3125,In_1275,In_1096);
and U3126 (N_3126,In_1331,In_2465);
or U3127 (N_3127,In_1256,In_1606);
xnor U3128 (N_3128,In_1571,In_1540);
xnor U3129 (N_3129,In_2419,In_936);
and U3130 (N_3130,In_779,In_1283);
nor U3131 (N_3131,In_2051,In_0);
and U3132 (N_3132,In_715,In_544);
xnor U3133 (N_3133,In_2479,In_664);
and U3134 (N_3134,In_99,In_1831);
xnor U3135 (N_3135,In_1308,In_2041);
nor U3136 (N_3136,In_1340,In_1948);
nor U3137 (N_3137,In_392,In_293);
nor U3138 (N_3138,In_741,In_846);
and U3139 (N_3139,In_463,In_2194);
and U3140 (N_3140,In_1416,In_2105);
nand U3141 (N_3141,In_39,In_1869);
and U3142 (N_3142,In_1967,In_187);
and U3143 (N_3143,In_2434,In_2442);
or U3144 (N_3144,In_2298,In_82);
nand U3145 (N_3145,In_1961,In_1981);
xor U3146 (N_3146,In_1861,In_2499);
nor U3147 (N_3147,In_754,In_179);
or U3148 (N_3148,In_2142,In_1566);
nand U3149 (N_3149,In_1962,In_1954);
nor U3150 (N_3150,In_840,In_903);
and U3151 (N_3151,In_68,In_2237);
xnor U3152 (N_3152,In_111,In_153);
nand U3153 (N_3153,In_438,In_1087);
or U3154 (N_3154,In_2316,In_734);
nor U3155 (N_3155,In_561,In_1204);
nand U3156 (N_3156,In_1030,In_1750);
nor U3157 (N_3157,In_2184,In_1506);
nand U3158 (N_3158,In_478,In_1221);
or U3159 (N_3159,In_1260,In_1598);
or U3160 (N_3160,In_1483,In_2200);
nor U3161 (N_3161,In_2332,In_2400);
nand U3162 (N_3162,In_478,In_1997);
nand U3163 (N_3163,In_819,In_906);
and U3164 (N_3164,In_1605,In_329);
and U3165 (N_3165,In_2186,In_1903);
and U3166 (N_3166,In_1714,In_184);
nand U3167 (N_3167,In_675,In_2087);
nor U3168 (N_3168,In_836,In_453);
nand U3169 (N_3169,In_1405,In_1145);
nor U3170 (N_3170,In_150,In_1259);
nor U3171 (N_3171,In_2128,In_866);
nand U3172 (N_3172,In_945,In_1065);
nand U3173 (N_3173,In_850,In_1039);
nand U3174 (N_3174,In_1431,In_1514);
nand U3175 (N_3175,In_1244,In_1038);
nor U3176 (N_3176,In_2230,In_608);
and U3177 (N_3177,In_193,In_138);
and U3178 (N_3178,In_2490,In_422);
and U3179 (N_3179,In_1534,In_231);
nand U3180 (N_3180,In_2075,In_129);
and U3181 (N_3181,In_656,In_928);
and U3182 (N_3182,In_690,In_1605);
nor U3183 (N_3183,In_1425,In_1865);
nand U3184 (N_3184,In_1171,In_1656);
or U3185 (N_3185,In_1961,In_790);
or U3186 (N_3186,In_313,In_1016);
or U3187 (N_3187,In_465,In_2076);
xor U3188 (N_3188,In_1679,In_1308);
nor U3189 (N_3189,In_297,In_841);
or U3190 (N_3190,In_1948,In_2464);
nand U3191 (N_3191,In_2189,In_919);
or U3192 (N_3192,In_599,In_1293);
or U3193 (N_3193,In_1338,In_1489);
nand U3194 (N_3194,In_239,In_1001);
and U3195 (N_3195,In_1268,In_2116);
or U3196 (N_3196,In_204,In_186);
xnor U3197 (N_3197,In_278,In_170);
nand U3198 (N_3198,In_1948,In_901);
and U3199 (N_3199,In_2240,In_774);
or U3200 (N_3200,In_420,In_1847);
and U3201 (N_3201,In_99,In_1859);
and U3202 (N_3202,In_2097,In_123);
or U3203 (N_3203,In_120,In_253);
and U3204 (N_3204,In_304,In_974);
nand U3205 (N_3205,In_10,In_875);
or U3206 (N_3206,In_573,In_1378);
nand U3207 (N_3207,In_2388,In_150);
nand U3208 (N_3208,In_2441,In_1643);
or U3209 (N_3209,In_2143,In_1393);
and U3210 (N_3210,In_1642,In_890);
nand U3211 (N_3211,In_2281,In_322);
nand U3212 (N_3212,In_2366,In_1727);
and U3213 (N_3213,In_2091,In_299);
or U3214 (N_3214,In_780,In_2415);
or U3215 (N_3215,In_1414,In_2247);
nor U3216 (N_3216,In_754,In_2027);
or U3217 (N_3217,In_2049,In_944);
nor U3218 (N_3218,In_2379,In_1863);
and U3219 (N_3219,In_2224,In_2419);
nor U3220 (N_3220,In_2267,In_1716);
nor U3221 (N_3221,In_1,In_2370);
nor U3222 (N_3222,In_1731,In_501);
nand U3223 (N_3223,In_144,In_1856);
and U3224 (N_3224,In_1902,In_430);
nand U3225 (N_3225,In_569,In_1572);
nor U3226 (N_3226,In_2239,In_810);
nor U3227 (N_3227,In_556,In_1305);
or U3228 (N_3228,In_1323,In_1213);
and U3229 (N_3229,In_2490,In_908);
nor U3230 (N_3230,In_2057,In_2350);
nand U3231 (N_3231,In_20,In_1959);
and U3232 (N_3232,In_1668,In_1515);
xor U3233 (N_3233,In_2288,In_1670);
and U3234 (N_3234,In_502,In_2416);
nand U3235 (N_3235,In_631,In_1744);
or U3236 (N_3236,In_2030,In_1908);
and U3237 (N_3237,In_1772,In_1589);
nor U3238 (N_3238,In_1539,In_523);
or U3239 (N_3239,In_406,In_1379);
or U3240 (N_3240,In_581,In_765);
or U3241 (N_3241,In_2300,In_1196);
nor U3242 (N_3242,In_2177,In_1795);
or U3243 (N_3243,In_288,In_1480);
nand U3244 (N_3244,In_952,In_2390);
nor U3245 (N_3245,In_769,In_454);
and U3246 (N_3246,In_1497,In_1028);
and U3247 (N_3247,In_1815,In_548);
and U3248 (N_3248,In_1956,In_912);
and U3249 (N_3249,In_623,In_2222);
nor U3250 (N_3250,In_2211,In_349);
nand U3251 (N_3251,In_877,In_1583);
nor U3252 (N_3252,In_1801,In_2013);
nor U3253 (N_3253,In_2426,In_1524);
or U3254 (N_3254,In_1383,In_1099);
and U3255 (N_3255,In_1147,In_2430);
or U3256 (N_3256,In_670,In_1154);
nand U3257 (N_3257,In_609,In_873);
or U3258 (N_3258,In_1679,In_2092);
or U3259 (N_3259,In_1573,In_971);
and U3260 (N_3260,In_1470,In_286);
or U3261 (N_3261,In_988,In_1000);
xnor U3262 (N_3262,In_1580,In_1800);
nand U3263 (N_3263,In_1260,In_1617);
nand U3264 (N_3264,In_383,In_203);
and U3265 (N_3265,In_1133,In_78);
nand U3266 (N_3266,In_2402,In_460);
and U3267 (N_3267,In_709,In_1487);
and U3268 (N_3268,In_1444,In_1155);
nor U3269 (N_3269,In_2015,In_711);
nand U3270 (N_3270,In_36,In_2153);
nand U3271 (N_3271,In_1489,In_1267);
nand U3272 (N_3272,In_1955,In_1794);
or U3273 (N_3273,In_1072,In_1688);
nand U3274 (N_3274,In_892,In_2201);
and U3275 (N_3275,In_1031,In_1773);
or U3276 (N_3276,In_374,In_925);
or U3277 (N_3277,In_2115,In_192);
and U3278 (N_3278,In_2225,In_2118);
nand U3279 (N_3279,In_454,In_2485);
or U3280 (N_3280,In_1976,In_1966);
or U3281 (N_3281,In_194,In_1761);
nor U3282 (N_3282,In_1641,In_1302);
nor U3283 (N_3283,In_1706,In_1251);
nor U3284 (N_3284,In_1545,In_1429);
and U3285 (N_3285,In_353,In_1952);
nor U3286 (N_3286,In_885,In_344);
and U3287 (N_3287,In_556,In_61);
or U3288 (N_3288,In_560,In_1165);
nor U3289 (N_3289,In_494,In_1036);
nor U3290 (N_3290,In_2242,In_1788);
and U3291 (N_3291,In_838,In_2337);
nand U3292 (N_3292,In_186,In_1205);
nor U3293 (N_3293,In_556,In_251);
nand U3294 (N_3294,In_917,In_2483);
nor U3295 (N_3295,In_723,In_233);
nand U3296 (N_3296,In_184,In_1620);
or U3297 (N_3297,In_2322,In_2219);
and U3298 (N_3298,In_950,In_570);
and U3299 (N_3299,In_662,In_2428);
and U3300 (N_3300,In_1008,In_694);
or U3301 (N_3301,In_197,In_1300);
nand U3302 (N_3302,In_655,In_1672);
nand U3303 (N_3303,In_1945,In_2024);
nand U3304 (N_3304,In_886,In_1499);
nor U3305 (N_3305,In_265,In_2413);
nor U3306 (N_3306,In_1958,In_2443);
and U3307 (N_3307,In_2282,In_2417);
or U3308 (N_3308,In_2485,In_299);
and U3309 (N_3309,In_915,In_1002);
nand U3310 (N_3310,In_710,In_2020);
nand U3311 (N_3311,In_1931,In_1176);
nand U3312 (N_3312,In_736,In_957);
nor U3313 (N_3313,In_2042,In_171);
or U3314 (N_3314,In_50,In_2073);
nand U3315 (N_3315,In_99,In_404);
or U3316 (N_3316,In_515,In_2320);
or U3317 (N_3317,In_1053,In_606);
and U3318 (N_3318,In_1527,In_1041);
and U3319 (N_3319,In_276,In_333);
nand U3320 (N_3320,In_943,In_1221);
nand U3321 (N_3321,In_199,In_397);
nor U3322 (N_3322,In_381,In_1002);
and U3323 (N_3323,In_2181,In_983);
nand U3324 (N_3324,In_312,In_2256);
nand U3325 (N_3325,In_1624,In_2301);
or U3326 (N_3326,In_381,In_1628);
or U3327 (N_3327,In_1233,In_1853);
nor U3328 (N_3328,In_602,In_1194);
nor U3329 (N_3329,In_1220,In_1447);
or U3330 (N_3330,In_791,In_1861);
or U3331 (N_3331,In_1198,In_1353);
or U3332 (N_3332,In_1879,In_121);
or U3333 (N_3333,In_596,In_1560);
or U3334 (N_3334,In_1764,In_524);
nor U3335 (N_3335,In_2407,In_1049);
nor U3336 (N_3336,In_459,In_668);
nor U3337 (N_3337,In_360,In_2438);
or U3338 (N_3338,In_1676,In_1855);
nor U3339 (N_3339,In_336,In_246);
and U3340 (N_3340,In_885,In_1476);
nor U3341 (N_3341,In_1681,In_582);
and U3342 (N_3342,In_735,In_644);
or U3343 (N_3343,In_1402,In_906);
or U3344 (N_3344,In_2231,In_647);
or U3345 (N_3345,In_2191,In_1459);
and U3346 (N_3346,In_1369,In_440);
or U3347 (N_3347,In_2113,In_125);
nand U3348 (N_3348,In_79,In_2188);
nor U3349 (N_3349,In_434,In_2250);
or U3350 (N_3350,In_1219,In_91);
nor U3351 (N_3351,In_486,In_805);
or U3352 (N_3352,In_28,In_2002);
and U3353 (N_3353,In_1858,In_415);
or U3354 (N_3354,In_2494,In_816);
nor U3355 (N_3355,In_1701,In_208);
or U3356 (N_3356,In_1071,In_279);
nand U3357 (N_3357,In_492,In_2281);
or U3358 (N_3358,In_1642,In_999);
and U3359 (N_3359,In_826,In_357);
or U3360 (N_3360,In_1374,In_691);
or U3361 (N_3361,In_1346,In_1402);
nor U3362 (N_3362,In_1170,In_2071);
nor U3363 (N_3363,In_2105,In_301);
nand U3364 (N_3364,In_296,In_559);
or U3365 (N_3365,In_2223,In_2390);
and U3366 (N_3366,In_395,In_2484);
nor U3367 (N_3367,In_309,In_34);
nand U3368 (N_3368,In_45,In_356);
and U3369 (N_3369,In_2359,In_1412);
and U3370 (N_3370,In_1749,In_1017);
or U3371 (N_3371,In_1176,In_1591);
nor U3372 (N_3372,In_1385,In_1517);
and U3373 (N_3373,In_239,In_1011);
and U3374 (N_3374,In_311,In_2310);
nand U3375 (N_3375,In_2173,In_1295);
and U3376 (N_3376,In_1257,In_2209);
or U3377 (N_3377,In_1608,In_379);
nand U3378 (N_3378,In_1078,In_250);
and U3379 (N_3379,In_1225,In_2389);
nand U3380 (N_3380,In_2122,In_50);
and U3381 (N_3381,In_726,In_917);
nor U3382 (N_3382,In_106,In_937);
xnor U3383 (N_3383,In_2393,In_2230);
nand U3384 (N_3384,In_1035,In_1403);
nor U3385 (N_3385,In_1223,In_2017);
nand U3386 (N_3386,In_1770,In_1898);
or U3387 (N_3387,In_2028,In_1081);
nand U3388 (N_3388,In_2144,In_521);
nand U3389 (N_3389,In_2420,In_1417);
or U3390 (N_3390,In_2324,In_2441);
xnor U3391 (N_3391,In_858,In_272);
xor U3392 (N_3392,In_1267,In_1472);
xor U3393 (N_3393,In_1412,In_2408);
or U3394 (N_3394,In_1823,In_1652);
nand U3395 (N_3395,In_1321,In_1817);
nor U3396 (N_3396,In_230,In_960);
nor U3397 (N_3397,In_2136,In_519);
nor U3398 (N_3398,In_2056,In_2173);
or U3399 (N_3399,In_47,In_2305);
nor U3400 (N_3400,In_1685,In_788);
nand U3401 (N_3401,In_2295,In_609);
and U3402 (N_3402,In_2091,In_1757);
nor U3403 (N_3403,In_210,In_458);
or U3404 (N_3404,In_369,In_1060);
nand U3405 (N_3405,In_2123,In_378);
or U3406 (N_3406,In_1395,In_2405);
nor U3407 (N_3407,In_1328,In_923);
or U3408 (N_3408,In_76,In_2172);
or U3409 (N_3409,In_208,In_2308);
and U3410 (N_3410,In_240,In_1025);
nor U3411 (N_3411,In_296,In_1207);
nor U3412 (N_3412,In_168,In_767);
nand U3413 (N_3413,In_2241,In_632);
or U3414 (N_3414,In_1886,In_2003);
and U3415 (N_3415,In_352,In_860);
nand U3416 (N_3416,In_2290,In_394);
or U3417 (N_3417,In_2299,In_1477);
or U3418 (N_3418,In_688,In_1311);
and U3419 (N_3419,In_1085,In_2301);
or U3420 (N_3420,In_998,In_928);
xnor U3421 (N_3421,In_2214,In_2318);
or U3422 (N_3422,In_614,In_1881);
nand U3423 (N_3423,In_385,In_2385);
or U3424 (N_3424,In_1035,In_2480);
and U3425 (N_3425,In_331,In_2099);
nor U3426 (N_3426,In_931,In_255);
nand U3427 (N_3427,In_2118,In_2228);
nor U3428 (N_3428,In_14,In_795);
or U3429 (N_3429,In_357,In_562);
or U3430 (N_3430,In_591,In_487);
nand U3431 (N_3431,In_962,In_491);
nand U3432 (N_3432,In_1114,In_696);
and U3433 (N_3433,In_2040,In_2005);
nor U3434 (N_3434,In_671,In_340);
nand U3435 (N_3435,In_698,In_1906);
nand U3436 (N_3436,In_855,In_648);
nor U3437 (N_3437,In_588,In_1271);
or U3438 (N_3438,In_1493,In_140);
nor U3439 (N_3439,In_139,In_1636);
and U3440 (N_3440,In_1643,In_1730);
nand U3441 (N_3441,In_1823,In_573);
nor U3442 (N_3442,In_1892,In_1056);
or U3443 (N_3443,In_1579,In_1187);
nand U3444 (N_3444,In_807,In_894);
nor U3445 (N_3445,In_120,In_2077);
and U3446 (N_3446,In_1994,In_1946);
nor U3447 (N_3447,In_1472,In_249);
or U3448 (N_3448,In_2193,In_1025);
or U3449 (N_3449,In_1199,In_1613);
nand U3450 (N_3450,In_1937,In_1704);
xnor U3451 (N_3451,In_1962,In_743);
nand U3452 (N_3452,In_921,In_1746);
and U3453 (N_3453,In_106,In_1178);
xor U3454 (N_3454,In_1639,In_149);
and U3455 (N_3455,In_1459,In_1449);
nand U3456 (N_3456,In_450,In_129);
nand U3457 (N_3457,In_430,In_638);
nor U3458 (N_3458,In_2254,In_1243);
nor U3459 (N_3459,In_1353,In_661);
or U3460 (N_3460,In_1646,In_2197);
or U3461 (N_3461,In_701,In_82);
nand U3462 (N_3462,In_1063,In_1065);
and U3463 (N_3463,In_1595,In_805);
nand U3464 (N_3464,In_1961,In_1971);
nand U3465 (N_3465,In_1050,In_748);
nor U3466 (N_3466,In_85,In_1604);
nand U3467 (N_3467,In_2228,In_832);
nor U3468 (N_3468,In_1831,In_2052);
and U3469 (N_3469,In_2094,In_576);
nor U3470 (N_3470,In_2039,In_985);
or U3471 (N_3471,In_1159,In_1320);
or U3472 (N_3472,In_1397,In_2237);
and U3473 (N_3473,In_1884,In_8);
and U3474 (N_3474,In_727,In_1391);
or U3475 (N_3475,In_421,In_2368);
nor U3476 (N_3476,In_1416,In_2341);
nor U3477 (N_3477,In_2164,In_429);
or U3478 (N_3478,In_125,In_1529);
nand U3479 (N_3479,In_95,In_1552);
nand U3480 (N_3480,In_1530,In_351);
or U3481 (N_3481,In_947,In_1581);
or U3482 (N_3482,In_607,In_2389);
and U3483 (N_3483,In_978,In_1948);
nor U3484 (N_3484,In_1700,In_1838);
or U3485 (N_3485,In_26,In_167);
or U3486 (N_3486,In_1182,In_1896);
nor U3487 (N_3487,In_727,In_64);
and U3488 (N_3488,In_1689,In_1943);
nor U3489 (N_3489,In_1850,In_1310);
nand U3490 (N_3490,In_2051,In_1284);
nand U3491 (N_3491,In_1549,In_2343);
nor U3492 (N_3492,In_1510,In_304);
and U3493 (N_3493,In_1163,In_2254);
nand U3494 (N_3494,In_2124,In_1128);
or U3495 (N_3495,In_606,In_1513);
nor U3496 (N_3496,In_163,In_71);
or U3497 (N_3497,In_437,In_156);
nand U3498 (N_3498,In_240,In_37);
nand U3499 (N_3499,In_700,In_1453);
or U3500 (N_3500,In_1505,In_794);
xnor U3501 (N_3501,In_775,In_2267);
and U3502 (N_3502,In_534,In_1471);
and U3503 (N_3503,In_457,In_154);
nand U3504 (N_3504,In_85,In_1779);
or U3505 (N_3505,In_739,In_196);
nor U3506 (N_3506,In_178,In_261);
and U3507 (N_3507,In_914,In_1324);
nand U3508 (N_3508,In_1633,In_1191);
and U3509 (N_3509,In_2075,In_1000);
or U3510 (N_3510,In_1486,In_2169);
nand U3511 (N_3511,In_1329,In_1832);
nor U3512 (N_3512,In_468,In_615);
and U3513 (N_3513,In_732,In_353);
and U3514 (N_3514,In_1097,In_2204);
or U3515 (N_3515,In_1133,In_1483);
nor U3516 (N_3516,In_1251,In_470);
nand U3517 (N_3517,In_2476,In_1421);
nor U3518 (N_3518,In_98,In_436);
or U3519 (N_3519,In_1097,In_46);
and U3520 (N_3520,In_1556,In_294);
nor U3521 (N_3521,In_1272,In_694);
xnor U3522 (N_3522,In_781,In_596);
nand U3523 (N_3523,In_1392,In_711);
nor U3524 (N_3524,In_610,In_2057);
and U3525 (N_3525,In_1131,In_941);
or U3526 (N_3526,In_909,In_1077);
or U3527 (N_3527,In_1185,In_1126);
and U3528 (N_3528,In_2222,In_116);
nand U3529 (N_3529,In_1625,In_1850);
and U3530 (N_3530,In_303,In_1475);
or U3531 (N_3531,In_741,In_4);
nand U3532 (N_3532,In_118,In_2424);
nor U3533 (N_3533,In_1399,In_1428);
nand U3534 (N_3534,In_74,In_204);
nor U3535 (N_3535,In_1339,In_1337);
or U3536 (N_3536,In_1753,In_1090);
nor U3537 (N_3537,In_482,In_1231);
and U3538 (N_3538,In_2235,In_1540);
nand U3539 (N_3539,In_987,In_506);
or U3540 (N_3540,In_2380,In_1083);
and U3541 (N_3541,In_431,In_2413);
nand U3542 (N_3542,In_1104,In_1457);
nor U3543 (N_3543,In_541,In_2092);
nand U3544 (N_3544,In_1921,In_859);
xnor U3545 (N_3545,In_1707,In_1191);
nor U3546 (N_3546,In_2454,In_1475);
nand U3547 (N_3547,In_747,In_1078);
and U3548 (N_3548,In_2300,In_2411);
nor U3549 (N_3549,In_666,In_1453);
nand U3550 (N_3550,In_1850,In_1972);
and U3551 (N_3551,In_871,In_1220);
or U3552 (N_3552,In_837,In_1619);
xor U3553 (N_3553,In_727,In_96);
nand U3554 (N_3554,In_2113,In_1763);
nand U3555 (N_3555,In_2312,In_114);
or U3556 (N_3556,In_1968,In_1024);
or U3557 (N_3557,In_465,In_112);
nor U3558 (N_3558,In_43,In_1403);
nor U3559 (N_3559,In_2306,In_2088);
nand U3560 (N_3560,In_859,In_1293);
nor U3561 (N_3561,In_2232,In_1761);
or U3562 (N_3562,In_1968,In_58);
or U3563 (N_3563,In_430,In_2314);
nor U3564 (N_3564,In_1849,In_53);
and U3565 (N_3565,In_442,In_1792);
or U3566 (N_3566,In_438,In_1392);
and U3567 (N_3567,In_2127,In_1615);
or U3568 (N_3568,In_226,In_1279);
nor U3569 (N_3569,In_779,In_1485);
nand U3570 (N_3570,In_163,In_2433);
nor U3571 (N_3571,In_922,In_983);
nand U3572 (N_3572,In_716,In_1301);
or U3573 (N_3573,In_1822,In_1699);
nor U3574 (N_3574,In_2298,In_422);
xnor U3575 (N_3575,In_1678,In_1217);
xor U3576 (N_3576,In_949,In_1489);
or U3577 (N_3577,In_2112,In_2070);
or U3578 (N_3578,In_2253,In_1117);
nor U3579 (N_3579,In_1281,In_871);
nor U3580 (N_3580,In_56,In_2419);
or U3581 (N_3581,In_2151,In_1431);
nor U3582 (N_3582,In_32,In_818);
nand U3583 (N_3583,In_450,In_1721);
and U3584 (N_3584,In_2175,In_1392);
nor U3585 (N_3585,In_597,In_982);
xor U3586 (N_3586,In_442,In_1003);
and U3587 (N_3587,In_206,In_1638);
nor U3588 (N_3588,In_367,In_1807);
and U3589 (N_3589,In_1158,In_1844);
and U3590 (N_3590,In_1478,In_1115);
or U3591 (N_3591,In_2489,In_463);
or U3592 (N_3592,In_2058,In_166);
or U3593 (N_3593,In_1382,In_2351);
or U3594 (N_3594,In_24,In_1555);
nor U3595 (N_3595,In_2081,In_630);
or U3596 (N_3596,In_91,In_2130);
and U3597 (N_3597,In_1694,In_346);
nor U3598 (N_3598,In_2446,In_329);
or U3599 (N_3599,In_107,In_2442);
nand U3600 (N_3600,In_326,In_1911);
nor U3601 (N_3601,In_863,In_980);
nand U3602 (N_3602,In_2144,In_2246);
nand U3603 (N_3603,In_417,In_1999);
or U3604 (N_3604,In_468,In_2006);
nor U3605 (N_3605,In_308,In_25);
nand U3606 (N_3606,In_1396,In_877);
nand U3607 (N_3607,In_229,In_877);
or U3608 (N_3608,In_245,In_281);
or U3609 (N_3609,In_147,In_858);
nand U3610 (N_3610,In_479,In_2409);
nor U3611 (N_3611,In_1228,In_1096);
nand U3612 (N_3612,In_879,In_2178);
or U3613 (N_3613,In_1386,In_522);
or U3614 (N_3614,In_608,In_1535);
and U3615 (N_3615,In_532,In_505);
or U3616 (N_3616,In_1501,In_1419);
and U3617 (N_3617,In_2324,In_1073);
nand U3618 (N_3618,In_1752,In_2076);
nor U3619 (N_3619,In_231,In_858);
nand U3620 (N_3620,In_1995,In_990);
or U3621 (N_3621,In_1947,In_1513);
nor U3622 (N_3622,In_2013,In_662);
or U3623 (N_3623,In_372,In_2356);
and U3624 (N_3624,In_1010,In_742);
nand U3625 (N_3625,In_110,In_2492);
nor U3626 (N_3626,In_773,In_460);
and U3627 (N_3627,In_958,In_1053);
nand U3628 (N_3628,In_931,In_595);
xor U3629 (N_3629,In_38,In_125);
xnor U3630 (N_3630,In_314,In_1805);
nor U3631 (N_3631,In_516,In_128);
nand U3632 (N_3632,In_1394,In_317);
and U3633 (N_3633,In_704,In_1045);
xor U3634 (N_3634,In_1064,In_1643);
or U3635 (N_3635,In_1428,In_1644);
and U3636 (N_3636,In_145,In_2102);
nor U3637 (N_3637,In_1994,In_1126);
nand U3638 (N_3638,In_1517,In_235);
and U3639 (N_3639,In_379,In_2030);
and U3640 (N_3640,In_1774,In_945);
and U3641 (N_3641,In_1521,In_1128);
nor U3642 (N_3642,In_1408,In_1102);
nand U3643 (N_3643,In_67,In_106);
nand U3644 (N_3644,In_277,In_17);
and U3645 (N_3645,In_782,In_528);
or U3646 (N_3646,In_175,In_1100);
nand U3647 (N_3647,In_1093,In_1048);
and U3648 (N_3648,In_1733,In_2277);
nand U3649 (N_3649,In_391,In_2132);
nand U3650 (N_3650,In_1618,In_2301);
nor U3651 (N_3651,In_1123,In_1158);
or U3652 (N_3652,In_1510,In_547);
and U3653 (N_3653,In_1608,In_1742);
and U3654 (N_3654,In_467,In_2221);
or U3655 (N_3655,In_480,In_246);
nand U3656 (N_3656,In_788,In_1130);
xor U3657 (N_3657,In_895,In_1283);
and U3658 (N_3658,In_578,In_608);
or U3659 (N_3659,In_1303,In_671);
and U3660 (N_3660,In_950,In_2012);
or U3661 (N_3661,In_1497,In_2433);
and U3662 (N_3662,In_610,In_1223);
or U3663 (N_3663,In_1057,In_1516);
nor U3664 (N_3664,In_1867,In_1457);
and U3665 (N_3665,In_53,In_1411);
nand U3666 (N_3666,In_1582,In_425);
nand U3667 (N_3667,In_1402,In_320);
and U3668 (N_3668,In_2372,In_318);
or U3669 (N_3669,In_1870,In_1864);
or U3670 (N_3670,In_1894,In_1020);
or U3671 (N_3671,In_1010,In_328);
and U3672 (N_3672,In_1272,In_1933);
nand U3673 (N_3673,In_1072,In_1543);
or U3674 (N_3674,In_2339,In_1485);
nor U3675 (N_3675,In_2130,In_2091);
or U3676 (N_3676,In_1344,In_1825);
and U3677 (N_3677,In_172,In_2316);
nor U3678 (N_3678,In_491,In_1787);
nor U3679 (N_3679,In_1170,In_2068);
nand U3680 (N_3680,In_692,In_1715);
nor U3681 (N_3681,In_1017,In_566);
nand U3682 (N_3682,In_2016,In_410);
and U3683 (N_3683,In_2437,In_1788);
nand U3684 (N_3684,In_1869,In_1896);
or U3685 (N_3685,In_2402,In_1439);
or U3686 (N_3686,In_1753,In_460);
and U3687 (N_3687,In_2259,In_483);
and U3688 (N_3688,In_2003,In_1367);
nand U3689 (N_3689,In_425,In_1053);
xnor U3690 (N_3690,In_1184,In_560);
or U3691 (N_3691,In_1901,In_948);
nand U3692 (N_3692,In_738,In_2370);
and U3693 (N_3693,In_268,In_1247);
nand U3694 (N_3694,In_837,In_764);
and U3695 (N_3695,In_2138,In_619);
or U3696 (N_3696,In_897,In_1043);
and U3697 (N_3697,In_667,In_854);
nor U3698 (N_3698,In_27,In_182);
nor U3699 (N_3699,In_1430,In_68);
or U3700 (N_3700,In_109,In_771);
and U3701 (N_3701,In_160,In_920);
and U3702 (N_3702,In_753,In_765);
or U3703 (N_3703,In_328,In_109);
nor U3704 (N_3704,In_491,In_2497);
nor U3705 (N_3705,In_73,In_2253);
nand U3706 (N_3706,In_1351,In_2353);
and U3707 (N_3707,In_1420,In_1574);
nor U3708 (N_3708,In_2227,In_814);
nor U3709 (N_3709,In_2313,In_431);
or U3710 (N_3710,In_1254,In_1777);
or U3711 (N_3711,In_953,In_1597);
nor U3712 (N_3712,In_1982,In_1738);
and U3713 (N_3713,In_655,In_1722);
or U3714 (N_3714,In_977,In_630);
nor U3715 (N_3715,In_2495,In_1234);
nand U3716 (N_3716,In_1462,In_1811);
and U3717 (N_3717,In_2412,In_936);
nand U3718 (N_3718,In_1596,In_1552);
nand U3719 (N_3719,In_2340,In_2302);
nand U3720 (N_3720,In_1749,In_16);
or U3721 (N_3721,In_438,In_2276);
or U3722 (N_3722,In_340,In_216);
nand U3723 (N_3723,In_2411,In_2297);
or U3724 (N_3724,In_330,In_1537);
and U3725 (N_3725,In_168,In_1875);
and U3726 (N_3726,In_1182,In_1492);
or U3727 (N_3727,In_166,In_959);
nand U3728 (N_3728,In_778,In_1848);
or U3729 (N_3729,In_350,In_1288);
or U3730 (N_3730,In_945,In_475);
or U3731 (N_3731,In_122,In_646);
and U3732 (N_3732,In_1747,In_246);
nor U3733 (N_3733,In_1612,In_1750);
xnor U3734 (N_3734,In_2226,In_1775);
nand U3735 (N_3735,In_2167,In_622);
nand U3736 (N_3736,In_296,In_2091);
nand U3737 (N_3737,In_1991,In_1524);
nand U3738 (N_3738,In_1282,In_964);
and U3739 (N_3739,In_1435,In_560);
and U3740 (N_3740,In_1848,In_2042);
or U3741 (N_3741,In_1324,In_2182);
or U3742 (N_3742,In_2492,In_2067);
nand U3743 (N_3743,In_358,In_231);
and U3744 (N_3744,In_744,In_2042);
or U3745 (N_3745,In_2479,In_364);
or U3746 (N_3746,In_473,In_418);
or U3747 (N_3747,In_976,In_1267);
and U3748 (N_3748,In_2420,In_884);
and U3749 (N_3749,In_128,In_2032);
and U3750 (N_3750,In_843,In_359);
or U3751 (N_3751,In_548,In_797);
nand U3752 (N_3752,In_869,In_241);
or U3753 (N_3753,In_1024,In_713);
or U3754 (N_3754,In_2421,In_1193);
nor U3755 (N_3755,In_1438,In_1208);
and U3756 (N_3756,In_626,In_744);
and U3757 (N_3757,In_1886,In_1687);
or U3758 (N_3758,In_286,In_799);
and U3759 (N_3759,In_2277,In_362);
nor U3760 (N_3760,In_1384,In_516);
or U3761 (N_3761,In_2427,In_1053);
nand U3762 (N_3762,In_390,In_2462);
nor U3763 (N_3763,In_2162,In_2210);
and U3764 (N_3764,In_2007,In_2421);
nor U3765 (N_3765,In_1213,In_608);
nor U3766 (N_3766,In_1463,In_1031);
or U3767 (N_3767,In_2054,In_1884);
nand U3768 (N_3768,In_674,In_1686);
or U3769 (N_3769,In_94,In_2211);
nand U3770 (N_3770,In_178,In_1731);
nand U3771 (N_3771,In_1349,In_1750);
or U3772 (N_3772,In_1530,In_498);
or U3773 (N_3773,In_2486,In_518);
nand U3774 (N_3774,In_2161,In_1027);
or U3775 (N_3775,In_214,In_1681);
nor U3776 (N_3776,In_813,In_119);
and U3777 (N_3777,In_1614,In_716);
nand U3778 (N_3778,In_898,In_2191);
or U3779 (N_3779,In_2325,In_1179);
nand U3780 (N_3780,In_146,In_2471);
nor U3781 (N_3781,In_2075,In_2436);
and U3782 (N_3782,In_2406,In_2239);
or U3783 (N_3783,In_125,In_89);
nor U3784 (N_3784,In_458,In_1294);
nand U3785 (N_3785,In_712,In_808);
nand U3786 (N_3786,In_888,In_1329);
or U3787 (N_3787,In_24,In_1818);
or U3788 (N_3788,In_839,In_2296);
or U3789 (N_3789,In_184,In_265);
nor U3790 (N_3790,In_917,In_115);
nor U3791 (N_3791,In_700,In_1502);
and U3792 (N_3792,In_1063,In_173);
nand U3793 (N_3793,In_215,In_1907);
nand U3794 (N_3794,In_1541,In_1176);
nor U3795 (N_3795,In_1393,In_1559);
nand U3796 (N_3796,In_1252,In_1277);
nor U3797 (N_3797,In_625,In_1875);
nand U3798 (N_3798,In_605,In_1752);
and U3799 (N_3799,In_1341,In_315);
and U3800 (N_3800,In_1463,In_1805);
or U3801 (N_3801,In_1580,In_516);
and U3802 (N_3802,In_867,In_1226);
nor U3803 (N_3803,In_552,In_2291);
or U3804 (N_3804,In_1051,In_1990);
and U3805 (N_3805,In_1191,In_966);
and U3806 (N_3806,In_2139,In_2029);
nor U3807 (N_3807,In_2269,In_960);
nand U3808 (N_3808,In_1979,In_1440);
or U3809 (N_3809,In_2463,In_2287);
nand U3810 (N_3810,In_2090,In_2116);
and U3811 (N_3811,In_1618,In_990);
nor U3812 (N_3812,In_2344,In_34);
and U3813 (N_3813,In_1057,In_566);
nor U3814 (N_3814,In_1635,In_817);
nand U3815 (N_3815,In_1649,In_783);
nor U3816 (N_3816,In_1861,In_354);
and U3817 (N_3817,In_1180,In_1082);
nand U3818 (N_3818,In_212,In_574);
and U3819 (N_3819,In_1492,In_1293);
nand U3820 (N_3820,In_271,In_431);
nand U3821 (N_3821,In_320,In_1015);
nor U3822 (N_3822,In_1344,In_1105);
nand U3823 (N_3823,In_2045,In_1026);
nand U3824 (N_3824,In_1399,In_239);
or U3825 (N_3825,In_1867,In_2154);
nand U3826 (N_3826,In_2105,In_1477);
nand U3827 (N_3827,In_802,In_629);
nand U3828 (N_3828,In_962,In_1670);
nor U3829 (N_3829,In_1142,In_145);
xor U3830 (N_3830,In_1439,In_1649);
nand U3831 (N_3831,In_835,In_2343);
nor U3832 (N_3832,In_2305,In_204);
nand U3833 (N_3833,In_262,In_2315);
or U3834 (N_3834,In_53,In_367);
nand U3835 (N_3835,In_77,In_204);
or U3836 (N_3836,In_1239,In_2046);
nand U3837 (N_3837,In_579,In_756);
or U3838 (N_3838,In_1504,In_191);
or U3839 (N_3839,In_2100,In_1856);
nand U3840 (N_3840,In_2385,In_166);
nand U3841 (N_3841,In_1904,In_617);
or U3842 (N_3842,In_1969,In_1968);
or U3843 (N_3843,In_90,In_1443);
xor U3844 (N_3844,In_1499,In_694);
nor U3845 (N_3845,In_1869,In_419);
and U3846 (N_3846,In_554,In_123);
nand U3847 (N_3847,In_560,In_2180);
nand U3848 (N_3848,In_2021,In_1796);
nor U3849 (N_3849,In_2022,In_430);
or U3850 (N_3850,In_821,In_1944);
nor U3851 (N_3851,In_2426,In_2153);
nor U3852 (N_3852,In_682,In_1564);
nor U3853 (N_3853,In_898,In_1699);
nand U3854 (N_3854,In_839,In_1343);
and U3855 (N_3855,In_1747,In_2109);
nand U3856 (N_3856,In_1759,In_580);
and U3857 (N_3857,In_1432,In_1612);
nand U3858 (N_3858,In_682,In_1151);
or U3859 (N_3859,In_1323,In_932);
nor U3860 (N_3860,In_1754,In_2339);
or U3861 (N_3861,In_1913,In_2314);
or U3862 (N_3862,In_1795,In_554);
or U3863 (N_3863,In_2119,In_1500);
and U3864 (N_3864,In_1616,In_1498);
nand U3865 (N_3865,In_1279,In_2481);
or U3866 (N_3866,In_878,In_818);
or U3867 (N_3867,In_858,In_2205);
and U3868 (N_3868,In_2120,In_1938);
nand U3869 (N_3869,In_137,In_920);
and U3870 (N_3870,In_1405,In_436);
nand U3871 (N_3871,In_822,In_1151);
nand U3872 (N_3872,In_554,In_2186);
or U3873 (N_3873,In_1143,In_2307);
or U3874 (N_3874,In_1711,In_653);
nor U3875 (N_3875,In_214,In_84);
and U3876 (N_3876,In_1447,In_2276);
and U3877 (N_3877,In_1376,In_2296);
or U3878 (N_3878,In_2478,In_410);
and U3879 (N_3879,In_784,In_2392);
nor U3880 (N_3880,In_438,In_591);
nor U3881 (N_3881,In_247,In_1523);
and U3882 (N_3882,In_2028,In_779);
and U3883 (N_3883,In_201,In_438);
and U3884 (N_3884,In_2257,In_1501);
and U3885 (N_3885,In_166,In_105);
nand U3886 (N_3886,In_817,In_1703);
nor U3887 (N_3887,In_1208,In_1849);
and U3888 (N_3888,In_1281,In_2163);
nor U3889 (N_3889,In_1614,In_1203);
nand U3890 (N_3890,In_1947,In_2316);
nand U3891 (N_3891,In_2451,In_1051);
nand U3892 (N_3892,In_426,In_1804);
xnor U3893 (N_3893,In_1854,In_1908);
or U3894 (N_3894,In_1858,In_502);
and U3895 (N_3895,In_2137,In_2256);
or U3896 (N_3896,In_1047,In_370);
and U3897 (N_3897,In_1055,In_1947);
nand U3898 (N_3898,In_719,In_2438);
nand U3899 (N_3899,In_1692,In_1508);
nand U3900 (N_3900,In_28,In_2365);
xnor U3901 (N_3901,In_1898,In_2137);
nor U3902 (N_3902,In_881,In_1940);
nand U3903 (N_3903,In_2289,In_2403);
or U3904 (N_3904,In_107,In_462);
or U3905 (N_3905,In_2277,In_2021);
nand U3906 (N_3906,In_488,In_670);
and U3907 (N_3907,In_892,In_2412);
nand U3908 (N_3908,In_1838,In_2013);
and U3909 (N_3909,In_406,In_2183);
nand U3910 (N_3910,In_2092,In_1791);
or U3911 (N_3911,In_2273,In_653);
or U3912 (N_3912,In_2370,In_451);
or U3913 (N_3913,In_715,In_187);
and U3914 (N_3914,In_1069,In_2309);
nand U3915 (N_3915,In_2150,In_2118);
nor U3916 (N_3916,In_1481,In_279);
nor U3917 (N_3917,In_391,In_427);
nor U3918 (N_3918,In_2458,In_2031);
nand U3919 (N_3919,In_1475,In_853);
and U3920 (N_3920,In_1954,In_2131);
nor U3921 (N_3921,In_65,In_282);
or U3922 (N_3922,In_1782,In_2451);
nand U3923 (N_3923,In_1705,In_445);
and U3924 (N_3924,In_1987,In_1464);
nand U3925 (N_3925,In_1196,In_743);
and U3926 (N_3926,In_776,In_491);
nand U3927 (N_3927,In_1310,In_655);
nor U3928 (N_3928,In_1181,In_435);
nor U3929 (N_3929,In_2241,In_2329);
nand U3930 (N_3930,In_2001,In_2442);
or U3931 (N_3931,In_1578,In_526);
or U3932 (N_3932,In_1814,In_2167);
nand U3933 (N_3933,In_1950,In_1356);
nor U3934 (N_3934,In_2408,In_368);
or U3935 (N_3935,In_2361,In_258);
nor U3936 (N_3936,In_661,In_492);
nor U3937 (N_3937,In_1156,In_2056);
nor U3938 (N_3938,In_2085,In_687);
or U3939 (N_3939,In_2448,In_263);
nor U3940 (N_3940,In_140,In_278);
or U3941 (N_3941,In_1874,In_1580);
or U3942 (N_3942,In_801,In_1428);
nor U3943 (N_3943,In_1960,In_201);
nor U3944 (N_3944,In_251,In_1932);
or U3945 (N_3945,In_740,In_1761);
nor U3946 (N_3946,In_1419,In_840);
nand U3947 (N_3947,In_1909,In_2243);
nor U3948 (N_3948,In_749,In_2080);
nor U3949 (N_3949,In_1666,In_2117);
or U3950 (N_3950,In_2276,In_2017);
nor U3951 (N_3951,In_1977,In_1773);
xnor U3952 (N_3952,In_2014,In_514);
and U3953 (N_3953,In_1064,In_2159);
nand U3954 (N_3954,In_2274,In_758);
and U3955 (N_3955,In_1934,In_2055);
nand U3956 (N_3956,In_1757,In_164);
or U3957 (N_3957,In_3,In_771);
xor U3958 (N_3958,In_2259,In_2200);
nor U3959 (N_3959,In_830,In_375);
or U3960 (N_3960,In_2296,In_1416);
nand U3961 (N_3961,In_578,In_512);
nor U3962 (N_3962,In_527,In_1174);
or U3963 (N_3963,In_2336,In_2011);
or U3964 (N_3964,In_1553,In_1307);
nor U3965 (N_3965,In_851,In_821);
nor U3966 (N_3966,In_90,In_1586);
nand U3967 (N_3967,In_1450,In_986);
nor U3968 (N_3968,In_862,In_541);
or U3969 (N_3969,In_25,In_987);
nand U3970 (N_3970,In_1642,In_58);
xor U3971 (N_3971,In_939,In_1444);
and U3972 (N_3972,In_615,In_1726);
nor U3973 (N_3973,In_2019,In_2315);
xor U3974 (N_3974,In_248,In_867);
or U3975 (N_3975,In_2327,In_1477);
nor U3976 (N_3976,In_48,In_2155);
or U3977 (N_3977,In_562,In_1268);
nor U3978 (N_3978,In_1535,In_2410);
nand U3979 (N_3979,In_1487,In_721);
nor U3980 (N_3980,In_2004,In_1775);
nand U3981 (N_3981,In_2287,In_1112);
or U3982 (N_3982,In_1674,In_1032);
nand U3983 (N_3983,In_1449,In_851);
nor U3984 (N_3984,In_1635,In_1576);
nand U3985 (N_3985,In_875,In_95);
nor U3986 (N_3986,In_25,In_1641);
nor U3987 (N_3987,In_809,In_904);
nand U3988 (N_3988,In_2034,In_1905);
nor U3989 (N_3989,In_105,In_1218);
or U3990 (N_3990,In_1379,In_2313);
nor U3991 (N_3991,In_2445,In_637);
or U3992 (N_3992,In_2185,In_1763);
nor U3993 (N_3993,In_626,In_2492);
or U3994 (N_3994,In_749,In_1920);
and U3995 (N_3995,In_1339,In_1969);
or U3996 (N_3996,In_981,In_1415);
xnor U3997 (N_3997,In_1112,In_1071);
or U3998 (N_3998,In_696,In_2233);
and U3999 (N_3999,In_316,In_1668);
and U4000 (N_4000,In_1936,In_591);
nand U4001 (N_4001,In_706,In_2321);
nand U4002 (N_4002,In_972,In_2001);
nand U4003 (N_4003,In_1228,In_999);
nor U4004 (N_4004,In_37,In_1337);
nand U4005 (N_4005,In_2041,In_816);
and U4006 (N_4006,In_2247,In_2052);
nor U4007 (N_4007,In_934,In_1703);
nand U4008 (N_4008,In_2255,In_2154);
or U4009 (N_4009,In_2454,In_1163);
or U4010 (N_4010,In_1939,In_1732);
and U4011 (N_4011,In_713,In_426);
nor U4012 (N_4012,In_903,In_1064);
nor U4013 (N_4013,In_1023,In_802);
or U4014 (N_4014,In_188,In_730);
and U4015 (N_4015,In_1876,In_756);
nand U4016 (N_4016,In_1355,In_1344);
and U4017 (N_4017,In_1091,In_957);
nor U4018 (N_4018,In_860,In_603);
or U4019 (N_4019,In_1682,In_1227);
or U4020 (N_4020,In_1335,In_2473);
or U4021 (N_4021,In_1105,In_587);
and U4022 (N_4022,In_508,In_1938);
nand U4023 (N_4023,In_2275,In_673);
nand U4024 (N_4024,In_2362,In_373);
or U4025 (N_4025,In_1296,In_48);
or U4026 (N_4026,In_1314,In_1062);
nor U4027 (N_4027,In_462,In_630);
nor U4028 (N_4028,In_1782,In_1962);
and U4029 (N_4029,In_1691,In_798);
xnor U4030 (N_4030,In_235,In_187);
and U4031 (N_4031,In_900,In_341);
nand U4032 (N_4032,In_1314,In_2211);
nand U4033 (N_4033,In_2007,In_1998);
or U4034 (N_4034,In_249,In_2220);
or U4035 (N_4035,In_2041,In_1311);
and U4036 (N_4036,In_1470,In_712);
nand U4037 (N_4037,In_2412,In_2040);
nand U4038 (N_4038,In_607,In_499);
nor U4039 (N_4039,In_202,In_1931);
or U4040 (N_4040,In_193,In_650);
and U4041 (N_4041,In_473,In_1954);
and U4042 (N_4042,In_448,In_1413);
or U4043 (N_4043,In_479,In_1616);
nand U4044 (N_4044,In_361,In_700);
and U4045 (N_4045,In_2488,In_493);
and U4046 (N_4046,In_35,In_1471);
and U4047 (N_4047,In_1455,In_1494);
and U4048 (N_4048,In_58,In_674);
and U4049 (N_4049,In_2265,In_1770);
nand U4050 (N_4050,In_1719,In_98);
nand U4051 (N_4051,In_657,In_427);
nand U4052 (N_4052,In_1758,In_1198);
or U4053 (N_4053,In_1157,In_345);
nor U4054 (N_4054,In_1455,In_2008);
nor U4055 (N_4055,In_440,In_79);
nand U4056 (N_4056,In_1591,In_430);
nor U4057 (N_4057,In_1372,In_615);
nand U4058 (N_4058,In_814,In_357);
nor U4059 (N_4059,In_2317,In_1776);
xor U4060 (N_4060,In_930,In_1986);
and U4061 (N_4061,In_471,In_98);
or U4062 (N_4062,In_964,In_972);
nor U4063 (N_4063,In_2494,In_483);
nand U4064 (N_4064,In_1881,In_793);
nor U4065 (N_4065,In_2244,In_65);
and U4066 (N_4066,In_2327,In_1863);
and U4067 (N_4067,In_991,In_2469);
nand U4068 (N_4068,In_382,In_1876);
and U4069 (N_4069,In_1766,In_1751);
nor U4070 (N_4070,In_2359,In_955);
nor U4071 (N_4071,In_1055,In_942);
and U4072 (N_4072,In_242,In_95);
and U4073 (N_4073,In_1545,In_1361);
nand U4074 (N_4074,In_2209,In_2208);
and U4075 (N_4075,In_741,In_51);
nand U4076 (N_4076,In_1717,In_554);
or U4077 (N_4077,In_1764,In_650);
or U4078 (N_4078,In_2352,In_769);
or U4079 (N_4079,In_1704,In_2159);
and U4080 (N_4080,In_2347,In_1837);
or U4081 (N_4081,In_1112,In_777);
nand U4082 (N_4082,In_898,In_449);
nor U4083 (N_4083,In_2145,In_1677);
or U4084 (N_4084,In_1828,In_1877);
nand U4085 (N_4085,In_1065,In_1425);
or U4086 (N_4086,In_1580,In_570);
nor U4087 (N_4087,In_2385,In_1710);
or U4088 (N_4088,In_1845,In_1426);
nand U4089 (N_4089,In_673,In_1226);
nand U4090 (N_4090,In_1286,In_1961);
and U4091 (N_4091,In_1909,In_564);
or U4092 (N_4092,In_660,In_550);
and U4093 (N_4093,In_2485,In_1511);
nor U4094 (N_4094,In_1067,In_208);
nand U4095 (N_4095,In_840,In_1624);
xnor U4096 (N_4096,In_310,In_156);
nor U4097 (N_4097,In_511,In_355);
nor U4098 (N_4098,In_1665,In_2064);
nand U4099 (N_4099,In_1753,In_527);
nor U4100 (N_4100,In_144,In_1851);
or U4101 (N_4101,In_817,In_611);
xor U4102 (N_4102,In_2294,In_504);
or U4103 (N_4103,In_707,In_1213);
nand U4104 (N_4104,In_2226,In_2281);
and U4105 (N_4105,In_1901,In_125);
nand U4106 (N_4106,In_22,In_492);
or U4107 (N_4107,In_1695,In_1635);
and U4108 (N_4108,In_600,In_102);
nor U4109 (N_4109,In_2010,In_2094);
nand U4110 (N_4110,In_213,In_1139);
or U4111 (N_4111,In_829,In_1859);
and U4112 (N_4112,In_795,In_803);
or U4113 (N_4113,In_2208,In_1758);
nand U4114 (N_4114,In_1573,In_775);
or U4115 (N_4115,In_2422,In_1147);
nand U4116 (N_4116,In_1768,In_1292);
and U4117 (N_4117,In_536,In_518);
nand U4118 (N_4118,In_1511,In_1124);
and U4119 (N_4119,In_2227,In_2015);
nand U4120 (N_4120,In_2310,In_53);
nor U4121 (N_4121,In_115,In_1048);
and U4122 (N_4122,In_2389,In_1384);
nand U4123 (N_4123,In_690,In_564);
and U4124 (N_4124,In_1826,In_1222);
xnor U4125 (N_4125,In_157,In_1289);
or U4126 (N_4126,In_866,In_316);
nor U4127 (N_4127,In_87,In_1517);
nand U4128 (N_4128,In_462,In_1694);
or U4129 (N_4129,In_2178,In_1847);
nand U4130 (N_4130,In_1339,In_1106);
nor U4131 (N_4131,In_2252,In_1390);
nor U4132 (N_4132,In_1116,In_2147);
or U4133 (N_4133,In_2395,In_583);
and U4134 (N_4134,In_988,In_68);
nor U4135 (N_4135,In_1289,In_709);
nand U4136 (N_4136,In_1373,In_2410);
nor U4137 (N_4137,In_542,In_1614);
nor U4138 (N_4138,In_1389,In_1326);
nor U4139 (N_4139,In_585,In_482);
nor U4140 (N_4140,In_2064,In_750);
nor U4141 (N_4141,In_1364,In_2276);
or U4142 (N_4142,In_1536,In_1042);
and U4143 (N_4143,In_1840,In_1428);
nor U4144 (N_4144,In_2232,In_695);
and U4145 (N_4145,In_71,In_1333);
or U4146 (N_4146,In_1600,In_1752);
xor U4147 (N_4147,In_2053,In_1302);
or U4148 (N_4148,In_257,In_360);
or U4149 (N_4149,In_1987,In_1465);
or U4150 (N_4150,In_2342,In_1760);
nor U4151 (N_4151,In_121,In_1023);
nand U4152 (N_4152,In_2106,In_231);
or U4153 (N_4153,In_442,In_1114);
nand U4154 (N_4154,In_1897,In_1942);
nand U4155 (N_4155,In_1227,In_495);
nand U4156 (N_4156,In_705,In_270);
nor U4157 (N_4157,In_107,In_2235);
nor U4158 (N_4158,In_2103,In_1492);
and U4159 (N_4159,In_756,In_1513);
nand U4160 (N_4160,In_221,In_575);
nor U4161 (N_4161,In_588,In_1329);
nor U4162 (N_4162,In_288,In_477);
nor U4163 (N_4163,In_1664,In_1646);
and U4164 (N_4164,In_1122,In_1311);
nor U4165 (N_4165,In_337,In_884);
and U4166 (N_4166,In_1687,In_1252);
and U4167 (N_4167,In_2175,In_847);
nor U4168 (N_4168,In_1461,In_2344);
nand U4169 (N_4169,In_253,In_2249);
or U4170 (N_4170,In_1322,In_100);
and U4171 (N_4171,In_1925,In_118);
nand U4172 (N_4172,In_812,In_2439);
and U4173 (N_4173,In_29,In_1118);
or U4174 (N_4174,In_1053,In_718);
and U4175 (N_4175,In_1746,In_1303);
or U4176 (N_4176,In_2287,In_1452);
nor U4177 (N_4177,In_1405,In_2090);
and U4178 (N_4178,In_734,In_936);
nand U4179 (N_4179,In_90,In_2285);
or U4180 (N_4180,In_1426,In_930);
and U4181 (N_4181,In_753,In_299);
nor U4182 (N_4182,In_804,In_1653);
or U4183 (N_4183,In_1923,In_2235);
nor U4184 (N_4184,In_715,In_2043);
or U4185 (N_4185,In_964,In_380);
nand U4186 (N_4186,In_29,In_920);
nor U4187 (N_4187,In_1830,In_1654);
nor U4188 (N_4188,In_138,In_2222);
and U4189 (N_4189,In_407,In_1443);
nand U4190 (N_4190,In_756,In_2113);
or U4191 (N_4191,In_2395,In_2078);
and U4192 (N_4192,In_1723,In_1110);
nand U4193 (N_4193,In_1151,In_313);
or U4194 (N_4194,In_1196,In_2333);
nand U4195 (N_4195,In_163,In_1581);
xnor U4196 (N_4196,In_653,In_24);
and U4197 (N_4197,In_986,In_1215);
and U4198 (N_4198,In_97,In_1587);
nor U4199 (N_4199,In_1000,In_1516);
or U4200 (N_4200,In_1750,In_1);
and U4201 (N_4201,In_2353,In_2398);
nand U4202 (N_4202,In_487,In_573);
nor U4203 (N_4203,In_1109,In_4);
and U4204 (N_4204,In_1489,In_899);
nor U4205 (N_4205,In_1178,In_2335);
and U4206 (N_4206,In_387,In_121);
and U4207 (N_4207,In_401,In_45);
or U4208 (N_4208,In_1026,In_1346);
or U4209 (N_4209,In_1664,In_111);
nor U4210 (N_4210,In_964,In_630);
and U4211 (N_4211,In_2398,In_795);
and U4212 (N_4212,In_286,In_2302);
or U4213 (N_4213,In_1341,In_1197);
and U4214 (N_4214,In_602,In_1238);
nand U4215 (N_4215,In_1001,In_921);
nor U4216 (N_4216,In_588,In_2087);
and U4217 (N_4217,In_1337,In_2026);
nand U4218 (N_4218,In_813,In_2327);
or U4219 (N_4219,In_1868,In_827);
or U4220 (N_4220,In_1013,In_218);
xnor U4221 (N_4221,In_83,In_32);
nor U4222 (N_4222,In_290,In_1494);
or U4223 (N_4223,In_1866,In_1477);
and U4224 (N_4224,In_1424,In_2378);
nand U4225 (N_4225,In_2372,In_653);
nor U4226 (N_4226,In_2420,In_1600);
or U4227 (N_4227,In_1602,In_1257);
and U4228 (N_4228,In_1820,In_998);
nor U4229 (N_4229,In_1889,In_1251);
and U4230 (N_4230,In_442,In_1873);
xor U4231 (N_4231,In_1262,In_106);
nor U4232 (N_4232,In_1876,In_1525);
nand U4233 (N_4233,In_2118,In_1473);
or U4234 (N_4234,In_2251,In_308);
or U4235 (N_4235,In_532,In_1480);
or U4236 (N_4236,In_1515,In_88);
nor U4237 (N_4237,In_1535,In_2438);
and U4238 (N_4238,In_410,In_1430);
nor U4239 (N_4239,In_1891,In_471);
nor U4240 (N_4240,In_1257,In_2176);
and U4241 (N_4241,In_2130,In_1287);
and U4242 (N_4242,In_210,In_1219);
nor U4243 (N_4243,In_333,In_633);
and U4244 (N_4244,In_691,In_2411);
and U4245 (N_4245,In_208,In_716);
or U4246 (N_4246,In_2033,In_1273);
or U4247 (N_4247,In_1069,In_924);
and U4248 (N_4248,In_1195,In_2177);
and U4249 (N_4249,In_348,In_672);
nor U4250 (N_4250,In_2278,In_1558);
nand U4251 (N_4251,In_1784,In_970);
or U4252 (N_4252,In_3,In_407);
or U4253 (N_4253,In_1282,In_1212);
and U4254 (N_4254,In_1114,In_1051);
nand U4255 (N_4255,In_1383,In_2378);
and U4256 (N_4256,In_244,In_2026);
or U4257 (N_4257,In_1211,In_293);
nor U4258 (N_4258,In_528,In_742);
and U4259 (N_4259,In_892,In_1560);
nor U4260 (N_4260,In_1410,In_1111);
or U4261 (N_4261,In_621,In_2456);
nand U4262 (N_4262,In_1489,In_573);
and U4263 (N_4263,In_1125,In_2411);
nor U4264 (N_4264,In_214,In_1960);
and U4265 (N_4265,In_1508,In_423);
nand U4266 (N_4266,In_772,In_2134);
nand U4267 (N_4267,In_1124,In_1715);
nand U4268 (N_4268,In_746,In_849);
nor U4269 (N_4269,In_2254,In_1473);
nor U4270 (N_4270,In_2247,In_1857);
xnor U4271 (N_4271,In_1317,In_574);
and U4272 (N_4272,In_952,In_94);
nand U4273 (N_4273,In_753,In_2354);
nand U4274 (N_4274,In_440,In_1604);
and U4275 (N_4275,In_2220,In_1648);
nand U4276 (N_4276,In_924,In_138);
or U4277 (N_4277,In_411,In_2427);
nand U4278 (N_4278,In_1472,In_1546);
and U4279 (N_4279,In_938,In_2123);
nand U4280 (N_4280,In_528,In_205);
nand U4281 (N_4281,In_813,In_2308);
nand U4282 (N_4282,In_1999,In_769);
nor U4283 (N_4283,In_298,In_2358);
and U4284 (N_4284,In_1546,In_2267);
and U4285 (N_4285,In_780,In_2218);
nand U4286 (N_4286,In_1451,In_475);
nand U4287 (N_4287,In_2378,In_226);
nand U4288 (N_4288,In_678,In_1003);
nand U4289 (N_4289,In_286,In_2355);
xor U4290 (N_4290,In_1851,In_2014);
xor U4291 (N_4291,In_2101,In_1899);
nor U4292 (N_4292,In_777,In_104);
and U4293 (N_4293,In_14,In_2188);
nor U4294 (N_4294,In_1408,In_1090);
or U4295 (N_4295,In_2217,In_1986);
nor U4296 (N_4296,In_625,In_2194);
nand U4297 (N_4297,In_676,In_401);
nand U4298 (N_4298,In_2290,In_1267);
nand U4299 (N_4299,In_1119,In_683);
and U4300 (N_4300,In_127,In_462);
nand U4301 (N_4301,In_976,In_2327);
nand U4302 (N_4302,In_1686,In_2040);
nand U4303 (N_4303,In_1034,In_1145);
nand U4304 (N_4304,In_2257,In_997);
nor U4305 (N_4305,In_2305,In_2133);
nor U4306 (N_4306,In_1712,In_880);
and U4307 (N_4307,In_873,In_306);
nor U4308 (N_4308,In_16,In_264);
nand U4309 (N_4309,In_1322,In_2029);
and U4310 (N_4310,In_1472,In_197);
and U4311 (N_4311,In_1017,In_1134);
or U4312 (N_4312,In_250,In_1933);
and U4313 (N_4313,In_2319,In_1048);
nand U4314 (N_4314,In_460,In_1809);
and U4315 (N_4315,In_941,In_934);
and U4316 (N_4316,In_1108,In_1184);
nand U4317 (N_4317,In_331,In_39);
nor U4318 (N_4318,In_117,In_2124);
nor U4319 (N_4319,In_1791,In_1112);
and U4320 (N_4320,In_930,In_1813);
or U4321 (N_4321,In_1295,In_2198);
or U4322 (N_4322,In_441,In_1923);
and U4323 (N_4323,In_1110,In_418);
or U4324 (N_4324,In_860,In_255);
and U4325 (N_4325,In_82,In_262);
nand U4326 (N_4326,In_2223,In_742);
and U4327 (N_4327,In_633,In_326);
or U4328 (N_4328,In_2110,In_613);
nand U4329 (N_4329,In_1568,In_979);
nand U4330 (N_4330,In_801,In_613);
nor U4331 (N_4331,In_1047,In_424);
nand U4332 (N_4332,In_1358,In_469);
nor U4333 (N_4333,In_666,In_449);
or U4334 (N_4334,In_2247,In_296);
or U4335 (N_4335,In_530,In_2259);
and U4336 (N_4336,In_677,In_1874);
nand U4337 (N_4337,In_1554,In_403);
and U4338 (N_4338,In_1493,In_816);
or U4339 (N_4339,In_1030,In_1770);
or U4340 (N_4340,In_574,In_1575);
nor U4341 (N_4341,In_45,In_617);
and U4342 (N_4342,In_523,In_1856);
nand U4343 (N_4343,In_372,In_2023);
and U4344 (N_4344,In_800,In_1096);
or U4345 (N_4345,In_2434,In_1005);
or U4346 (N_4346,In_1148,In_2286);
nand U4347 (N_4347,In_1592,In_390);
xor U4348 (N_4348,In_508,In_1056);
nor U4349 (N_4349,In_1135,In_1887);
nand U4350 (N_4350,In_393,In_2438);
nand U4351 (N_4351,In_1624,In_1527);
nor U4352 (N_4352,In_1514,In_1623);
or U4353 (N_4353,In_628,In_779);
nand U4354 (N_4354,In_1989,In_623);
or U4355 (N_4355,In_964,In_667);
nor U4356 (N_4356,In_234,In_1318);
and U4357 (N_4357,In_1749,In_487);
and U4358 (N_4358,In_2119,In_1342);
or U4359 (N_4359,In_460,In_1779);
or U4360 (N_4360,In_2320,In_310);
xor U4361 (N_4361,In_2275,In_1926);
nand U4362 (N_4362,In_965,In_2046);
nand U4363 (N_4363,In_1994,In_2038);
nor U4364 (N_4364,In_280,In_1992);
and U4365 (N_4365,In_1231,In_827);
and U4366 (N_4366,In_2104,In_1213);
or U4367 (N_4367,In_2328,In_2231);
nand U4368 (N_4368,In_1805,In_1336);
and U4369 (N_4369,In_2447,In_327);
or U4370 (N_4370,In_1362,In_2280);
nand U4371 (N_4371,In_1593,In_1710);
nand U4372 (N_4372,In_886,In_2126);
and U4373 (N_4373,In_220,In_1024);
nor U4374 (N_4374,In_1744,In_546);
and U4375 (N_4375,In_2024,In_1025);
and U4376 (N_4376,In_525,In_1325);
nand U4377 (N_4377,In_679,In_489);
nor U4378 (N_4378,In_1655,In_2404);
and U4379 (N_4379,In_719,In_1925);
nand U4380 (N_4380,In_2226,In_312);
and U4381 (N_4381,In_1982,In_308);
nor U4382 (N_4382,In_2262,In_2218);
and U4383 (N_4383,In_148,In_2007);
and U4384 (N_4384,In_1975,In_1412);
nand U4385 (N_4385,In_1986,In_1347);
or U4386 (N_4386,In_1835,In_990);
and U4387 (N_4387,In_1706,In_2220);
and U4388 (N_4388,In_1587,In_2242);
nor U4389 (N_4389,In_1597,In_763);
and U4390 (N_4390,In_182,In_1411);
or U4391 (N_4391,In_396,In_855);
nand U4392 (N_4392,In_2312,In_507);
or U4393 (N_4393,In_92,In_762);
or U4394 (N_4394,In_1950,In_1294);
nand U4395 (N_4395,In_412,In_1237);
or U4396 (N_4396,In_1423,In_800);
or U4397 (N_4397,In_205,In_1329);
nor U4398 (N_4398,In_1456,In_1980);
or U4399 (N_4399,In_1991,In_252);
nand U4400 (N_4400,In_1659,In_696);
and U4401 (N_4401,In_1391,In_1661);
nand U4402 (N_4402,In_237,In_1513);
or U4403 (N_4403,In_2093,In_1033);
nor U4404 (N_4404,In_810,In_2425);
or U4405 (N_4405,In_34,In_777);
nor U4406 (N_4406,In_684,In_2241);
and U4407 (N_4407,In_1034,In_550);
nor U4408 (N_4408,In_1234,In_1879);
nor U4409 (N_4409,In_641,In_1288);
or U4410 (N_4410,In_2412,In_2276);
and U4411 (N_4411,In_662,In_2133);
nand U4412 (N_4412,In_565,In_2001);
nand U4413 (N_4413,In_272,In_2253);
nand U4414 (N_4414,In_470,In_82);
and U4415 (N_4415,In_1899,In_11);
nand U4416 (N_4416,In_324,In_27);
nor U4417 (N_4417,In_94,In_1231);
nor U4418 (N_4418,In_1125,In_821);
nand U4419 (N_4419,In_2433,In_537);
or U4420 (N_4420,In_353,In_721);
and U4421 (N_4421,In_1021,In_2137);
or U4422 (N_4422,In_2146,In_1822);
xor U4423 (N_4423,In_924,In_2444);
nor U4424 (N_4424,In_1663,In_2415);
nand U4425 (N_4425,In_1696,In_4);
and U4426 (N_4426,In_1454,In_1764);
and U4427 (N_4427,In_327,In_2084);
and U4428 (N_4428,In_2097,In_928);
nor U4429 (N_4429,In_2224,In_1883);
nand U4430 (N_4430,In_1888,In_782);
nor U4431 (N_4431,In_826,In_1801);
or U4432 (N_4432,In_710,In_1974);
and U4433 (N_4433,In_889,In_1104);
and U4434 (N_4434,In_809,In_1243);
nor U4435 (N_4435,In_1583,In_709);
nor U4436 (N_4436,In_987,In_522);
and U4437 (N_4437,In_1907,In_1971);
and U4438 (N_4438,In_672,In_2273);
nand U4439 (N_4439,In_1462,In_1705);
and U4440 (N_4440,In_1572,In_2250);
nor U4441 (N_4441,In_395,In_1875);
nand U4442 (N_4442,In_1645,In_241);
or U4443 (N_4443,In_943,In_2484);
nor U4444 (N_4444,In_919,In_283);
nor U4445 (N_4445,In_1374,In_2158);
and U4446 (N_4446,In_704,In_57);
or U4447 (N_4447,In_29,In_609);
nand U4448 (N_4448,In_907,In_1913);
or U4449 (N_4449,In_946,In_1323);
xor U4450 (N_4450,In_1120,In_1979);
nand U4451 (N_4451,In_1515,In_1661);
nor U4452 (N_4452,In_1490,In_278);
or U4453 (N_4453,In_1988,In_1938);
and U4454 (N_4454,In_1258,In_630);
nor U4455 (N_4455,In_1195,In_2479);
or U4456 (N_4456,In_1289,In_1511);
nor U4457 (N_4457,In_884,In_2120);
nand U4458 (N_4458,In_1647,In_2042);
nor U4459 (N_4459,In_1677,In_2311);
nand U4460 (N_4460,In_1123,In_1374);
nor U4461 (N_4461,In_104,In_2200);
nor U4462 (N_4462,In_1757,In_781);
nand U4463 (N_4463,In_1261,In_660);
nor U4464 (N_4464,In_511,In_371);
nor U4465 (N_4465,In_2103,In_1956);
and U4466 (N_4466,In_2076,In_1122);
nor U4467 (N_4467,In_2417,In_527);
nand U4468 (N_4468,In_2035,In_38);
and U4469 (N_4469,In_1322,In_787);
nor U4470 (N_4470,In_1175,In_1610);
xnor U4471 (N_4471,In_1991,In_91);
xnor U4472 (N_4472,In_93,In_1079);
and U4473 (N_4473,In_1138,In_1857);
and U4474 (N_4474,In_705,In_289);
or U4475 (N_4475,In_615,In_2470);
nor U4476 (N_4476,In_217,In_1652);
and U4477 (N_4477,In_558,In_943);
and U4478 (N_4478,In_796,In_762);
nand U4479 (N_4479,In_565,In_2325);
nor U4480 (N_4480,In_1885,In_615);
nor U4481 (N_4481,In_2456,In_606);
or U4482 (N_4482,In_2319,In_2246);
nand U4483 (N_4483,In_317,In_2316);
and U4484 (N_4484,In_165,In_1134);
and U4485 (N_4485,In_1239,In_2445);
or U4486 (N_4486,In_494,In_2288);
or U4487 (N_4487,In_195,In_625);
nand U4488 (N_4488,In_2239,In_854);
or U4489 (N_4489,In_1101,In_64);
nor U4490 (N_4490,In_898,In_356);
nor U4491 (N_4491,In_1001,In_2289);
or U4492 (N_4492,In_1761,In_1294);
and U4493 (N_4493,In_526,In_301);
and U4494 (N_4494,In_1468,In_792);
nor U4495 (N_4495,In_2236,In_1820);
nand U4496 (N_4496,In_792,In_527);
nand U4497 (N_4497,In_794,In_1337);
and U4498 (N_4498,In_8,In_1837);
or U4499 (N_4499,In_86,In_2182);
xor U4500 (N_4500,In_19,In_1827);
or U4501 (N_4501,In_1605,In_1415);
nand U4502 (N_4502,In_1525,In_864);
or U4503 (N_4503,In_845,In_22);
nand U4504 (N_4504,In_2204,In_1810);
nand U4505 (N_4505,In_2369,In_2293);
nor U4506 (N_4506,In_1270,In_2240);
nand U4507 (N_4507,In_1117,In_2264);
nor U4508 (N_4508,In_565,In_2098);
or U4509 (N_4509,In_1049,In_207);
nand U4510 (N_4510,In_2284,In_1972);
nand U4511 (N_4511,In_2238,In_75);
nand U4512 (N_4512,In_2453,In_1057);
nand U4513 (N_4513,In_1149,In_1009);
nor U4514 (N_4514,In_344,In_364);
nand U4515 (N_4515,In_294,In_147);
and U4516 (N_4516,In_2378,In_1486);
nand U4517 (N_4517,In_1798,In_1374);
nor U4518 (N_4518,In_1024,In_1157);
and U4519 (N_4519,In_1442,In_910);
nor U4520 (N_4520,In_382,In_1671);
or U4521 (N_4521,In_2178,In_539);
nor U4522 (N_4522,In_1461,In_1304);
nor U4523 (N_4523,In_1313,In_2408);
nor U4524 (N_4524,In_2443,In_1210);
and U4525 (N_4525,In_672,In_1143);
and U4526 (N_4526,In_864,In_1327);
xor U4527 (N_4527,In_1973,In_1037);
or U4528 (N_4528,In_2369,In_1539);
nand U4529 (N_4529,In_1289,In_922);
or U4530 (N_4530,In_1153,In_1899);
nand U4531 (N_4531,In_1282,In_1890);
or U4532 (N_4532,In_2112,In_718);
or U4533 (N_4533,In_987,In_1675);
or U4534 (N_4534,In_2188,In_267);
nor U4535 (N_4535,In_1745,In_168);
or U4536 (N_4536,In_1799,In_20);
nor U4537 (N_4537,In_363,In_1835);
nor U4538 (N_4538,In_2498,In_1580);
or U4539 (N_4539,In_523,In_939);
nor U4540 (N_4540,In_2046,In_1200);
and U4541 (N_4541,In_144,In_2346);
nor U4542 (N_4542,In_513,In_2174);
and U4543 (N_4543,In_1365,In_1788);
and U4544 (N_4544,In_1865,In_537);
nor U4545 (N_4545,In_2163,In_1520);
or U4546 (N_4546,In_2429,In_2386);
nor U4547 (N_4547,In_656,In_1449);
and U4548 (N_4548,In_640,In_2054);
nand U4549 (N_4549,In_2020,In_1707);
nor U4550 (N_4550,In_887,In_1046);
and U4551 (N_4551,In_1811,In_1479);
or U4552 (N_4552,In_2210,In_300);
or U4553 (N_4553,In_891,In_581);
nor U4554 (N_4554,In_455,In_1988);
nor U4555 (N_4555,In_1433,In_2341);
or U4556 (N_4556,In_1394,In_1853);
nand U4557 (N_4557,In_722,In_834);
nand U4558 (N_4558,In_455,In_1685);
or U4559 (N_4559,In_2277,In_1488);
and U4560 (N_4560,In_1801,In_580);
nand U4561 (N_4561,In_372,In_548);
nand U4562 (N_4562,In_910,In_1427);
nor U4563 (N_4563,In_897,In_2395);
nor U4564 (N_4564,In_499,In_1153);
nand U4565 (N_4565,In_1017,In_1176);
or U4566 (N_4566,In_837,In_2495);
and U4567 (N_4567,In_148,In_1980);
nor U4568 (N_4568,In_1735,In_1151);
nor U4569 (N_4569,In_744,In_66);
nor U4570 (N_4570,In_787,In_825);
or U4571 (N_4571,In_1104,In_334);
nand U4572 (N_4572,In_880,In_2288);
nor U4573 (N_4573,In_1400,In_821);
or U4574 (N_4574,In_1898,In_2233);
nor U4575 (N_4575,In_1147,In_2245);
and U4576 (N_4576,In_1203,In_2100);
or U4577 (N_4577,In_1857,In_1260);
nor U4578 (N_4578,In_938,In_987);
and U4579 (N_4579,In_444,In_1906);
and U4580 (N_4580,In_1937,In_1071);
nand U4581 (N_4581,In_2311,In_738);
nor U4582 (N_4582,In_122,In_239);
or U4583 (N_4583,In_777,In_2404);
nand U4584 (N_4584,In_2168,In_328);
and U4585 (N_4585,In_39,In_672);
and U4586 (N_4586,In_108,In_1056);
nor U4587 (N_4587,In_2035,In_2168);
and U4588 (N_4588,In_1357,In_1488);
nand U4589 (N_4589,In_1943,In_2134);
and U4590 (N_4590,In_28,In_2252);
nor U4591 (N_4591,In_1520,In_1557);
and U4592 (N_4592,In_1128,In_1173);
and U4593 (N_4593,In_2226,In_2465);
nand U4594 (N_4594,In_908,In_950);
or U4595 (N_4595,In_888,In_1456);
nand U4596 (N_4596,In_2443,In_122);
xor U4597 (N_4597,In_2416,In_44);
or U4598 (N_4598,In_533,In_2322);
and U4599 (N_4599,In_1391,In_96);
nor U4600 (N_4600,In_1388,In_48);
nor U4601 (N_4601,In_1943,In_117);
nor U4602 (N_4602,In_1745,In_1916);
nor U4603 (N_4603,In_498,In_1040);
xnor U4604 (N_4604,In_2198,In_1366);
or U4605 (N_4605,In_372,In_596);
nand U4606 (N_4606,In_210,In_554);
or U4607 (N_4607,In_962,In_2084);
and U4608 (N_4608,In_440,In_126);
nand U4609 (N_4609,In_2296,In_1890);
nor U4610 (N_4610,In_1921,In_1348);
nor U4611 (N_4611,In_290,In_1818);
and U4612 (N_4612,In_1097,In_208);
or U4613 (N_4613,In_539,In_1969);
and U4614 (N_4614,In_2197,In_350);
nor U4615 (N_4615,In_759,In_1638);
nor U4616 (N_4616,In_1928,In_2301);
nand U4617 (N_4617,In_1274,In_16);
or U4618 (N_4618,In_1364,In_1357);
nand U4619 (N_4619,In_560,In_431);
or U4620 (N_4620,In_1878,In_2099);
or U4621 (N_4621,In_26,In_1361);
xnor U4622 (N_4622,In_526,In_2260);
or U4623 (N_4623,In_1914,In_133);
or U4624 (N_4624,In_376,In_1314);
or U4625 (N_4625,In_282,In_565);
nand U4626 (N_4626,In_77,In_711);
and U4627 (N_4627,In_1684,In_1037);
nand U4628 (N_4628,In_1364,In_951);
nor U4629 (N_4629,In_587,In_977);
and U4630 (N_4630,In_1372,In_1938);
and U4631 (N_4631,In_2088,In_2163);
or U4632 (N_4632,In_2354,In_1129);
nand U4633 (N_4633,In_153,In_411);
or U4634 (N_4634,In_2412,In_305);
nand U4635 (N_4635,In_1560,In_1105);
and U4636 (N_4636,In_2430,In_738);
nand U4637 (N_4637,In_1024,In_1317);
nor U4638 (N_4638,In_1231,In_2191);
nor U4639 (N_4639,In_1932,In_892);
and U4640 (N_4640,In_1170,In_2076);
or U4641 (N_4641,In_1260,In_1771);
nor U4642 (N_4642,In_100,In_1233);
nand U4643 (N_4643,In_459,In_1220);
nor U4644 (N_4644,In_518,In_1279);
and U4645 (N_4645,In_586,In_1291);
and U4646 (N_4646,In_2121,In_293);
nand U4647 (N_4647,In_2357,In_1527);
and U4648 (N_4648,In_1653,In_1354);
nand U4649 (N_4649,In_2470,In_1502);
and U4650 (N_4650,In_293,In_1067);
nand U4651 (N_4651,In_392,In_1297);
nand U4652 (N_4652,In_706,In_2092);
and U4653 (N_4653,In_393,In_2127);
nand U4654 (N_4654,In_320,In_30);
nor U4655 (N_4655,In_552,In_1082);
nand U4656 (N_4656,In_263,In_1754);
or U4657 (N_4657,In_450,In_2);
or U4658 (N_4658,In_1803,In_153);
or U4659 (N_4659,In_1127,In_1984);
nand U4660 (N_4660,In_1031,In_1848);
nor U4661 (N_4661,In_524,In_1062);
or U4662 (N_4662,In_408,In_1157);
nor U4663 (N_4663,In_465,In_139);
and U4664 (N_4664,In_1477,In_638);
and U4665 (N_4665,In_508,In_1496);
or U4666 (N_4666,In_2138,In_1906);
nand U4667 (N_4667,In_244,In_1831);
nor U4668 (N_4668,In_1838,In_1287);
and U4669 (N_4669,In_1442,In_484);
or U4670 (N_4670,In_1379,In_1450);
or U4671 (N_4671,In_362,In_864);
or U4672 (N_4672,In_1385,In_2380);
nand U4673 (N_4673,In_2340,In_369);
nor U4674 (N_4674,In_793,In_2424);
and U4675 (N_4675,In_2017,In_143);
xor U4676 (N_4676,In_2387,In_1196);
nor U4677 (N_4677,In_850,In_1680);
nand U4678 (N_4678,In_563,In_1744);
or U4679 (N_4679,In_682,In_1556);
xnor U4680 (N_4680,In_802,In_2079);
and U4681 (N_4681,In_1473,In_1974);
or U4682 (N_4682,In_810,In_1320);
nor U4683 (N_4683,In_2169,In_40);
nor U4684 (N_4684,In_393,In_2286);
nor U4685 (N_4685,In_1055,In_1854);
and U4686 (N_4686,In_1863,In_903);
and U4687 (N_4687,In_451,In_63);
xor U4688 (N_4688,In_193,In_1567);
nand U4689 (N_4689,In_330,In_998);
and U4690 (N_4690,In_1468,In_904);
nand U4691 (N_4691,In_568,In_1835);
and U4692 (N_4692,In_1550,In_1311);
and U4693 (N_4693,In_1787,In_923);
and U4694 (N_4694,In_593,In_1699);
nor U4695 (N_4695,In_1102,In_366);
nand U4696 (N_4696,In_813,In_554);
or U4697 (N_4697,In_879,In_1715);
nor U4698 (N_4698,In_285,In_187);
and U4699 (N_4699,In_1454,In_2066);
nor U4700 (N_4700,In_1746,In_1330);
or U4701 (N_4701,In_1727,In_170);
or U4702 (N_4702,In_2204,In_435);
nand U4703 (N_4703,In_2233,In_689);
and U4704 (N_4704,In_988,In_1546);
and U4705 (N_4705,In_522,In_890);
nor U4706 (N_4706,In_1087,In_1990);
nor U4707 (N_4707,In_684,In_283);
nand U4708 (N_4708,In_1047,In_1541);
nor U4709 (N_4709,In_981,In_1877);
and U4710 (N_4710,In_2461,In_1528);
and U4711 (N_4711,In_2493,In_2066);
nand U4712 (N_4712,In_357,In_1304);
nand U4713 (N_4713,In_1935,In_1876);
or U4714 (N_4714,In_718,In_1517);
or U4715 (N_4715,In_725,In_1462);
xor U4716 (N_4716,In_1428,In_2221);
nand U4717 (N_4717,In_1772,In_770);
nor U4718 (N_4718,In_1616,In_1630);
or U4719 (N_4719,In_289,In_954);
and U4720 (N_4720,In_622,In_856);
nand U4721 (N_4721,In_1564,In_899);
or U4722 (N_4722,In_1355,In_1529);
and U4723 (N_4723,In_776,In_1384);
nor U4724 (N_4724,In_214,In_152);
nor U4725 (N_4725,In_2234,In_2377);
and U4726 (N_4726,In_646,In_367);
nor U4727 (N_4727,In_1467,In_2403);
nand U4728 (N_4728,In_1222,In_1817);
or U4729 (N_4729,In_643,In_1126);
or U4730 (N_4730,In_1986,In_1275);
nor U4731 (N_4731,In_2476,In_557);
or U4732 (N_4732,In_2202,In_692);
and U4733 (N_4733,In_807,In_2017);
and U4734 (N_4734,In_53,In_589);
and U4735 (N_4735,In_317,In_2283);
and U4736 (N_4736,In_1587,In_1029);
nand U4737 (N_4737,In_117,In_1842);
nand U4738 (N_4738,In_220,In_1828);
and U4739 (N_4739,In_2029,In_868);
or U4740 (N_4740,In_1325,In_545);
nand U4741 (N_4741,In_474,In_1307);
or U4742 (N_4742,In_1662,In_826);
nor U4743 (N_4743,In_1996,In_681);
xnor U4744 (N_4744,In_2119,In_1195);
nor U4745 (N_4745,In_1131,In_658);
and U4746 (N_4746,In_2177,In_2383);
or U4747 (N_4747,In_2320,In_1847);
nand U4748 (N_4748,In_1850,In_305);
nand U4749 (N_4749,In_1476,In_2091);
or U4750 (N_4750,In_1014,In_9);
or U4751 (N_4751,In_1682,In_1592);
and U4752 (N_4752,In_697,In_1138);
or U4753 (N_4753,In_1982,In_2336);
and U4754 (N_4754,In_53,In_592);
nor U4755 (N_4755,In_1961,In_154);
nand U4756 (N_4756,In_944,In_1662);
nor U4757 (N_4757,In_530,In_241);
nand U4758 (N_4758,In_624,In_408);
nand U4759 (N_4759,In_870,In_85);
nor U4760 (N_4760,In_1314,In_2224);
nor U4761 (N_4761,In_97,In_1978);
nor U4762 (N_4762,In_31,In_881);
or U4763 (N_4763,In_1988,In_700);
or U4764 (N_4764,In_570,In_2202);
and U4765 (N_4765,In_149,In_1034);
and U4766 (N_4766,In_500,In_682);
nor U4767 (N_4767,In_1064,In_1848);
nor U4768 (N_4768,In_575,In_2399);
and U4769 (N_4769,In_1990,In_552);
or U4770 (N_4770,In_1638,In_369);
nor U4771 (N_4771,In_289,In_723);
nor U4772 (N_4772,In_1109,In_59);
or U4773 (N_4773,In_1799,In_1174);
and U4774 (N_4774,In_1148,In_872);
nand U4775 (N_4775,In_849,In_536);
and U4776 (N_4776,In_1070,In_423);
nor U4777 (N_4777,In_781,In_286);
nor U4778 (N_4778,In_1952,In_525);
and U4779 (N_4779,In_1305,In_1356);
or U4780 (N_4780,In_479,In_209);
and U4781 (N_4781,In_1497,In_1449);
or U4782 (N_4782,In_442,In_36);
nand U4783 (N_4783,In_2075,In_1938);
nor U4784 (N_4784,In_2034,In_932);
nand U4785 (N_4785,In_1454,In_157);
nand U4786 (N_4786,In_2142,In_1845);
nor U4787 (N_4787,In_196,In_448);
nand U4788 (N_4788,In_365,In_2243);
xnor U4789 (N_4789,In_488,In_2033);
nor U4790 (N_4790,In_2206,In_23);
nor U4791 (N_4791,In_349,In_2405);
nand U4792 (N_4792,In_2256,In_32);
nand U4793 (N_4793,In_1017,In_1617);
nand U4794 (N_4794,In_1682,In_853);
and U4795 (N_4795,In_2298,In_830);
nor U4796 (N_4796,In_2232,In_2063);
nand U4797 (N_4797,In_2378,In_1763);
and U4798 (N_4798,In_296,In_1700);
nor U4799 (N_4799,In_2,In_609);
nand U4800 (N_4800,In_1338,In_1875);
and U4801 (N_4801,In_443,In_1353);
nand U4802 (N_4802,In_174,In_125);
or U4803 (N_4803,In_20,In_532);
or U4804 (N_4804,In_2060,In_381);
nand U4805 (N_4805,In_296,In_2205);
and U4806 (N_4806,In_2268,In_309);
or U4807 (N_4807,In_1660,In_1019);
nand U4808 (N_4808,In_1873,In_2297);
xor U4809 (N_4809,In_2367,In_1905);
nand U4810 (N_4810,In_1599,In_591);
and U4811 (N_4811,In_2370,In_113);
or U4812 (N_4812,In_987,In_391);
and U4813 (N_4813,In_1000,In_1279);
nand U4814 (N_4814,In_1172,In_138);
xnor U4815 (N_4815,In_1510,In_895);
and U4816 (N_4816,In_1510,In_2125);
xor U4817 (N_4817,In_801,In_1280);
and U4818 (N_4818,In_2080,In_2326);
xnor U4819 (N_4819,In_1346,In_1933);
nand U4820 (N_4820,In_680,In_724);
and U4821 (N_4821,In_2179,In_87);
nand U4822 (N_4822,In_2382,In_2287);
nand U4823 (N_4823,In_778,In_454);
nand U4824 (N_4824,In_2477,In_1585);
and U4825 (N_4825,In_553,In_2423);
nor U4826 (N_4826,In_1169,In_1319);
nor U4827 (N_4827,In_1347,In_2318);
or U4828 (N_4828,In_498,In_726);
nand U4829 (N_4829,In_1137,In_1080);
and U4830 (N_4830,In_880,In_288);
and U4831 (N_4831,In_1588,In_1052);
and U4832 (N_4832,In_1886,In_1099);
nand U4833 (N_4833,In_1571,In_2486);
and U4834 (N_4834,In_2359,In_174);
xor U4835 (N_4835,In_81,In_464);
and U4836 (N_4836,In_935,In_738);
nand U4837 (N_4837,In_813,In_1936);
or U4838 (N_4838,In_259,In_2424);
or U4839 (N_4839,In_500,In_1838);
nor U4840 (N_4840,In_470,In_0);
nand U4841 (N_4841,In_963,In_1200);
and U4842 (N_4842,In_803,In_1416);
nand U4843 (N_4843,In_2265,In_1493);
xnor U4844 (N_4844,In_464,In_473);
nand U4845 (N_4845,In_356,In_437);
nor U4846 (N_4846,In_1281,In_2239);
nor U4847 (N_4847,In_1529,In_190);
or U4848 (N_4848,In_450,In_1237);
and U4849 (N_4849,In_404,In_207);
and U4850 (N_4850,In_698,In_1597);
nor U4851 (N_4851,In_137,In_558);
nor U4852 (N_4852,In_757,In_931);
or U4853 (N_4853,In_1153,In_1828);
and U4854 (N_4854,In_1482,In_199);
or U4855 (N_4855,In_984,In_758);
nand U4856 (N_4856,In_2266,In_742);
and U4857 (N_4857,In_2001,In_1525);
and U4858 (N_4858,In_1787,In_1786);
nand U4859 (N_4859,In_1430,In_186);
or U4860 (N_4860,In_1889,In_1688);
nor U4861 (N_4861,In_1584,In_1179);
nand U4862 (N_4862,In_1036,In_1948);
or U4863 (N_4863,In_238,In_1901);
nand U4864 (N_4864,In_576,In_2389);
nor U4865 (N_4865,In_1669,In_129);
and U4866 (N_4866,In_2275,In_717);
nand U4867 (N_4867,In_2293,In_295);
nand U4868 (N_4868,In_1272,In_2288);
and U4869 (N_4869,In_690,In_627);
or U4870 (N_4870,In_1471,In_1615);
or U4871 (N_4871,In_1055,In_2070);
nand U4872 (N_4872,In_763,In_2053);
nor U4873 (N_4873,In_1810,In_48);
nand U4874 (N_4874,In_1367,In_1415);
and U4875 (N_4875,In_613,In_582);
nand U4876 (N_4876,In_938,In_2382);
or U4877 (N_4877,In_729,In_71);
nor U4878 (N_4878,In_1461,In_1424);
nand U4879 (N_4879,In_882,In_1100);
nor U4880 (N_4880,In_898,In_1708);
nand U4881 (N_4881,In_1901,In_2406);
and U4882 (N_4882,In_432,In_2049);
nor U4883 (N_4883,In_865,In_1878);
nor U4884 (N_4884,In_112,In_1145);
nor U4885 (N_4885,In_843,In_1870);
or U4886 (N_4886,In_2090,In_2370);
nand U4887 (N_4887,In_877,In_551);
nor U4888 (N_4888,In_637,In_1138);
and U4889 (N_4889,In_1028,In_2217);
and U4890 (N_4890,In_2311,In_953);
nand U4891 (N_4891,In_1137,In_2329);
nand U4892 (N_4892,In_2343,In_483);
nand U4893 (N_4893,In_34,In_1493);
nor U4894 (N_4894,In_2042,In_647);
nand U4895 (N_4895,In_2376,In_2224);
and U4896 (N_4896,In_252,In_2040);
and U4897 (N_4897,In_838,In_2150);
nand U4898 (N_4898,In_2227,In_697);
and U4899 (N_4899,In_1450,In_1912);
nand U4900 (N_4900,In_888,In_218);
nor U4901 (N_4901,In_1214,In_2373);
or U4902 (N_4902,In_1180,In_1477);
or U4903 (N_4903,In_287,In_2206);
or U4904 (N_4904,In_473,In_2164);
nor U4905 (N_4905,In_1072,In_1892);
nor U4906 (N_4906,In_305,In_38);
nand U4907 (N_4907,In_1752,In_2312);
and U4908 (N_4908,In_1101,In_1068);
and U4909 (N_4909,In_896,In_747);
nand U4910 (N_4910,In_1487,In_219);
and U4911 (N_4911,In_924,In_605);
nand U4912 (N_4912,In_1848,In_2320);
nor U4913 (N_4913,In_1565,In_68);
or U4914 (N_4914,In_1906,In_1176);
nor U4915 (N_4915,In_1152,In_1306);
or U4916 (N_4916,In_322,In_1835);
or U4917 (N_4917,In_1516,In_2012);
or U4918 (N_4918,In_207,In_2435);
and U4919 (N_4919,In_990,In_1634);
and U4920 (N_4920,In_231,In_1212);
nor U4921 (N_4921,In_1699,In_827);
nor U4922 (N_4922,In_1174,In_2154);
and U4923 (N_4923,In_2127,In_1504);
nand U4924 (N_4924,In_861,In_2264);
nand U4925 (N_4925,In_1710,In_1509);
xnor U4926 (N_4926,In_222,In_1936);
nor U4927 (N_4927,In_1438,In_1315);
or U4928 (N_4928,In_2175,In_1616);
and U4929 (N_4929,In_960,In_1519);
or U4930 (N_4930,In_2277,In_859);
and U4931 (N_4931,In_1592,In_160);
nor U4932 (N_4932,In_1848,In_574);
or U4933 (N_4933,In_740,In_757);
or U4934 (N_4934,In_323,In_620);
nor U4935 (N_4935,In_2329,In_2170);
nor U4936 (N_4936,In_1482,In_1649);
nand U4937 (N_4937,In_1102,In_70);
nand U4938 (N_4938,In_1197,In_1306);
nor U4939 (N_4939,In_184,In_2131);
nand U4940 (N_4940,In_2377,In_2351);
and U4941 (N_4941,In_2182,In_2351);
or U4942 (N_4942,In_1522,In_1905);
or U4943 (N_4943,In_572,In_819);
and U4944 (N_4944,In_1289,In_1270);
nand U4945 (N_4945,In_1450,In_917);
nand U4946 (N_4946,In_1265,In_1192);
nand U4947 (N_4947,In_199,In_534);
or U4948 (N_4948,In_1834,In_928);
nor U4949 (N_4949,In_998,In_2293);
and U4950 (N_4950,In_132,In_2296);
nor U4951 (N_4951,In_695,In_1439);
or U4952 (N_4952,In_1107,In_926);
nor U4953 (N_4953,In_574,In_174);
and U4954 (N_4954,In_2114,In_2414);
or U4955 (N_4955,In_109,In_1010);
nand U4956 (N_4956,In_1532,In_497);
nor U4957 (N_4957,In_175,In_1098);
and U4958 (N_4958,In_1221,In_544);
nor U4959 (N_4959,In_2457,In_402);
nand U4960 (N_4960,In_2457,In_1559);
or U4961 (N_4961,In_1677,In_1399);
or U4962 (N_4962,In_367,In_1122);
or U4963 (N_4963,In_1226,In_2152);
and U4964 (N_4964,In_161,In_151);
nor U4965 (N_4965,In_1578,In_10);
and U4966 (N_4966,In_1289,In_1540);
and U4967 (N_4967,In_202,In_1511);
and U4968 (N_4968,In_1907,In_2264);
nand U4969 (N_4969,In_467,In_1681);
or U4970 (N_4970,In_974,In_953);
and U4971 (N_4971,In_819,In_1191);
or U4972 (N_4972,In_515,In_1647);
and U4973 (N_4973,In_1153,In_2382);
nor U4974 (N_4974,In_323,In_1160);
nand U4975 (N_4975,In_826,In_988);
or U4976 (N_4976,In_1628,In_838);
nor U4977 (N_4977,In_438,In_753);
or U4978 (N_4978,In_1962,In_669);
nor U4979 (N_4979,In_429,In_1399);
nor U4980 (N_4980,In_1676,In_2344);
and U4981 (N_4981,In_1853,In_1711);
and U4982 (N_4982,In_661,In_2202);
and U4983 (N_4983,In_1012,In_1170);
nor U4984 (N_4984,In_1085,In_2013);
nand U4985 (N_4985,In_2406,In_1402);
xnor U4986 (N_4986,In_832,In_1745);
and U4987 (N_4987,In_1447,In_1964);
xnor U4988 (N_4988,In_1550,In_2454);
nor U4989 (N_4989,In_1627,In_1769);
and U4990 (N_4990,In_401,In_997);
or U4991 (N_4991,In_1057,In_941);
nand U4992 (N_4992,In_1674,In_1446);
and U4993 (N_4993,In_531,In_1123);
nor U4994 (N_4994,In_2081,In_773);
nor U4995 (N_4995,In_1675,In_2192);
nor U4996 (N_4996,In_1491,In_1321);
and U4997 (N_4997,In_2129,In_1104);
nor U4998 (N_4998,In_168,In_404);
or U4999 (N_4999,In_709,In_1891);
nor U5000 (N_5000,N_3310,N_4936);
or U5001 (N_5001,N_343,N_1347);
and U5002 (N_5002,N_1148,N_2614);
nand U5003 (N_5003,N_359,N_2315);
nor U5004 (N_5004,N_3302,N_4001);
nor U5005 (N_5005,N_4005,N_2513);
and U5006 (N_5006,N_2394,N_4416);
and U5007 (N_5007,N_586,N_138);
nand U5008 (N_5008,N_2542,N_430);
or U5009 (N_5009,N_4914,N_498);
and U5010 (N_5010,N_2543,N_3349);
and U5011 (N_5011,N_4349,N_340);
or U5012 (N_5012,N_1774,N_4368);
and U5013 (N_5013,N_4760,N_3535);
and U5014 (N_5014,N_912,N_3386);
or U5015 (N_5015,N_2926,N_568);
nor U5016 (N_5016,N_2971,N_3093);
and U5017 (N_5017,N_2324,N_3517);
nand U5018 (N_5018,N_1573,N_1010);
and U5019 (N_5019,N_4500,N_297);
nand U5020 (N_5020,N_3172,N_2725);
and U5021 (N_5021,N_3278,N_2400);
nand U5022 (N_5022,N_3836,N_36);
or U5023 (N_5023,N_3473,N_1337);
nor U5024 (N_5024,N_780,N_1380);
or U5025 (N_5025,N_3231,N_4950);
or U5026 (N_5026,N_3770,N_602);
or U5027 (N_5027,N_3890,N_3225);
or U5028 (N_5028,N_4387,N_4877);
nor U5029 (N_5029,N_2135,N_441);
nand U5030 (N_5030,N_537,N_3718);
and U5031 (N_5031,N_2960,N_933);
and U5032 (N_5032,N_290,N_1439);
xor U5033 (N_5033,N_2270,N_1957);
and U5034 (N_5034,N_3686,N_2667);
and U5035 (N_5035,N_104,N_4076);
nand U5036 (N_5036,N_581,N_3105);
and U5037 (N_5037,N_860,N_2418);
and U5038 (N_5038,N_4614,N_949);
nand U5039 (N_5039,N_3226,N_2829);
nor U5040 (N_5040,N_4596,N_1084);
and U5041 (N_5041,N_2250,N_1053);
and U5042 (N_5042,N_1560,N_110);
nor U5043 (N_5043,N_4243,N_1801);
and U5044 (N_5044,N_3173,N_52);
or U5045 (N_5045,N_3229,N_194);
nand U5046 (N_5046,N_3014,N_4549);
or U5047 (N_5047,N_468,N_4627);
or U5048 (N_5048,N_1875,N_4136);
and U5049 (N_5049,N_4528,N_3889);
or U5050 (N_5050,N_4605,N_2658);
nand U5051 (N_5051,N_852,N_1836);
or U5052 (N_5052,N_2824,N_1041);
nand U5053 (N_5053,N_3394,N_91);
nor U5054 (N_5054,N_1477,N_1061);
nand U5055 (N_5055,N_4283,N_3722);
nor U5056 (N_5056,N_4172,N_3498);
and U5057 (N_5057,N_78,N_257);
nand U5058 (N_5058,N_1945,N_3725);
xor U5059 (N_5059,N_2225,N_2556);
nor U5060 (N_5060,N_4372,N_240);
and U5061 (N_5061,N_1189,N_3994);
or U5062 (N_5062,N_1808,N_416);
and U5063 (N_5063,N_3500,N_1014);
or U5064 (N_5064,N_3511,N_220);
nor U5065 (N_5065,N_2395,N_3233);
nand U5066 (N_5066,N_4809,N_2622);
and U5067 (N_5067,N_4742,N_2771);
nand U5068 (N_5068,N_95,N_1604);
nand U5069 (N_5069,N_3094,N_527);
nor U5070 (N_5070,N_2252,N_1640);
nand U5071 (N_5071,N_1228,N_3887);
xnor U5072 (N_5072,N_3631,N_559);
and U5073 (N_5073,N_2657,N_2372);
and U5074 (N_5074,N_945,N_2274);
nand U5075 (N_5075,N_4872,N_3230);
nor U5076 (N_5076,N_4466,N_767);
nand U5077 (N_5077,N_3973,N_34);
nand U5078 (N_5078,N_1071,N_812);
nand U5079 (N_5079,N_1113,N_254);
nor U5080 (N_5080,N_2902,N_1270);
nor U5081 (N_5081,N_2433,N_2010);
nor U5082 (N_5082,N_3204,N_2473);
nor U5083 (N_5083,N_2592,N_3030);
nand U5084 (N_5084,N_590,N_944);
nand U5085 (N_5085,N_510,N_3934);
nor U5086 (N_5086,N_1466,N_3313);
nor U5087 (N_5087,N_2936,N_490);
and U5088 (N_5088,N_1981,N_3541);
nand U5089 (N_5089,N_1078,N_3086);
xnor U5090 (N_5090,N_4770,N_4677);
or U5091 (N_5091,N_378,N_205);
nand U5092 (N_5092,N_2665,N_982);
and U5093 (N_5093,N_2790,N_2647);
and U5094 (N_5094,N_2442,N_4850);
or U5095 (N_5095,N_2033,N_3301);
nor U5096 (N_5096,N_3685,N_315);
nand U5097 (N_5097,N_4274,N_2819);
and U5098 (N_5098,N_4735,N_769);
and U5099 (N_5099,N_4488,N_2110);
and U5100 (N_5100,N_4719,N_473);
and U5101 (N_5101,N_1138,N_4137);
and U5102 (N_5102,N_3041,N_4984);
nand U5103 (N_5103,N_2758,N_2890);
nand U5104 (N_5104,N_1177,N_2438);
or U5105 (N_5105,N_1795,N_4712);
or U5106 (N_5106,N_1326,N_1844);
nor U5107 (N_5107,N_1388,N_4553);
nor U5108 (N_5108,N_4412,N_520);
and U5109 (N_5109,N_310,N_425);
nor U5110 (N_5110,N_1658,N_2077);
and U5111 (N_5111,N_4434,N_2288);
nor U5112 (N_5112,N_2554,N_1351);
and U5113 (N_5113,N_4916,N_3788);
nor U5114 (N_5114,N_2152,N_4278);
nor U5115 (N_5115,N_3491,N_2440);
or U5116 (N_5116,N_4004,N_2413);
and U5117 (N_5117,N_1026,N_19);
or U5118 (N_5118,N_329,N_3650);
nor U5119 (N_5119,N_3830,N_3923);
nor U5120 (N_5120,N_2741,N_364);
xnor U5121 (N_5121,N_267,N_3104);
and U5122 (N_5122,N_3780,N_3234);
and U5123 (N_5123,N_4143,N_3360);
nand U5124 (N_5124,N_3243,N_1058);
xnor U5125 (N_5125,N_1419,N_715);
xnor U5126 (N_5126,N_696,N_127);
or U5127 (N_5127,N_4887,N_4542);
nand U5128 (N_5128,N_2251,N_39);
nor U5129 (N_5129,N_253,N_2661);
and U5130 (N_5130,N_3678,N_2880);
or U5131 (N_5131,N_1108,N_4366);
nor U5132 (N_5132,N_4604,N_875);
nor U5133 (N_5133,N_4418,N_4805);
xor U5134 (N_5134,N_2978,N_604);
nand U5135 (N_5135,N_1778,N_407);
and U5136 (N_5136,N_1623,N_3122);
and U5137 (N_5137,N_4775,N_193);
and U5138 (N_5138,N_1846,N_4721);
and U5139 (N_5139,N_1015,N_2654);
nor U5140 (N_5140,N_139,N_474);
nor U5141 (N_5141,N_2017,N_3010);
nand U5142 (N_5142,N_819,N_1833);
nor U5143 (N_5143,N_2500,N_4360);
or U5144 (N_5144,N_229,N_841);
and U5145 (N_5145,N_989,N_1710);
xor U5146 (N_5146,N_293,N_1780);
nand U5147 (N_5147,N_4700,N_3680);
nor U5148 (N_5148,N_4122,N_3139);
nand U5149 (N_5149,N_2302,N_1669);
or U5150 (N_5150,N_585,N_4580);
or U5151 (N_5151,N_1476,N_4864);
nor U5152 (N_5152,N_993,N_2720);
and U5153 (N_5153,N_3540,N_3411);
and U5154 (N_5154,N_437,N_825);
nor U5155 (N_5155,N_4455,N_4388);
nand U5156 (N_5156,N_4990,N_4014);
and U5157 (N_5157,N_3213,N_3670);
nor U5158 (N_5158,N_4726,N_3177);
and U5159 (N_5159,N_4876,N_1223);
nand U5160 (N_5160,N_2334,N_2600);
and U5161 (N_5161,N_3857,N_1902);
nor U5162 (N_5162,N_4968,N_4408);
nand U5163 (N_5163,N_3152,N_2745);
and U5164 (N_5164,N_3991,N_2316);
and U5165 (N_5165,N_2740,N_2211);
nand U5166 (N_5166,N_1158,N_41);
nor U5167 (N_5167,N_2703,N_4428);
or U5168 (N_5168,N_3572,N_3833);
nand U5169 (N_5169,N_4903,N_3646);
and U5170 (N_5170,N_879,N_3098);
or U5171 (N_5171,N_4093,N_1204);
nor U5172 (N_5172,N_446,N_641);
nor U5173 (N_5173,N_1164,N_2276);
nand U5174 (N_5174,N_2519,N_4);
nor U5175 (N_5175,N_1564,N_260);
and U5176 (N_5176,N_496,N_157);
or U5177 (N_5177,N_4295,N_4287);
nor U5178 (N_5178,N_3866,N_3180);
nand U5179 (N_5179,N_4685,N_3194);
nor U5180 (N_5180,N_3927,N_832);
xor U5181 (N_5181,N_4730,N_3146);
nand U5182 (N_5182,N_1149,N_3912);
nor U5183 (N_5183,N_1978,N_1589);
nor U5184 (N_5184,N_1184,N_4406);
or U5185 (N_5185,N_1211,N_2392);
or U5186 (N_5186,N_1430,N_4346);
or U5187 (N_5187,N_1673,N_1815);
or U5188 (N_5188,N_4884,N_1511);
nor U5189 (N_5189,N_1356,N_3885);
and U5190 (N_5190,N_1565,N_3902);
nand U5191 (N_5191,N_301,N_1517);
nor U5192 (N_5192,N_2924,N_1112);
and U5193 (N_5193,N_370,N_4858);
nand U5194 (N_5194,N_4329,N_1865);
or U5195 (N_5195,N_1441,N_4407);
and U5196 (N_5196,N_4907,N_1130);
nor U5197 (N_5197,N_1412,N_4253);
nand U5198 (N_5198,N_3892,N_4139);
nor U5199 (N_5199,N_1697,N_3043);
and U5200 (N_5200,N_3075,N_4110);
nor U5201 (N_5201,N_1965,N_3948);
nor U5202 (N_5202,N_3615,N_2635);
nor U5203 (N_5203,N_271,N_186);
nand U5204 (N_5204,N_4281,N_3412);
and U5205 (N_5205,N_3121,N_3297);
nand U5206 (N_5206,N_939,N_4906);
nand U5207 (N_5207,N_4559,N_984);
or U5208 (N_5208,N_4327,N_2626);
xor U5209 (N_5209,N_2037,N_4495);
and U5210 (N_5210,N_752,N_3416);
or U5211 (N_5211,N_2688,N_125);
or U5212 (N_5212,N_94,N_4121);
and U5213 (N_5213,N_3006,N_2130);
or U5214 (N_5214,N_3215,N_3537);
nand U5215 (N_5215,N_1037,N_4856);
nand U5216 (N_5216,N_2406,N_797);
nand U5217 (N_5217,N_623,N_753);
nand U5218 (N_5218,N_3971,N_4870);
nor U5219 (N_5219,N_4019,N_2532);
nor U5220 (N_5220,N_4954,N_4167);
and U5221 (N_5221,N_942,N_679);
nand U5222 (N_5222,N_1044,N_4361);
nor U5223 (N_5223,N_123,N_433);
nand U5224 (N_5224,N_2985,N_4022);
nor U5225 (N_5225,N_4953,N_2835);
and U5226 (N_5226,N_2687,N_2646);
and U5227 (N_5227,N_3112,N_1977);
and U5228 (N_5228,N_1295,N_3931);
or U5229 (N_5229,N_3848,N_2948);
or U5230 (N_5230,N_1721,N_3381);
nand U5231 (N_5231,N_2774,N_3831);
nor U5232 (N_5232,N_3283,N_3672);
or U5233 (N_5233,N_2853,N_4904);
and U5234 (N_5234,N_282,N_4128);
nand U5235 (N_5235,N_2128,N_488);
or U5236 (N_5236,N_3626,N_1153);
and U5237 (N_5237,N_3363,N_3271);
nand U5238 (N_5238,N_4741,N_734);
xor U5239 (N_5239,N_1332,N_1552);
nor U5240 (N_5240,N_4105,N_3758);
nand U5241 (N_5241,N_2139,N_1145);
nor U5242 (N_5242,N_1373,N_3026);
and U5243 (N_5243,N_2846,N_1747);
or U5244 (N_5244,N_636,N_2942);
nand U5245 (N_5245,N_3087,N_375);
nand U5246 (N_5246,N_674,N_2709);
and U5247 (N_5247,N_429,N_2845);
nor U5248 (N_5248,N_2927,N_2675);
xor U5249 (N_5249,N_3554,N_2263);
or U5250 (N_5250,N_516,N_4077);
nand U5251 (N_5251,N_4066,N_3577);
xor U5252 (N_5252,N_402,N_3368);
nor U5253 (N_5253,N_589,N_1689);
and U5254 (N_5254,N_2430,N_836);
nor U5255 (N_5255,N_4912,N_4308);
or U5256 (N_5256,N_3628,N_591);
nor U5257 (N_5257,N_32,N_955);
nor U5258 (N_5258,N_3940,N_1948);
or U5259 (N_5259,N_398,N_3551);
and U5260 (N_5260,N_1251,N_1767);
nand U5261 (N_5261,N_1793,N_1591);
and U5262 (N_5262,N_3322,N_2203);
and U5263 (N_5263,N_318,N_3961);
nand U5264 (N_5264,N_519,N_2022);
nand U5265 (N_5265,N_4572,N_3235);
nand U5266 (N_5266,N_422,N_4744);
and U5267 (N_5267,N_4170,N_4225);
and U5268 (N_5268,N_1907,N_4797);
nand U5269 (N_5269,N_671,N_2634);
and U5270 (N_5270,N_612,N_911);
and U5271 (N_5271,N_2950,N_3896);
nor U5272 (N_5272,N_2455,N_3657);
or U5273 (N_5273,N_4727,N_2059);
and U5274 (N_5274,N_2855,N_4922);
nor U5275 (N_5275,N_2050,N_4010);
nor U5276 (N_5276,N_3189,N_351);
nand U5277 (N_5277,N_2861,N_470);
nor U5278 (N_5278,N_4835,N_2478);
and U5279 (N_5279,N_642,N_4588);
nand U5280 (N_5280,N_639,N_320);
or U5281 (N_5281,N_4030,N_4567);
or U5282 (N_5282,N_3712,N_2764);
nand U5283 (N_5283,N_1416,N_1513);
nor U5284 (N_5284,N_3175,N_2312);
or U5285 (N_5285,N_3339,N_920);
or U5286 (N_5286,N_4717,N_4213);
nand U5287 (N_5287,N_4338,N_3861);
nand U5288 (N_5288,N_4198,N_1630);
or U5289 (N_5289,N_3398,N_3096);
nor U5290 (N_5290,N_544,N_1855);
nand U5291 (N_5291,N_1512,N_2322);
nand U5292 (N_5292,N_122,N_4385);
nor U5293 (N_5293,N_4980,N_563);
nor U5294 (N_5294,N_1989,N_2876);
nor U5295 (N_5295,N_3683,N_2627);
or U5296 (N_5296,N_1216,N_4740);
nor U5297 (N_5297,N_2599,N_1843);
or U5298 (N_5298,N_22,N_1849);
and U5299 (N_5299,N_1881,N_1825);
nand U5300 (N_5300,N_3395,N_4271);
nor U5301 (N_5301,N_2120,N_1996);
or U5302 (N_5302,N_3478,N_1156);
nor U5303 (N_5303,N_2265,N_1209);
nand U5304 (N_5304,N_3065,N_975);
nor U5305 (N_5305,N_4692,N_2159);
and U5306 (N_5306,N_1374,N_4080);
nor U5307 (N_5307,N_2154,N_2437);
or U5308 (N_5308,N_4736,N_515);
or U5309 (N_5309,N_1804,N_2264);
xnor U5310 (N_5310,N_3151,N_1414);
nor U5311 (N_5311,N_795,N_4475);
nor U5312 (N_5312,N_2759,N_3655);
and U5313 (N_5313,N_807,N_1530);
nand U5314 (N_5314,N_314,N_1398);
or U5315 (N_5315,N_4516,N_2466);
nand U5316 (N_5316,N_1862,N_3978);
nor U5317 (N_5317,N_2097,N_2648);
or U5318 (N_5318,N_1915,N_864);
and U5319 (N_5319,N_2974,N_779);
nor U5320 (N_5320,N_2522,N_856);
and U5321 (N_5321,N_2769,N_2713);
and U5322 (N_5322,N_724,N_1773);
nand U5323 (N_5323,N_3490,N_2305);
nand U5324 (N_5324,N_565,N_2539);
nor U5325 (N_5325,N_2078,N_4160);
nand U5326 (N_5326,N_3079,N_412);
nand U5327 (N_5327,N_2357,N_1242);
nand U5328 (N_5328,N_2218,N_367);
and U5329 (N_5329,N_3786,N_4836);
nor U5330 (N_5330,N_289,N_3674);
and U5331 (N_5331,N_609,N_3950);
nand U5332 (N_5332,N_3164,N_2307);
and U5333 (N_5333,N_890,N_774);
nor U5334 (N_5334,N_816,N_4205);
or U5335 (N_5335,N_4843,N_2506);
or U5336 (N_5336,N_517,N_2184);
nor U5337 (N_5337,N_213,N_698);
and U5338 (N_5338,N_245,N_4514);
and U5339 (N_5339,N_4060,N_449);
or U5340 (N_5340,N_3980,N_4266);
or U5341 (N_5341,N_2823,N_332);
nor U5342 (N_5342,N_2416,N_4085);
or U5343 (N_5343,N_4831,N_4078);
nor U5344 (N_5344,N_4071,N_2236);
nor U5345 (N_5345,N_4923,N_4895);
nor U5346 (N_5346,N_116,N_1188);
and U5347 (N_5347,N_3936,N_2202);
nor U5348 (N_5348,N_2089,N_1066);
nor U5349 (N_5349,N_3983,N_4427);
nand U5350 (N_5350,N_4917,N_4367);
nand U5351 (N_5351,N_941,N_4787);
nand U5352 (N_5352,N_4557,N_76);
nor U5353 (N_5353,N_3762,N_1447);
or U5354 (N_5354,N_1803,N_4460);
and U5355 (N_5355,N_2517,N_2621);
nor U5356 (N_5356,N_3543,N_3208);
nand U5357 (N_5357,N_179,N_3544);
and U5358 (N_5358,N_3633,N_931);
nor U5359 (N_5359,N_45,N_459);
nand U5360 (N_5360,N_3291,N_1488);
or U5361 (N_5361,N_614,N_2140);
or U5362 (N_5362,N_140,N_4355);
and U5363 (N_5363,N_418,N_4467);
nor U5364 (N_5364,N_1614,N_3843);
xor U5365 (N_5365,N_1578,N_2768);
nand U5366 (N_5366,N_1282,N_409);
or U5367 (N_5367,N_3601,N_4020);
nand U5368 (N_5368,N_3749,N_3299);
and U5369 (N_5369,N_2802,N_714);
nor U5370 (N_5370,N_4034,N_562);
nor U5371 (N_5371,N_2718,N_2964);
nor U5372 (N_5372,N_1340,N_2286);
and U5373 (N_5373,N_4555,N_4182);
nand U5374 (N_5374,N_834,N_4072);
nand U5375 (N_5375,N_708,N_2669);
and U5376 (N_5376,N_738,N_1093);
nor U5377 (N_5377,N_3364,N_1147);
or U5378 (N_5378,N_4468,N_1999);
xnor U5379 (N_5379,N_3400,N_1303);
nor U5380 (N_5380,N_2629,N_2460);
or U5381 (N_5381,N_762,N_1940);
nor U5382 (N_5382,N_2535,N_3501);
and U5383 (N_5383,N_1453,N_1302);
or U5384 (N_5384,N_1612,N_4017);
nand U5385 (N_5385,N_3461,N_523);
or U5386 (N_5386,N_3277,N_353);
nor U5387 (N_5387,N_4403,N_1493);
or U5388 (N_5388,N_115,N_3066);
and U5389 (N_5389,N_4669,N_1615);
or U5390 (N_5390,N_3521,N_2239);
and U5391 (N_5391,N_4657,N_4834);
nor U5392 (N_5392,N_3997,N_403);
nor U5393 (N_5393,N_4280,N_4963);
and U5394 (N_5394,N_4796,N_2071);
nor U5395 (N_5395,N_2194,N_2219);
nor U5396 (N_5396,N_1923,N_967);
or U5397 (N_5397,N_4344,N_69);
nor U5398 (N_5398,N_152,N_4714);
and U5399 (N_5399,N_4556,N_1943);
and U5400 (N_5400,N_3150,N_851);
or U5401 (N_5401,N_507,N_828);
and U5402 (N_5402,N_2570,N_1092);
nor U5403 (N_5403,N_1482,N_4039);
nor U5404 (N_5404,N_2951,N_3254);
nor U5405 (N_5405,N_54,N_3688);
and U5406 (N_5406,N_4286,N_185);
or U5407 (N_5407,N_3426,N_234);
nor U5408 (N_5408,N_4548,N_2388);
and U5409 (N_5409,N_3047,N_4675);
xor U5410 (N_5410,N_2333,N_1639);
nor U5411 (N_5411,N_4840,N_1101);
and U5412 (N_5412,N_3850,N_4301);
nand U5413 (N_5413,N_1961,N_1269);
nor U5414 (N_5414,N_2373,N_4148);
nand U5415 (N_5415,N_3789,N_3974);
xnor U5416 (N_5416,N_4636,N_1764);
and U5417 (N_5417,N_2705,N_2178);
or U5418 (N_5418,N_4441,N_3945);
nor U5419 (N_5419,N_2216,N_951);
nor U5420 (N_5420,N_2121,N_13);
and U5421 (N_5421,N_3436,N_184);
nor U5422 (N_5422,N_1911,N_1763);
nor U5423 (N_5423,N_680,N_569);
and U5424 (N_5424,N_4720,N_3358);
and U5425 (N_5425,N_1850,N_3908);
or U5426 (N_5426,N_3734,N_4369);
or U5427 (N_5427,N_2243,N_2679);
nor U5428 (N_5428,N_3329,N_1962);
or U5429 (N_5429,N_1759,N_2509);
nor U5430 (N_5430,N_4165,N_2403);
nor U5431 (N_5431,N_649,N_393);
nand U5432 (N_5432,N_1403,N_495);
nor U5433 (N_5433,N_298,N_597);
or U5434 (N_5434,N_1879,N_2054);
nand U5435 (N_5435,N_2484,N_2083);
or U5436 (N_5436,N_728,N_295);
nand U5437 (N_5437,N_3001,N_3131);
and U5438 (N_5438,N_3594,N_2761);
and U5439 (N_5439,N_4611,N_4353);
nor U5440 (N_5440,N_1884,N_3032);
and U5441 (N_5441,N_4728,N_2786);
and U5442 (N_5442,N_1896,N_2092);
and U5443 (N_5443,N_570,N_1685);
or U5444 (N_5444,N_557,N_1152);
or U5445 (N_5445,N_3220,N_4395);
and U5446 (N_5446,N_4890,N_2280);
nor U5447 (N_5447,N_1777,N_247);
and U5448 (N_5448,N_1516,N_3922);
nand U5449 (N_5449,N_143,N_742);
or U5450 (N_5450,N_3567,N_4003);
nand U5451 (N_5451,N_2704,N_1947);
nand U5452 (N_5452,N_1040,N_216);
nor U5453 (N_5453,N_2356,N_4392);
or U5454 (N_5454,N_2602,N_1527);
or U5455 (N_5455,N_3883,N_1901);
or U5456 (N_5456,N_3727,N_1549);
or U5457 (N_5457,N_1814,N_4325);
nand U5458 (N_5458,N_3196,N_3750);
or U5459 (N_5459,N_2272,N_4849);
or U5460 (N_5460,N_1226,N_1135);
nand U5461 (N_5461,N_560,N_4846);
nand U5462 (N_5462,N_103,N_801);
nor U5463 (N_5463,N_721,N_3565);
and U5464 (N_5464,N_1910,N_4848);
nand U5465 (N_5465,N_1871,N_2246);
nor U5466 (N_5466,N_356,N_1963);
nor U5467 (N_5467,N_4432,N_1249);
nand U5468 (N_5468,N_3592,N_4144);
nor U5469 (N_5469,N_1821,N_889);
and U5470 (N_5470,N_735,N_1574);
nand U5471 (N_5471,N_3487,N_2125);
nand U5472 (N_5472,N_3099,N_3120);
nor U5473 (N_5473,N_1913,N_4818);
or U5474 (N_5474,N_3257,N_2997);
or U5475 (N_5475,N_2215,N_3101);
nand U5476 (N_5476,N_992,N_776);
nor U5477 (N_5477,N_2736,N_2751);
nor U5478 (N_5478,N_197,N_3351);
or U5479 (N_5479,N_2448,N_4245);
nor U5480 (N_5480,N_3656,N_2963);
or U5481 (N_5481,N_1118,N_3449);
nand U5482 (N_5482,N_2454,N_4610);
and U5483 (N_5483,N_1726,N_3095);
nor U5484 (N_5484,N_3083,N_4153);
or U5485 (N_5485,N_2006,N_1768);
nor U5486 (N_5486,N_1796,N_3787);
or U5487 (N_5487,N_4859,N_3856);
or U5488 (N_5488,N_83,N_866);
and U5489 (N_5489,N_656,N_4209);
nand U5490 (N_5490,N_1823,N_3044);
nor U5491 (N_5491,N_2283,N_1123);
or U5492 (N_5492,N_455,N_3796);
and U5493 (N_5493,N_4011,N_1238);
nand U5494 (N_5494,N_2151,N_117);
nor U5495 (N_5495,N_3659,N_2267);
and U5496 (N_5496,N_2979,N_3259);
and U5497 (N_5497,N_4342,N_2422);
nand U5498 (N_5498,N_2463,N_1459);
nand U5499 (N_5499,N_688,N_2756);
nand U5500 (N_5500,N_4667,N_3415);
and U5501 (N_5501,N_1765,N_82);
nand U5502 (N_5502,N_86,N_4647);
nand U5503 (N_5503,N_102,N_3179);
xnor U5504 (N_5504,N_4315,N_669);
nor U5505 (N_5505,N_4289,N_3085);
or U5506 (N_5506,N_1504,N_387);
or U5507 (N_5507,N_4634,N_414);
or U5508 (N_5508,N_4979,N_3706);
nand U5509 (N_5509,N_3295,N_2107);
nand U5510 (N_5510,N_2337,N_147);
and U5511 (N_5511,N_2342,N_2160);
nand U5512 (N_5512,N_2608,N_3452);
nor U5513 (N_5513,N_215,N_3274);
xnor U5514 (N_5514,N_361,N_3137);
xnor U5515 (N_5515,N_685,N_2652);
or U5516 (N_5516,N_3546,N_227);
or U5517 (N_5517,N_2256,N_4814);
and U5518 (N_5518,N_2177,N_4648);
or U5519 (N_5519,N_3964,N_1567);
nor U5520 (N_5520,N_121,N_4762);
nor U5521 (N_5521,N_716,N_2591);
nor U5522 (N_5522,N_1581,N_3728);
nand U5523 (N_5523,N_2959,N_3935);
or U5524 (N_5524,N_4929,N_3880);
nor U5525 (N_5525,N_2817,N_1621);
and U5526 (N_5526,N_377,N_1059);
and U5527 (N_5527,N_2335,N_1045);
nor U5528 (N_5528,N_2628,N_3050);
nand U5529 (N_5529,N_3485,N_859);
or U5530 (N_5530,N_3975,N_1982);
and U5531 (N_5531,N_2707,N_3939);
and U5532 (N_5532,N_1737,N_1007);
or U5533 (N_5533,N_145,N_4226);
and U5534 (N_5534,N_3807,N_4920);
and U5535 (N_5535,N_3744,N_4911);
and U5536 (N_5536,N_871,N_2401);
and U5537 (N_5537,N_2459,N_2573);
or U5538 (N_5538,N_610,N_2623);
nor U5539 (N_5539,N_3015,N_2914);
and U5540 (N_5540,N_2788,N_1062);
xor U5541 (N_5541,N_4633,N_9);
nor U5542 (N_5542,N_3970,N_4925);
and U5543 (N_5543,N_542,N_111);
or U5544 (N_5544,N_44,N_2765);
nand U5545 (N_5545,N_2701,N_3153);
or U5546 (N_5546,N_1976,N_4737);
or U5547 (N_5547,N_2516,N_1840);
or U5548 (N_5548,N_3860,N_1636);
nand U5549 (N_5549,N_2115,N_1695);
and U5550 (N_5550,N_1528,N_4302);
or U5551 (N_5551,N_4048,N_2631);
or U5552 (N_5552,N_4759,N_1468);
nor U5553 (N_5553,N_3341,N_699);
or U5554 (N_5554,N_1676,N_3711);
nand U5555 (N_5555,N_2673,N_467);
nor U5556 (N_5556,N_3671,N_4552);
or U5557 (N_5557,N_3888,N_4099);
or U5558 (N_5558,N_3154,N_3766);
nand U5559 (N_5559,N_2984,N_4739);
and U5560 (N_5560,N_2712,N_43);
or U5561 (N_5561,N_1626,N_4674);
nand U5562 (N_5562,N_4970,N_3460);
and U5563 (N_5563,N_3365,N_199);
nor U5564 (N_5564,N_726,N_1139);
nor U5565 (N_5565,N_629,N_4352);
nand U5566 (N_5566,N_960,N_2088);
nand U5567 (N_5567,N_2040,N_1318);
or U5568 (N_5568,N_2515,N_2816);
or U5569 (N_5569,N_3507,N_2217);
nor U5570 (N_5570,N_4749,N_4520);
or U5571 (N_5571,N_2540,N_3924);
nand U5572 (N_5572,N_611,N_476);
or U5573 (N_5573,N_3996,N_1179);
nand U5574 (N_5574,N_3575,N_1401);
xor U5575 (N_5575,N_2548,N_3804);
and U5576 (N_5576,N_904,N_2352);
or U5577 (N_5577,N_675,N_2347);
nand U5578 (N_5578,N_766,N_2838);
and U5579 (N_5579,N_1917,N_3108);
and U5580 (N_5580,N_3082,N_615);
nand U5581 (N_5581,N_2803,N_2737);
nor U5582 (N_5582,N_3314,N_3012);
or U5583 (N_5583,N_2419,N_4507);
nor U5584 (N_5584,N_3817,N_3566);
nor U5585 (N_5585,N_4875,N_3417);
and U5586 (N_5586,N_1670,N_2052);
or U5587 (N_5587,N_3188,N_206);
and U5588 (N_5588,N_3782,N_800);
nor U5589 (N_5589,N_1886,N_258);
and U5590 (N_5590,N_3304,N_4813);
nand U5591 (N_5591,N_4002,N_225);
nor U5592 (N_5592,N_1109,N_4842);
nor U5593 (N_5593,N_3636,N_4800);
and U5594 (N_5594,N_3553,N_2757);
or U5595 (N_5595,N_2199,N_2461);
and U5596 (N_5596,N_108,N_818);
and U5597 (N_5597,N_3825,N_2794);
and U5598 (N_5598,N_743,N_2122);
or U5599 (N_5599,N_1106,N_2558);
and U5600 (N_5600,N_1806,N_2668);
and U5601 (N_5601,N_2491,N_2496);
nand U5602 (N_5602,N_3506,N_3210);
and U5603 (N_5603,N_1903,N_2474);
nor U5604 (N_5604,N_1172,N_4145);
nand U5605 (N_5605,N_613,N_3502);
or U5606 (N_5606,N_2176,N_2863);
nand U5607 (N_5607,N_162,N_3228);
nor U5608 (N_5608,N_1532,N_278);
or U5609 (N_5609,N_1348,N_644);
nand U5610 (N_5610,N_4220,N_4415);
nand U5611 (N_5611,N_4777,N_4297);
and U5612 (N_5612,N_4939,N_1449);
nor U5613 (N_5613,N_1541,N_999);
and U5614 (N_5614,N_1233,N_457);
or U5615 (N_5615,N_813,N_2826);
and U5616 (N_5616,N_2070,N_481);
nor U5617 (N_5617,N_3118,N_3024);
nand U5618 (N_5618,N_4442,N_4622);
and U5619 (N_5619,N_3928,N_67);
or U5620 (N_5620,N_894,N_4161);
and U5621 (N_5621,N_4752,N_758);
nor U5622 (N_5622,N_1568,N_3703);
or U5623 (N_5623,N_1741,N_107);
nor U5624 (N_5624,N_4879,N_3769);
and U5625 (N_5625,N_2467,N_1192);
nand U5626 (N_5626,N_4828,N_3019);
nand U5627 (N_5627,N_4486,N_1570);
nand U5628 (N_5628,N_4267,N_3458);
and U5629 (N_5629,N_1448,N_2941);
nor U5630 (N_5630,N_153,N_655);
and U5631 (N_5631,N_3191,N_3754);
nand U5632 (N_5632,N_2165,N_1959);
xor U5633 (N_5633,N_3472,N_1444);
nand U5634 (N_5634,N_988,N_1324);
nand U5635 (N_5635,N_4587,N_2339);
nor U5636 (N_5636,N_2501,N_4313);
or U5637 (N_5637,N_3263,N_4340);
nand U5638 (N_5638,N_798,N_1809);
nor U5639 (N_5639,N_149,N_2364);
nor U5640 (N_5640,N_2641,N_4637);
nor U5641 (N_5641,N_1433,N_1807);
or U5642 (N_5642,N_48,N_2399);
and U5643 (N_5643,N_529,N_631);
and U5644 (N_5644,N_3946,N_2451);
or U5645 (N_5645,N_163,N_1960);
and U5646 (N_5646,N_4974,N_1052);
nand U5647 (N_5647,N_907,N_4661);
and U5648 (N_5648,N_4680,N_479);
nor U5649 (N_5649,N_3677,N_3503);
nor U5650 (N_5650,N_4256,N_4565);
or U5651 (N_5651,N_4630,N_3186);
and U5652 (N_5652,N_1606,N_246);
nor U5653 (N_5653,N_3649,N_2381);
nor U5654 (N_5654,N_2079,N_2007);
nand U5655 (N_5655,N_524,N_3480);
and U5656 (N_5656,N_1334,N_2389);
nor U5657 (N_5657,N_759,N_1703);
nand U5658 (N_5658,N_1550,N_1688);
or U5659 (N_5659,N_256,N_3018);
or U5660 (N_5660,N_3696,N_2989);
nand U5661 (N_5661,N_71,N_3951);
nand U5662 (N_5662,N_4487,N_1175);
nand U5663 (N_5663,N_1497,N_1684);
and U5664 (N_5664,N_3570,N_2343);
nor U5665 (N_5665,N_2489,N_150);
and U5666 (N_5666,N_4866,N_2594);
nor U5667 (N_5667,N_4789,N_4560);
nor U5668 (N_5668,N_3054,N_399);
and U5669 (N_5669,N_1155,N_1485);
or U5670 (N_5670,N_2505,N_1027);
nor U5671 (N_5671,N_970,N_4829);
or U5672 (N_5672,N_1285,N_388);
nor U5673 (N_5673,N_815,N_4683);
nand U5674 (N_5674,N_1271,N_1758);
or U5675 (N_5675,N_2962,N_4328);
and U5676 (N_5676,N_4164,N_3826);
or U5677 (N_5677,N_3011,N_1994);
or U5678 (N_5678,N_3170,N_1986);
or U5679 (N_5679,N_3697,N_624);
nor U5680 (N_5680,N_3124,N_1748);
or U5681 (N_5681,N_209,N_2586);
or U5682 (N_5682,N_3926,N_1022);
nand U5683 (N_5683,N_584,N_4566);
nand U5684 (N_5684,N_3042,N_1891);
nor U5685 (N_5685,N_4106,N_548);
or U5686 (N_5686,N_2262,N_128);
or U5687 (N_5687,N_2014,N_3009);
nor U5688 (N_5688,N_3740,N_419);
nor U5689 (N_5689,N_3237,N_1544);
and U5690 (N_5690,N_1257,N_3619);
nor U5691 (N_5691,N_4900,N_3123);
or U5692 (N_5692,N_2783,N_3576);
nor U5693 (N_5693,N_804,N_577);
and U5694 (N_5694,N_587,N_4778);
and U5695 (N_5695,N_1545,N_4397);
and U5696 (N_5696,N_63,N_4766);
or U5697 (N_5697,N_1297,N_1031);
nand U5698 (N_5698,N_390,N_3055);
nor U5699 (N_5699,N_486,N_793);
or U5700 (N_5700,N_2966,N_4390);
and U5701 (N_5701,N_3462,N_2980);
and U5702 (N_5702,N_4378,N_657);
and U5703 (N_5703,N_2806,N_1312);
and U5704 (N_5704,N_4053,N_3737);
and U5705 (N_5705,N_1237,N_4331);
nand U5706 (N_5706,N_1735,N_1125);
or U5707 (N_5707,N_4386,N_770);
nand U5708 (N_5708,N_518,N_3855);
and U5709 (N_5709,N_4090,N_2977);
xor U5710 (N_5710,N_1665,N_1719);
xnor U5711 (N_5711,N_3838,N_2671);
nor U5712 (N_5712,N_3088,N_3867);
nor U5713 (N_5713,N_1043,N_4628);
and U5714 (N_5714,N_552,N_2770);
and U5715 (N_5715,N_2113,N_2257);
and U5716 (N_5716,N_1694,N_1766);
nor U5717 (N_5717,N_4481,N_1955);
nor U5718 (N_5718,N_2541,N_2084);
and U5719 (N_5719,N_3547,N_1478);
or U5720 (N_5720,N_3067,N_4748);
nand U5721 (N_5721,N_1370,N_1868);
nand U5722 (N_5722,N_465,N_2993);
nand U5723 (N_5723,N_4196,N_3362);
nor U5724 (N_5724,N_1013,N_1951);
nor U5725 (N_5725,N_11,N_1218);
nor U5726 (N_5726,N_4104,N_3586);
and U5727 (N_5727,N_4975,N_3070);
nor U5728 (N_5728,N_3031,N_4476);
nor U5729 (N_5729,N_4234,N_690);
nor U5730 (N_5730,N_2739,N_3111);
or U5731 (N_5731,N_3422,N_2224);
nand U5732 (N_5732,N_1278,N_2638);
and U5733 (N_5733,N_966,N_2005);
nor U5734 (N_5734,N_2818,N_1207);
nand U5735 (N_5735,N_169,N_4526);
xor U5736 (N_5736,N_2730,N_2240);
or U5737 (N_5737,N_4931,N_1258);
nand U5738 (N_5738,N_2995,N_3824);
or U5739 (N_5739,N_4827,N_2587);
and U5740 (N_5740,N_1446,N_1341);
or U5741 (N_5741,N_3569,N_4092);
xor U5742 (N_5742,N_619,N_1610);
nor U5743 (N_5743,N_4731,N_4158);
or U5744 (N_5744,N_494,N_338);
nand U5745 (N_5745,N_1255,N_3248);
xor U5746 (N_5746,N_287,N_1105);
or U5747 (N_5747,N_1693,N_1789);
or U5748 (N_5748,N_4469,N_608);
or U5749 (N_5749,N_4293,N_1739);
nand U5750 (N_5750,N_2295,N_2061);
nand U5751 (N_5751,N_658,N_3470);
and U5752 (N_5752,N_3802,N_1034);
nand U5753 (N_5753,N_3539,N_3721);
nor U5754 (N_5754,N_2021,N_1590);
and U5755 (N_5755,N_4532,N_4988);
and U5756 (N_5756,N_3020,N_2385);
nand U5757 (N_5757,N_2436,N_3906);
nand U5758 (N_5758,N_1983,N_2141);
and U5759 (N_5759,N_1895,N_2133);
nand U5760 (N_5760,N_1056,N_2677);
and U5761 (N_5761,N_1929,N_3909);
nor U5762 (N_5762,N_858,N_2625);
or U5763 (N_5763,N_1716,N_1301);
or U5764 (N_5764,N_3585,N_218);
nand U5765 (N_5765,N_2574,N_594);
or U5766 (N_5766,N_3692,N_791);
or U5767 (N_5767,N_17,N_1704);
or U5768 (N_5768,N_4180,N_3907);
and U5769 (N_5769,N_3600,N_4356);
nor U5770 (N_5770,N_1064,N_3495);
or U5771 (N_5771,N_1317,N_3654);
nand U5772 (N_5772,N_180,N_2805);
nand U5773 (N_5773,N_3367,N_4188);
nor U5774 (N_5774,N_413,N_3486);
nand U5775 (N_5775,N_1648,N_1176);
nand U5776 (N_5776,N_4554,N_1714);
xor U5777 (N_5777,N_59,N_1445);
nand U5778 (N_5778,N_1906,N_4782);
nor U5779 (N_5779,N_4291,N_934);
and U5780 (N_5780,N_1121,N_2411);
nand U5781 (N_5781,N_2732,N_1494);
nand U5782 (N_5782,N_778,N_1274);
or U5783 (N_5783,N_4676,N_1760);
or U5784 (N_5784,N_2642,N_3582);
or U5785 (N_5785,N_2192,N_4659);
nand U5786 (N_5786,N_4803,N_3777);
nand U5787 (N_5787,N_872,N_1365);
and U5788 (N_5788,N_4175,N_324);
nor U5789 (N_5789,N_3076,N_4584);
nor U5790 (N_5790,N_2371,N_3057);
and U5791 (N_5791,N_1909,N_3579);
nand U5792 (N_5792,N_4247,N_3138);
nand U5793 (N_5793,N_2056,N_4269);
nor U5794 (N_5794,N_305,N_3645);
nand U5795 (N_5795,N_913,N_1141);
xnor U5796 (N_5796,N_4694,N_2020);
nor U5797 (N_5797,N_4952,N_782);
or U5798 (N_5798,N_3060,N_4631);
or U5799 (N_5799,N_3803,N_3181);
or U5800 (N_5800,N_1094,N_4448);
or U5801 (N_5801,N_4898,N_3901);
nor U5802 (N_5802,N_722,N_214);
and U5803 (N_5803,N_2242,N_25);
or U5804 (N_5804,N_2872,N_4309);
or U5805 (N_5805,N_1263,N_2476);
nor U5806 (N_5806,N_4045,N_1140);
nor U5807 (N_5807,N_3581,N_1097);
and U5808 (N_5808,N_389,N_3174);
or U5809 (N_5809,N_396,N_694);
nor U5810 (N_5810,N_4945,N_909);
or U5811 (N_5811,N_2193,N_3508);
or U5812 (N_5812,N_2791,N_3315);
nor U5813 (N_5813,N_4658,N_2205);
nor U5814 (N_5814,N_2624,N_1854);
or U5815 (N_5815,N_1456,N_3493);
nor U5816 (N_5816,N_1547,N_3262);
and U5817 (N_5817,N_1784,N_1397);
or U5818 (N_5818,N_4038,N_1616);
and U5819 (N_5819,N_1234,N_4453);
or U5820 (N_5820,N_2362,N_3350);
nor U5821 (N_5821,N_1786,N_2723);
and U5822 (N_5822,N_3716,N_3063);
nand U5823 (N_5823,N_3915,N_2445);
or U5824 (N_5824,N_555,N_3115);
or U5825 (N_5825,N_3348,N_3038);
nand U5826 (N_5826,N_4063,N_2375);
nor U5827 (N_5827,N_223,N_3512);
or U5828 (N_5828,N_2923,N_3224);
nor U5829 (N_5829,N_2544,N_411);
or U5830 (N_5830,N_1486,N_2369);
nand U5831 (N_5831,N_1089,N_1425);
nor U5832 (N_5832,N_4229,N_595);
or U5833 (N_5833,N_4211,N_3209);
and U5834 (N_5834,N_635,N_29);
or U5835 (N_5835,N_4823,N_4100);
nor U5836 (N_5836,N_336,N_2710);
nand U5837 (N_5837,N_2498,N_1382);
nand U5838 (N_5838,N_3028,N_1872);
or U5839 (N_5839,N_1316,N_1632);
nor U5840 (N_5840,N_2822,N_4707);
nor U5841 (N_5841,N_294,N_2439);
or U5842 (N_5842,N_4521,N_3819);
or U5843 (N_5843,N_3751,N_1405);
or U5844 (N_5844,N_3783,N_4508);
or U5845 (N_5845,N_573,N_3200);
and U5846 (N_5846,N_3285,N_2650);
and U5847 (N_5847,N_1025,N_881);
or U5848 (N_5848,N_4844,N_2026);
or U5849 (N_5849,N_335,N_4124);
nand U5850 (N_5850,N_617,N_1338);
nor U5851 (N_5851,N_2408,N_3952);
nor U5852 (N_5852,N_2158,N_2038);
nand U5853 (N_5853,N_4204,N_2031);
xnor U5854 (N_5854,N_822,N_2905);
nand U5855 (N_5855,N_1557,N_1818);
nand U5856 (N_5856,N_275,N_3081);
nor U5857 (N_5857,N_2878,N_1283);
and U5858 (N_5858,N_833,N_3286);
and U5859 (N_5859,N_2747,N_3805);
nand U5860 (N_5860,N_2609,N_68);
nor U5861 (N_5861,N_1841,N_835);
or U5862 (N_5862,N_4915,N_3919);
nor U5863 (N_5863,N_3614,N_1864);
xnor U5864 (N_5864,N_2809,N_1831);
and U5865 (N_5865,N_668,N_3201);
and U5866 (N_5866,N_2117,N_2415);
nand U5867 (N_5867,N_1921,N_2190);
xnor U5868 (N_5868,N_513,N_2842);
nor U5869 (N_5869,N_1099,N_1953);
and U5870 (N_5870,N_3427,N_1586);
nor U5871 (N_5871,N_1131,N_97);
and U5872 (N_5872,N_1136,N_148);
and U5873 (N_5873,N_1411,N_1196);
nand U5874 (N_5874,N_1827,N_2983);
nand U5875 (N_5875,N_3823,N_4678);
nand U5876 (N_5876,N_2615,N_2967);
or U5877 (N_5877,N_1867,N_3840);
and U5878 (N_5878,N_4696,N_1335);
nor U5879 (N_5879,N_4558,N_2990);
and U5880 (N_5880,N_903,N_963);
or U5881 (N_5881,N_4222,N_1899);
nor U5882 (N_5882,N_4461,N_4185);
or U5883 (N_5883,N_90,N_2828);
and U5884 (N_5884,N_200,N_3431);
nor U5885 (N_5885,N_4248,N_3355);
and U5886 (N_5886,N_4235,N_57);
nand U5887 (N_5887,N_3324,N_3642);
or U5888 (N_5888,N_1353,N_4522);
nand U5889 (N_5889,N_634,N_3133);
nand U5890 (N_5890,N_3763,N_4880);
and U5891 (N_5891,N_133,N_3726);
and U5892 (N_5892,N_876,N_1775);
or U5893 (N_5893,N_2180,N_2992);
nor U5894 (N_5894,N_1117,N_1157);
or U5895 (N_5895,N_1160,N_4270);
or U5896 (N_5896,N_1385,N_3625);
or U5897 (N_5897,N_4709,N_1950);
nor U5898 (N_5898,N_2834,N_1644);
nor U5899 (N_5899,N_3735,N_4081);
nor U5900 (N_5900,N_3207,N_1667);
or U5901 (N_5901,N_3812,N_748);
nor U5902 (N_5902,N_2074,N_1559);
nor U5903 (N_5903,N_4817,N_1344);
nand U5904 (N_5904,N_2865,N_3616);
or U5905 (N_5905,N_1284,N_4337);
nor U5906 (N_5906,N_1931,N_355);
nand U5907 (N_5907,N_56,N_2559);
and U5908 (N_5908,N_4771,N_2189);
nor U5909 (N_5909,N_1487,N_2493);
or U5910 (N_5910,N_4489,N_2494);
and U5911 (N_5911,N_3155,N_4194);
and U5912 (N_5912,N_4690,N_4947);
and U5913 (N_5913,N_1733,N_4451);
nor U5914 (N_5914,N_4471,N_1465);
nand U5915 (N_5915,N_366,N_4918);
nor U5916 (N_5916,N_983,N_3910);
nand U5917 (N_5917,N_3612,N_2894);
nand U5918 (N_5918,N_3618,N_4938);
or U5919 (N_5919,N_2046,N_4036);
and U5920 (N_5920,N_1054,N_4056);
nor U5921 (N_5921,N_3305,N_4967);
nand U5922 (N_5922,N_4259,N_2098);
nor U5923 (N_5923,N_2321,N_3222);
nor U5924 (N_5924,N_1191,N_3296);
nor U5925 (N_5925,N_605,N_4825);
nor U5926 (N_5926,N_4094,N_2167);
nor U5927 (N_5927,N_4792,N_72);
or U5928 (N_5928,N_4282,N_2);
nor U5929 (N_5929,N_937,N_1077);
and U5930 (N_5930,N_1769,N_475);
or U5931 (N_5931,N_654,N_1474);
or U5932 (N_5932,N_354,N_3068);
nand U5933 (N_5933,N_4433,N_3666);
and U5934 (N_5934,N_4962,N_2595);
xor U5935 (N_5935,N_2655,N_2547);
nand U5936 (N_5936,N_2424,N_1933);
nand U5937 (N_5937,N_2379,N_3559);
nor U5938 (N_5938,N_4635,N_1535);
and U5939 (N_5939,N_2820,N_3317);
or U5940 (N_5940,N_2528,N_3447);
or U5941 (N_5941,N_2597,N_3736);
and U5942 (N_5942,N_1576,N_3448);
nor U5943 (N_5943,N_3662,N_1299);
or U5944 (N_5944,N_236,N_2472);
nand U5945 (N_5945,N_2188,N_1096);
and U5946 (N_5946,N_670,N_70);
and U5947 (N_5947,N_3166,N_434);
nor U5948 (N_5948,N_1049,N_3724);
and U5949 (N_5949,N_1776,N_2186);
nand U5950 (N_5950,N_321,N_3477);
or U5951 (N_5951,N_3545,N_1048);
or U5952 (N_5952,N_2358,N_3933);
and U5953 (N_5953,N_1230,N_1551);
or U5954 (N_5954,N_4251,N_3602);
nand U5955 (N_5955,N_424,N_2175);
nor U5956 (N_5956,N_3264,N_3205);
nand U5957 (N_5957,N_4992,N_736);
nor U5958 (N_5958,N_906,N_3148);
nand U5959 (N_5959,N_3800,N_817);
nor U5960 (N_5960,N_4783,N_4421);
and U5961 (N_5961,N_4541,N_3282);
nand U5962 (N_5962,N_2452,N_3815);
or U5963 (N_5963,N_3005,N_2187);
nand U5964 (N_5964,N_2279,N_3388);
or U5965 (N_5965,N_522,N_4681);
and U5966 (N_5966,N_3483,N_2804);
or U5967 (N_5967,N_313,N_823);
and U5968 (N_5968,N_2248,N_2664);
and U5969 (N_5969,N_3818,N_3145);
and U5970 (N_5970,N_1239,N_3813);
nor U5971 (N_5971,N_796,N_4494);
or U5972 (N_5972,N_307,N_4551);
nor U5973 (N_5973,N_3168,N_2477);
xnor U5974 (N_5974,N_1087,N_4013);
nand U5975 (N_5975,N_1057,N_182);
nor U5976 (N_5976,N_2633,N_1674);
nand U5977 (N_5977,N_1180,N_1319);
nand U5978 (N_5978,N_2886,N_607);
and U5979 (N_5979,N_3925,N_1235);
nand U5980 (N_5980,N_453,N_2883);
or U5981 (N_5981,N_2551,N_640);
or U5982 (N_5982,N_3917,N_2915);
nand U5983 (N_5983,N_916,N_3456);
and U5984 (N_5984,N_3899,N_4300);
and U5985 (N_5985,N_2197,N_697);
nand U5986 (N_5986,N_1536,N_4064);
xor U5987 (N_5987,N_3705,N_2144);
nor U5988 (N_5988,N_2377,N_1490);
or U5989 (N_5989,N_1393,N_4944);
nand U5990 (N_5990,N_1558,N_1024);
nand U5991 (N_5991,N_4819,N_84);
and U5992 (N_5992,N_4496,N_707);
nor U5993 (N_5993,N_1873,N_333);
or U5994 (N_5994,N_3211,N_710);
nor U5995 (N_5995,N_3077,N_2832);
and U5996 (N_5996,N_4391,N_3467);
or U5997 (N_5997,N_1617,N_3184);
and U5998 (N_5998,N_645,N_492);
nand U5999 (N_5999,N_952,N_2755);
or U6000 (N_6000,N_3611,N_676);
nor U6001 (N_6001,N_1366,N_4969);
nand U6002 (N_6002,N_1711,N_1666);
nand U6003 (N_6003,N_423,N_264);
nor U6004 (N_6004,N_2453,N_1129);
or U6005 (N_6005,N_4393,N_3630);
or U6006 (N_6006,N_938,N_2301);
and U6007 (N_6007,N_2260,N_2601);
nor U6008 (N_6008,N_4163,N_1245);
and U6009 (N_6009,N_4802,N_4190);
nand U6010 (N_6010,N_4320,N_4224);
and U6011 (N_6011,N_1984,N_3027);
nor U6012 (N_6012,N_672,N_1201);
and U6013 (N_6013,N_296,N_814);
or U6014 (N_6014,N_65,N_2446);
or U6015 (N_6015,N_4798,N_489);
and U6016 (N_6016,N_621,N_1143);
or U6017 (N_6017,N_3943,N_695);
or U6018 (N_6018,N_1838,N_2281);
nand U6019 (N_6019,N_1525,N_1304);
or U6020 (N_6020,N_1645,N_665);
nand U6021 (N_6021,N_3929,N_785);
nor U6022 (N_6022,N_347,N_3176);
and U6023 (N_6023,N_2091,N_96);
xnor U6024 (N_6024,N_1904,N_3089);
or U6025 (N_6025,N_554,N_4671);
nand U6026 (N_6026,N_1229,N_4029);
and U6027 (N_6027,N_2214,N_3976);
nand U6028 (N_6028,N_1095,N_3732);
nor U6029 (N_6029,N_2840,N_2030);
or U6030 (N_6030,N_1067,N_1602);
or U6031 (N_6031,N_4438,N_1522);
nand U6032 (N_6032,N_417,N_1501);
nand U6033 (N_6033,N_3438,N_2220);
nand U6034 (N_6034,N_3284,N_1571);
or U6035 (N_6035,N_3900,N_4563);
and U6036 (N_6036,N_4780,N_88);
nand U6037 (N_6037,N_1731,N_4430);
nand U6038 (N_6038,N_921,N_885);
nand U6039 (N_6039,N_1609,N_3613);
nand U6040 (N_6040,N_3466,N_3798);
nor U6041 (N_6041,N_1378,N_786);
or U6042 (N_6042,N_2549,N_3558);
or U6043 (N_6043,N_4097,N_965);
nand U6044 (N_6044,N_4534,N_4695);
and U6045 (N_6045,N_2511,N_23);
nand U6046 (N_6046,N_1169,N_1390);
nor U6047 (N_6047,N_3245,N_491);
and U6048 (N_6048,N_2428,N_1509);
or U6049 (N_6049,N_3522,N_1692);
and U6050 (N_6050,N_1655,N_4547);
nand U6051 (N_6051,N_4515,N_173);
nand U6052 (N_6052,N_849,N_1481);
and U6053 (N_6053,N_719,N_2887);
or U6054 (N_6054,N_3795,N_3739);
nor U6055 (N_6055,N_142,N_1781);
and U6056 (N_6056,N_1457,N_1751);
or U6057 (N_6057,N_4474,N_2314);
nand U6058 (N_6058,N_978,N_827);
and U6059 (N_6059,N_3597,N_2368);
or U6060 (N_6060,N_737,N_1114);
nor U6061 (N_6061,N_3275,N_3977);
xor U6062 (N_6062,N_853,N_2132);
or U6063 (N_6063,N_3663,N_3990);
nand U6064 (N_6064,N_2976,N_3599);
nor U6065 (N_6065,N_3185,N_1975);
and U6066 (N_6066,N_3482,N_4924);
and U6067 (N_6067,N_2940,N_4983);
nand U6068 (N_6068,N_3759,N_1280);
nand U6069 (N_6069,N_512,N_932);
or U6070 (N_6070,N_3938,N_1020);
nand U6071 (N_6071,N_729,N_1734);
and U6072 (N_6072,N_1343,N_2432);
nor U6073 (N_6073,N_1594,N_601);
or U6074 (N_6074,N_1681,N_2727);
or U6075 (N_6075,N_2920,N_1675);
nor U6076 (N_6076,N_401,N_1051);
nand U6077 (N_6077,N_170,N_3143);
and U6078 (N_6078,N_1320,N_869);
nand U6079 (N_6079,N_1935,N_2808);
nand U6080 (N_6080,N_948,N_1208);
and U6081 (N_6081,N_1287,N_979);
or U6082 (N_6082,N_2423,N_224);
and U6083 (N_6083,N_196,N_4377);
nand U6084 (N_6084,N_2954,N_3287);
nor U6085 (N_6085,N_3268,N_4111);
or U6086 (N_6086,N_1625,N_1736);
or U6087 (N_6087,N_4223,N_2487);
nor U6088 (N_6088,N_3621,N_132);
nand U6089 (N_6089,N_3319,N_3335);
or U6090 (N_6090,N_463,N_902);
nand U6091 (N_6091,N_1743,N_2210);
and U6092 (N_6092,N_4419,N_4075);
or U6093 (N_6093,N_1442,N_1829);
nor U6094 (N_6094,N_4608,N_4946);
or U6095 (N_6095,N_1210,N_4612);
nor U6096 (N_6096,N_2481,N_821);
and U6097 (N_6097,N_3859,N_2018);
xnor U6098 (N_6098,N_4159,N_3169);
nor U6099 (N_6099,N_3035,N_3420);
nand U6100 (N_6100,N_4119,N_1213);
or U6101 (N_6101,N_1012,N_3419);
nand U6102 (N_6102,N_421,N_4793);
nor U6103 (N_6103,N_4987,N_3713);
and U6104 (N_6104,N_4051,N_3610);
and U6105 (N_6105,N_3167,N_3793);
or U6106 (N_6106,N_2156,N_3911);
and U6107 (N_6107,N_4285,N_1732);
nand U6108 (N_6108,N_4733,N_4125);
and U6109 (N_6109,N_1364,N_1839);
or U6110 (N_6110,N_2365,N_4638);
nor U6111 (N_6111,N_4140,N_1392);
nor U6112 (N_6112,N_3423,N_2907);
and U6113 (N_6113,N_2700,N_3531);
xor U6114 (N_6114,N_1384,N_342);
or U6115 (N_6115,N_2660,N_3058);
nor U6116 (N_6116,N_2434,N_4724);
and U6117 (N_6117,N_3634,N_848);
xnor U6118 (N_6118,N_4973,N_4994);
and U6119 (N_6119,N_4199,N_4443);
or U6120 (N_6120,N_3049,N_4756);
or U6121 (N_6121,N_2630,N_547);
and U6122 (N_6122,N_1691,N_21);
or U6123 (N_6123,N_4429,N_1820);
and U6124 (N_6124,N_4156,N_1779);
or U6125 (N_6125,N_2716,N_395);
nand U6126 (N_6126,N_1349,N_4607);
nand U6127 (N_6127,N_2781,N_4573);
nor U6128 (N_6128,N_188,N_3604);
nor U6129 (N_6129,N_4743,N_1247);
or U6130 (N_6130,N_1597,N_958);
or U6131 (N_6131,N_4881,N_892);
or U6132 (N_6132,N_3383,N_4239);
or U6133 (N_6133,N_3920,N_2427);
or U6134 (N_6134,N_1548,N_3988);
xor U6135 (N_6135,N_2854,N_2998);
nand U6136 (N_6136,N_867,N_2041);
nand U6137 (N_6137,N_136,N_3187);
or U6138 (N_6138,N_1068,N_651);
or U6139 (N_6139,N_2693,N_1534);
nor U6140 (N_6140,N_1272,N_1918);
nand U6141 (N_6141,N_846,N_576);
and U6142 (N_6142,N_1260,N_809);
xnor U6143 (N_6143,N_633,N_3464);
or U6144 (N_6144,N_3129,N_174);
nand U6145 (N_6145,N_3870,N_4147);
or U6146 (N_6146,N_4162,N_4454);
and U6147 (N_6147,N_1336,N_4538);
or U6148 (N_6148,N_1934,N_4268);
nor U6149 (N_6149,N_327,N_3045);
or U6150 (N_6150,N_4257,N_533);
nor U6151 (N_6151,N_781,N_1613);
nand U6152 (N_6152,N_2277,N_3114);
and U6153 (N_6153,N_897,N_308);
or U6154 (N_6154,N_681,N_3918);
or U6155 (N_6155,N_4103,N_4847);
nand U6156 (N_6156,N_156,N_4763);
and U6157 (N_6157,N_2172,N_1810);
nand U6158 (N_6158,N_4277,N_1729);
nand U6159 (N_6159,N_3359,N_92);
or U6160 (N_6160,N_2576,N_3781);
or U6161 (N_6161,N_2825,N_870);
or U6162 (N_6162,N_908,N_1042);
nand U6163 (N_6163,N_4867,N_4978);
and U6164 (N_6164,N_4799,N_1170);
and U6165 (N_6165,N_4624,N_3755);
or U6166 (N_6166,N_1252,N_4298);
and U6167 (N_6167,N_750,N_3999);
or U6168 (N_6168,N_4919,N_2603);
nor U6169 (N_6169,N_435,N_261);
and U6170 (N_6170,N_3704,N_1174);
nand U6171 (N_6171,N_1728,N_3834);
or U6172 (N_6172,N_3794,N_87);
nand U6173 (N_6173,N_3239,N_1660);
nor U6174 (N_6174,N_3841,N_4027);
nor U6175 (N_6175,N_4444,N_1718);
or U6176 (N_6176,N_4784,N_2605);
and U6177 (N_6177,N_3249,N_830);
and U6178 (N_6178,N_4606,N_647);
and U6179 (N_6179,N_2670,N_3773);
nand U6180 (N_6180,N_4512,N_3965);
or U6181 (N_6181,N_1944,N_4462);
or U6182 (N_6182,N_2168,N_3061);
and U6183 (N_6183,N_720,N_3624);
nor U6184 (N_6184,N_2311,N_3474);
and U6185 (N_6185,N_4601,N_1104);
nand U6186 (N_6186,N_1757,N_1937);
or U6187 (N_6187,N_2813,N_4643);
nor U6188 (N_6188,N_3519,N_230);
nand U6189 (N_6189,N_3514,N_1954);
nand U6190 (N_6190,N_4830,N_1254);
nand U6191 (N_6191,N_1754,N_4178);
nor U6192 (N_6192,N_4999,N_2093);
xor U6193 (N_6193,N_2049,N_363);
nor U6194 (N_6194,N_3748,N_755);
and U6195 (N_6195,N_3279,N_783);
or U6196 (N_6196,N_4942,N_3303);
or U6197 (N_6197,N_3622,N_2684);
or U6198 (N_6198,N_4394,N_898);
nand U6199 (N_6199,N_1091,N_2526);
nor U6200 (N_6200,N_579,N_1787);
and U6201 (N_6201,N_3142,N_497);
or U6202 (N_6202,N_4061,N_3008);
xor U6203 (N_6203,N_3407,N_588);
and U6204 (N_6204,N_159,N_600);
nand U6205 (N_6205,N_1584,N_368);
or U6206 (N_6206,N_2510,N_888);
nand U6207 (N_6207,N_2228,N_3580);
and U6208 (N_6208,N_4102,N_3203);
and U6209 (N_6209,N_3389,N_3764);
or U6210 (N_6210,N_1890,N_279);
nor U6211 (N_6211,N_1050,N_350);
and U6212 (N_6212,N_339,N_1742);
nor U6213 (N_6213,N_4853,N_408);
nor U6214 (N_6214,N_2767,N_1914);
and U6215 (N_6215,N_2499,N_3532);
or U6216 (N_6216,N_1791,N_344);
or U6217 (N_6217,N_4117,N_3097);
xor U6218 (N_6218,N_2520,N_3344);
nor U6219 (N_6219,N_1154,N_482);
nor U6220 (N_6220,N_772,N_2386);
nor U6221 (N_6221,N_2932,N_928);
nor U6222 (N_6222,N_243,N_1790);
nor U6223 (N_6223,N_2546,N_3471);
nor U6224 (N_6224,N_183,N_4399);
and U6225 (N_6225,N_3003,N_357);
and U6226 (N_6226,N_3144,N_3809);
nor U6227 (N_6227,N_1115,N_3664);
nor U6228 (N_6228,N_99,N_2956);
and U6229 (N_6229,N_704,N_1098);
or U6230 (N_6230,N_4350,N_2611);
nand U6231 (N_6231,N_160,N_3513);
and U6232 (N_6232,N_1389,N_525);
nor U6233 (N_6233,N_4413,N_3316);
nor U6234 (N_6234,N_3930,N_420);
nand U6235 (N_6235,N_144,N_1046);
nand U6236 (N_6236,N_1822,N_4951);
and U6237 (N_6237,N_583,N_3430);
nor U6238 (N_6238,N_1124,N_1892);
and U6239 (N_6239,N_2157,N_1346);
and U6240 (N_6240,N_2397,N_4303);
and U6241 (N_6241,N_79,N_646);
and U6242 (N_6242,N_3300,N_2917);
or U6243 (N_6243,N_3992,N_3895);
nand U6244 (N_6244,N_3942,N_3865);
nand U6245 (N_6245,N_4592,N_1863);
nor U6246 (N_6246,N_4791,N_4354);
nand U6247 (N_6247,N_2579,N_652);
nand U6248 (N_6248,N_124,N_4098);
or U6249 (N_6249,N_1969,N_2285);
nand U6250 (N_6250,N_228,N_4120);
nor U6251 (N_6251,N_1725,N_3864);
nor U6252 (N_6252,N_1859,N_915);
or U6253 (N_6253,N_1253,N_806);
nor U6254 (N_6254,N_477,N_3216);
nand U6255 (N_6255,N_3799,N_1120);
and U6256 (N_6256,N_1467,N_4664);
or U6257 (N_6257,N_2801,N_1897);
or U6258 (N_6258,N_0,N_3607);
or U6259 (N_6259,N_2972,N_1217);
or U6260 (N_6260,N_2807,N_3573);
nand U6261 (N_6261,N_3852,N_2457);
nor U6262 (N_6262,N_1205,N_2482);
nor U6263 (N_6263,N_2748,N_3439);
nor U6264 (N_6264,N_1083,N_1178);
nand U6265 (N_6265,N_3403,N_4492);
xnor U6266 (N_6266,N_485,N_4860);
nor U6267 (N_6267,N_4768,N_536);
and U6268 (N_6268,N_2470,N_4632);
or U6269 (N_6269,N_283,N_4570);
nor U6270 (N_6270,N_1480,N_3667);
and U6271 (N_6271,N_3261,N_4718);
and U6272 (N_6272,N_3714,N_1502);
and U6273 (N_6273,N_2095,N_2728);
and U6274 (N_6274,N_1227,N_2036);
and U6275 (N_6275,N_239,N_784);
nor U6276 (N_6276,N_4781,N_2080);
nor U6277 (N_6277,N_4166,N_1503);
or U6278 (N_6278,N_1722,N_4294);
nand U6279 (N_6279,N_4232,N_4663);
nand U6280 (N_6280,N_4116,N_155);
nor U6281 (N_6281,N_3451,N_4909);
and U6282 (N_6282,N_2722,N_826);
nand U6283 (N_6283,N_1585,N_987);
or U6284 (N_6284,N_1321,N_808);
nand U6285 (N_6285,N_2085,N_3198);
nor U6286 (N_6286,N_3687,N_768);
or U6287 (N_6287,N_3768,N_4321);
nand U6288 (N_6288,N_2785,N_930);
or U6289 (N_6289,N_3443,N_1019);
nor U6290 (N_6290,N_2961,N_4943);
nor U6291 (N_6291,N_1127,N_3258);
and U6292 (N_6292,N_3465,N_2338);
nor U6293 (N_6293,N_4578,N_3206);
and U6294 (N_6294,N_2483,N_1452);
or U6295 (N_6295,N_2148,N_358);
and U6296 (N_6296,N_3958,N_4794);
nand U6297 (N_6297,N_4210,N_1792);
nor U6298 (N_6298,N_3916,N_3102);
xnor U6299 (N_6299,N_3306,N_771);
or U6300 (N_6300,N_222,N_840);
or U6301 (N_6301,N_1952,N_1654);
or U6302 (N_6302,N_666,N_126);
xnor U6303 (N_6303,N_2024,N_4183);
and U6304 (N_6304,N_4761,N_4697);
nand U6305 (N_6305,N_251,N_4998);
and U6306 (N_6306,N_747,N_1858);
nor U6307 (N_6307,N_1432,N_391);
nand U6308 (N_6308,N_3183,N_1618);
nand U6309 (N_6309,N_4832,N_4482);
or U6310 (N_6310,N_2076,N_4882);
nand U6311 (N_6311,N_2359,N_2367);
or U6312 (N_6312,N_4389,N_312);
and U6313 (N_6313,N_4646,N_943);
and U6314 (N_6314,N_47,N_2512);
or U6315 (N_6315,N_109,N_392);
and U6316 (N_6316,N_4620,N_4189);
and U6317 (N_6317,N_4233,N_2746);
and U6318 (N_6318,N_4333,N_4208);
or U6319 (N_6319,N_2620,N_4824);
nor U6320 (N_6320,N_1167,N_3247);
or U6321 (N_6321,N_596,N_2800);
xor U6322 (N_6322,N_2572,N_3125);
and U6323 (N_6323,N_3979,N_4472);
nand U6324 (N_6324,N_1599,N_2814);
nor U6325 (N_6325,N_371,N_3158);
and U6326 (N_6326,N_381,N_2291);
nor U6327 (N_6327,N_3874,N_4575);
nor U6328 (N_6328,N_2968,N_1361);
nor U6329 (N_6329,N_3292,N_2409);
nor U6330 (N_6330,N_2869,N_4841);
nor U6331 (N_6331,N_693,N_2057);
or U6332 (N_6332,N_112,N_3550);
or U6333 (N_6333,N_328,N_4738);
nor U6334 (N_6334,N_4024,N_1404);
nand U6335 (N_6335,N_514,N_4186);
and U6336 (N_6336,N_436,N_1438);
nor U6337 (N_6337,N_1744,N_4016);
nor U6338 (N_6338,N_2468,N_3455);
and U6339 (N_6339,N_4041,N_1159);
or U6340 (N_6340,N_1600,N_4131);
nand U6341 (N_6341,N_3881,N_3854);
or U6342 (N_6342,N_386,N_1579);
xor U6343 (N_6343,N_2174,N_74);
and U6344 (N_6344,N_1690,N_3147);
and U6345 (N_6345,N_4458,N_2545);
or U6346 (N_6346,N_1797,N_2987);
and U6347 (N_6347,N_450,N_4398);
and U6348 (N_6348,N_1647,N_1635);
or U6349 (N_6349,N_1866,N_114);
and U6350 (N_6350,N_1848,N_2719);
nand U6351 (N_6351,N_4237,N_1603);
or U6352 (N_6352,N_630,N_1785);
nand U6353 (N_6353,N_545,N_311);
or U6354 (N_6354,N_3858,N_3891);
nand U6355 (N_6355,N_4668,N_3676);
or U6356 (N_6356,N_4540,N_4642);
and U6357 (N_6357,N_2928,N_3556);
and U6358 (N_6358,N_2330,N_1073);
nand U6359 (N_6359,N_1889,N_4660);
nand U6360 (N_6360,N_3563,N_2042);
nand U6361 (N_6361,N_4411,N_2284);
and U6362 (N_6362,N_3475,N_3217);
and U6363 (N_6363,N_24,N_2185);
nor U6364 (N_6364,N_235,N_120);
nand U6365 (N_6365,N_1883,N_723);
and U6366 (N_6366,N_438,N_4949);
nor U6367 (N_6367,N_3719,N_4790);
and U6368 (N_6368,N_4527,N_325);
nand U6369 (N_6369,N_4238,N_4273);
nand U6370 (N_6370,N_4854,N_4219);
or U6371 (N_6371,N_2253,N_1151);
nand U6372 (N_6372,N_2208,N_4202);
or U6373 (N_6373,N_2827,N_745);
or U6374 (N_6374,N_2331,N_4626);
nand U6375 (N_6375,N_4993,N_201);
and U6376 (N_6376,N_4753,N_1709);
or U6377 (N_6377,N_2147,N_369);
nand U6378 (N_6378,N_4307,N_28);
nand U6379 (N_6379,N_4324,N_3080);
or U6380 (N_6380,N_1637,N_2245);
or U6381 (N_6381,N_3141,N_2207);
nand U6382 (N_6382,N_895,N_3779);
and U6383 (N_6383,N_905,N_3801);
or U6384 (N_6384,N_1293,N_1958);
xnor U6385 (N_6385,N_349,N_3036);
and U6386 (N_6386,N_4810,N_1396);
and U6387 (N_6387,N_4425,N_2536);
or U6388 (N_6388,N_3694,N_3591);
nor U6389 (N_6389,N_2729,N_1507);
or U6390 (N_6390,N_2944,N_2161);
xnor U6391 (N_6391,N_3742,N_2724);
and U6392 (N_6392,N_1329,N_1266);
nand U6393 (N_6393,N_1060,N_3822);
nor U6394 (N_6394,N_2507,N_3637);
and U6395 (N_6395,N_1296,N_1461);
or U6396 (N_6396,N_1298,N_4806);
nand U6397 (N_6397,N_1500,N_2326);
or U6398 (N_6398,N_1069,N_1506);
nor U6399 (N_6399,N_1627,N_3898);
or U6400 (N_6400,N_2426,N_2435);
or U6401 (N_6401,N_4044,N_2906);
or U6402 (N_6402,N_1638,N_380);
nor U6403 (N_6403,N_1116,N_4035);
or U6404 (N_6404,N_1753,N_42);
nand U6405 (N_6405,N_2261,N_4703);
nand U6406 (N_6406,N_2011,N_4318);
and U6407 (N_6407,N_1055,N_4304);
nand U6408 (N_6408,N_3022,N_787);
or U6409 (N_6409,N_1119,N_4195);
nor U6410 (N_6410,N_3775,N_1771);
nand U6411 (N_6411,N_2815,N_2497);
and U6412 (N_6412,N_4976,N_4905);
or U6413 (N_6413,N_3002,N_2683);
and U6414 (N_6414,N_3260,N_1643);
or U6415 (N_6415,N_2678,N_1679);
nand U6416 (N_6416,N_4621,N_663);
and U6417 (N_6417,N_1491,N_3957);
nor U6418 (N_6418,N_1150,N_2738);
and U6419 (N_6419,N_4523,N_309);
nor U6420 (N_6420,N_4129,N_168);
or U6421 (N_6421,N_2862,N_4597);
or U6422 (N_6422,N_2821,N_1161);
and U6423 (N_6423,N_1483,N_4296);
nor U6424 (N_6424,N_883,N_3428);
nor U6425 (N_6425,N_1355,N_2514);
nor U6426 (N_6426,N_3767,N_2255);
xnor U6427 (N_6427,N_3309,N_1798);
and U6428 (N_6428,N_2898,N_291);
and U6429 (N_6429,N_2674,N_2345);
and U6430 (N_6430,N_662,N_3312);
and U6431 (N_6431,N_2970,N_3523);
nand U6432 (N_6432,N_3290,N_3620);
or U6433 (N_6433,N_3110,N_2206);
and U6434 (N_6434,N_1537,N_2444);
and U6435 (N_6435,N_231,N_2259);
nor U6436 (N_6436,N_158,N_4123);
and U6437 (N_6437,N_3760,N_466);
and U6438 (N_6438,N_1988,N_3331);
nand U6439 (N_6439,N_3134,N_811);
nand U6440 (N_6440,N_2734,N_2012);
nor U6441 (N_6441,N_1555,N_345);
or U6442 (N_6442,N_4883,N_1186);
nand U6443 (N_6443,N_3453,N_2860);
nor U6444 (N_6444,N_4723,N_2644);
nor U6445 (N_6445,N_1998,N_799);
nand U6446 (N_6446,N_4940,N_383);
and U6447 (N_6447,N_3835,N_925);
nand U6448 (N_6448,N_4114,N_300);
nand U6449 (N_6449,N_842,N_4937);
or U6450 (N_6450,N_4958,N_1755);
or U6451 (N_6451,N_2798,N_2733);
and U6452 (N_6452,N_2058,N_31);
nor U6453 (N_6453,N_3969,N_3375);
and U6454 (N_6454,N_1653,N_2953);
or U6455 (N_6455,N_3214,N_4241);
and U6456 (N_6456,N_844,N_896);
or U6457 (N_6457,N_250,N_857);
and U6458 (N_6458,N_4525,N_4716);
xnor U6459 (N_6459,N_4133,N_1900);
or U6460 (N_6460,N_3814,N_1715);
nand U6461 (N_6461,N_4031,N_1942);
nand U6462 (N_6462,N_4279,N_4625);
nand U6463 (N_6463,N_4594,N_3227);
and U6464 (N_6464,N_718,N_3433);
and U6465 (N_6465,N_2051,N_4941);
and U6466 (N_6466,N_4672,N_2233);
or U6467 (N_6467,N_2696,N_1427);
or U6468 (N_6468,N_277,N_4142);
and U6469 (N_6469,N_1357,N_4546);
and U6470 (N_6470,N_3385,N_1383);
or U6471 (N_6471,N_2221,N_838);
nor U6472 (N_6472,N_712,N_3847);
and U6473 (N_6473,N_373,N_1783);
nor U6474 (N_6474,N_4754,N_893);
or U6475 (N_6475,N_2695,N_3691);
and U6476 (N_6476,N_2028,N_431);
or U6477 (N_6477,N_1372,N_4478);
nor U6478 (N_6478,N_3492,N_2275);
and U6479 (N_6479,N_1799,N_4152);
and U6480 (N_6480,N_4228,N_4264);
nor U6481 (N_6481,N_3090,N_3778);
xor U6482 (N_6482,N_1912,N_4446);
and U6483 (N_6483,N_3256,N_2173);
and U6484 (N_6484,N_346,N_2223);
and U6485 (N_6485,N_3100,N_526);
or U6486 (N_6486,N_3690,N_2839);
nand U6487 (N_6487,N_1469,N_1402);
nor U6488 (N_6488,N_1275,N_3772);
nand U6489 (N_6489,N_4861,N_3413);
and U6490 (N_6490,N_4459,N_1713);
nor U6491 (N_6491,N_4529,N_4215);
nor U6492 (N_6492,N_873,N_2874);
nor U6493 (N_6493,N_3192,N_85);
and U6494 (N_6494,N_2584,N_4896);
or U6495 (N_6495,N_3463,N_3361);
or U6496 (N_6496,N_1081,N_4376);
or U6497 (N_6497,N_4910,N_3162);
nand U6498 (N_6498,N_3530,N_1649);
and U6499 (N_6499,N_1422,N_2929);
or U6500 (N_6500,N_4275,N_3877);
and U6501 (N_6501,N_2680,N_1359);
and U6502 (N_6502,N_3729,N_2557);
or U6503 (N_6503,N_3966,N_1458);
nand U6504 (N_6504,N_472,N_4535);
or U6505 (N_6505,N_3827,N_2666);
and U6506 (N_6506,N_274,N_1971);
nand U6507 (N_6507,N_765,N_276);
nand U6508 (N_6508,N_2637,N_532);
nand U6509 (N_6509,N_3197,N_1499);
nand U6510 (N_6510,N_4656,N_1428);
nand U6511 (N_6511,N_1451,N_4855);
nor U6512 (N_6512,N_1633,N_1706);
nand U6513 (N_6513,N_3564,N_1575);
and U6514 (N_6514,N_4593,N_1946);
and U6515 (N_6515,N_4913,N_3052);
nand U6516 (N_6516,N_847,N_2916);
or U6517 (N_6517,N_1847,N_1880);
or U6518 (N_6518,N_4420,N_2981);
or U6519 (N_6519,N_1065,N_1212);
nand U6520 (N_6520,N_4473,N_4290);
nand U6521 (N_6521,N_2772,N_3745);
nor U6522 (N_6522,N_272,N_4057);
and U6523 (N_6523,N_113,N_4348);
or U6524 (N_6524,N_880,N_3034);
and U6525 (N_6525,N_4046,N_1028);
nand U6526 (N_6526,N_1696,N_38);
or U6527 (N_6527,N_3444,N_3527);
nor U6528 (N_6528,N_1805,N_3025);
nand U6529 (N_6529,N_1857,N_2486);
or U6530 (N_6530,N_1938,N_2831);
and U6531 (N_6531,N_1342,N_701);
nand U6532 (N_6532,N_8,N_2116);
and U6533 (N_6533,N_2060,N_1330);
nand U6534 (N_6534,N_757,N_3072);
and U6535 (N_6535,N_4322,N_4240);
and U6536 (N_6536,N_506,N_4569);
nor U6537 (N_6537,N_175,N_3069);
or U6538 (N_6538,N_4207,N_1195);
and U6539 (N_6539,N_4491,N_165);
and U6540 (N_6540,N_4533,N_3171);
or U6541 (N_6541,N_2762,N_1852);
or U6542 (N_6542,N_49,N_692);
and U6543 (N_6543,N_1523,N_4961);
and U6544 (N_6544,N_3792,N_2269);
or U6545 (N_6545,N_3059,N_2851);
or U6546 (N_6546,N_1082,N_1193);
nand U6547 (N_6547,N_2640,N_1286);
nand U6548 (N_6548,N_4808,N_868);
and U6549 (N_6549,N_775,N_4086);
nor U6550 (N_6550,N_829,N_317);
and U6551 (N_6551,N_2896,N_1072);
nand U6552 (N_6552,N_4524,N_1489);
nand U6553 (N_6553,N_691,N_4684);
and U6554 (N_6554,N_1995,N_2166);
nor U6555 (N_6555,N_189,N_865);
nor U6556 (N_6556,N_4497,N_1707);
or U6557 (N_6557,N_1001,N_1762);
nand U6558 (N_6558,N_2885,N_824);
nor U6559 (N_6559,N_1972,N_3281);
xor U6560 (N_6560,N_756,N_4452);
and U6561 (N_6561,N_1770,N_1698);
nor U6562 (N_6562,N_2590,N_1265);
and U6563 (N_6563,N_3525,N_1974);
and U6564 (N_6564,N_2163,N_2908);
nand U6565 (N_6565,N_2425,N_4539);
nor U6566 (N_6566,N_3377,N_964);
and U6567 (N_6567,N_664,N_3294);
nand U6568 (N_6568,N_2032,N_3821);
nand U6569 (N_6569,N_2273,N_3369);
nor U6570 (N_6570,N_4138,N_2429);
nor U6571 (N_6571,N_129,N_2523);
or U6572 (N_6572,N_1243,N_1622);
or U6573 (N_6573,N_4288,N_4701);
or U6574 (N_6574,N_439,N_3963);
nor U6575 (N_6575,N_2581,N_4370);
nor U6576 (N_6576,N_444,N_4263);
nand U6577 (N_6577,N_382,N_2811);
and U6578 (N_6578,N_3232,N_4897);
and U6579 (N_6579,N_2114,N_4230);
or U6580 (N_6580,N_3328,N_270);
or U6581 (N_6581,N_733,N_900);
or U6582 (N_6582,N_3408,N_1307);
or U6583 (N_6583,N_1074,N_58);
and U6584 (N_6584,N_2043,N_1225);
nor U6585 (N_6585,N_1413,N_1746);
nand U6586 (N_6586,N_4901,N_2181);
and U6587 (N_6587,N_4699,N_886);
and U6588 (N_6588,N_1290,N_2656);
and U6589 (N_6589,N_2900,N_3549);
and U6590 (N_6590,N_374,N_3689);
and U6591 (N_6591,N_2323,N_3828);
or U6592 (N_6592,N_3372,N_16);
nand U6593 (N_6593,N_500,N_326);
or U6594 (N_6594,N_14,N_4191);
and U6595 (N_6595,N_4465,N_4603);
nand U6596 (N_6596,N_1011,N_1851);
nand U6597 (N_6597,N_1111,N_4868);
nor U6598 (N_6598,N_4242,N_3693);
and U6599 (N_6599,N_3557,N_406);
xnor U6600 (N_6600,N_4710,N_4617);
and U6601 (N_6601,N_877,N_4564);
nand U6602 (N_6602,N_3882,N_802);
and U6603 (N_6603,N_4184,N_4227);
or U6604 (N_6604,N_2731,N_1292);
nor U6605 (N_6605,N_2383,N_4590);
xnor U6606 (N_6606,N_1350,N_4589);
nor U6607 (N_6607,N_540,N_4972);
nand U6608 (N_6608,N_1566,N_177);
nor U6609 (N_6609,N_998,N_3873);
nor U6610 (N_6610,N_3846,N_2354);
nand U6611 (N_6611,N_1197,N_3366);
or U6612 (N_6612,N_3113,N_1203);
nor U6613 (N_6613,N_2065,N_2023);
nor U6614 (N_6614,N_3536,N_2612);
nor U6615 (N_6615,N_3241,N_969);
nand U6616 (N_6616,N_3280,N_4422);
and U6617 (N_6617,N_4623,N_4640);
nor U6618 (N_6618,N_1017,N_1607);
and U6619 (N_6619,N_1580,N_1005);
nor U6620 (N_6620,N_4040,N_1730);
or U6621 (N_6621,N_4401,N_3505);
nor U6622 (N_6622,N_2155,N_3832);
or U6623 (N_6623,N_1276,N_2282);
and U6624 (N_6624,N_1246,N_4067);
and U6625 (N_6625,N_323,N_1926);
and U6626 (N_6626,N_1834,N_4688);
or U6627 (N_6627,N_2577,N_4284);
nor U6628 (N_6628,N_2034,N_1070);
or U6629 (N_6629,N_1874,N_3178);
nor U6630 (N_6630,N_684,N_1569);
nand U6631 (N_6631,N_4651,N_4310);
nor U6632 (N_6632,N_2241,N_2789);
or U6633 (N_6633,N_1454,N_3298);
or U6634 (N_6634,N_1531,N_2899);
nor U6635 (N_6635,N_3357,N_914);
or U6636 (N_6636,N_348,N_1583);
or U6637 (N_6637,N_2303,N_2965);
or U6638 (N_6638,N_2414,N_2753);
or U6639 (N_6639,N_2396,N_73);
or U6640 (N_6640,N_2714,N_2810);
nor U6641 (N_6641,N_4069,N_404);
nand U6642 (N_6642,N_1387,N_2934);
nand U6643 (N_6643,N_511,N_2232);
nor U6644 (N_6644,N_462,N_3390);
nand U6645 (N_6645,N_3510,N_2320);
nor U6646 (N_6646,N_1992,N_4732);
nand U6647 (N_6647,N_3488,N_4863);
nor U6648 (N_6648,N_977,N_1888);
nand U6649 (N_6649,N_2142,N_461);
nor U6650 (N_6650,N_940,N_2502);
nand U6651 (N_6651,N_2913,N_648);
and U6652 (N_6652,N_763,N_957);
nand U6653 (N_6653,N_1455,N_1678);
nand U6654 (N_6654,N_3743,N_4602);
and U6655 (N_6655,N_3774,N_4511);
nand U6656 (N_6656,N_2462,N_2348);
or U6657 (N_6657,N_2891,N_1166);
or U6658 (N_6658,N_4801,N_244);
and U6659 (N_6659,N_2986,N_4874);
or U6660 (N_6660,N_198,N_2027);
and U6661 (N_6661,N_2258,N_677);
nor U6662 (N_6662,N_2398,N_3747);
nor U6663 (N_6663,N_4236,N_427);
nand U6664 (N_6664,N_2227,N_2164);
nand U6665 (N_6665,N_4347,N_1437);
nor U6666 (N_6666,N_3504,N_4498);
and U6667 (N_6667,N_2799,N_171);
nand U6668 (N_6668,N_717,N_2618);
or U6669 (N_6669,N_2471,N_1708);
and U6670 (N_6670,N_861,N_4435);
xor U6671 (N_6671,N_4821,N_2308);
nand U6672 (N_6672,N_1429,N_3479);
nand U6673 (N_6673,N_4323,N_4691);
or U6674 (N_6674,N_4052,N_1122);
or U6675 (N_6675,N_2310,N_2055);
nor U6676 (N_6676,N_3791,N_530);
nand U6677 (N_6677,N_1628,N_4568);
nand U6678 (N_6678,N_3518,N_1920);
nor U6679 (N_6679,N_2196,N_2309);
nor U6680 (N_6680,N_1313,N_616);
or U6681 (N_6681,N_2534,N_976);
nand U6682 (N_6682,N_1273,N_4869);
and U6683 (N_6683,N_4666,N_4586);
or U6684 (N_6684,N_4772,N_1782);
xor U6685 (N_6685,N_3578,N_3236);
or U6686 (N_6686,N_1039,N_451);
or U6687 (N_6687,N_2123,N_62);
or U6688 (N_6688,N_4682,N_4928);
nand U6689 (N_6689,N_3251,N_242);
or U6690 (N_6690,N_4181,N_4639);
nand U6691 (N_6691,N_3698,N_917);
and U6692 (N_6692,N_204,N_4026);
nor U6693 (N_6693,N_2957,N_1004);
and U6694 (N_6694,N_4345,N_3336);
or U6695 (N_6695,N_1288,N_1990);
nor U6696 (N_6696,N_1611,N_3163);
nor U6697 (N_6697,N_2571,N_262);
xor U6698 (N_6698,N_273,N_4702);
nand U6699 (N_6699,N_4244,N_119);
or U6700 (N_6700,N_3409,N_3524);
or U6701 (N_6701,N_3810,N_1595);
or U6702 (N_6702,N_508,N_2402);
xnor U6703 (N_6703,N_3325,N_2882);
or U6704 (N_6704,N_2450,N_1250);
nor U6705 (N_6705,N_534,N_269);
nor U6706 (N_6706,N_4070,N_3489);
nand U6707 (N_6707,N_3875,N_2568);
nor U6708 (N_6708,N_4679,N_1939);
and U6709 (N_6709,N_2893,N_2111);
nor U6710 (N_6710,N_1426,N_632);
and U6711 (N_6711,N_850,N_3609);
and U6712 (N_6712,N_4499,N_3404);
or U6713 (N_6713,N_2754,N_5);
nor U6714 (N_6714,N_447,N_2580);
nor U6715 (N_6715,N_2697,N_226);
or U6716 (N_6716,N_3393,N_3590);
and U6717 (N_6717,N_1345,N_2875);
or U6718 (N_6718,N_4405,N_4025);
or U6719 (N_6719,N_2449,N_1090);
and U6720 (N_6720,N_3273,N_4734);
or U6721 (N_6721,N_3862,N_1553);
and U6722 (N_6722,N_3311,N_4074);
nand U6723 (N_6723,N_266,N_2930);
or U6724 (N_6724,N_3103,N_4380);
nand U6725 (N_6725,N_1198,N_4965);
and U6726 (N_6726,N_4885,N_3868);
and U6727 (N_6727,N_3459,N_4330);
nand U6728 (N_6728,N_2212,N_4964);
nor U6729 (N_6729,N_1376,N_2170);
or U6730 (N_6730,N_46,N_4221);
and U6731 (N_6731,N_1185,N_4115);
nor U6732 (N_6732,N_3212,N_2346);
nor U6733 (N_6733,N_2234,N_4955);
nor U6734 (N_6734,N_1264,N_3160);
nand U6735 (N_6735,N_3842,N_4431);
nor U6736 (N_6736,N_1752,N_2495);
or U6737 (N_6737,N_3476,N_2895);
or U6738 (N_6738,N_2858,N_2382);
or U6739 (N_6739,N_1659,N_4820);
or U6740 (N_6740,N_1811,N_1424);
nand U6741 (N_6741,N_2336,N_1309);
nand U6742 (N_6742,N_1508,N_3720);
and U6743 (N_6743,N_1956,N_4711);
nor U6744 (N_6744,N_2289,N_3402);
nor U6745 (N_6745,N_2016,N_1702);
nor U6746 (N_6746,N_1967,N_1492);
nor U6747 (N_6747,N_141,N_2393);
nand U6748 (N_6748,N_4893,N_3334);
nor U6749 (N_6749,N_3884,N_3071);
and U6750 (N_6750,N_98,N_3913);
nor U6751 (N_6751,N_2857,N_901);
nand U6752 (N_6752,N_543,N_968);
nor U6753 (N_6753,N_2458,N_4670);
nor U6754 (N_6754,N_3893,N_1608);
nand U6755 (N_6755,N_2127,N_4862);
nor U6756 (N_6756,N_384,N_2412);
nand U6757 (N_6757,N_1826,N_1588);
or U6758 (N_6758,N_1705,N_1861);
or U6759 (N_6759,N_2153,N_4981);
and U6760 (N_6760,N_3454,N_3332);
nor U6761 (N_6761,N_1289,N_839);
or U6762 (N_6762,N_1664,N_1518);
nand U6763 (N_6763,N_678,N_1876);
or U6764 (N_6764,N_3555,N_26);
nand U6765 (N_6765,N_3989,N_1837);
and U6766 (N_6766,N_1828,N_1168);
nand U6767 (N_6767,N_4506,N_1587);
or U6768 (N_6768,N_3343,N_3242);
and U6769 (N_6769,N_2793,N_4618);
nor U6770 (N_6770,N_3308,N_4960);
nor U6771 (N_6771,N_3074,N_4410);
and U6772 (N_6772,N_1519,N_4402);
nor U6773 (N_6773,N_2773,N_4956);
or U6774 (N_6774,N_3998,N_3021);
nor U6775 (N_6775,N_4837,N_2565);
or U6776 (N_6776,N_3469,N_874);
and U6777 (N_6777,N_2527,N_2937);
and U6778 (N_6778,N_2881,N_622);
and U6779 (N_6779,N_1377,N_4561);
or U6780 (N_6780,N_3342,N_4576);
nor U6781 (N_6781,N_2691,N_2969);
or U6782 (N_6782,N_4966,N_3048);
nand U6783 (N_6783,N_2552,N_4047);
and U6784 (N_6784,N_1562,N_61);
nor U6785 (N_6785,N_161,N_521);
or U6786 (N_6786,N_2796,N_4440);
or U6787 (N_6787,N_4141,N_990);
nor U6788 (N_6788,N_1598,N_929);
and U6789 (N_6789,N_4384,N_1076);
nor U6790 (N_6790,N_2344,N_4653);
nand U6791 (N_6791,N_2118,N_3560);
and U6792 (N_6792,N_4615,N_4852);
xnor U6793 (N_6793,N_4574,N_2777);
nand U6794 (N_6794,N_2480,N_3255);
xnor U6795 (N_6795,N_3165,N_1450);
nand U6796 (N_6796,N_4149,N_2053);
nor U6797 (N_6797,N_394,N_686);
or U6798 (N_6798,N_1700,N_3140);
or U6799 (N_6799,N_820,N_1200);
nand U6800 (N_6800,N_3440,N_4706);
xnor U6801 (N_6801,N_3668,N_3741);
nor U6802 (N_6802,N_3318,N_4212);
nor U6803 (N_6803,N_3135,N_2298);
or U6804 (N_6804,N_2112,N_2935);
or U6805 (N_6805,N_2639,N_2304);
or U6806 (N_6806,N_3878,N_1515);
nor U6807 (N_6807,N_764,N_1561);
xor U6808 (N_6808,N_580,N_352);
nand U6809 (N_6809,N_3346,N_3288);
nor U6810 (N_6810,N_3699,N_1830);
nand U6811 (N_6811,N_1,N_1723);
nand U6812 (N_6812,N_4400,N_3051);
or U6813 (N_6813,N_4250,N_1788);
or U6814 (N_6814,N_4436,N_1761);
and U6815 (N_6815,N_2582,N_790);
nand U6816 (N_6816,N_4262,N_3130);
nor U6817 (N_6817,N_2100,N_1063);
nor U6818 (N_6818,N_4088,N_1870);
nor U6819 (N_6819,N_2145,N_1727);
or U6820 (N_6820,N_2296,N_4673);
nand U6821 (N_6821,N_1464,N_3595);
and U6822 (N_6822,N_1323,N_233);
or U6823 (N_6823,N_4033,N_4113);
nand U6824 (N_6824,N_3265,N_1268);
nand U6825 (N_6825,N_4336,N_1262);
nor U6826 (N_6826,N_3562,N_4157);
and U6827 (N_6827,N_2994,N_1592);
nand U6828 (N_6828,N_238,N_3869);
and U6829 (N_6829,N_37,N_3509);
nand U6830 (N_6830,N_3091,N_2949);
nor U6831 (N_6831,N_2859,N_1856);
or U6832 (N_6832,N_3391,N_1291);
nand U6833 (N_6833,N_950,N_1885);
and U6834 (N_6834,N_1701,N_4686);
or U6835 (N_6835,N_1712,N_4127);
and U6836 (N_6836,N_1311,N_1980);
nor U6837 (N_6837,N_1936,N_4764);
and U6838 (N_6838,N_878,N_2931);
nor U6839 (N_6839,N_2431,N_794);
nand U6840 (N_6840,N_3534,N_1368);
or U6841 (N_6841,N_2538,N_4833);
and U6842 (N_6842,N_66,N_2229);
nor U6843 (N_6843,N_2596,N_1431);
nor U6844 (N_6844,N_1315,N_4276);
nand U6845 (N_6845,N_4358,N_3159);
nor U6846 (N_6846,N_659,N_2562);
xor U6847 (N_6847,N_706,N_918);
or U6848 (N_6848,N_725,N_4083);
and U6849 (N_6849,N_3829,N_2529);
nor U6850 (N_6850,N_3202,N_4650);
nor U6851 (N_6851,N_1495,N_4470);
nor U6852 (N_6852,N_4058,N_4959);
nand U6853 (N_6853,N_4655,N_2632);
xnor U6854 (N_6854,N_3752,N_4977);
nand U6855 (N_6855,N_2743,N_3053);
or U6856 (N_6856,N_3684,N_3723);
and U6857 (N_6857,N_2200,N_2327);
nor U6858 (N_6858,N_4996,N_4091);
and U6859 (N_6859,N_4130,N_4725);
nand U6860 (N_6860,N_3953,N_3806);
and U6861 (N_6861,N_1352,N_1964);
nand U6862 (N_6862,N_1463,N_3161);
and U6863 (N_6863,N_2780,N_440);
nor U6864 (N_6864,N_191,N_2649);
and U6865 (N_6865,N_2955,N_3661);
nor U6866 (N_6866,N_2465,N_284);
nand U6867 (N_6867,N_1869,N_249);
and U6868 (N_6868,N_3960,N_1657);
or U6869 (N_6869,N_4151,N_1949);
nor U6870 (N_6870,N_2877,N_4934);
or U6871 (N_6871,N_2340,N_2108);
nor U6872 (N_6872,N_4107,N_443);
and U6873 (N_6873,N_3397,N_961);
nor U6874 (N_6874,N_1279,N_3330);
nand U6875 (N_6875,N_452,N_4745);
or U6876 (N_6876,N_4351,N_1720);
or U6877 (N_6877,N_2146,N_4873);
nand U6878 (N_6878,N_3643,N_3323);
or U6879 (N_6879,N_3598,N_2039);
nand U6880 (N_6880,N_164,N_4933);
nor U6881 (N_6881,N_1893,N_4042);
and U6882 (N_6882,N_2844,N_2000);
and U6883 (N_6883,N_2129,N_4464);
nor U6884 (N_6884,N_1310,N_4306);
or U6885 (N_6885,N_1845,N_3040);
nor U6886 (N_6886,N_154,N_974);
nand U6887 (N_6887,N_302,N_3715);
nor U6888 (N_6888,N_1248,N_1473);
or U6889 (N_6889,N_4363,N_2134);
nand U6890 (N_6890,N_4109,N_176);
and U6891 (N_6891,N_2833,N_2002);
nor U6892 (N_6892,N_2776,N_1215);
nand U6893 (N_6893,N_2082,N_2182);
nor U6894 (N_6894,N_1146,N_4032);
or U6895 (N_6895,N_2717,N_2475);
nand U6896 (N_6896,N_899,N_2569);
and U6897 (N_6897,N_705,N_1369);
or U6898 (N_6898,N_1038,N_3944);
nor U6899 (N_6899,N_4037,N_2420);
nor U6900 (N_6900,N_1756,N_3608);
nand U6901 (N_6901,N_30,N_316);
or U6902 (N_6902,N_3272,N_2567);
and U6903 (N_6903,N_4490,N_2812);
nor U6904 (N_6904,N_1656,N_2991);
or U6905 (N_6905,N_2198,N_3276);
or U6906 (N_6906,N_653,N_53);
nor U6907 (N_6907,N_3701,N_2830);
nor U6908 (N_6908,N_1000,N_2533);
or U6909 (N_6909,N_855,N_1008);
and U6910 (N_6910,N_3984,N_2171);
or U6911 (N_6911,N_2191,N_4543);
nand U6912 (N_6912,N_7,N_2131);
nand U6913 (N_6913,N_319,N_146);
or U6914 (N_6914,N_1406,N_882);
nor U6915 (N_6915,N_80,N_773);
nor U6916 (N_6916,N_3033,N_2892);
and U6917 (N_6917,N_2564,N_3641);
and U6918 (N_6918,N_1002,N_3240);
or U6919 (N_6919,N_341,N_181);
nor U6920 (N_6920,N_195,N_2589);
and U6921 (N_6921,N_27,N_954);
or U6922 (N_6922,N_509,N_3401);
or U6923 (N_6923,N_503,N_618);
xnor U6924 (N_6924,N_4292,N_501);
or U6925 (N_6925,N_3520,N_2300);
nand U6926 (N_6926,N_3987,N_3106);
and U6927 (N_6927,N_3326,N_484);
and U6928 (N_6928,N_4255,N_4341);
or U6929 (N_6929,N_3914,N_1144);
nand U6930 (N_6930,N_2235,N_4424);
nor U6931 (N_6931,N_1894,N_3808);
or U6932 (N_6932,N_603,N_4169);
or U6933 (N_6933,N_730,N_2387);
and U6934 (N_6934,N_3321,N_4654);
xnor U6935 (N_6935,N_1103,N_1079);
and U6936 (N_6936,N_4218,N_4299);
or U6937 (N_6937,N_2101,N_1671);
xor U6938 (N_6938,N_3446,N_4456);
nor U6939 (N_6939,N_2918,N_2328);
nor U6940 (N_6940,N_3753,N_442);
nand U6941 (N_6941,N_936,N_2169);
and U6942 (N_6942,N_2910,N_620);
or U6943 (N_6943,N_3638,N_2318);
nand U6944 (N_6944,N_1214,N_172);
nand U6945 (N_6945,N_1498,N_946);
xnor U6946 (N_6946,N_3849,N_4343);
and U6947 (N_6947,N_4902,N_2179);
nand U6948 (N_6948,N_428,N_1749);
and U6949 (N_6949,N_4006,N_566);
nand U6950 (N_6950,N_118,N_4373);
nor U6951 (N_6951,N_4249,N_448);
or U6952 (N_6952,N_2063,N_1968);
and U6953 (N_6953,N_241,N_4028);
nor U6954 (N_6954,N_4414,N_212);
nand U6955 (N_6955,N_4927,N_1520);
xnor U6956 (N_6956,N_1367,N_703);
nand U6957 (N_6957,N_1163,N_4704);
nand U6958 (N_6958,N_1661,N_971);
nand U6959 (N_6959,N_1206,N_4985);
nand U6960 (N_6960,N_3731,N_337);
nand U6961 (N_6961,N_1699,N_3700);
or U6962 (N_6962,N_1877,N_3356);
and U6963 (N_6963,N_3627,N_93);
xor U6964 (N_6964,N_2686,N_4054);
nor U6965 (N_6965,N_751,N_538);
and U6966 (N_6966,N_4693,N_2797);
nand U6967 (N_6967,N_2659,N_3771);
xor U6968 (N_6968,N_4079,N_1533);
nand U6969 (N_6969,N_1259,N_1802);
nand U6970 (N_6970,N_3499,N_1882);
and U6971 (N_6971,N_15,N_3374);
and U6972 (N_6972,N_2226,N_1102);
xor U6973 (N_6973,N_626,N_3396);
nor U6974 (N_6974,N_1496,N_2332);
and U6975 (N_6975,N_3947,N_2366);
nor U6976 (N_6976,N_667,N_3496);
and U6977 (N_6977,N_3589,N_2029);
nand U6978 (N_6978,N_962,N_77);
nand U6979 (N_6979,N_376,N_4609);
and U6980 (N_6980,N_1277,N_2390);
nand U6981 (N_6981,N_4049,N_166);
or U6982 (N_6982,N_4007,N_3955);
nand U6983 (N_6983,N_1540,N_4921);
nor U6984 (N_6984,N_2008,N_3293);
nor U6985 (N_6985,N_4501,N_2706);
and U6986 (N_6986,N_4272,N_4513);
nor U6987 (N_6987,N_178,N_4641);
or U6988 (N_6988,N_1930,N_3993);
nand U6989 (N_6989,N_2488,N_3132);
or U6990 (N_6990,N_926,N_3640);
or U6991 (N_6991,N_4822,N_2555);
nand U6992 (N_6992,N_1652,N_1354);
xor U6993 (N_6993,N_3289,N_4059);
nor U6994 (N_6994,N_2973,N_3653);
and U6995 (N_6995,N_2616,N_4312);
or U6996 (N_6996,N_2843,N_740);
and U6997 (N_6997,N_4445,N_739);
or U6998 (N_6998,N_2421,N_4375);
or U6999 (N_6999,N_2742,N_2067);
nand U7000 (N_7000,N_4767,N_1021);
nor U7001 (N_7001,N_564,N_1308);
and U7002 (N_7002,N_2766,N_2779);
and U7003 (N_7003,N_3921,N_3876);
or U7004 (N_7004,N_3223,N_1925);
nand U7005 (N_7005,N_4807,N_1086);
nor U7006 (N_7006,N_2952,N_101);
nor U7007 (N_7007,N_4087,N_972);
nor U7008 (N_7008,N_3119,N_1941);
or U7009 (N_7009,N_4838,N_2925);
nor U7010 (N_7010,N_464,N_3450);
or U7011 (N_7011,N_4591,N_1572);
xnor U7012 (N_7012,N_3149,N_2537);
or U7013 (N_7013,N_4112,N_1294);
or U7014 (N_7014,N_1526,N_1542);
nor U7015 (N_7015,N_4023,N_2643);
or U7016 (N_7016,N_4311,N_1173);
and U7017 (N_7017,N_3985,N_207);
or U7018 (N_7018,N_3218,N_4265);
or U7019 (N_7019,N_3538,N_1543);
and U7020 (N_7020,N_3708,N_4096);
nand U7021 (N_7021,N_994,N_4816);
nor U7022 (N_7022,N_3516,N_3660);
and U7023 (N_7023,N_2068,N_2852);
xor U7024 (N_7024,N_3707,N_3384);
and U7025 (N_7025,N_3894,N_299);
nand U7026 (N_7026,N_843,N_3320);
and U7027 (N_7027,N_2784,N_3445);
nor U7028 (N_7028,N_60,N_4217);
nand U7029 (N_7029,N_2866,N_1524);
or U7030 (N_7030,N_2361,N_2329);
or U7031 (N_7031,N_996,N_4000);
or U7032 (N_7032,N_2066,N_2441);
and U7033 (N_7033,N_2137,N_4463);
and U7034 (N_7034,N_4357,N_3596);
nand U7035 (N_7035,N_1985,N_1546);
or U7036 (N_7036,N_2035,N_731);
nor U7037 (N_7037,N_1134,N_777);
nand U7038 (N_7038,N_4426,N_2604);
or U7039 (N_7039,N_1538,N_1328);
nand U7040 (N_7040,N_2752,N_1505);
and U7041 (N_7041,N_232,N_2598);
nand U7042 (N_7042,N_1556,N_4171);
and U7043 (N_7043,N_1381,N_2015);
xnor U7044 (N_7044,N_4447,N_3084);
nor U7045 (N_7045,N_1819,N_1029);
and U7046 (N_7046,N_2201,N_1339);
nand U7047 (N_7047,N_2636,N_502);
and U7048 (N_7048,N_3959,N_2380);
or U7049 (N_7049,N_2561,N_4786);
nand U7050 (N_7050,N_2313,N_187);
nand U7051 (N_7051,N_2204,N_673);
or U7052 (N_7052,N_1333,N_281);
nor U7053 (N_7053,N_2873,N_1800);
nand U7054 (N_7054,N_2945,N_151);
and U7055 (N_7055,N_4483,N_2350);
nand U7056 (N_7056,N_4774,N_2504);
nand U7057 (N_7057,N_4176,N_3886);
nor U7058 (N_7058,N_792,N_4479);
nand U7059 (N_7059,N_1395,N_803);
or U7060 (N_7060,N_2702,N_1231);
or U7061 (N_7061,N_4396,N_3644);
or U7062 (N_7062,N_2195,N_4505);
nor U7063 (N_7063,N_379,N_1165);
and U7064 (N_7064,N_2001,N_1651);
nand U7065 (N_7065,N_304,N_2231);
nor U7066 (N_7066,N_1479,N_4989);
and U7067 (N_7067,N_661,N_1440);
or U7068 (N_7068,N_2062,N_3307);
and U7069 (N_7069,N_4146,N_4457);
nand U7070 (N_7070,N_997,N_106);
nor U7071 (N_7071,N_2735,N_4629);
nor U7072 (N_7072,N_2715,N_1916);
nor U7073 (N_7073,N_1860,N_2939);
nor U7074 (N_7074,N_741,N_582);
and U7075 (N_7075,N_4537,N_2868);
nor U7076 (N_7076,N_2384,N_2864);
nor U7077 (N_7077,N_2143,N_4530);
nand U7078 (N_7078,N_947,N_4751);
nor U7079 (N_7079,N_286,N_248);
nor U7080 (N_7080,N_1908,N_956);
xnor U7081 (N_7081,N_3406,N_3623);
and U7082 (N_7082,N_268,N_1126);
nor U7083 (N_7083,N_4334,N_1738);
nor U7084 (N_7084,N_4544,N_1030);
nor U7085 (N_7085,N_2138,N_4314);
nand U7086 (N_7086,N_3897,N_3007);
and U7087 (N_7087,N_2370,N_4705);
or U7088 (N_7088,N_4359,N_2982);
or U7089 (N_7089,N_1646,N_1794);
nor U7090 (N_7090,N_4504,N_4062);
nor U7091 (N_7091,N_3949,N_4503);
and U7092 (N_7092,N_3382,N_2404);
and U7093 (N_7093,N_1202,N_3765);
nand U7094 (N_7094,N_3266,N_2849);
nor U7095 (N_7095,N_4132,N_1835);
nor U7096 (N_7096,N_744,N_4216);
nor U7097 (N_7097,N_2662,N_2410);
xnor U7098 (N_7098,N_2293,N_1928);
and U7099 (N_7099,N_1199,N_985);
or U7100 (N_7100,N_2763,N_1853);
nor U7101 (N_7101,N_3574,N_2317);
nor U7102 (N_7102,N_1035,N_4851);
or U7103 (N_7103,N_2685,N_1187);
nand U7104 (N_7104,N_1088,N_4891);
nor U7105 (N_7105,N_2087,N_3046);
nand U7106 (N_7106,N_561,N_1371);
and U7107 (N_7107,N_3932,N_4785);
nand U7108 (N_7108,N_2266,N_3785);
nor U7109 (N_7109,N_3972,N_2867);
nor U7110 (N_7110,N_1241,N_2073);
xnor U7111 (N_7111,N_288,N_2004);
and U7112 (N_7112,N_3629,N_3717);
nand U7113 (N_7113,N_1817,N_1582);
nor U7114 (N_7114,N_2921,N_593);
or U7115 (N_7115,N_3584,N_2047);
xnor U7116 (N_7116,N_713,N_2209);
nor U7117 (N_7117,N_4134,N_2524);
nand U7118 (N_7118,N_4246,N_643);
nand U7119 (N_7119,N_1436,N_3405);
nor U7120 (N_7120,N_3136,N_1672);
nor U7121 (N_7121,N_2306,N_4260);
and U7122 (N_7122,N_1182,N_650);
and U7123 (N_7123,N_4082,N_2943);
or U7124 (N_7124,N_4957,N_2297);
nand U7125 (N_7125,N_3879,N_2254);
or U7126 (N_7126,N_4750,N_18);
xnor U7127 (N_7127,N_2848,N_3037);
xor U7128 (N_7128,N_2183,N_1997);
and U7129 (N_7129,N_285,N_1322);
or U7130 (N_7130,N_4485,N_3981);
nand U7131 (N_7131,N_2349,N_959);
and U7132 (N_7132,N_203,N_130);
nand U7133 (N_7133,N_1662,N_3195);
or U7134 (N_7134,N_927,N_2721);
nor U7135 (N_7135,N_2271,N_3529);
nand U7136 (N_7136,N_592,N_50);
and U7137 (N_7137,N_2075,N_4050);
nand U7138 (N_7138,N_1887,N_4480);
nor U7139 (N_7139,N_3,N_3333);
nor U7140 (N_7140,N_3526,N_1236);
nand U7141 (N_7141,N_4150,N_1816);
or U7142 (N_7142,N_4715,N_4179);
or U7143 (N_7143,N_3837,N_3588);
and U7144 (N_7144,N_2405,N_3571);
nor U7145 (N_7145,N_2376,N_1629);
nand U7146 (N_7146,N_687,N_3709);
and U7147 (N_7147,N_3078,N_1267);
and U7148 (N_7148,N_3432,N_4948);
or U7149 (N_7149,N_1824,N_1593);
or U7150 (N_7150,N_3542,N_2578);
and U7151 (N_7151,N_4583,N_1306);
and U7152 (N_7152,N_1128,N_1400);
or U7153 (N_7153,N_1171,N_4662);
nor U7154 (N_7154,N_3871,N_599);
or U7155 (N_7155,N_1137,N_4687);
and U7156 (N_7156,N_2645,N_4174);
nor U7157 (N_7157,N_2351,N_259);
nand U7158 (N_7158,N_334,N_4582);
nor U7159 (N_7159,N_2525,N_1745);
nand U7160 (N_7160,N_1363,N_2889);
or U7161 (N_7161,N_1033,N_4930);
nand U7162 (N_7162,N_922,N_3679);
nand U7163 (N_7163,N_549,N_2287);
nand U7164 (N_7164,N_2996,N_2518);
nand U7165 (N_7165,N_2663,N_3995);
nor U7166 (N_7166,N_3904,N_4200);
nor U7167 (N_7167,N_1399,N_2947);
nor U7168 (N_7168,N_3250,N_2508);
or U7169 (N_7169,N_89,N_3127);
or U7170 (N_7170,N_134,N_4055);
nand U7171 (N_7171,N_4316,N_995);
and U7172 (N_7172,N_3347,N_2909);
or U7173 (N_7173,N_1100,N_3182);
or U7174 (N_7174,N_1032,N_3658);
or U7175 (N_7175,N_3515,N_746);
nand U7176 (N_7176,N_3116,N_3238);
or U7177 (N_7177,N_4450,N_2792);
nor U7178 (N_7178,N_887,N_546);
xnor U7179 (N_7179,N_1375,N_2613);
nor U7180 (N_7180,N_2019,N_1222);
nand U7181 (N_7181,N_2521,N_2699);
or U7182 (N_7182,N_2319,N_4126);
or U7183 (N_7183,N_3784,N_1417);
xnor U7184 (N_7184,N_3605,N_919);
and U7185 (N_7185,N_2104,N_1314);
and U7186 (N_7186,N_1620,N_3380);
and U7187 (N_7187,N_2922,N_4332);
nand U7188 (N_7188,N_891,N_2069);
nand U7189 (N_7189,N_167,N_845);
and U7190 (N_7190,N_1261,N_4335);
or U7191 (N_7191,N_4857,N_924);
nand U7192 (N_7192,N_1360,N_3387);
and U7193 (N_7193,N_322,N_3267);
nor U7194 (N_7194,N_1421,N_1472);
nand U7195 (N_7195,N_6,N_3193);
nand U7196 (N_7196,N_397,N_2531);
nor U7197 (N_7197,N_4765,N_2692);
or U7198 (N_7198,N_3373,N_1510);
and U7199 (N_7199,N_3632,N_574);
and U7200 (N_7200,N_2162,N_2290);
and U7201 (N_7201,N_2836,N_2025);
or U7202 (N_7202,N_3424,N_3023);
nand U7203 (N_7203,N_2689,N_2485);
and U7204 (N_7204,N_732,N_2150);
nand U7205 (N_7205,N_3905,N_192);
nor U7206 (N_7206,N_4317,N_4991);
nand U7207 (N_7207,N_2676,N_1075);
and U7208 (N_7208,N_2013,N_365);
or U7209 (N_7209,N_1619,N_2149);
nor U7210 (N_7210,N_3219,N_3738);
nor U7211 (N_7211,N_3647,N_4995);
nor U7212 (N_7212,N_3982,N_2560);
nand U7213 (N_7213,N_1539,N_3253);
nor U7214 (N_7214,N_3399,N_2690);
nor U7215 (N_7215,N_4746,N_4519);
nand U7216 (N_7216,N_75,N_1391);
nor U7217 (N_7217,N_4747,N_4252);
and U7218 (N_7218,N_4484,N_3352);
nor U7219 (N_7219,N_3378,N_4935);
nor U7220 (N_7220,N_4197,N_3376);
xor U7221 (N_7221,N_749,N_1717);
nand U7222 (N_7222,N_4043,N_2294);
nor U7223 (N_7223,N_789,N_3481);
nor U7224 (N_7224,N_4187,N_4908);
nand U7225 (N_7225,N_1410,N_953);
and U7226 (N_7226,N_2094,N_3954);
nand U7227 (N_7227,N_1408,N_1650);
nand U7228 (N_7228,N_483,N_2988);
xnor U7229 (N_7229,N_2103,N_1683);
and U7230 (N_7230,N_4095,N_1677);
and U7231 (N_7231,N_2048,N_2750);
or U7232 (N_7232,N_935,N_981);
nor U7233 (N_7233,N_3548,N_689);
or U7234 (N_7234,N_4089,N_1142);
nand U7235 (N_7235,N_4839,N_4889);
xor U7236 (N_7236,N_1415,N_2575);
nor U7237 (N_7237,N_2299,N_3863);
nor U7238 (N_7238,N_3056,N_2694);
nor U7239 (N_7239,N_3733,N_805);
xor U7240 (N_7240,N_405,N_4595);
nor U7241 (N_7241,N_2238,N_2045);
or U7242 (N_7242,N_3903,N_1394);
or U7243 (N_7243,N_458,N_3853);
or U7244 (N_7244,N_1194,N_131);
nand U7245 (N_7245,N_567,N_1471);
nand U7246 (N_7246,N_1973,N_2938);
nand U7247 (N_7247,N_292,N_837);
or U7248 (N_7248,N_1634,N_504);
and U7249 (N_7249,N_3552,N_3441);
and U7250 (N_7250,N_2698,N_2222);
and U7251 (N_7251,N_709,N_638);
or U7252 (N_7252,N_2099,N_2237);
and U7253 (N_7253,N_2353,N_40);
nor U7254 (N_7254,N_3986,N_1443);
nand U7255 (N_7255,N_1221,N_578);
nor U7256 (N_7256,N_454,N_2136);
nor U7257 (N_7257,N_2447,N_2841);
or U7258 (N_7258,N_4201,N_4804);
nand U7259 (N_7259,N_1514,N_1305);
nand U7260 (N_7260,N_330,N_1842);
nand U7261 (N_7261,N_3354,N_3730);
and U7262 (N_7262,N_4118,N_2278);
and U7263 (N_7263,N_4619,N_3702);
and U7264 (N_7264,N_3593,N_660);
nor U7265 (N_7265,N_2553,N_3337);
or U7266 (N_7266,N_331,N_4084);
nand U7267 (N_7267,N_4982,N_2563);
nor U7268 (N_7268,N_3029,N_3811);
nor U7269 (N_7269,N_4598,N_761);
and U7270 (N_7270,N_1006,N_1624);
and U7271 (N_7271,N_3761,N_2325);
or U7272 (N_7272,N_426,N_4708);
or U7273 (N_7273,N_456,N_4788);
nand U7274 (N_7274,N_1162,N_2443);
nor U7275 (N_7275,N_1018,N_1641);
and U7276 (N_7276,N_4155,N_385);
nand U7277 (N_7277,N_3652,N_4021);
and U7278 (N_7278,N_1521,N_831);
and U7279 (N_7279,N_2492,N_4135);
or U7280 (N_7280,N_1300,N_493);
nor U7281 (N_7281,N_551,N_1927);
and U7282 (N_7282,N_2374,N_4757);
nor U7283 (N_7283,N_3199,N_4510);
or U7284 (N_7284,N_3156,N_2230);
and U7285 (N_7285,N_4865,N_3494);
and U7286 (N_7286,N_2268,N_2072);
nor U7287 (N_7287,N_3004,N_711);
and U7288 (N_7288,N_1470,N_4795);
nor U7289 (N_7289,N_280,N_1554);
and U7290 (N_7290,N_973,N_2407);
nand U7291 (N_7291,N_1772,N_1682);
and U7292 (N_7292,N_3340,N_4769);
xor U7293 (N_7293,N_4015,N_3345);
nand U7294 (N_7294,N_3695,N_3776);
and U7295 (N_7295,N_4811,N_1224);
and U7296 (N_7296,N_3533,N_2360);
or U7297 (N_7297,N_2651,N_3675);
nand U7298 (N_7298,N_3418,N_3425);
or U7299 (N_7299,N_51,N_2593);
nor U7300 (N_7300,N_252,N_3844);
nor U7301 (N_7301,N_1418,N_3587);
or U7302 (N_7302,N_1036,N_2355);
nand U7303 (N_7303,N_4649,N_4652);
or U7304 (N_7304,N_1181,N_2081);
nand U7305 (N_7305,N_1642,N_1484);
nor U7306 (N_7306,N_64,N_3648);
nor U7307 (N_7307,N_4326,N_3457);
nand U7308 (N_7308,N_4644,N_410);
and U7309 (N_7309,N_3244,N_1812);
nor U7310 (N_7310,N_3442,N_2378);
or U7311 (N_7311,N_2244,N_3528);
nor U7312 (N_7312,N_3872,N_487);
nand U7313 (N_7313,N_2106,N_219);
nor U7314 (N_7314,N_2726,N_3379);
nand U7315 (N_7315,N_3353,N_1596);
nand U7316 (N_7316,N_3157,N_2911);
and U7317 (N_7317,N_2109,N_683);
xnor U7318 (N_7318,N_4886,N_1529);
nand U7319 (N_7319,N_1631,N_1420);
nor U7320 (N_7320,N_2653,N_1132);
and U7321 (N_7321,N_1898,N_4177);
nand U7322 (N_7322,N_3421,N_627);
and U7323 (N_7323,N_4173,N_1932);
nand U7324 (N_7324,N_480,N_3190);
or U7325 (N_7325,N_884,N_1563);
xnor U7326 (N_7326,N_1663,N_2681);
and U7327 (N_7327,N_4729,N_991);
nor U7328 (N_7328,N_1003,N_760);
and U7329 (N_7329,N_2782,N_4364);
nand U7330 (N_7330,N_3937,N_910);
nor U7331 (N_7331,N_535,N_217);
and U7332 (N_7332,N_2044,N_1016);
nor U7333 (N_7333,N_4439,N_4509);
nand U7334 (N_7334,N_33,N_3429);
nand U7335 (N_7335,N_4562,N_4892);
nor U7336 (N_7336,N_3845,N_2795);
nor U7337 (N_7337,N_2126,N_2503);
nor U7338 (N_7338,N_4997,N_682);
xnor U7339 (N_7339,N_4698,N_1183);
and U7340 (N_7340,N_1281,N_3790);
or U7341 (N_7341,N_2888,N_4971);
and U7342 (N_7342,N_372,N_135);
or U7343 (N_7343,N_2946,N_863);
nand U7344 (N_7344,N_3437,N_1668);
nor U7345 (N_7345,N_2585,N_3568);
nor U7346 (N_7346,N_1023,N_3338);
or U7347 (N_7347,N_2856,N_2850);
nand U7348 (N_7348,N_2490,N_4888);
and U7349 (N_7349,N_202,N_4409);
and U7350 (N_7350,N_263,N_4899);
or U7351 (N_7351,N_3956,N_2009);
nand U7352 (N_7352,N_1577,N_986);
and U7353 (N_7353,N_3392,N_4613);
nand U7354 (N_7354,N_2456,N_4779);
nand U7355 (N_7355,N_303,N_2837);
nand U7356 (N_7356,N_1987,N_1085);
and U7357 (N_7357,N_4894,N_10);
nand U7358 (N_7358,N_4261,N_2760);
xor U7359 (N_7359,N_2583,N_105);
or U7360 (N_7360,N_1724,N_2903);
and U7361 (N_7361,N_3117,N_4417);
nor U7362 (N_7362,N_3603,N_2904);
and U7363 (N_7363,N_2775,N_3583);
and U7364 (N_7364,N_2933,N_1190);
and U7365 (N_7365,N_1327,N_3270);
or U7366 (N_7366,N_2566,N_4362);
nor U7367 (N_7367,N_4713,N_211);
nor U7368 (N_7368,N_4108,N_1435);
or U7369 (N_7369,N_208,N_1970);
nand U7370 (N_7370,N_2550,N_3617);
or U7371 (N_7371,N_362,N_2479);
and U7372 (N_7372,N_2999,N_4154);
nand U7373 (N_7373,N_221,N_4381);
nor U7374 (N_7374,N_4616,N_2213);
nor U7375 (N_7375,N_3435,N_980);
nand U7376 (N_7376,N_2124,N_1219);
or U7377 (N_7377,N_1680,N_2871);
and U7378 (N_7378,N_3269,N_4305);
nand U7379 (N_7379,N_4101,N_556);
nand U7380 (N_7380,N_4168,N_3941);
nor U7381 (N_7381,N_3062,N_1462);
nand U7382 (N_7382,N_3746,N_3816);
and U7383 (N_7383,N_1331,N_4009);
nand U7384 (N_7384,N_360,N_478);
nand U7385 (N_7385,N_4722,N_4579);
xor U7386 (N_7386,N_499,N_3107);
and U7387 (N_7387,N_460,N_1256);
nand U7388 (N_7388,N_4008,N_469);
and U7389 (N_7389,N_400,N_2363);
or U7390 (N_7390,N_3606,N_4383);
and U7391 (N_7391,N_4371,N_2341);
and U7392 (N_7392,N_4550,N_3126);
nor U7393 (N_7393,N_3016,N_2749);
and U7394 (N_7394,N_3851,N_2897);
or U7395 (N_7395,N_3635,N_1107);
xor U7396 (N_7396,N_4776,N_3414);
and U7397 (N_7397,N_598,N_1409);
nand U7398 (N_7398,N_4423,N_1407);
nor U7399 (N_7399,N_2682,N_3039);
nand U7400 (N_7400,N_2588,N_539);
or U7401 (N_7401,N_700,N_1240);
nor U7402 (N_7402,N_862,N_4812);
nand U7403 (N_7403,N_3797,N_4878);
or U7404 (N_7404,N_4518,N_1687);
and U7405 (N_7405,N_2787,N_4502);
and U7406 (N_7406,N_575,N_1905);
and U7407 (N_7407,N_3681,N_1220);
and U7408 (N_7408,N_3092,N_3434);
and U7409 (N_7409,N_1362,N_4065);
nor U7410 (N_7410,N_4536,N_4206);
or U7411 (N_7411,N_4231,N_1325);
and U7412 (N_7412,N_531,N_4449);
or U7413 (N_7413,N_4599,N_1423);
or U7414 (N_7414,N_3109,N_3669);
nand U7415 (N_7415,N_2975,N_1750);
xor U7416 (N_7416,N_4339,N_1460);
and U7417 (N_7417,N_432,N_4437);
and U7418 (N_7418,N_3757,N_2105);
nor U7419 (N_7419,N_4214,N_3665);
and U7420 (N_7420,N_541,N_3128);
nor U7421 (N_7421,N_4689,N_1386);
or U7422 (N_7422,N_628,N_1009);
nand U7423 (N_7423,N_4871,N_2919);
nor U7424 (N_7424,N_1110,N_81);
nand U7425 (N_7425,N_727,N_3246);
and U7426 (N_7426,N_3484,N_1686);
or U7427 (N_7427,N_4319,N_1047);
or U7428 (N_7428,N_4531,N_12);
nor U7429 (N_7429,N_1358,N_4926);
nor U7430 (N_7430,N_1991,N_3673);
nor U7431 (N_7431,N_2778,N_3013);
nand U7432 (N_7432,N_3962,N_137);
and U7433 (N_7433,N_190,N_2464);
nand U7434 (N_7434,N_3000,N_3682);
nand U7435 (N_7435,N_3327,N_210);
nor U7436 (N_7436,N_4545,N_4571);
and U7437 (N_7437,N_4382,N_702);
and U7438 (N_7438,N_3967,N_4773);
nor U7439 (N_7439,N_854,N_4577);
nand U7440 (N_7440,N_1832,N_4665);
nor U7441 (N_7441,N_1740,N_3410);
or U7442 (N_7442,N_3497,N_3651);
nor U7443 (N_7443,N_55,N_2879);
nand U7444 (N_7444,N_1922,N_2610);
or U7445 (N_7445,N_2096,N_2086);
nand U7446 (N_7446,N_2119,N_4755);
and U7447 (N_7447,N_4073,N_4254);
nor U7448 (N_7448,N_1979,N_415);
or U7449 (N_7449,N_528,N_265);
nor U7450 (N_7450,N_3221,N_1919);
nand U7451 (N_7451,N_1232,N_2606);
and U7452 (N_7452,N_2672,N_3820);
and U7453 (N_7453,N_606,N_4600);
or U7454 (N_7454,N_4758,N_4845);
nand U7455 (N_7455,N_2711,N_4193);
and U7456 (N_7456,N_3371,N_4379);
nor U7457 (N_7457,N_1966,N_2958);
nand U7458 (N_7458,N_471,N_35);
and U7459 (N_7459,N_4932,N_2003);
nand U7460 (N_7460,N_100,N_4374);
nor U7461 (N_7461,N_2391,N_20);
or U7462 (N_7462,N_306,N_4203);
nor U7463 (N_7463,N_4581,N_1475);
or U7464 (N_7464,N_625,N_3073);
or U7465 (N_7465,N_3639,N_3839);
or U7466 (N_7466,N_2884,N_3756);
nor U7467 (N_7467,N_2417,N_4068);
nor U7468 (N_7468,N_4493,N_3252);
and U7469 (N_7469,N_558,N_1605);
nand U7470 (N_7470,N_2744,N_3968);
nor U7471 (N_7471,N_4365,N_4477);
or U7472 (N_7472,N_3017,N_1878);
or U7473 (N_7473,N_445,N_2247);
nor U7474 (N_7474,N_572,N_2607);
nand U7475 (N_7475,N_2102,N_2708);
nand U7476 (N_7476,N_1813,N_3064);
or U7477 (N_7477,N_4404,N_4018);
nand U7478 (N_7478,N_4645,N_4258);
and U7479 (N_7479,N_505,N_4826);
nor U7480 (N_7480,N_3370,N_2847);
nor U7481 (N_7481,N_2901,N_550);
or U7482 (N_7482,N_1924,N_2870);
nand U7483 (N_7483,N_1993,N_1601);
xor U7484 (N_7484,N_571,N_1379);
nor U7485 (N_7485,N_3710,N_3468);
nand U7486 (N_7486,N_810,N_4012);
nor U7487 (N_7487,N_1244,N_4986);
or U7488 (N_7488,N_2249,N_788);
nor U7489 (N_7489,N_2530,N_237);
or U7490 (N_7490,N_1434,N_2090);
nor U7491 (N_7491,N_754,N_4517);
and U7492 (N_7492,N_3561,N_1080);
nor U7493 (N_7493,N_4585,N_4815);
nor U7494 (N_7494,N_553,N_923);
nand U7495 (N_7495,N_2617,N_4192);
nand U7496 (N_7496,N_2292,N_1133);
nor U7497 (N_7497,N_2912,N_2619);
nor U7498 (N_7498,N_2469,N_255);
or U7499 (N_7499,N_637,N_2064);
nor U7500 (N_7500,N_3476,N_243);
nand U7501 (N_7501,N_1415,N_2717);
or U7502 (N_7502,N_143,N_2549);
nand U7503 (N_7503,N_1494,N_58);
and U7504 (N_7504,N_850,N_228);
nand U7505 (N_7505,N_2089,N_1508);
or U7506 (N_7506,N_3904,N_1991);
or U7507 (N_7507,N_4579,N_979);
or U7508 (N_7508,N_1422,N_1283);
nand U7509 (N_7509,N_1595,N_4925);
and U7510 (N_7510,N_1129,N_3083);
or U7511 (N_7511,N_801,N_2430);
and U7512 (N_7512,N_4552,N_1596);
nand U7513 (N_7513,N_4609,N_3361);
or U7514 (N_7514,N_2250,N_4660);
and U7515 (N_7515,N_2557,N_2337);
nor U7516 (N_7516,N_3300,N_3368);
or U7517 (N_7517,N_668,N_4931);
or U7518 (N_7518,N_2048,N_210);
or U7519 (N_7519,N_1348,N_1947);
and U7520 (N_7520,N_1467,N_2245);
nor U7521 (N_7521,N_900,N_4879);
nor U7522 (N_7522,N_4413,N_3138);
nor U7523 (N_7523,N_756,N_228);
nor U7524 (N_7524,N_4239,N_3197);
or U7525 (N_7525,N_4749,N_2057);
and U7526 (N_7526,N_993,N_4990);
and U7527 (N_7527,N_3312,N_2155);
nor U7528 (N_7528,N_4900,N_1032);
or U7529 (N_7529,N_478,N_1383);
nor U7530 (N_7530,N_3183,N_4751);
and U7531 (N_7531,N_855,N_2970);
nor U7532 (N_7532,N_2284,N_4452);
nand U7533 (N_7533,N_3618,N_4184);
xnor U7534 (N_7534,N_1215,N_3485);
nand U7535 (N_7535,N_3484,N_25);
nor U7536 (N_7536,N_3845,N_3918);
or U7537 (N_7537,N_2055,N_3454);
nor U7538 (N_7538,N_3910,N_955);
and U7539 (N_7539,N_3707,N_4541);
nand U7540 (N_7540,N_2670,N_3641);
nand U7541 (N_7541,N_4565,N_100);
nand U7542 (N_7542,N_4759,N_2515);
or U7543 (N_7543,N_2242,N_255);
nor U7544 (N_7544,N_872,N_192);
nor U7545 (N_7545,N_902,N_4212);
xnor U7546 (N_7546,N_1372,N_2712);
nand U7547 (N_7547,N_1350,N_3056);
nand U7548 (N_7548,N_2295,N_196);
nor U7549 (N_7549,N_1354,N_3043);
or U7550 (N_7550,N_1011,N_4572);
nand U7551 (N_7551,N_1439,N_2493);
nand U7552 (N_7552,N_2918,N_3752);
nor U7553 (N_7553,N_4204,N_3419);
or U7554 (N_7554,N_4073,N_3114);
and U7555 (N_7555,N_3052,N_1151);
and U7556 (N_7556,N_3449,N_3995);
nand U7557 (N_7557,N_3407,N_2110);
nand U7558 (N_7558,N_3206,N_4643);
and U7559 (N_7559,N_3461,N_3475);
nand U7560 (N_7560,N_2987,N_4380);
or U7561 (N_7561,N_2165,N_825);
nor U7562 (N_7562,N_566,N_765);
nor U7563 (N_7563,N_1592,N_2594);
nand U7564 (N_7564,N_3989,N_1101);
and U7565 (N_7565,N_3390,N_3303);
nor U7566 (N_7566,N_2271,N_148);
nand U7567 (N_7567,N_91,N_3162);
or U7568 (N_7568,N_794,N_3379);
or U7569 (N_7569,N_1358,N_2199);
nand U7570 (N_7570,N_4802,N_2492);
nand U7571 (N_7571,N_3461,N_4754);
nand U7572 (N_7572,N_3447,N_4429);
nand U7573 (N_7573,N_1541,N_452);
nor U7574 (N_7574,N_3170,N_2152);
and U7575 (N_7575,N_4017,N_4567);
or U7576 (N_7576,N_1900,N_333);
nand U7577 (N_7577,N_2443,N_470);
nor U7578 (N_7578,N_4201,N_4700);
and U7579 (N_7579,N_1079,N_4608);
nor U7580 (N_7580,N_393,N_799);
or U7581 (N_7581,N_1736,N_1026);
or U7582 (N_7582,N_1434,N_1429);
nor U7583 (N_7583,N_3048,N_1651);
or U7584 (N_7584,N_3934,N_1221);
or U7585 (N_7585,N_4505,N_1347);
nand U7586 (N_7586,N_4481,N_1917);
nand U7587 (N_7587,N_3522,N_2581);
or U7588 (N_7588,N_4329,N_4269);
xor U7589 (N_7589,N_481,N_316);
nor U7590 (N_7590,N_1545,N_2965);
and U7591 (N_7591,N_3648,N_3447);
nand U7592 (N_7592,N_2760,N_1808);
and U7593 (N_7593,N_4243,N_854);
or U7594 (N_7594,N_2586,N_3515);
xnor U7595 (N_7595,N_2538,N_3296);
or U7596 (N_7596,N_1059,N_379);
nand U7597 (N_7597,N_3834,N_4151);
and U7598 (N_7598,N_3153,N_1830);
nor U7599 (N_7599,N_1571,N_3458);
nor U7600 (N_7600,N_2986,N_2796);
nor U7601 (N_7601,N_514,N_1836);
nor U7602 (N_7602,N_2386,N_1311);
nand U7603 (N_7603,N_4014,N_3808);
nor U7604 (N_7604,N_2457,N_3885);
nand U7605 (N_7605,N_3829,N_4959);
or U7606 (N_7606,N_3252,N_1081);
nand U7607 (N_7607,N_4148,N_2573);
nor U7608 (N_7608,N_1547,N_440);
and U7609 (N_7609,N_4509,N_2296);
nor U7610 (N_7610,N_1694,N_2610);
or U7611 (N_7611,N_3737,N_2737);
nand U7612 (N_7612,N_2768,N_4073);
nand U7613 (N_7613,N_4890,N_1774);
or U7614 (N_7614,N_3615,N_2060);
nor U7615 (N_7615,N_2407,N_4327);
and U7616 (N_7616,N_4184,N_2283);
and U7617 (N_7617,N_2683,N_3034);
and U7618 (N_7618,N_3903,N_4661);
nor U7619 (N_7619,N_1904,N_3628);
and U7620 (N_7620,N_1318,N_4585);
and U7621 (N_7621,N_2933,N_80);
nand U7622 (N_7622,N_2701,N_2388);
or U7623 (N_7623,N_2307,N_4599);
nand U7624 (N_7624,N_61,N_3278);
nand U7625 (N_7625,N_3065,N_3954);
nand U7626 (N_7626,N_4152,N_2752);
and U7627 (N_7627,N_1487,N_4773);
nor U7628 (N_7628,N_460,N_4709);
nor U7629 (N_7629,N_3686,N_4159);
or U7630 (N_7630,N_964,N_1138);
or U7631 (N_7631,N_4503,N_4842);
nand U7632 (N_7632,N_3641,N_1177);
nand U7633 (N_7633,N_3102,N_4353);
and U7634 (N_7634,N_1472,N_1384);
nand U7635 (N_7635,N_1599,N_3117);
nor U7636 (N_7636,N_3726,N_1024);
or U7637 (N_7637,N_338,N_282);
nand U7638 (N_7638,N_4884,N_1024);
and U7639 (N_7639,N_748,N_2285);
nand U7640 (N_7640,N_3057,N_1607);
and U7641 (N_7641,N_3526,N_4443);
or U7642 (N_7642,N_2464,N_3775);
or U7643 (N_7643,N_622,N_230);
nor U7644 (N_7644,N_3048,N_3670);
nand U7645 (N_7645,N_2115,N_3481);
or U7646 (N_7646,N_2222,N_144);
and U7647 (N_7647,N_3401,N_1666);
and U7648 (N_7648,N_3803,N_253);
nand U7649 (N_7649,N_1732,N_3558);
or U7650 (N_7650,N_1837,N_3354);
and U7651 (N_7651,N_670,N_3506);
nand U7652 (N_7652,N_2081,N_1767);
nand U7653 (N_7653,N_171,N_4188);
and U7654 (N_7654,N_4567,N_2836);
nor U7655 (N_7655,N_2979,N_2765);
or U7656 (N_7656,N_389,N_3739);
nand U7657 (N_7657,N_4982,N_2585);
nor U7658 (N_7658,N_621,N_1582);
nand U7659 (N_7659,N_3878,N_4842);
and U7660 (N_7660,N_2145,N_1175);
nand U7661 (N_7661,N_3207,N_2954);
or U7662 (N_7662,N_3520,N_2724);
nor U7663 (N_7663,N_500,N_1584);
and U7664 (N_7664,N_1630,N_1285);
or U7665 (N_7665,N_570,N_3899);
nand U7666 (N_7666,N_3665,N_2436);
nor U7667 (N_7667,N_1102,N_3638);
or U7668 (N_7668,N_4106,N_3544);
nand U7669 (N_7669,N_620,N_4315);
or U7670 (N_7670,N_2570,N_3847);
or U7671 (N_7671,N_922,N_3296);
nor U7672 (N_7672,N_4581,N_3551);
or U7673 (N_7673,N_4190,N_867);
nor U7674 (N_7674,N_3540,N_454);
nand U7675 (N_7675,N_553,N_2485);
nand U7676 (N_7676,N_1043,N_3295);
nor U7677 (N_7677,N_2123,N_810);
xnor U7678 (N_7678,N_4517,N_4270);
and U7679 (N_7679,N_3758,N_554);
nand U7680 (N_7680,N_385,N_3852);
or U7681 (N_7681,N_1085,N_2412);
nor U7682 (N_7682,N_1971,N_2308);
and U7683 (N_7683,N_2629,N_4863);
or U7684 (N_7684,N_4421,N_3999);
nand U7685 (N_7685,N_2096,N_2195);
nor U7686 (N_7686,N_969,N_4331);
nor U7687 (N_7687,N_3394,N_4929);
nand U7688 (N_7688,N_4973,N_1769);
or U7689 (N_7689,N_1562,N_2307);
or U7690 (N_7690,N_4919,N_2317);
or U7691 (N_7691,N_2535,N_1295);
or U7692 (N_7692,N_1210,N_1977);
nor U7693 (N_7693,N_131,N_4664);
and U7694 (N_7694,N_211,N_816);
and U7695 (N_7695,N_2925,N_2059);
nor U7696 (N_7696,N_4317,N_3285);
nand U7697 (N_7697,N_3348,N_640);
and U7698 (N_7698,N_4949,N_2312);
and U7699 (N_7699,N_2188,N_1573);
nor U7700 (N_7700,N_498,N_359);
or U7701 (N_7701,N_4749,N_931);
or U7702 (N_7702,N_794,N_3490);
or U7703 (N_7703,N_1659,N_2198);
and U7704 (N_7704,N_781,N_4932);
nor U7705 (N_7705,N_970,N_4936);
and U7706 (N_7706,N_2826,N_3874);
or U7707 (N_7707,N_3560,N_630);
and U7708 (N_7708,N_2882,N_3219);
xnor U7709 (N_7709,N_4136,N_676);
nor U7710 (N_7710,N_3326,N_1164);
nand U7711 (N_7711,N_2532,N_2499);
nor U7712 (N_7712,N_181,N_3965);
nor U7713 (N_7713,N_4687,N_783);
nor U7714 (N_7714,N_4855,N_620);
nor U7715 (N_7715,N_850,N_2995);
nand U7716 (N_7716,N_3829,N_2176);
nand U7717 (N_7717,N_3128,N_2381);
nand U7718 (N_7718,N_2189,N_1620);
or U7719 (N_7719,N_341,N_1317);
nand U7720 (N_7720,N_1704,N_2959);
or U7721 (N_7721,N_4532,N_3650);
or U7722 (N_7722,N_1735,N_3989);
and U7723 (N_7723,N_3055,N_2005);
nand U7724 (N_7724,N_4524,N_2294);
or U7725 (N_7725,N_3793,N_4276);
nand U7726 (N_7726,N_2656,N_3537);
or U7727 (N_7727,N_4576,N_4176);
nor U7728 (N_7728,N_3358,N_4993);
xor U7729 (N_7729,N_1764,N_2277);
nor U7730 (N_7730,N_4698,N_3104);
nand U7731 (N_7731,N_1756,N_3988);
and U7732 (N_7732,N_1956,N_2512);
or U7733 (N_7733,N_276,N_2286);
nor U7734 (N_7734,N_1259,N_3826);
nor U7735 (N_7735,N_3761,N_3849);
nor U7736 (N_7736,N_2220,N_3497);
nor U7737 (N_7737,N_134,N_2155);
or U7738 (N_7738,N_4680,N_2946);
or U7739 (N_7739,N_4383,N_4149);
and U7740 (N_7740,N_3870,N_3278);
nand U7741 (N_7741,N_1109,N_2177);
or U7742 (N_7742,N_1485,N_2050);
nor U7743 (N_7743,N_4460,N_4881);
and U7744 (N_7744,N_1664,N_3663);
and U7745 (N_7745,N_351,N_3422);
or U7746 (N_7746,N_4119,N_1754);
and U7747 (N_7747,N_2787,N_1548);
and U7748 (N_7748,N_4210,N_3019);
nand U7749 (N_7749,N_909,N_328);
or U7750 (N_7750,N_2555,N_3689);
xor U7751 (N_7751,N_3507,N_2393);
and U7752 (N_7752,N_4424,N_1005);
and U7753 (N_7753,N_3600,N_4348);
nand U7754 (N_7754,N_1614,N_3013);
and U7755 (N_7755,N_53,N_395);
and U7756 (N_7756,N_4426,N_377);
or U7757 (N_7757,N_2557,N_4279);
nand U7758 (N_7758,N_2200,N_1662);
or U7759 (N_7759,N_1525,N_1527);
nor U7760 (N_7760,N_3886,N_3057);
or U7761 (N_7761,N_2150,N_1506);
nor U7762 (N_7762,N_3052,N_2025);
nand U7763 (N_7763,N_1156,N_2416);
nor U7764 (N_7764,N_2225,N_1680);
xor U7765 (N_7765,N_137,N_3665);
and U7766 (N_7766,N_1072,N_3786);
and U7767 (N_7767,N_4883,N_14);
or U7768 (N_7768,N_3415,N_728);
nor U7769 (N_7769,N_1046,N_1404);
or U7770 (N_7770,N_3004,N_3177);
and U7771 (N_7771,N_2050,N_524);
and U7772 (N_7772,N_3284,N_963);
nor U7773 (N_7773,N_2078,N_3877);
and U7774 (N_7774,N_2213,N_3383);
nor U7775 (N_7775,N_4161,N_4814);
and U7776 (N_7776,N_2603,N_4323);
and U7777 (N_7777,N_1779,N_4512);
nor U7778 (N_7778,N_4635,N_1393);
nand U7779 (N_7779,N_2453,N_1850);
or U7780 (N_7780,N_1589,N_3391);
or U7781 (N_7781,N_132,N_577);
nor U7782 (N_7782,N_4911,N_2394);
nand U7783 (N_7783,N_4094,N_1872);
and U7784 (N_7784,N_4607,N_1033);
nor U7785 (N_7785,N_3930,N_4063);
and U7786 (N_7786,N_38,N_2184);
or U7787 (N_7787,N_214,N_3356);
nand U7788 (N_7788,N_1311,N_2203);
nor U7789 (N_7789,N_3374,N_2827);
and U7790 (N_7790,N_332,N_2104);
nor U7791 (N_7791,N_106,N_4228);
nand U7792 (N_7792,N_1948,N_2347);
or U7793 (N_7793,N_403,N_4176);
nor U7794 (N_7794,N_1078,N_3758);
and U7795 (N_7795,N_688,N_3766);
and U7796 (N_7796,N_3075,N_4419);
and U7797 (N_7797,N_3825,N_2587);
or U7798 (N_7798,N_585,N_977);
nand U7799 (N_7799,N_2396,N_2036);
or U7800 (N_7800,N_4521,N_1963);
and U7801 (N_7801,N_1373,N_1744);
or U7802 (N_7802,N_191,N_4024);
nand U7803 (N_7803,N_881,N_4654);
and U7804 (N_7804,N_3130,N_2199);
and U7805 (N_7805,N_1944,N_1605);
or U7806 (N_7806,N_3047,N_2254);
nand U7807 (N_7807,N_4354,N_1202);
nand U7808 (N_7808,N_4052,N_4207);
or U7809 (N_7809,N_98,N_1939);
nand U7810 (N_7810,N_4923,N_4170);
nand U7811 (N_7811,N_3354,N_4766);
nand U7812 (N_7812,N_39,N_2699);
nand U7813 (N_7813,N_4206,N_3431);
nor U7814 (N_7814,N_1064,N_1395);
or U7815 (N_7815,N_3346,N_127);
nor U7816 (N_7816,N_3160,N_3519);
and U7817 (N_7817,N_3708,N_1548);
xnor U7818 (N_7818,N_4827,N_4989);
nand U7819 (N_7819,N_1584,N_4166);
nand U7820 (N_7820,N_2966,N_3244);
and U7821 (N_7821,N_845,N_2307);
nand U7822 (N_7822,N_175,N_295);
or U7823 (N_7823,N_4574,N_1298);
and U7824 (N_7824,N_4581,N_1560);
and U7825 (N_7825,N_4832,N_1294);
nand U7826 (N_7826,N_3465,N_2820);
or U7827 (N_7827,N_3510,N_2676);
nand U7828 (N_7828,N_3107,N_4712);
nand U7829 (N_7829,N_2127,N_1498);
nand U7830 (N_7830,N_1075,N_4886);
nor U7831 (N_7831,N_853,N_3955);
xnor U7832 (N_7832,N_4979,N_1981);
nand U7833 (N_7833,N_60,N_3433);
or U7834 (N_7834,N_4801,N_1767);
or U7835 (N_7835,N_3118,N_292);
xnor U7836 (N_7836,N_2902,N_3403);
nor U7837 (N_7837,N_2889,N_1007);
and U7838 (N_7838,N_2642,N_2067);
and U7839 (N_7839,N_4091,N_3186);
and U7840 (N_7840,N_378,N_3083);
or U7841 (N_7841,N_4318,N_1837);
nor U7842 (N_7842,N_3692,N_4319);
nand U7843 (N_7843,N_133,N_685);
and U7844 (N_7844,N_4647,N_2006);
nor U7845 (N_7845,N_3255,N_2575);
and U7846 (N_7846,N_94,N_447);
nor U7847 (N_7847,N_4243,N_3793);
nor U7848 (N_7848,N_4848,N_1270);
or U7849 (N_7849,N_929,N_3375);
nand U7850 (N_7850,N_4829,N_2736);
and U7851 (N_7851,N_773,N_1009);
or U7852 (N_7852,N_2659,N_3693);
or U7853 (N_7853,N_3347,N_3972);
nand U7854 (N_7854,N_3677,N_4258);
and U7855 (N_7855,N_589,N_2758);
or U7856 (N_7856,N_1830,N_4214);
and U7857 (N_7857,N_330,N_1037);
or U7858 (N_7858,N_2746,N_2748);
nand U7859 (N_7859,N_2208,N_1359);
and U7860 (N_7860,N_2487,N_3061);
nor U7861 (N_7861,N_2004,N_3216);
nor U7862 (N_7862,N_510,N_3425);
nand U7863 (N_7863,N_2171,N_4245);
nor U7864 (N_7864,N_4432,N_3344);
or U7865 (N_7865,N_546,N_1250);
and U7866 (N_7866,N_2582,N_778);
nand U7867 (N_7867,N_2774,N_2230);
or U7868 (N_7868,N_3311,N_2497);
or U7869 (N_7869,N_3480,N_4131);
nand U7870 (N_7870,N_4349,N_3340);
and U7871 (N_7871,N_2476,N_3331);
and U7872 (N_7872,N_2538,N_452);
nor U7873 (N_7873,N_3614,N_1810);
or U7874 (N_7874,N_2565,N_2864);
nor U7875 (N_7875,N_1400,N_4791);
nor U7876 (N_7876,N_3545,N_2969);
nor U7877 (N_7877,N_2316,N_8);
and U7878 (N_7878,N_1520,N_442);
and U7879 (N_7879,N_434,N_2201);
nand U7880 (N_7880,N_2905,N_4177);
and U7881 (N_7881,N_2630,N_495);
nand U7882 (N_7882,N_4678,N_166);
nand U7883 (N_7883,N_3482,N_3608);
or U7884 (N_7884,N_104,N_98);
nor U7885 (N_7885,N_1315,N_2500);
and U7886 (N_7886,N_4234,N_3359);
and U7887 (N_7887,N_286,N_304);
xor U7888 (N_7888,N_1753,N_2470);
nor U7889 (N_7889,N_1060,N_286);
nor U7890 (N_7890,N_708,N_4033);
nor U7891 (N_7891,N_4113,N_4225);
and U7892 (N_7892,N_444,N_3479);
nand U7893 (N_7893,N_904,N_714);
nor U7894 (N_7894,N_4353,N_774);
nand U7895 (N_7895,N_1550,N_3298);
or U7896 (N_7896,N_568,N_4624);
and U7897 (N_7897,N_2091,N_720);
and U7898 (N_7898,N_355,N_2304);
nand U7899 (N_7899,N_364,N_2835);
nor U7900 (N_7900,N_4149,N_4882);
nand U7901 (N_7901,N_1513,N_3910);
nand U7902 (N_7902,N_550,N_4515);
or U7903 (N_7903,N_2533,N_876);
nand U7904 (N_7904,N_1589,N_4523);
nor U7905 (N_7905,N_1707,N_2784);
and U7906 (N_7906,N_1141,N_427);
nor U7907 (N_7907,N_3928,N_4010);
nor U7908 (N_7908,N_2250,N_4762);
xor U7909 (N_7909,N_2251,N_2656);
and U7910 (N_7910,N_1558,N_2767);
or U7911 (N_7911,N_4439,N_1508);
or U7912 (N_7912,N_4447,N_3724);
or U7913 (N_7913,N_3274,N_4115);
and U7914 (N_7914,N_3418,N_1232);
nand U7915 (N_7915,N_3674,N_3640);
nand U7916 (N_7916,N_4338,N_1536);
nor U7917 (N_7917,N_12,N_4773);
nand U7918 (N_7918,N_3947,N_1240);
and U7919 (N_7919,N_3637,N_3652);
and U7920 (N_7920,N_4812,N_3576);
nand U7921 (N_7921,N_141,N_3495);
nor U7922 (N_7922,N_84,N_632);
nand U7923 (N_7923,N_4261,N_810);
nand U7924 (N_7924,N_2369,N_1295);
nor U7925 (N_7925,N_1097,N_318);
nor U7926 (N_7926,N_3018,N_4295);
and U7927 (N_7927,N_3651,N_4635);
and U7928 (N_7928,N_4655,N_4723);
nor U7929 (N_7929,N_4971,N_2304);
or U7930 (N_7930,N_1392,N_4080);
nand U7931 (N_7931,N_1933,N_142);
nand U7932 (N_7932,N_1935,N_2782);
or U7933 (N_7933,N_899,N_632);
nand U7934 (N_7934,N_3616,N_3461);
nand U7935 (N_7935,N_292,N_327);
nor U7936 (N_7936,N_4448,N_1697);
nor U7937 (N_7937,N_2066,N_4968);
or U7938 (N_7938,N_1330,N_4871);
nor U7939 (N_7939,N_2560,N_4082);
and U7940 (N_7940,N_3716,N_2824);
nor U7941 (N_7941,N_3223,N_2968);
nor U7942 (N_7942,N_1550,N_384);
and U7943 (N_7943,N_4736,N_3637);
and U7944 (N_7944,N_4843,N_3600);
nor U7945 (N_7945,N_2172,N_3449);
nor U7946 (N_7946,N_3706,N_1536);
nand U7947 (N_7947,N_1366,N_2193);
or U7948 (N_7948,N_877,N_4703);
and U7949 (N_7949,N_2592,N_3267);
nor U7950 (N_7950,N_3966,N_3610);
nand U7951 (N_7951,N_78,N_4468);
and U7952 (N_7952,N_1683,N_3656);
or U7953 (N_7953,N_2898,N_1514);
nor U7954 (N_7954,N_2931,N_4364);
nor U7955 (N_7955,N_1873,N_286);
xnor U7956 (N_7956,N_2972,N_1946);
and U7957 (N_7957,N_2724,N_259);
nand U7958 (N_7958,N_4878,N_2220);
and U7959 (N_7959,N_531,N_1189);
and U7960 (N_7960,N_39,N_478);
and U7961 (N_7961,N_1266,N_4493);
nand U7962 (N_7962,N_4440,N_3205);
nand U7963 (N_7963,N_1097,N_2938);
and U7964 (N_7964,N_4583,N_2789);
nand U7965 (N_7965,N_2098,N_4166);
or U7966 (N_7966,N_9,N_1564);
nand U7967 (N_7967,N_3971,N_2185);
nor U7968 (N_7968,N_3055,N_1850);
nand U7969 (N_7969,N_4330,N_282);
or U7970 (N_7970,N_509,N_1698);
and U7971 (N_7971,N_3272,N_4552);
or U7972 (N_7972,N_2412,N_2675);
nor U7973 (N_7973,N_1244,N_281);
and U7974 (N_7974,N_2522,N_4614);
nand U7975 (N_7975,N_2467,N_2313);
and U7976 (N_7976,N_2783,N_3046);
or U7977 (N_7977,N_1507,N_4735);
nor U7978 (N_7978,N_2865,N_1928);
or U7979 (N_7979,N_872,N_3159);
nor U7980 (N_7980,N_3648,N_4414);
or U7981 (N_7981,N_721,N_2561);
xnor U7982 (N_7982,N_2911,N_2746);
or U7983 (N_7983,N_3046,N_409);
nand U7984 (N_7984,N_1758,N_3140);
nor U7985 (N_7985,N_4603,N_2198);
xnor U7986 (N_7986,N_4812,N_3014);
and U7987 (N_7987,N_2252,N_3471);
nand U7988 (N_7988,N_177,N_1654);
nor U7989 (N_7989,N_2343,N_451);
nor U7990 (N_7990,N_3604,N_4320);
and U7991 (N_7991,N_1185,N_749);
or U7992 (N_7992,N_4916,N_72);
or U7993 (N_7993,N_3198,N_1557);
nand U7994 (N_7994,N_2505,N_378);
or U7995 (N_7995,N_3892,N_2608);
nand U7996 (N_7996,N_3447,N_732);
or U7997 (N_7997,N_1537,N_2369);
or U7998 (N_7998,N_3057,N_2353);
or U7999 (N_7999,N_1850,N_1262);
or U8000 (N_8000,N_1181,N_1052);
and U8001 (N_8001,N_2501,N_355);
nor U8002 (N_8002,N_4581,N_3054);
nand U8003 (N_8003,N_2348,N_3399);
or U8004 (N_8004,N_1603,N_4834);
and U8005 (N_8005,N_242,N_3383);
nand U8006 (N_8006,N_3211,N_1307);
and U8007 (N_8007,N_4755,N_192);
or U8008 (N_8008,N_3260,N_411);
nand U8009 (N_8009,N_4879,N_983);
nor U8010 (N_8010,N_3526,N_1240);
or U8011 (N_8011,N_1490,N_2297);
and U8012 (N_8012,N_2167,N_3067);
nor U8013 (N_8013,N_2580,N_4444);
nor U8014 (N_8014,N_4726,N_4052);
nor U8015 (N_8015,N_2666,N_2711);
and U8016 (N_8016,N_3148,N_3352);
or U8017 (N_8017,N_3051,N_3998);
or U8018 (N_8018,N_4465,N_1606);
or U8019 (N_8019,N_1457,N_2472);
nand U8020 (N_8020,N_1135,N_898);
or U8021 (N_8021,N_1766,N_1688);
nor U8022 (N_8022,N_2418,N_1778);
nor U8023 (N_8023,N_38,N_2801);
or U8024 (N_8024,N_3000,N_4365);
nor U8025 (N_8025,N_1119,N_2860);
nor U8026 (N_8026,N_1835,N_3092);
nor U8027 (N_8027,N_3540,N_1728);
nand U8028 (N_8028,N_2790,N_2964);
nand U8029 (N_8029,N_982,N_46);
nand U8030 (N_8030,N_688,N_1542);
and U8031 (N_8031,N_4516,N_1846);
and U8032 (N_8032,N_934,N_2440);
nand U8033 (N_8033,N_3721,N_3693);
nor U8034 (N_8034,N_4841,N_3669);
or U8035 (N_8035,N_4013,N_4332);
nor U8036 (N_8036,N_1018,N_3085);
nand U8037 (N_8037,N_1770,N_2971);
nand U8038 (N_8038,N_3094,N_4514);
and U8039 (N_8039,N_4705,N_4823);
nor U8040 (N_8040,N_4536,N_3192);
or U8041 (N_8041,N_4458,N_3026);
and U8042 (N_8042,N_4755,N_2692);
or U8043 (N_8043,N_1760,N_1407);
and U8044 (N_8044,N_2573,N_215);
or U8045 (N_8045,N_477,N_648);
xor U8046 (N_8046,N_2040,N_3073);
or U8047 (N_8047,N_4269,N_944);
nand U8048 (N_8048,N_2735,N_1761);
nand U8049 (N_8049,N_962,N_4206);
nor U8050 (N_8050,N_236,N_943);
or U8051 (N_8051,N_3126,N_3891);
nand U8052 (N_8052,N_222,N_3688);
and U8053 (N_8053,N_1547,N_1916);
and U8054 (N_8054,N_4717,N_4267);
nor U8055 (N_8055,N_2509,N_2642);
and U8056 (N_8056,N_1739,N_2059);
or U8057 (N_8057,N_2598,N_4221);
nor U8058 (N_8058,N_2870,N_4279);
nor U8059 (N_8059,N_2753,N_1182);
nor U8060 (N_8060,N_4987,N_1945);
nand U8061 (N_8061,N_4338,N_4119);
nand U8062 (N_8062,N_210,N_4835);
and U8063 (N_8063,N_1934,N_2955);
or U8064 (N_8064,N_3147,N_2328);
or U8065 (N_8065,N_4569,N_1868);
or U8066 (N_8066,N_1622,N_1706);
nor U8067 (N_8067,N_3894,N_3251);
nor U8068 (N_8068,N_3394,N_1847);
and U8069 (N_8069,N_1867,N_2042);
nor U8070 (N_8070,N_1893,N_3082);
and U8071 (N_8071,N_2170,N_3299);
nand U8072 (N_8072,N_3863,N_2771);
or U8073 (N_8073,N_522,N_3526);
nor U8074 (N_8074,N_1296,N_2572);
and U8075 (N_8075,N_2504,N_1391);
nor U8076 (N_8076,N_4841,N_4063);
nor U8077 (N_8077,N_315,N_791);
or U8078 (N_8078,N_942,N_2074);
nand U8079 (N_8079,N_3353,N_1997);
or U8080 (N_8080,N_595,N_4755);
or U8081 (N_8081,N_44,N_2946);
or U8082 (N_8082,N_1501,N_2946);
and U8083 (N_8083,N_4908,N_1810);
and U8084 (N_8084,N_788,N_232);
nor U8085 (N_8085,N_3889,N_1970);
and U8086 (N_8086,N_3745,N_2679);
nor U8087 (N_8087,N_3474,N_3478);
nand U8088 (N_8088,N_2737,N_3375);
and U8089 (N_8089,N_4687,N_4210);
or U8090 (N_8090,N_1404,N_4569);
nand U8091 (N_8091,N_2506,N_371);
or U8092 (N_8092,N_4985,N_3770);
and U8093 (N_8093,N_4825,N_3400);
nand U8094 (N_8094,N_4518,N_4711);
and U8095 (N_8095,N_2083,N_2244);
or U8096 (N_8096,N_4168,N_2439);
or U8097 (N_8097,N_1329,N_3535);
and U8098 (N_8098,N_3450,N_503);
and U8099 (N_8099,N_2927,N_2246);
nor U8100 (N_8100,N_4871,N_1599);
nand U8101 (N_8101,N_2193,N_1415);
or U8102 (N_8102,N_3533,N_2186);
or U8103 (N_8103,N_2143,N_2717);
and U8104 (N_8104,N_2985,N_2082);
nand U8105 (N_8105,N_3423,N_838);
and U8106 (N_8106,N_2353,N_3538);
and U8107 (N_8107,N_3104,N_4265);
or U8108 (N_8108,N_581,N_4890);
and U8109 (N_8109,N_4282,N_491);
and U8110 (N_8110,N_3671,N_4878);
nand U8111 (N_8111,N_2118,N_302);
nor U8112 (N_8112,N_1894,N_4567);
nand U8113 (N_8113,N_3603,N_1449);
or U8114 (N_8114,N_659,N_4473);
or U8115 (N_8115,N_1833,N_260);
or U8116 (N_8116,N_4138,N_1888);
or U8117 (N_8117,N_4986,N_3188);
and U8118 (N_8118,N_3929,N_4740);
nor U8119 (N_8119,N_1665,N_662);
nand U8120 (N_8120,N_2733,N_1164);
nor U8121 (N_8121,N_1886,N_4059);
nor U8122 (N_8122,N_264,N_4141);
nand U8123 (N_8123,N_2903,N_2533);
and U8124 (N_8124,N_2677,N_1368);
nand U8125 (N_8125,N_820,N_2639);
xnor U8126 (N_8126,N_4206,N_3348);
nand U8127 (N_8127,N_2063,N_3358);
or U8128 (N_8128,N_4477,N_3588);
nor U8129 (N_8129,N_1168,N_1214);
nand U8130 (N_8130,N_23,N_3522);
or U8131 (N_8131,N_994,N_3116);
nor U8132 (N_8132,N_4519,N_2298);
or U8133 (N_8133,N_2261,N_4650);
nor U8134 (N_8134,N_67,N_2410);
xor U8135 (N_8135,N_1316,N_3403);
or U8136 (N_8136,N_2875,N_3859);
or U8137 (N_8137,N_4152,N_4367);
nor U8138 (N_8138,N_13,N_4240);
nor U8139 (N_8139,N_645,N_3868);
nand U8140 (N_8140,N_3856,N_1949);
nand U8141 (N_8141,N_3314,N_405);
nand U8142 (N_8142,N_2727,N_4096);
or U8143 (N_8143,N_1816,N_2958);
or U8144 (N_8144,N_4229,N_2354);
nand U8145 (N_8145,N_3287,N_3047);
nor U8146 (N_8146,N_4162,N_3036);
or U8147 (N_8147,N_1998,N_2081);
nand U8148 (N_8148,N_3025,N_1070);
nand U8149 (N_8149,N_4030,N_277);
or U8150 (N_8150,N_930,N_2410);
nand U8151 (N_8151,N_3954,N_746);
and U8152 (N_8152,N_2584,N_2801);
or U8153 (N_8153,N_4104,N_1247);
nand U8154 (N_8154,N_3173,N_1163);
or U8155 (N_8155,N_318,N_180);
and U8156 (N_8156,N_2377,N_756);
or U8157 (N_8157,N_1686,N_3510);
nand U8158 (N_8158,N_1799,N_2434);
nand U8159 (N_8159,N_3691,N_3420);
and U8160 (N_8160,N_2633,N_2913);
nor U8161 (N_8161,N_3969,N_482);
and U8162 (N_8162,N_1835,N_4028);
or U8163 (N_8163,N_4309,N_2567);
nand U8164 (N_8164,N_2407,N_3202);
and U8165 (N_8165,N_749,N_2921);
nor U8166 (N_8166,N_4242,N_4287);
and U8167 (N_8167,N_952,N_2115);
nand U8168 (N_8168,N_146,N_238);
nor U8169 (N_8169,N_4482,N_2877);
nand U8170 (N_8170,N_909,N_2703);
or U8171 (N_8171,N_4738,N_702);
nand U8172 (N_8172,N_1268,N_3268);
nand U8173 (N_8173,N_175,N_3074);
or U8174 (N_8174,N_41,N_1993);
nand U8175 (N_8175,N_2457,N_1218);
nand U8176 (N_8176,N_1074,N_2733);
nor U8177 (N_8177,N_894,N_3852);
and U8178 (N_8178,N_865,N_4910);
and U8179 (N_8179,N_1740,N_3013);
and U8180 (N_8180,N_2992,N_3408);
and U8181 (N_8181,N_3279,N_2027);
nor U8182 (N_8182,N_2389,N_4500);
nor U8183 (N_8183,N_2278,N_290);
nor U8184 (N_8184,N_4502,N_210);
or U8185 (N_8185,N_2912,N_581);
nor U8186 (N_8186,N_4828,N_3564);
nand U8187 (N_8187,N_1159,N_4956);
or U8188 (N_8188,N_3313,N_4928);
or U8189 (N_8189,N_3969,N_294);
nor U8190 (N_8190,N_708,N_4279);
xnor U8191 (N_8191,N_2361,N_569);
and U8192 (N_8192,N_919,N_2431);
or U8193 (N_8193,N_4528,N_2513);
nand U8194 (N_8194,N_300,N_4867);
nor U8195 (N_8195,N_4302,N_4899);
nor U8196 (N_8196,N_401,N_4774);
nor U8197 (N_8197,N_4288,N_3245);
nand U8198 (N_8198,N_167,N_1858);
or U8199 (N_8199,N_2029,N_570);
nand U8200 (N_8200,N_1747,N_2682);
or U8201 (N_8201,N_663,N_1576);
or U8202 (N_8202,N_3849,N_799);
or U8203 (N_8203,N_1849,N_4330);
nor U8204 (N_8204,N_4373,N_2796);
or U8205 (N_8205,N_3241,N_3657);
nor U8206 (N_8206,N_3348,N_1887);
nand U8207 (N_8207,N_2950,N_2776);
nor U8208 (N_8208,N_4631,N_1124);
nor U8209 (N_8209,N_1706,N_4700);
nor U8210 (N_8210,N_4007,N_4097);
nand U8211 (N_8211,N_4609,N_4805);
nand U8212 (N_8212,N_956,N_1080);
and U8213 (N_8213,N_4345,N_2668);
and U8214 (N_8214,N_2230,N_1457);
and U8215 (N_8215,N_2240,N_938);
nor U8216 (N_8216,N_26,N_3035);
nor U8217 (N_8217,N_1524,N_4141);
or U8218 (N_8218,N_4896,N_1473);
and U8219 (N_8219,N_685,N_752);
and U8220 (N_8220,N_687,N_3688);
nand U8221 (N_8221,N_1172,N_1424);
nand U8222 (N_8222,N_3202,N_2208);
nand U8223 (N_8223,N_187,N_275);
and U8224 (N_8224,N_1615,N_70);
or U8225 (N_8225,N_1455,N_1464);
nand U8226 (N_8226,N_402,N_1903);
or U8227 (N_8227,N_2760,N_1902);
or U8228 (N_8228,N_2969,N_3365);
nor U8229 (N_8229,N_3185,N_1870);
or U8230 (N_8230,N_3516,N_1457);
nand U8231 (N_8231,N_4352,N_4278);
nand U8232 (N_8232,N_391,N_4022);
and U8233 (N_8233,N_100,N_2263);
or U8234 (N_8234,N_3182,N_3395);
nor U8235 (N_8235,N_4056,N_3471);
nand U8236 (N_8236,N_4369,N_2098);
nand U8237 (N_8237,N_3212,N_4968);
or U8238 (N_8238,N_4834,N_252);
and U8239 (N_8239,N_949,N_2733);
and U8240 (N_8240,N_3895,N_1719);
nand U8241 (N_8241,N_3812,N_3807);
nand U8242 (N_8242,N_823,N_1461);
nor U8243 (N_8243,N_3366,N_1924);
and U8244 (N_8244,N_1657,N_3931);
nand U8245 (N_8245,N_922,N_2315);
nand U8246 (N_8246,N_2940,N_3332);
nor U8247 (N_8247,N_1467,N_98);
or U8248 (N_8248,N_1594,N_3794);
nand U8249 (N_8249,N_3475,N_2193);
nand U8250 (N_8250,N_1717,N_1685);
and U8251 (N_8251,N_4385,N_4409);
or U8252 (N_8252,N_793,N_1965);
and U8253 (N_8253,N_3291,N_4471);
or U8254 (N_8254,N_3330,N_3358);
xnor U8255 (N_8255,N_2805,N_3627);
nor U8256 (N_8256,N_4406,N_2477);
nor U8257 (N_8257,N_1014,N_4466);
nor U8258 (N_8258,N_525,N_3306);
nor U8259 (N_8259,N_3600,N_1302);
or U8260 (N_8260,N_956,N_3605);
or U8261 (N_8261,N_4090,N_1114);
and U8262 (N_8262,N_4411,N_1040);
and U8263 (N_8263,N_4559,N_3936);
and U8264 (N_8264,N_2404,N_704);
nand U8265 (N_8265,N_138,N_615);
nor U8266 (N_8266,N_4725,N_2915);
nor U8267 (N_8267,N_140,N_4833);
or U8268 (N_8268,N_754,N_1723);
or U8269 (N_8269,N_301,N_2307);
nand U8270 (N_8270,N_2663,N_2887);
nor U8271 (N_8271,N_3069,N_3929);
and U8272 (N_8272,N_4885,N_1253);
and U8273 (N_8273,N_2540,N_4239);
nor U8274 (N_8274,N_766,N_1654);
and U8275 (N_8275,N_769,N_2030);
or U8276 (N_8276,N_3159,N_765);
or U8277 (N_8277,N_4641,N_4776);
nor U8278 (N_8278,N_4704,N_628);
nand U8279 (N_8279,N_2014,N_2367);
and U8280 (N_8280,N_4653,N_885);
nor U8281 (N_8281,N_671,N_3640);
nand U8282 (N_8282,N_4282,N_3825);
and U8283 (N_8283,N_4651,N_32);
nand U8284 (N_8284,N_4534,N_526);
and U8285 (N_8285,N_4040,N_3976);
and U8286 (N_8286,N_3792,N_3858);
nor U8287 (N_8287,N_2098,N_1749);
and U8288 (N_8288,N_4877,N_170);
or U8289 (N_8289,N_1193,N_2563);
nor U8290 (N_8290,N_2568,N_2647);
nand U8291 (N_8291,N_676,N_693);
nand U8292 (N_8292,N_3951,N_2963);
or U8293 (N_8293,N_2678,N_1594);
and U8294 (N_8294,N_3554,N_2372);
and U8295 (N_8295,N_333,N_4673);
nor U8296 (N_8296,N_1299,N_3512);
nor U8297 (N_8297,N_4515,N_638);
xnor U8298 (N_8298,N_1796,N_589);
nor U8299 (N_8299,N_606,N_2942);
and U8300 (N_8300,N_2174,N_1101);
and U8301 (N_8301,N_4682,N_691);
and U8302 (N_8302,N_1659,N_997);
nand U8303 (N_8303,N_949,N_1787);
nand U8304 (N_8304,N_2496,N_2328);
nand U8305 (N_8305,N_1126,N_1894);
nand U8306 (N_8306,N_2426,N_711);
and U8307 (N_8307,N_4696,N_2611);
or U8308 (N_8308,N_2963,N_414);
nand U8309 (N_8309,N_2399,N_2791);
and U8310 (N_8310,N_815,N_4915);
or U8311 (N_8311,N_2674,N_1847);
and U8312 (N_8312,N_1101,N_4983);
nor U8313 (N_8313,N_2108,N_1959);
nor U8314 (N_8314,N_1884,N_1966);
nor U8315 (N_8315,N_3218,N_1741);
and U8316 (N_8316,N_2701,N_487);
and U8317 (N_8317,N_2007,N_3694);
nor U8318 (N_8318,N_3273,N_4042);
xor U8319 (N_8319,N_3386,N_2933);
and U8320 (N_8320,N_4614,N_1612);
nand U8321 (N_8321,N_4596,N_1200);
nor U8322 (N_8322,N_2209,N_1281);
nand U8323 (N_8323,N_937,N_1342);
nor U8324 (N_8324,N_3470,N_287);
and U8325 (N_8325,N_998,N_4971);
nand U8326 (N_8326,N_415,N_808);
nor U8327 (N_8327,N_1231,N_3730);
or U8328 (N_8328,N_1332,N_3278);
or U8329 (N_8329,N_1258,N_4825);
or U8330 (N_8330,N_2101,N_4451);
nand U8331 (N_8331,N_848,N_2427);
nor U8332 (N_8332,N_172,N_827);
nor U8333 (N_8333,N_2291,N_3373);
nand U8334 (N_8334,N_1432,N_47);
or U8335 (N_8335,N_539,N_3419);
xor U8336 (N_8336,N_4100,N_373);
or U8337 (N_8337,N_1025,N_4087);
or U8338 (N_8338,N_2606,N_215);
and U8339 (N_8339,N_4615,N_2419);
nor U8340 (N_8340,N_4738,N_2547);
nor U8341 (N_8341,N_3105,N_922);
nor U8342 (N_8342,N_2613,N_1772);
nand U8343 (N_8343,N_4594,N_1076);
nand U8344 (N_8344,N_506,N_3032);
or U8345 (N_8345,N_1768,N_1522);
and U8346 (N_8346,N_1258,N_4237);
nand U8347 (N_8347,N_4672,N_4267);
and U8348 (N_8348,N_4227,N_3046);
or U8349 (N_8349,N_3490,N_1898);
or U8350 (N_8350,N_4161,N_3545);
nor U8351 (N_8351,N_2539,N_1046);
xnor U8352 (N_8352,N_3826,N_2229);
nand U8353 (N_8353,N_1219,N_1676);
nand U8354 (N_8354,N_4336,N_2842);
xnor U8355 (N_8355,N_3632,N_1285);
and U8356 (N_8356,N_944,N_1101);
nor U8357 (N_8357,N_4662,N_2724);
nand U8358 (N_8358,N_3194,N_1515);
or U8359 (N_8359,N_4920,N_1651);
and U8360 (N_8360,N_4091,N_850);
and U8361 (N_8361,N_4937,N_2827);
or U8362 (N_8362,N_910,N_2482);
and U8363 (N_8363,N_4754,N_1215);
or U8364 (N_8364,N_1822,N_3575);
nand U8365 (N_8365,N_935,N_1859);
and U8366 (N_8366,N_4577,N_3379);
nor U8367 (N_8367,N_253,N_400);
nand U8368 (N_8368,N_4036,N_3066);
and U8369 (N_8369,N_3261,N_4049);
and U8370 (N_8370,N_1822,N_3165);
and U8371 (N_8371,N_650,N_841);
nor U8372 (N_8372,N_3414,N_4805);
and U8373 (N_8373,N_952,N_1649);
or U8374 (N_8374,N_2953,N_2905);
nor U8375 (N_8375,N_2986,N_3429);
nor U8376 (N_8376,N_4613,N_3148);
nor U8377 (N_8377,N_4772,N_951);
or U8378 (N_8378,N_3718,N_1367);
or U8379 (N_8379,N_1493,N_4318);
and U8380 (N_8380,N_2583,N_2719);
nor U8381 (N_8381,N_4756,N_1691);
nand U8382 (N_8382,N_4755,N_169);
nand U8383 (N_8383,N_3374,N_2714);
or U8384 (N_8384,N_2371,N_2272);
or U8385 (N_8385,N_1670,N_3397);
or U8386 (N_8386,N_3634,N_3392);
nor U8387 (N_8387,N_2546,N_4264);
or U8388 (N_8388,N_2821,N_740);
nor U8389 (N_8389,N_1551,N_3084);
nor U8390 (N_8390,N_2642,N_2332);
nor U8391 (N_8391,N_2917,N_415);
and U8392 (N_8392,N_2583,N_1496);
or U8393 (N_8393,N_4414,N_127);
or U8394 (N_8394,N_3422,N_3148);
nand U8395 (N_8395,N_2822,N_4128);
nand U8396 (N_8396,N_1275,N_2176);
nor U8397 (N_8397,N_4774,N_4632);
nand U8398 (N_8398,N_1985,N_2194);
or U8399 (N_8399,N_4356,N_4793);
nor U8400 (N_8400,N_1473,N_384);
or U8401 (N_8401,N_1326,N_4993);
nand U8402 (N_8402,N_1104,N_3031);
or U8403 (N_8403,N_2107,N_1609);
nor U8404 (N_8404,N_15,N_3251);
and U8405 (N_8405,N_3024,N_2453);
nand U8406 (N_8406,N_1831,N_2404);
nand U8407 (N_8407,N_1458,N_1642);
nor U8408 (N_8408,N_3891,N_124);
or U8409 (N_8409,N_4394,N_781);
and U8410 (N_8410,N_2237,N_4461);
and U8411 (N_8411,N_4364,N_2737);
and U8412 (N_8412,N_2564,N_2249);
or U8413 (N_8413,N_287,N_2102);
nor U8414 (N_8414,N_269,N_4864);
and U8415 (N_8415,N_507,N_1659);
or U8416 (N_8416,N_1508,N_1887);
and U8417 (N_8417,N_1734,N_1975);
nand U8418 (N_8418,N_4964,N_3052);
nor U8419 (N_8419,N_1110,N_1345);
nor U8420 (N_8420,N_723,N_3344);
nor U8421 (N_8421,N_2594,N_3128);
or U8422 (N_8422,N_113,N_1248);
and U8423 (N_8423,N_627,N_4935);
and U8424 (N_8424,N_3712,N_784);
nor U8425 (N_8425,N_1815,N_4721);
nor U8426 (N_8426,N_3184,N_3821);
and U8427 (N_8427,N_724,N_2068);
and U8428 (N_8428,N_919,N_3212);
nor U8429 (N_8429,N_3612,N_4766);
nor U8430 (N_8430,N_1273,N_1413);
or U8431 (N_8431,N_4761,N_910);
nand U8432 (N_8432,N_1022,N_4214);
or U8433 (N_8433,N_3929,N_2080);
nand U8434 (N_8434,N_2947,N_2251);
and U8435 (N_8435,N_1224,N_4362);
and U8436 (N_8436,N_157,N_3979);
or U8437 (N_8437,N_77,N_199);
and U8438 (N_8438,N_73,N_2941);
and U8439 (N_8439,N_2442,N_314);
or U8440 (N_8440,N_1009,N_2373);
nand U8441 (N_8441,N_4167,N_3756);
nand U8442 (N_8442,N_715,N_2917);
nor U8443 (N_8443,N_3333,N_2701);
nand U8444 (N_8444,N_3335,N_3203);
nand U8445 (N_8445,N_1267,N_3300);
nand U8446 (N_8446,N_2112,N_3991);
or U8447 (N_8447,N_603,N_2440);
and U8448 (N_8448,N_4406,N_2549);
or U8449 (N_8449,N_3777,N_4364);
nor U8450 (N_8450,N_3763,N_4964);
and U8451 (N_8451,N_3543,N_983);
nand U8452 (N_8452,N_737,N_3432);
or U8453 (N_8453,N_106,N_636);
and U8454 (N_8454,N_96,N_2414);
and U8455 (N_8455,N_4216,N_1048);
and U8456 (N_8456,N_3442,N_722);
or U8457 (N_8457,N_4263,N_1625);
nand U8458 (N_8458,N_4755,N_3049);
and U8459 (N_8459,N_4443,N_3653);
xnor U8460 (N_8460,N_4737,N_1347);
nand U8461 (N_8461,N_3195,N_2774);
nor U8462 (N_8462,N_2284,N_4791);
and U8463 (N_8463,N_3582,N_3615);
nand U8464 (N_8464,N_1644,N_3819);
nor U8465 (N_8465,N_2428,N_3625);
and U8466 (N_8466,N_87,N_3427);
and U8467 (N_8467,N_3726,N_4402);
xnor U8468 (N_8468,N_2589,N_2825);
and U8469 (N_8469,N_445,N_1380);
and U8470 (N_8470,N_3250,N_478);
nor U8471 (N_8471,N_464,N_1762);
nand U8472 (N_8472,N_1643,N_1256);
nand U8473 (N_8473,N_3564,N_501);
and U8474 (N_8474,N_1891,N_4714);
nor U8475 (N_8475,N_386,N_3506);
or U8476 (N_8476,N_3359,N_4053);
or U8477 (N_8477,N_135,N_1848);
nor U8478 (N_8478,N_2214,N_115);
or U8479 (N_8479,N_3428,N_2288);
and U8480 (N_8480,N_1219,N_525);
xor U8481 (N_8481,N_948,N_939);
and U8482 (N_8482,N_515,N_3006);
xnor U8483 (N_8483,N_4666,N_822);
nor U8484 (N_8484,N_3305,N_2232);
nor U8485 (N_8485,N_560,N_572);
or U8486 (N_8486,N_3244,N_3581);
nor U8487 (N_8487,N_3679,N_546);
nand U8488 (N_8488,N_309,N_4318);
nand U8489 (N_8489,N_4537,N_4435);
and U8490 (N_8490,N_248,N_1722);
nand U8491 (N_8491,N_3962,N_3130);
nor U8492 (N_8492,N_4311,N_1629);
or U8493 (N_8493,N_4412,N_2033);
nand U8494 (N_8494,N_2698,N_3693);
nand U8495 (N_8495,N_2958,N_4672);
nand U8496 (N_8496,N_2921,N_1024);
nand U8497 (N_8497,N_4166,N_4722);
nand U8498 (N_8498,N_299,N_4498);
nand U8499 (N_8499,N_4064,N_1443);
nor U8500 (N_8500,N_91,N_3544);
xor U8501 (N_8501,N_3666,N_2157);
and U8502 (N_8502,N_2360,N_3035);
nor U8503 (N_8503,N_4288,N_3278);
or U8504 (N_8504,N_961,N_1001);
nor U8505 (N_8505,N_3469,N_3065);
nand U8506 (N_8506,N_2949,N_2625);
or U8507 (N_8507,N_1351,N_4519);
nand U8508 (N_8508,N_4702,N_3836);
or U8509 (N_8509,N_2127,N_3170);
nand U8510 (N_8510,N_1541,N_1290);
nand U8511 (N_8511,N_1857,N_2140);
xor U8512 (N_8512,N_3131,N_1960);
and U8513 (N_8513,N_3705,N_3959);
nand U8514 (N_8514,N_1871,N_501);
nand U8515 (N_8515,N_4018,N_1003);
nand U8516 (N_8516,N_1579,N_794);
nor U8517 (N_8517,N_3967,N_2092);
and U8518 (N_8518,N_932,N_54);
nand U8519 (N_8519,N_2322,N_3730);
nand U8520 (N_8520,N_557,N_1046);
and U8521 (N_8521,N_4630,N_2073);
or U8522 (N_8522,N_2125,N_3980);
nor U8523 (N_8523,N_664,N_3360);
nor U8524 (N_8524,N_1319,N_3174);
nand U8525 (N_8525,N_4127,N_3831);
nor U8526 (N_8526,N_4118,N_375);
nor U8527 (N_8527,N_686,N_4304);
nand U8528 (N_8528,N_66,N_4850);
or U8529 (N_8529,N_1801,N_2213);
nand U8530 (N_8530,N_2642,N_2513);
or U8531 (N_8531,N_802,N_1398);
nand U8532 (N_8532,N_2868,N_181);
and U8533 (N_8533,N_1906,N_558);
nand U8534 (N_8534,N_1159,N_2293);
and U8535 (N_8535,N_2212,N_267);
or U8536 (N_8536,N_2620,N_246);
and U8537 (N_8537,N_1458,N_2254);
or U8538 (N_8538,N_562,N_2261);
xor U8539 (N_8539,N_3888,N_3708);
nand U8540 (N_8540,N_1938,N_3072);
nor U8541 (N_8541,N_146,N_4122);
nand U8542 (N_8542,N_3599,N_2994);
and U8543 (N_8543,N_262,N_1922);
and U8544 (N_8544,N_1764,N_2270);
or U8545 (N_8545,N_1005,N_1345);
and U8546 (N_8546,N_3500,N_4452);
or U8547 (N_8547,N_1444,N_1445);
xnor U8548 (N_8548,N_1846,N_2178);
nor U8549 (N_8549,N_1059,N_2432);
or U8550 (N_8550,N_823,N_625);
nor U8551 (N_8551,N_260,N_1824);
nand U8552 (N_8552,N_3215,N_558);
nand U8553 (N_8553,N_1748,N_2853);
nor U8554 (N_8554,N_855,N_3965);
nor U8555 (N_8555,N_3477,N_1349);
and U8556 (N_8556,N_2271,N_1113);
nor U8557 (N_8557,N_2113,N_2063);
nor U8558 (N_8558,N_465,N_635);
or U8559 (N_8559,N_2530,N_961);
xor U8560 (N_8560,N_4960,N_3570);
nor U8561 (N_8561,N_746,N_1376);
nor U8562 (N_8562,N_1525,N_3433);
or U8563 (N_8563,N_3210,N_1409);
nand U8564 (N_8564,N_2200,N_1003);
nor U8565 (N_8565,N_2229,N_4041);
nor U8566 (N_8566,N_4576,N_2300);
and U8567 (N_8567,N_1107,N_337);
nor U8568 (N_8568,N_749,N_4443);
and U8569 (N_8569,N_4836,N_1158);
or U8570 (N_8570,N_2210,N_1971);
nand U8571 (N_8571,N_1625,N_309);
nor U8572 (N_8572,N_3115,N_3183);
nand U8573 (N_8573,N_2171,N_2918);
or U8574 (N_8574,N_3621,N_3565);
or U8575 (N_8575,N_687,N_195);
or U8576 (N_8576,N_80,N_1816);
nand U8577 (N_8577,N_638,N_2159);
and U8578 (N_8578,N_3555,N_1304);
nand U8579 (N_8579,N_4863,N_4606);
or U8580 (N_8580,N_853,N_3517);
or U8581 (N_8581,N_534,N_2520);
and U8582 (N_8582,N_4741,N_2709);
nor U8583 (N_8583,N_653,N_2963);
nor U8584 (N_8584,N_808,N_1360);
nor U8585 (N_8585,N_4163,N_4617);
nor U8586 (N_8586,N_4415,N_2223);
and U8587 (N_8587,N_2224,N_4085);
nand U8588 (N_8588,N_513,N_1376);
and U8589 (N_8589,N_2163,N_929);
nor U8590 (N_8590,N_3328,N_822);
or U8591 (N_8591,N_3408,N_3079);
or U8592 (N_8592,N_448,N_4972);
and U8593 (N_8593,N_874,N_1236);
or U8594 (N_8594,N_4171,N_3144);
and U8595 (N_8595,N_4378,N_1193);
nand U8596 (N_8596,N_4356,N_2095);
nand U8597 (N_8597,N_4532,N_4443);
xnor U8598 (N_8598,N_3220,N_2656);
and U8599 (N_8599,N_4002,N_3577);
nor U8600 (N_8600,N_1643,N_2948);
nand U8601 (N_8601,N_78,N_4466);
and U8602 (N_8602,N_258,N_2185);
or U8603 (N_8603,N_3652,N_1843);
nand U8604 (N_8604,N_3578,N_3917);
nand U8605 (N_8605,N_461,N_573);
nand U8606 (N_8606,N_1214,N_2759);
nor U8607 (N_8607,N_3341,N_80);
nand U8608 (N_8608,N_297,N_1018);
and U8609 (N_8609,N_4748,N_3677);
or U8610 (N_8610,N_4563,N_1357);
or U8611 (N_8611,N_4834,N_1954);
nor U8612 (N_8612,N_2967,N_1594);
xnor U8613 (N_8613,N_932,N_841);
and U8614 (N_8614,N_4876,N_4038);
or U8615 (N_8615,N_4080,N_1076);
nand U8616 (N_8616,N_4030,N_498);
nor U8617 (N_8617,N_4832,N_2462);
and U8618 (N_8618,N_4828,N_555);
or U8619 (N_8619,N_1070,N_4752);
xor U8620 (N_8620,N_3971,N_2758);
nor U8621 (N_8621,N_948,N_4759);
and U8622 (N_8622,N_4100,N_3888);
or U8623 (N_8623,N_3032,N_4252);
or U8624 (N_8624,N_323,N_4322);
xnor U8625 (N_8625,N_4978,N_105);
nor U8626 (N_8626,N_114,N_1081);
and U8627 (N_8627,N_1394,N_3402);
or U8628 (N_8628,N_2195,N_2688);
nor U8629 (N_8629,N_1222,N_4880);
nand U8630 (N_8630,N_2877,N_2367);
nor U8631 (N_8631,N_3647,N_2741);
or U8632 (N_8632,N_4554,N_1194);
nor U8633 (N_8633,N_2942,N_432);
or U8634 (N_8634,N_1531,N_4760);
nor U8635 (N_8635,N_370,N_4320);
nor U8636 (N_8636,N_1591,N_4494);
nor U8637 (N_8637,N_1814,N_3681);
and U8638 (N_8638,N_1861,N_1624);
nor U8639 (N_8639,N_3379,N_2792);
or U8640 (N_8640,N_3681,N_592);
nor U8641 (N_8641,N_3073,N_525);
or U8642 (N_8642,N_4343,N_985);
or U8643 (N_8643,N_3213,N_2842);
nand U8644 (N_8644,N_926,N_1731);
or U8645 (N_8645,N_3969,N_4797);
nor U8646 (N_8646,N_168,N_3833);
and U8647 (N_8647,N_4064,N_100);
nand U8648 (N_8648,N_3178,N_220);
or U8649 (N_8649,N_4077,N_4520);
nor U8650 (N_8650,N_4005,N_1811);
or U8651 (N_8651,N_1642,N_747);
and U8652 (N_8652,N_2905,N_4566);
nand U8653 (N_8653,N_978,N_3064);
or U8654 (N_8654,N_1135,N_3762);
nand U8655 (N_8655,N_3840,N_4382);
or U8656 (N_8656,N_330,N_4318);
or U8657 (N_8657,N_4738,N_2728);
nor U8658 (N_8658,N_3662,N_2897);
nand U8659 (N_8659,N_4027,N_4553);
nand U8660 (N_8660,N_2986,N_2808);
nand U8661 (N_8661,N_692,N_3480);
or U8662 (N_8662,N_2179,N_1453);
or U8663 (N_8663,N_2556,N_4654);
and U8664 (N_8664,N_2801,N_3337);
or U8665 (N_8665,N_121,N_2953);
nand U8666 (N_8666,N_604,N_4143);
nand U8667 (N_8667,N_2666,N_142);
and U8668 (N_8668,N_2221,N_3972);
xnor U8669 (N_8669,N_1952,N_3508);
or U8670 (N_8670,N_4628,N_208);
nor U8671 (N_8671,N_3716,N_1868);
and U8672 (N_8672,N_1032,N_2292);
nand U8673 (N_8673,N_3054,N_8);
or U8674 (N_8674,N_2545,N_3172);
or U8675 (N_8675,N_379,N_4269);
nor U8676 (N_8676,N_3077,N_2387);
nand U8677 (N_8677,N_47,N_3738);
xor U8678 (N_8678,N_4918,N_2015);
nand U8679 (N_8679,N_3694,N_4500);
and U8680 (N_8680,N_2467,N_460);
and U8681 (N_8681,N_2175,N_707);
nor U8682 (N_8682,N_4293,N_4177);
and U8683 (N_8683,N_3635,N_4253);
or U8684 (N_8684,N_786,N_1326);
nand U8685 (N_8685,N_1691,N_2684);
or U8686 (N_8686,N_3561,N_665);
or U8687 (N_8687,N_3418,N_194);
and U8688 (N_8688,N_4428,N_2874);
nor U8689 (N_8689,N_2579,N_3878);
nor U8690 (N_8690,N_1544,N_2846);
nand U8691 (N_8691,N_4573,N_432);
and U8692 (N_8692,N_100,N_4915);
nor U8693 (N_8693,N_2047,N_3401);
and U8694 (N_8694,N_1588,N_464);
or U8695 (N_8695,N_1167,N_1310);
nor U8696 (N_8696,N_130,N_1548);
nand U8697 (N_8697,N_4874,N_2261);
or U8698 (N_8698,N_3840,N_3387);
and U8699 (N_8699,N_4339,N_3893);
and U8700 (N_8700,N_49,N_2020);
and U8701 (N_8701,N_2002,N_746);
or U8702 (N_8702,N_785,N_1698);
nor U8703 (N_8703,N_1100,N_4162);
and U8704 (N_8704,N_3948,N_977);
or U8705 (N_8705,N_999,N_4637);
or U8706 (N_8706,N_906,N_946);
and U8707 (N_8707,N_4328,N_1911);
nor U8708 (N_8708,N_2713,N_4438);
nand U8709 (N_8709,N_3074,N_2639);
and U8710 (N_8710,N_1353,N_2915);
or U8711 (N_8711,N_2573,N_2925);
nor U8712 (N_8712,N_3320,N_2761);
or U8713 (N_8713,N_2708,N_3741);
nor U8714 (N_8714,N_4452,N_2955);
nand U8715 (N_8715,N_2032,N_3009);
nand U8716 (N_8716,N_4228,N_3833);
or U8717 (N_8717,N_3820,N_3770);
nor U8718 (N_8718,N_3506,N_2740);
nand U8719 (N_8719,N_2294,N_2982);
and U8720 (N_8720,N_3883,N_976);
or U8721 (N_8721,N_3412,N_4195);
nor U8722 (N_8722,N_4423,N_3759);
and U8723 (N_8723,N_4159,N_3986);
and U8724 (N_8724,N_836,N_1077);
nand U8725 (N_8725,N_265,N_4347);
nand U8726 (N_8726,N_2349,N_1835);
nand U8727 (N_8727,N_2992,N_1662);
nor U8728 (N_8728,N_4974,N_538);
nand U8729 (N_8729,N_4003,N_3623);
nand U8730 (N_8730,N_3585,N_2388);
or U8731 (N_8731,N_3939,N_1119);
nand U8732 (N_8732,N_2542,N_2465);
nor U8733 (N_8733,N_4649,N_359);
nand U8734 (N_8734,N_1012,N_3953);
and U8735 (N_8735,N_2974,N_98);
nor U8736 (N_8736,N_642,N_4961);
nand U8737 (N_8737,N_4733,N_427);
nand U8738 (N_8738,N_2626,N_3157);
nand U8739 (N_8739,N_1991,N_280);
or U8740 (N_8740,N_2835,N_4526);
and U8741 (N_8741,N_3531,N_2755);
nand U8742 (N_8742,N_1010,N_2272);
and U8743 (N_8743,N_4434,N_166);
nand U8744 (N_8744,N_2465,N_3756);
nor U8745 (N_8745,N_4957,N_4665);
or U8746 (N_8746,N_2200,N_4499);
nor U8747 (N_8747,N_1418,N_588);
or U8748 (N_8748,N_4629,N_4653);
or U8749 (N_8749,N_2947,N_1967);
nand U8750 (N_8750,N_48,N_4487);
and U8751 (N_8751,N_1052,N_4802);
nand U8752 (N_8752,N_3967,N_1184);
nand U8753 (N_8753,N_4780,N_4760);
or U8754 (N_8754,N_2396,N_2658);
or U8755 (N_8755,N_739,N_4252);
nand U8756 (N_8756,N_1635,N_2256);
nor U8757 (N_8757,N_4365,N_3316);
and U8758 (N_8758,N_3841,N_3128);
xnor U8759 (N_8759,N_3881,N_3690);
nand U8760 (N_8760,N_2140,N_104);
nand U8761 (N_8761,N_1931,N_1230);
nand U8762 (N_8762,N_1580,N_2979);
nor U8763 (N_8763,N_2032,N_3800);
or U8764 (N_8764,N_1587,N_1664);
nor U8765 (N_8765,N_452,N_1427);
nand U8766 (N_8766,N_2220,N_4489);
or U8767 (N_8767,N_2386,N_2889);
or U8768 (N_8768,N_4435,N_29);
nand U8769 (N_8769,N_1310,N_2299);
nand U8770 (N_8770,N_2797,N_3920);
nand U8771 (N_8771,N_25,N_4327);
and U8772 (N_8772,N_1775,N_2705);
and U8773 (N_8773,N_3905,N_2443);
nor U8774 (N_8774,N_1215,N_466);
nor U8775 (N_8775,N_3915,N_3333);
or U8776 (N_8776,N_3638,N_3032);
or U8777 (N_8777,N_4394,N_3618);
and U8778 (N_8778,N_2900,N_892);
nand U8779 (N_8779,N_1273,N_3343);
nand U8780 (N_8780,N_4267,N_1131);
or U8781 (N_8781,N_3818,N_4869);
nand U8782 (N_8782,N_3852,N_883);
nand U8783 (N_8783,N_2457,N_4830);
nor U8784 (N_8784,N_3696,N_1183);
or U8785 (N_8785,N_3101,N_3124);
nand U8786 (N_8786,N_2784,N_2396);
or U8787 (N_8787,N_4129,N_2438);
nor U8788 (N_8788,N_1970,N_1734);
or U8789 (N_8789,N_3957,N_4174);
nand U8790 (N_8790,N_2463,N_4867);
and U8791 (N_8791,N_2278,N_901);
nor U8792 (N_8792,N_3172,N_2452);
nand U8793 (N_8793,N_1853,N_3206);
and U8794 (N_8794,N_4200,N_3293);
nor U8795 (N_8795,N_4034,N_2661);
nand U8796 (N_8796,N_856,N_1720);
or U8797 (N_8797,N_4556,N_2717);
nand U8798 (N_8798,N_2868,N_2166);
nand U8799 (N_8799,N_542,N_4772);
nand U8800 (N_8800,N_905,N_2256);
nor U8801 (N_8801,N_4644,N_4208);
or U8802 (N_8802,N_1865,N_3716);
nand U8803 (N_8803,N_2298,N_3819);
xnor U8804 (N_8804,N_2151,N_1476);
and U8805 (N_8805,N_2156,N_2651);
and U8806 (N_8806,N_4308,N_4387);
or U8807 (N_8807,N_4032,N_38);
nand U8808 (N_8808,N_4724,N_1716);
or U8809 (N_8809,N_4765,N_2243);
or U8810 (N_8810,N_3690,N_3407);
xnor U8811 (N_8811,N_2647,N_1426);
and U8812 (N_8812,N_3859,N_1028);
nor U8813 (N_8813,N_4925,N_3322);
and U8814 (N_8814,N_2246,N_4177);
nor U8815 (N_8815,N_2300,N_2180);
or U8816 (N_8816,N_2782,N_3478);
and U8817 (N_8817,N_4288,N_114);
xor U8818 (N_8818,N_4654,N_106);
and U8819 (N_8819,N_4118,N_4320);
and U8820 (N_8820,N_268,N_3210);
and U8821 (N_8821,N_1208,N_1674);
nor U8822 (N_8822,N_1712,N_4420);
and U8823 (N_8823,N_4723,N_1615);
and U8824 (N_8824,N_2727,N_1362);
nand U8825 (N_8825,N_4863,N_4103);
nand U8826 (N_8826,N_2217,N_1829);
nand U8827 (N_8827,N_4865,N_3517);
nand U8828 (N_8828,N_1469,N_2415);
xnor U8829 (N_8829,N_4858,N_1126);
or U8830 (N_8830,N_767,N_2625);
nand U8831 (N_8831,N_1602,N_2556);
or U8832 (N_8832,N_3323,N_1946);
or U8833 (N_8833,N_1531,N_1163);
nor U8834 (N_8834,N_1612,N_4023);
nor U8835 (N_8835,N_2829,N_838);
or U8836 (N_8836,N_3019,N_2072);
nor U8837 (N_8837,N_3074,N_2631);
and U8838 (N_8838,N_1134,N_145);
and U8839 (N_8839,N_1304,N_4769);
or U8840 (N_8840,N_4241,N_4611);
nand U8841 (N_8841,N_2685,N_2827);
nor U8842 (N_8842,N_1728,N_3428);
and U8843 (N_8843,N_2396,N_4688);
and U8844 (N_8844,N_1278,N_1164);
and U8845 (N_8845,N_3591,N_3556);
nor U8846 (N_8846,N_2506,N_3668);
nand U8847 (N_8847,N_451,N_3536);
and U8848 (N_8848,N_3812,N_4688);
nand U8849 (N_8849,N_4130,N_4816);
nand U8850 (N_8850,N_1367,N_3842);
or U8851 (N_8851,N_1971,N_4812);
nand U8852 (N_8852,N_2135,N_4915);
nand U8853 (N_8853,N_1592,N_1078);
or U8854 (N_8854,N_171,N_1222);
nor U8855 (N_8855,N_2360,N_4277);
and U8856 (N_8856,N_1739,N_4348);
nand U8857 (N_8857,N_1688,N_1169);
and U8858 (N_8858,N_3489,N_3751);
or U8859 (N_8859,N_972,N_1580);
nand U8860 (N_8860,N_4962,N_3038);
nand U8861 (N_8861,N_602,N_3707);
nand U8862 (N_8862,N_3353,N_3792);
nor U8863 (N_8863,N_3561,N_4642);
nor U8864 (N_8864,N_1932,N_4402);
or U8865 (N_8865,N_3724,N_1113);
or U8866 (N_8866,N_714,N_4770);
and U8867 (N_8867,N_4956,N_566);
and U8868 (N_8868,N_2698,N_4880);
and U8869 (N_8869,N_2366,N_811);
or U8870 (N_8870,N_1647,N_2924);
and U8871 (N_8871,N_3981,N_3002);
or U8872 (N_8872,N_3608,N_936);
and U8873 (N_8873,N_2143,N_46);
and U8874 (N_8874,N_4056,N_2199);
or U8875 (N_8875,N_4597,N_4084);
or U8876 (N_8876,N_3994,N_111);
nor U8877 (N_8877,N_1900,N_1073);
and U8878 (N_8878,N_4605,N_1240);
or U8879 (N_8879,N_4559,N_2811);
and U8880 (N_8880,N_4636,N_4793);
or U8881 (N_8881,N_2573,N_2052);
and U8882 (N_8882,N_1441,N_3139);
or U8883 (N_8883,N_3379,N_3753);
and U8884 (N_8884,N_1214,N_1892);
and U8885 (N_8885,N_4888,N_3021);
nor U8886 (N_8886,N_1415,N_2174);
nor U8887 (N_8887,N_4928,N_3966);
nand U8888 (N_8888,N_1507,N_3431);
nor U8889 (N_8889,N_9,N_3371);
or U8890 (N_8890,N_2255,N_3621);
nand U8891 (N_8891,N_2101,N_1103);
and U8892 (N_8892,N_2488,N_3765);
and U8893 (N_8893,N_4737,N_2645);
nor U8894 (N_8894,N_4730,N_3183);
nand U8895 (N_8895,N_2727,N_379);
and U8896 (N_8896,N_983,N_1242);
and U8897 (N_8897,N_4299,N_553);
nand U8898 (N_8898,N_3885,N_1786);
nor U8899 (N_8899,N_1904,N_4449);
or U8900 (N_8900,N_3517,N_1081);
and U8901 (N_8901,N_1848,N_3108);
nor U8902 (N_8902,N_3645,N_2867);
and U8903 (N_8903,N_1123,N_369);
and U8904 (N_8904,N_1096,N_3345);
and U8905 (N_8905,N_3656,N_1938);
and U8906 (N_8906,N_1908,N_4714);
and U8907 (N_8907,N_4245,N_1327);
or U8908 (N_8908,N_3695,N_443);
xor U8909 (N_8909,N_2307,N_1618);
or U8910 (N_8910,N_1794,N_921);
or U8911 (N_8911,N_1121,N_4243);
and U8912 (N_8912,N_2772,N_4307);
nor U8913 (N_8913,N_2015,N_2008);
and U8914 (N_8914,N_4406,N_371);
nor U8915 (N_8915,N_1943,N_1547);
and U8916 (N_8916,N_31,N_3360);
or U8917 (N_8917,N_4296,N_3910);
and U8918 (N_8918,N_2608,N_2331);
nand U8919 (N_8919,N_1108,N_2195);
nand U8920 (N_8920,N_3376,N_2456);
xor U8921 (N_8921,N_169,N_406);
or U8922 (N_8922,N_2309,N_82);
nand U8923 (N_8923,N_2009,N_4482);
nand U8924 (N_8924,N_1260,N_2800);
and U8925 (N_8925,N_1852,N_558);
nand U8926 (N_8926,N_260,N_1466);
nand U8927 (N_8927,N_1222,N_1704);
nor U8928 (N_8928,N_3201,N_203);
or U8929 (N_8929,N_500,N_3493);
or U8930 (N_8930,N_351,N_3853);
or U8931 (N_8931,N_3391,N_1041);
and U8932 (N_8932,N_884,N_4746);
nand U8933 (N_8933,N_4703,N_3444);
nand U8934 (N_8934,N_3002,N_80);
nor U8935 (N_8935,N_2333,N_3695);
or U8936 (N_8936,N_4085,N_640);
nor U8937 (N_8937,N_4103,N_3008);
nand U8938 (N_8938,N_2360,N_4506);
or U8939 (N_8939,N_2578,N_3200);
nor U8940 (N_8940,N_535,N_1025);
or U8941 (N_8941,N_3570,N_1010);
nor U8942 (N_8942,N_1779,N_1265);
or U8943 (N_8943,N_404,N_3726);
or U8944 (N_8944,N_2468,N_1565);
nand U8945 (N_8945,N_3167,N_2188);
nor U8946 (N_8946,N_1789,N_2710);
nor U8947 (N_8947,N_1185,N_4558);
nor U8948 (N_8948,N_3269,N_2760);
or U8949 (N_8949,N_2109,N_1900);
or U8950 (N_8950,N_4949,N_4197);
and U8951 (N_8951,N_3711,N_689);
nor U8952 (N_8952,N_1300,N_1412);
nor U8953 (N_8953,N_4363,N_760);
nor U8954 (N_8954,N_4215,N_4648);
or U8955 (N_8955,N_2334,N_4227);
nor U8956 (N_8956,N_1654,N_1233);
and U8957 (N_8957,N_393,N_4345);
nand U8958 (N_8958,N_1148,N_790);
or U8959 (N_8959,N_3521,N_3714);
and U8960 (N_8960,N_3673,N_3526);
nand U8961 (N_8961,N_22,N_1078);
nand U8962 (N_8962,N_1102,N_1996);
nor U8963 (N_8963,N_3369,N_3952);
or U8964 (N_8964,N_2723,N_2219);
nand U8965 (N_8965,N_691,N_2073);
nor U8966 (N_8966,N_1977,N_3125);
or U8967 (N_8967,N_887,N_3956);
nand U8968 (N_8968,N_4213,N_827);
nand U8969 (N_8969,N_3115,N_2483);
or U8970 (N_8970,N_3634,N_2674);
or U8971 (N_8971,N_1432,N_66);
nand U8972 (N_8972,N_3257,N_4098);
nand U8973 (N_8973,N_103,N_159);
nor U8974 (N_8974,N_3955,N_2257);
and U8975 (N_8975,N_3724,N_3079);
nor U8976 (N_8976,N_1266,N_2579);
or U8977 (N_8977,N_3392,N_1757);
and U8978 (N_8978,N_4916,N_4242);
xor U8979 (N_8979,N_4291,N_3947);
or U8980 (N_8980,N_90,N_667);
nor U8981 (N_8981,N_1761,N_3233);
nor U8982 (N_8982,N_2190,N_1439);
nand U8983 (N_8983,N_4386,N_90);
nor U8984 (N_8984,N_1328,N_2431);
nand U8985 (N_8985,N_875,N_1390);
and U8986 (N_8986,N_4807,N_3774);
nor U8987 (N_8987,N_3220,N_1303);
nand U8988 (N_8988,N_3819,N_1686);
and U8989 (N_8989,N_4357,N_3633);
nand U8990 (N_8990,N_3831,N_3602);
or U8991 (N_8991,N_376,N_2626);
nand U8992 (N_8992,N_1841,N_1211);
nor U8993 (N_8993,N_449,N_4848);
nand U8994 (N_8994,N_4245,N_242);
and U8995 (N_8995,N_1735,N_2779);
or U8996 (N_8996,N_295,N_1630);
or U8997 (N_8997,N_4214,N_1941);
nand U8998 (N_8998,N_3273,N_3134);
and U8999 (N_8999,N_1690,N_2690);
nor U9000 (N_9000,N_273,N_3324);
nor U9001 (N_9001,N_1810,N_3077);
and U9002 (N_9002,N_2006,N_1818);
nor U9003 (N_9003,N_1297,N_1780);
and U9004 (N_9004,N_2927,N_4599);
nor U9005 (N_9005,N_403,N_4262);
nand U9006 (N_9006,N_671,N_493);
or U9007 (N_9007,N_3989,N_756);
or U9008 (N_9008,N_4600,N_3705);
and U9009 (N_9009,N_4353,N_709);
nand U9010 (N_9010,N_1024,N_4258);
nand U9011 (N_9011,N_674,N_3551);
and U9012 (N_9012,N_3093,N_4494);
and U9013 (N_9013,N_2648,N_2286);
nand U9014 (N_9014,N_1283,N_2527);
or U9015 (N_9015,N_1491,N_3970);
or U9016 (N_9016,N_3235,N_3860);
or U9017 (N_9017,N_4132,N_173);
or U9018 (N_9018,N_2677,N_1530);
or U9019 (N_9019,N_646,N_3428);
nand U9020 (N_9020,N_1518,N_975);
and U9021 (N_9021,N_4534,N_4424);
and U9022 (N_9022,N_1731,N_2697);
or U9023 (N_9023,N_2250,N_3776);
nor U9024 (N_9024,N_4543,N_4336);
or U9025 (N_9025,N_1449,N_2322);
nand U9026 (N_9026,N_4110,N_2159);
or U9027 (N_9027,N_600,N_495);
nand U9028 (N_9028,N_2581,N_2173);
or U9029 (N_9029,N_2146,N_1862);
nand U9030 (N_9030,N_1525,N_2550);
and U9031 (N_9031,N_2878,N_600);
and U9032 (N_9032,N_4193,N_1189);
or U9033 (N_9033,N_4095,N_592);
or U9034 (N_9034,N_3327,N_3276);
and U9035 (N_9035,N_287,N_3833);
nand U9036 (N_9036,N_4089,N_703);
nand U9037 (N_9037,N_1387,N_1563);
nor U9038 (N_9038,N_3599,N_3167);
and U9039 (N_9039,N_1139,N_2178);
and U9040 (N_9040,N_868,N_3057);
and U9041 (N_9041,N_1996,N_4760);
nor U9042 (N_9042,N_4996,N_4109);
or U9043 (N_9043,N_3931,N_1385);
nor U9044 (N_9044,N_1264,N_1133);
nor U9045 (N_9045,N_3874,N_2339);
or U9046 (N_9046,N_226,N_4033);
nand U9047 (N_9047,N_4161,N_429);
or U9048 (N_9048,N_4034,N_2079);
nand U9049 (N_9049,N_2615,N_2504);
nand U9050 (N_9050,N_1080,N_2062);
and U9051 (N_9051,N_1397,N_3819);
or U9052 (N_9052,N_891,N_1434);
and U9053 (N_9053,N_2136,N_216);
and U9054 (N_9054,N_4136,N_3342);
xor U9055 (N_9055,N_466,N_2758);
nor U9056 (N_9056,N_37,N_2918);
nor U9057 (N_9057,N_3467,N_1892);
nand U9058 (N_9058,N_3060,N_4638);
or U9059 (N_9059,N_4728,N_4599);
nand U9060 (N_9060,N_234,N_1921);
nand U9061 (N_9061,N_3135,N_2273);
nand U9062 (N_9062,N_414,N_4518);
nand U9063 (N_9063,N_1259,N_3108);
nand U9064 (N_9064,N_3645,N_39);
or U9065 (N_9065,N_912,N_802);
and U9066 (N_9066,N_2209,N_3462);
or U9067 (N_9067,N_4696,N_3447);
or U9068 (N_9068,N_699,N_4298);
xnor U9069 (N_9069,N_919,N_4457);
xnor U9070 (N_9070,N_1185,N_718);
nand U9071 (N_9071,N_1064,N_1665);
nor U9072 (N_9072,N_800,N_4279);
nand U9073 (N_9073,N_3905,N_15);
or U9074 (N_9074,N_4754,N_3527);
nor U9075 (N_9075,N_1561,N_788);
nor U9076 (N_9076,N_1652,N_1247);
and U9077 (N_9077,N_3196,N_3812);
nand U9078 (N_9078,N_3185,N_613);
nand U9079 (N_9079,N_4048,N_4466);
and U9080 (N_9080,N_3489,N_202);
or U9081 (N_9081,N_642,N_4279);
nand U9082 (N_9082,N_4865,N_4986);
and U9083 (N_9083,N_4048,N_4515);
nand U9084 (N_9084,N_1077,N_4141);
or U9085 (N_9085,N_1719,N_3461);
or U9086 (N_9086,N_4384,N_4479);
nand U9087 (N_9087,N_4879,N_3237);
and U9088 (N_9088,N_3680,N_4845);
nor U9089 (N_9089,N_2414,N_985);
nand U9090 (N_9090,N_2526,N_4606);
or U9091 (N_9091,N_1974,N_4106);
and U9092 (N_9092,N_879,N_1452);
or U9093 (N_9093,N_1684,N_4643);
xor U9094 (N_9094,N_1799,N_112);
nand U9095 (N_9095,N_2463,N_4510);
and U9096 (N_9096,N_345,N_1780);
and U9097 (N_9097,N_4463,N_1713);
and U9098 (N_9098,N_3423,N_4857);
or U9099 (N_9099,N_4824,N_4694);
nand U9100 (N_9100,N_1973,N_2224);
and U9101 (N_9101,N_1985,N_3859);
nor U9102 (N_9102,N_1590,N_2631);
nor U9103 (N_9103,N_1832,N_3704);
or U9104 (N_9104,N_921,N_1461);
nand U9105 (N_9105,N_4792,N_326);
nand U9106 (N_9106,N_3173,N_689);
or U9107 (N_9107,N_1186,N_1107);
or U9108 (N_9108,N_990,N_3994);
or U9109 (N_9109,N_1237,N_3590);
or U9110 (N_9110,N_4875,N_4686);
and U9111 (N_9111,N_1708,N_4923);
nand U9112 (N_9112,N_4735,N_1619);
or U9113 (N_9113,N_3268,N_4550);
nor U9114 (N_9114,N_1795,N_3314);
nand U9115 (N_9115,N_1311,N_3836);
nand U9116 (N_9116,N_628,N_4765);
or U9117 (N_9117,N_31,N_497);
nand U9118 (N_9118,N_1265,N_3285);
nor U9119 (N_9119,N_1376,N_4578);
or U9120 (N_9120,N_949,N_1427);
nor U9121 (N_9121,N_1924,N_2047);
or U9122 (N_9122,N_508,N_4921);
nand U9123 (N_9123,N_193,N_1328);
nand U9124 (N_9124,N_1473,N_581);
nor U9125 (N_9125,N_3412,N_982);
and U9126 (N_9126,N_2693,N_2813);
and U9127 (N_9127,N_3968,N_4348);
or U9128 (N_9128,N_4593,N_3399);
nand U9129 (N_9129,N_542,N_651);
nor U9130 (N_9130,N_4049,N_2144);
xor U9131 (N_9131,N_2091,N_4807);
or U9132 (N_9132,N_813,N_2782);
and U9133 (N_9133,N_183,N_4113);
and U9134 (N_9134,N_4901,N_396);
nor U9135 (N_9135,N_2157,N_4341);
nand U9136 (N_9136,N_1385,N_4850);
nor U9137 (N_9137,N_1551,N_388);
nor U9138 (N_9138,N_3205,N_2055);
nand U9139 (N_9139,N_1268,N_4467);
nand U9140 (N_9140,N_4035,N_1072);
nand U9141 (N_9141,N_3547,N_1949);
and U9142 (N_9142,N_1514,N_4745);
nand U9143 (N_9143,N_2076,N_4733);
or U9144 (N_9144,N_1725,N_2537);
nand U9145 (N_9145,N_975,N_2894);
nand U9146 (N_9146,N_1557,N_3586);
nand U9147 (N_9147,N_4270,N_1739);
and U9148 (N_9148,N_2301,N_4437);
and U9149 (N_9149,N_1260,N_2209);
nand U9150 (N_9150,N_494,N_1115);
and U9151 (N_9151,N_2291,N_1398);
nor U9152 (N_9152,N_4689,N_1269);
and U9153 (N_9153,N_1550,N_3748);
and U9154 (N_9154,N_544,N_4340);
nand U9155 (N_9155,N_952,N_2386);
nand U9156 (N_9156,N_739,N_4064);
or U9157 (N_9157,N_4839,N_1896);
or U9158 (N_9158,N_4630,N_164);
nor U9159 (N_9159,N_2747,N_2005);
and U9160 (N_9160,N_2686,N_121);
and U9161 (N_9161,N_2796,N_2661);
or U9162 (N_9162,N_1983,N_786);
nor U9163 (N_9163,N_3603,N_3196);
nor U9164 (N_9164,N_3170,N_4627);
or U9165 (N_9165,N_4441,N_3133);
nand U9166 (N_9166,N_4603,N_2093);
and U9167 (N_9167,N_4465,N_385);
and U9168 (N_9168,N_3357,N_1166);
or U9169 (N_9169,N_3936,N_2);
or U9170 (N_9170,N_2381,N_423);
nand U9171 (N_9171,N_4945,N_3700);
or U9172 (N_9172,N_4414,N_4154);
and U9173 (N_9173,N_171,N_3008);
or U9174 (N_9174,N_2569,N_783);
nand U9175 (N_9175,N_2751,N_437);
or U9176 (N_9176,N_2484,N_2782);
nand U9177 (N_9177,N_132,N_3124);
and U9178 (N_9178,N_1738,N_862);
or U9179 (N_9179,N_795,N_907);
nand U9180 (N_9180,N_4267,N_718);
and U9181 (N_9181,N_1771,N_2017);
or U9182 (N_9182,N_1714,N_684);
or U9183 (N_9183,N_4605,N_318);
nand U9184 (N_9184,N_2643,N_3246);
and U9185 (N_9185,N_2372,N_836);
and U9186 (N_9186,N_2741,N_2081);
nor U9187 (N_9187,N_2200,N_652);
nor U9188 (N_9188,N_1224,N_3613);
and U9189 (N_9189,N_181,N_2079);
nor U9190 (N_9190,N_3666,N_1738);
xnor U9191 (N_9191,N_483,N_1651);
and U9192 (N_9192,N_2103,N_2442);
nor U9193 (N_9193,N_3539,N_4417);
and U9194 (N_9194,N_901,N_1903);
or U9195 (N_9195,N_740,N_2807);
and U9196 (N_9196,N_1597,N_81);
nand U9197 (N_9197,N_1337,N_4474);
nor U9198 (N_9198,N_2974,N_4606);
nor U9199 (N_9199,N_748,N_583);
xor U9200 (N_9200,N_698,N_3826);
and U9201 (N_9201,N_4226,N_3263);
and U9202 (N_9202,N_3446,N_3969);
and U9203 (N_9203,N_2876,N_451);
xor U9204 (N_9204,N_766,N_4237);
nand U9205 (N_9205,N_2174,N_3034);
nand U9206 (N_9206,N_2608,N_2368);
and U9207 (N_9207,N_695,N_3210);
nand U9208 (N_9208,N_4947,N_4386);
nor U9209 (N_9209,N_3349,N_2873);
nand U9210 (N_9210,N_6,N_4718);
nand U9211 (N_9211,N_1630,N_3892);
nand U9212 (N_9212,N_611,N_1997);
nand U9213 (N_9213,N_447,N_3849);
nand U9214 (N_9214,N_236,N_1596);
nand U9215 (N_9215,N_1553,N_2);
nand U9216 (N_9216,N_1670,N_1893);
nand U9217 (N_9217,N_4126,N_4180);
or U9218 (N_9218,N_4849,N_3299);
or U9219 (N_9219,N_358,N_3480);
or U9220 (N_9220,N_3142,N_835);
nor U9221 (N_9221,N_1611,N_3175);
nor U9222 (N_9222,N_2850,N_3319);
nand U9223 (N_9223,N_4393,N_4327);
nand U9224 (N_9224,N_2339,N_1053);
nand U9225 (N_9225,N_2492,N_1532);
and U9226 (N_9226,N_3697,N_2029);
or U9227 (N_9227,N_2847,N_2948);
nor U9228 (N_9228,N_4605,N_3476);
and U9229 (N_9229,N_312,N_1181);
or U9230 (N_9230,N_800,N_2418);
or U9231 (N_9231,N_481,N_1940);
and U9232 (N_9232,N_279,N_1610);
xnor U9233 (N_9233,N_1691,N_1249);
or U9234 (N_9234,N_1411,N_4236);
nor U9235 (N_9235,N_2136,N_837);
or U9236 (N_9236,N_1371,N_4351);
nand U9237 (N_9237,N_2941,N_2020);
and U9238 (N_9238,N_4580,N_4539);
and U9239 (N_9239,N_4328,N_3737);
nand U9240 (N_9240,N_361,N_3519);
and U9241 (N_9241,N_969,N_1804);
or U9242 (N_9242,N_1049,N_2312);
and U9243 (N_9243,N_936,N_1179);
nor U9244 (N_9244,N_1249,N_3088);
nand U9245 (N_9245,N_4866,N_1787);
nor U9246 (N_9246,N_1234,N_934);
xor U9247 (N_9247,N_3083,N_3542);
nor U9248 (N_9248,N_4643,N_4117);
or U9249 (N_9249,N_2034,N_4747);
nor U9250 (N_9250,N_3963,N_1921);
nand U9251 (N_9251,N_2978,N_887);
or U9252 (N_9252,N_330,N_1565);
and U9253 (N_9253,N_68,N_920);
nand U9254 (N_9254,N_3935,N_3860);
nand U9255 (N_9255,N_1441,N_470);
nor U9256 (N_9256,N_2538,N_4029);
and U9257 (N_9257,N_716,N_328);
or U9258 (N_9258,N_686,N_904);
or U9259 (N_9259,N_2956,N_3693);
or U9260 (N_9260,N_1679,N_4059);
and U9261 (N_9261,N_369,N_4295);
nand U9262 (N_9262,N_3949,N_2865);
nor U9263 (N_9263,N_2741,N_485);
or U9264 (N_9264,N_2674,N_2618);
and U9265 (N_9265,N_1109,N_1666);
and U9266 (N_9266,N_3409,N_1912);
and U9267 (N_9267,N_1537,N_3578);
and U9268 (N_9268,N_2832,N_4251);
nor U9269 (N_9269,N_2748,N_1316);
nor U9270 (N_9270,N_1171,N_1175);
nand U9271 (N_9271,N_2424,N_3023);
and U9272 (N_9272,N_2660,N_4753);
or U9273 (N_9273,N_1243,N_3748);
and U9274 (N_9274,N_2966,N_51);
or U9275 (N_9275,N_4370,N_3491);
or U9276 (N_9276,N_182,N_734);
nand U9277 (N_9277,N_1381,N_3368);
nor U9278 (N_9278,N_1397,N_2998);
nand U9279 (N_9279,N_135,N_2546);
nor U9280 (N_9280,N_4043,N_4153);
nor U9281 (N_9281,N_643,N_2089);
and U9282 (N_9282,N_1461,N_2550);
nor U9283 (N_9283,N_1398,N_55);
and U9284 (N_9284,N_1993,N_4676);
or U9285 (N_9285,N_1319,N_4157);
and U9286 (N_9286,N_2888,N_4327);
nand U9287 (N_9287,N_4413,N_2084);
and U9288 (N_9288,N_771,N_3135);
and U9289 (N_9289,N_3492,N_4155);
and U9290 (N_9290,N_1100,N_4173);
nand U9291 (N_9291,N_4306,N_2501);
and U9292 (N_9292,N_1575,N_207);
or U9293 (N_9293,N_121,N_427);
nor U9294 (N_9294,N_1074,N_466);
or U9295 (N_9295,N_3429,N_180);
nor U9296 (N_9296,N_1807,N_2229);
and U9297 (N_9297,N_2230,N_4405);
or U9298 (N_9298,N_60,N_4590);
or U9299 (N_9299,N_1428,N_4440);
nand U9300 (N_9300,N_54,N_4681);
nand U9301 (N_9301,N_3091,N_3008);
nand U9302 (N_9302,N_2783,N_3854);
or U9303 (N_9303,N_2581,N_3755);
or U9304 (N_9304,N_4500,N_1034);
and U9305 (N_9305,N_2129,N_2532);
nand U9306 (N_9306,N_1054,N_4900);
nor U9307 (N_9307,N_2612,N_4755);
or U9308 (N_9308,N_466,N_367);
nor U9309 (N_9309,N_2733,N_2182);
or U9310 (N_9310,N_148,N_3875);
nand U9311 (N_9311,N_4008,N_1967);
or U9312 (N_9312,N_4733,N_569);
nand U9313 (N_9313,N_2492,N_382);
and U9314 (N_9314,N_2339,N_51);
and U9315 (N_9315,N_2931,N_4784);
nand U9316 (N_9316,N_1032,N_2076);
or U9317 (N_9317,N_3773,N_2248);
and U9318 (N_9318,N_1122,N_3283);
nor U9319 (N_9319,N_2424,N_3838);
or U9320 (N_9320,N_3772,N_389);
nor U9321 (N_9321,N_4759,N_2754);
nor U9322 (N_9322,N_16,N_3563);
nor U9323 (N_9323,N_3842,N_4975);
or U9324 (N_9324,N_4089,N_3756);
nor U9325 (N_9325,N_156,N_4078);
nand U9326 (N_9326,N_959,N_4963);
and U9327 (N_9327,N_1221,N_4614);
and U9328 (N_9328,N_4488,N_2853);
or U9329 (N_9329,N_2798,N_4232);
or U9330 (N_9330,N_1245,N_341);
nand U9331 (N_9331,N_2090,N_1177);
and U9332 (N_9332,N_1397,N_3027);
or U9333 (N_9333,N_367,N_2341);
and U9334 (N_9334,N_538,N_3183);
nor U9335 (N_9335,N_3020,N_4673);
and U9336 (N_9336,N_1400,N_2359);
nand U9337 (N_9337,N_4946,N_1379);
nand U9338 (N_9338,N_639,N_3348);
xor U9339 (N_9339,N_3060,N_4164);
or U9340 (N_9340,N_2895,N_1639);
nand U9341 (N_9341,N_2250,N_3087);
and U9342 (N_9342,N_3407,N_2670);
and U9343 (N_9343,N_3520,N_110);
xnor U9344 (N_9344,N_3493,N_1032);
nor U9345 (N_9345,N_405,N_1507);
or U9346 (N_9346,N_937,N_1715);
nor U9347 (N_9347,N_3663,N_3719);
or U9348 (N_9348,N_3151,N_11);
nand U9349 (N_9349,N_330,N_1023);
nand U9350 (N_9350,N_1803,N_3591);
and U9351 (N_9351,N_4094,N_1662);
or U9352 (N_9352,N_3231,N_1501);
nand U9353 (N_9353,N_2722,N_3473);
nor U9354 (N_9354,N_549,N_2852);
nor U9355 (N_9355,N_4932,N_1492);
or U9356 (N_9356,N_2294,N_3051);
and U9357 (N_9357,N_1830,N_332);
or U9358 (N_9358,N_148,N_2001);
nand U9359 (N_9359,N_3536,N_253);
or U9360 (N_9360,N_4157,N_15);
nor U9361 (N_9361,N_4156,N_447);
and U9362 (N_9362,N_961,N_1750);
nand U9363 (N_9363,N_1014,N_1514);
and U9364 (N_9364,N_2599,N_2503);
or U9365 (N_9365,N_956,N_2431);
xnor U9366 (N_9366,N_4615,N_4286);
and U9367 (N_9367,N_3386,N_1551);
or U9368 (N_9368,N_1791,N_2326);
nor U9369 (N_9369,N_2203,N_1026);
or U9370 (N_9370,N_4458,N_2774);
or U9371 (N_9371,N_1473,N_1871);
nand U9372 (N_9372,N_4769,N_2340);
nor U9373 (N_9373,N_1751,N_3488);
nor U9374 (N_9374,N_3642,N_2022);
and U9375 (N_9375,N_1270,N_2879);
and U9376 (N_9376,N_4326,N_3227);
nor U9377 (N_9377,N_741,N_4248);
and U9378 (N_9378,N_2928,N_2514);
nand U9379 (N_9379,N_3717,N_2205);
nor U9380 (N_9380,N_3717,N_771);
nor U9381 (N_9381,N_2159,N_119);
nand U9382 (N_9382,N_550,N_4568);
nor U9383 (N_9383,N_1355,N_3997);
or U9384 (N_9384,N_431,N_3649);
nand U9385 (N_9385,N_3308,N_865);
nor U9386 (N_9386,N_4851,N_1049);
nor U9387 (N_9387,N_2731,N_4831);
or U9388 (N_9388,N_184,N_3865);
xor U9389 (N_9389,N_351,N_2098);
nor U9390 (N_9390,N_889,N_3778);
nand U9391 (N_9391,N_3188,N_578);
or U9392 (N_9392,N_3243,N_284);
and U9393 (N_9393,N_2372,N_655);
and U9394 (N_9394,N_1334,N_2759);
and U9395 (N_9395,N_3266,N_4208);
nor U9396 (N_9396,N_561,N_1036);
nand U9397 (N_9397,N_2973,N_2782);
and U9398 (N_9398,N_4543,N_3514);
or U9399 (N_9399,N_3518,N_675);
or U9400 (N_9400,N_4629,N_1570);
nor U9401 (N_9401,N_1918,N_2798);
nor U9402 (N_9402,N_4351,N_2274);
and U9403 (N_9403,N_1824,N_136);
or U9404 (N_9404,N_4633,N_841);
nor U9405 (N_9405,N_637,N_4161);
nand U9406 (N_9406,N_3452,N_2244);
and U9407 (N_9407,N_4748,N_2767);
or U9408 (N_9408,N_1317,N_2129);
nand U9409 (N_9409,N_226,N_1368);
nand U9410 (N_9410,N_4558,N_1830);
or U9411 (N_9411,N_3803,N_599);
and U9412 (N_9412,N_3584,N_2013);
nor U9413 (N_9413,N_1199,N_3542);
nand U9414 (N_9414,N_3821,N_38);
nor U9415 (N_9415,N_1299,N_2159);
nor U9416 (N_9416,N_4447,N_2275);
or U9417 (N_9417,N_1363,N_3532);
nand U9418 (N_9418,N_2797,N_2140);
nand U9419 (N_9419,N_2621,N_749);
nor U9420 (N_9420,N_1915,N_3790);
nor U9421 (N_9421,N_1960,N_4635);
or U9422 (N_9422,N_3512,N_101);
and U9423 (N_9423,N_1292,N_419);
nand U9424 (N_9424,N_3776,N_2453);
nor U9425 (N_9425,N_4732,N_1695);
and U9426 (N_9426,N_197,N_2279);
or U9427 (N_9427,N_4430,N_680);
nand U9428 (N_9428,N_152,N_941);
and U9429 (N_9429,N_1514,N_2131);
or U9430 (N_9430,N_2259,N_1221);
nand U9431 (N_9431,N_2329,N_215);
nor U9432 (N_9432,N_1130,N_1585);
or U9433 (N_9433,N_331,N_3448);
or U9434 (N_9434,N_1052,N_3180);
and U9435 (N_9435,N_801,N_3261);
nand U9436 (N_9436,N_4266,N_2556);
or U9437 (N_9437,N_4552,N_3542);
and U9438 (N_9438,N_3856,N_155);
or U9439 (N_9439,N_2293,N_4391);
nand U9440 (N_9440,N_2867,N_1026);
and U9441 (N_9441,N_255,N_2363);
and U9442 (N_9442,N_2906,N_1673);
and U9443 (N_9443,N_1044,N_3656);
and U9444 (N_9444,N_3020,N_4750);
nor U9445 (N_9445,N_2541,N_4591);
nor U9446 (N_9446,N_4800,N_2335);
and U9447 (N_9447,N_1604,N_3561);
or U9448 (N_9448,N_1331,N_4927);
and U9449 (N_9449,N_753,N_3875);
and U9450 (N_9450,N_2718,N_1344);
nand U9451 (N_9451,N_2078,N_796);
nand U9452 (N_9452,N_611,N_401);
or U9453 (N_9453,N_3678,N_2144);
or U9454 (N_9454,N_2411,N_3964);
nand U9455 (N_9455,N_1710,N_2217);
or U9456 (N_9456,N_3212,N_3611);
or U9457 (N_9457,N_452,N_663);
nand U9458 (N_9458,N_2074,N_1085);
and U9459 (N_9459,N_4547,N_1676);
nand U9460 (N_9460,N_2002,N_3627);
nor U9461 (N_9461,N_2194,N_318);
nor U9462 (N_9462,N_524,N_4401);
xnor U9463 (N_9463,N_3612,N_1155);
and U9464 (N_9464,N_3174,N_4873);
and U9465 (N_9465,N_3382,N_1029);
nand U9466 (N_9466,N_3616,N_3491);
or U9467 (N_9467,N_3741,N_4741);
or U9468 (N_9468,N_1539,N_4371);
nand U9469 (N_9469,N_459,N_3501);
or U9470 (N_9470,N_2373,N_698);
nand U9471 (N_9471,N_893,N_3746);
nor U9472 (N_9472,N_448,N_4831);
nand U9473 (N_9473,N_565,N_856);
and U9474 (N_9474,N_2880,N_363);
nor U9475 (N_9475,N_3551,N_3259);
nand U9476 (N_9476,N_2069,N_478);
and U9477 (N_9477,N_4563,N_521);
nor U9478 (N_9478,N_3978,N_4540);
or U9479 (N_9479,N_3876,N_63);
nand U9480 (N_9480,N_2552,N_4517);
or U9481 (N_9481,N_4989,N_2994);
and U9482 (N_9482,N_704,N_3272);
and U9483 (N_9483,N_197,N_116);
or U9484 (N_9484,N_3596,N_3546);
and U9485 (N_9485,N_1031,N_1386);
nand U9486 (N_9486,N_4822,N_2821);
nor U9487 (N_9487,N_2697,N_339);
or U9488 (N_9488,N_103,N_374);
or U9489 (N_9489,N_2075,N_3315);
or U9490 (N_9490,N_4616,N_1995);
nand U9491 (N_9491,N_1103,N_857);
or U9492 (N_9492,N_1272,N_1444);
nor U9493 (N_9493,N_3476,N_1346);
and U9494 (N_9494,N_2053,N_1804);
or U9495 (N_9495,N_437,N_3105);
or U9496 (N_9496,N_4232,N_1795);
or U9497 (N_9497,N_4079,N_1861);
and U9498 (N_9498,N_3372,N_4783);
or U9499 (N_9499,N_3134,N_3672);
and U9500 (N_9500,N_3746,N_1818);
nand U9501 (N_9501,N_682,N_471);
nand U9502 (N_9502,N_3274,N_396);
and U9503 (N_9503,N_3526,N_1817);
xor U9504 (N_9504,N_417,N_2465);
and U9505 (N_9505,N_3017,N_1788);
and U9506 (N_9506,N_3168,N_1145);
nand U9507 (N_9507,N_2561,N_1992);
or U9508 (N_9508,N_2415,N_770);
or U9509 (N_9509,N_3269,N_2732);
xnor U9510 (N_9510,N_797,N_443);
or U9511 (N_9511,N_578,N_524);
nor U9512 (N_9512,N_3062,N_2025);
nand U9513 (N_9513,N_1766,N_2568);
nor U9514 (N_9514,N_4389,N_615);
and U9515 (N_9515,N_148,N_1893);
nor U9516 (N_9516,N_1729,N_2583);
nor U9517 (N_9517,N_808,N_2928);
nor U9518 (N_9518,N_368,N_3396);
or U9519 (N_9519,N_4983,N_2732);
or U9520 (N_9520,N_3106,N_3799);
nand U9521 (N_9521,N_2322,N_471);
or U9522 (N_9522,N_2537,N_1129);
nand U9523 (N_9523,N_1580,N_4053);
or U9524 (N_9524,N_1964,N_3244);
nand U9525 (N_9525,N_1874,N_1519);
and U9526 (N_9526,N_4358,N_2990);
nand U9527 (N_9527,N_3601,N_4023);
or U9528 (N_9528,N_119,N_1554);
nor U9529 (N_9529,N_3109,N_1849);
xor U9530 (N_9530,N_4662,N_3746);
nand U9531 (N_9531,N_3019,N_4273);
nor U9532 (N_9532,N_3054,N_2333);
nor U9533 (N_9533,N_2026,N_1593);
or U9534 (N_9534,N_1287,N_3680);
nor U9535 (N_9535,N_1282,N_3848);
nor U9536 (N_9536,N_2333,N_4263);
nand U9537 (N_9537,N_1692,N_2394);
and U9538 (N_9538,N_3919,N_4380);
nand U9539 (N_9539,N_2831,N_4404);
nor U9540 (N_9540,N_2334,N_4289);
nor U9541 (N_9541,N_4293,N_4219);
or U9542 (N_9542,N_485,N_4532);
nor U9543 (N_9543,N_4005,N_396);
nand U9544 (N_9544,N_4416,N_2515);
or U9545 (N_9545,N_4842,N_3640);
nor U9546 (N_9546,N_3582,N_85);
and U9547 (N_9547,N_1591,N_3135);
or U9548 (N_9548,N_3880,N_3787);
nor U9549 (N_9549,N_3998,N_2984);
and U9550 (N_9550,N_2772,N_4686);
nand U9551 (N_9551,N_4848,N_2191);
nand U9552 (N_9552,N_3307,N_3312);
nand U9553 (N_9553,N_3010,N_1852);
and U9554 (N_9554,N_2677,N_4843);
nand U9555 (N_9555,N_2811,N_2054);
nand U9556 (N_9556,N_2549,N_2324);
and U9557 (N_9557,N_2054,N_1183);
nand U9558 (N_9558,N_1404,N_4231);
xnor U9559 (N_9559,N_1785,N_2973);
nand U9560 (N_9560,N_4115,N_3709);
nor U9561 (N_9561,N_1084,N_3489);
or U9562 (N_9562,N_1008,N_4413);
nor U9563 (N_9563,N_419,N_131);
nand U9564 (N_9564,N_3890,N_1780);
and U9565 (N_9565,N_3504,N_1023);
nand U9566 (N_9566,N_1947,N_444);
nand U9567 (N_9567,N_3205,N_2089);
nand U9568 (N_9568,N_2181,N_3474);
or U9569 (N_9569,N_4681,N_360);
nor U9570 (N_9570,N_4067,N_1144);
or U9571 (N_9571,N_4388,N_788);
or U9572 (N_9572,N_4513,N_3537);
and U9573 (N_9573,N_209,N_1050);
or U9574 (N_9574,N_3894,N_1743);
and U9575 (N_9575,N_3981,N_769);
nand U9576 (N_9576,N_4805,N_291);
nor U9577 (N_9577,N_2267,N_1342);
nand U9578 (N_9578,N_4596,N_2383);
nor U9579 (N_9579,N_1921,N_908);
or U9580 (N_9580,N_1253,N_1601);
and U9581 (N_9581,N_725,N_2916);
nand U9582 (N_9582,N_300,N_2363);
and U9583 (N_9583,N_3043,N_4630);
nand U9584 (N_9584,N_4249,N_83);
nor U9585 (N_9585,N_2379,N_3387);
nand U9586 (N_9586,N_3118,N_4850);
or U9587 (N_9587,N_4371,N_242);
xnor U9588 (N_9588,N_1047,N_4998);
and U9589 (N_9589,N_4799,N_2455);
or U9590 (N_9590,N_2590,N_1071);
nor U9591 (N_9591,N_4202,N_986);
nor U9592 (N_9592,N_161,N_1268);
nand U9593 (N_9593,N_4305,N_2031);
or U9594 (N_9594,N_989,N_425);
nand U9595 (N_9595,N_687,N_1028);
or U9596 (N_9596,N_1908,N_4559);
or U9597 (N_9597,N_2905,N_780);
nand U9598 (N_9598,N_3468,N_2390);
nor U9599 (N_9599,N_3775,N_2855);
nand U9600 (N_9600,N_1680,N_1900);
nand U9601 (N_9601,N_4057,N_1298);
nand U9602 (N_9602,N_3304,N_1881);
nand U9603 (N_9603,N_3428,N_3223);
nand U9604 (N_9604,N_2099,N_2474);
and U9605 (N_9605,N_2315,N_1797);
or U9606 (N_9606,N_4202,N_1938);
nor U9607 (N_9607,N_4552,N_3557);
or U9608 (N_9608,N_2859,N_1191);
nand U9609 (N_9609,N_3811,N_1072);
and U9610 (N_9610,N_1103,N_4765);
nand U9611 (N_9611,N_3557,N_1652);
and U9612 (N_9612,N_1906,N_3208);
and U9613 (N_9613,N_2318,N_4996);
nor U9614 (N_9614,N_3532,N_1761);
or U9615 (N_9615,N_926,N_234);
or U9616 (N_9616,N_4904,N_1711);
nand U9617 (N_9617,N_2273,N_3583);
nor U9618 (N_9618,N_1199,N_3934);
nor U9619 (N_9619,N_3055,N_3327);
nor U9620 (N_9620,N_4578,N_1720);
nand U9621 (N_9621,N_3560,N_4648);
and U9622 (N_9622,N_1501,N_2000);
nor U9623 (N_9623,N_4768,N_1393);
nand U9624 (N_9624,N_2296,N_1642);
nand U9625 (N_9625,N_1246,N_3250);
or U9626 (N_9626,N_461,N_1260);
and U9627 (N_9627,N_4961,N_2713);
nand U9628 (N_9628,N_2903,N_3047);
or U9629 (N_9629,N_3352,N_3304);
or U9630 (N_9630,N_1564,N_4664);
xnor U9631 (N_9631,N_4354,N_3396);
or U9632 (N_9632,N_3788,N_3637);
and U9633 (N_9633,N_1447,N_3628);
nor U9634 (N_9634,N_3667,N_4330);
nand U9635 (N_9635,N_4119,N_899);
and U9636 (N_9636,N_4527,N_1555);
or U9637 (N_9637,N_2742,N_2515);
and U9638 (N_9638,N_1583,N_4871);
nand U9639 (N_9639,N_554,N_3412);
nor U9640 (N_9640,N_4818,N_2187);
nor U9641 (N_9641,N_2021,N_3150);
nand U9642 (N_9642,N_1916,N_2105);
nor U9643 (N_9643,N_2636,N_2470);
and U9644 (N_9644,N_4761,N_969);
and U9645 (N_9645,N_1050,N_608);
nand U9646 (N_9646,N_1862,N_2453);
nand U9647 (N_9647,N_797,N_2714);
and U9648 (N_9648,N_1795,N_4149);
and U9649 (N_9649,N_4023,N_733);
nand U9650 (N_9650,N_2380,N_1887);
and U9651 (N_9651,N_2159,N_793);
or U9652 (N_9652,N_860,N_3036);
nor U9653 (N_9653,N_1450,N_1713);
nand U9654 (N_9654,N_4322,N_4302);
nor U9655 (N_9655,N_1405,N_660);
and U9656 (N_9656,N_787,N_1561);
nand U9657 (N_9657,N_3878,N_4829);
and U9658 (N_9658,N_2049,N_906);
nand U9659 (N_9659,N_1315,N_3628);
or U9660 (N_9660,N_4087,N_3746);
or U9661 (N_9661,N_3681,N_601);
nor U9662 (N_9662,N_4380,N_2058);
nor U9663 (N_9663,N_552,N_3737);
nor U9664 (N_9664,N_3382,N_4927);
or U9665 (N_9665,N_623,N_362);
or U9666 (N_9666,N_4352,N_100);
or U9667 (N_9667,N_1250,N_107);
nor U9668 (N_9668,N_3138,N_2520);
nand U9669 (N_9669,N_2229,N_2121);
nand U9670 (N_9670,N_2424,N_483);
or U9671 (N_9671,N_802,N_3407);
nor U9672 (N_9672,N_1063,N_3320);
and U9673 (N_9673,N_4377,N_4564);
or U9674 (N_9674,N_3237,N_3756);
nor U9675 (N_9675,N_2450,N_3913);
nor U9676 (N_9676,N_2563,N_359);
nand U9677 (N_9677,N_2724,N_3063);
nor U9678 (N_9678,N_2979,N_3593);
nor U9679 (N_9679,N_4824,N_3863);
or U9680 (N_9680,N_1935,N_2779);
nand U9681 (N_9681,N_3057,N_148);
nand U9682 (N_9682,N_1222,N_2233);
and U9683 (N_9683,N_4835,N_1423);
nand U9684 (N_9684,N_1576,N_1314);
nand U9685 (N_9685,N_1603,N_4306);
or U9686 (N_9686,N_3286,N_4123);
or U9687 (N_9687,N_2782,N_931);
or U9688 (N_9688,N_2105,N_2464);
nand U9689 (N_9689,N_2792,N_3085);
and U9690 (N_9690,N_656,N_4318);
and U9691 (N_9691,N_4788,N_4290);
and U9692 (N_9692,N_1205,N_4745);
nand U9693 (N_9693,N_2781,N_3360);
and U9694 (N_9694,N_295,N_1890);
and U9695 (N_9695,N_436,N_1305);
xnor U9696 (N_9696,N_3951,N_3458);
nor U9697 (N_9697,N_2422,N_2125);
xnor U9698 (N_9698,N_3030,N_2445);
nand U9699 (N_9699,N_3304,N_1452);
or U9700 (N_9700,N_4684,N_3151);
nor U9701 (N_9701,N_3520,N_4098);
or U9702 (N_9702,N_3746,N_4477);
or U9703 (N_9703,N_1732,N_4248);
or U9704 (N_9704,N_4028,N_288);
and U9705 (N_9705,N_977,N_1107);
nor U9706 (N_9706,N_3783,N_4579);
xnor U9707 (N_9707,N_490,N_708);
nor U9708 (N_9708,N_599,N_3098);
xor U9709 (N_9709,N_1845,N_1518);
nand U9710 (N_9710,N_4203,N_1348);
or U9711 (N_9711,N_2268,N_2381);
nor U9712 (N_9712,N_601,N_2922);
or U9713 (N_9713,N_1012,N_4037);
and U9714 (N_9714,N_1764,N_2421);
nor U9715 (N_9715,N_1487,N_1733);
or U9716 (N_9716,N_322,N_3966);
nand U9717 (N_9717,N_1950,N_394);
nor U9718 (N_9718,N_4083,N_4579);
and U9719 (N_9719,N_2885,N_3447);
or U9720 (N_9720,N_179,N_4684);
or U9721 (N_9721,N_1193,N_2444);
and U9722 (N_9722,N_2921,N_3607);
and U9723 (N_9723,N_3382,N_1544);
nor U9724 (N_9724,N_4370,N_2855);
or U9725 (N_9725,N_4586,N_1290);
nor U9726 (N_9726,N_3481,N_3596);
and U9727 (N_9727,N_2521,N_3933);
or U9728 (N_9728,N_1678,N_2988);
nand U9729 (N_9729,N_461,N_2790);
or U9730 (N_9730,N_60,N_388);
xor U9731 (N_9731,N_739,N_1183);
nor U9732 (N_9732,N_1292,N_3961);
or U9733 (N_9733,N_4591,N_54);
or U9734 (N_9734,N_3417,N_3284);
and U9735 (N_9735,N_3332,N_252);
nand U9736 (N_9736,N_2226,N_3435);
and U9737 (N_9737,N_2720,N_667);
nand U9738 (N_9738,N_3388,N_2171);
nor U9739 (N_9739,N_3381,N_3547);
nor U9740 (N_9740,N_1770,N_2068);
or U9741 (N_9741,N_356,N_395);
nand U9742 (N_9742,N_3760,N_2152);
or U9743 (N_9743,N_2138,N_4449);
nor U9744 (N_9744,N_3471,N_3882);
and U9745 (N_9745,N_546,N_3193);
or U9746 (N_9746,N_1881,N_4875);
or U9747 (N_9747,N_3865,N_3577);
nand U9748 (N_9748,N_2431,N_1441);
or U9749 (N_9749,N_1184,N_4325);
and U9750 (N_9750,N_2950,N_4749);
and U9751 (N_9751,N_2005,N_4626);
nor U9752 (N_9752,N_2699,N_4067);
nand U9753 (N_9753,N_2144,N_4030);
and U9754 (N_9754,N_1355,N_2868);
nand U9755 (N_9755,N_4906,N_1909);
nand U9756 (N_9756,N_425,N_341);
and U9757 (N_9757,N_4543,N_1576);
nor U9758 (N_9758,N_1121,N_3435);
nand U9759 (N_9759,N_207,N_1134);
and U9760 (N_9760,N_1834,N_4137);
xor U9761 (N_9761,N_4440,N_4112);
and U9762 (N_9762,N_2488,N_4012);
nor U9763 (N_9763,N_1819,N_4244);
or U9764 (N_9764,N_2169,N_92);
nand U9765 (N_9765,N_3833,N_3138);
nand U9766 (N_9766,N_3174,N_1916);
nor U9767 (N_9767,N_3543,N_4333);
and U9768 (N_9768,N_1129,N_1664);
nand U9769 (N_9769,N_3004,N_3250);
or U9770 (N_9770,N_751,N_4378);
nor U9771 (N_9771,N_1082,N_4708);
nand U9772 (N_9772,N_4354,N_3);
and U9773 (N_9773,N_1863,N_4024);
nor U9774 (N_9774,N_1309,N_1497);
xor U9775 (N_9775,N_4434,N_3210);
or U9776 (N_9776,N_3452,N_339);
xor U9777 (N_9777,N_1031,N_1414);
and U9778 (N_9778,N_3671,N_2514);
nor U9779 (N_9779,N_3825,N_926);
nor U9780 (N_9780,N_3026,N_2832);
and U9781 (N_9781,N_3508,N_4896);
nand U9782 (N_9782,N_4471,N_4204);
nand U9783 (N_9783,N_409,N_4336);
nand U9784 (N_9784,N_3353,N_3438);
nor U9785 (N_9785,N_4510,N_2656);
or U9786 (N_9786,N_2186,N_207);
nand U9787 (N_9787,N_164,N_3720);
nor U9788 (N_9788,N_183,N_4619);
nand U9789 (N_9789,N_4276,N_685);
and U9790 (N_9790,N_3021,N_4816);
or U9791 (N_9791,N_1074,N_2388);
xor U9792 (N_9792,N_779,N_3785);
nand U9793 (N_9793,N_1783,N_2489);
or U9794 (N_9794,N_2147,N_4405);
and U9795 (N_9795,N_326,N_3488);
nand U9796 (N_9796,N_987,N_572);
nand U9797 (N_9797,N_97,N_3592);
nor U9798 (N_9798,N_777,N_886);
nand U9799 (N_9799,N_2886,N_3549);
or U9800 (N_9800,N_1694,N_2036);
nor U9801 (N_9801,N_1920,N_3955);
nand U9802 (N_9802,N_3266,N_4030);
nand U9803 (N_9803,N_1228,N_463);
nor U9804 (N_9804,N_4278,N_4843);
and U9805 (N_9805,N_4241,N_122);
or U9806 (N_9806,N_1058,N_985);
and U9807 (N_9807,N_150,N_36);
and U9808 (N_9808,N_405,N_2998);
nand U9809 (N_9809,N_3299,N_1704);
or U9810 (N_9810,N_1038,N_494);
nor U9811 (N_9811,N_2764,N_2416);
or U9812 (N_9812,N_2940,N_1039);
nor U9813 (N_9813,N_4414,N_4420);
nand U9814 (N_9814,N_1574,N_3116);
and U9815 (N_9815,N_4241,N_3332);
or U9816 (N_9816,N_453,N_3940);
nor U9817 (N_9817,N_714,N_492);
nor U9818 (N_9818,N_1282,N_2893);
nand U9819 (N_9819,N_1075,N_3227);
nand U9820 (N_9820,N_1251,N_4603);
and U9821 (N_9821,N_851,N_4230);
or U9822 (N_9822,N_1900,N_3925);
and U9823 (N_9823,N_337,N_2216);
nand U9824 (N_9824,N_1647,N_3150);
nor U9825 (N_9825,N_2746,N_209);
nor U9826 (N_9826,N_1860,N_1361);
nor U9827 (N_9827,N_1109,N_1887);
or U9828 (N_9828,N_895,N_3327);
or U9829 (N_9829,N_1109,N_2251);
or U9830 (N_9830,N_4864,N_3266);
or U9831 (N_9831,N_803,N_4569);
or U9832 (N_9832,N_3147,N_4140);
nand U9833 (N_9833,N_3515,N_4724);
or U9834 (N_9834,N_3583,N_2959);
nor U9835 (N_9835,N_1674,N_2);
nor U9836 (N_9836,N_1005,N_438);
and U9837 (N_9837,N_1797,N_2279);
or U9838 (N_9838,N_748,N_3346);
and U9839 (N_9839,N_3386,N_3345);
or U9840 (N_9840,N_813,N_4280);
nand U9841 (N_9841,N_1451,N_1572);
nor U9842 (N_9842,N_3876,N_4063);
nand U9843 (N_9843,N_1027,N_3052);
nor U9844 (N_9844,N_2144,N_2681);
nand U9845 (N_9845,N_4238,N_214);
nor U9846 (N_9846,N_4860,N_4523);
nand U9847 (N_9847,N_742,N_3599);
nor U9848 (N_9848,N_2811,N_2326);
nor U9849 (N_9849,N_3245,N_2976);
nand U9850 (N_9850,N_263,N_1452);
nor U9851 (N_9851,N_1810,N_2191);
or U9852 (N_9852,N_2664,N_385);
nor U9853 (N_9853,N_2935,N_4162);
nor U9854 (N_9854,N_2425,N_186);
nand U9855 (N_9855,N_3632,N_4387);
nor U9856 (N_9856,N_651,N_1022);
nor U9857 (N_9857,N_3242,N_1442);
or U9858 (N_9858,N_3463,N_3801);
nand U9859 (N_9859,N_1535,N_1859);
or U9860 (N_9860,N_1248,N_836);
nor U9861 (N_9861,N_2084,N_4139);
or U9862 (N_9862,N_1332,N_4000);
or U9863 (N_9863,N_2611,N_4357);
nor U9864 (N_9864,N_714,N_216);
nand U9865 (N_9865,N_3235,N_2840);
nor U9866 (N_9866,N_320,N_4906);
and U9867 (N_9867,N_607,N_2855);
and U9868 (N_9868,N_525,N_3971);
or U9869 (N_9869,N_4954,N_2808);
or U9870 (N_9870,N_3926,N_2656);
or U9871 (N_9871,N_4176,N_3648);
xor U9872 (N_9872,N_2988,N_3827);
or U9873 (N_9873,N_4069,N_2505);
nor U9874 (N_9874,N_4105,N_1970);
and U9875 (N_9875,N_1600,N_614);
nand U9876 (N_9876,N_3151,N_3973);
and U9877 (N_9877,N_193,N_3891);
or U9878 (N_9878,N_2472,N_1666);
or U9879 (N_9879,N_2227,N_4406);
or U9880 (N_9880,N_2293,N_1262);
nor U9881 (N_9881,N_334,N_2137);
or U9882 (N_9882,N_2069,N_496);
nand U9883 (N_9883,N_1908,N_2812);
and U9884 (N_9884,N_2561,N_1873);
or U9885 (N_9885,N_4989,N_444);
and U9886 (N_9886,N_4668,N_2599);
nor U9887 (N_9887,N_4373,N_1430);
and U9888 (N_9888,N_1578,N_3904);
and U9889 (N_9889,N_431,N_89);
nor U9890 (N_9890,N_4537,N_2424);
and U9891 (N_9891,N_4174,N_2787);
nor U9892 (N_9892,N_969,N_137);
or U9893 (N_9893,N_843,N_782);
or U9894 (N_9894,N_368,N_2203);
xnor U9895 (N_9895,N_4989,N_2837);
and U9896 (N_9896,N_4397,N_3346);
nand U9897 (N_9897,N_4445,N_2068);
nor U9898 (N_9898,N_33,N_2707);
xor U9899 (N_9899,N_4568,N_1209);
nor U9900 (N_9900,N_930,N_4260);
nor U9901 (N_9901,N_4424,N_1621);
or U9902 (N_9902,N_4458,N_1317);
and U9903 (N_9903,N_3879,N_942);
or U9904 (N_9904,N_1876,N_1280);
or U9905 (N_9905,N_4447,N_187);
and U9906 (N_9906,N_133,N_3174);
nor U9907 (N_9907,N_4148,N_523);
or U9908 (N_9908,N_228,N_2300);
nor U9909 (N_9909,N_377,N_213);
and U9910 (N_9910,N_2975,N_2379);
nor U9911 (N_9911,N_1532,N_2122);
nand U9912 (N_9912,N_1276,N_4528);
nor U9913 (N_9913,N_873,N_2835);
and U9914 (N_9914,N_2997,N_4633);
nand U9915 (N_9915,N_1699,N_1281);
and U9916 (N_9916,N_2589,N_4826);
nand U9917 (N_9917,N_4630,N_2202);
nand U9918 (N_9918,N_3450,N_2373);
or U9919 (N_9919,N_4247,N_3101);
and U9920 (N_9920,N_1547,N_930);
nand U9921 (N_9921,N_4095,N_4931);
or U9922 (N_9922,N_586,N_2769);
or U9923 (N_9923,N_3263,N_1714);
nand U9924 (N_9924,N_4893,N_258);
nand U9925 (N_9925,N_1181,N_3053);
nand U9926 (N_9926,N_246,N_2217);
and U9927 (N_9927,N_3281,N_4204);
nand U9928 (N_9928,N_3988,N_4291);
nand U9929 (N_9929,N_4555,N_2822);
nand U9930 (N_9930,N_2596,N_1312);
nor U9931 (N_9931,N_4758,N_4373);
nor U9932 (N_9932,N_4125,N_3626);
nand U9933 (N_9933,N_4040,N_2265);
nor U9934 (N_9934,N_3602,N_3848);
nand U9935 (N_9935,N_1849,N_4423);
nor U9936 (N_9936,N_1803,N_3181);
nand U9937 (N_9937,N_2949,N_3716);
or U9938 (N_9938,N_617,N_2448);
nand U9939 (N_9939,N_746,N_4741);
nor U9940 (N_9940,N_3106,N_4456);
nand U9941 (N_9941,N_2171,N_3694);
and U9942 (N_9942,N_4346,N_269);
nand U9943 (N_9943,N_2622,N_3209);
and U9944 (N_9944,N_4143,N_3287);
nor U9945 (N_9945,N_3097,N_168);
nor U9946 (N_9946,N_3901,N_573);
nor U9947 (N_9947,N_4369,N_3948);
nand U9948 (N_9948,N_1774,N_3588);
nand U9949 (N_9949,N_1935,N_4427);
nor U9950 (N_9950,N_240,N_3700);
and U9951 (N_9951,N_1539,N_4654);
or U9952 (N_9952,N_1748,N_3668);
and U9953 (N_9953,N_1260,N_350);
nand U9954 (N_9954,N_1004,N_290);
nand U9955 (N_9955,N_559,N_4230);
and U9956 (N_9956,N_806,N_2056);
or U9957 (N_9957,N_4412,N_1225);
or U9958 (N_9958,N_37,N_4095);
nand U9959 (N_9959,N_3148,N_355);
nor U9960 (N_9960,N_3821,N_3964);
nand U9961 (N_9961,N_3216,N_1284);
nor U9962 (N_9962,N_2176,N_1344);
nor U9963 (N_9963,N_4578,N_2052);
nor U9964 (N_9964,N_4125,N_237);
nand U9965 (N_9965,N_3586,N_4634);
and U9966 (N_9966,N_1595,N_1853);
nor U9967 (N_9967,N_3211,N_3253);
and U9968 (N_9968,N_3868,N_4391);
nor U9969 (N_9969,N_3247,N_1683);
or U9970 (N_9970,N_325,N_1660);
nand U9971 (N_9971,N_4835,N_1805);
nor U9972 (N_9972,N_776,N_3071);
and U9973 (N_9973,N_4774,N_338);
nor U9974 (N_9974,N_2480,N_4438);
and U9975 (N_9975,N_1989,N_923);
and U9976 (N_9976,N_3604,N_1474);
nor U9977 (N_9977,N_3458,N_1296);
and U9978 (N_9978,N_1127,N_289);
and U9979 (N_9979,N_2688,N_1595);
nand U9980 (N_9980,N_3868,N_2803);
nor U9981 (N_9981,N_791,N_2187);
and U9982 (N_9982,N_2347,N_2721);
nand U9983 (N_9983,N_4238,N_860);
nor U9984 (N_9984,N_4073,N_2505);
or U9985 (N_9985,N_1867,N_610);
and U9986 (N_9986,N_1485,N_2915);
nor U9987 (N_9987,N_2925,N_2376);
nor U9988 (N_9988,N_4625,N_567);
nor U9989 (N_9989,N_4224,N_2639);
or U9990 (N_9990,N_2364,N_1311);
xor U9991 (N_9991,N_4997,N_1367);
and U9992 (N_9992,N_453,N_247);
nand U9993 (N_9993,N_1735,N_2647);
and U9994 (N_9994,N_1919,N_3368);
and U9995 (N_9995,N_1959,N_3496);
nand U9996 (N_9996,N_3624,N_4849);
and U9997 (N_9997,N_514,N_4075);
nor U9998 (N_9998,N_2739,N_3425);
or U9999 (N_9999,N_3102,N_3483);
and U10000 (N_10000,N_6513,N_5283);
or U10001 (N_10001,N_7641,N_5628);
and U10002 (N_10002,N_7766,N_8936);
and U10003 (N_10003,N_6687,N_6112);
or U10004 (N_10004,N_7532,N_5607);
nand U10005 (N_10005,N_7578,N_7243);
or U10006 (N_10006,N_6878,N_7807);
nand U10007 (N_10007,N_7471,N_6138);
nor U10008 (N_10008,N_6604,N_6169);
nand U10009 (N_10009,N_5205,N_9496);
or U10010 (N_10010,N_9492,N_9775);
nand U10011 (N_10011,N_6275,N_6538);
or U10012 (N_10012,N_5106,N_7299);
and U10013 (N_10013,N_9653,N_5510);
and U10014 (N_10014,N_6299,N_9230);
or U10015 (N_10015,N_8991,N_5137);
nor U10016 (N_10016,N_9886,N_5162);
nand U10017 (N_10017,N_8228,N_5877);
and U10018 (N_10018,N_6623,N_7417);
and U10019 (N_10019,N_5164,N_5840);
and U10020 (N_10020,N_7403,N_8575);
and U10021 (N_10021,N_9415,N_7287);
nand U10022 (N_10022,N_6931,N_5751);
nand U10023 (N_10023,N_9452,N_7272);
nand U10024 (N_10024,N_7358,N_6759);
nor U10025 (N_10025,N_8609,N_7452);
nand U10026 (N_10026,N_7431,N_5631);
or U10027 (N_10027,N_7362,N_9229);
or U10028 (N_10028,N_9550,N_5854);
and U10029 (N_10029,N_9377,N_7119);
xor U10030 (N_10030,N_8368,N_7945);
nor U10031 (N_10031,N_9833,N_7900);
nor U10032 (N_10032,N_9036,N_6692);
nor U10033 (N_10033,N_7803,N_8824);
or U10034 (N_10034,N_5421,N_9661);
and U10035 (N_10035,N_8344,N_7921);
nor U10036 (N_10036,N_6755,N_5154);
or U10037 (N_10037,N_7124,N_6395);
and U10038 (N_10038,N_5839,N_9147);
or U10039 (N_10039,N_7639,N_9395);
or U10040 (N_10040,N_8295,N_7042);
nor U10041 (N_10041,N_6521,N_8735);
or U10042 (N_10042,N_7758,N_7721);
nand U10043 (N_10043,N_7208,N_6379);
nand U10044 (N_10044,N_5379,N_8202);
and U10045 (N_10045,N_7582,N_6718);
and U10046 (N_10046,N_5117,N_8549);
or U10047 (N_10047,N_9509,N_6573);
xnor U10048 (N_10048,N_6296,N_8263);
and U10049 (N_10049,N_5515,N_9828);
nand U10050 (N_10050,N_5770,N_5655);
nor U10051 (N_10051,N_7810,N_7646);
nor U10052 (N_10052,N_7987,N_7581);
nand U10053 (N_10053,N_6602,N_9345);
and U10054 (N_10054,N_6688,N_8853);
or U10055 (N_10055,N_7034,N_7770);
and U10056 (N_10056,N_7603,N_7269);
and U10057 (N_10057,N_9453,N_8501);
and U10058 (N_10058,N_9614,N_9787);
and U10059 (N_10059,N_5139,N_5358);
and U10060 (N_10060,N_9236,N_7896);
nand U10061 (N_10061,N_6305,N_6029);
nand U10062 (N_10062,N_5938,N_5698);
or U10063 (N_10063,N_7478,N_6807);
or U10064 (N_10064,N_7301,N_8893);
and U10065 (N_10065,N_9458,N_8543);
nor U10066 (N_10066,N_6348,N_7214);
or U10067 (N_10067,N_9414,N_9923);
nor U10068 (N_10068,N_6276,N_6376);
and U10069 (N_10069,N_7405,N_5375);
and U10070 (N_10070,N_6202,N_6765);
or U10071 (N_10071,N_6026,N_9922);
nor U10072 (N_10072,N_5058,N_8724);
nand U10073 (N_10073,N_8426,N_5883);
nand U10074 (N_10074,N_6754,N_8156);
nor U10075 (N_10075,N_9276,N_9843);
xnor U10076 (N_10076,N_8270,N_5925);
nand U10077 (N_10077,N_6283,N_5913);
nor U10078 (N_10078,N_8705,N_9440);
nand U10079 (N_10079,N_8029,N_8173);
nor U10080 (N_10080,N_5753,N_6634);
and U10081 (N_10081,N_9356,N_9609);
nor U10082 (N_10082,N_8244,N_6678);
or U10083 (N_10083,N_5734,N_8178);
nor U10084 (N_10084,N_9920,N_9026);
nand U10085 (N_10085,N_6076,N_7497);
nand U10086 (N_10086,N_6815,N_7412);
nor U10087 (N_10087,N_8036,N_5987);
nand U10088 (N_10088,N_7141,N_5048);
nand U10089 (N_10089,N_6811,N_9016);
or U10090 (N_10090,N_7796,N_5397);
and U10091 (N_10091,N_5612,N_5077);
nand U10092 (N_10092,N_6371,N_7589);
nand U10093 (N_10093,N_5694,N_5714);
nand U10094 (N_10094,N_7442,N_6748);
nand U10095 (N_10095,N_6546,N_7339);
and U10096 (N_10096,N_5941,N_9112);
and U10097 (N_10097,N_8455,N_6410);
and U10098 (N_10098,N_9839,N_6558);
nor U10099 (N_10099,N_7284,N_9433);
nand U10100 (N_10100,N_9785,N_6819);
or U10101 (N_10101,N_8741,N_8261);
and U10102 (N_10102,N_5282,N_5492);
and U10103 (N_10103,N_9547,N_6812);
nor U10104 (N_10104,N_6857,N_6825);
nand U10105 (N_10105,N_5614,N_8334);
nand U10106 (N_10106,N_6249,N_5231);
nor U10107 (N_10107,N_6928,N_7942);
or U10108 (N_10108,N_9817,N_8820);
and U10109 (N_10109,N_7003,N_8767);
and U10110 (N_10110,N_5999,N_9949);
nor U10111 (N_10111,N_5656,N_5210);
nor U10112 (N_10112,N_9362,N_7677);
or U10113 (N_10113,N_6971,N_5452);
and U10114 (N_10114,N_5788,N_5316);
and U10115 (N_10115,N_6566,N_7701);
and U10116 (N_10116,N_9764,N_5616);
or U10117 (N_10117,N_9318,N_5769);
nand U10118 (N_10118,N_6149,N_5519);
nand U10119 (N_10119,N_5838,N_5212);
and U10120 (N_10120,N_7157,N_6702);
and U10121 (N_10121,N_6981,N_9611);
nand U10122 (N_10122,N_5223,N_8372);
and U10123 (N_10123,N_9728,N_9089);
nor U10124 (N_10124,N_5267,N_8114);
nor U10125 (N_10125,N_7710,N_9140);
or U10126 (N_10126,N_7767,N_6116);
nand U10127 (N_10127,N_7369,N_9536);
nand U10128 (N_10128,N_9128,N_7467);
nor U10129 (N_10129,N_7436,N_7391);
nor U10130 (N_10130,N_5356,N_8191);
nor U10131 (N_10131,N_7837,N_6552);
nor U10132 (N_10132,N_7748,N_8307);
nand U10133 (N_10133,N_7516,N_7464);
nor U10134 (N_10134,N_8214,N_6631);
and U10135 (N_10135,N_5449,N_6096);
nor U10136 (N_10136,N_6586,N_9867);
and U10137 (N_10137,N_7112,N_5026);
nand U10138 (N_10138,N_6427,N_8355);
nand U10139 (N_10139,N_8409,N_7712);
xor U10140 (N_10140,N_6053,N_8971);
and U10141 (N_10141,N_5665,N_6961);
and U10142 (N_10142,N_7596,N_5398);
nand U10143 (N_10143,N_7222,N_9371);
nand U10144 (N_10144,N_7585,N_5371);
nor U10145 (N_10145,N_8927,N_7292);
nor U10146 (N_10146,N_9392,N_5443);
and U10147 (N_10147,N_9824,N_8618);
nor U10148 (N_10148,N_9664,N_8034);
or U10149 (N_10149,N_5095,N_5464);
nand U10150 (N_10150,N_7021,N_6663);
xnor U10151 (N_10151,N_5150,N_6821);
and U10152 (N_10152,N_9635,N_8189);
and U10153 (N_10153,N_9482,N_9374);
nor U10154 (N_10154,N_8364,N_5457);
or U10155 (N_10155,N_5257,N_9790);
and U10156 (N_10156,N_7859,N_6469);
nor U10157 (N_10157,N_8674,N_9028);
nor U10158 (N_10158,N_5730,N_8155);
nor U10159 (N_10159,N_7634,N_9658);
nand U10160 (N_10160,N_7909,N_8584);
nor U10161 (N_10161,N_6592,N_9760);
and U10162 (N_10162,N_9270,N_9917);
or U10163 (N_10163,N_8693,N_6222);
or U10164 (N_10164,N_8947,N_9302);
nor U10165 (N_10165,N_5045,N_5046);
nor U10166 (N_10166,N_7763,N_5721);
or U10167 (N_10167,N_7819,N_5486);
nor U10168 (N_10168,N_7468,N_9445);
or U10169 (N_10169,N_8143,N_8630);
or U10170 (N_10170,N_5991,N_7813);
nand U10171 (N_10171,N_9424,N_7308);
and U10172 (N_10172,N_9514,N_9666);
nor U10173 (N_10173,N_6040,N_5467);
nand U10174 (N_10174,N_5794,N_8049);
or U10175 (N_10175,N_6715,N_7707);
or U10176 (N_10176,N_7876,N_9731);
and U10177 (N_10177,N_9282,N_9934);
nand U10178 (N_10178,N_8287,N_8386);
or U10179 (N_10179,N_6813,N_6417);
or U10180 (N_10180,N_6695,N_9122);
nand U10181 (N_10181,N_9014,N_7061);
or U10182 (N_10182,N_8210,N_7620);
xor U10183 (N_10183,N_7475,N_5374);
or U10184 (N_10184,N_8788,N_6262);
and U10185 (N_10185,N_6062,N_7298);
nor U10186 (N_10186,N_7846,N_7345);
xnor U10187 (N_10187,N_8476,N_9132);
nand U10188 (N_10188,N_5044,N_7450);
and U10189 (N_10189,N_9589,N_8774);
nand U10190 (N_10190,N_5113,N_8753);
nor U10191 (N_10191,N_8236,N_6609);
nand U10192 (N_10192,N_5797,N_7420);
nand U10193 (N_10193,N_5448,N_8614);
and U10194 (N_10194,N_6508,N_6805);
nand U10195 (N_10195,N_8610,N_9491);
nand U10196 (N_10196,N_8134,N_8598);
nor U10197 (N_10197,N_9891,N_5100);
nand U10198 (N_10198,N_9111,N_5388);
and U10199 (N_10199,N_8954,N_8527);
nor U10200 (N_10200,N_5440,N_5891);
nor U10201 (N_10201,N_8812,N_8994);
and U10202 (N_10202,N_7444,N_5109);
nand U10203 (N_10203,N_7191,N_7280);
nor U10204 (N_10204,N_9357,N_6505);
or U10205 (N_10205,N_6545,N_7249);
nand U10206 (N_10206,N_9504,N_8343);
or U10207 (N_10207,N_7576,N_7728);
nor U10208 (N_10208,N_6480,N_7381);
or U10209 (N_10209,N_8387,N_7289);
nor U10210 (N_10210,N_6921,N_9237);
and U10211 (N_10211,N_9621,N_8897);
nand U10212 (N_10212,N_7938,N_7167);
or U10213 (N_10213,N_6372,N_8212);
xor U10214 (N_10214,N_6297,N_8463);
nor U10215 (N_10215,N_7519,N_5034);
nand U10216 (N_10216,N_6129,N_6881);
and U10217 (N_10217,N_6122,N_6132);
and U10218 (N_10218,N_6875,N_6436);
or U10219 (N_10219,N_9720,N_5285);
and U10220 (N_10220,N_9681,N_8608);
nand U10221 (N_10221,N_5686,N_9263);
or U10222 (N_10222,N_7015,N_8567);
nand U10223 (N_10223,N_9960,N_5272);
nor U10224 (N_10224,N_7103,N_6996);
nor U10225 (N_10225,N_6041,N_5343);
or U10226 (N_10226,N_8417,N_8923);
nor U10227 (N_10227,N_7773,N_8087);
and U10228 (N_10228,N_5323,N_7880);
nor U10229 (N_10229,N_9228,N_8699);
or U10230 (N_10230,N_6253,N_6445);
or U10231 (N_10231,N_7919,N_8999);
nor U10232 (N_10232,N_6488,N_9094);
or U10233 (N_10233,N_7703,N_8206);
or U10234 (N_10234,N_5978,N_8806);
nor U10235 (N_10235,N_7194,N_7418);
and U10236 (N_10236,N_6413,N_7877);
nand U10237 (N_10237,N_7072,N_5597);
nand U10238 (N_10238,N_8321,N_7833);
and U10239 (N_10239,N_9042,N_6017);
nand U10240 (N_10240,N_9644,N_6037);
xnor U10241 (N_10241,N_7386,N_8815);
and U10242 (N_10242,N_8542,N_8240);
or U10243 (N_10243,N_5057,N_7598);
nor U10244 (N_10244,N_8733,N_6817);
nand U10245 (N_10245,N_6452,N_6373);
or U10246 (N_10246,N_7500,N_9900);
or U10247 (N_10247,N_9989,N_9770);
or U10248 (N_10248,N_7951,N_7943);
nor U10249 (N_10249,N_7740,N_5477);
and U10250 (N_10250,N_5684,N_6824);
nor U10251 (N_10251,N_5277,N_8827);
nor U10252 (N_10252,N_8057,N_7346);
nor U10253 (N_10253,N_8835,N_8989);
or U10254 (N_10254,N_6635,N_9544);
nand U10255 (N_10255,N_6318,N_8085);
and U10256 (N_10256,N_5293,N_8770);
and U10257 (N_10257,N_7563,N_7929);
and U10258 (N_10258,N_5939,N_5031);
nand U10259 (N_10259,N_8582,N_6031);
nor U10260 (N_10260,N_5561,N_6752);
nand U10261 (N_10261,N_8775,N_9078);
xor U10262 (N_10262,N_8934,N_6871);
or U10263 (N_10263,N_5707,N_7676);
and U10264 (N_10264,N_9901,N_7507);
nor U10265 (N_10265,N_7889,N_9224);
or U10266 (N_10266,N_8347,N_6482);
nor U10267 (N_10267,N_5042,N_9805);
nor U10268 (N_10268,N_6915,N_5322);
nand U10269 (N_10269,N_9397,N_7761);
or U10270 (N_10270,N_6081,N_5787);
xor U10271 (N_10271,N_9197,N_6330);
nor U10272 (N_10272,N_7648,N_6650);
and U10273 (N_10273,N_9876,N_8447);
nor U10274 (N_10274,N_7808,N_9628);
and U10275 (N_10275,N_7658,N_5529);
nor U10276 (N_10276,N_5158,N_6048);
or U10277 (N_10277,N_7526,N_5481);
or U10278 (N_10278,N_8219,N_8249);
xor U10279 (N_10279,N_5260,N_6851);
nor U10280 (N_10280,N_8916,N_5414);
or U10281 (N_10281,N_9388,N_7623);
or U10282 (N_10282,N_5600,N_6547);
and U10283 (N_10283,N_6137,N_5014);
xnor U10284 (N_10284,N_8856,N_9921);
nand U10285 (N_10285,N_9455,N_9725);
nor U10286 (N_10286,N_6704,N_8140);
or U10287 (N_10287,N_7057,N_8793);
nor U10288 (N_10288,N_5670,N_9002);
nor U10289 (N_10289,N_6610,N_7499);
xnor U10290 (N_10290,N_6432,N_9716);
nand U10291 (N_10291,N_6437,N_5276);
or U10292 (N_10292,N_5613,N_5965);
nor U10293 (N_10293,N_7357,N_8292);
nand U10294 (N_10294,N_8064,N_9786);
nor U10295 (N_10295,N_7739,N_8404);
and U10296 (N_10296,N_7400,N_8267);
nor U10297 (N_10297,N_7262,N_6574);
and U10298 (N_10298,N_8102,N_9209);
and U10299 (N_10299,N_8412,N_6839);
or U10300 (N_10300,N_6886,N_8425);
nor U10301 (N_10301,N_6594,N_7312);
or U10302 (N_10302,N_6016,N_8318);
nand U10303 (N_10303,N_5022,N_5903);
and U10304 (N_10304,N_9640,N_5653);
nand U10305 (N_10305,N_6233,N_6471);
or U10306 (N_10306,N_8520,N_5220);
nor U10307 (N_10307,N_5270,N_8510);
nor U10308 (N_10308,N_5855,N_7679);
and U10309 (N_10309,N_6158,N_8957);
nor U10310 (N_10310,N_8588,N_7363);
and U10311 (N_10311,N_6911,N_8866);
and U10312 (N_10312,N_6294,N_9470);
nand U10313 (N_10313,N_8784,N_8148);
and U10314 (N_10314,N_7433,N_7466);
nor U10315 (N_10315,N_8833,N_6385);
nand U10316 (N_10316,N_5327,N_5722);
nand U10317 (N_10317,N_9821,N_6674);
or U10318 (N_10318,N_8882,N_5630);
and U10319 (N_10319,N_5284,N_9849);
and U10320 (N_10320,N_9338,N_7040);
and U10321 (N_10321,N_7958,N_9620);
nand U10322 (N_10322,N_9796,N_8319);
nor U10323 (N_10323,N_7046,N_8294);
or U10324 (N_10324,N_5354,N_8738);
nand U10325 (N_10325,N_5920,N_5782);
or U10326 (N_10326,N_8621,N_6406);
nand U10327 (N_10327,N_7760,N_7538);
nand U10328 (N_10328,N_5326,N_8063);
nand U10329 (N_10329,N_7399,N_6567);
nor U10330 (N_10330,N_6734,N_8717);
and U10331 (N_10331,N_5271,N_7528);
nand U10332 (N_10332,N_7008,N_9826);
nor U10333 (N_10333,N_9518,N_7587);
nor U10334 (N_10334,N_8782,N_9004);
or U10335 (N_10335,N_5640,N_5689);
nor U10336 (N_10336,N_8496,N_9659);
nand U10337 (N_10337,N_6421,N_5344);
nor U10338 (N_10338,N_6738,N_5501);
xor U10339 (N_10339,N_8227,N_5902);
nor U10340 (N_10340,N_8495,N_5054);
nand U10341 (N_10341,N_8781,N_9945);
and U10342 (N_10342,N_5017,N_9800);
xnor U10343 (N_10343,N_6142,N_7931);
and U10344 (N_10344,N_9473,N_8195);
nand U10345 (N_10345,N_5625,N_5914);
nand U10346 (N_10346,N_8459,N_8975);
nand U10347 (N_10347,N_7747,N_9866);
nand U10348 (N_10348,N_9349,N_5424);
and U10349 (N_10349,N_5065,N_6953);
or U10350 (N_10350,N_6948,N_7274);
or U10351 (N_10351,N_9296,N_7695);
and U10352 (N_10352,N_8314,N_9510);
nor U10353 (N_10353,N_8253,N_5837);
and U10354 (N_10354,N_9757,N_9535);
and U10355 (N_10355,N_5248,N_5079);
nor U10356 (N_10356,N_5678,N_5831);
and U10357 (N_10357,N_7470,N_9006);
and U10358 (N_10358,N_8059,N_8291);
nand U10359 (N_10359,N_9558,N_6221);
nand U10360 (N_10360,N_8147,N_6994);
nor U10361 (N_10361,N_5559,N_7861);
and U10362 (N_10362,N_7210,N_9878);
nand U10363 (N_10363,N_8084,N_9950);
and U10364 (N_10364,N_8054,N_9802);
or U10365 (N_10365,N_9673,N_6232);
and U10366 (N_10366,N_5055,N_9501);
or U10367 (N_10367,N_5222,N_8904);
nand U10368 (N_10368,N_8963,N_7074);
nand U10369 (N_10369,N_9836,N_6295);
and U10370 (N_10370,N_5206,N_7177);
xor U10371 (N_10371,N_7447,N_6743);
or U10372 (N_10372,N_9413,N_7937);
nor U10373 (N_10373,N_8657,N_5971);
nand U10374 (N_10374,N_7899,N_8732);
nand U10375 (N_10375,N_5850,N_6761);
or U10376 (N_10376,N_7370,N_5554);
or U10377 (N_10377,N_6261,N_8796);
nand U10378 (N_10378,N_5273,N_5660);
and U10379 (N_10379,N_6106,N_7028);
nor U10380 (N_10380,N_5713,N_7195);
or U10381 (N_10381,N_5442,N_9541);
or U10382 (N_10382,N_8902,N_9292);
or U10383 (N_10383,N_8697,N_9751);
and U10384 (N_10384,N_7482,N_5899);
nand U10385 (N_10385,N_8356,N_5986);
nor U10386 (N_10386,N_6159,N_7957);
nand U10387 (N_10387,N_7781,N_7041);
nor U10388 (N_10388,N_6357,N_6783);
nand U10389 (N_10389,N_7635,N_6331);
and U10390 (N_10390,N_5310,N_6234);
or U10391 (N_10391,N_5423,N_8216);
or U10392 (N_10392,N_9148,N_5256);
and U10393 (N_10393,N_6840,N_9598);
or U10394 (N_10394,N_8576,N_5595);
nor U10395 (N_10395,N_6684,N_6887);
or U10396 (N_10396,N_8174,N_7973);
and U10397 (N_10397,N_8864,N_5916);
and U10398 (N_10398,N_9762,N_8324);
nand U10399 (N_10399,N_5428,N_6309);
or U10400 (N_10400,N_6900,N_5433);
or U10401 (N_10401,N_7114,N_5926);
nand U10402 (N_10402,N_7137,N_9521);
nor U10403 (N_10403,N_6367,N_8199);
and U10404 (N_10404,N_5191,N_9506);
and U10405 (N_10405,N_6278,N_9688);
or U10406 (N_10406,N_6272,N_8393);
nand U10407 (N_10407,N_5781,N_5008);
or U10408 (N_10408,N_9394,N_5437);
nor U10409 (N_10409,N_6866,N_8286);
nor U10410 (N_10410,N_9604,N_7533);
and U10411 (N_10411,N_8505,N_6519);
nor U10412 (N_10412,N_9743,N_8467);
nor U10413 (N_10413,N_6174,N_8096);
nor U10414 (N_10414,N_7671,N_5967);
nor U10415 (N_10415,N_6838,N_6771);
or U10416 (N_10416,N_7784,N_9410);
and U10417 (N_10417,N_9571,N_7465);
nor U10418 (N_10418,N_7058,N_7534);
or U10419 (N_10419,N_7488,N_5497);
nand U10420 (N_10420,N_6263,N_6798);
nor U10421 (N_10421,N_8332,N_8370);
nand U10422 (N_10422,N_6269,N_9141);
or U10423 (N_10423,N_7143,N_7787);
or U10424 (N_10424,N_8785,N_8497);
or U10425 (N_10425,N_5247,N_6700);
or U10426 (N_10426,N_9380,N_6560);
or U10427 (N_10427,N_8573,N_5199);
xnor U10428 (N_10428,N_9336,N_6117);
nand U10429 (N_10429,N_7811,N_8534);
nor U10430 (N_10430,N_8335,N_9534);
nor U10431 (N_10431,N_7515,N_6633);
or U10432 (N_10432,N_8254,N_6997);
nand U10433 (N_10433,N_7368,N_6032);
nand U10434 (N_10434,N_8560,N_7304);
nand U10435 (N_10435,N_5943,N_6920);
nor U10436 (N_10436,N_6964,N_8099);
nand U10437 (N_10437,N_9530,N_8132);
nor U10438 (N_10438,N_9119,N_5330);
nand U10439 (N_10439,N_9246,N_9031);
or U10440 (N_10440,N_8969,N_9074);
or U10441 (N_10441,N_7316,N_8622);
nor U10442 (N_10442,N_9293,N_6936);
or U10443 (N_10443,N_5380,N_5708);
nor U10444 (N_10444,N_5063,N_7204);
or U10445 (N_10445,N_5025,N_8456);
nor U10446 (N_10446,N_6532,N_7564);
or U10447 (N_10447,N_9647,N_7759);
or U10448 (N_10448,N_8648,N_8293);
nand U10449 (N_10449,N_9733,N_6027);
or U10450 (N_10450,N_9166,N_6459);
or U10451 (N_10451,N_7798,N_5833);
nand U10452 (N_10452,N_8973,N_9918);
nand U10453 (N_10453,N_8278,N_5579);
or U10454 (N_10454,N_7451,N_8358);
and U10455 (N_10455,N_9971,N_5626);
nand U10456 (N_10456,N_7215,N_9245);
nand U10457 (N_10457,N_6760,N_9158);
and U10458 (N_10458,N_9581,N_6615);
and U10459 (N_10459,N_8751,N_7799);
nand U10460 (N_10460,N_6717,N_7014);
or U10461 (N_10461,N_8929,N_9093);
or U10462 (N_10462,N_6462,N_7754);
or U10463 (N_10463,N_5824,N_7786);
nor U10464 (N_10464,N_7012,N_8110);
nor U10465 (N_10465,N_8094,N_6796);
nor U10466 (N_10466,N_7199,N_9761);
and U10467 (N_10467,N_8488,N_8400);
or U10468 (N_10468,N_9970,N_7537);
nand U10469 (N_10469,N_9966,N_8274);
nor U10470 (N_10470,N_9386,N_9864);
nand U10471 (N_10471,N_6491,N_6876);
or U10472 (N_10472,N_7925,N_5802);
and U10473 (N_10473,N_7725,N_6618);
and U10474 (N_10474,N_7765,N_9870);
or U10475 (N_10475,N_9124,N_7100);
xor U10476 (N_10476,N_5551,N_7340);
and U10477 (N_10477,N_6596,N_9788);
nor U10478 (N_10478,N_5750,N_9241);
and U10479 (N_10479,N_7002,N_8982);
and U10480 (N_10480,N_8153,N_8887);
nor U10481 (N_10481,N_9634,N_6733);
nand U10482 (N_10482,N_7764,N_8097);
nand U10483 (N_10483,N_6528,N_5923);
nor U10484 (N_10484,N_9701,N_8689);
or U10485 (N_10485,N_6914,N_6083);
or U10486 (N_10486,N_9759,N_9645);
nand U10487 (N_10487,N_5078,N_6363);
nor U10488 (N_10488,N_7329,N_8823);
nand U10489 (N_10489,N_7966,N_6844);
and U10490 (N_10490,N_6526,N_7715);
nand U10491 (N_10491,N_7377,N_9330);
nand U10492 (N_10492,N_9834,N_7752);
or U10493 (N_10493,N_9915,N_5495);
nand U10494 (N_10494,N_7353,N_7882);
nor U10495 (N_10495,N_8531,N_9744);
and U10496 (N_10496,N_7347,N_7731);
nand U10497 (N_10497,N_9846,N_7897);
or U10498 (N_10498,N_7780,N_7873);
nand U10499 (N_10499,N_8707,N_5606);
nor U10500 (N_10500,N_9676,N_8915);
nand U10501 (N_10501,N_6856,N_5460);
nand U10502 (N_10502,N_8678,N_8894);
nand U10503 (N_10503,N_5545,N_7930);
nand U10504 (N_10504,N_7556,N_9531);
or U10505 (N_10505,N_5856,N_6312);
or U10506 (N_10506,N_5834,N_8439);
nand U10507 (N_10507,N_7278,N_8627);
nand U10508 (N_10508,N_7256,N_9425);
nor U10509 (N_10509,N_9056,N_8040);
or U10510 (N_10510,N_8419,N_8848);
nor U10511 (N_10511,N_9144,N_8427);
or U10512 (N_10512,N_9264,N_8171);
nand U10513 (N_10513,N_7883,N_9832);
nor U10514 (N_10514,N_9961,N_7890);
nand U10515 (N_10515,N_5860,N_5615);
and U10516 (N_10516,N_7484,N_7914);
nand U10517 (N_10517,N_8960,N_9643);
nor U10518 (N_10518,N_5325,N_8571);
and U10519 (N_10519,N_8048,N_5441);
and U10520 (N_10520,N_6319,N_5146);
and U10521 (N_10521,N_6321,N_5992);
nor U10522 (N_10522,N_6778,N_8093);
nor U10523 (N_10523,N_5890,N_8625);
nand U10524 (N_10524,N_7800,N_6183);
and U10525 (N_10525,N_9485,N_8250);
nor U10526 (N_10526,N_5413,N_7672);
or U10527 (N_10527,N_6861,N_7423);
nand U10528 (N_10528,N_9472,N_5588);
nor U10529 (N_10529,N_9239,N_5024);
or U10530 (N_10530,N_7115,N_8892);
nand U10531 (N_10531,N_5970,N_9650);
and U10532 (N_10532,N_9909,N_7501);
nor U10533 (N_10533,N_5634,N_7239);
and U10534 (N_10534,N_9953,N_8329);
nor U10535 (N_10535,N_6584,N_8695);
or U10536 (N_10536,N_9792,N_9546);
or U10537 (N_10537,N_5532,N_6885);
and U10538 (N_10538,N_5308,N_8222);
or U10539 (N_10539,N_5124,N_6624);
nand U10540 (N_10540,N_6972,N_9622);
and U10541 (N_10541,N_8819,N_5743);
nor U10542 (N_10542,N_9125,N_8655);
or U10543 (N_10543,N_5604,N_9668);
or U10544 (N_10544,N_5863,N_9862);
and U10545 (N_10545,N_5204,N_6454);
xnor U10546 (N_10546,N_8579,N_8925);
and U10547 (N_10547,N_8095,N_5956);
or U10548 (N_10548,N_5530,N_8685);
or U10549 (N_10549,N_7597,N_8883);
nand U10550 (N_10550,N_5426,N_6003);
nor U10551 (N_10551,N_8224,N_5773);
nor U10552 (N_10552,N_9010,N_7974);
xnor U10553 (N_10553,N_8503,N_9454);
and U10554 (N_10554,N_7742,N_8818);
nand U10555 (N_10555,N_8844,N_5183);
nand U10556 (N_10556,N_7180,N_9977);
nand U10557 (N_10557,N_9020,N_5471);
and U10558 (N_10558,N_7644,N_5864);
and U10559 (N_10559,N_9273,N_7457);
and U10560 (N_10560,N_6335,N_7290);
xor U10561 (N_10561,N_5816,N_7797);
or U10562 (N_10562,N_8440,N_9586);
and U10563 (N_10563,N_5072,N_8638);
or U10564 (N_10564,N_5382,N_7489);
nor U10565 (N_10565,N_9131,N_9777);
nand U10566 (N_10566,N_7078,N_8703);
nand U10567 (N_10567,N_9767,N_7314);
nor U10568 (N_10568,N_9747,N_8792);
xnor U10569 (N_10569,N_7995,N_9769);
nand U10570 (N_10570,N_6493,N_6223);
or U10571 (N_10571,N_8421,N_9557);
and U10572 (N_10572,N_8354,N_6365);
nand U10573 (N_10573,N_8995,N_6342);
nor U10574 (N_10574,N_8450,N_5447);
nand U10575 (N_10575,N_5915,N_8232);
xnor U10576 (N_10576,N_8185,N_8310);
and U10577 (N_10577,N_9317,N_5861);
nor U10578 (N_10578,N_8757,N_7776);
and U10579 (N_10579,N_5214,N_9930);
or U10580 (N_10580,N_8470,N_6176);
and U10581 (N_10581,N_8039,N_6448);
or U10582 (N_10582,N_7536,N_8581);
nor U10583 (N_10583,N_8032,N_7173);
and U10584 (N_10584,N_5372,N_6642);
nand U10585 (N_10585,N_5583,N_9297);
or U10586 (N_10586,N_5098,N_5667);
nor U10587 (N_10587,N_5683,N_8945);
nand U10588 (N_10588,N_6781,N_6240);
nand U10589 (N_10589,N_5238,N_6962);
nand U10590 (N_10590,N_7300,N_6197);
nor U10591 (N_10591,N_5829,N_7430);
and U10592 (N_10592,N_7548,N_9913);
and U10593 (N_10593,N_8700,N_6793);
or U10594 (N_10594,N_9639,N_8223);
nor U10595 (N_10595,N_8037,N_6523);
nand U10596 (N_10596,N_7011,N_8763);
nand U10597 (N_10597,N_5114,N_6719);
and U10598 (N_10598,N_8772,N_6849);
nor U10599 (N_10599,N_6264,N_5439);
or U10600 (N_10600,N_6346,N_9965);
nand U10601 (N_10601,N_9321,N_8789);
and U10602 (N_10602,N_7091,N_8895);
nor U10603 (N_10603,N_5489,N_9696);
or U10604 (N_10604,N_8390,N_8100);
nand U10605 (N_10605,N_7558,N_5985);
nand U10606 (N_10606,N_9218,N_5982);
or U10607 (N_10607,N_6585,N_9520);
nand U10608 (N_10608,N_9987,N_9754);
nor U10609 (N_10609,N_8388,N_8682);
and U10610 (N_10610,N_9258,N_9607);
nand U10611 (N_10611,N_9164,N_6338);
nor U10612 (N_10612,N_8420,N_5280);
or U10613 (N_10613,N_7888,N_7678);
or U10614 (N_10614,N_7654,N_7685);
xor U10615 (N_10615,N_7474,N_9809);
xnor U10616 (N_10616,N_5043,N_6588);
nand U10617 (N_10617,N_6470,N_7621);
nor U10618 (N_10618,N_7149,N_5576);
and U10619 (N_10619,N_8233,N_8055);
nand U10620 (N_10620,N_7700,N_6208);
nand U10621 (N_10621,N_8525,N_8157);
and U10622 (N_10622,N_6792,N_7202);
nor U10623 (N_10623,N_9061,N_8027);
xor U10624 (N_10624,N_8117,N_8288);
nor U10625 (N_10625,N_8996,N_7082);
and U10626 (N_10626,N_6616,N_7096);
nor U10627 (N_10627,N_8964,N_8997);
and U10628 (N_10628,N_8677,N_8911);
and U10629 (N_10629,N_6724,N_5051);
or U10630 (N_10630,N_7540,N_7681);
and U10631 (N_10631,N_5337,N_6123);
and U10632 (N_10632,N_7379,N_6113);
or U10633 (N_10633,N_5658,N_7116);
nand U10634 (N_10634,N_7265,N_6230);
and U10635 (N_10635,N_7662,N_5185);
nor U10636 (N_10636,N_6658,N_9339);
nor U10637 (N_10637,N_5544,N_9116);
xor U10638 (N_10638,N_8512,N_6510);
and U10639 (N_10639,N_5400,N_7660);
xor U10640 (N_10640,N_8940,N_9980);
nand U10641 (N_10641,N_8540,N_5018);
xor U10642 (N_10642,N_8080,N_7240);
nand U10643 (N_10643,N_8652,N_9772);
nand U10644 (N_10644,N_7517,N_9789);
xor U10645 (N_10645,N_7230,N_6457);
nand U10646 (N_10646,N_6621,N_5701);
or U10647 (N_10647,N_6091,N_8198);
or U10648 (N_10648,N_7860,N_6200);
nor U10649 (N_10649,N_7858,N_7086);
nor U10650 (N_10650,N_6682,N_9156);
and U10651 (N_10651,N_5153,N_6891);
nor U10652 (N_10652,N_6386,N_5716);
and U10653 (N_10653,N_9955,N_8771);
or U10654 (N_10654,N_6101,N_5141);
nand U10655 (N_10655,N_8880,N_8868);
nand U10656 (N_10656,N_5216,N_7331);
xor U10657 (N_10657,N_5618,N_8740);
nand U10658 (N_10658,N_5674,N_8901);
xnor U10659 (N_10659,N_7997,N_6729);
nor U10660 (N_10660,N_7427,N_7750);
nand U10661 (N_10661,N_5994,N_7454);
nor U10662 (N_10662,N_7940,N_5633);
or U10663 (N_10663,N_6038,N_8395);
nor U10664 (N_10664,N_9615,N_8007);
or U10665 (N_10665,N_9206,N_9034);
or U10666 (N_10666,N_6351,N_7605);
or U10667 (N_10667,N_9637,N_7244);
nand U10668 (N_10668,N_8300,N_8385);
or U10669 (N_10669,N_9449,N_6217);
nor U10670 (N_10670,N_8941,N_9669);
or U10671 (N_10671,N_9269,N_7372);
or U10672 (N_10672,N_9177,N_8203);
nand U10673 (N_10673,N_5881,N_8838);
nand U10674 (N_10674,N_5907,N_5953);
and U10675 (N_10675,N_5240,N_7123);
nor U10676 (N_10676,N_7874,N_6426);
nor U10677 (N_10677,N_6736,N_6192);
nor U10678 (N_10678,N_7777,N_5898);
or U10679 (N_10679,N_5748,N_5422);
or U10680 (N_10680,N_8177,N_7458);
or U10681 (N_10681,N_6071,N_7348);
or U10682 (N_10682,N_8051,N_8704);
or U10683 (N_10683,N_7025,N_5720);
and U10684 (N_10684,N_5523,N_8137);
and U10685 (N_10685,N_7090,N_5800);
nor U10686 (N_10686,N_8825,N_9712);
or U10687 (N_10687,N_9327,N_9049);
nand U10688 (N_10688,N_8946,N_5798);
and U10689 (N_10689,N_5619,N_5807);
nand U10690 (N_10690,N_6257,N_9268);
or U10691 (N_10691,N_5636,N_5693);
nand U10692 (N_10692,N_9422,N_9667);
or U10693 (N_10693,N_8266,N_7030);
xor U10694 (N_10694,N_8176,N_9243);
nor U10695 (N_10695,N_5680,N_5858);
and U10696 (N_10696,N_9212,N_9606);
nand U10697 (N_10697,N_6134,N_6237);
and U10698 (N_10698,N_8443,N_6355);
nor U10699 (N_10699,N_8026,N_6362);
and U10700 (N_10700,N_6506,N_9978);
nand U10701 (N_10701,N_5430,N_5386);
nor U10702 (N_10702,N_8229,N_8626);
nand U10703 (N_10703,N_9648,N_9279);
nor U10704 (N_10704,N_8912,N_6884);
nand U10705 (N_10705,N_9163,N_8754);
nor U10706 (N_10706,N_5200,N_9979);
and U10707 (N_10707,N_5521,N_9505);
xor U10708 (N_10708,N_9159,N_6265);
nor U10709 (N_10709,N_8637,N_5377);
and U10710 (N_10710,N_6917,N_6476);
or U10711 (N_10711,N_6098,N_7665);
nor U10712 (N_10712,N_6643,N_8494);
or U10713 (N_10713,N_9024,N_6830);
nor U10714 (N_10714,N_8323,N_5389);
nand U10715 (N_10715,N_8342,N_5446);
or U10716 (N_10716,N_6286,N_8664);
xnor U10717 (N_10717,N_8245,N_8888);
or U10718 (N_10718,N_9407,N_9182);
or U10719 (N_10719,N_5983,N_8641);
or U10720 (N_10720,N_5110,N_6568);
and U10721 (N_10721,N_5852,N_6483);
nor U10722 (N_10722,N_5202,N_8116);
xnor U10723 (N_10723,N_9522,N_8200);
nand U10724 (N_10724,N_9333,N_6720);
nor U10725 (N_10725,N_8264,N_8131);
and U10726 (N_10726,N_8829,N_7064);
and U10727 (N_10727,N_5391,N_9068);
nand U10728 (N_10728,N_9564,N_5569);
nand U10729 (N_10729,N_9393,N_9179);
xor U10730 (N_10730,N_5350,N_5115);
nand U10731 (N_10731,N_9779,N_8668);
or U10732 (N_10732,N_8003,N_8949);
and U10733 (N_10733,N_6382,N_6021);
or U10734 (N_10734,N_6051,N_9512);
and U10735 (N_10735,N_8725,N_9959);
xor U10736 (N_10736,N_5312,N_8862);
and U10737 (N_10737,N_5681,N_9352);
nor U10738 (N_10738,N_9680,N_9823);
or U10739 (N_10739,N_7118,N_5929);
or U10740 (N_10740,N_9483,N_9682);
or U10741 (N_10741,N_5764,N_8811);
and U10742 (N_10742,N_5092,N_5811);
or U10743 (N_10743,N_6140,N_8720);
or U10744 (N_10744,N_7147,N_9887);
nor U10745 (N_10745,N_7908,N_8507);
nand U10746 (N_10746,N_7663,N_5696);
nor U10747 (N_10747,N_7511,N_8490);
or U10748 (N_10748,N_7647,N_5755);
nand U10749 (N_10749,N_5425,N_7145);
nand U10750 (N_10750,N_6974,N_5972);
nor U10751 (N_10751,N_5036,N_7069);
or U10752 (N_10752,N_9175,N_9882);
and U10753 (N_10753,N_9039,N_6554);
or U10754 (N_10754,N_7065,N_6337);
nor U10755 (N_10755,N_7734,N_7033);
or U10756 (N_10756,N_6608,N_8316);
and U10757 (N_10757,N_9850,N_8403);
xor U10758 (N_10758,N_9314,N_8898);
or U10759 (N_10759,N_5482,N_7378);
or U10760 (N_10760,N_5944,N_9717);
and U10761 (N_10761,N_6154,N_8710);
and U10762 (N_10762,N_9381,N_8489);
xor U10763 (N_10763,N_9765,N_7218);
nor U10764 (N_10764,N_5418,N_6306);
nand U10765 (N_10765,N_5575,N_7736);
nand U10766 (N_10766,N_6291,N_5932);
or U10767 (N_10767,N_7505,N_7738);
nand U10768 (N_10768,N_5432,N_5657);
and U10769 (N_10769,N_9154,N_8952);
or U10770 (N_10770,N_9599,N_8736);
nand U10771 (N_10771,N_5596,N_7146);
and U10772 (N_10772,N_9627,N_9137);
and U10773 (N_10773,N_9626,N_7407);
nand U10774 (N_10774,N_6600,N_7313);
nand U10775 (N_10775,N_6789,N_6213);
or U10776 (N_10776,N_6387,N_9860);
or U10777 (N_10777,N_6749,N_7980);
and U10778 (N_10778,N_5242,N_6499);
and U10779 (N_10779,N_9935,N_8362);
nand U10780 (N_10780,N_9525,N_6103);
or U10781 (N_10781,N_9117,N_5704);
nor U10782 (N_10782,N_5947,N_7968);
or U10783 (N_10783,N_8120,N_9191);
nor U10784 (N_10784,N_6619,N_9255);
or U10785 (N_10785,N_5784,N_8761);
and U10786 (N_10786,N_9291,N_6168);
nand U10787 (N_10787,N_7223,N_6683);
nand U10788 (N_10788,N_7506,N_8908);
and U10789 (N_10789,N_6529,N_6475);
or U10790 (N_10790,N_5218,N_6777);
and U10791 (N_10791,N_9706,N_5977);
nand U10792 (N_10792,N_5084,N_6977);
or U10793 (N_10793,N_6082,N_9799);
or U10794 (N_10794,N_9881,N_5771);
nor U10795 (N_10795,N_5221,N_5862);
or U10796 (N_10796,N_9011,N_8675);
or U10797 (N_10797,N_9723,N_7277);
nand U10798 (N_10798,N_6019,N_8146);
or U10799 (N_10799,N_5629,N_8666);
or U10800 (N_10800,N_8277,N_8142);
nand U10801 (N_10801,N_7893,N_6162);
and U10802 (N_10802,N_7371,N_9109);
or U10803 (N_10803,N_5962,N_8410);
and U10804 (N_10804,N_8089,N_9551);
or U10805 (N_10805,N_6520,N_9524);
and U10806 (N_10806,N_7863,N_6245);
and U10807 (N_10807,N_5805,N_8069);
and U10808 (N_10808,N_7054,N_9994);
nor U10809 (N_10809,N_5030,N_5080);
and U10810 (N_10810,N_7826,N_9385);
or U10811 (N_10811,N_5167,N_6442);
nor U10812 (N_10812,N_6853,N_9108);
or U10813 (N_10813,N_8884,N_7514);
nand U10814 (N_10814,N_8587,N_5478);
nor U10815 (N_10815,N_6009,N_9618);
and U10816 (N_10816,N_9331,N_5339);
and U10817 (N_10817,N_5127,N_6206);
or U10818 (N_10818,N_8128,N_9988);
or U10819 (N_10819,N_5699,N_7560);
nand U10820 (N_10820,N_6220,N_8061);
and U10821 (N_10821,N_6108,N_6046);
or U10822 (N_10822,N_8047,N_6077);
xor U10823 (N_10823,N_8516,N_9813);
xor U10824 (N_10824,N_6629,N_9563);
nor U10825 (N_10825,N_9748,N_7198);
nand U10826 (N_10826,N_6723,N_6923);
xor U10827 (N_10827,N_5644,N_9795);
or U10828 (N_10828,N_7852,N_6478);
nand U10829 (N_10829,N_5076,N_8746);
and U10830 (N_10830,N_5360,N_8688);
nand U10831 (N_10831,N_9012,N_6652);
nor U10832 (N_10832,N_8673,N_8568);
nor U10833 (N_10833,N_9610,N_9065);
and U10834 (N_10834,N_9201,N_5847);
nand U10835 (N_10835,N_7886,N_6002);
and U10836 (N_10836,N_8481,N_5754);
nor U10837 (N_10837,N_9262,N_7821);
or U10838 (N_10838,N_7018,N_7258);
or U10839 (N_10839,N_6207,N_5333);
and U10840 (N_10840,N_6525,N_7211);
or U10841 (N_10841,N_5233,N_5669);
and U10842 (N_10842,N_8716,N_7148);
and U10843 (N_10843,N_9105,N_8553);
nor U10844 (N_10844,N_9914,N_7073);
or U10845 (N_10845,N_5165,N_5465);
nand U10846 (N_10846,N_6601,N_8234);
nor U10847 (N_10847,N_9516,N_8983);
nor U10848 (N_10848,N_6366,N_5866);
nand U10849 (N_10849,N_7960,N_7779);
nand U10850 (N_10850,N_9138,N_6214);
and U10851 (N_10851,N_8193,N_9560);
nand U10852 (N_10852,N_9502,N_8526);
or U10853 (N_10853,N_7668,N_9387);
nand U10854 (N_10854,N_6512,N_6314);
or U10855 (N_10855,N_9176,N_5688);
or U10856 (N_10856,N_6255,N_6186);
nor U10857 (N_10857,N_9543,N_5082);
nand U10858 (N_10858,N_5219,N_5821);
and U10859 (N_10859,N_6463,N_5589);
nor U10860 (N_10860,N_9456,N_7203);
nor U10861 (N_10861,N_7959,N_6419);
and U10862 (N_10862,N_6912,N_8405);
or U10863 (N_10863,N_6534,N_5450);
or U10864 (N_10864,N_7093,N_5853);
or U10865 (N_10865,N_5598,N_6906);
or U10866 (N_10866,N_8965,N_5969);
or U10867 (N_10867,N_8423,N_5010);
and U10868 (N_10868,N_5016,N_7594);
or U10869 (N_10869,N_9025,N_5960);
nand U10870 (N_10870,N_9383,N_7875);
and U10871 (N_10871,N_5181,N_9974);
and U10872 (N_10872,N_8418,N_5516);
nand U10873 (N_10873,N_7424,N_5873);
nand U10874 (N_10874,N_5407,N_6023);
nor U10875 (N_10875,N_7855,N_8943);
nand U10876 (N_10876,N_8152,N_8221);
nor U10877 (N_10877,N_8302,N_8551);
nand U10878 (N_10878,N_8926,N_5461);
nand U10879 (N_10879,N_8024,N_5578);
nand U10880 (N_10880,N_7949,N_5235);
nor U10881 (N_10881,N_5517,N_7075);
nor U10882 (N_10882,N_6675,N_8615);
nor U10883 (N_10883,N_7267,N_6648);
or U10884 (N_10884,N_6196,N_7865);
nor U10885 (N_10885,N_8474,N_6256);
nand U10886 (N_10886,N_9829,N_9250);
and U10887 (N_10887,N_8956,N_8309);
nand U10888 (N_10888,N_5332,N_6711);
and U10889 (N_10889,N_7985,N_7017);
nor U10890 (N_10890,N_8847,N_6740);
nand U10891 (N_10891,N_6531,N_6980);
nand U10892 (N_10892,N_7535,N_5289);
nor U10893 (N_10893,N_6638,N_5091);
nand U10894 (N_10894,N_7394,N_6938);
or U10895 (N_10895,N_6440,N_8283);
nand U10896 (N_10896,N_6425,N_9677);
or U10897 (N_10897,N_7844,N_5135);
nand U10898 (N_10898,N_7753,N_9041);
nand U10899 (N_10899,N_7022,N_6831);
or U10900 (N_10900,N_5385,N_5968);
nor U10901 (N_10901,N_7970,N_5419);
nand U10902 (N_10902,N_6418,N_7224);
and U10903 (N_10903,N_6553,N_8905);
and U10904 (N_10904,N_5336,N_9632);
and U10905 (N_10905,N_5319,N_9157);
nand U10906 (N_10906,N_5294,N_6247);
and U10907 (N_10907,N_7910,N_8282);
or U10908 (N_10908,N_6210,N_7016);
nor U10909 (N_10909,N_7083,N_5119);
nand U10910 (N_10910,N_9150,N_7225);
nand U10911 (N_10911,N_6075,N_9675);
nand U10912 (N_10912,N_8633,N_8313);
or U10913 (N_10913,N_8062,N_8826);
nor U10914 (N_10914,N_9244,N_8477);
nor U10915 (N_10915,N_8091,N_5955);
or U10916 (N_10916,N_8890,N_9325);
nand U10917 (N_10917,N_8706,N_6967);
or U10918 (N_10918,N_9556,N_7186);
nand U10919 (N_10919,N_5290,N_5288);
nor U10920 (N_10920,N_7305,N_6467);
nor U10921 (N_10921,N_5528,N_5911);
and U10922 (N_10922,N_7510,N_9685);
nand U10923 (N_10923,N_8671,N_5621);
nor U10924 (N_10924,N_7176,N_5691);
nor U10925 (N_10925,N_8435,N_5408);
or U10926 (N_10926,N_7954,N_9252);
or U10927 (N_10927,N_7095,N_5817);
nand U10928 (N_10928,N_5412,N_8268);
nor U10929 (N_10929,N_9438,N_5959);
and U10930 (N_10930,N_6823,N_7248);
nand U10931 (N_10931,N_6659,N_6164);
nor U10932 (N_10932,N_8758,N_5803);
xnor U10933 (N_10933,N_5571,N_6637);
and U10934 (N_10934,N_8656,N_5320);
and U10935 (N_10935,N_9507,N_7401);
and U10936 (N_10936,N_9369,N_8436);
xnor U10937 (N_10937,N_6438,N_6978);
nor U10938 (N_10938,N_5946,N_8658);
nand U10939 (N_10939,N_8723,N_7912);
or U10940 (N_10940,N_8119,N_6909);
and U10941 (N_10941,N_9037,N_5549);
nor U10942 (N_10942,N_6579,N_7553);
or U10943 (N_10943,N_5826,N_7250);
nor U10944 (N_10944,N_7652,N_5211);
and U10945 (N_10945,N_9391,N_5786);
nand U10946 (N_10946,N_6287,N_9596);
nor U10947 (N_10947,N_9075,N_6956);
or U10948 (N_10948,N_9488,N_7988);
or U10949 (N_10949,N_7101,N_8462);
or U10950 (N_10950,N_6145,N_7629);
and U10951 (N_10951,N_7429,N_5638);
and U10952 (N_10952,N_7050,N_8265);
nand U10953 (N_10953,N_6721,N_6025);
or U10954 (N_10954,N_8284,N_9023);
xor U10955 (N_10955,N_5537,N_8341);
nor U10956 (N_10956,N_9842,N_6045);
nor U10957 (N_10957,N_9686,N_8980);
or U10958 (N_10958,N_8365,N_9873);
nor U10959 (N_10959,N_7964,N_9332);
and U10960 (N_10960,N_5744,N_9737);
nand U10961 (N_10961,N_5775,N_9083);
or U10962 (N_10962,N_8138,N_9288);
or U10963 (N_10963,N_9328,N_9114);
nor U10964 (N_10964,N_5910,N_8126);
or U10965 (N_10965,N_8207,N_9811);
nor U10966 (N_10966,N_8554,N_6411);
xor U10967 (N_10967,N_7013,N_9466);
nor U10968 (N_10968,N_8998,N_8121);
nor U10969 (N_10969,N_9248,N_5580);
or U10970 (N_10970,N_7673,N_6388);
and U10971 (N_10971,N_8552,N_6693);
nand U10972 (N_10972,N_8513,N_5778);
and U10973 (N_10973,N_9202,N_8303);
nand U10974 (N_10974,N_7561,N_9411);
nor U10975 (N_10975,N_8752,N_8645);
nor U10976 (N_10976,N_8182,N_9638);
or U10977 (N_10977,N_6273,N_5259);
and U10978 (N_10978,N_7502,N_9337);
nor U10979 (N_10979,N_5846,N_9408);
nor U10980 (N_10980,N_6827,N_7184);
nor U10981 (N_10981,N_8896,N_8511);
and U10982 (N_10982,N_6178,N_6044);
nor U10983 (N_10983,N_6167,N_9178);
nor U10984 (N_10984,N_9569,N_7229);
or U10985 (N_10985,N_7816,N_9816);
nor U10986 (N_10986,N_6067,N_7288);
nor U10987 (N_10987,N_5958,N_5193);
or U10988 (N_10988,N_8589,N_6985);
or U10989 (N_10989,N_6960,N_6352);
nor U10990 (N_10990,N_5307,N_6479);
nand U10991 (N_10991,N_8378,N_6919);
and U10992 (N_10992,N_9665,N_9630);
nor U10993 (N_10993,N_7885,N_5239);
nor U10994 (N_10994,N_6785,N_8506);
and U10995 (N_10995,N_6580,N_9465);
and U10996 (N_10996,N_8935,N_6869);
xnor U10997 (N_10997,N_7872,N_7696);
nand U10998 (N_10998,N_5366,N_6092);
nor U10999 (N_10999,N_7448,N_8079);
nor U11000 (N_11000,N_7898,N_7614);
nor U11001 (N_11001,N_8159,N_5702);
or U11002 (N_11002,N_8776,N_8981);
nor U11003 (N_11003,N_7293,N_5488);
and U11004 (N_11004,N_5927,N_9129);
nor U11005 (N_11005,N_5496,N_6959);
or U11006 (N_11006,N_8602,N_7469);
or U11007 (N_11007,N_5514,N_5059);
nand U11008 (N_11008,N_6069,N_9284);
nor U11009 (N_11009,N_8843,N_5392);
nor U11010 (N_11010,N_7321,N_9835);
nand U11011 (N_11011,N_7549,N_5318);
xor U11012 (N_11012,N_7911,N_6500);
nor U11013 (N_11013,N_5049,N_5402);
and U11014 (N_11014,N_9441,N_7642);
and U11015 (N_11015,N_8469,N_6243);
nand U11016 (N_11016,N_7979,N_6864);
nand U11017 (N_11017,N_9574,N_5364);
nor U11018 (N_11018,N_5887,N_5175);
nor U11019 (N_11019,N_7178,N_5705);
or U11020 (N_11020,N_9810,N_8643);
nor U11021 (N_11021,N_5512,N_5313);
xnor U11022 (N_11022,N_9207,N_9845);
nand U11023 (N_11023,N_9319,N_8555);
or U11024 (N_11024,N_9732,N_8879);
nor U11025 (N_11025,N_7933,N_5315);
nand U11026 (N_11026,N_7162,N_9919);
xnor U11027 (N_11027,N_6189,N_7946);
or U11028 (N_11028,N_5573,N_6036);
and U11029 (N_11029,N_9259,N_6260);
or U11030 (N_11030,N_5226,N_9047);
and U11031 (N_11031,N_9186,N_9278);
nor U11032 (N_11032,N_5083,N_9568);
or U11033 (N_11033,N_5813,N_6361);
nor U11034 (N_11034,N_8580,N_8528);
nand U11035 (N_11035,N_5995,N_8330);
nor U11036 (N_11036,N_9067,N_7487);
nor U11037 (N_11037,N_6944,N_6191);
and U11038 (N_11038,N_7741,N_9893);
nor U11039 (N_11039,N_7383,N_5836);
nand U11040 (N_11040,N_7939,N_7432);
nand U11041 (N_11041,N_7092,N_6157);
or U11042 (N_11042,N_6252,N_5225);
nand U11043 (N_11043,N_6515,N_6603);
or U11044 (N_11044,N_7847,N_6908);
nand U11045 (N_11045,N_6569,N_8530);
and U11046 (N_11046,N_5201,N_9360);
xnor U11047 (N_11047,N_5642,N_5513);
or U11048 (N_11048,N_5093,N_8259);
or U11049 (N_11049,N_8854,N_8478);
nor U11050 (N_11050,N_6378,N_6498);
and U11051 (N_11051,N_6874,N_5468);
nand U11052 (N_11052,N_9942,N_8433);
nand U11053 (N_11053,N_6267,N_8086);
nor U11054 (N_11054,N_7052,N_5000);
and U11055 (N_11055,N_6422,N_8446);
nor U11056 (N_11056,N_5870,N_8098);
nor U11057 (N_11057,N_8906,N_8593);
nand U11058 (N_11058,N_7972,N_8665);
and U11059 (N_11059,N_9936,N_6668);
and U11060 (N_11060,N_9776,N_6161);
nor U11061 (N_11061,N_8369,N_5254);
nor U11062 (N_11062,N_6929,N_6622);
nor U11063 (N_11063,N_5627,N_9007);
or U11064 (N_11064,N_8842,N_6611);
nand U11065 (N_11065,N_9721,N_6329);
and U11066 (N_11066,N_6872,N_5013);
nor U11067 (N_11067,N_7557,N_5799);
nor U11068 (N_11068,N_7268,N_7406);
nand U11069 (N_11069,N_9838,N_8779);
and U11070 (N_11070,N_5675,N_6070);
and U11071 (N_11071,N_5808,N_9057);
or U11072 (N_11072,N_8948,N_7716);
nor U11073 (N_11073,N_6084,N_8247);
and U11074 (N_11074,N_5399,N_9857);
nand U11075 (N_11075,N_9498,N_7131);
nor U11076 (N_11076,N_6598,N_7486);
and U11077 (N_11077,N_5845,N_6973);
and U11078 (N_11078,N_9820,N_5746);
nand U11079 (N_11079,N_9926,N_6492);
nor U11080 (N_11080,N_8984,N_7056);
xor U11081 (N_11081,N_6770,N_8398);
nand U11082 (N_11082,N_9964,N_9727);
xor U11083 (N_11083,N_9092,N_5037);
or U11084 (N_11084,N_6008,N_9313);
or U11085 (N_11085,N_6004,N_7729);
nor U11086 (N_11086,N_5404,N_8914);
or U11087 (N_11087,N_5666,N_8828);
nand U11088 (N_11088,N_5148,N_9734);
nor U11089 (N_11089,N_8179,N_6905);
or U11090 (N_11090,N_6397,N_9888);
or U11091 (N_11091,N_7251,N_8105);
nor U11092 (N_11092,N_9085,N_5456);
and U11093 (N_11093,N_5922,N_6163);
xor U11094 (N_11094,N_5264,N_8337);
nand U11095 (N_11095,N_6641,N_5352);
and U11096 (N_11096,N_8340,N_6495);
and U11097 (N_11097,N_6065,N_8876);
nand U11098 (N_11098,N_7285,N_5867);
nand U11099 (N_11099,N_6089,N_6481);
nand U11100 (N_11100,N_9277,N_7920);
nor U11101 (N_11101,N_9804,N_6311);
nand U11102 (N_11102,N_8424,N_8181);
xnor U11103 (N_11103,N_7830,N_9084);
nor U11104 (N_11104,N_5526,N_5857);
xor U11105 (N_11105,N_8289,N_7252);
and U11106 (N_11106,N_9825,N_8647);
nand U11107 (N_11107,N_8246,N_6446);
xnor U11108 (N_11108,N_9553,N_5173);
or U11109 (N_11109,N_5487,N_5314);
and U11110 (N_11110,N_9528,N_7077);
xor U11111 (N_11111,N_8280,N_7613);
and U11112 (N_11112,N_7573,N_9997);
or U11113 (N_11113,N_8517,N_7438);
xnor U11114 (N_11114,N_8239,N_8466);
nor U11115 (N_11115,N_7374,N_6727);
nand U11116 (N_11116,N_7881,N_7541);
or U11117 (N_11117,N_5033,N_8413);
nor U11118 (N_11118,N_8106,N_9299);
and U11119 (N_11119,N_7171,N_5396);
and U11120 (N_11120,N_8379,N_8667);
nand U11121 (N_11121,N_5435,N_7627);
nand U11122 (N_11122,N_5089,N_7496);
nand U11123 (N_11123,N_6058,N_5601);
nor U11124 (N_11124,N_9578,N_9948);
and U11125 (N_11125,N_5828,N_6540);
nor U11126 (N_11126,N_6341,N_6453);
nand U11127 (N_11127,N_5373,N_6896);
xnor U11128 (N_11128,N_9871,N_8359);
nor U11129 (N_11129,N_8441,N_8713);
or U11130 (N_11130,N_6332,N_8885);
and U11131 (N_11131,N_7991,N_5801);
nand U11132 (N_11132,N_9365,N_5820);
and U11133 (N_11133,N_8204,N_6826);
nand U11134 (N_11134,N_8750,N_8150);
nand U11135 (N_11135,N_9461,N_7004);
or U11136 (N_11136,N_5176,N_9070);
or U11137 (N_11137,N_8113,N_5649);
nand U11138 (N_11138,N_7828,N_9697);
or U11139 (N_11139,N_5780,N_6539);
or U11140 (N_11140,N_9879,N_8361);
and U11141 (N_11141,N_7924,N_6801);
nand U11142 (N_11142,N_7404,N_6583);
and U11143 (N_11143,N_9593,N_6227);
or U11144 (N_11144,N_8539,N_9812);
nand U11145 (N_11145,N_8351,N_6219);
xor U11146 (N_11146,N_5728,N_8006);
nor U11147 (N_11147,N_5331,N_6431);
nor U11148 (N_11148,N_9435,N_9794);
nor U11149 (N_11149,N_6632,N_6490);
nor U11150 (N_11150,N_7276,N_9937);
nand U11151 (N_11151,N_9402,N_7569);
nor U11152 (N_11152,N_6013,N_8078);
nand U11153 (N_11153,N_7601,N_6590);
and U11154 (N_11154,N_9654,N_7664);
and U11155 (N_11155,N_8686,N_8502);
nor U11156 (N_11156,N_7866,N_6788);
nor U11157 (N_11157,N_7529,N_8640);
or U11158 (N_11158,N_6151,N_8194);
or U11159 (N_11159,N_7396,N_5709);
and U11160 (N_11160,N_8764,N_6509);
xnor U11161 (N_11161,N_7410,N_5729);
xnor U11162 (N_11162,N_8160,N_6456);
or U11163 (N_11163,N_7854,N_7698);
nand U11164 (N_11164,N_7503,N_9249);
nand U11165 (N_11165,N_9999,N_6072);
nor U11166 (N_11166,N_5002,N_5476);
or U11167 (N_11167,N_9781,N_5690);
nor U11168 (N_11168,N_9464,N_5246);
nor U11169 (N_11169,N_8020,N_6258);
or U11170 (N_11170,N_9705,N_7309);
nand U11171 (N_11171,N_6970,N_8399);
and U11172 (N_11172,N_7163,N_5329);
xor U11173 (N_11173,N_9631,N_6039);
nand U11174 (N_11174,N_5023,N_6399);
or U11175 (N_11175,N_7590,N_7791);
nand U11176 (N_11176,N_9286,N_8930);
nor U11177 (N_11177,N_7579,N_5546);
nor U11178 (N_11178,N_9013,N_7455);
nand U11179 (N_11179,N_5261,N_8910);
or U11180 (N_11180,N_6745,N_9232);
nand U11181 (N_11181,N_6224,N_8196);
or U11182 (N_11182,N_7026,N_9355);
nand U11183 (N_11183,N_8454,N_8515);
nor U11184 (N_11184,N_8471,N_5912);
nand U11185 (N_11185,N_5493,N_6360);
nor U11186 (N_11186,N_9242,N_9718);
xor U11187 (N_11187,N_9847,N_9471);
nor U11188 (N_11188,N_6859,N_8760);
nand U11189 (N_11189,N_6800,N_8805);
or U11190 (N_11190,N_7546,N_7719);
or U11191 (N_11191,N_5145,N_8397);
or U11192 (N_11192,N_8005,N_8709);
nor U11193 (N_11193,N_7156,N_9431);
or U11194 (N_11194,N_8011,N_7326);
or U11195 (N_11195,N_8273,N_6895);
or U11196 (N_11196,N_6686,N_6466);
nand U11197 (N_11197,N_7822,N_6860);
nand U11198 (N_11198,N_7155,N_8201);
nand U11199 (N_11199,N_8251,N_9312);
or U11200 (N_11200,N_9907,N_9868);
nand U11201 (N_11201,N_8676,N_5557);
nor U11202 (N_11202,N_6180,N_9973);
nor U11203 (N_11203,N_8415,N_7209);
nor U11204 (N_11204,N_9591,N_5603);
nor U11205 (N_11205,N_8013,N_8670);
and U11206 (N_11206,N_7508,N_9662);
nand U11207 (N_11207,N_6808,N_7834);
nor U11208 (N_11208,N_5742,N_5198);
nor U11209 (N_11209,N_8068,N_5126);
nor U11210 (N_11210,N_7755,N_7127);
nor U11211 (N_11211,N_7170,N_7032);
nor U11212 (N_11212,N_7574,N_8111);
or U11213 (N_11213,N_8822,N_9646);
or U11214 (N_11214,N_7637,N_9830);
and U11215 (N_11215,N_6292,N_9110);
and U11216 (N_11216,N_6301,N_6472);
nand U11217 (N_11217,N_8722,N_7389);
and U11218 (N_11218,N_8978,N_5706);
xnor U11219 (N_11219,N_6185,N_9694);
and U11220 (N_11220,N_5265,N_5804);
nand U11221 (N_11221,N_6976,N_8325);
xor U11222 (N_11222,N_9859,N_8684);
or U11223 (N_11223,N_8889,N_8659);
nand U11224 (N_11224,N_5305,N_8872);
or U11225 (N_11225,N_9602,N_7068);
nand U11226 (N_11226,N_6548,N_5556);
nand U11227 (N_11227,N_7094,N_7387);
nand U11228 (N_11228,N_6402,N_6455);
nand U11229 (N_11229,N_6706,N_6556);
or U11230 (N_11230,N_7317,N_7655);
nand U11231 (N_11231,N_9992,N_9925);
and U11232 (N_11232,N_7666,N_7320);
nand U11233 (N_11233,N_7261,N_8056);
and U11234 (N_11234,N_7183,N_9486);
and U11235 (N_11235,N_9972,N_7730);
nand U11236 (N_11236,N_8972,N_7479);
and U11237 (N_11237,N_8366,N_8428);
nor U11238 (N_11238,N_7053,N_7047);
xor U11239 (N_11239,N_5005,N_9872);
nand U11240 (N_11240,N_6880,N_7070);
nand U11241 (N_11241,N_8238,N_9619);
nor U11242 (N_11242,N_9684,N_7472);
and U11243 (N_11243,N_8730,N_9693);
xnor U11244 (N_11244,N_5768,N_6190);
nand U11245 (N_11245,N_9982,N_5494);
and U11246 (N_11246,N_7271,N_9540);
nor U11247 (N_11247,N_7916,N_5930);
nand U11248 (N_11248,N_9136,N_5438);
or U11249 (N_11249,N_7081,N_9063);
nand U11250 (N_11250,N_8951,N_6551);
and U11251 (N_11251,N_9566,N_5712);
or U11252 (N_11252,N_5763,N_7783);
or U11253 (N_11253,N_5723,N_7670);
nand U11254 (N_11254,N_7045,N_6726);
nor U11255 (N_11255,N_6903,N_8687);
or U11256 (N_11256,N_8783,N_8976);
or U11257 (N_11257,N_6187,N_5752);
and U11258 (N_11258,N_9095,N_5384);
nand U11259 (N_11259,N_8802,N_7948);
and U11260 (N_11260,N_5552,N_6732);
and U11261 (N_11261,N_6841,N_6503);
and U11262 (N_11262,N_5192,N_7619);
nand U11263 (N_11263,N_6969,N_6102);
nor U11264 (N_11264,N_7757,N_7790);
and U11265 (N_11265,N_8777,N_7831);
or U11266 (N_11266,N_8357,N_8021);
nand U11267 (N_11267,N_9052,N_7242);
or U11268 (N_11268,N_8928,N_6465);
nand U11269 (N_11269,N_9265,N_9096);
xor U11270 (N_11270,N_7152,N_7947);
or U11271 (N_11271,N_8742,N_7841);
nor U11272 (N_11272,N_5169,N_7392);
or U11273 (N_11273,N_8498,N_5297);
nor U11274 (N_11274,N_5727,N_5209);
and U11275 (N_11275,N_8275,N_9120);
or U11276 (N_11276,N_7723,N_7393);
or U11277 (N_11277,N_5156,N_8073);
nor U11278 (N_11278,N_9985,N_7936);
nand U11279 (N_11279,N_7720,N_8535);
nor U11280 (N_11280,N_8650,N_6172);
nor U11281 (N_11281,N_9517,N_8363);
or U11282 (N_11282,N_7071,N_9652);
or U11283 (N_11283,N_6317,N_5009);
or U11284 (N_11284,N_8491,N_8600);
nand U11285 (N_11285,N_9719,N_6393);
or U11286 (N_11286,N_9780,N_5187);
nand U11287 (N_11287,N_5558,N_8791);
nor U11288 (N_11288,N_9861,N_5370);
nor U11289 (N_11289,N_5885,N_9885);
or U11290 (N_11290,N_6228,N_9040);
and U11291 (N_11291,N_9134,N_6701);
xor U11292 (N_11292,N_5711,N_9001);
or U11293 (N_11293,N_9554,N_9848);
nand U11294 (N_11294,N_8558,N_5668);
nand U11295 (N_11295,N_7989,N_5203);
xnor U11296 (N_11296,N_6772,N_7690);
nor U11297 (N_11297,N_9308,N_8749);
nand U11298 (N_11298,N_9298,N_6940);
nand U11299 (N_11299,N_9170,N_7459);
and U11300 (N_11300,N_9929,N_9071);
or U11301 (N_11301,N_6205,N_9021);
and U11302 (N_11302,N_5952,N_6883);
nor U11303 (N_11303,N_8919,N_5085);
or U11304 (N_11304,N_5924,N_8125);
nand U11305 (N_11305,N_6315,N_5901);
nor U11306 (N_11306,N_7434,N_7060);
and U11307 (N_11307,N_6290,N_6088);
nor U11308 (N_11308,N_6888,N_9753);
xnor U11309 (N_11309,N_7283,N_6156);
or U11310 (N_11310,N_8961,N_9434);
and U11311 (N_11311,N_6949,N_9983);
nor U11312 (N_11312,N_7932,N_9755);
nor U11313 (N_11313,N_6430,N_8124);
or U11314 (N_11314,N_6390,N_9469);
and U11315 (N_11315,N_8164,N_5361);
or U11316 (N_11316,N_8312,N_5311);
and U11317 (N_11317,N_7688,N_9444);
nand U11318 (N_11318,N_7001,N_5302);
nor U11319 (N_11319,N_8272,N_5368);
nor U11320 (N_11320,N_7704,N_6945);
nor U11321 (N_11321,N_9367,N_7555);
nand U11322 (N_11322,N_6119,N_7718);
nand U11323 (N_11323,N_8747,N_7551);
nor U11324 (N_11324,N_7626,N_6450);
or U11325 (N_11325,N_7915,N_7311);
nand U11326 (N_11326,N_7840,N_6555);
or U11327 (N_11327,N_9161,N_9213);
nor U11328 (N_11328,N_7439,N_6052);
nand U11329 (N_11329,N_5996,N_5566);
and U11330 (N_11330,N_5632,N_8692);
nand U11331 (N_11331,N_7724,N_6613);
or U11332 (N_11332,N_6617,N_7153);
nor U11333 (N_11333,N_7918,N_8015);
nand U11334 (N_11334,N_6429,N_8023);
or U11335 (N_11335,N_6474,N_9490);
and U11336 (N_11336,N_9474,N_8702);
nand U11337 (N_11337,N_5677,N_8564);
or U11338 (N_11338,N_9745,N_6775);
or U11339 (N_11339,N_8852,N_6672);
or U11340 (N_11340,N_8909,N_6685);
nand U11341 (N_11341,N_9340,N_5635);
nand U11342 (N_11342,N_9542,N_8484);
nand U11343 (N_11343,N_9030,N_6597);
nand U11344 (N_11344,N_9174,N_8141);
nand U11345 (N_11345,N_8644,N_8458);
or U11346 (N_11346,N_6696,N_6441);
or U11347 (N_11347,N_5570,N_9335);
or U11348 (N_11348,N_7107,N_9981);
and U11349 (N_11349,N_7492,N_8953);
nor U11350 (N_11350,N_8168,N_6383);
and U11351 (N_11351,N_9890,N_5767);
nand U11352 (N_11352,N_6359,N_7428);
nor U11353 (N_11353,N_6576,N_8840);
or U11354 (N_11354,N_6712,N_7850);
nand U11355 (N_11355,N_5759,N_8696);
nand U11356 (N_11356,N_5118,N_7994);
and U11357 (N_11357,N_9149,N_7993);
nor U11358 (N_11358,N_9768,N_6932);
nand U11359 (N_11359,N_8144,N_8859);
nor U11360 (N_11360,N_8374,N_5876);
nand U11361 (N_11361,N_6527,N_8215);
or U11362 (N_11362,N_8955,N_6582);
nand U11363 (N_11363,N_7571,N_9570);
nor U11364 (N_11364,N_8205,N_7691);
and U11365 (N_11365,N_7168,N_5121);
and U11366 (N_11366,N_9436,N_7182);
or U11367 (N_11367,N_6141,N_6254);
nand U11368 (N_11368,N_5357,N_9005);
nor U11369 (N_11369,N_5581,N_9304);
nor U11370 (N_11370,N_9798,N_5416);
nand U11371 (N_11371,N_9181,N_6060);
or U11372 (N_11372,N_6707,N_5524);
or U11373 (N_11373,N_8402,N_9484);
and U11374 (N_11374,N_9738,N_9351);
or U11375 (N_11375,N_7969,N_9672);
or U11376 (N_11376,N_5490,N_8508);
and U11377 (N_11377,N_7027,N_8353);
nor U11378 (N_11378,N_8162,N_9169);
nand U11379 (N_11379,N_7411,N_6744);
and U11380 (N_11380,N_7682,N_7775);
nor U11381 (N_11381,N_9526,N_6339);
nand U11382 (N_11382,N_8076,N_5848);
nand U11383 (N_11383,N_5733,N_9043);
nand U11384 (N_11384,N_9489,N_8448);
nand U11385 (N_11385,N_9220,N_9139);
nand U11386 (N_11386,N_8765,N_9763);
nand U11387 (N_11387,N_8122,N_8315);
nand U11388 (N_11388,N_7440,N_8518);
xor U11389 (N_11389,N_5096,N_5703);
or U11390 (N_11390,N_6848,N_8449);
and U11391 (N_11391,N_7217,N_9709);
nor U11392 (N_11392,N_7226,N_6304);
nand U11393 (N_11393,N_7693,N_7981);
nand U11394 (N_11394,N_7699,N_8151);
or U11395 (N_11395,N_8169,N_7437);
and U11396 (N_11396,N_5395,N_7680);
nand U11397 (N_11397,N_7711,N_8786);
and U11398 (N_11398,N_7870,N_9572);
nor U11399 (N_11399,N_7593,N_7577);
nor U11400 (N_11400,N_7600,N_7524);
and U11401 (N_11401,N_9657,N_5774);
or U11402 (N_11402,N_9584,N_8900);
or U11403 (N_11403,N_6660,N_6862);
nand U11404 (N_11404,N_9532,N_8857);
and U11405 (N_11405,N_7659,N_7006);
or U11406 (N_11406,N_7122,N_7200);
and U11407 (N_11407,N_9468,N_5262);
nor U11408 (N_11408,N_8311,N_8523);
xor U11409 (N_11409,N_6750,N_7632);
xor U11410 (N_11410,N_6517,N_6175);
or U11411 (N_11411,N_7525,N_7849);
nor U11412 (N_11412,N_6439,N_9749);
nor U11413 (N_11413,N_7282,N_5303);
and U11414 (N_11414,N_9479,N_6165);
nor U11415 (N_11415,N_8338,N_7616);
nor U11416 (N_11416,N_7023,N_8808);
and U11417 (N_11417,N_6514,N_5228);
nor U11418 (N_11418,N_7234,N_8886);
xnor U11419 (N_11419,N_7446,N_5735);
and U11420 (N_11420,N_7130,N_9290);
or U11421 (N_11421,N_9939,N_7306);
xnor U11422 (N_11422,N_5904,N_7318);
or U11423 (N_11423,N_8165,N_9133);
or U11424 (N_11424,N_7868,N_8592);
or U11425 (N_11425,N_8123,N_7669);
nand U11426 (N_11426,N_6879,N_5940);
xor U11427 (N_11427,N_7233,N_8950);
nand U11428 (N_11428,N_7480,N_7640);
and U11429 (N_11429,N_9741,N_5140);
nand U11430 (N_11430,N_7238,N_8519);
nor U11431 (N_11431,N_7904,N_7325);
nand U11432 (N_11432,N_7697,N_7207);
nor U11433 (N_11433,N_6496,N_8453);
or U11434 (N_11434,N_7185,N_7373);
and U11435 (N_11435,N_7193,N_5682);
nand U11436 (N_11436,N_6767,N_5586);
and U11437 (N_11437,N_6835,N_5129);
and U11438 (N_11438,N_5585,N_8591);
and U11439 (N_11439,N_9600,N_8537);
or U11440 (N_11440,N_5321,N_5793);
and U11441 (N_11441,N_6014,N_5736);
and U11442 (N_11442,N_6757,N_5155);
nand U11443 (N_11443,N_7667,N_5789);
and U11444 (N_11444,N_6656,N_9363);
nand U11445 (N_11445,N_7892,N_7247);
nor U11446 (N_11446,N_6458,N_9223);
nand U11447 (N_11447,N_5473,N_9736);
or U11448 (N_11448,N_7089,N_5086);
and U11449 (N_11449,N_6662,N_7771);
nand U11450 (N_11450,N_7809,N_6572);
nand U11451 (N_11451,N_6957,N_5342);
and U11452 (N_11452,N_8988,N_7902);
nor U11453 (N_11453,N_9219,N_5133);
nand U11454 (N_11454,N_5275,N_8661);
and U11455 (N_11455,N_8595,N_8679);
and U11456 (N_11456,N_8377,N_7361);
nor U11457 (N_11457,N_5806,N_7815);
nand U11458 (N_11458,N_8654,N_8074);
or U11459 (N_11459,N_5673,N_9519);
nand U11460 (N_11460,N_6148,N_7035);
and U11461 (N_11461,N_7140,N_5623);
and U11462 (N_11462,N_6999,N_7303);
nor U11463 (N_11463,N_5692,N_9594);
nor U11464 (N_11464,N_7324,N_8406);
nand U11465 (N_11465,N_8090,N_6780);
nor U11466 (N_11466,N_7159,N_7187);
or U11467 (N_11467,N_6100,N_8492);
or U11468 (N_11468,N_7829,N_8331);
or U11469 (N_11469,N_8350,N_6204);
nand U11470 (N_11470,N_6925,N_8058);
xnor U11471 (N_11471,N_9724,N_8163);
and U11472 (N_11472,N_5536,N_9015);
nand U11473 (N_11473,N_6877,N_6852);
or U11474 (N_11474,N_8317,N_7864);
nand U11475 (N_11475,N_6416,N_6389);
nor U11476 (N_11476,N_8262,N_9416);
or U11477 (N_11477,N_6730,N_6943);
nand U11478 (N_11478,N_5931,N_9151);
or U11479 (N_11479,N_5459,N_6677);
or U11480 (N_11480,N_9446,N_7259);
nor U11481 (N_11481,N_7144,N_7132);
nor U11482 (N_11482,N_7610,N_5090);
and U11483 (N_11483,N_8504,N_6028);
or U11484 (N_11484,N_7802,N_9118);
or U11485 (N_11485,N_9633,N_8959);
and U11486 (N_11486,N_6281,N_7901);
nand U11487 (N_11487,N_5679,N_5966);
nor U11488 (N_11488,N_9975,N_6279);
nand U11489 (N_11489,N_5533,N_7559);
nor U11490 (N_11490,N_5249,N_5362);
nand U11491 (N_11491,N_6722,N_8304);
nor U11492 (N_11492,N_6022,N_5324);
nand U11493 (N_11493,N_6673,N_9226);
nand U11494 (N_11494,N_5236,N_7636);
nand U11495 (N_11495,N_8218,N_8127);
nand U11496 (N_11496,N_5123,N_5134);
and U11497 (N_11497,N_5809,N_5111);
nand U11498 (N_11498,N_8257,N_6047);
nand U11499 (N_11499,N_5292,N_6639);
or U11500 (N_11500,N_7566,N_7477);
nand U11501 (N_11501,N_5919,N_9420);
nor U11502 (N_11502,N_6288,N_5470);
nor U11503 (N_11503,N_6334,N_9695);
and U11504 (N_11504,N_8187,N_8790);
nand U11505 (N_11505,N_6787,N_7602);
nor U11506 (N_11506,N_9991,N_5157);
and U11507 (N_11507,N_5172,N_8437);
and U11508 (N_11508,N_5166,N_9399);
nor U11509 (N_11509,N_8565,N_6728);
nor U11510 (N_11510,N_7684,N_7827);
nand U11511 (N_11511,N_8987,N_7445);
and U11512 (N_11512,N_8012,N_8460);
nand U11513 (N_11513,N_8631,N_5525);
or U11514 (N_11514,N_5749,N_9261);
nor U11515 (N_11515,N_7281,N_6502);
and U11516 (N_11516,N_5541,N_5232);
nor U11517 (N_11517,N_9062,N_5563);
nand U11518 (N_11518,N_9806,N_8577);
nand U11519 (N_11519,N_8968,N_6893);
or U11520 (N_11520,N_6114,N_6676);
and U11521 (N_11521,N_6209,N_6226);
and U11522 (N_11522,N_6188,N_5039);
or U11523 (N_11523,N_7817,N_5593);
or U11524 (N_11524,N_9577,N_9896);
nor U11525 (N_11525,N_6782,N_9924);
and U11526 (N_11526,N_9671,N_7336);
nor U11527 (N_11527,N_7172,N_5957);
nand U11528 (N_11528,N_9165,N_5099);
and U11529 (N_11529,N_5822,N_5599);
xor U11530 (N_11530,N_5745,N_8780);
or U11531 (N_11531,N_6725,N_9858);
nand U11532 (N_11532,N_5281,N_7063);
xnor U11533 (N_11533,N_7206,N_7649);
and U11534 (N_11534,N_8932,N_8616);
nand U11535 (N_11535,N_9500,N_9803);
and U11536 (N_11536,N_6913,N_9406);
and U11537 (N_11537,N_9567,N_6394);
nand U11538 (N_11538,N_9194,N_8499);
nor U11539 (N_11539,N_6739,N_5105);
and U11540 (N_11540,N_9323,N_9801);
and U11541 (N_11541,N_8649,N_5605);
nor U11542 (N_11542,N_9869,N_9295);
or U11543 (N_11543,N_7113,N_6144);
xor U11544 (N_11544,N_9649,N_7814);
nor U11545 (N_11545,N_9899,N_8380);
or U11546 (N_11546,N_8586,N_5747);
and U11547 (N_11547,N_5504,N_6270);
nand U11548 (N_11548,N_9863,N_9107);
nand U11549 (N_11549,N_5087,N_9561);
and U11550 (N_11550,N_9623,N_6110);
nand U11551 (N_11551,N_9853,N_8653);
or U11552 (N_11552,N_9529,N_5609);
or U11553 (N_11553,N_7151,N_7848);
and U11554 (N_11554,N_5453,N_9275);
and U11555 (N_11555,N_9032,N_6563);
nor U11556 (N_11556,N_7583,N_5568);
nand U11557 (N_11557,N_6130,N_7572);
and U11558 (N_11558,N_7842,N_5884);
nor U11559 (N_11559,N_5469,N_8830);
and U11560 (N_11560,N_7609,N_6313);
nand U11561 (N_11561,N_6460,N_9060);
or U11562 (N_11562,N_6010,N_9791);
nor U11563 (N_11563,N_9099,N_7624);
nor U11564 (N_11564,N_7990,N_7337);
or U11565 (N_11565,N_6986,N_5954);
nor U11566 (N_11566,N_6343,N_8166);
xor U11567 (N_11567,N_6147,N_5879);
nand U11568 (N_11568,N_9947,N_8050);
nor U11569 (N_11569,N_6832,N_5186);
nor U11570 (N_11570,N_5376,N_5015);
or U11571 (N_11571,N_7425,N_8237);
nor U11572 (N_11572,N_7804,N_7350);
and U11573 (N_11573,N_8184,N_6742);
nor U11574 (N_11574,N_6535,N_8620);
nor U11575 (N_11575,N_9460,N_7108);
nor U11576 (N_11576,N_8809,N_9642);
or U11577 (N_11577,N_8136,N_7513);
nor U11578 (N_11578,N_7953,N_8041);
nand U11579 (N_11579,N_6620,N_8524);
nor U11580 (N_11580,N_7291,N_8944);
nand U11581 (N_11581,N_6713,N_5250);
nand U11582 (N_11582,N_7871,N_5245);
or U11583 (N_11583,N_8831,N_8101);
nor U11584 (N_11584,N_9044,N_7611);
or U11585 (N_11585,N_9494,N_7169);
nor U11586 (N_11586,N_8628,N_8672);
nor U11587 (N_11587,N_7935,N_5761);
or U11588 (N_11588,N_8018,N_8798);
nand U11589 (N_11589,N_5948,N_9698);
or U11590 (N_11590,N_5149,N_7481);
nand U11591 (N_11591,N_8800,N_6375);
nand U11592 (N_11592,N_9774,N_6143);
nand U11593 (N_11593,N_6628,N_9819);
or U11594 (N_11594,N_8993,N_9066);
or U11595 (N_11595,N_6194,N_9773);
and U11596 (N_11596,N_6537,N_6992);
nand U11597 (N_11597,N_5921,N_5534);
nor U11598 (N_11598,N_6391,N_7820);
nand U11599 (N_11599,N_5540,N_8241);
nand U11600 (N_11600,N_6284,N_5003);
and U11601 (N_11601,N_5882,N_5454);
nor U11602 (N_11602,N_7650,N_5012);
or U11603 (N_11603,N_8010,N_9310);
or U11604 (N_11604,N_5762,N_7575);
nor U11605 (N_11605,N_9343,N_6384);
and U11606 (N_11606,N_8958,N_5758);
nand U11607 (N_11607,N_8271,N_9088);
and U11608 (N_11608,N_7595,N_8025);
nand U11609 (N_11609,N_5338,N_5842);
nor U11610 (N_11610,N_8837,N_8756);
nand U11611 (N_11611,N_6955,N_9417);
nor U11612 (N_11612,N_8924,N_9320);
or U11613 (N_11613,N_6412,N_5511);
and U11614 (N_11614,N_7102,N_8907);
or U11615 (N_11615,N_5019,N_9233);
or U11616 (N_11616,N_5650,N_9612);
and U11617 (N_11617,N_7228,N_7512);
nand U11618 (N_11618,N_6630,N_5785);
and U11619 (N_11619,N_9815,N_6484);
and U11620 (N_11620,N_5643,N_5178);
and U11621 (N_11621,N_9086,N_9069);
or U11622 (N_11622,N_5444,N_8475);
and U11623 (N_11623,N_7166,N_5215);
or U11624 (N_11624,N_7241,N_5387);
or U11625 (N_11625,N_9180,N_7062);
and U11626 (N_11626,N_7733,N_7106);
or U11627 (N_11627,N_5403,N_9102);
nand U11628 (N_11628,N_7307,N_9579);
or U11629 (N_11629,N_8070,N_7962);
nand U11630 (N_11630,N_6599,N_8922);
xnor U11631 (N_11631,N_7785,N_9146);
nand U11632 (N_11632,N_8623,N_9448);
or U11633 (N_11633,N_9691,N_7622);
or U11634 (N_11634,N_9984,N_6086);
nand U11635 (N_11635,N_7197,N_8017);
and U11636 (N_11636,N_8985,N_9405);
nand U11637 (N_11637,N_9267,N_6873);
nor U11638 (N_11638,N_5976,N_5886);
and U11639 (N_11639,N_6991,N_9347);
nand U11640 (N_11640,N_9375,N_6661);
nor U11641 (N_11641,N_7031,N_5268);
or U11642 (N_11642,N_6935,N_8180);
and U11643 (N_11643,N_5194,N_7708);
and U11644 (N_11644,N_9418,N_5335);
and U11645 (N_11645,N_9889,N_6710);
xor U11646 (N_11646,N_7539,N_9636);
or U11647 (N_11647,N_5485,N_9715);
and U11648 (N_11648,N_8801,N_7310);
nand U11649 (N_11649,N_8739,N_7580);
nand U11650 (N_11650,N_8533,N_5182);
nor U11651 (N_11651,N_6184,N_7952);
nor U11652 (N_11652,N_5029,N_6820);
and U11653 (N_11653,N_7845,N_9009);
or U11654 (N_11654,N_9189,N_8190);
and U11655 (N_11655,N_7286,N_7485);
nand U11656 (N_11656,N_7562,N_5740);
and U11657 (N_11657,N_9253,N_9766);
and U11658 (N_11658,N_9902,N_8186);
nand U11659 (N_11659,N_9358,N_7079);
or U11660 (N_11660,N_7397,N_9854);
and U11661 (N_11661,N_6170,N_8617);
and U11662 (N_11662,N_8937,N_8849);
nand U11663 (N_11663,N_5564,N_7727);
nor U11664 (N_11664,N_9018,N_6012);
nand U11665 (N_11665,N_6035,N_7782);
and U11666 (N_11666,N_5378,N_6795);
nand U11667 (N_11667,N_7544,N_5917);
or U11668 (N_11668,N_7722,N_9663);
nor U11669 (N_11669,N_9904,N_8548);
and U11670 (N_11670,N_9523,N_9476);
nand U11671 (N_11671,N_6698,N_9808);
nor U11672 (N_11672,N_7360,N_7944);
nand U11673 (N_11673,N_7443,N_9752);
and U11674 (N_11674,N_5455,N_6408);
nand U11675 (N_11675,N_6381,N_6951);
or U11676 (N_11676,N_9707,N_6323);
nand U11677 (N_11677,N_8858,N_6239);
and U11678 (N_11678,N_6587,N_9442);
and U11679 (N_11679,N_7388,N_6836);
or U11680 (N_11680,N_6501,N_8422);
nor U11681 (N_11681,N_5081,N_6099);
xor U11682 (N_11682,N_9100,N_9421);
or U11683 (N_11683,N_8243,N_5132);
nor U11684 (N_11684,N_8033,N_6345);
or U11685 (N_11685,N_7694,N_9439);
or U11686 (N_11686,N_7319,N_5349);
nand U11687 (N_11687,N_5715,N_6612);
and U11688 (N_11688,N_9274,N_5830);
nor U11689 (N_11689,N_8797,N_6054);
xor U11690 (N_11690,N_5934,N_9951);
or U11691 (N_11691,N_6697,N_6664);
nor U11692 (N_11692,N_6068,N_8044);
nor U11693 (N_11693,N_6423,N_5286);
xor U11694 (N_11694,N_6890,N_5122);
nor U11695 (N_11695,N_6855,N_9527);
and U11696 (N_11696,N_8081,N_5427);
and U11697 (N_11697,N_5472,N_9874);
nor U11698 (N_11698,N_9595,N_9240);
and U11699 (N_11699,N_5128,N_6109);
nand U11700 (N_11700,N_9778,N_8841);
and U11701 (N_11701,N_6115,N_7375);
nand U11702 (N_11702,N_5075,N_5843);
and U11703 (N_11703,N_9995,N_8821);
nor U11704 (N_11704,N_7999,N_6401);
nor U11705 (N_11705,N_6177,N_7302);
nand U11706 (N_11706,N_7020,N_7133);
xnor U11707 (N_11707,N_6589,N_8712);
or U11708 (N_11708,N_6333,N_8465);
or U11709 (N_11709,N_7384,N_6681);
nand U11710 (N_11710,N_8183,N_6902);
nor U11711 (N_11711,N_7462,N_9587);
nand U11712 (N_11712,N_6211,N_7851);
nand U11713 (N_11713,N_8408,N_7037);
nand U11714 (N_11714,N_9285,N_5542);
nand U11715 (N_11715,N_7188,N_5792);
nor U11716 (N_11716,N_5484,N_5950);
nor U11717 (N_11717,N_5878,N_6093);
or U11718 (N_11718,N_5710,N_6863);
or U11719 (N_11719,N_7705,N_7570);
and U11720 (N_11720,N_8867,N_5732);
nor U11721 (N_11721,N_7266,N_6447);
nor U11722 (N_11722,N_7907,N_5654);
nand U11723 (N_11723,N_8479,N_9508);
nand U11724 (N_11724,N_6173,N_9674);
and U11725 (N_11725,N_8869,N_5981);
and U11726 (N_11726,N_5945,N_7565);
and U11727 (N_11727,N_9576,N_8766);
or U11728 (N_11728,N_5295,N_9324);
and U11729 (N_11729,N_5351,N_5610);
nor U11730 (N_11730,N_9827,N_7567);
nand U11731 (N_11731,N_5565,N_5102);
nor U11732 (N_11732,N_5143,N_5503);
or U11733 (N_11733,N_8158,N_9499);
nand U11734 (N_11734,N_5582,N_7110);
nor U11735 (N_11735,N_7853,N_7212);
or U11736 (N_11736,N_6104,N_8578);
or U11737 (N_11737,N_8817,N_9481);
and U11738 (N_11738,N_7836,N_6690);
nand U11739 (N_11739,N_8226,N_5279);
nand U11740 (N_11740,N_7976,N_8014);
nand U11741 (N_11741,N_6998,N_9954);
and U11742 (N_11742,N_6370,N_7205);
nand U11743 (N_11743,N_8605,N_6049);
nand U11744 (N_11744,N_5224,N_5159);
nand U11745 (N_11745,N_6776,N_7894);
nor U11746 (N_11746,N_9952,N_8851);
nand U11747 (N_11747,N_7419,N_8167);
and U11748 (N_11748,N_6193,N_7135);
and U11749 (N_11749,N_6056,N_7421);
nor U11750 (N_11750,N_5725,N_8734);
xnor U11751 (N_11751,N_6236,N_8493);
nand U11752 (N_11752,N_5662,N_5116);
nor U11753 (N_11753,N_5346,N_5241);
or U11754 (N_11754,N_6250,N_7376);
or U11755 (N_11755,N_8170,N_8787);
or U11756 (N_11756,N_7867,N_9726);
nand U11757 (N_11757,N_9123,N_5035);
and U11758 (N_11758,N_9539,N_6784);
or U11759 (N_11759,N_6654,N_9503);
or U11760 (N_11760,N_7409,N_6006);
or U11761 (N_11761,N_6424,N_9059);
nor U11762 (N_11762,N_9616,N_6504);
and U11763 (N_11763,N_9103,N_8104);
and U11764 (N_11764,N_8597,N_8532);
or U11765 (N_11765,N_9162,N_7245);
nand U11766 (N_11766,N_5353,N_6244);
nand U11767 (N_11767,N_7961,N_6644);
and U11768 (N_11768,N_5498,N_6665);
and U11769 (N_11769,N_7253,N_9429);
nor U11770 (N_11770,N_5230,N_7142);
xnor U11771 (N_11771,N_5553,N_7903);
or U11772 (N_11772,N_6645,N_5480);
and U11773 (N_11773,N_8038,N_7380);
and U11774 (N_11774,N_5500,N_8231);
or U11775 (N_11775,N_5908,N_5406);
xor U11776 (N_11776,N_7257,N_5849);
and U11777 (N_11777,N_7036,N_6990);
and U11778 (N_11778,N_9875,N_9990);
nand U11779 (N_11779,N_5973,N_5458);
nor U11780 (N_11780,N_7633,N_5125);
nand U11781 (N_11781,N_6415,N_9361);
or U11782 (N_11782,N_6271,N_5810);
nand U11783 (N_11783,N_5988,N_6042);
nand U11784 (N_11784,N_8053,N_5518);
nand U11785 (N_11785,N_6809,N_5052);
or U11786 (N_11786,N_6061,N_7737);
nor U11787 (N_11787,N_8345,N_8561);
or U11788 (N_11788,N_5064,N_5401);
or U11789 (N_11789,N_8514,N_7656);
or U11790 (N_11790,N_9730,N_6420);
nand U11791 (N_11791,N_7612,N_7769);
nand U11792 (N_11792,N_6816,N_9072);
nand U11793 (N_11793,N_7109,N_6121);
or U11794 (N_11794,N_5687,N_5897);
nor U11795 (N_11795,N_5841,N_9941);
nor U11796 (N_11796,N_5047,N_5527);
and U11797 (N_11797,N_5263,N_8804);
nor U11798 (N_11798,N_9537,N_7884);
and U11799 (N_11799,N_6846,N_9427);
nor U11800 (N_11800,N_6073,N_9477);
or U11801 (N_11801,N_8035,N_7657);
nand U11802 (N_11802,N_5138,N_7653);
nand U11803 (N_11803,N_6593,N_5617);
or U11804 (N_11804,N_6764,N_8596);
nor U11805 (N_11805,N_6434,N_6443);
nand U11806 (N_11806,N_8009,N_8149);
or U11807 (N_11807,N_7201,N_5266);
and U11808 (N_11808,N_7509,N_7413);
or U11809 (N_11809,N_5935,N_7246);
or U11810 (N_11810,N_6899,N_6055);
or U11811 (N_11811,N_5641,N_6655);
and U11812 (N_11812,N_6238,N_8071);
nor U11813 (N_11813,N_7150,N_6536);
nor U11814 (N_11814,N_5892,N_5974);
nand U11815 (N_11815,N_5462,N_9462);
nand U11816 (N_11816,N_5975,N_8083);
or U11817 (N_11817,N_8962,N_8701);
nand U11818 (N_11818,N_7521,N_8762);
or U11819 (N_11819,N_9115,N_5555);
and U11820 (N_11820,N_9396,N_8108);
or U11821 (N_11821,N_6215,N_8875);
and U11822 (N_11822,N_8376,N_9341);
nor U11823 (N_11823,N_5900,N_7522);
or U11824 (N_11824,N_9538,N_6942);
and U11825 (N_11825,N_5060,N_8557);
or U11826 (N_11826,N_9487,N_9641);
and U11827 (N_11827,N_6064,N_9969);
nand U11828 (N_11828,N_7048,N_7158);
nand U11829 (N_11829,N_9326,N_5196);
and U11830 (N_11830,N_9171,N_8850);
and U11831 (N_11831,N_7689,N_7706);
nor U11832 (N_11832,N_7843,N_8464);
or U11833 (N_11833,N_5038,N_5007);
nand U11834 (N_11834,N_9389,N_5942);
nor U11835 (N_11835,N_5818,N_7630);
and U11836 (N_11836,N_9079,N_9051);
nor U11837 (N_11837,N_8445,N_5872);
or U11838 (N_11838,N_5685,N_5300);
nor U11839 (N_11839,N_5814,N_7778);
nand U11840 (N_11840,N_9758,N_6524);
and U11841 (N_11841,N_7586,N_5522);
nor U11842 (N_11842,N_9463,N_8130);
and U11843 (N_11843,N_8429,N_6409);
and U11844 (N_11844,N_7295,N_5719);
or U11845 (N_11845,N_5334,N_8604);
nor U11846 (N_11846,N_5131,N_9559);
nand U11847 (N_11847,N_7527,N_9703);
nand U11848 (N_11848,N_9656,N_5304);
or U11849 (N_11849,N_6259,N_5567);
nor U11850 (N_11850,N_9035,N_7255);
or U11851 (N_11851,N_8728,N_6414);
or U11852 (N_11852,N_5760,N_9368);
and U11853 (N_11853,N_6461,N_5451);
or U11854 (N_11854,N_9017,N_9348);
nand U11855 (N_11855,N_7332,N_6918);
nor U11856 (N_11856,N_8255,N_9702);
and U11857 (N_11857,N_6802,N_8726);
and U11858 (N_11858,N_5671,N_7599);
or U11859 (N_11859,N_6125,N_5980);
and U11860 (N_11860,N_7554,N_6449);
and U11861 (N_11861,N_6769,N_6377);
xnor U11862 (N_11862,N_8260,N_5796);
nand U11863 (N_11863,N_7066,N_5548);
or U11864 (N_11864,N_6577,N_8016);
nand U11865 (N_11865,N_7221,N_5217);
nand U11866 (N_11866,N_5097,N_9687);
nand U11867 (N_11867,N_8873,N_8719);
nor U11868 (N_11868,N_9898,N_5056);
nor U11869 (N_11869,N_8001,N_7279);
or U11870 (N_11870,N_6937,N_9903);
or U11871 (N_11871,N_8298,N_6570);
or U11872 (N_11872,N_6762,N_9683);
and U11873 (N_11873,N_5041,N_6000);
nor U11874 (N_11874,N_9437,N_6828);
nor U11875 (N_11875,N_9722,N_6120);
nand U11876 (N_11876,N_9511,N_7366);
and U11877 (N_11877,N_8727,N_7628);
nand U11878 (N_11878,N_7543,N_6591);
nand U11879 (N_11879,N_7491,N_9222);
nand U11880 (N_11880,N_6057,N_8487);
and U11881 (N_11881,N_7732,N_6575);
or U11882 (N_11882,N_8546,N_5253);
or U11883 (N_11883,N_6845,N_5738);
or U11884 (N_11884,N_8816,N_6094);
nand U11885 (N_11885,N_8279,N_5298);
nor U11886 (N_11886,N_6562,N_5591);
nor U11887 (N_11887,N_9933,N_9451);
nor U11888 (N_11888,N_6640,N_8903);
or U11889 (N_11889,N_5507,N_9247);
or U11890 (N_11890,N_6882,N_9038);
nand U11891 (N_11891,N_7584,N_9382);
or U11892 (N_11892,N_7365,N_8680);
nor U11893 (N_11893,N_7735,N_5237);
and U11894 (N_11894,N_7098,N_9597);
and U11895 (N_11895,N_9655,N_8662);
nor U11896 (N_11896,N_9585,N_8721);
or U11897 (N_11897,N_6979,N_5463);
or U11898 (N_11898,N_6403,N_9841);
and U11899 (N_11899,N_7029,N_5050);
or U11900 (N_11900,N_6277,N_9208);
nor U11901 (N_11901,N_7164,N_8745);
or U11902 (N_11902,N_9306,N_9582);
nor U11903 (N_11903,N_7879,N_8570);
nand U11904 (N_11904,N_6246,N_8599);
and U11905 (N_11905,N_9256,N_5410);
nand U11906 (N_11906,N_8714,N_9588);
and U11907 (N_11907,N_9746,N_5731);
xnor U11908 (N_11908,N_9077,N_8414);
or U11909 (N_11909,N_7051,N_5756);
nand U11910 (N_11910,N_6870,N_9580);
nor U11911 (N_11911,N_7138,N_9740);
or U11912 (N_11912,N_7856,N_6892);
and U11913 (N_11913,N_9739,N_7297);
nor U11914 (N_11914,N_6522,N_6059);
nand U11915 (N_11915,N_8642,N_8461);
and U11916 (N_11916,N_5296,N_6756);
and U11917 (N_11917,N_9027,N_7236);
or U11918 (N_11918,N_5608,N_6818);
or U11919 (N_11919,N_9996,N_6507);
nand U11920 (N_11920,N_5112,N_9364);
nor U11921 (N_11921,N_9426,N_7523);
or U11922 (N_11922,N_8836,N_5479);
nand U11923 (N_11923,N_6405,N_6679);
and U11924 (N_11924,N_6074,N_9121);
nor U11925 (N_11925,N_5234,N_7878);
and U11926 (N_11926,N_8432,N_6018);
nor U11927 (N_11927,N_7839,N_7950);
and U11928 (N_11928,N_9195,N_5602);
and U11929 (N_11929,N_5409,N_5963);
and U11930 (N_11930,N_7996,N_6398);
nor U11931 (N_11931,N_5071,N_5101);
or U11932 (N_11932,N_9822,N_8918);
and U11933 (N_11933,N_6324,N_5108);
and U11934 (N_11934,N_7165,N_5104);
nor U11935 (N_11935,N_9608,N_9058);
nor U11936 (N_11936,N_8301,N_9127);
nor U11937 (N_11937,N_9495,N_6549);
and U11938 (N_11938,N_9289,N_8891);
nand U11939 (N_11939,N_7174,N_9513);
or U11940 (N_11940,N_9254,N_8795);
nand U11941 (N_11941,N_5152,N_6975);
and U11942 (N_11942,N_6336,N_8855);
nand U11943 (N_11943,N_9216,N_9305);
nand U11944 (N_11944,N_6930,N_5538);
and U11945 (N_11945,N_9398,N_7354);
nand U11946 (N_11946,N_7097,N_7504);
or U11947 (N_11947,N_6968,N_7476);
xnor U11948 (N_11948,N_8729,N_9840);
nand U11949 (N_11949,N_7352,N_8211);
nand U11950 (N_11950,N_8931,N_6653);
nor U11951 (N_11951,N_6958,N_9235);
nand U11952 (N_11952,N_8529,N_6799);
nand U11953 (N_11953,N_5505,N_7125);
and U11954 (N_11954,N_9877,N_6020);
and U11955 (N_11955,N_9153,N_9565);
or U11956 (N_11956,N_8799,N_7390);
and U11957 (N_11957,N_8392,N_6353);
nand U11958 (N_11958,N_5347,N_9266);
nor U11959 (N_11959,N_8217,N_8544);
nor U11960 (N_11960,N_8327,N_9467);
xnor U11961 (N_11961,N_9143,N_8803);
nand U11962 (N_11962,N_8992,N_9098);
and U11963 (N_11963,N_8252,N_5851);
nor U11964 (N_11964,N_8077,N_7067);
nand U11965 (N_11965,N_7161,N_5672);
or U11966 (N_11966,N_7824,N_9670);
or U11967 (N_11967,N_8813,N_6497);
and U11968 (N_11968,N_7743,N_7709);
or U11969 (N_11969,N_7364,N_8336);
nor U11970 (N_11970,N_6989,N_7625);
or U11971 (N_11971,N_9183,N_9409);
and U11972 (N_11972,N_6689,N_6485);
and U11973 (N_11973,N_6922,N_7111);
nor U11974 (N_11974,N_5993,N_8624);
nor U11975 (N_11975,N_5620,N_5989);
nand U11976 (N_11976,N_7449,N_8870);
and U11977 (N_11977,N_9378,N_9203);
and U11978 (N_11978,N_6166,N_6298);
nor U11979 (N_11979,N_8651,N_7772);
nand U11980 (N_11980,N_7992,N_6307);
or U11981 (N_11981,N_5168,N_8213);
nand U11982 (N_11982,N_6435,N_9190);
nor U11983 (N_11983,N_9172,N_6533);
xnor U11984 (N_11984,N_9583,N_7905);
nor U11985 (N_11985,N_5509,N_9549);
and U11986 (N_11986,N_9459,N_5070);
or U11987 (N_11987,N_8072,N_5664);
or U11988 (N_11988,N_7341,N_6834);
nand U11989 (N_11989,N_7039,N_7887);
nor U11990 (N_11990,N_6181,N_6487);
or U11991 (N_11991,N_8986,N_7213);
nor U11992 (N_11992,N_6606,N_7335);
or U11993 (N_11993,N_7080,N_5436);
and U11994 (N_11994,N_6451,N_8921);
or U11995 (N_11995,N_5170,N_7978);
nor U11996 (N_11996,N_7604,N_6195);
nor U11997 (N_11997,N_9605,N_6714);
nor U11998 (N_11998,N_7835,N_9894);
nor U11999 (N_11999,N_6565,N_6518);
or U12000 (N_12000,N_7461,N_7010);
and U12001 (N_12001,N_8899,N_6571);
nor U12002 (N_12002,N_6651,N_5646);
nand U12003 (N_12003,N_7275,N_9280);
nand U12004 (N_12004,N_8042,N_9029);
or U12005 (N_12005,N_7683,N_7745);
nor U12006 (N_12006,N_9690,N_9390);
or U12007 (N_12007,N_9234,N_6127);
or U12008 (N_12008,N_9814,N_8172);
and U12009 (N_12009,N_9575,N_5560);
and U12010 (N_12010,N_5431,N_8559);
nand U12011 (N_12011,N_6952,N_5611);
or U12012 (N_12012,N_8550,N_7338);
nand U12013 (N_12013,N_6153,N_8938);
or U12014 (N_12014,N_7435,N_8242);
xnor U12015 (N_12015,N_6737,N_9784);
nand U12016 (N_12016,N_7963,N_6316);
nor U12017 (N_12017,N_7323,N_9366);
nor U12018 (N_12018,N_9019,N_9101);
nand U12019 (N_12019,N_8208,N_9497);
or U12020 (N_12020,N_5648,N_6995);
and U12021 (N_12021,N_5647,N_9053);
nor U12022 (N_12022,N_6494,N_8563);
nand U12023 (N_12023,N_7923,N_9679);
nor U12024 (N_12024,N_6303,N_5278);
or U12025 (N_12025,N_6095,N_9782);
nor U12026 (N_12026,N_5574,N_9742);
nand U12027 (N_12027,N_9562,N_7498);
nand U12028 (N_12028,N_6946,N_9046);
nor U12029 (N_12029,N_5197,N_5726);
nor U12030 (N_12030,N_9185,N_6988);
nand U12031 (N_12031,N_5411,N_9211);
nand U12032 (N_12032,N_8339,N_5584);
nor U12033 (N_12033,N_7862,N_9750);
and U12034 (N_12034,N_6779,N_8451);
and U12035 (N_12035,N_7117,N_6709);
nand U12036 (N_12036,N_6626,N_8743);
nor U12037 (N_12037,N_8639,N_7227);
xor U12038 (N_12038,N_9423,N_5562);
or U12039 (N_12039,N_6139,N_5011);
and U12040 (N_12040,N_5531,N_8522);
nor U12041 (N_12041,N_8197,N_5577);
nor U12042 (N_12042,N_9054,N_7530);
nand U12043 (N_12043,N_5645,N_9097);
or U12044 (N_12044,N_7768,N_7342);
and U12045 (N_12045,N_6965,N_6011);
or U12046 (N_12046,N_7007,N_9545);
or U12047 (N_12047,N_9081,N_6155);
or U12048 (N_12048,N_7975,N_6797);
nor U12049 (N_12049,N_6578,N_6694);
and U12050 (N_12050,N_6300,N_9344);
nand U12051 (N_12051,N_7382,N_7592);
nor U12052 (N_12052,N_9142,N_7190);
and U12053 (N_12053,N_8296,N_8175);
or U12054 (N_12054,N_5161,N_9892);
and U12055 (N_12055,N_8438,N_8480);
nor U12056 (N_12056,N_8603,N_8718);
and U12057 (N_12057,N_6947,N_7983);
nor U12058 (N_12058,N_8299,N_7196);
nor U12059 (N_12059,N_9711,N_9708);
or U12060 (N_12060,N_8384,N_9956);
and U12061 (N_12061,N_9350,N_9311);
and U12062 (N_12062,N_8326,N_8349);
xnor U12063 (N_12063,N_5144,N_7134);
nor U12064 (N_12064,N_5951,N_7717);
and U12065 (N_12065,N_8794,N_6131);
or U12066 (N_12066,N_5868,N_5790);
and U12067 (N_12067,N_5718,N_6595);
and U12068 (N_12068,N_9354,N_5171);
nor U12069 (N_12069,N_8942,N_6268);
or U12070 (N_12070,N_5252,N_9126);
and U12071 (N_12071,N_9837,N_9271);
and U12072 (N_12072,N_8634,N_5815);
or U12073 (N_12073,N_8103,N_8629);
or U12074 (N_12074,N_5893,N_9573);
and U12075 (N_12075,N_9797,N_8878);
nor U12076 (N_12076,N_7344,N_7956);
or U12077 (N_12077,N_6708,N_6751);
and U12078 (N_12078,N_6837,N_5572);
and U12079 (N_12079,N_6746,N_6794);
nand U12080 (N_12080,N_6561,N_8046);
nor U12081 (N_12081,N_6814,N_9309);
and U12082 (N_12082,N_9895,N_8030);
nand U12083 (N_12083,N_5652,N_8632);
or U12084 (N_12084,N_5027,N_9210);
nor U12085 (N_12085,N_6274,N_5434);
and U12086 (N_12086,N_6774,N_5306);
nor U12087 (N_12087,N_8711,N_5068);
nor U12088 (N_12088,N_6489,N_7270);
nor U12089 (N_12089,N_8861,N_5213);
nand U12090 (N_12090,N_8256,N_8874);
nand U12091 (N_12091,N_5823,N_6078);
nand U12092 (N_12092,N_8698,N_5369);
nor U12093 (N_12093,N_7774,N_8683);
or U12094 (N_12094,N_6605,N_9851);
nor U12095 (N_12095,N_9130,N_7986);
and U12096 (N_12096,N_7139,N_6627);
and U12097 (N_12097,N_8367,N_9104);
or U12098 (N_12098,N_5420,N_5949);
nand U12099 (N_12099,N_6235,N_6927);
or U12100 (N_12100,N_7675,N_6218);
nor U12101 (N_12101,N_8373,N_7746);
and U12102 (N_12102,N_8281,N_5766);
or U12103 (N_12103,N_8572,N_5590);
and U12104 (N_12104,N_6647,N_5348);
and U12105 (N_12105,N_9048,N_7895);
and U12106 (N_12106,N_8065,N_5550);
nor U12107 (N_12107,N_5151,N_9196);
and U12108 (N_12108,N_9963,N_6079);
or U12109 (N_12109,N_9160,N_7367);
or U12110 (N_12110,N_7714,N_9928);
nor U12111 (N_12111,N_9205,N_6198);
or U12112 (N_12112,N_9322,N_5906);
nand U12113 (N_12113,N_5547,N_6842);
and U12114 (N_12114,N_7456,N_6804);
and U12115 (N_12115,N_8235,N_6542);
nor U12116 (N_12116,N_7926,N_6934);
nor U12117 (N_12117,N_8411,N_5624);
and U12118 (N_12118,N_9412,N_8500);
and U12119 (N_12119,N_8556,N_5094);
or U12120 (N_12120,N_5502,N_6282);
or U12121 (N_12121,N_5697,N_8613);
nand U12122 (N_12122,N_8845,N_7349);
or U12123 (N_12123,N_8297,N_6763);
and U12124 (N_12124,N_7490,N_6581);
nor U12125 (N_12125,N_5363,N_9090);
or U12126 (N_12126,N_7801,N_7917);
or U12127 (N_12127,N_6670,N_9603);
nor U12128 (N_12128,N_5466,N_6199);
nor U12129 (N_12129,N_6649,N_6858);
and U12130 (N_12130,N_7643,N_6486);
or U12131 (N_12131,N_5535,N_9428);
nand U12132 (N_12132,N_5208,N_9342);
and U12133 (N_12133,N_8748,N_6843);
nor U12134 (N_12134,N_5777,N_9353);
nor U12135 (N_12135,N_6201,N_7327);
nand U12136 (N_12136,N_5880,N_6097);
and U12137 (N_12137,N_7260,N_8452);
or U12138 (N_12138,N_9227,N_8269);
or U12139 (N_12139,N_7415,N_6667);
and U12140 (N_12140,N_5032,N_5328);
nand U12141 (N_12141,N_5520,N_9783);
and U12142 (N_12142,N_7120,N_7441);
or U12143 (N_12143,N_5984,N_7088);
and U12144 (N_12144,N_5964,N_5062);
nor U12145 (N_12145,N_7617,N_5474);
or U12146 (N_12146,N_8979,N_6152);
and U12147 (N_12147,N_5103,N_5163);
nor U12148 (N_12148,N_6080,N_6926);
nand U12149 (N_12149,N_9856,N_5001);
and U12150 (N_12150,N_9231,N_5179);
nor U12151 (N_12151,N_6543,N_5301);
nand U12152 (N_12152,N_5174,N_6229);
nor U12153 (N_12153,N_9906,N_5405);
nor U12154 (N_12154,N_8768,N_7385);
or U12155 (N_12155,N_6786,N_8002);
nor U12156 (N_12156,N_8871,N_6933);
nand U12157 (N_12157,N_6087,N_5073);
nand U12158 (N_12158,N_6544,N_7922);
nor U12159 (N_12159,N_8562,N_8755);
and U12160 (N_12160,N_6328,N_6691);
or U12161 (N_12161,N_5394,N_7104);
nand U12162 (N_12162,N_8737,N_8308);
nor U12163 (N_12163,N_6007,N_6407);
nand U12164 (N_12164,N_6966,N_8348);
or U12165 (N_12165,N_7315,N_9307);
nor U12166 (N_12166,N_6464,N_6559);
and U12167 (N_12167,N_8509,N_6806);
nand U12168 (N_12168,N_7674,N_7402);
xnor U12169 (N_12169,N_9533,N_6666);
nand U12170 (N_12170,N_5795,N_8569);
or U12171 (N_12171,N_5227,N_6212);
or U12172 (N_12172,N_6646,N_6680);
and U12173 (N_12173,N_9003,N_9376);
nand U12174 (N_12174,N_6669,N_5142);
and U12175 (N_12175,N_6428,N_6358);
and U12176 (N_12176,N_6248,N_9967);
or U12177 (N_12177,N_6867,N_7296);
nand U12178 (N_12178,N_9283,N_8486);
and U12179 (N_12179,N_5367,N_7913);
or U12180 (N_12180,N_6984,N_5888);
nand U12181 (N_12181,N_5835,N_8306);
nor U12182 (N_12182,N_7588,N_8067);
and U12183 (N_12183,N_6135,N_6322);
nor U12184 (N_12184,N_5355,N_8863);
nor U12185 (N_12185,N_7416,N_8472);
nand U12186 (N_12186,N_8401,N_9660);
nor U12187 (N_12187,N_6916,N_5274);
or U12188 (N_12188,N_8457,N_5383);
and U12189 (N_12189,N_7971,N_5136);
or U12190 (N_12190,N_5832,N_6251);
and U12191 (N_12191,N_7105,N_6015);
nand U12192 (N_12192,N_9315,N_8225);
and U12193 (N_12193,N_7608,N_6225);
or U12194 (N_12194,N_9932,N_8209);
nand U12195 (N_12195,N_9221,N_8276);
or U12196 (N_12196,N_7941,N_8583);
or U12197 (N_12197,N_7055,N_6541);
nand U12198 (N_12198,N_6671,N_8129);
nor U12199 (N_12199,N_6369,N_8636);
nand U12200 (N_12200,N_9372,N_7351);
nor U12201 (N_12201,N_8601,N_7906);
or U12202 (N_12202,N_7084,N_6766);
nand U12203 (N_12203,N_7087,N_6146);
or U12204 (N_12204,N_8154,N_5998);
nand U12205 (N_12205,N_7483,N_8977);
nor U12206 (N_12206,N_7531,N_7687);
nand U12207 (N_12207,N_9905,N_6829);
nand U12208 (N_12208,N_6380,N_9359);
and U12209 (N_12209,N_8442,N_5508);
nor U12210 (N_12210,N_8371,N_6477);
or U12211 (N_12211,N_7264,N_7019);
nor U12212 (N_12212,N_6404,N_8161);
or U12213 (N_12213,N_6444,N_5812);
nand U12214 (N_12214,N_5130,N_9493);
nand U12215 (N_12215,N_5622,N_9225);
nor U12216 (N_12216,N_8545,N_6868);
or U12217 (N_12217,N_8538,N_5189);
nor U12218 (N_12218,N_9401,N_8846);
and U12219 (N_12219,N_7473,N_7121);
or U12220 (N_12220,N_8230,N_8485);
nand U12221 (N_12221,N_8966,N_8967);
or U12222 (N_12222,N_5909,N_8066);
or U12223 (N_12223,N_6889,N_6349);
and U12224 (N_12224,N_9831,N_7049);
or U12225 (N_12225,N_8482,N_5190);
and U12226 (N_12226,N_7328,N_9908);
nor U12227 (N_12227,N_6356,N_5067);
xnor U12228 (N_12228,N_5255,N_5587);
or U12229 (N_12229,N_9303,N_8004);
nor U12230 (N_12230,N_8585,N_9033);
or U12231 (N_12231,N_9962,N_9880);
nand U12232 (N_12232,N_7618,N_7806);
nand U12233 (N_12233,N_7805,N_5739);
nand U12234 (N_12234,N_6326,N_6865);
nor U12235 (N_12235,N_7273,N_5061);
nand U12236 (N_12236,N_8694,N_6085);
nand U12237 (N_12237,N_9272,N_8536);
nand U12238 (N_12238,N_5299,N_6320);
nand U12239 (N_12239,N_9771,N_8635);
or U12240 (N_12240,N_6160,N_8612);
and U12241 (N_12241,N_6907,N_9251);
and U12242 (N_12242,N_9601,N_7175);
nand U12243 (N_12243,N_7651,N_5180);
or U12244 (N_12244,N_6901,N_6773);
nor U12245 (N_12245,N_6910,N_9714);
nor U12246 (N_12246,N_7645,N_7408);
nand U12247 (N_12247,N_9173,N_9590);
nand U12248 (N_12248,N_7005,N_8660);
nand U12249 (N_12249,N_9884,N_5195);
nand U12250 (N_12250,N_9300,N_8416);
or U12251 (N_12251,N_9076,N_7356);
or U12252 (N_12252,N_8832,N_8913);
and U12253 (N_12253,N_6327,N_7422);
nand U12254 (N_12254,N_9091,N_8382);
nand U12255 (N_12255,N_5700,N_9735);
nor U12256 (N_12256,N_8881,N_8112);
nor U12257 (N_12257,N_6368,N_7495);
or U12258 (N_12258,N_6043,N_5088);
nand U12259 (N_12259,N_6550,N_8468);
nor U12260 (N_12260,N_5251,N_9008);
and U12261 (N_12261,N_5188,N_5475);
and U12262 (N_12262,N_6791,N_9912);
and U12263 (N_12263,N_5415,N_9316);
and U12264 (N_12264,N_6310,N_6374);
and U12265 (N_12265,N_6293,N_5928);
and U12266 (N_12266,N_6179,N_9214);
nor U12267 (N_12267,N_9419,N_7099);
and U12268 (N_12268,N_6747,N_9082);
nor U12269 (N_12269,N_9087,N_7832);
nor U12270 (N_12270,N_7869,N_7044);
nand U12271 (N_12271,N_7453,N_5896);
nand U12272 (N_12272,N_6111,N_6904);
or U12273 (N_12273,N_9167,N_7542);
nand U12274 (N_12274,N_8594,N_8619);
and U12275 (N_12275,N_5390,N_6939);
or U12276 (N_12276,N_6473,N_8773);
or U12277 (N_12277,N_7520,N_9193);
or U12278 (N_12278,N_9204,N_8814);
and U12279 (N_12279,N_7638,N_6400);
nor U12280 (N_12280,N_6833,N_7615);
and U12281 (N_12281,N_9329,N_9944);
or U12282 (N_12282,N_5184,N_6105);
or U12283 (N_12283,N_6280,N_7220);
or U12284 (N_12284,N_9199,N_5825);
xnor U12285 (N_12285,N_5317,N_6340);
nand U12286 (N_12286,N_9927,N_6241);
or U12287 (N_12287,N_5269,N_9400);
or U12288 (N_12288,N_9883,N_8407);
and U12289 (N_12289,N_9238,N_8810);
nor U12290 (N_12290,N_5074,N_9334);
nor U12291 (N_12291,N_5918,N_7818);
nand U12292 (N_12292,N_8391,N_8135);
and U12293 (N_12293,N_5869,N_5894);
or U12294 (N_12294,N_7189,N_7661);
nor U12295 (N_12295,N_5865,N_6614);
and U12296 (N_12296,N_8483,N_7059);
or U12297 (N_12297,N_7085,N_7789);
nor U12298 (N_12298,N_9617,N_8646);
nand U12299 (N_12299,N_8192,N_5417);
and U12300 (N_12300,N_6468,N_7631);
or U12301 (N_12301,N_7463,N_7744);
and U12302 (N_12302,N_7568,N_5695);
and U12303 (N_12303,N_5757,N_7794);
nor U12304 (N_12304,N_6308,N_6983);
nand U12305 (N_12305,N_5979,N_7263);
nand U12306 (N_12306,N_9943,N_6124);
and U12307 (N_12307,N_8000,N_8285);
or U12308 (N_12308,N_8839,N_7128);
or U12309 (N_12309,N_9370,N_7414);
xor U12310 (N_12310,N_6758,N_7333);
or U12311 (N_12311,N_5340,N_7460);
nand U12312 (N_12312,N_7788,N_9404);
nor U12313 (N_12313,N_5345,N_6242);
nor U12314 (N_12314,N_8691,N_7955);
nor U12315 (N_12315,N_6033,N_9198);
xnor U12316 (N_12316,N_6005,N_8681);
and U12317 (N_12317,N_7607,N_6847);
or U12318 (N_12318,N_7024,N_8690);
nand U12319 (N_12319,N_5483,N_7977);
nor U12320 (N_12320,N_5875,N_7518);
nand U12321 (N_12321,N_7606,N_8381);
and U12322 (N_12322,N_7426,N_5160);
xnor U12323 (N_12323,N_8375,N_8759);
nand U12324 (N_12324,N_9301,N_9625);
nand U12325 (N_12325,N_5905,N_5053);
nand U12326 (N_12326,N_5506,N_7076);
or U12327 (N_12327,N_8031,N_6063);
nor U12328 (N_12328,N_6133,N_9379);
or U12329 (N_12329,N_7000,N_7756);
xor U12330 (N_12330,N_9432,N_5539);
and U12331 (N_12331,N_6557,N_6941);
nor U12332 (N_12332,N_9916,N_5997);
nand U12333 (N_12333,N_5717,N_6266);
or U12334 (N_12334,N_8430,N_9155);
and U12335 (N_12335,N_8109,N_9629);
nand U12336 (N_12336,N_7181,N_5243);
nand U12337 (N_12337,N_6753,N_8052);
nor U12338 (N_12338,N_9818,N_9865);
nand U12339 (N_12339,N_7334,N_9055);
nand U12340 (N_12340,N_5772,N_5659);
nor U12341 (N_12341,N_9187,N_7713);
and U12342 (N_12342,N_5309,N_9447);
nand U12343 (N_12343,N_7795,N_8333);
and U12344 (N_12344,N_9403,N_5229);
and U12345 (N_12345,N_5827,N_9807);
nor U12346 (N_12346,N_9294,N_7984);
nor U12347 (N_12347,N_8188,N_6302);
nor U12348 (N_12348,N_7547,N_7294);
and U12349 (N_12349,N_5594,N_5341);
nor U12350 (N_12350,N_7812,N_6150);
nand U12351 (N_12351,N_7136,N_8970);
or U12352 (N_12352,N_9450,N_7751);
nand U12353 (N_12353,N_8444,N_5889);
xor U12354 (N_12354,N_9678,N_9346);
nor U12355 (N_12355,N_6699,N_9976);
or U12356 (N_12356,N_8394,N_9957);
and U12357 (N_12357,N_8521,N_8917);
or U12358 (N_12358,N_8139,N_6433);
and U12359 (N_12359,N_6898,N_7793);
nor U12360 (N_12360,N_8019,N_9986);
nand U12361 (N_12361,N_9946,N_6703);
nor U12362 (N_12362,N_9281,N_8145);
and U12363 (N_12363,N_7686,N_9592);
or U12364 (N_12364,N_5006,N_6118);
or U12365 (N_12365,N_9145,N_5147);
nor U12366 (N_12366,N_6950,N_8933);
or U12367 (N_12367,N_9188,N_8320);
and U12368 (N_12368,N_9080,N_8115);
nand U12369 (N_12369,N_6136,N_9938);
nor U12370 (N_12370,N_9384,N_8744);
nor U12371 (N_12371,N_6564,N_5741);
or U12372 (N_12372,N_7398,N_9931);
nand U12373 (N_12373,N_6894,N_5783);
and U12374 (N_12374,N_5021,N_6803);
nand U12375 (N_12375,N_9152,N_8092);
or U12376 (N_12376,N_8606,N_9729);
nand U12377 (N_12377,N_8396,N_8769);
or U12378 (N_12378,N_8877,N_7355);
and U12379 (N_12379,N_8389,N_6128);
or U12380 (N_12380,N_8060,N_8865);
nor U12381 (N_12381,N_5724,N_6107);
and U12382 (N_12382,N_6741,N_9050);
or U12383 (N_12383,N_5663,N_5543);
nand U12384 (N_12384,N_8360,N_7550);
nand U12385 (N_12385,N_5874,N_9700);
and U12386 (N_12386,N_6924,N_7126);
nand U12387 (N_12387,N_7129,N_9704);
nand U12388 (N_12388,N_6993,N_6350);
nand U12389 (N_12389,N_5020,N_9480);
nand U12390 (N_12390,N_6050,N_7891);
nand U12391 (N_12391,N_6810,N_7160);
nand U12392 (N_12392,N_6735,N_7322);
nand U12393 (N_12393,N_7237,N_9215);
nor U12394 (N_12394,N_9692,N_8383);
nor U12395 (N_12395,N_9713,N_6982);
nor U12396 (N_12396,N_7726,N_5819);
nor U12397 (N_12397,N_6954,N_7216);
or U12398 (N_12398,N_5028,N_6285);
nor U12399 (N_12399,N_9651,N_7231);
or U12400 (N_12400,N_6354,N_6716);
or U12401 (N_12401,N_7009,N_9548);
nor U12402 (N_12402,N_7154,N_5258);
nand U12403 (N_12403,N_6607,N_5859);
nor U12404 (N_12404,N_8346,N_7395);
xor U12405 (N_12405,N_9217,N_5651);
or U12406 (N_12406,N_6850,N_8715);
xor U12407 (N_12407,N_5177,N_9897);
nand U12408 (N_12408,N_6182,N_6289);
or U12409 (N_12409,N_7232,N_9457);
and U12410 (N_12410,N_9958,N_6347);
xor U12411 (N_12411,N_6625,N_9475);
nand U12412 (N_12412,N_5499,N_6396);
xor U12413 (N_12413,N_9940,N_7792);
and U12414 (N_12414,N_8328,N_9430);
nor U12415 (N_12415,N_9000,N_9113);
or U12416 (N_12416,N_6344,N_8590);
nand U12417 (N_12417,N_8807,N_6325);
nor U12418 (N_12418,N_7934,N_7192);
nand U12419 (N_12419,N_5737,N_9689);
nand U12420 (N_12420,N_9993,N_8248);
or U12421 (N_12421,N_8990,N_7857);
nand U12422 (N_12422,N_7179,N_6126);
or U12423 (N_12423,N_5961,N_9910);
or U12424 (N_12424,N_9793,N_8008);
or U12425 (N_12425,N_5069,N_9852);
nor U12426 (N_12426,N_5661,N_9756);
nand U12427 (N_12427,N_8611,N_6768);
and U12428 (N_12428,N_5676,N_5937);
nand U12429 (N_12429,N_9073,N_7359);
or U12430 (N_12430,N_5776,N_6731);
nor U12431 (N_12431,N_9552,N_6790);
nand U12432 (N_12432,N_8290,N_8133);
and U12433 (N_12433,N_7702,N_8607);
and U12434 (N_12434,N_5291,N_6001);
nand U12435 (N_12435,N_9200,N_7235);
and U12436 (N_12436,N_5120,N_9373);
nor U12437 (N_12437,N_7591,N_7838);
or U12438 (N_12438,N_5207,N_9911);
nor U12439 (N_12439,N_7749,N_6705);
nor U12440 (N_12440,N_5040,N_6034);
and U12441 (N_12441,N_6963,N_6511);
nand U12442 (N_12442,N_8352,N_9045);
and U12443 (N_12443,N_8322,N_5244);
and U12444 (N_12444,N_9844,N_9968);
nand U12445 (N_12445,N_6030,N_9699);
or U12446 (N_12446,N_9184,N_7998);
or U12447 (N_12447,N_9855,N_7254);
nor U12448 (N_12448,N_8043,N_8107);
nand U12449 (N_12449,N_6822,N_9192);
nand U12450 (N_12450,N_5287,N_8860);
or U12451 (N_12451,N_9443,N_7825);
and U12452 (N_12452,N_9260,N_6392);
nor U12453 (N_12453,N_7494,N_6171);
and U12454 (N_12454,N_8088,N_8118);
or U12455 (N_12455,N_6231,N_6657);
xnor U12456 (N_12456,N_8022,N_6066);
and U12457 (N_12457,N_7928,N_8082);
or U12458 (N_12458,N_5445,N_5004);
or U12459 (N_12459,N_9613,N_8834);
nand U12460 (N_12460,N_5393,N_5429);
and U12461 (N_12461,N_6854,N_8045);
nand U12462 (N_12462,N_7043,N_5779);
and U12463 (N_12463,N_8939,N_8541);
nand U12464 (N_12464,N_8473,N_6203);
or U12465 (N_12465,N_5365,N_8920);
nand U12466 (N_12466,N_9257,N_8974);
nor U12467 (N_12467,N_6530,N_5791);
and U12468 (N_12468,N_5765,N_7982);
nor U12469 (N_12469,N_5359,N_6516);
nor U12470 (N_12470,N_6364,N_7552);
and U12471 (N_12471,N_6987,N_8669);
nor U12472 (N_12472,N_5895,N_5491);
nor U12473 (N_12473,N_7493,N_9064);
nand U12474 (N_12474,N_7219,N_7545);
nand U12475 (N_12475,N_9624,N_8431);
and U12476 (N_12476,N_8778,N_5844);
nor U12477 (N_12477,N_8305,N_9998);
nand U12478 (N_12478,N_8708,N_5637);
nand U12479 (N_12479,N_7330,N_9168);
or U12480 (N_12480,N_5990,N_7823);
nor U12481 (N_12481,N_5066,N_8258);
nand U12482 (N_12482,N_9022,N_8574);
or U12483 (N_12483,N_5936,N_9555);
or U12484 (N_12484,N_7343,N_8220);
and U12485 (N_12485,N_9710,N_7692);
nor U12486 (N_12486,N_6636,N_9106);
nand U12487 (N_12487,N_9287,N_8663);
or U12488 (N_12488,N_6897,N_8566);
and U12489 (N_12489,N_7038,N_8731);
nor U12490 (N_12490,N_5592,N_7967);
or U12491 (N_12491,N_5871,N_8547);
and U12492 (N_12492,N_5107,N_6090);
and U12493 (N_12493,N_7965,N_9478);
nor U12494 (N_12494,N_6024,N_8028);
nor U12495 (N_12495,N_9135,N_5639);
or U12496 (N_12496,N_8434,N_5381);
or U12497 (N_12497,N_7927,N_7762);
and U12498 (N_12498,N_8075,N_5933);
xor U12499 (N_12499,N_9515,N_6216);
nand U12500 (N_12500,N_5356,N_8636);
nor U12501 (N_12501,N_8395,N_7946);
or U12502 (N_12502,N_5935,N_9142);
nand U12503 (N_12503,N_5844,N_6735);
and U12504 (N_12504,N_8777,N_6971);
or U12505 (N_12505,N_8762,N_6974);
nor U12506 (N_12506,N_5643,N_9202);
nor U12507 (N_12507,N_7311,N_5316);
and U12508 (N_12508,N_5318,N_7153);
or U12509 (N_12509,N_6016,N_6969);
or U12510 (N_12510,N_9238,N_7880);
and U12511 (N_12511,N_9324,N_8325);
nand U12512 (N_12512,N_5679,N_6843);
nand U12513 (N_12513,N_9336,N_5956);
or U12514 (N_12514,N_5126,N_7468);
or U12515 (N_12515,N_6652,N_8059);
and U12516 (N_12516,N_6210,N_9502);
and U12517 (N_12517,N_6420,N_5453);
or U12518 (N_12518,N_7358,N_7565);
nand U12519 (N_12519,N_8416,N_7008);
nor U12520 (N_12520,N_8494,N_7332);
nor U12521 (N_12521,N_9450,N_9050);
nor U12522 (N_12522,N_9040,N_5647);
nand U12523 (N_12523,N_7383,N_5831);
and U12524 (N_12524,N_6028,N_5074);
nor U12525 (N_12525,N_9579,N_7219);
nand U12526 (N_12526,N_8127,N_8105);
nand U12527 (N_12527,N_9666,N_5076);
xor U12528 (N_12528,N_6302,N_6172);
nor U12529 (N_12529,N_7329,N_9183);
nor U12530 (N_12530,N_6386,N_5392);
or U12531 (N_12531,N_6929,N_5197);
nor U12532 (N_12532,N_7277,N_9672);
or U12533 (N_12533,N_8195,N_9800);
and U12534 (N_12534,N_5579,N_9826);
nor U12535 (N_12535,N_5338,N_9481);
nor U12536 (N_12536,N_7028,N_8734);
nand U12537 (N_12537,N_8971,N_9788);
nand U12538 (N_12538,N_8877,N_7455);
and U12539 (N_12539,N_8491,N_9493);
and U12540 (N_12540,N_6450,N_9161);
nand U12541 (N_12541,N_5236,N_9824);
nor U12542 (N_12542,N_5109,N_8773);
nor U12543 (N_12543,N_9504,N_6759);
and U12544 (N_12544,N_6083,N_5527);
nor U12545 (N_12545,N_8349,N_7533);
and U12546 (N_12546,N_9009,N_7784);
nand U12547 (N_12547,N_8970,N_8588);
xor U12548 (N_12548,N_8139,N_5194);
nor U12549 (N_12549,N_8886,N_6869);
nand U12550 (N_12550,N_5718,N_5801);
nand U12551 (N_12551,N_8188,N_5719);
and U12552 (N_12552,N_5133,N_7904);
or U12553 (N_12553,N_6134,N_7499);
nor U12554 (N_12554,N_7598,N_7100);
and U12555 (N_12555,N_8084,N_6327);
or U12556 (N_12556,N_5300,N_7346);
or U12557 (N_12557,N_9561,N_6275);
and U12558 (N_12558,N_7360,N_7704);
and U12559 (N_12559,N_6123,N_9442);
and U12560 (N_12560,N_6971,N_5311);
nand U12561 (N_12561,N_6176,N_7940);
nor U12562 (N_12562,N_8842,N_9062);
nand U12563 (N_12563,N_9377,N_8268);
nor U12564 (N_12564,N_7333,N_8919);
xor U12565 (N_12565,N_6084,N_7558);
xnor U12566 (N_12566,N_9483,N_6425);
or U12567 (N_12567,N_7090,N_9187);
or U12568 (N_12568,N_8591,N_7765);
nor U12569 (N_12569,N_9606,N_9720);
nand U12570 (N_12570,N_7299,N_8556);
or U12571 (N_12571,N_9641,N_9279);
nand U12572 (N_12572,N_7130,N_9454);
nand U12573 (N_12573,N_8241,N_5347);
and U12574 (N_12574,N_5414,N_9527);
nand U12575 (N_12575,N_9855,N_5908);
and U12576 (N_12576,N_9445,N_5500);
nor U12577 (N_12577,N_8515,N_6290);
nor U12578 (N_12578,N_9611,N_5283);
and U12579 (N_12579,N_6417,N_6420);
nand U12580 (N_12580,N_9030,N_5833);
nand U12581 (N_12581,N_6385,N_9822);
xor U12582 (N_12582,N_8340,N_8930);
or U12583 (N_12583,N_9112,N_7837);
or U12584 (N_12584,N_6626,N_5853);
and U12585 (N_12585,N_6529,N_7518);
nand U12586 (N_12586,N_9104,N_9053);
and U12587 (N_12587,N_7692,N_6406);
and U12588 (N_12588,N_6891,N_8925);
nor U12589 (N_12589,N_8415,N_7976);
and U12590 (N_12590,N_5032,N_7727);
or U12591 (N_12591,N_7889,N_7225);
and U12592 (N_12592,N_9858,N_6753);
nor U12593 (N_12593,N_5897,N_6630);
nand U12594 (N_12594,N_7779,N_6088);
nand U12595 (N_12595,N_7807,N_5315);
nor U12596 (N_12596,N_9704,N_9714);
nand U12597 (N_12597,N_8098,N_9224);
and U12598 (N_12598,N_6492,N_6191);
or U12599 (N_12599,N_7390,N_9903);
and U12600 (N_12600,N_8750,N_6824);
nor U12601 (N_12601,N_9737,N_6702);
nor U12602 (N_12602,N_9981,N_6286);
nor U12603 (N_12603,N_9196,N_9699);
or U12604 (N_12604,N_9788,N_5834);
and U12605 (N_12605,N_9476,N_6981);
and U12606 (N_12606,N_6725,N_9181);
nor U12607 (N_12607,N_6525,N_8017);
and U12608 (N_12608,N_8961,N_8558);
or U12609 (N_12609,N_7783,N_8433);
nor U12610 (N_12610,N_8052,N_6896);
and U12611 (N_12611,N_8875,N_7282);
and U12612 (N_12612,N_5483,N_5014);
nand U12613 (N_12613,N_9716,N_8893);
or U12614 (N_12614,N_8650,N_8429);
and U12615 (N_12615,N_8059,N_7174);
nand U12616 (N_12616,N_7130,N_8352);
or U12617 (N_12617,N_5093,N_9469);
and U12618 (N_12618,N_9160,N_5014);
and U12619 (N_12619,N_7470,N_8450);
nand U12620 (N_12620,N_7297,N_6118);
or U12621 (N_12621,N_7647,N_6717);
nand U12622 (N_12622,N_7920,N_7404);
xnor U12623 (N_12623,N_6002,N_9975);
and U12624 (N_12624,N_9882,N_7180);
nand U12625 (N_12625,N_5858,N_8504);
and U12626 (N_12626,N_5483,N_5623);
nor U12627 (N_12627,N_6027,N_5402);
or U12628 (N_12628,N_8164,N_5261);
and U12629 (N_12629,N_5103,N_5866);
xnor U12630 (N_12630,N_9239,N_5523);
nand U12631 (N_12631,N_5104,N_7502);
nor U12632 (N_12632,N_8102,N_9964);
xnor U12633 (N_12633,N_5221,N_6616);
and U12634 (N_12634,N_7809,N_7792);
nand U12635 (N_12635,N_5236,N_5777);
nor U12636 (N_12636,N_6556,N_5252);
or U12637 (N_12637,N_8775,N_9356);
and U12638 (N_12638,N_5996,N_5668);
nor U12639 (N_12639,N_9762,N_6810);
and U12640 (N_12640,N_7651,N_7520);
or U12641 (N_12641,N_7421,N_7466);
xnor U12642 (N_12642,N_5034,N_9447);
nand U12643 (N_12643,N_6610,N_6770);
and U12644 (N_12644,N_7454,N_6232);
nand U12645 (N_12645,N_7759,N_7618);
nor U12646 (N_12646,N_5073,N_7878);
and U12647 (N_12647,N_5097,N_9372);
or U12648 (N_12648,N_8400,N_8618);
nand U12649 (N_12649,N_5886,N_9255);
and U12650 (N_12650,N_5562,N_5641);
or U12651 (N_12651,N_6782,N_8400);
or U12652 (N_12652,N_6924,N_5237);
nor U12653 (N_12653,N_5632,N_7882);
nor U12654 (N_12654,N_6898,N_6469);
nor U12655 (N_12655,N_9450,N_9543);
or U12656 (N_12656,N_7688,N_6943);
or U12657 (N_12657,N_9262,N_5505);
nor U12658 (N_12658,N_8395,N_7634);
and U12659 (N_12659,N_9838,N_5559);
nor U12660 (N_12660,N_6013,N_5387);
nand U12661 (N_12661,N_5541,N_8709);
and U12662 (N_12662,N_8243,N_9406);
and U12663 (N_12663,N_6069,N_9421);
nor U12664 (N_12664,N_9658,N_9504);
nand U12665 (N_12665,N_9513,N_7515);
or U12666 (N_12666,N_5890,N_8707);
nand U12667 (N_12667,N_8970,N_5004);
and U12668 (N_12668,N_7726,N_9823);
nor U12669 (N_12669,N_6333,N_6628);
nor U12670 (N_12670,N_6780,N_5970);
nand U12671 (N_12671,N_7381,N_8699);
nor U12672 (N_12672,N_7904,N_7750);
or U12673 (N_12673,N_6477,N_9039);
or U12674 (N_12674,N_6444,N_8263);
and U12675 (N_12675,N_7145,N_9728);
nor U12676 (N_12676,N_6673,N_9379);
or U12677 (N_12677,N_5646,N_5334);
and U12678 (N_12678,N_6404,N_5507);
nand U12679 (N_12679,N_9186,N_5065);
nand U12680 (N_12680,N_8654,N_7154);
nor U12681 (N_12681,N_7600,N_6651);
and U12682 (N_12682,N_7959,N_5305);
nor U12683 (N_12683,N_8047,N_5610);
nor U12684 (N_12684,N_5078,N_6948);
nand U12685 (N_12685,N_9827,N_6530);
and U12686 (N_12686,N_6482,N_7024);
or U12687 (N_12687,N_7577,N_7900);
or U12688 (N_12688,N_6180,N_9317);
or U12689 (N_12689,N_9755,N_5897);
nand U12690 (N_12690,N_7810,N_8344);
or U12691 (N_12691,N_5150,N_8849);
nor U12692 (N_12692,N_5893,N_9969);
nor U12693 (N_12693,N_6844,N_7532);
nand U12694 (N_12694,N_7269,N_6165);
or U12695 (N_12695,N_6103,N_5497);
nand U12696 (N_12696,N_6146,N_6485);
or U12697 (N_12697,N_9532,N_9112);
nand U12698 (N_12698,N_7504,N_7491);
nand U12699 (N_12699,N_8669,N_8780);
nor U12700 (N_12700,N_8297,N_5724);
and U12701 (N_12701,N_5480,N_7695);
and U12702 (N_12702,N_6948,N_6604);
and U12703 (N_12703,N_5414,N_5364);
nand U12704 (N_12704,N_9187,N_9669);
nor U12705 (N_12705,N_8834,N_7575);
nand U12706 (N_12706,N_6955,N_9836);
nor U12707 (N_12707,N_7231,N_8287);
or U12708 (N_12708,N_6221,N_6562);
and U12709 (N_12709,N_9589,N_6391);
nor U12710 (N_12710,N_9143,N_6226);
nand U12711 (N_12711,N_5807,N_6290);
or U12712 (N_12712,N_7934,N_6837);
and U12713 (N_12713,N_9022,N_6232);
nand U12714 (N_12714,N_5671,N_9249);
and U12715 (N_12715,N_9961,N_9298);
nand U12716 (N_12716,N_7207,N_9834);
nand U12717 (N_12717,N_5711,N_7697);
or U12718 (N_12718,N_9540,N_6150);
nand U12719 (N_12719,N_5289,N_9033);
and U12720 (N_12720,N_9964,N_9820);
and U12721 (N_12721,N_8362,N_8553);
and U12722 (N_12722,N_7452,N_9292);
or U12723 (N_12723,N_9428,N_9706);
and U12724 (N_12724,N_9526,N_7140);
nor U12725 (N_12725,N_5749,N_6367);
nor U12726 (N_12726,N_9236,N_6236);
nor U12727 (N_12727,N_6143,N_8297);
or U12728 (N_12728,N_5485,N_9271);
or U12729 (N_12729,N_7101,N_5323);
nand U12730 (N_12730,N_5160,N_7859);
nor U12731 (N_12731,N_6760,N_9055);
or U12732 (N_12732,N_5902,N_7964);
nor U12733 (N_12733,N_9221,N_6349);
nor U12734 (N_12734,N_8832,N_7255);
nor U12735 (N_12735,N_5497,N_8064);
and U12736 (N_12736,N_6411,N_5897);
or U12737 (N_12737,N_5617,N_6288);
nand U12738 (N_12738,N_9313,N_7926);
xnor U12739 (N_12739,N_6939,N_7563);
nor U12740 (N_12740,N_8353,N_6120);
nor U12741 (N_12741,N_5630,N_8656);
nand U12742 (N_12742,N_8219,N_7215);
or U12743 (N_12743,N_5654,N_9338);
or U12744 (N_12744,N_6706,N_9542);
nand U12745 (N_12745,N_9587,N_5623);
and U12746 (N_12746,N_5654,N_8215);
nand U12747 (N_12747,N_8558,N_8965);
or U12748 (N_12748,N_5978,N_9990);
nand U12749 (N_12749,N_8831,N_5411);
nand U12750 (N_12750,N_8596,N_9736);
and U12751 (N_12751,N_9828,N_8633);
nand U12752 (N_12752,N_5387,N_6923);
nor U12753 (N_12753,N_9583,N_9394);
nand U12754 (N_12754,N_5238,N_9729);
nor U12755 (N_12755,N_7030,N_5027);
or U12756 (N_12756,N_7539,N_6352);
nand U12757 (N_12757,N_7435,N_9489);
nand U12758 (N_12758,N_8927,N_5882);
xor U12759 (N_12759,N_7829,N_6545);
or U12760 (N_12760,N_8332,N_8992);
nand U12761 (N_12761,N_9495,N_8460);
and U12762 (N_12762,N_5592,N_6805);
nor U12763 (N_12763,N_6007,N_9724);
nand U12764 (N_12764,N_7169,N_5933);
and U12765 (N_12765,N_8526,N_6777);
nand U12766 (N_12766,N_9621,N_8862);
or U12767 (N_12767,N_6544,N_8642);
xnor U12768 (N_12768,N_9501,N_5804);
nand U12769 (N_12769,N_9826,N_6974);
and U12770 (N_12770,N_8417,N_7408);
nor U12771 (N_12771,N_9406,N_6598);
nand U12772 (N_12772,N_8071,N_8833);
nand U12773 (N_12773,N_5554,N_7979);
nor U12774 (N_12774,N_6951,N_8570);
nand U12775 (N_12775,N_6056,N_9724);
and U12776 (N_12776,N_6651,N_5236);
nand U12777 (N_12777,N_5032,N_9953);
nor U12778 (N_12778,N_6802,N_7161);
nand U12779 (N_12779,N_9300,N_6882);
nand U12780 (N_12780,N_8274,N_8482);
nand U12781 (N_12781,N_7473,N_6174);
nand U12782 (N_12782,N_5296,N_5369);
nand U12783 (N_12783,N_8063,N_9441);
and U12784 (N_12784,N_7650,N_8109);
nor U12785 (N_12785,N_6184,N_7254);
xnor U12786 (N_12786,N_7180,N_6091);
nor U12787 (N_12787,N_9608,N_6095);
nor U12788 (N_12788,N_7847,N_6836);
or U12789 (N_12789,N_9703,N_9756);
nand U12790 (N_12790,N_6216,N_5168);
or U12791 (N_12791,N_6316,N_7006);
xnor U12792 (N_12792,N_7543,N_5494);
or U12793 (N_12793,N_7018,N_8344);
or U12794 (N_12794,N_9596,N_8923);
nand U12795 (N_12795,N_5878,N_7193);
and U12796 (N_12796,N_6481,N_7759);
nor U12797 (N_12797,N_6354,N_5750);
nand U12798 (N_12798,N_7079,N_9427);
nor U12799 (N_12799,N_9321,N_8252);
xnor U12800 (N_12800,N_9222,N_7736);
nor U12801 (N_12801,N_6210,N_8180);
or U12802 (N_12802,N_9964,N_7809);
xor U12803 (N_12803,N_8429,N_6936);
nand U12804 (N_12804,N_6205,N_5391);
or U12805 (N_12805,N_8944,N_7862);
nand U12806 (N_12806,N_7304,N_8744);
nor U12807 (N_12807,N_6951,N_5834);
nand U12808 (N_12808,N_9863,N_6444);
nor U12809 (N_12809,N_7694,N_9112);
and U12810 (N_12810,N_9883,N_9050);
or U12811 (N_12811,N_9983,N_7218);
and U12812 (N_12812,N_7873,N_9425);
nor U12813 (N_12813,N_9917,N_7407);
nor U12814 (N_12814,N_8236,N_5155);
nand U12815 (N_12815,N_7001,N_6778);
or U12816 (N_12816,N_5820,N_7011);
and U12817 (N_12817,N_8504,N_5903);
or U12818 (N_12818,N_8877,N_5005);
nand U12819 (N_12819,N_5582,N_8273);
and U12820 (N_12820,N_5424,N_8374);
nor U12821 (N_12821,N_9699,N_9697);
nor U12822 (N_12822,N_7320,N_9542);
nor U12823 (N_12823,N_7296,N_5249);
and U12824 (N_12824,N_5977,N_7305);
or U12825 (N_12825,N_9748,N_6348);
and U12826 (N_12826,N_6181,N_6786);
and U12827 (N_12827,N_7607,N_5178);
nor U12828 (N_12828,N_5002,N_5205);
and U12829 (N_12829,N_7455,N_6442);
or U12830 (N_12830,N_5386,N_8522);
and U12831 (N_12831,N_5525,N_6877);
xnor U12832 (N_12832,N_7008,N_9612);
or U12833 (N_12833,N_7349,N_5209);
nand U12834 (N_12834,N_5280,N_6277);
nand U12835 (N_12835,N_8973,N_9864);
nand U12836 (N_12836,N_8120,N_9926);
or U12837 (N_12837,N_6445,N_8177);
and U12838 (N_12838,N_6425,N_6938);
nand U12839 (N_12839,N_8453,N_9683);
nor U12840 (N_12840,N_5307,N_8368);
nand U12841 (N_12841,N_8512,N_7105);
and U12842 (N_12842,N_8427,N_8650);
or U12843 (N_12843,N_8195,N_8548);
and U12844 (N_12844,N_8369,N_5330);
nand U12845 (N_12845,N_6221,N_6185);
nand U12846 (N_12846,N_5155,N_9546);
nand U12847 (N_12847,N_8506,N_5728);
nor U12848 (N_12848,N_8828,N_7022);
nor U12849 (N_12849,N_8157,N_9511);
or U12850 (N_12850,N_7749,N_8913);
or U12851 (N_12851,N_5154,N_7989);
and U12852 (N_12852,N_9886,N_5949);
nand U12853 (N_12853,N_7911,N_9588);
nand U12854 (N_12854,N_9333,N_6158);
nand U12855 (N_12855,N_7339,N_6394);
nor U12856 (N_12856,N_7332,N_8853);
xnor U12857 (N_12857,N_7983,N_6319);
or U12858 (N_12858,N_6090,N_8851);
or U12859 (N_12859,N_5752,N_9746);
or U12860 (N_12860,N_7457,N_8711);
nand U12861 (N_12861,N_6644,N_8142);
and U12862 (N_12862,N_8985,N_9339);
or U12863 (N_12863,N_5335,N_5224);
nor U12864 (N_12864,N_8869,N_7118);
and U12865 (N_12865,N_8114,N_6066);
and U12866 (N_12866,N_6714,N_9566);
nor U12867 (N_12867,N_6067,N_5452);
nand U12868 (N_12868,N_7626,N_5149);
or U12869 (N_12869,N_9994,N_9933);
and U12870 (N_12870,N_9366,N_9604);
nand U12871 (N_12871,N_7503,N_5334);
nor U12872 (N_12872,N_7164,N_6648);
or U12873 (N_12873,N_6632,N_5836);
and U12874 (N_12874,N_9254,N_9057);
xnor U12875 (N_12875,N_8413,N_7061);
or U12876 (N_12876,N_8020,N_5005);
and U12877 (N_12877,N_9621,N_5052);
nand U12878 (N_12878,N_6368,N_5075);
nor U12879 (N_12879,N_7389,N_6548);
nand U12880 (N_12880,N_6643,N_5145);
nand U12881 (N_12881,N_6928,N_6496);
and U12882 (N_12882,N_9779,N_9034);
and U12883 (N_12883,N_7875,N_5842);
and U12884 (N_12884,N_9958,N_8330);
nand U12885 (N_12885,N_9006,N_7564);
nand U12886 (N_12886,N_6649,N_9461);
nor U12887 (N_12887,N_7660,N_8118);
and U12888 (N_12888,N_6015,N_9450);
nor U12889 (N_12889,N_5640,N_5420);
nor U12890 (N_12890,N_8145,N_7510);
nor U12891 (N_12891,N_8907,N_6959);
nand U12892 (N_12892,N_9202,N_9324);
or U12893 (N_12893,N_5617,N_5098);
nor U12894 (N_12894,N_8028,N_8258);
nor U12895 (N_12895,N_6130,N_9821);
and U12896 (N_12896,N_9341,N_9313);
or U12897 (N_12897,N_5245,N_9676);
and U12898 (N_12898,N_8271,N_8679);
nand U12899 (N_12899,N_8755,N_5920);
nand U12900 (N_12900,N_8821,N_7027);
or U12901 (N_12901,N_5701,N_8045);
nand U12902 (N_12902,N_9926,N_8981);
xnor U12903 (N_12903,N_9779,N_8016);
nand U12904 (N_12904,N_9977,N_9428);
xor U12905 (N_12905,N_5131,N_6478);
and U12906 (N_12906,N_5655,N_8316);
nor U12907 (N_12907,N_6696,N_8888);
xnor U12908 (N_12908,N_6837,N_8474);
nand U12909 (N_12909,N_9441,N_8401);
or U12910 (N_12910,N_7536,N_8625);
and U12911 (N_12911,N_8006,N_7675);
and U12912 (N_12912,N_5836,N_8439);
and U12913 (N_12913,N_9460,N_7256);
nand U12914 (N_12914,N_6700,N_9712);
and U12915 (N_12915,N_5919,N_6876);
or U12916 (N_12916,N_6055,N_5380);
or U12917 (N_12917,N_8754,N_8368);
or U12918 (N_12918,N_8998,N_5725);
or U12919 (N_12919,N_6602,N_8779);
nor U12920 (N_12920,N_5258,N_9092);
nand U12921 (N_12921,N_7245,N_7490);
or U12922 (N_12922,N_5857,N_9197);
and U12923 (N_12923,N_9183,N_6879);
nand U12924 (N_12924,N_7539,N_5757);
nand U12925 (N_12925,N_9881,N_6348);
nand U12926 (N_12926,N_8819,N_7557);
nor U12927 (N_12927,N_7322,N_9827);
or U12928 (N_12928,N_8543,N_7653);
xor U12929 (N_12929,N_8284,N_7710);
and U12930 (N_12930,N_7354,N_6999);
nand U12931 (N_12931,N_5061,N_8280);
and U12932 (N_12932,N_8680,N_5849);
nand U12933 (N_12933,N_5828,N_8020);
or U12934 (N_12934,N_9299,N_7171);
or U12935 (N_12935,N_9549,N_9233);
or U12936 (N_12936,N_5710,N_8097);
nand U12937 (N_12937,N_5413,N_5829);
or U12938 (N_12938,N_7350,N_5082);
or U12939 (N_12939,N_9542,N_5681);
or U12940 (N_12940,N_9638,N_9410);
or U12941 (N_12941,N_7358,N_5332);
or U12942 (N_12942,N_6203,N_6244);
or U12943 (N_12943,N_6448,N_9216);
or U12944 (N_12944,N_9980,N_6141);
nor U12945 (N_12945,N_7343,N_6467);
nor U12946 (N_12946,N_7962,N_7493);
nand U12947 (N_12947,N_8935,N_5910);
or U12948 (N_12948,N_5585,N_5801);
nor U12949 (N_12949,N_8121,N_7397);
nor U12950 (N_12950,N_5155,N_9794);
and U12951 (N_12951,N_5280,N_7741);
and U12952 (N_12952,N_5061,N_7231);
nor U12953 (N_12953,N_7923,N_6959);
or U12954 (N_12954,N_9016,N_9189);
nor U12955 (N_12955,N_7987,N_7137);
nand U12956 (N_12956,N_6864,N_7941);
and U12957 (N_12957,N_6686,N_9521);
nand U12958 (N_12958,N_8060,N_8408);
or U12959 (N_12959,N_5958,N_9677);
nand U12960 (N_12960,N_8014,N_8386);
nor U12961 (N_12961,N_5386,N_8542);
nand U12962 (N_12962,N_5653,N_9477);
nor U12963 (N_12963,N_9249,N_6244);
xnor U12964 (N_12964,N_9594,N_7216);
nand U12965 (N_12965,N_5519,N_8742);
nand U12966 (N_12966,N_7475,N_9101);
nand U12967 (N_12967,N_7158,N_9817);
nand U12968 (N_12968,N_6038,N_5101);
nand U12969 (N_12969,N_9267,N_5650);
nand U12970 (N_12970,N_9478,N_7881);
or U12971 (N_12971,N_5165,N_5790);
xor U12972 (N_12972,N_6686,N_6462);
nand U12973 (N_12973,N_8075,N_6214);
or U12974 (N_12974,N_8649,N_5737);
nand U12975 (N_12975,N_8866,N_6890);
nor U12976 (N_12976,N_8202,N_7231);
nor U12977 (N_12977,N_6452,N_8261);
or U12978 (N_12978,N_5296,N_8201);
nand U12979 (N_12979,N_8438,N_8429);
or U12980 (N_12980,N_5029,N_6565);
nor U12981 (N_12981,N_5679,N_6841);
nand U12982 (N_12982,N_7678,N_5820);
nor U12983 (N_12983,N_9595,N_6548);
and U12984 (N_12984,N_9476,N_7529);
or U12985 (N_12985,N_8428,N_7754);
and U12986 (N_12986,N_5486,N_7042);
or U12987 (N_12987,N_8857,N_7919);
or U12988 (N_12988,N_9861,N_9657);
nor U12989 (N_12989,N_8839,N_8069);
nand U12990 (N_12990,N_5120,N_5742);
nand U12991 (N_12991,N_7071,N_6180);
and U12992 (N_12992,N_7462,N_5783);
nor U12993 (N_12993,N_7533,N_5233);
and U12994 (N_12994,N_7442,N_6322);
nor U12995 (N_12995,N_9032,N_5554);
nand U12996 (N_12996,N_8186,N_5853);
and U12997 (N_12997,N_5556,N_6850);
nand U12998 (N_12998,N_8265,N_5225);
nor U12999 (N_12999,N_8310,N_9574);
and U13000 (N_13000,N_8622,N_9600);
nor U13001 (N_13001,N_6267,N_5260);
nor U13002 (N_13002,N_6482,N_7970);
and U13003 (N_13003,N_7714,N_8817);
or U13004 (N_13004,N_6408,N_9562);
nand U13005 (N_13005,N_5438,N_6958);
and U13006 (N_13006,N_7842,N_6454);
and U13007 (N_13007,N_7807,N_6697);
nand U13008 (N_13008,N_5947,N_6086);
xor U13009 (N_13009,N_9258,N_7730);
or U13010 (N_13010,N_7688,N_8849);
and U13011 (N_13011,N_9670,N_5269);
or U13012 (N_13012,N_5440,N_6173);
nor U13013 (N_13013,N_8612,N_6977);
or U13014 (N_13014,N_8524,N_7651);
and U13015 (N_13015,N_7802,N_7441);
nor U13016 (N_13016,N_6482,N_5220);
or U13017 (N_13017,N_6055,N_5404);
xnor U13018 (N_13018,N_8707,N_8904);
or U13019 (N_13019,N_8383,N_9470);
nand U13020 (N_13020,N_9654,N_9789);
and U13021 (N_13021,N_9624,N_8528);
and U13022 (N_13022,N_5778,N_7921);
nand U13023 (N_13023,N_8182,N_9579);
nand U13024 (N_13024,N_6095,N_5126);
and U13025 (N_13025,N_5242,N_7711);
and U13026 (N_13026,N_9750,N_9120);
nand U13027 (N_13027,N_9643,N_8017);
nor U13028 (N_13028,N_9946,N_8254);
nor U13029 (N_13029,N_9905,N_9839);
nand U13030 (N_13030,N_7308,N_8207);
and U13031 (N_13031,N_6471,N_7078);
or U13032 (N_13032,N_6108,N_7953);
or U13033 (N_13033,N_5999,N_6001);
nor U13034 (N_13034,N_5970,N_5842);
nand U13035 (N_13035,N_6496,N_9429);
or U13036 (N_13036,N_9716,N_9310);
nand U13037 (N_13037,N_9523,N_7200);
nand U13038 (N_13038,N_9978,N_9182);
nor U13039 (N_13039,N_7159,N_8431);
or U13040 (N_13040,N_9282,N_6051);
nand U13041 (N_13041,N_7252,N_5154);
or U13042 (N_13042,N_9629,N_9384);
and U13043 (N_13043,N_5336,N_9116);
and U13044 (N_13044,N_9121,N_9791);
and U13045 (N_13045,N_6795,N_7563);
and U13046 (N_13046,N_7203,N_7182);
nor U13047 (N_13047,N_6999,N_6234);
and U13048 (N_13048,N_6662,N_5659);
and U13049 (N_13049,N_8616,N_8260);
and U13050 (N_13050,N_5892,N_9346);
xnor U13051 (N_13051,N_8755,N_7676);
nor U13052 (N_13052,N_9852,N_7304);
nor U13053 (N_13053,N_5458,N_9670);
or U13054 (N_13054,N_5011,N_5830);
nand U13055 (N_13055,N_9921,N_8945);
nand U13056 (N_13056,N_7287,N_8574);
or U13057 (N_13057,N_8152,N_9494);
nor U13058 (N_13058,N_8348,N_8833);
or U13059 (N_13059,N_8484,N_8252);
nand U13060 (N_13060,N_7002,N_6085);
and U13061 (N_13061,N_7056,N_8965);
or U13062 (N_13062,N_6255,N_7688);
nand U13063 (N_13063,N_6964,N_6214);
nor U13064 (N_13064,N_5664,N_5111);
and U13065 (N_13065,N_6314,N_9141);
xor U13066 (N_13066,N_8835,N_7376);
nor U13067 (N_13067,N_9855,N_5136);
nor U13068 (N_13068,N_7838,N_5091);
and U13069 (N_13069,N_9713,N_8084);
nor U13070 (N_13070,N_5174,N_9617);
nand U13071 (N_13071,N_5295,N_9450);
and U13072 (N_13072,N_5046,N_8549);
or U13073 (N_13073,N_6685,N_8048);
nand U13074 (N_13074,N_7929,N_6898);
and U13075 (N_13075,N_6130,N_7491);
or U13076 (N_13076,N_7645,N_6346);
nor U13077 (N_13077,N_6941,N_7965);
and U13078 (N_13078,N_6710,N_9713);
or U13079 (N_13079,N_9591,N_5974);
or U13080 (N_13080,N_8260,N_6876);
nor U13081 (N_13081,N_8444,N_5446);
or U13082 (N_13082,N_6533,N_9311);
or U13083 (N_13083,N_9627,N_8218);
and U13084 (N_13084,N_6110,N_5258);
or U13085 (N_13085,N_8567,N_5950);
nor U13086 (N_13086,N_5229,N_9365);
nand U13087 (N_13087,N_8879,N_9012);
nand U13088 (N_13088,N_5066,N_9907);
and U13089 (N_13089,N_7036,N_5679);
nand U13090 (N_13090,N_9657,N_8571);
nor U13091 (N_13091,N_8264,N_6490);
xnor U13092 (N_13092,N_9019,N_7155);
and U13093 (N_13093,N_8958,N_8734);
nand U13094 (N_13094,N_8072,N_8116);
and U13095 (N_13095,N_5627,N_5535);
xnor U13096 (N_13096,N_7747,N_8806);
nand U13097 (N_13097,N_9818,N_8022);
or U13098 (N_13098,N_8713,N_8747);
xor U13099 (N_13099,N_8597,N_6088);
xor U13100 (N_13100,N_6624,N_9078);
or U13101 (N_13101,N_9313,N_7039);
and U13102 (N_13102,N_9163,N_7463);
or U13103 (N_13103,N_6480,N_8508);
or U13104 (N_13104,N_9913,N_5057);
or U13105 (N_13105,N_6625,N_5761);
nor U13106 (N_13106,N_5394,N_8277);
nor U13107 (N_13107,N_8836,N_5636);
or U13108 (N_13108,N_8754,N_6456);
nand U13109 (N_13109,N_7667,N_9602);
or U13110 (N_13110,N_6571,N_6096);
or U13111 (N_13111,N_9357,N_5993);
and U13112 (N_13112,N_6690,N_8780);
nor U13113 (N_13113,N_8106,N_8049);
or U13114 (N_13114,N_9140,N_7713);
and U13115 (N_13115,N_9288,N_6046);
nor U13116 (N_13116,N_8054,N_9318);
or U13117 (N_13117,N_7858,N_8165);
or U13118 (N_13118,N_8531,N_9179);
nor U13119 (N_13119,N_5050,N_8471);
nand U13120 (N_13120,N_9409,N_7511);
nor U13121 (N_13121,N_8043,N_5349);
and U13122 (N_13122,N_5499,N_7079);
nor U13123 (N_13123,N_6570,N_9705);
or U13124 (N_13124,N_5810,N_8410);
or U13125 (N_13125,N_9082,N_6623);
and U13126 (N_13126,N_5657,N_9930);
or U13127 (N_13127,N_7309,N_6725);
nand U13128 (N_13128,N_7459,N_5786);
nand U13129 (N_13129,N_5863,N_6961);
or U13130 (N_13130,N_8416,N_6594);
or U13131 (N_13131,N_9388,N_7258);
nor U13132 (N_13132,N_5347,N_9203);
xor U13133 (N_13133,N_8096,N_6859);
nor U13134 (N_13134,N_8565,N_7765);
nor U13135 (N_13135,N_9313,N_8167);
and U13136 (N_13136,N_7617,N_7753);
and U13137 (N_13137,N_7419,N_5756);
and U13138 (N_13138,N_9118,N_7429);
nor U13139 (N_13139,N_7006,N_8333);
and U13140 (N_13140,N_6770,N_5716);
nor U13141 (N_13141,N_7687,N_5975);
or U13142 (N_13142,N_6852,N_8231);
nor U13143 (N_13143,N_8315,N_9895);
and U13144 (N_13144,N_8811,N_5683);
and U13145 (N_13145,N_9923,N_9504);
nor U13146 (N_13146,N_7811,N_9807);
and U13147 (N_13147,N_7253,N_7709);
nand U13148 (N_13148,N_9403,N_7820);
nor U13149 (N_13149,N_9585,N_8815);
and U13150 (N_13150,N_8305,N_9979);
nor U13151 (N_13151,N_8886,N_7927);
nor U13152 (N_13152,N_7156,N_6578);
or U13153 (N_13153,N_5232,N_8287);
nor U13154 (N_13154,N_6699,N_8544);
nand U13155 (N_13155,N_7085,N_7216);
nor U13156 (N_13156,N_9159,N_6524);
xor U13157 (N_13157,N_6590,N_9431);
or U13158 (N_13158,N_9164,N_8299);
nor U13159 (N_13159,N_8138,N_5644);
or U13160 (N_13160,N_8622,N_5907);
or U13161 (N_13161,N_9786,N_9404);
nor U13162 (N_13162,N_9647,N_6307);
nor U13163 (N_13163,N_8005,N_7219);
nor U13164 (N_13164,N_5059,N_6067);
nand U13165 (N_13165,N_6365,N_6776);
nor U13166 (N_13166,N_6646,N_9037);
and U13167 (N_13167,N_5886,N_7074);
xor U13168 (N_13168,N_9592,N_6865);
xor U13169 (N_13169,N_5084,N_5890);
or U13170 (N_13170,N_7726,N_7292);
and U13171 (N_13171,N_8961,N_5453);
and U13172 (N_13172,N_8780,N_7500);
or U13173 (N_13173,N_8480,N_9082);
and U13174 (N_13174,N_5995,N_9247);
or U13175 (N_13175,N_5411,N_9707);
nor U13176 (N_13176,N_7317,N_8985);
and U13177 (N_13177,N_6953,N_8569);
and U13178 (N_13178,N_6364,N_7597);
nand U13179 (N_13179,N_6769,N_7232);
and U13180 (N_13180,N_6201,N_5977);
and U13181 (N_13181,N_7341,N_9290);
and U13182 (N_13182,N_9667,N_8255);
and U13183 (N_13183,N_5333,N_8195);
nor U13184 (N_13184,N_9934,N_5690);
nor U13185 (N_13185,N_7757,N_6896);
and U13186 (N_13186,N_6613,N_8605);
and U13187 (N_13187,N_8977,N_9162);
nor U13188 (N_13188,N_6414,N_7911);
nand U13189 (N_13189,N_8732,N_6546);
nand U13190 (N_13190,N_6683,N_6888);
nor U13191 (N_13191,N_9844,N_9132);
nor U13192 (N_13192,N_6769,N_9650);
nor U13193 (N_13193,N_8821,N_5926);
and U13194 (N_13194,N_9435,N_8573);
nand U13195 (N_13195,N_5932,N_9837);
and U13196 (N_13196,N_8957,N_7774);
and U13197 (N_13197,N_8174,N_9704);
xor U13198 (N_13198,N_9844,N_6050);
nor U13199 (N_13199,N_8760,N_8090);
xor U13200 (N_13200,N_5524,N_9128);
nor U13201 (N_13201,N_8935,N_6531);
nor U13202 (N_13202,N_6904,N_8674);
xnor U13203 (N_13203,N_7617,N_8393);
or U13204 (N_13204,N_7490,N_6847);
nand U13205 (N_13205,N_6747,N_9617);
nand U13206 (N_13206,N_6307,N_9702);
nand U13207 (N_13207,N_8563,N_5318);
nor U13208 (N_13208,N_7315,N_7152);
nor U13209 (N_13209,N_6183,N_9537);
or U13210 (N_13210,N_9256,N_5628);
nand U13211 (N_13211,N_8561,N_5038);
nand U13212 (N_13212,N_6805,N_5867);
and U13213 (N_13213,N_7784,N_7965);
or U13214 (N_13214,N_6697,N_5303);
xor U13215 (N_13215,N_7040,N_9350);
nor U13216 (N_13216,N_6110,N_9417);
nand U13217 (N_13217,N_6656,N_6342);
or U13218 (N_13218,N_6659,N_6121);
nor U13219 (N_13219,N_9784,N_8560);
and U13220 (N_13220,N_7151,N_8673);
and U13221 (N_13221,N_8695,N_5549);
and U13222 (N_13222,N_9641,N_5178);
nand U13223 (N_13223,N_7105,N_8016);
or U13224 (N_13224,N_7182,N_8893);
and U13225 (N_13225,N_9661,N_8202);
nor U13226 (N_13226,N_9806,N_5766);
and U13227 (N_13227,N_9102,N_7370);
nand U13228 (N_13228,N_9779,N_8374);
nand U13229 (N_13229,N_9442,N_8949);
nor U13230 (N_13230,N_7481,N_7953);
and U13231 (N_13231,N_7608,N_6484);
and U13232 (N_13232,N_9882,N_8741);
nand U13233 (N_13233,N_9982,N_6713);
nand U13234 (N_13234,N_5995,N_6732);
nor U13235 (N_13235,N_9819,N_7497);
or U13236 (N_13236,N_7133,N_9642);
xnor U13237 (N_13237,N_8921,N_6151);
nor U13238 (N_13238,N_9104,N_8697);
nor U13239 (N_13239,N_7883,N_9673);
and U13240 (N_13240,N_8219,N_5998);
or U13241 (N_13241,N_5207,N_7040);
nand U13242 (N_13242,N_6840,N_7522);
nand U13243 (N_13243,N_8695,N_6151);
nand U13244 (N_13244,N_6337,N_8563);
nand U13245 (N_13245,N_7103,N_5820);
nor U13246 (N_13246,N_6980,N_8591);
nand U13247 (N_13247,N_5132,N_7495);
or U13248 (N_13248,N_8983,N_6865);
nand U13249 (N_13249,N_6180,N_8883);
or U13250 (N_13250,N_9414,N_8852);
or U13251 (N_13251,N_7315,N_8133);
and U13252 (N_13252,N_7425,N_8772);
or U13253 (N_13253,N_8269,N_6372);
and U13254 (N_13254,N_7081,N_6636);
and U13255 (N_13255,N_6849,N_9327);
or U13256 (N_13256,N_7588,N_8986);
nand U13257 (N_13257,N_6119,N_6326);
and U13258 (N_13258,N_9049,N_8352);
or U13259 (N_13259,N_6959,N_6230);
or U13260 (N_13260,N_8960,N_5916);
and U13261 (N_13261,N_6706,N_9324);
or U13262 (N_13262,N_8475,N_9629);
xnor U13263 (N_13263,N_6218,N_6117);
or U13264 (N_13264,N_7703,N_9064);
or U13265 (N_13265,N_5147,N_9666);
and U13266 (N_13266,N_5342,N_7808);
or U13267 (N_13267,N_7683,N_9380);
nor U13268 (N_13268,N_8063,N_5677);
and U13269 (N_13269,N_6683,N_5303);
or U13270 (N_13270,N_8757,N_6783);
or U13271 (N_13271,N_8406,N_8977);
nor U13272 (N_13272,N_8748,N_8036);
or U13273 (N_13273,N_6825,N_9464);
nand U13274 (N_13274,N_9913,N_7511);
or U13275 (N_13275,N_9116,N_5059);
or U13276 (N_13276,N_8553,N_7838);
nand U13277 (N_13277,N_6232,N_6526);
nand U13278 (N_13278,N_9997,N_6986);
nor U13279 (N_13279,N_8078,N_7241);
or U13280 (N_13280,N_9763,N_6233);
nand U13281 (N_13281,N_9959,N_7154);
nor U13282 (N_13282,N_8548,N_7870);
nand U13283 (N_13283,N_5040,N_5379);
or U13284 (N_13284,N_5433,N_6466);
nand U13285 (N_13285,N_5701,N_8199);
and U13286 (N_13286,N_6346,N_8586);
nor U13287 (N_13287,N_7405,N_9347);
and U13288 (N_13288,N_8093,N_8347);
and U13289 (N_13289,N_8814,N_9106);
and U13290 (N_13290,N_7399,N_8168);
or U13291 (N_13291,N_8857,N_5041);
nor U13292 (N_13292,N_9038,N_9617);
and U13293 (N_13293,N_6183,N_8376);
nor U13294 (N_13294,N_7997,N_6492);
or U13295 (N_13295,N_5034,N_6219);
or U13296 (N_13296,N_7645,N_5778);
and U13297 (N_13297,N_8677,N_6303);
nand U13298 (N_13298,N_8130,N_5875);
nand U13299 (N_13299,N_9973,N_7665);
and U13300 (N_13300,N_8083,N_7546);
nand U13301 (N_13301,N_9794,N_6712);
nor U13302 (N_13302,N_9195,N_9288);
nand U13303 (N_13303,N_8090,N_9855);
nor U13304 (N_13304,N_7170,N_7764);
and U13305 (N_13305,N_9150,N_8466);
nand U13306 (N_13306,N_8671,N_6835);
or U13307 (N_13307,N_8143,N_6457);
nand U13308 (N_13308,N_9255,N_5720);
nand U13309 (N_13309,N_7283,N_8593);
or U13310 (N_13310,N_5645,N_8020);
or U13311 (N_13311,N_8416,N_6968);
nor U13312 (N_13312,N_9152,N_5587);
nor U13313 (N_13313,N_9864,N_7408);
nor U13314 (N_13314,N_6630,N_5614);
nand U13315 (N_13315,N_6643,N_7562);
or U13316 (N_13316,N_6559,N_5413);
xor U13317 (N_13317,N_7053,N_8763);
nand U13318 (N_13318,N_7416,N_8358);
nor U13319 (N_13319,N_9575,N_9279);
nand U13320 (N_13320,N_5603,N_7320);
and U13321 (N_13321,N_5489,N_5352);
nand U13322 (N_13322,N_8799,N_6484);
or U13323 (N_13323,N_5637,N_9885);
nor U13324 (N_13324,N_8599,N_7634);
nor U13325 (N_13325,N_9958,N_6971);
or U13326 (N_13326,N_8711,N_6443);
and U13327 (N_13327,N_8109,N_6149);
nand U13328 (N_13328,N_5009,N_6603);
and U13329 (N_13329,N_7805,N_6849);
and U13330 (N_13330,N_7239,N_7422);
and U13331 (N_13331,N_8261,N_5154);
nand U13332 (N_13332,N_7564,N_9446);
nor U13333 (N_13333,N_7158,N_7387);
nor U13334 (N_13334,N_5167,N_5978);
nor U13335 (N_13335,N_7067,N_7404);
and U13336 (N_13336,N_6813,N_7543);
or U13337 (N_13337,N_6574,N_9183);
and U13338 (N_13338,N_5791,N_7541);
and U13339 (N_13339,N_6170,N_6587);
nor U13340 (N_13340,N_6233,N_7564);
nor U13341 (N_13341,N_8431,N_6399);
and U13342 (N_13342,N_5819,N_6123);
nor U13343 (N_13343,N_6903,N_8487);
or U13344 (N_13344,N_7848,N_6719);
and U13345 (N_13345,N_8538,N_6085);
nand U13346 (N_13346,N_8270,N_9562);
nor U13347 (N_13347,N_8380,N_5804);
nor U13348 (N_13348,N_7672,N_5777);
nor U13349 (N_13349,N_6731,N_9313);
nor U13350 (N_13350,N_9363,N_5137);
or U13351 (N_13351,N_6834,N_8962);
or U13352 (N_13352,N_5810,N_9719);
and U13353 (N_13353,N_7929,N_6380);
and U13354 (N_13354,N_9745,N_6124);
and U13355 (N_13355,N_9149,N_6348);
and U13356 (N_13356,N_5971,N_9153);
and U13357 (N_13357,N_7997,N_5554);
nand U13358 (N_13358,N_6341,N_5855);
or U13359 (N_13359,N_6079,N_5620);
nor U13360 (N_13360,N_6509,N_9064);
and U13361 (N_13361,N_6011,N_5520);
or U13362 (N_13362,N_7694,N_9152);
or U13363 (N_13363,N_7805,N_8416);
nand U13364 (N_13364,N_7982,N_5681);
nor U13365 (N_13365,N_9177,N_8432);
nor U13366 (N_13366,N_7564,N_7804);
nor U13367 (N_13367,N_6031,N_9452);
and U13368 (N_13368,N_9464,N_8040);
and U13369 (N_13369,N_6357,N_8648);
or U13370 (N_13370,N_7192,N_8828);
nand U13371 (N_13371,N_8343,N_9779);
and U13372 (N_13372,N_7004,N_6950);
nand U13373 (N_13373,N_8427,N_5799);
nor U13374 (N_13374,N_5271,N_6420);
nor U13375 (N_13375,N_6018,N_6739);
or U13376 (N_13376,N_9694,N_9276);
nand U13377 (N_13377,N_5494,N_6773);
or U13378 (N_13378,N_9249,N_8783);
and U13379 (N_13379,N_6374,N_6122);
nand U13380 (N_13380,N_5684,N_8782);
nand U13381 (N_13381,N_7967,N_6690);
nor U13382 (N_13382,N_6054,N_7989);
nand U13383 (N_13383,N_5475,N_9125);
or U13384 (N_13384,N_5827,N_8766);
nand U13385 (N_13385,N_9891,N_8565);
or U13386 (N_13386,N_5334,N_7034);
or U13387 (N_13387,N_9069,N_5610);
nand U13388 (N_13388,N_6906,N_9339);
or U13389 (N_13389,N_9653,N_7256);
or U13390 (N_13390,N_5216,N_8733);
nor U13391 (N_13391,N_6934,N_9009);
and U13392 (N_13392,N_6928,N_7016);
nor U13393 (N_13393,N_5195,N_6977);
nor U13394 (N_13394,N_7034,N_9156);
nor U13395 (N_13395,N_9435,N_9868);
nor U13396 (N_13396,N_9864,N_9256);
nor U13397 (N_13397,N_7301,N_8165);
nor U13398 (N_13398,N_8627,N_7066);
nand U13399 (N_13399,N_9394,N_9823);
nand U13400 (N_13400,N_5662,N_8004);
and U13401 (N_13401,N_9546,N_9695);
or U13402 (N_13402,N_9960,N_6169);
and U13403 (N_13403,N_5265,N_7484);
or U13404 (N_13404,N_5851,N_9838);
and U13405 (N_13405,N_6005,N_5452);
or U13406 (N_13406,N_7618,N_5889);
and U13407 (N_13407,N_5666,N_5526);
and U13408 (N_13408,N_9282,N_9449);
nand U13409 (N_13409,N_8318,N_8059);
xnor U13410 (N_13410,N_6645,N_9889);
nor U13411 (N_13411,N_6411,N_5216);
or U13412 (N_13412,N_9834,N_8945);
or U13413 (N_13413,N_6999,N_5656);
and U13414 (N_13414,N_8923,N_6879);
and U13415 (N_13415,N_5567,N_9202);
nor U13416 (N_13416,N_9393,N_7782);
nor U13417 (N_13417,N_6699,N_8954);
nand U13418 (N_13418,N_7062,N_8136);
or U13419 (N_13419,N_6205,N_6849);
nor U13420 (N_13420,N_6001,N_9101);
or U13421 (N_13421,N_8747,N_5405);
nand U13422 (N_13422,N_8652,N_7927);
nand U13423 (N_13423,N_6280,N_7178);
or U13424 (N_13424,N_8728,N_6065);
nand U13425 (N_13425,N_7221,N_6583);
nand U13426 (N_13426,N_7637,N_6384);
nand U13427 (N_13427,N_5906,N_7626);
and U13428 (N_13428,N_7271,N_5440);
and U13429 (N_13429,N_7740,N_8415);
nor U13430 (N_13430,N_5182,N_7668);
nand U13431 (N_13431,N_8292,N_9915);
nand U13432 (N_13432,N_5602,N_6810);
and U13433 (N_13433,N_8015,N_9060);
nand U13434 (N_13434,N_6446,N_5439);
and U13435 (N_13435,N_7328,N_7095);
or U13436 (N_13436,N_8806,N_5632);
nand U13437 (N_13437,N_8810,N_9347);
and U13438 (N_13438,N_9626,N_6347);
nor U13439 (N_13439,N_6709,N_8218);
nor U13440 (N_13440,N_7496,N_6571);
or U13441 (N_13441,N_8311,N_5945);
nand U13442 (N_13442,N_9636,N_7212);
nor U13443 (N_13443,N_8071,N_7448);
or U13444 (N_13444,N_7708,N_8269);
nand U13445 (N_13445,N_8818,N_9060);
nor U13446 (N_13446,N_9908,N_8038);
or U13447 (N_13447,N_8906,N_7954);
or U13448 (N_13448,N_7299,N_9677);
nor U13449 (N_13449,N_7821,N_7753);
nor U13450 (N_13450,N_6892,N_9624);
or U13451 (N_13451,N_5863,N_8890);
nor U13452 (N_13452,N_7868,N_5584);
or U13453 (N_13453,N_6993,N_8273);
xnor U13454 (N_13454,N_6115,N_5322);
nor U13455 (N_13455,N_5286,N_8563);
or U13456 (N_13456,N_8602,N_6880);
nor U13457 (N_13457,N_5791,N_9698);
nor U13458 (N_13458,N_5597,N_7425);
or U13459 (N_13459,N_6689,N_5470);
nor U13460 (N_13460,N_5090,N_8065);
or U13461 (N_13461,N_7352,N_8093);
nor U13462 (N_13462,N_8621,N_5814);
nand U13463 (N_13463,N_8314,N_7792);
nor U13464 (N_13464,N_8119,N_9854);
or U13465 (N_13465,N_8690,N_6912);
and U13466 (N_13466,N_9860,N_9156);
and U13467 (N_13467,N_7028,N_8992);
or U13468 (N_13468,N_8545,N_5384);
or U13469 (N_13469,N_5453,N_5116);
nand U13470 (N_13470,N_7971,N_5107);
nor U13471 (N_13471,N_8953,N_8222);
nand U13472 (N_13472,N_6949,N_7580);
nand U13473 (N_13473,N_5018,N_7942);
nor U13474 (N_13474,N_6977,N_8571);
or U13475 (N_13475,N_8803,N_8083);
and U13476 (N_13476,N_8856,N_8861);
and U13477 (N_13477,N_7503,N_5180);
or U13478 (N_13478,N_5553,N_7437);
nor U13479 (N_13479,N_6259,N_8218);
and U13480 (N_13480,N_6302,N_6319);
nand U13481 (N_13481,N_8903,N_5306);
nor U13482 (N_13482,N_8606,N_8262);
or U13483 (N_13483,N_5816,N_5076);
and U13484 (N_13484,N_8048,N_5769);
and U13485 (N_13485,N_5639,N_7156);
and U13486 (N_13486,N_6397,N_5197);
nand U13487 (N_13487,N_6161,N_5517);
and U13488 (N_13488,N_9802,N_9818);
and U13489 (N_13489,N_8017,N_7650);
nor U13490 (N_13490,N_6829,N_5553);
nand U13491 (N_13491,N_9857,N_5852);
nand U13492 (N_13492,N_7399,N_9497);
nand U13493 (N_13493,N_7377,N_6747);
nor U13494 (N_13494,N_8256,N_6065);
or U13495 (N_13495,N_5541,N_8067);
nand U13496 (N_13496,N_7923,N_5423);
nand U13497 (N_13497,N_8358,N_7713);
and U13498 (N_13498,N_7369,N_9302);
or U13499 (N_13499,N_5133,N_6238);
nor U13500 (N_13500,N_5569,N_5643);
xor U13501 (N_13501,N_6460,N_6753);
nand U13502 (N_13502,N_5853,N_9965);
nor U13503 (N_13503,N_6720,N_7862);
and U13504 (N_13504,N_6139,N_5762);
and U13505 (N_13505,N_6262,N_5308);
and U13506 (N_13506,N_5581,N_6077);
and U13507 (N_13507,N_6642,N_8000);
nor U13508 (N_13508,N_9779,N_8017);
nor U13509 (N_13509,N_6043,N_9677);
nand U13510 (N_13510,N_8251,N_9295);
and U13511 (N_13511,N_5835,N_7889);
nand U13512 (N_13512,N_7399,N_7184);
xor U13513 (N_13513,N_7855,N_5104);
nor U13514 (N_13514,N_7396,N_8628);
nor U13515 (N_13515,N_7468,N_5011);
and U13516 (N_13516,N_6875,N_5570);
and U13517 (N_13517,N_8306,N_7818);
nor U13518 (N_13518,N_9592,N_5457);
and U13519 (N_13519,N_6855,N_5070);
and U13520 (N_13520,N_8116,N_6104);
nor U13521 (N_13521,N_6133,N_8398);
or U13522 (N_13522,N_7664,N_5589);
or U13523 (N_13523,N_5901,N_8317);
nor U13524 (N_13524,N_6487,N_6706);
nor U13525 (N_13525,N_9228,N_6563);
xnor U13526 (N_13526,N_9633,N_7197);
nand U13527 (N_13527,N_8957,N_5842);
nor U13528 (N_13528,N_8995,N_8429);
nor U13529 (N_13529,N_5984,N_9285);
nor U13530 (N_13530,N_9176,N_6003);
or U13531 (N_13531,N_7826,N_6364);
and U13532 (N_13532,N_5447,N_7218);
nor U13533 (N_13533,N_7155,N_8333);
nor U13534 (N_13534,N_6861,N_9022);
and U13535 (N_13535,N_9049,N_8542);
nand U13536 (N_13536,N_5616,N_8280);
or U13537 (N_13537,N_5752,N_9526);
and U13538 (N_13538,N_7569,N_6156);
and U13539 (N_13539,N_7837,N_7960);
nand U13540 (N_13540,N_9134,N_7871);
nor U13541 (N_13541,N_8914,N_6480);
or U13542 (N_13542,N_7479,N_5810);
and U13543 (N_13543,N_9590,N_6148);
nor U13544 (N_13544,N_5162,N_8517);
or U13545 (N_13545,N_6099,N_7490);
nand U13546 (N_13546,N_9807,N_6238);
and U13547 (N_13547,N_7620,N_5358);
or U13548 (N_13548,N_5992,N_5292);
xor U13549 (N_13549,N_9702,N_9109);
nor U13550 (N_13550,N_8503,N_7304);
nor U13551 (N_13551,N_6114,N_8877);
nor U13552 (N_13552,N_7492,N_5994);
and U13553 (N_13553,N_9282,N_6386);
nand U13554 (N_13554,N_7456,N_6415);
or U13555 (N_13555,N_9435,N_6630);
nand U13556 (N_13556,N_9702,N_7722);
nor U13557 (N_13557,N_9393,N_9389);
nand U13558 (N_13558,N_8586,N_9586);
or U13559 (N_13559,N_7554,N_9020);
nand U13560 (N_13560,N_8903,N_6015);
nor U13561 (N_13561,N_7692,N_6587);
or U13562 (N_13562,N_9248,N_5624);
and U13563 (N_13563,N_6856,N_7518);
and U13564 (N_13564,N_8941,N_7156);
and U13565 (N_13565,N_9137,N_6582);
and U13566 (N_13566,N_7311,N_6221);
or U13567 (N_13567,N_5176,N_9436);
and U13568 (N_13568,N_6028,N_7718);
or U13569 (N_13569,N_6241,N_5362);
and U13570 (N_13570,N_7761,N_8476);
nor U13571 (N_13571,N_5480,N_9534);
or U13572 (N_13572,N_7089,N_5198);
xnor U13573 (N_13573,N_9332,N_9539);
and U13574 (N_13574,N_5556,N_8923);
xor U13575 (N_13575,N_6953,N_6409);
or U13576 (N_13576,N_8611,N_7007);
or U13577 (N_13577,N_8069,N_8383);
and U13578 (N_13578,N_8866,N_8459);
nor U13579 (N_13579,N_5268,N_6209);
and U13580 (N_13580,N_6093,N_8832);
nor U13581 (N_13581,N_5847,N_9161);
nand U13582 (N_13582,N_6795,N_9832);
nor U13583 (N_13583,N_5794,N_9092);
xnor U13584 (N_13584,N_8862,N_6378);
or U13585 (N_13585,N_8092,N_8837);
nand U13586 (N_13586,N_8942,N_8017);
nor U13587 (N_13587,N_5015,N_5810);
xor U13588 (N_13588,N_7950,N_9134);
nor U13589 (N_13589,N_9790,N_9067);
or U13590 (N_13590,N_7644,N_7233);
nand U13591 (N_13591,N_6303,N_6824);
nor U13592 (N_13592,N_8883,N_5027);
or U13593 (N_13593,N_8073,N_8553);
nand U13594 (N_13594,N_6587,N_8679);
and U13595 (N_13595,N_9646,N_7474);
and U13596 (N_13596,N_8528,N_8937);
nor U13597 (N_13597,N_8866,N_5529);
and U13598 (N_13598,N_5535,N_8613);
nor U13599 (N_13599,N_7691,N_5741);
nand U13600 (N_13600,N_6139,N_6561);
or U13601 (N_13601,N_5504,N_8726);
nand U13602 (N_13602,N_9855,N_6767);
xnor U13603 (N_13603,N_7863,N_6237);
nand U13604 (N_13604,N_7755,N_8926);
nor U13605 (N_13605,N_9032,N_9488);
and U13606 (N_13606,N_6914,N_8576);
or U13607 (N_13607,N_9592,N_6298);
and U13608 (N_13608,N_9373,N_9888);
or U13609 (N_13609,N_9044,N_8304);
and U13610 (N_13610,N_8071,N_7388);
and U13611 (N_13611,N_7528,N_6981);
and U13612 (N_13612,N_6514,N_5248);
nand U13613 (N_13613,N_7227,N_5709);
nor U13614 (N_13614,N_8640,N_5638);
and U13615 (N_13615,N_7549,N_9725);
or U13616 (N_13616,N_5576,N_6508);
or U13617 (N_13617,N_7027,N_5321);
or U13618 (N_13618,N_7002,N_6071);
or U13619 (N_13619,N_7919,N_5932);
nand U13620 (N_13620,N_7956,N_8671);
nand U13621 (N_13621,N_8530,N_8384);
or U13622 (N_13622,N_7694,N_5239);
or U13623 (N_13623,N_7604,N_7599);
or U13624 (N_13624,N_7333,N_6143);
nor U13625 (N_13625,N_7994,N_6306);
nand U13626 (N_13626,N_8368,N_6894);
and U13627 (N_13627,N_5036,N_7331);
and U13628 (N_13628,N_5101,N_5378);
and U13629 (N_13629,N_8857,N_9163);
nor U13630 (N_13630,N_5384,N_7347);
nand U13631 (N_13631,N_5117,N_9697);
nor U13632 (N_13632,N_8558,N_9214);
nor U13633 (N_13633,N_8772,N_9141);
nand U13634 (N_13634,N_5007,N_5105);
or U13635 (N_13635,N_7619,N_7744);
xor U13636 (N_13636,N_8021,N_5578);
nand U13637 (N_13637,N_5798,N_7161);
xor U13638 (N_13638,N_7799,N_8945);
and U13639 (N_13639,N_5877,N_6123);
nand U13640 (N_13640,N_6422,N_6938);
nor U13641 (N_13641,N_8406,N_9156);
nor U13642 (N_13642,N_9262,N_7546);
nor U13643 (N_13643,N_8820,N_9312);
or U13644 (N_13644,N_8015,N_5628);
or U13645 (N_13645,N_9734,N_7133);
and U13646 (N_13646,N_6422,N_7491);
xor U13647 (N_13647,N_7382,N_9009);
and U13648 (N_13648,N_8572,N_7932);
xor U13649 (N_13649,N_5413,N_5770);
or U13650 (N_13650,N_9198,N_6610);
nand U13651 (N_13651,N_6242,N_7754);
or U13652 (N_13652,N_6217,N_9566);
nand U13653 (N_13653,N_9253,N_7809);
nand U13654 (N_13654,N_8229,N_8164);
nor U13655 (N_13655,N_7716,N_7245);
and U13656 (N_13656,N_5304,N_7539);
nand U13657 (N_13657,N_5563,N_8494);
or U13658 (N_13658,N_7767,N_9279);
nand U13659 (N_13659,N_5865,N_6288);
nand U13660 (N_13660,N_8124,N_7721);
or U13661 (N_13661,N_6196,N_7504);
and U13662 (N_13662,N_7796,N_7004);
xor U13663 (N_13663,N_8404,N_8254);
and U13664 (N_13664,N_9709,N_6596);
xor U13665 (N_13665,N_5866,N_8890);
or U13666 (N_13666,N_8778,N_7587);
or U13667 (N_13667,N_5445,N_7438);
nor U13668 (N_13668,N_5531,N_9069);
and U13669 (N_13669,N_9234,N_7506);
nor U13670 (N_13670,N_6467,N_8598);
nand U13671 (N_13671,N_6474,N_5300);
nand U13672 (N_13672,N_9490,N_8609);
or U13673 (N_13673,N_8068,N_9223);
nand U13674 (N_13674,N_7303,N_6825);
nor U13675 (N_13675,N_6413,N_7438);
nand U13676 (N_13676,N_8556,N_7182);
and U13677 (N_13677,N_5081,N_6081);
nor U13678 (N_13678,N_6401,N_6737);
nand U13679 (N_13679,N_6584,N_7963);
or U13680 (N_13680,N_5688,N_6986);
and U13681 (N_13681,N_8880,N_8100);
and U13682 (N_13682,N_6742,N_8495);
nor U13683 (N_13683,N_6551,N_5172);
nand U13684 (N_13684,N_5650,N_8025);
nor U13685 (N_13685,N_5118,N_6485);
nor U13686 (N_13686,N_8841,N_7949);
nand U13687 (N_13687,N_7788,N_7282);
or U13688 (N_13688,N_8830,N_6408);
nand U13689 (N_13689,N_8839,N_8406);
nand U13690 (N_13690,N_9165,N_8110);
nand U13691 (N_13691,N_9491,N_8228);
or U13692 (N_13692,N_5474,N_6603);
and U13693 (N_13693,N_7658,N_8166);
and U13694 (N_13694,N_8880,N_6556);
and U13695 (N_13695,N_6729,N_5449);
and U13696 (N_13696,N_9603,N_5165);
or U13697 (N_13697,N_9593,N_9314);
nor U13698 (N_13698,N_6308,N_7141);
or U13699 (N_13699,N_7579,N_8035);
and U13700 (N_13700,N_9937,N_9086);
or U13701 (N_13701,N_7508,N_7548);
and U13702 (N_13702,N_8662,N_8606);
nand U13703 (N_13703,N_8699,N_8724);
nor U13704 (N_13704,N_6464,N_8636);
nor U13705 (N_13705,N_6815,N_9138);
or U13706 (N_13706,N_6720,N_7476);
xor U13707 (N_13707,N_7503,N_7703);
or U13708 (N_13708,N_7849,N_5042);
and U13709 (N_13709,N_5604,N_5454);
and U13710 (N_13710,N_7976,N_5645);
nor U13711 (N_13711,N_6005,N_5774);
nor U13712 (N_13712,N_8227,N_5049);
and U13713 (N_13713,N_8598,N_6231);
and U13714 (N_13714,N_7265,N_8773);
nand U13715 (N_13715,N_7012,N_9081);
nor U13716 (N_13716,N_5218,N_5578);
nand U13717 (N_13717,N_9565,N_9245);
nand U13718 (N_13718,N_5745,N_8603);
or U13719 (N_13719,N_8739,N_7004);
xnor U13720 (N_13720,N_6640,N_9638);
nand U13721 (N_13721,N_6138,N_9976);
or U13722 (N_13722,N_7452,N_7287);
and U13723 (N_13723,N_9866,N_7820);
or U13724 (N_13724,N_7441,N_8412);
or U13725 (N_13725,N_6357,N_6044);
or U13726 (N_13726,N_6831,N_8029);
nor U13727 (N_13727,N_6046,N_8061);
nor U13728 (N_13728,N_6964,N_6087);
xnor U13729 (N_13729,N_5705,N_5545);
nand U13730 (N_13730,N_9760,N_9202);
and U13731 (N_13731,N_9351,N_5051);
or U13732 (N_13732,N_7214,N_9572);
nand U13733 (N_13733,N_8379,N_7617);
nor U13734 (N_13734,N_8504,N_9724);
nand U13735 (N_13735,N_9904,N_7805);
or U13736 (N_13736,N_6988,N_8739);
nand U13737 (N_13737,N_6574,N_6595);
or U13738 (N_13738,N_9906,N_8354);
nand U13739 (N_13739,N_9262,N_8360);
and U13740 (N_13740,N_8168,N_8103);
and U13741 (N_13741,N_6599,N_9875);
and U13742 (N_13742,N_6960,N_9899);
and U13743 (N_13743,N_6270,N_5399);
nand U13744 (N_13744,N_7106,N_7494);
nand U13745 (N_13745,N_6200,N_5409);
nor U13746 (N_13746,N_8796,N_8963);
and U13747 (N_13747,N_5092,N_8266);
and U13748 (N_13748,N_7523,N_7724);
and U13749 (N_13749,N_7966,N_5455);
nor U13750 (N_13750,N_7012,N_9866);
nand U13751 (N_13751,N_5695,N_6666);
nand U13752 (N_13752,N_5786,N_6617);
nand U13753 (N_13753,N_5216,N_8946);
and U13754 (N_13754,N_7647,N_7294);
and U13755 (N_13755,N_5071,N_8803);
or U13756 (N_13756,N_9300,N_7262);
or U13757 (N_13757,N_9309,N_6559);
or U13758 (N_13758,N_8327,N_7632);
nand U13759 (N_13759,N_6711,N_5372);
or U13760 (N_13760,N_5593,N_8400);
nor U13761 (N_13761,N_9483,N_9428);
and U13762 (N_13762,N_8110,N_5638);
and U13763 (N_13763,N_7275,N_7180);
or U13764 (N_13764,N_5382,N_8604);
and U13765 (N_13765,N_6080,N_5507);
or U13766 (N_13766,N_6550,N_6313);
or U13767 (N_13767,N_9186,N_9155);
nand U13768 (N_13768,N_8258,N_5077);
and U13769 (N_13769,N_9204,N_9482);
and U13770 (N_13770,N_7648,N_6188);
and U13771 (N_13771,N_5606,N_6325);
nand U13772 (N_13772,N_9235,N_8170);
and U13773 (N_13773,N_9215,N_5727);
and U13774 (N_13774,N_7966,N_8569);
nor U13775 (N_13775,N_9391,N_5768);
and U13776 (N_13776,N_7336,N_7078);
nand U13777 (N_13777,N_7850,N_9115);
and U13778 (N_13778,N_7321,N_8741);
nor U13779 (N_13779,N_9794,N_8179);
and U13780 (N_13780,N_5672,N_6958);
or U13781 (N_13781,N_5949,N_8132);
xnor U13782 (N_13782,N_7006,N_7848);
and U13783 (N_13783,N_9969,N_9300);
nand U13784 (N_13784,N_6945,N_6057);
nor U13785 (N_13785,N_6216,N_6681);
nor U13786 (N_13786,N_5908,N_6965);
nand U13787 (N_13787,N_5205,N_7111);
and U13788 (N_13788,N_6302,N_9668);
nand U13789 (N_13789,N_6187,N_8018);
nand U13790 (N_13790,N_8555,N_7249);
and U13791 (N_13791,N_6139,N_8138);
or U13792 (N_13792,N_8710,N_8554);
and U13793 (N_13793,N_9557,N_9739);
nor U13794 (N_13794,N_6982,N_5374);
and U13795 (N_13795,N_8573,N_7809);
or U13796 (N_13796,N_5371,N_7692);
or U13797 (N_13797,N_9132,N_7020);
or U13798 (N_13798,N_9550,N_6210);
and U13799 (N_13799,N_7667,N_6616);
nand U13800 (N_13800,N_5877,N_5207);
or U13801 (N_13801,N_7235,N_9028);
nand U13802 (N_13802,N_5623,N_8622);
and U13803 (N_13803,N_6737,N_6752);
and U13804 (N_13804,N_8673,N_8769);
nor U13805 (N_13805,N_9967,N_6287);
or U13806 (N_13806,N_5929,N_8654);
nand U13807 (N_13807,N_6415,N_9406);
nand U13808 (N_13808,N_9426,N_7776);
or U13809 (N_13809,N_5971,N_5637);
or U13810 (N_13810,N_8774,N_6256);
nand U13811 (N_13811,N_6692,N_7605);
nor U13812 (N_13812,N_8266,N_8148);
nand U13813 (N_13813,N_6264,N_7225);
nand U13814 (N_13814,N_9916,N_6240);
or U13815 (N_13815,N_6357,N_8633);
nor U13816 (N_13816,N_7205,N_9312);
nand U13817 (N_13817,N_8846,N_9517);
nand U13818 (N_13818,N_5772,N_5514);
nand U13819 (N_13819,N_7210,N_9208);
and U13820 (N_13820,N_9298,N_7368);
and U13821 (N_13821,N_7513,N_7541);
or U13822 (N_13822,N_9152,N_7087);
nor U13823 (N_13823,N_7338,N_5941);
or U13824 (N_13824,N_5190,N_9036);
xnor U13825 (N_13825,N_8774,N_6834);
or U13826 (N_13826,N_6593,N_5839);
and U13827 (N_13827,N_9036,N_6263);
nand U13828 (N_13828,N_9097,N_5006);
nor U13829 (N_13829,N_9543,N_7100);
and U13830 (N_13830,N_5335,N_8766);
nand U13831 (N_13831,N_9477,N_8329);
and U13832 (N_13832,N_8698,N_7267);
nand U13833 (N_13833,N_8632,N_6712);
or U13834 (N_13834,N_7706,N_5563);
nor U13835 (N_13835,N_7482,N_9809);
and U13836 (N_13836,N_7368,N_9748);
and U13837 (N_13837,N_9133,N_9613);
and U13838 (N_13838,N_5362,N_8719);
or U13839 (N_13839,N_8731,N_8985);
or U13840 (N_13840,N_5470,N_5650);
and U13841 (N_13841,N_9962,N_5496);
nor U13842 (N_13842,N_7507,N_8556);
nor U13843 (N_13843,N_8025,N_6996);
xnor U13844 (N_13844,N_7586,N_9392);
nand U13845 (N_13845,N_6697,N_9978);
xor U13846 (N_13846,N_8648,N_7730);
and U13847 (N_13847,N_9203,N_5482);
nor U13848 (N_13848,N_6357,N_7719);
and U13849 (N_13849,N_8692,N_8877);
or U13850 (N_13850,N_7486,N_7671);
nand U13851 (N_13851,N_7931,N_5849);
or U13852 (N_13852,N_9199,N_8170);
and U13853 (N_13853,N_7250,N_8947);
nand U13854 (N_13854,N_5721,N_9692);
nor U13855 (N_13855,N_6633,N_7590);
nor U13856 (N_13856,N_5661,N_5431);
or U13857 (N_13857,N_5925,N_5756);
xor U13858 (N_13858,N_8035,N_6887);
or U13859 (N_13859,N_5581,N_7652);
nand U13860 (N_13860,N_5501,N_7787);
and U13861 (N_13861,N_5902,N_6333);
nor U13862 (N_13862,N_7857,N_5672);
and U13863 (N_13863,N_6625,N_5515);
nor U13864 (N_13864,N_7827,N_9605);
nor U13865 (N_13865,N_5739,N_7764);
nor U13866 (N_13866,N_9756,N_8045);
and U13867 (N_13867,N_6821,N_8333);
and U13868 (N_13868,N_5030,N_6462);
nor U13869 (N_13869,N_6328,N_8994);
and U13870 (N_13870,N_8437,N_7611);
or U13871 (N_13871,N_9792,N_5947);
nand U13872 (N_13872,N_6660,N_9286);
xnor U13873 (N_13873,N_7839,N_7108);
or U13874 (N_13874,N_7598,N_8740);
nand U13875 (N_13875,N_6218,N_5714);
xor U13876 (N_13876,N_5885,N_9741);
or U13877 (N_13877,N_5100,N_5856);
nand U13878 (N_13878,N_8996,N_6497);
or U13879 (N_13879,N_6578,N_6478);
nand U13880 (N_13880,N_9019,N_7559);
or U13881 (N_13881,N_6294,N_5818);
nor U13882 (N_13882,N_9884,N_6270);
and U13883 (N_13883,N_6700,N_6013);
or U13884 (N_13884,N_8476,N_6145);
and U13885 (N_13885,N_9530,N_8506);
and U13886 (N_13886,N_5397,N_6672);
nor U13887 (N_13887,N_9115,N_8118);
and U13888 (N_13888,N_9226,N_8296);
nor U13889 (N_13889,N_7037,N_8118);
or U13890 (N_13890,N_8644,N_9309);
nor U13891 (N_13891,N_9172,N_5976);
nand U13892 (N_13892,N_6325,N_8070);
or U13893 (N_13893,N_7081,N_5629);
nor U13894 (N_13894,N_9258,N_6004);
nand U13895 (N_13895,N_7283,N_7589);
nand U13896 (N_13896,N_9646,N_9049);
nor U13897 (N_13897,N_5754,N_9562);
nor U13898 (N_13898,N_6060,N_6705);
or U13899 (N_13899,N_6518,N_6295);
nand U13900 (N_13900,N_8547,N_7322);
nand U13901 (N_13901,N_7913,N_7202);
or U13902 (N_13902,N_6196,N_6640);
or U13903 (N_13903,N_7153,N_5875);
nand U13904 (N_13904,N_6309,N_6367);
or U13905 (N_13905,N_9601,N_8041);
or U13906 (N_13906,N_7723,N_7772);
or U13907 (N_13907,N_5391,N_9952);
and U13908 (N_13908,N_9148,N_5786);
nand U13909 (N_13909,N_6420,N_9178);
and U13910 (N_13910,N_7344,N_6199);
xor U13911 (N_13911,N_9192,N_5797);
or U13912 (N_13912,N_6692,N_8627);
nor U13913 (N_13913,N_7656,N_8115);
and U13914 (N_13914,N_6558,N_6765);
and U13915 (N_13915,N_6987,N_7263);
nor U13916 (N_13916,N_7155,N_9550);
xor U13917 (N_13917,N_9289,N_7684);
nor U13918 (N_13918,N_9577,N_6617);
and U13919 (N_13919,N_5851,N_5299);
nand U13920 (N_13920,N_5215,N_9984);
nand U13921 (N_13921,N_6149,N_9595);
or U13922 (N_13922,N_9492,N_9713);
nand U13923 (N_13923,N_5228,N_5790);
xor U13924 (N_13924,N_6276,N_7085);
nor U13925 (N_13925,N_8669,N_6201);
and U13926 (N_13926,N_5686,N_6478);
and U13927 (N_13927,N_9570,N_7682);
and U13928 (N_13928,N_7208,N_9460);
or U13929 (N_13929,N_8349,N_8478);
nor U13930 (N_13930,N_9107,N_9470);
or U13931 (N_13931,N_7621,N_8613);
and U13932 (N_13932,N_5275,N_9699);
nand U13933 (N_13933,N_8102,N_8904);
and U13934 (N_13934,N_7821,N_9785);
and U13935 (N_13935,N_6801,N_8229);
nand U13936 (N_13936,N_5110,N_8997);
nor U13937 (N_13937,N_6192,N_7162);
nand U13938 (N_13938,N_7652,N_7733);
or U13939 (N_13939,N_7026,N_6026);
nand U13940 (N_13940,N_7795,N_6780);
nand U13941 (N_13941,N_7411,N_6052);
nand U13942 (N_13942,N_5054,N_6416);
or U13943 (N_13943,N_9756,N_8667);
or U13944 (N_13944,N_8834,N_6008);
and U13945 (N_13945,N_7804,N_9989);
nor U13946 (N_13946,N_7235,N_5129);
and U13947 (N_13947,N_8682,N_7251);
and U13948 (N_13948,N_7873,N_6973);
or U13949 (N_13949,N_6172,N_5399);
nor U13950 (N_13950,N_8704,N_8748);
nand U13951 (N_13951,N_8889,N_7811);
or U13952 (N_13952,N_7121,N_9516);
and U13953 (N_13953,N_7075,N_7193);
or U13954 (N_13954,N_9146,N_7375);
nor U13955 (N_13955,N_7082,N_8106);
and U13956 (N_13956,N_8077,N_6856);
or U13957 (N_13957,N_6060,N_5983);
nand U13958 (N_13958,N_8250,N_9183);
nor U13959 (N_13959,N_8146,N_5650);
nand U13960 (N_13960,N_9927,N_8047);
nor U13961 (N_13961,N_6797,N_6083);
nor U13962 (N_13962,N_9486,N_8416);
nor U13963 (N_13963,N_9726,N_9175);
nor U13964 (N_13964,N_8043,N_9675);
nand U13965 (N_13965,N_9836,N_5545);
nor U13966 (N_13966,N_5370,N_9218);
nor U13967 (N_13967,N_8731,N_8631);
or U13968 (N_13968,N_6548,N_9924);
nand U13969 (N_13969,N_8616,N_5511);
nor U13970 (N_13970,N_6036,N_5361);
and U13971 (N_13971,N_9559,N_9172);
nand U13972 (N_13972,N_5492,N_8806);
or U13973 (N_13973,N_9098,N_9560);
xor U13974 (N_13974,N_5129,N_7447);
nand U13975 (N_13975,N_7449,N_6486);
or U13976 (N_13976,N_7587,N_6475);
and U13977 (N_13977,N_8224,N_7563);
nand U13978 (N_13978,N_6987,N_6736);
nand U13979 (N_13979,N_7003,N_6830);
nor U13980 (N_13980,N_9797,N_7198);
and U13981 (N_13981,N_7686,N_7181);
nor U13982 (N_13982,N_5219,N_5022);
and U13983 (N_13983,N_5899,N_9627);
and U13984 (N_13984,N_5639,N_6791);
nand U13985 (N_13985,N_6737,N_6109);
nor U13986 (N_13986,N_8201,N_9629);
and U13987 (N_13987,N_6031,N_5634);
or U13988 (N_13988,N_5369,N_7860);
and U13989 (N_13989,N_6395,N_6578);
nand U13990 (N_13990,N_6827,N_5406);
or U13991 (N_13991,N_6922,N_5862);
and U13992 (N_13992,N_5125,N_9746);
nor U13993 (N_13993,N_6904,N_8837);
nor U13994 (N_13994,N_8145,N_7758);
nor U13995 (N_13995,N_8515,N_7736);
and U13996 (N_13996,N_8570,N_5303);
and U13997 (N_13997,N_6316,N_5887);
and U13998 (N_13998,N_6317,N_7070);
or U13999 (N_13999,N_9203,N_9659);
and U14000 (N_14000,N_6168,N_9292);
nor U14001 (N_14001,N_5077,N_9401);
or U14002 (N_14002,N_7884,N_8958);
nor U14003 (N_14003,N_8949,N_5085);
nand U14004 (N_14004,N_7223,N_5893);
or U14005 (N_14005,N_9025,N_6991);
nand U14006 (N_14006,N_8452,N_7934);
or U14007 (N_14007,N_9017,N_8033);
or U14008 (N_14008,N_6785,N_9551);
or U14009 (N_14009,N_9290,N_7715);
nor U14010 (N_14010,N_5719,N_5731);
or U14011 (N_14011,N_8290,N_6275);
nor U14012 (N_14012,N_5296,N_6830);
nor U14013 (N_14013,N_8799,N_7048);
or U14014 (N_14014,N_5634,N_9648);
and U14015 (N_14015,N_5618,N_8614);
and U14016 (N_14016,N_8414,N_5710);
and U14017 (N_14017,N_5981,N_8169);
and U14018 (N_14018,N_6625,N_7603);
nor U14019 (N_14019,N_9337,N_7930);
or U14020 (N_14020,N_7407,N_5363);
nand U14021 (N_14021,N_6297,N_7485);
nor U14022 (N_14022,N_6776,N_8200);
or U14023 (N_14023,N_6305,N_8732);
and U14024 (N_14024,N_9459,N_8520);
nand U14025 (N_14025,N_5680,N_5655);
and U14026 (N_14026,N_5427,N_8303);
nand U14027 (N_14027,N_8475,N_8198);
nor U14028 (N_14028,N_8028,N_8352);
and U14029 (N_14029,N_8705,N_5605);
nor U14030 (N_14030,N_8532,N_7582);
nor U14031 (N_14031,N_7274,N_7863);
or U14032 (N_14032,N_7477,N_9064);
xor U14033 (N_14033,N_7139,N_9207);
or U14034 (N_14034,N_9278,N_5266);
xnor U14035 (N_14035,N_8817,N_8108);
or U14036 (N_14036,N_9526,N_5627);
nand U14037 (N_14037,N_6659,N_6039);
nor U14038 (N_14038,N_7476,N_8147);
or U14039 (N_14039,N_9286,N_8758);
and U14040 (N_14040,N_7173,N_6859);
or U14041 (N_14041,N_9980,N_8597);
xnor U14042 (N_14042,N_6891,N_6541);
or U14043 (N_14043,N_8623,N_9969);
nor U14044 (N_14044,N_8235,N_9557);
nor U14045 (N_14045,N_7527,N_7273);
nand U14046 (N_14046,N_8710,N_5976);
nor U14047 (N_14047,N_8435,N_8907);
nand U14048 (N_14048,N_8473,N_6446);
nor U14049 (N_14049,N_9551,N_6676);
nor U14050 (N_14050,N_9042,N_9734);
and U14051 (N_14051,N_5094,N_7569);
nand U14052 (N_14052,N_5416,N_8720);
and U14053 (N_14053,N_7837,N_9729);
nor U14054 (N_14054,N_5643,N_7283);
xnor U14055 (N_14055,N_8811,N_7293);
nor U14056 (N_14056,N_8464,N_6143);
and U14057 (N_14057,N_8064,N_9698);
or U14058 (N_14058,N_5307,N_8151);
nand U14059 (N_14059,N_7557,N_6810);
nand U14060 (N_14060,N_6608,N_9296);
or U14061 (N_14061,N_7718,N_6002);
nor U14062 (N_14062,N_8934,N_5330);
nor U14063 (N_14063,N_8696,N_7728);
nor U14064 (N_14064,N_7343,N_7466);
or U14065 (N_14065,N_9039,N_5417);
xor U14066 (N_14066,N_5464,N_7168);
nand U14067 (N_14067,N_7854,N_5932);
or U14068 (N_14068,N_9736,N_9701);
and U14069 (N_14069,N_6024,N_9961);
nand U14070 (N_14070,N_5289,N_6239);
nand U14071 (N_14071,N_7056,N_8359);
or U14072 (N_14072,N_5362,N_5893);
nor U14073 (N_14073,N_6655,N_7533);
nand U14074 (N_14074,N_8322,N_6798);
nor U14075 (N_14075,N_9372,N_5323);
nor U14076 (N_14076,N_5767,N_5380);
and U14077 (N_14077,N_5911,N_7157);
and U14078 (N_14078,N_9149,N_5589);
nand U14079 (N_14079,N_6903,N_5312);
and U14080 (N_14080,N_8214,N_5317);
nand U14081 (N_14081,N_6955,N_8178);
nand U14082 (N_14082,N_9331,N_7235);
and U14083 (N_14083,N_5441,N_7822);
nor U14084 (N_14084,N_7770,N_9356);
and U14085 (N_14085,N_6262,N_7464);
or U14086 (N_14086,N_8810,N_8408);
and U14087 (N_14087,N_5214,N_6771);
and U14088 (N_14088,N_6237,N_5358);
and U14089 (N_14089,N_8039,N_5701);
or U14090 (N_14090,N_6443,N_9067);
or U14091 (N_14091,N_8229,N_5334);
or U14092 (N_14092,N_5558,N_5716);
nand U14093 (N_14093,N_6988,N_9189);
nor U14094 (N_14094,N_6118,N_8110);
nor U14095 (N_14095,N_9675,N_7201);
nor U14096 (N_14096,N_9090,N_8812);
nor U14097 (N_14097,N_8741,N_6743);
and U14098 (N_14098,N_7860,N_9618);
nand U14099 (N_14099,N_9107,N_7423);
nand U14100 (N_14100,N_8240,N_7440);
nor U14101 (N_14101,N_6802,N_7518);
nand U14102 (N_14102,N_7603,N_7700);
nor U14103 (N_14103,N_9730,N_5076);
or U14104 (N_14104,N_7419,N_7282);
or U14105 (N_14105,N_6441,N_8034);
nor U14106 (N_14106,N_5789,N_6073);
or U14107 (N_14107,N_5862,N_6468);
or U14108 (N_14108,N_5100,N_8234);
nand U14109 (N_14109,N_6289,N_6021);
or U14110 (N_14110,N_9896,N_7155);
nand U14111 (N_14111,N_8119,N_8657);
nand U14112 (N_14112,N_7303,N_8393);
nand U14113 (N_14113,N_9818,N_6948);
and U14114 (N_14114,N_8314,N_5266);
nand U14115 (N_14115,N_9720,N_7910);
nand U14116 (N_14116,N_6755,N_8689);
nor U14117 (N_14117,N_7002,N_5571);
nor U14118 (N_14118,N_9108,N_5048);
nor U14119 (N_14119,N_9205,N_5426);
nand U14120 (N_14120,N_9185,N_7231);
and U14121 (N_14121,N_7661,N_6551);
nand U14122 (N_14122,N_8451,N_5494);
nand U14123 (N_14123,N_5629,N_8574);
or U14124 (N_14124,N_8831,N_6527);
or U14125 (N_14125,N_6141,N_5084);
nand U14126 (N_14126,N_8842,N_7585);
nand U14127 (N_14127,N_9488,N_7718);
or U14128 (N_14128,N_5239,N_5900);
and U14129 (N_14129,N_7073,N_9404);
and U14130 (N_14130,N_8156,N_8461);
nor U14131 (N_14131,N_9621,N_6923);
and U14132 (N_14132,N_7321,N_5162);
nand U14133 (N_14133,N_7724,N_9573);
nand U14134 (N_14134,N_7753,N_8087);
nor U14135 (N_14135,N_6480,N_7096);
and U14136 (N_14136,N_8950,N_7025);
nand U14137 (N_14137,N_6459,N_6346);
nor U14138 (N_14138,N_8267,N_5161);
and U14139 (N_14139,N_6175,N_8150);
and U14140 (N_14140,N_6434,N_6229);
or U14141 (N_14141,N_8308,N_7607);
or U14142 (N_14142,N_8475,N_8347);
nor U14143 (N_14143,N_6192,N_6457);
or U14144 (N_14144,N_8215,N_5956);
nor U14145 (N_14145,N_7059,N_7038);
nor U14146 (N_14146,N_7519,N_6306);
or U14147 (N_14147,N_6359,N_8750);
nor U14148 (N_14148,N_9892,N_9223);
and U14149 (N_14149,N_7310,N_6318);
and U14150 (N_14150,N_6329,N_7135);
nor U14151 (N_14151,N_7323,N_6858);
nand U14152 (N_14152,N_9081,N_9794);
nor U14153 (N_14153,N_5789,N_8047);
nor U14154 (N_14154,N_9768,N_7801);
or U14155 (N_14155,N_7747,N_5879);
nor U14156 (N_14156,N_6380,N_5500);
xnor U14157 (N_14157,N_9559,N_6098);
nand U14158 (N_14158,N_5182,N_5383);
nor U14159 (N_14159,N_8678,N_9864);
nand U14160 (N_14160,N_6955,N_5404);
or U14161 (N_14161,N_9480,N_6347);
xnor U14162 (N_14162,N_7579,N_9988);
nor U14163 (N_14163,N_9827,N_7263);
and U14164 (N_14164,N_6506,N_6257);
nor U14165 (N_14165,N_9150,N_7673);
nand U14166 (N_14166,N_5404,N_5998);
or U14167 (N_14167,N_6808,N_8109);
xnor U14168 (N_14168,N_7893,N_5218);
nor U14169 (N_14169,N_8363,N_7844);
nor U14170 (N_14170,N_6018,N_7558);
and U14171 (N_14171,N_5106,N_6162);
nor U14172 (N_14172,N_9148,N_7585);
or U14173 (N_14173,N_9477,N_9123);
nand U14174 (N_14174,N_7654,N_6626);
nor U14175 (N_14175,N_5414,N_9796);
or U14176 (N_14176,N_5263,N_8875);
nand U14177 (N_14177,N_9214,N_6982);
and U14178 (N_14178,N_5414,N_7941);
nor U14179 (N_14179,N_8005,N_5817);
and U14180 (N_14180,N_7262,N_9753);
and U14181 (N_14181,N_5761,N_9244);
nor U14182 (N_14182,N_6563,N_7384);
and U14183 (N_14183,N_6759,N_5341);
and U14184 (N_14184,N_9858,N_7254);
nand U14185 (N_14185,N_5450,N_8772);
nand U14186 (N_14186,N_9238,N_5930);
nor U14187 (N_14187,N_9608,N_7452);
or U14188 (N_14188,N_7487,N_7131);
nor U14189 (N_14189,N_8393,N_9524);
nand U14190 (N_14190,N_8898,N_9853);
or U14191 (N_14191,N_7525,N_6545);
and U14192 (N_14192,N_9778,N_7210);
nand U14193 (N_14193,N_6566,N_6517);
nor U14194 (N_14194,N_8148,N_9348);
nor U14195 (N_14195,N_5900,N_9562);
or U14196 (N_14196,N_6818,N_8674);
or U14197 (N_14197,N_9131,N_7977);
nor U14198 (N_14198,N_9711,N_6572);
or U14199 (N_14199,N_5355,N_8966);
or U14200 (N_14200,N_7385,N_5433);
nand U14201 (N_14201,N_5531,N_5951);
and U14202 (N_14202,N_9890,N_8934);
or U14203 (N_14203,N_8844,N_6581);
nor U14204 (N_14204,N_6629,N_5029);
nor U14205 (N_14205,N_9391,N_9252);
and U14206 (N_14206,N_6220,N_6026);
nand U14207 (N_14207,N_7661,N_9158);
nor U14208 (N_14208,N_7123,N_5410);
or U14209 (N_14209,N_8649,N_5472);
and U14210 (N_14210,N_5504,N_6245);
and U14211 (N_14211,N_6103,N_8016);
or U14212 (N_14212,N_8951,N_7097);
nor U14213 (N_14213,N_8120,N_7331);
nor U14214 (N_14214,N_9202,N_8502);
nand U14215 (N_14215,N_8061,N_7202);
nand U14216 (N_14216,N_9532,N_6114);
nor U14217 (N_14217,N_7409,N_8125);
and U14218 (N_14218,N_6514,N_9822);
nand U14219 (N_14219,N_7361,N_6862);
nor U14220 (N_14220,N_5631,N_5433);
nand U14221 (N_14221,N_9282,N_6385);
nor U14222 (N_14222,N_9357,N_5878);
nor U14223 (N_14223,N_8206,N_6502);
nor U14224 (N_14224,N_5569,N_9046);
or U14225 (N_14225,N_6714,N_6197);
or U14226 (N_14226,N_7736,N_9561);
or U14227 (N_14227,N_5660,N_5816);
nand U14228 (N_14228,N_7249,N_9602);
or U14229 (N_14229,N_8799,N_5046);
nor U14230 (N_14230,N_9321,N_8943);
and U14231 (N_14231,N_8717,N_6893);
and U14232 (N_14232,N_7554,N_5089);
and U14233 (N_14233,N_8274,N_5242);
or U14234 (N_14234,N_6288,N_5973);
nor U14235 (N_14235,N_9608,N_6792);
or U14236 (N_14236,N_8130,N_9569);
nand U14237 (N_14237,N_5198,N_7826);
or U14238 (N_14238,N_6844,N_9103);
or U14239 (N_14239,N_6417,N_6655);
nand U14240 (N_14240,N_7656,N_9469);
or U14241 (N_14241,N_9169,N_6812);
nor U14242 (N_14242,N_7841,N_5574);
nand U14243 (N_14243,N_7198,N_8716);
or U14244 (N_14244,N_7237,N_8445);
and U14245 (N_14245,N_6290,N_8832);
and U14246 (N_14246,N_8352,N_6394);
and U14247 (N_14247,N_5022,N_8874);
or U14248 (N_14248,N_5443,N_6514);
and U14249 (N_14249,N_6819,N_5145);
or U14250 (N_14250,N_7347,N_8611);
or U14251 (N_14251,N_7674,N_9207);
or U14252 (N_14252,N_9199,N_6568);
and U14253 (N_14253,N_6855,N_9545);
nor U14254 (N_14254,N_8056,N_5210);
xor U14255 (N_14255,N_6126,N_8832);
nor U14256 (N_14256,N_7084,N_7984);
nand U14257 (N_14257,N_5952,N_8178);
or U14258 (N_14258,N_7769,N_7069);
or U14259 (N_14259,N_7645,N_6182);
or U14260 (N_14260,N_5768,N_5187);
and U14261 (N_14261,N_9561,N_8043);
nor U14262 (N_14262,N_7433,N_9707);
and U14263 (N_14263,N_7207,N_5910);
nor U14264 (N_14264,N_9849,N_6439);
and U14265 (N_14265,N_6557,N_7962);
nand U14266 (N_14266,N_7389,N_8479);
or U14267 (N_14267,N_8001,N_6401);
nand U14268 (N_14268,N_8538,N_8882);
or U14269 (N_14269,N_8290,N_7104);
or U14270 (N_14270,N_6893,N_7126);
xnor U14271 (N_14271,N_6136,N_7580);
and U14272 (N_14272,N_8632,N_9736);
and U14273 (N_14273,N_9162,N_6035);
and U14274 (N_14274,N_5558,N_6534);
nor U14275 (N_14275,N_6236,N_7378);
and U14276 (N_14276,N_6840,N_9745);
nor U14277 (N_14277,N_6079,N_7868);
xnor U14278 (N_14278,N_6343,N_6122);
and U14279 (N_14279,N_6247,N_7991);
and U14280 (N_14280,N_6071,N_7189);
nand U14281 (N_14281,N_6809,N_6143);
nand U14282 (N_14282,N_9335,N_5118);
and U14283 (N_14283,N_7440,N_6590);
or U14284 (N_14284,N_8625,N_5721);
nand U14285 (N_14285,N_9962,N_6343);
nand U14286 (N_14286,N_9637,N_6934);
nand U14287 (N_14287,N_5949,N_9839);
nor U14288 (N_14288,N_7939,N_5689);
nor U14289 (N_14289,N_6513,N_9505);
xnor U14290 (N_14290,N_7809,N_6763);
and U14291 (N_14291,N_9153,N_7096);
nand U14292 (N_14292,N_8082,N_5677);
and U14293 (N_14293,N_6879,N_5314);
nand U14294 (N_14294,N_5568,N_5079);
or U14295 (N_14295,N_9542,N_5335);
and U14296 (N_14296,N_6823,N_6722);
or U14297 (N_14297,N_6594,N_6957);
or U14298 (N_14298,N_7026,N_5660);
or U14299 (N_14299,N_5334,N_6843);
xnor U14300 (N_14300,N_9034,N_6469);
nand U14301 (N_14301,N_7139,N_7776);
or U14302 (N_14302,N_6491,N_7243);
xnor U14303 (N_14303,N_6022,N_7794);
and U14304 (N_14304,N_6578,N_5421);
or U14305 (N_14305,N_8313,N_5152);
and U14306 (N_14306,N_5719,N_5263);
nor U14307 (N_14307,N_7072,N_7603);
and U14308 (N_14308,N_7860,N_5728);
nand U14309 (N_14309,N_7736,N_9815);
or U14310 (N_14310,N_7192,N_8855);
and U14311 (N_14311,N_7750,N_7717);
or U14312 (N_14312,N_6670,N_5945);
or U14313 (N_14313,N_9950,N_5959);
or U14314 (N_14314,N_8313,N_8607);
nand U14315 (N_14315,N_7156,N_8518);
nor U14316 (N_14316,N_6022,N_8582);
and U14317 (N_14317,N_8464,N_9675);
nand U14318 (N_14318,N_5776,N_8788);
nand U14319 (N_14319,N_6866,N_7552);
nand U14320 (N_14320,N_5653,N_6585);
nor U14321 (N_14321,N_7258,N_5356);
or U14322 (N_14322,N_6233,N_5998);
and U14323 (N_14323,N_9601,N_9667);
and U14324 (N_14324,N_9121,N_8878);
nor U14325 (N_14325,N_9297,N_7165);
nand U14326 (N_14326,N_9309,N_6196);
nor U14327 (N_14327,N_6038,N_5550);
nand U14328 (N_14328,N_9076,N_8165);
and U14329 (N_14329,N_8807,N_9363);
and U14330 (N_14330,N_6279,N_6123);
nand U14331 (N_14331,N_8841,N_7824);
and U14332 (N_14332,N_9412,N_5301);
or U14333 (N_14333,N_7621,N_6869);
or U14334 (N_14334,N_7682,N_8131);
and U14335 (N_14335,N_5118,N_6824);
and U14336 (N_14336,N_6596,N_5208);
or U14337 (N_14337,N_6521,N_5600);
and U14338 (N_14338,N_9985,N_8674);
and U14339 (N_14339,N_7397,N_6207);
and U14340 (N_14340,N_5087,N_6547);
and U14341 (N_14341,N_6414,N_6637);
nand U14342 (N_14342,N_7589,N_5314);
or U14343 (N_14343,N_7268,N_8767);
nand U14344 (N_14344,N_5815,N_5329);
or U14345 (N_14345,N_6438,N_5984);
nor U14346 (N_14346,N_7655,N_9340);
or U14347 (N_14347,N_8396,N_9569);
or U14348 (N_14348,N_5015,N_8615);
or U14349 (N_14349,N_9033,N_9190);
or U14350 (N_14350,N_8403,N_5273);
nor U14351 (N_14351,N_5825,N_5571);
and U14352 (N_14352,N_7386,N_8389);
or U14353 (N_14353,N_9796,N_5216);
and U14354 (N_14354,N_6681,N_5209);
and U14355 (N_14355,N_7067,N_6886);
and U14356 (N_14356,N_6563,N_8710);
nor U14357 (N_14357,N_5459,N_8133);
nor U14358 (N_14358,N_9661,N_5723);
and U14359 (N_14359,N_8643,N_8070);
or U14360 (N_14360,N_9619,N_6397);
nor U14361 (N_14361,N_7431,N_5954);
and U14362 (N_14362,N_6485,N_7360);
nand U14363 (N_14363,N_9895,N_8005);
and U14364 (N_14364,N_5085,N_5019);
and U14365 (N_14365,N_6816,N_7337);
or U14366 (N_14366,N_9963,N_8716);
or U14367 (N_14367,N_5372,N_9222);
nor U14368 (N_14368,N_7692,N_5772);
nor U14369 (N_14369,N_5482,N_9520);
or U14370 (N_14370,N_7771,N_9516);
nor U14371 (N_14371,N_6871,N_6699);
or U14372 (N_14372,N_9247,N_6000);
nor U14373 (N_14373,N_9411,N_5009);
nand U14374 (N_14374,N_6980,N_6615);
and U14375 (N_14375,N_5075,N_9176);
and U14376 (N_14376,N_5148,N_5502);
or U14377 (N_14377,N_6687,N_8551);
nor U14378 (N_14378,N_8810,N_7487);
nand U14379 (N_14379,N_8784,N_9178);
nand U14380 (N_14380,N_6293,N_9853);
and U14381 (N_14381,N_9246,N_8863);
nor U14382 (N_14382,N_9639,N_5111);
nand U14383 (N_14383,N_9301,N_9794);
nand U14384 (N_14384,N_9063,N_6215);
and U14385 (N_14385,N_6215,N_5778);
nor U14386 (N_14386,N_7290,N_7269);
and U14387 (N_14387,N_8117,N_9508);
nor U14388 (N_14388,N_9245,N_7321);
or U14389 (N_14389,N_7415,N_6292);
or U14390 (N_14390,N_6870,N_5352);
and U14391 (N_14391,N_9228,N_9856);
or U14392 (N_14392,N_9451,N_6545);
xor U14393 (N_14393,N_6844,N_9668);
or U14394 (N_14394,N_7412,N_5820);
and U14395 (N_14395,N_8761,N_7141);
and U14396 (N_14396,N_8568,N_5196);
and U14397 (N_14397,N_6080,N_5023);
nand U14398 (N_14398,N_7888,N_7874);
or U14399 (N_14399,N_8780,N_5035);
nor U14400 (N_14400,N_7404,N_8463);
nor U14401 (N_14401,N_9024,N_5311);
or U14402 (N_14402,N_8480,N_5460);
nor U14403 (N_14403,N_8139,N_5325);
nor U14404 (N_14404,N_5962,N_9627);
or U14405 (N_14405,N_9885,N_5431);
nand U14406 (N_14406,N_7198,N_5031);
nand U14407 (N_14407,N_5994,N_6685);
nor U14408 (N_14408,N_8129,N_7097);
or U14409 (N_14409,N_6786,N_8226);
or U14410 (N_14410,N_8176,N_8475);
and U14411 (N_14411,N_8912,N_5150);
nand U14412 (N_14412,N_8351,N_6861);
or U14413 (N_14413,N_7139,N_8433);
nor U14414 (N_14414,N_6740,N_9913);
or U14415 (N_14415,N_9405,N_5871);
nand U14416 (N_14416,N_5168,N_7371);
nand U14417 (N_14417,N_6548,N_9047);
and U14418 (N_14418,N_8700,N_8807);
or U14419 (N_14419,N_9009,N_7400);
nor U14420 (N_14420,N_9607,N_8625);
or U14421 (N_14421,N_5579,N_6612);
xnor U14422 (N_14422,N_9530,N_8701);
and U14423 (N_14423,N_9048,N_6670);
nor U14424 (N_14424,N_8773,N_5257);
and U14425 (N_14425,N_8471,N_6098);
nand U14426 (N_14426,N_9436,N_7279);
and U14427 (N_14427,N_5213,N_6523);
nor U14428 (N_14428,N_8961,N_6141);
and U14429 (N_14429,N_6410,N_9905);
nor U14430 (N_14430,N_9833,N_5512);
nand U14431 (N_14431,N_5731,N_9480);
nor U14432 (N_14432,N_8533,N_8671);
nor U14433 (N_14433,N_9039,N_7927);
and U14434 (N_14434,N_5567,N_8110);
or U14435 (N_14435,N_8868,N_6155);
nor U14436 (N_14436,N_6546,N_6746);
and U14437 (N_14437,N_6386,N_6080);
or U14438 (N_14438,N_8556,N_5824);
and U14439 (N_14439,N_6756,N_8710);
or U14440 (N_14440,N_5389,N_5084);
or U14441 (N_14441,N_9015,N_5904);
nor U14442 (N_14442,N_6939,N_5787);
nand U14443 (N_14443,N_8264,N_8030);
or U14444 (N_14444,N_7590,N_6037);
nor U14445 (N_14445,N_7941,N_6259);
or U14446 (N_14446,N_5046,N_5850);
nor U14447 (N_14447,N_9273,N_5173);
or U14448 (N_14448,N_5136,N_8254);
nand U14449 (N_14449,N_8751,N_9202);
nand U14450 (N_14450,N_9262,N_9177);
nand U14451 (N_14451,N_9584,N_5631);
nor U14452 (N_14452,N_8388,N_9656);
nand U14453 (N_14453,N_8993,N_7472);
or U14454 (N_14454,N_8718,N_9214);
nand U14455 (N_14455,N_9447,N_6867);
nor U14456 (N_14456,N_5952,N_9898);
and U14457 (N_14457,N_7666,N_5913);
nand U14458 (N_14458,N_9113,N_5198);
or U14459 (N_14459,N_6439,N_7477);
nor U14460 (N_14460,N_9510,N_7530);
and U14461 (N_14461,N_7507,N_8775);
nand U14462 (N_14462,N_6298,N_7270);
nor U14463 (N_14463,N_5603,N_6461);
or U14464 (N_14464,N_7188,N_7071);
or U14465 (N_14465,N_9023,N_6255);
or U14466 (N_14466,N_5053,N_8520);
or U14467 (N_14467,N_7185,N_7742);
nor U14468 (N_14468,N_6063,N_9641);
nor U14469 (N_14469,N_6835,N_7642);
nor U14470 (N_14470,N_6803,N_5891);
or U14471 (N_14471,N_6549,N_7546);
or U14472 (N_14472,N_8011,N_9192);
nor U14473 (N_14473,N_8460,N_5273);
or U14474 (N_14474,N_8274,N_9752);
nor U14475 (N_14475,N_8366,N_7304);
and U14476 (N_14476,N_7831,N_7022);
xnor U14477 (N_14477,N_8265,N_9230);
nor U14478 (N_14478,N_5911,N_8433);
or U14479 (N_14479,N_6847,N_9779);
and U14480 (N_14480,N_5348,N_5066);
nor U14481 (N_14481,N_5685,N_6254);
nand U14482 (N_14482,N_7999,N_8162);
nand U14483 (N_14483,N_5547,N_8246);
or U14484 (N_14484,N_6461,N_9700);
nor U14485 (N_14485,N_8738,N_5968);
and U14486 (N_14486,N_9398,N_8019);
and U14487 (N_14487,N_9999,N_7049);
or U14488 (N_14488,N_8945,N_7417);
or U14489 (N_14489,N_6159,N_6768);
nand U14490 (N_14490,N_5020,N_5421);
nor U14491 (N_14491,N_6052,N_8721);
and U14492 (N_14492,N_8834,N_5714);
and U14493 (N_14493,N_7025,N_7051);
nand U14494 (N_14494,N_5153,N_6888);
nand U14495 (N_14495,N_9842,N_8417);
nor U14496 (N_14496,N_9855,N_7231);
nor U14497 (N_14497,N_8640,N_7770);
nand U14498 (N_14498,N_8488,N_8924);
nor U14499 (N_14499,N_9943,N_5966);
and U14500 (N_14500,N_9151,N_7335);
nand U14501 (N_14501,N_7608,N_5547);
and U14502 (N_14502,N_7578,N_5415);
nand U14503 (N_14503,N_9746,N_6570);
or U14504 (N_14504,N_6139,N_9782);
nor U14505 (N_14505,N_6352,N_9435);
and U14506 (N_14506,N_8233,N_9089);
and U14507 (N_14507,N_8683,N_9827);
nor U14508 (N_14508,N_9357,N_9725);
nand U14509 (N_14509,N_6288,N_7699);
nand U14510 (N_14510,N_6495,N_8241);
or U14511 (N_14511,N_7284,N_7742);
and U14512 (N_14512,N_5553,N_9970);
nand U14513 (N_14513,N_5800,N_8350);
nand U14514 (N_14514,N_5844,N_7280);
nand U14515 (N_14515,N_6559,N_9099);
nor U14516 (N_14516,N_8052,N_6712);
nand U14517 (N_14517,N_7901,N_8970);
nand U14518 (N_14518,N_9831,N_7177);
or U14519 (N_14519,N_5576,N_8976);
xor U14520 (N_14520,N_7797,N_8311);
nand U14521 (N_14521,N_7883,N_7111);
nor U14522 (N_14522,N_8804,N_6991);
and U14523 (N_14523,N_8855,N_9205);
nand U14524 (N_14524,N_9291,N_5307);
nor U14525 (N_14525,N_5609,N_5058);
nor U14526 (N_14526,N_6210,N_9816);
nor U14527 (N_14527,N_8529,N_7512);
or U14528 (N_14528,N_8550,N_7089);
or U14529 (N_14529,N_9674,N_8491);
nor U14530 (N_14530,N_7787,N_8881);
or U14531 (N_14531,N_7409,N_7603);
nor U14532 (N_14532,N_8389,N_8721);
xnor U14533 (N_14533,N_6361,N_9325);
xnor U14534 (N_14534,N_7181,N_9764);
nor U14535 (N_14535,N_6010,N_9891);
and U14536 (N_14536,N_5510,N_6421);
or U14537 (N_14537,N_5758,N_5960);
nand U14538 (N_14538,N_7605,N_5993);
or U14539 (N_14539,N_7054,N_7199);
nand U14540 (N_14540,N_6506,N_6836);
nand U14541 (N_14541,N_5435,N_8985);
nand U14542 (N_14542,N_9529,N_7316);
and U14543 (N_14543,N_6702,N_9502);
and U14544 (N_14544,N_9165,N_8946);
nand U14545 (N_14545,N_7095,N_9638);
or U14546 (N_14546,N_9220,N_7213);
nand U14547 (N_14547,N_9254,N_8036);
nand U14548 (N_14548,N_8165,N_9138);
or U14549 (N_14549,N_5237,N_9972);
xor U14550 (N_14550,N_8399,N_5188);
nand U14551 (N_14551,N_7193,N_5391);
and U14552 (N_14552,N_6914,N_7208);
nor U14553 (N_14553,N_6436,N_8441);
nor U14554 (N_14554,N_8362,N_5702);
or U14555 (N_14555,N_9381,N_6839);
or U14556 (N_14556,N_6150,N_9991);
or U14557 (N_14557,N_7355,N_8256);
or U14558 (N_14558,N_6633,N_8473);
and U14559 (N_14559,N_7459,N_8027);
nor U14560 (N_14560,N_9719,N_7572);
nand U14561 (N_14561,N_8902,N_6494);
nand U14562 (N_14562,N_6311,N_5886);
nand U14563 (N_14563,N_6077,N_5250);
and U14564 (N_14564,N_6208,N_6561);
xnor U14565 (N_14565,N_7134,N_5092);
or U14566 (N_14566,N_9906,N_5742);
nand U14567 (N_14567,N_6757,N_6437);
nor U14568 (N_14568,N_9772,N_6867);
and U14569 (N_14569,N_9921,N_7351);
nor U14570 (N_14570,N_7143,N_8663);
and U14571 (N_14571,N_8614,N_6770);
or U14572 (N_14572,N_5943,N_6295);
nor U14573 (N_14573,N_9344,N_7589);
nor U14574 (N_14574,N_5116,N_9506);
nor U14575 (N_14575,N_9499,N_5927);
nor U14576 (N_14576,N_6536,N_6000);
nor U14577 (N_14577,N_5594,N_9893);
nor U14578 (N_14578,N_7494,N_6799);
or U14579 (N_14579,N_5235,N_8269);
or U14580 (N_14580,N_8792,N_9959);
or U14581 (N_14581,N_6890,N_9580);
and U14582 (N_14582,N_9601,N_8192);
or U14583 (N_14583,N_7670,N_7302);
nand U14584 (N_14584,N_5567,N_5589);
nand U14585 (N_14585,N_5470,N_9818);
and U14586 (N_14586,N_6649,N_6709);
nand U14587 (N_14587,N_7600,N_8704);
and U14588 (N_14588,N_9986,N_6566);
nor U14589 (N_14589,N_6633,N_6050);
nand U14590 (N_14590,N_5420,N_6092);
nand U14591 (N_14591,N_5541,N_7517);
nand U14592 (N_14592,N_5684,N_9444);
or U14593 (N_14593,N_5058,N_6927);
and U14594 (N_14594,N_9159,N_6243);
nor U14595 (N_14595,N_5998,N_9223);
xor U14596 (N_14596,N_5293,N_6272);
nand U14597 (N_14597,N_8522,N_8707);
or U14598 (N_14598,N_5001,N_5746);
or U14599 (N_14599,N_7907,N_7145);
nand U14600 (N_14600,N_9196,N_6496);
and U14601 (N_14601,N_5879,N_8577);
and U14602 (N_14602,N_7224,N_7738);
nor U14603 (N_14603,N_6575,N_7491);
xnor U14604 (N_14604,N_9141,N_9964);
or U14605 (N_14605,N_6238,N_5684);
nor U14606 (N_14606,N_7507,N_7483);
and U14607 (N_14607,N_7438,N_7111);
nand U14608 (N_14608,N_9604,N_8163);
or U14609 (N_14609,N_6435,N_7018);
nor U14610 (N_14610,N_8949,N_8984);
or U14611 (N_14611,N_7876,N_8563);
nand U14612 (N_14612,N_7073,N_8670);
or U14613 (N_14613,N_5945,N_8621);
xor U14614 (N_14614,N_9309,N_9381);
nand U14615 (N_14615,N_9674,N_6741);
or U14616 (N_14616,N_9303,N_5749);
nand U14617 (N_14617,N_6053,N_7600);
or U14618 (N_14618,N_9482,N_9893);
nand U14619 (N_14619,N_7697,N_5009);
nand U14620 (N_14620,N_8234,N_6506);
nand U14621 (N_14621,N_5383,N_8294);
and U14622 (N_14622,N_9887,N_8715);
nor U14623 (N_14623,N_9024,N_7447);
nand U14624 (N_14624,N_5797,N_8630);
nor U14625 (N_14625,N_5959,N_9802);
or U14626 (N_14626,N_7992,N_6871);
or U14627 (N_14627,N_8636,N_8957);
or U14628 (N_14628,N_6208,N_5972);
and U14629 (N_14629,N_8732,N_5301);
nand U14630 (N_14630,N_7803,N_6814);
nand U14631 (N_14631,N_5130,N_7339);
or U14632 (N_14632,N_6225,N_9450);
and U14633 (N_14633,N_8737,N_8204);
and U14634 (N_14634,N_6978,N_6829);
nand U14635 (N_14635,N_9285,N_7163);
or U14636 (N_14636,N_5582,N_8877);
nand U14637 (N_14637,N_5414,N_6782);
or U14638 (N_14638,N_8612,N_9635);
and U14639 (N_14639,N_7251,N_6818);
nand U14640 (N_14640,N_7490,N_9033);
or U14641 (N_14641,N_9457,N_6837);
or U14642 (N_14642,N_8895,N_8384);
and U14643 (N_14643,N_8302,N_5794);
xnor U14644 (N_14644,N_6617,N_5459);
nand U14645 (N_14645,N_6818,N_6996);
nand U14646 (N_14646,N_6608,N_9828);
and U14647 (N_14647,N_7412,N_7564);
and U14648 (N_14648,N_5935,N_5570);
xor U14649 (N_14649,N_9063,N_5999);
and U14650 (N_14650,N_8132,N_8699);
nor U14651 (N_14651,N_7418,N_5110);
or U14652 (N_14652,N_8548,N_5069);
nand U14653 (N_14653,N_6729,N_6973);
nor U14654 (N_14654,N_9607,N_9663);
nor U14655 (N_14655,N_6423,N_9287);
and U14656 (N_14656,N_9200,N_5757);
nand U14657 (N_14657,N_6807,N_7296);
and U14658 (N_14658,N_9327,N_8726);
nor U14659 (N_14659,N_5614,N_8719);
nand U14660 (N_14660,N_7892,N_8456);
nor U14661 (N_14661,N_5241,N_7503);
or U14662 (N_14662,N_9568,N_7714);
nor U14663 (N_14663,N_5532,N_5017);
nand U14664 (N_14664,N_6583,N_9723);
xnor U14665 (N_14665,N_9530,N_5374);
nor U14666 (N_14666,N_7841,N_9528);
nor U14667 (N_14667,N_9712,N_9515);
nand U14668 (N_14668,N_9133,N_9019);
and U14669 (N_14669,N_8190,N_5555);
nand U14670 (N_14670,N_6371,N_8776);
nand U14671 (N_14671,N_5446,N_7960);
or U14672 (N_14672,N_7827,N_8733);
and U14673 (N_14673,N_7440,N_7899);
or U14674 (N_14674,N_9771,N_8655);
or U14675 (N_14675,N_8924,N_8191);
nor U14676 (N_14676,N_7635,N_7509);
nor U14677 (N_14677,N_7107,N_6872);
and U14678 (N_14678,N_8615,N_7139);
nand U14679 (N_14679,N_6903,N_8801);
or U14680 (N_14680,N_7680,N_7367);
or U14681 (N_14681,N_6307,N_6792);
and U14682 (N_14682,N_9131,N_9054);
or U14683 (N_14683,N_6968,N_8596);
nand U14684 (N_14684,N_8429,N_8009);
nor U14685 (N_14685,N_5085,N_8348);
nand U14686 (N_14686,N_9292,N_9854);
nand U14687 (N_14687,N_8091,N_7112);
nand U14688 (N_14688,N_7437,N_8665);
nand U14689 (N_14689,N_6294,N_8933);
or U14690 (N_14690,N_5849,N_6555);
nor U14691 (N_14691,N_5731,N_8264);
and U14692 (N_14692,N_5492,N_9106);
or U14693 (N_14693,N_7266,N_6776);
nand U14694 (N_14694,N_9583,N_8496);
nand U14695 (N_14695,N_9724,N_9185);
nand U14696 (N_14696,N_8612,N_5448);
nor U14697 (N_14697,N_8758,N_6090);
and U14698 (N_14698,N_7750,N_8930);
and U14699 (N_14699,N_9135,N_8434);
and U14700 (N_14700,N_7261,N_7684);
and U14701 (N_14701,N_9317,N_9012);
nand U14702 (N_14702,N_9427,N_6890);
nand U14703 (N_14703,N_7758,N_5442);
or U14704 (N_14704,N_6595,N_8783);
nand U14705 (N_14705,N_6701,N_7500);
nor U14706 (N_14706,N_7760,N_7484);
and U14707 (N_14707,N_5887,N_6067);
or U14708 (N_14708,N_7348,N_9391);
and U14709 (N_14709,N_9268,N_7409);
nand U14710 (N_14710,N_6284,N_6616);
and U14711 (N_14711,N_5254,N_9028);
nand U14712 (N_14712,N_7730,N_7182);
nor U14713 (N_14713,N_6422,N_8768);
or U14714 (N_14714,N_5053,N_5117);
nand U14715 (N_14715,N_5081,N_6873);
nor U14716 (N_14716,N_5595,N_9977);
nor U14717 (N_14717,N_7988,N_5328);
nand U14718 (N_14718,N_8384,N_5391);
or U14719 (N_14719,N_6313,N_6745);
nor U14720 (N_14720,N_8245,N_8768);
and U14721 (N_14721,N_8773,N_8873);
or U14722 (N_14722,N_9573,N_7804);
or U14723 (N_14723,N_8428,N_9585);
and U14724 (N_14724,N_5982,N_9588);
and U14725 (N_14725,N_9214,N_8872);
nand U14726 (N_14726,N_5202,N_6832);
and U14727 (N_14727,N_6205,N_6362);
nand U14728 (N_14728,N_7977,N_6939);
or U14729 (N_14729,N_9100,N_6220);
nor U14730 (N_14730,N_9854,N_8249);
or U14731 (N_14731,N_9454,N_8613);
nor U14732 (N_14732,N_9260,N_8374);
or U14733 (N_14733,N_7587,N_7850);
nand U14734 (N_14734,N_6125,N_7865);
nor U14735 (N_14735,N_6098,N_6290);
nor U14736 (N_14736,N_5249,N_7299);
or U14737 (N_14737,N_5171,N_5309);
or U14738 (N_14738,N_7405,N_8195);
and U14739 (N_14739,N_6500,N_9936);
and U14740 (N_14740,N_6917,N_7061);
nand U14741 (N_14741,N_9863,N_6746);
nand U14742 (N_14742,N_8711,N_6687);
nor U14743 (N_14743,N_9966,N_5833);
nor U14744 (N_14744,N_9267,N_5044);
nor U14745 (N_14745,N_6671,N_7837);
xor U14746 (N_14746,N_6636,N_9584);
and U14747 (N_14747,N_9395,N_8834);
or U14748 (N_14748,N_7988,N_6949);
or U14749 (N_14749,N_6915,N_7429);
nand U14750 (N_14750,N_7948,N_9692);
nand U14751 (N_14751,N_7492,N_5403);
nand U14752 (N_14752,N_8452,N_8597);
nor U14753 (N_14753,N_7281,N_6898);
nand U14754 (N_14754,N_6322,N_8379);
and U14755 (N_14755,N_8565,N_5160);
nand U14756 (N_14756,N_5954,N_7918);
nor U14757 (N_14757,N_5493,N_5029);
nor U14758 (N_14758,N_5642,N_9596);
xor U14759 (N_14759,N_9405,N_7892);
or U14760 (N_14760,N_6494,N_8834);
nor U14761 (N_14761,N_6892,N_7861);
or U14762 (N_14762,N_9305,N_6777);
or U14763 (N_14763,N_9651,N_6592);
nor U14764 (N_14764,N_5786,N_9871);
nand U14765 (N_14765,N_8932,N_7227);
xor U14766 (N_14766,N_5360,N_7911);
nand U14767 (N_14767,N_9833,N_5786);
nand U14768 (N_14768,N_8562,N_9780);
nand U14769 (N_14769,N_9902,N_8642);
nand U14770 (N_14770,N_5888,N_5370);
and U14771 (N_14771,N_6797,N_6443);
nor U14772 (N_14772,N_5162,N_7437);
and U14773 (N_14773,N_6129,N_9941);
or U14774 (N_14774,N_7762,N_8701);
or U14775 (N_14775,N_9351,N_6041);
nand U14776 (N_14776,N_5037,N_6397);
and U14777 (N_14777,N_5057,N_5922);
nor U14778 (N_14778,N_9195,N_5112);
or U14779 (N_14779,N_8445,N_8861);
nand U14780 (N_14780,N_8355,N_5844);
and U14781 (N_14781,N_7406,N_7765);
nor U14782 (N_14782,N_6528,N_9393);
or U14783 (N_14783,N_8668,N_5549);
and U14784 (N_14784,N_6331,N_7020);
and U14785 (N_14785,N_7660,N_9591);
and U14786 (N_14786,N_8519,N_5937);
nand U14787 (N_14787,N_7983,N_5877);
or U14788 (N_14788,N_8546,N_9908);
and U14789 (N_14789,N_7359,N_6030);
and U14790 (N_14790,N_9707,N_9548);
nand U14791 (N_14791,N_7437,N_7814);
and U14792 (N_14792,N_6489,N_5588);
and U14793 (N_14793,N_8138,N_8890);
and U14794 (N_14794,N_7240,N_5610);
or U14795 (N_14795,N_9662,N_5077);
nand U14796 (N_14796,N_8524,N_7264);
and U14797 (N_14797,N_9019,N_5365);
nor U14798 (N_14798,N_6070,N_6307);
nor U14799 (N_14799,N_5278,N_5607);
nor U14800 (N_14800,N_8968,N_5794);
nand U14801 (N_14801,N_6928,N_9431);
nor U14802 (N_14802,N_8070,N_8724);
and U14803 (N_14803,N_8142,N_9468);
nand U14804 (N_14804,N_9809,N_9065);
and U14805 (N_14805,N_7262,N_8505);
nand U14806 (N_14806,N_6019,N_6270);
and U14807 (N_14807,N_7060,N_6384);
xor U14808 (N_14808,N_5633,N_7011);
or U14809 (N_14809,N_7565,N_9675);
or U14810 (N_14810,N_9269,N_5835);
and U14811 (N_14811,N_9385,N_5481);
nand U14812 (N_14812,N_7672,N_7070);
nand U14813 (N_14813,N_6816,N_6903);
nand U14814 (N_14814,N_6107,N_7115);
nor U14815 (N_14815,N_8290,N_5904);
or U14816 (N_14816,N_5211,N_5581);
and U14817 (N_14817,N_7337,N_6102);
nor U14818 (N_14818,N_9574,N_7702);
nand U14819 (N_14819,N_6785,N_8801);
nand U14820 (N_14820,N_6594,N_8043);
or U14821 (N_14821,N_5029,N_9913);
nor U14822 (N_14822,N_7609,N_7162);
nor U14823 (N_14823,N_8705,N_7821);
nand U14824 (N_14824,N_9262,N_9923);
or U14825 (N_14825,N_9855,N_9406);
nand U14826 (N_14826,N_9619,N_7597);
or U14827 (N_14827,N_8329,N_7107);
and U14828 (N_14828,N_5344,N_9426);
or U14829 (N_14829,N_5510,N_5570);
nand U14830 (N_14830,N_6442,N_6043);
nand U14831 (N_14831,N_7300,N_8972);
or U14832 (N_14832,N_9339,N_8723);
or U14833 (N_14833,N_5807,N_6021);
or U14834 (N_14834,N_9895,N_6932);
or U14835 (N_14835,N_6310,N_6135);
or U14836 (N_14836,N_7613,N_9314);
or U14837 (N_14837,N_8306,N_5153);
nand U14838 (N_14838,N_7446,N_5892);
and U14839 (N_14839,N_7863,N_5214);
nor U14840 (N_14840,N_9423,N_9854);
nor U14841 (N_14841,N_7362,N_7047);
or U14842 (N_14842,N_7103,N_6413);
nor U14843 (N_14843,N_9690,N_7659);
or U14844 (N_14844,N_6526,N_6473);
and U14845 (N_14845,N_9868,N_8130);
nor U14846 (N_14846,N_5519,N_8608);
or U14847 (N_14847,N_7125,N_8136);
nor U14848 (N_14848,N_8626,N_7598);
nor U14849 (N_14849,N_9385,N_6310);
nor U14850 (N_14850,N_5191,N_9296);
nor U14851 (N_14851,N_8682,N_8551);
and U14852 (N_14852,N_6106,N_8817);
and U14853 (N_14853,N_5323,N_8208);
or U14854 (N_14854,N_9165,N_8515);
and U14855 (N_14855,N_7092,N_7543);
or U14856 (N_14856,N_6454,N_9079);
nand U14857 (N_14857,N_9449,N_7994);
or U14858 (N_14858,N_6462,N_7329);
and U14859 (N_14859,N_5772,N_8973);
or U14860 (N_14860,N_6013,N_8380);
and U14861 (N_14861,N_5092,N_9922);
nand U14862 (N_14862,N_7957,N_9697);
nand U14863 (N_14863,N_8479,N_8304);
or U14864 (N_14864,N_5902,N_9219);
nand U14865 (N_14865,N_7948,N_9163);
or U14866 (N_14866,N_7264,N_8155);
xor U14867 (N_14867,N_9942,N_8884);
and U14868 (N_14868,N_7583,N_6173);
nor U14869 (N_14869,N_5099,N_5586);
nand U14870 (N_14870,N_7323,N_9831);
nand U14871 (N_14871,N_7321,N_8718);
nand U14872 (N_14872,N_6530,N_9018);
nor U14873 (N_14873,N_9654,N_6167);
nor U14874 (N_14874,N_9319,N_8596);
nor U14875 (N_14875,N_5243,N_7300);
or U14876 (N_14876,N_5843,N_5686);
or U14877 (N_14877,N_6503,N_5031);
or U14878 (N_14878,N_6023,N_8057);
or U14879 (N_14879,N_6641,N_7719);
nor U14880 (N_14880,N_6769,N_5873);
nor U14881 (N_14881,N_7549,N_8724);
nand U14882 (N_14882,N_5429,N_9946);
nor U14883 (N_14883,N_9318,N_6723);
nand U14884 (N_14884,N_5702,N_8335);
nor U14885 (N_14885,N_5992,N_5422);
nor U14886 (N_14886,N_5544,N_5024);
nand U14887 (N_14887,N_7932,N_8609);
nor U14888 (N_14888,N_6660,N_8608);
and U14889 (N_14889,N_7468,N_8138);
nand U14890 (N_14890,N_5468,N_6458);
nand U14891 (N_14891,N_9861,N_7511);
nand U14892 (N_14892,N_8862,N_7303);
and U14893 (N_14893,N_8240,N_8818);
nor U14894 (N_14894,N_7161,N_5078);
and U14895 (N_14895,N_5972,N_7886);
and U14896 (N_14896,N_5980,N_9153);
nor U14897 (N_14897,N_5702,N_7206);
and U14898 (N_14898,N_9190,N_6092);
nor U14899 (N_14899,N_9622,N_8280);
nand U14900 (N_14900,N_6816,N_9608);
nor U14901 (N_14901,N_7011,N_9384);
nor U14902 (N_14902,N_7025,N_8500);
nor U14903 (N_14903,N_7689,N_7424);
nor U14904 (N_14904,N_6183,N_7130);
nor U14905 (N_14905,N_8715,N_5185);
or U14906 (N_14906,N_9846,N_9374);
or U14907 (N_14907,N_6581,N_7879);
and U14908 (N_14908,N_5644,N_7386);
nor U14909 (N_14909,N_5885,N_9689);
nor U14910 (N_14910,N_8874,N_7030);
nor U14911 (N_14911,N_6033,N_7238);
nor U14912 (N_14912,N_9370,N_7234);
nor U14913 (N_14913,N_8970,N_5467);
or U14914 (N_14914,N_5271,N_8906);
or U14915 (N_14915,N_6878,N_6047);
and U14916 (N_14916,N_9449,N_7633);
or U14917 (N_14917,N_8633,N_8491);
or U14918 (N_14918,N_5153,N_6055);
or U14919 (N_14919,N_5783,N_8077);
nand U14920 (N_14920,N_6212,N_5028);
and U14921 (N_14921,N_7430,N_6840);
or U14922 (N_14922,N_8807,N_7223);
or U14923 (N_14923,N_8969,N_7791);
or U14924 (N_14924,N_7765,N_8336);
and U14925 (N_14925,N_6619,N_7234);
nand U14926 (N_14926,N_7491,N_5191);
nor U14927 (N_14927,N_8323,N_7985);
nand U14928 (N_14928,N_7320,N_5995);
nand U14929 (N_14929,N_5769,N_6625);
nor U14930 (N_14930,N_7593,N_8687);
or U14931 (N_14931,N_5970,N_8100);
nor U14932 (N_14932,N_9900,N_7454);
or U14933 (N_14933,N_5166,N_9847);
nand U14934 (N_14934,N_7860,N_8066);
or U14935 (N_14935,N_6814,N_7069);
or U14936 (N_14936,N_8211,N_8212);
nand U14937 (N_14937,N_5533,N_9316);
nand U14938 (N_14938,N_8604,N_7538);
nand U14939 (N_14939,N_5968,N_9585);
xnor U14940 (N_14940,N_8129,N_5239);
or U14941 (N_14941,N_5521,N_9311);
xor U14942 (N_14942,N_5488,N_8365);
or U14943 (N_14943,N_9580,N_8775);
nand U14944 (N_14944,N_7188,N_5116);
nand U14945 (N_14945,N_9817,N_9207);
nand U14946 (N_14946,N_7788,N_6806);
and U14947 (N_14947,N_8345,N_8310);
nand U14948 (N_14948,N_6644,N_7565);
xnor U14949 (N_14949,N_8871,N_5892);
xor U14950 (N_14950,N_8853,N_5647);
nor U14951 (N_14951,N_8309,N_7898);
nor U14952 (N_14952,N_8743,N_6152);
xnor U14953 (N_14953,N_5777,N_5075);
nand U14954 (N_14954,N_8521,N_6846);
and U14955 (N_14955,N_7810,N_5358);
nand U14956 (N_14956,N_6222,N_9698);
or U14957 (N_14957,N_8690,N_9759);
and U14958 (N_14958,N_9332,N_9726);
nor U14959 (N_14959,N_6363,N_6313);
and U14960 (N_14960,N_6660,N_9759);
nand U14961 (N_14961,N_6692,N_7250);
or U14962 (N_14962,N_6809,N_5866);
nand U14963 (N_14963,N_9476,N_8570);
nor U14964 (N_14964,N_7522,N_5208);
and U14965 (N_14965,N_9301,N_8181);
xnor U14966 (N_14966,N_9972,N_5893);
and U14967 (N_14967,N_8879,N_5728);
nor U14968 (N_14968,N_6483,N_6128);
nor U14969 (N_14969,N_8005,N_9994);
nor U14970 (N_14970,N_7531,N_9807);
nand U14971 (N_14971,N_7003,N_5520);
or U14972 (N_14972,N_8946,N_9964);
nor U14973 (N_14973,N_8938,N_6448);
nand U14974 (N_14974,N_9440,N_7552);
or U14975 (N_14975,N_6165,N_9029);
or U14976 (N_14976,N_8143,N_9974);
nand U14977 (N_14977,N_9948,N_8691);
or U14978 (N_14978,N_7411,N_7000);
nand U14979 (N_14979,N_5296,N_9027);
or U14980 (N_14980,N_8414,N_5725);
nor U14981 (N_14981,N_5604,N_5502);
nand U14982 (N_14982,N_8452,N_9389);
and U14983 (N_14983,N_8650,N_8583);
nand U14984 (N_14984,N_6777,N_9200);
or U14985 (N_14985,N_5159,N_9563);
xor U14986 (N_14986,N_6366,N_6954);
nand U14987 (N_14987,N_9765,N_6962);
nand U14988 (N_14988,N_9551,N_8599);
nand U14989 (N_14989,N_8755,N_7496);
or U14990 (N_14990,N_6131,N_6514);
or U14991 (N_14991,N_8091,N_5411);
nand U14992 (N_14992,N_5431,N_9487);
and U14993 (N_14993,N_7107,N_5262);
nand U14994 (N_14994,N_8005,N_5964);
or U14995 (N_14995,N_8056,N_6320);
nand U14996 (N_14996,N_7931,N_7137);
nand U14997 (N_14997,N_5131,N_8057);
or U14998 (N_14998,N_5984,N_9844);
or U14999 (N_14999,N_8526,N_5941);
nand U15000 (N_15000,N_10707,N_14846);
nor U15001 (N_15001,N_12882,N_13195);
or U15002 (N_15002,N_14165,N_10979);
or U15003 (N_15003,N_14881,N_11608);
or U15004 (N_15004,N_11079,N_10480);
and U15005 (N_15005,N_14925,N_11324);
nand U15006 (N_15006,N_13246,N_10539);
or U15007 (N_15007,N_13788,N_12884);
and U15008 (N_15008,N_11895,N_14632);
nor U15009 (N_15009,N_11007,N_12091);
and U15010 (N_15010,N_13652,N_13638);
and U15011 (N_15011,N_14038,N_13042);
nor U15012 (N_15012,N_13587,N_14416);
nand U15013 (N_15013,N_14849,N_10090);
nor U15014 (N_15014,N_12061,N_10178);
nor U15015 (N_15015,N_12660,N_10850);
nor U15016 (N_15016,N_11149,N_10011);
nor U15017 (N_15017,N_10896,N_10150);
nand U15018 (N_15018,N_13689,N_13987);
nand U15019 (N_15019,N_14321,N_10483);
nor U15020 (N_15020,N_11517,N_10425);
nand U15021 (N_15021,N_11877,N_10558);
nor U15022 (N_15022,N_11103,N_14275);
and U15023 (N_15023,N_10730,N_13301);
nand U15024 (N_15024,N_10103,N_11991);
or U15025 (N_15025,N_14917,N_10274);
and U15026 (N_15026,N_11425,N_12519);
nor U15027 (N_15027,N_13869,N_11232);
or U15028 (N_15028,N_11521,N_11761);
or U15029 (N_15029,N_13749,N_13339);
nand U15030 (N_15030,N_12532,N_12052);
nor U15031 (N_15031,N_10864,N_12078);
nor U15032 (N_15032,N_14337,N_11543);
nand U15033 (N_15033,N_13803,N_13441);
and U15034 (N_15034,N_10547,N_12798);
or U15035 (N_15035,N_12123,N_12819);
and U15036 (N_15036,N_10886,N_12845);
and U15037 (N_15037,N_14727,N_10384);
nand U15038 (N_15038,N_13244,N_10267);
nor U15039 (N_15039,N_10841,N_11474);
and U15040 (N_15040,N_11088,N_11575);
nand U15041 (N_15041,N_13561,N_14022);
nand U15042 (N_15042,N_10486,N_11797);
xnor U15043 (N_15043,N_14793,N_12531);
nor U15044 (N_15044,N_13527,N_14529);
or U15045 (N_15045,N_11479,N_13126);
and U15046 (N_15046,N_14500,N_10438);
and U15047 (N_15047,N_10755,N_14756);
nand U15048 (N_15048,N_11291,N_12975);
xor U15049 (N_15049,N_10917,N_12121);
nand U15050 (N_15050,N_10941,N_12471);
nor U15051 (N_15051,N_12535,N_14789);
and U15052 (N_15052,N_12460,N_10897);
nor U15053 (N_15053,N_12946,N_13818);
or U15054 (N_15054,N_13815,N_12469);
nand U15055 (N_15055,N_12404,N_10359);
nor U15056 (N_15056,N_14492,N_11097);
and U15057 (N_15057,N_14675,N_11189);
and U15058 (N_15058,N_12246,N_14992);
or U15059 (N_15059,N_14041,N_10708);
or U15060 (N_15060,N_13298,N_13308);
nand U15061 (N_15061,N_10676,N_10151);
and U15062 (N_15062,N_11994,N_11059);
nand U15063 (N_15063,N_14604,N_14641);
or U15064 (N_15064,N_13020,N_14884);
nand U15065 (N_15065,N_13490,N_14096);
nand U15066 (N_15066,N_13349,N_14322);
or U15067 (N_15067,N_13306,N_14119);
or U15068 (N_15068,N_13888,N_11857);
nand U15069 (N_15069,N_14306,N_12921);
or U15070 (N_15070,N_14611,N_10299);
nor U15071 (N_15071,N_11989,N_13555);
or U15072 (N_15072,N_12634,N_11932);
or U15073 (N_15073,N_12309,N_12089);
or U15074 (N_15074,N_12082,N_12978);
or U15075 (N_15075,N_11775,N_14344);
nand U15076 (N_15076,N_12232,N_14634);
xor U15077 (N_15077,N_14290,N_14628);
and U15078 (N_15078,N_11667,N_13178);
nor U15079 (N_15079,N_12964,N_10584);
and U15080 (N_15080,N_13105,N_11518);
and U15081 (N_15081,N_13094,N_14436);
nor U15082 (N_15082,N_13607,N_10024);
xnor U15083 (N_15083,N_14484,N_13680);
nor U15084 (N_15084,N_10382,N_12437);
or U15085 (N_15085,N_12735,N_10181);
nor U15086 (N_15086,N_11366,N_12979);
and U15087 (N_15087,N_11781,N_10732);
nand U15088 (N_15088,N_11592,N_12158);
or U15089 (N_15089,N_12347,N_14020);
nand U15090 (N_15090,N_13943,N_12777);
nand U15091 (N_15091,N_10750,N_12252);
nor U15092 (N_15092,N_11036,N_12141);
and U15093 (N_15093,N_11794,N_13789);
nand U15094 (N_15094,N_13808,N_11656);
nand U15095 (N_15095,N_11125,N_14482);
nand U15096 (N_15096,N_13725,N_10672);
nor U15097 (N_15097,N_13332,N_13025);
nor U15098 (N_15098,N_14470,N_12705);
nand U15099 (N_15099,N_14569,N_14490);
and U15100 (N_15100,N_12062,N_11185);
nor U15101 (N_15101,N_10350,N_10155);
or U15102 (N_15102,N_13731,N_14378);
nand U15103 (N_15103,N_12666,N_11420);
and U15104 (N_15104,N_10507,N_14832);
or U15105 (N_15105,N_12920,N_11634);
and U15106 (N_15106,N_12372,N_11936);
nor U15107 (N_15107,N_10461,N_14260);
nor U15108 (N_15108,N_10798,N_13641);
nor U15109 (N_15109,N_14230,N_12301);
or U15110 (N_15110,N_11198,N_10809);
nand U15111 (N_15111,N_13872,N_14910);
or U15112 (N_15112,N_12569,N_14718);
nor U15113 (N_15113,N_13068,N_13996);
nand U15114 (N_15114,N_12354,N_13820);
or U15115 (N_15115,N_14983,N_10124);
nor U15116 (N_15116,N_10948,N_11567);
and U15117 (N_15117,N_13035,N_14002);
or U15118 (N_15118,N_10981,N_10426);
nand U15119 (N_15119,N_12891,N_10143);
nand U15120 (N_15120,N_14764,N_14315);
nor U15121 (N_15121,N_12412,N_12813);
nor U15122 (N_15122,N_10934,N_11325);
xnor U15123 (N_15123,N_11524,N_10926);
nand U15124 (N_15124,N_13645,N_14562);
and U15125 (N_15125,N_13464,N_14738);
nor U15126 (N_15126,N_14618,N_10504);
nor U15127 (N_15127,N_13054,N_11942);
xnor U15128 (N_15128,N_13253,N_13959);
nand U15129 (N_15129,N_11636,N_12972);
or U15130 (N_15130,N_14352,N_13843);
or U15131 (N_15131,N_10806,N_11742);
nand U15132 (N_15132,N_13770,N_14144);
nor U15133 (N_15133,N_10451,N_11265);
and U15134 (N_15134,N_11744,N_14204);
nand U15135 (N_15135,N_10478,N_14769);
or U15136 (N_15136,N_11136,N_10751);
or U15137 (N_15137,N_13595,N_10249);
nand U15138 (N_15138,N_14535,N_12317);
nand U15139 (N_15139,N_12572,N_12299);
nand U15140 (N_15140,N_10420,N_12326);
or U15141 (N_15141,N_12425,N_10332);
nor U15142 (N_15142,N_14081,N_12983);
nor U15143 (N_15143,N_12403,N_14036);
nand U15144 (N_15144,N_12844,N_10639);
or U15145 (N_15145,N_10530,N_11838);
nor U15146 (N_15146,N_10235,N_10596);
and U15147 (N_15147,N_12654,N_11293);
nand U15148 (N_15148,N_14539,N_14148);
nor U15149 (N_15149,N_10745,N_11261);
nor U15150 (N_15150,N_11078,N_12609);
nor U15151 (N_15151,N_11555,N_10497);
nor U15152 (N_15152,N_12670,N_11760);
or U15153 (N_15153,N_13963,N_12594);
nand U15154 (N_15154,N_10920,N_12216);
and U15155 (N_15155,N_11464,N_12671);
nand U15156 (N_15156,N_10622,N_14391);
nand U15157 (N_15157,N_11536,N_13717);
or U15158 (N_15158,N_14737,N_13708);
xnor U15159 (N_15159,N_14661,N_12318);
nor U15160 (N_15160,N_11999,N_14596);
nor U15161 (N_15161,N_11685,N_14763);
or U15162 (N_15162,N_11066,N_10354);
nor U15163 (N_15163,N_11514,N_13227);
nor U15164 (N_15164,N_13915,N_14198);
nor U15165 (N_15165,N_14015,N_12218);
or U15166 (N_15166,N_13034,N_12831);
nor U15167 (N_15167,N_14307,N_12570);
nand U15168 (N_15168,N_12247,N_14221);
and U15169 (N_15169,N_11174,N_12533);
and U15170 (N_15170,N_10921,N_12868);
nand U15171 (N_15171,N_13406,N_12416);
or U15172 (N_15172,N_11746,N_13488);
or U15173 (N_15173,N_13416,N_14501);
and U15174 (N_15174,N_11154,N_11448);
nand U15175 (N_15175,N_14725,N_12370);
nor U15176 (N_15176,N_12643,N_11844);
and U15177 (N_15177,N_10375,N_11616);
nand U15178 (N_15178,N_11475,N_12626);
nand U15179 (N_15179,N_13209,N_10071);
nand U15180 (N_15180,N_12663,N_13995);
nor U15181 (N_15181,N_14220,N_14396);
and U15182 (N_15182,N_11571,N_10265);
nand U15183 (N_15183,N_12811,N_14493);
nor U15184 (N_15184,N_13266,N_10889);
nor U15185 (N_15185,N_14018,N_12342);
nor U15186 (N_15186,N_12542,N_12915);
nand U15187 (N_15187,N_14605,N_14049);
and U15188 (N_15188,N_12363,N_10070);
and U15189 (N_15189,N_10693,N_12615);
and U15190 (N_15190,N_12332,N_14991);
or U15191 (N_15191,N_11166,N_11032);
or U15192 (N_15192,N_14751,N_10187);
xor U15193 (N_15193,N_14229,N_11600);
nand U15194 (N_15194,N_12140,N_11723);
or U15195 (N_15195,N_12480,N_10522);
nand U15196 (N_15196,N_14366,N_14726);
and U15197 (N_15197,N_13117,N_12076);
or U15198 (N_15198,N_10300,N_11418);
nor U15199 (N_15199,N_12011,N_13955);
or U15200 (N_15200,N_13546,N_13424);
nand U15201 (N_15201,N_10524,N_11345);
nand U15202 (N_15202,N_11308,N_11453);
and U15203 (N_15203,N_10959,N_12970);
or U15204 (N_15204,N_11463,N_13296);
nand U15205 (N_15205,N_13316,N_12649);
or U15206 (N_15206,N_14948,N_13055);
and U15207 (N_15207,N_10797,N_10978);
or U15208 (N_15208,N_10456,N_10125);
nand U15209 (N_15209,N_13153,N_12652);
nand U15210 (N_15210,N_14570,N_12438);
and U15211 (N_15211,N_11181,N_12459);
or U15212 (N_15212,N_10554,N_11708);
nor U15213 (N_15213,N_13163,N_14234);
nor U15214 (N_15214,N_12830,N_11827);
nor U15215 (N_15215,N_12439,N_12719);
nor U15216 (N_15216,N_14784,N_11491);
nor U15217 (N_15217,N_14298,N_13685);
and U15218 (N_15218,N_12579,N_12406);
nor U15219 (N_15219,N_12548,N_10421);
nand U15220 (N_15220,N_14058,N_12431);
nand U15221 (N_15221,N_10092,N_14263);
nand U15222 (N_15222,N_13252,N_10469);
nor U15223 (N_15223,N_14467,N_10659);
or U15224 (N_15224,N_10073,N_12485);
nor U15225 (N_15225,N_12068,N_10351);
or U15226 (N_15226,N_13033,N_11916);
nand U15227 (N_15227,N_12717,N_11752);
and U15228 (N_15228,N_13567,N_10418);
nor U15229 (N_15229,N_12527,N_11573);
or U15230 (N_15230,N_12242,N_10966);
nor U15231 (N_15231,N_11964,N_11480);
and U15232 (N_15232,N_12185,N_10819);
nand U15233 (N_15233,N_14131,N_11043);
nand U15234 (N_15234,N_10410,N_13192);
or U15235 (N_15235,N_11628,N_14936);
and U15236 (N_15236,N_14888,N_13554);
nand U15237 (N_15237,N_11510,N_11559);
nand U15238 (N_15238,N_11651,N_12494);
nor U15239 (N_15239,N_10313,N_13081);
nor U15240 (N_15240,N_13695,N_11664);
nor U15241 (N_15241,N_12873,N_13201);
nor U15242 (N_15242,N_11386,N_14226);
and U15243 (N_15243,N_11789,N_13141);
nor U15244 (N_15244,N_11963,N_12487);
nand U15245 (N_15245,N_14214,N_12588);
nor U15246 (N_15246,N_14957,N_14410);
and U15247 (N_15247,N_13364,N_12266);
and U15248 (N_15248,N_14671,N_11210);
and U15249 (N_15249,N_14346,N_10029);
nor U15250 (N_15250,N_14816,N_12545);
nand U15251 (N_15251,N_13103,N_13040);
xnor U15252 (N_15252,N_11176,N_11428);
nand U15253 (N_15253,N_10520,N_11579);
or U15254 (N_15254,N_11186,N_11866);
and U15255 (N_15255,N_13707,N_14474);
and U15256 (N_15256,N_14944,N_13916);
nor U15257 (N_15257,N_12550,N_11973);
nand U15258 (N_15258,N_10457,N_10053);
nand U15259 (N_15259,N_14898,N_14614);
nor U15260 (N_15260,N_11143,N_12506);
nand U15261 (N_15261,N_12708,N_12781);
nor U15262 (N_15262,N_10165,N_11644);
nand U15263 (N_15263,N_10587,N_13484);
and U15264 (N_15264,N_11687,N_13357);
and U15265 (N_15265,N_14567,N_10996);
or U15266 (N_15266,N_11701,N_13615);
nor U15267 (N_15267,N_10719,N_12820);
or U15268 (N_15268,N_13966,N_10454);
and U15269 (N_15269,N_14664,N_12986);
nor U15270 (N_15270,N_12784,N_10314);
or U15271 (N_15271,N_14739,N_12623);
or U15272 (N_15272,N_10834,N_11710);
and U15273 (N_15273,N_10091,N_12380);
nand U15274 (N_15274,N_11669,N_10845);
nor U15275 (N_15275,N_14357,N_14340);
nand U15276 (N_15276,N_10813,N_13400);
and U15277 (N_15277,N_11019,N_14025);
or U15278 (N_15278,N_10127,N_13714);
nand U15279 (N_15279,N_11888,N_14033);
nand U15280 (N_15280,N_10684,N_10414);
and U15281 (N_15281,N_13097,N_10863);
or U15282 (N_15282,N_11676,N_11028);
nand U15283 (N_15283,N_14892,N_14358);
or U15284 (N_15284,N_14776,N_14172);
or U15285 (N_15285,N_12357,N_10177);
and U15286 (N_15286,N_14456,N_11828);
or U15287 (N_15287,N_10339,N_14120);
and U15288 (N_15288,N_11487,N_11894);
nor U15289 (N_15289,N_10213,N_12418);
nor U15290 (N_15290,N_10821,N_13350);
nor U15291 (N_15291,N_13190,N_12413);
nand U15292 (N_15292,N_11163,N_14981);
nor U15293 (N_15293,N_12286,N_13367);
and U15294 (N_15294,N_11605,N_13860);
xnor U15295 (N_15295,N_10573,N_11326);
nand U15296 (N_15296,N_14714,N_11422);
and U15297 (N_15297,N_13128,N_14394);
or U15298 (N_15298,N_13404,N_11743);
nor U15299 (N_15299,N_11037,N_12270);
or U15300 (N_15300,N_14415,N_10785);
nand U15301 (N_15301,N_12192,N_12573);
nand U15302 (N_15302,N_14259,N_11812);
nand U15303 (N_15303,N_11587,N_11411);
or U15304 (N_15304,N_14913,N_10439);
nor U15305 (N_15305,N_14195,N_12024);
or U15306 (N_15306,N_13620,N_10895);
nand U15307 (N_15307,N_10860,N_11945);
and U15308 (N_15308,N_11388,N_14463);
and U15309 (N_15309,N_10471,N_13745);
and U15310 (N_15310,N_13057,N_12990);
nor U15311 (N_15311,N_10188,N_13886);
nor U15312 (N_15312,N_12033,N_10197);
nand U15313 (N_15313,N_13239,N_14351);
or U15314 (N_15314,N_14046,N_14767);
nor U15315 (N_15315,N_11550,N_11279);
nand U15316 (N_15316,N_11909,N_13071);
or U15317 (N_15317,N_10361,N_12248);
and U15318 (N_15318,N_10973,N_12849);
nor U15319 (N_15319,N_14329,N_13011);
and U15320 (N_15320,N_10085,N_14543);
nor U15321 (N_15321,N_10328,N_13275);
nand U15322 (N_15322,N_12650,N_13323);
or U15323 (N_15323,N_10465,N_12441);
nand U15324 (N_15324,N_10319,N_13376);
nor U15325 (N_15325,N_13131,N_10556);
or U15326 (N_15326,N_14920,N_13841);
nand U15327 (N_15327,N_13670,N_12563);
nor U15328 (N_15328,N_10263,N_14274);
and U15329 (N_15329,N_10320,N_10799);
and U15330 (N_15330,N_12906,N_12848);
nor U15331 (N_15331,N_14194,N_14869);
nor U15332 (N_15332,N_10650,N_11852);
or U15333 (N_15333,N_14496,N_11635);
nand U15334 (N_15334,N_13315,N_11026);
nor U15335 (N_15335,N_14573,N_12585);
nand U15336 (N_15336,N_11488,N_13528);
or U15337 (N_15337,N_12835,N_14525);
nand U15338 (N_15338,N_12738,N_11531);
nor U15339 (N_15339,N_12327,N_10142);
xnor U15340 (N_15340,N_10336,N_11557);
nand U15341 (N_15341,N_12281,N_14222);
nor U15342 (N_15342,N_12751,N_14114);
nor U15343 (N_15343,N_14538,N_10972);
xor U15344 (N_15344,N_12324,N_13063);
and U15345 (N_15345,N_11642,N_11609);
nand U15346 (N_15346,N_10673,N_11251);
and U15347 (N_15347,N_11465,N_13372);
or U15348 (N_15348,N_11900,N_14365);
or U15349 (N_15349,N_14791,N_13050);
and U15350 (N_15350,N_11530,N_11489);
nand U15351 (N_15351,N_10166,N_10131);
or U15352 (N_15352,N_11823,N_14093);
nor U15353 (N_15353,N_11193,N_12925);
or U15354 (N_15354,N_14476,N_13876);
and U15355 (N_15355,N_10407,N_11572);
and U15356 (N_15356,N_13728,N_14199);
or U15357 (N_15357,N_11560,N_11100);
nor U15358 (N_15358,N_12178,N_12551);
or U15359 (N_15359,N_11228,N_13656);
and U15360 (N_15360,N_14838,N_14609);
or U15361 (N_15361,N_10731,N_14950);
and U15362 (N_15362,N_13145,N_13241);
or U15363 (N_15363,N_12050,N_12887);
nand U15364 (N_15364,N_13008,N_14963);
nand U15365 (N_15365,N_12116,N_10565);
or U15366 (N_15366,N_13973,N_14056);
and U15367 (N_15367,N_10932,N_13969);
nor U15368 (N_15368,N_13385,N_10066);
nand U15369 (N_15369,N_14061,N_10583);
and U15370 (N_15370,N_10180,N_13880);
and U15371 (N_15371,N_13526,N_12175);
nor U15372 (N_15372,N_14808,N_12361);
nor U15373 (N_15373,N_11309,N_10427);
nor U15374 (N_15374,N_12943,N_10893);
or U15375 (N_15375,N_13925,N_10710);
nor U15376 (N_15376,N_12904,N_13785);
and U15377 (N_15377,N_10153,N_14741);
nor U15378 (N_15378,N_13868,N_12228);
nor U15379 (N_15379,N_14548,N_11061);
or U15380 (N_15380,N_14746,N_10881);
nor U15381 (N_15381,N_10636,N_10511);
and U15382 (N_15382,N_12478,N_10723);
or U15383 (N_15383,N_14870,N_14108);
and U15384 (N_15384,N_12155,N_14680);
and U15385 (N_15385,N_12893,N_11498);
nor U15386 (N_15386,N_11564,N_12842);
or U15387 (N_15387,N_13511,N_10116);
nor U15388 (N_15388,N_14028,N_10388);
nor U15389 (N_15389,N_11358,N_12522);
and U15390 (N_15390,N_11831,N_14999);
nand U15391 (N_15391,N_12465,N_14742);
nor U15392 (N_15392,N_14928,N_12935);
nand U15393 (N_15393,N_11796,N_13061);
and U15394 (N_15394,N_12631,N_13148);
nand U15395 (N_15395,N_12992,N_14672);
or U15396 (N_15396,N_13550,N_13751);
nor U15397 (N_15397,N_13643,N_13772);
and U15398 (N_15398,N_12696,N_14778);
or U15399 (N_15399,N_13047,N_13510);
nor U15400 (N_15400,N_12768,N_14129);
nor U15401 (N_15401,N_11627,N_12422);
or U15402 (N_15402,N_10543,N_10324);
nand U15403 (N_15403,N_12463,N_11639);
or U15404 (N_15404,N_12328,N_11224);
or U15405 (N_15405,N_13090,N_12960);
or U15406 (N_15406,N_11933,N_14276);
nand U15407 (N_15407,N_10301,N_12368);
nand U15408 (N_15408,N_14123,N_14674);
or U15409 (N_15409,N_11834,N_10399);
nand U15410 (N_15410,N_14635,N_10744);
nand U15411 (N_15411,N_12190,N_13563);
nand U15412 (N_15412,N_13474,N_14430);
nand U15413 (N_15413,N_10276,N_10967);
or U15414 (N_15414,N_13478,N_13965);
or U15415 (N_15415,N_10129,N_12988);
nor U15416 (N_15416,N_13724,N_11859);
nor U15417 (N_15417,N_11092,N_10876);
nand U15418 (N_15418,N_13109,N_11268);
and U15419 (N_15419,N_13814,N_13476);
nor U15420 (N_15420,N_14524,N_11625);
nor U15421 (N_15421,N_11603,N_14942);
and U15422 (N_15422,N_10856,N_14255);
and U15423 (N_15423,N_13056,N_11696);
or U15424 (N_15424,N_12322,N_11034);
and U15425 (N_15425,N_12809,N_10479);
nor U15426 (N_15426,N_10431,N_13505);
or U15427 (N_15427,N_13425,N_13083);
and U15428 (N_15428,N_12343,N_11558);
nand U15429 (N_15429,N_13032,N_12795);
and U15430 (N_15430,N_13794,N_11093);
xor U15431 (N_15431,N_14853,N_14083);
or U15432 (N_15432,N_10588,N_13979);
nor U15433 (N_15433,N_13358,N_12118);
nand U15434 (N_15434,N_13375,N_10642);
nor U15435 (N_15435,N_13194,N_11926);
nand U15436 (N_15436,N_13233,N_14914);
nor U15437 (N_15437,N_14292,N_13447);
nor U15438 (N_15438,N_10904,N_12641);
nor U15439 (N_15439,N_10088,N_14821);
nand U15440 (N_15440,N_11009,N_11469);
nor U15441 (N_15441,N_12358,N_12423);
nor U15442 (N_15442,N_13743,N_13181);
or U15443 (N_15443,N_14937,N_12702);
nand U15444 (N_15444,N_13283,N_12310);
or U15445 (N_15445,N_14085,N_12307);
and U15446 (N_15446,N_12664,N_11912);
nand U15447 (N_15447,N_14115,N_12734);
or U15448 (N_15448,N_14440,N_13921);
nand U15449 (N_15449,N_14502,N_13512);
nand U15450 (N_15450,N_13041,N_12941);
or U15451 (N_15451,N_12231,N_10726);
nor U15452 (N_15452,N_12329,N_11306);
or U15453 (N_15453,N_10331,N_14972);
nor U15454 (N_15454,N_10849,N_10297);
nor U15455 (N_15455,N_10638,N_12775);
nor U15456 (N_15456,N_13417,N_13971);
nand U15457 (N_15457,N_12864,N_11731);
nand U15458 (N_15458,N_13154,N_11652);
nor U15459 (N_15459,N_13051,N_14062);
and U15460 (N_15460,N_11538,N_12040);
and U15461 (N_15461,N_13377,N_11956);
and U15462 (N_15462,N_12698,N_14241);
nor U15463 (N_15463,N_10575,N_12264);
nand U15464 (N_15464,N_11172,N_12790);
nor U15465 (N_15465,N_14556,N_13191);
nor U15466 (N_15466,N_11661,N_11599);
and U15467 (N_15467,N_12742,N_13562);
and U15468 (N_15468,N_13345,N_12337);
nand U15469 (N_15469,N_13968,N_10599);
or U15470 (N_15470,N_11363,N_14600);
nand U15471 (N_15471,N_10990,N_12740);
nor U15472 (N_15472,N_12818,N_12097);
xor U15473 (N_15473,N_12929,N_14079);
nand U15474 (N_15474,N_11180,N_12729);
or U15475 (N_15475,N_11212,N_10526);
or U15476 (N_15476,N_10112,N_13009);
nand U15477 (N_15477,N_12381,N_11131);
nand U15478 (N_15478,N_11348,N_13300);
and U15479 (N_15479,N_11004,N_10724);
or U15480 (N_15480,N_13104,N_12171);
and U15481 (N_15481,N_13964,N_14401);
nor U15482 (N_15482,N_11987,N_11606);
and U15483 (N_15483,N_11581,N_11076);
nor U15484 (N_15484,N_11477,N_11540);
nand U15485 (N_15485,N_13781,N_10488);
xnor U15486 (N_15486,N_11523,N_10464);
nor U15487 (N_15487,N_11449,N_14031);
nor U15488 (N_15488,N_10458,N_12184);
and U15489 (N_15489,N_14927,N_14954);
nand U15490 (N_15490,N_13100,N_13713);
nand U15491 (N_15491,N_13867,N_11774);
nand U15492 (N_15492,N_13204,N_11984);
nand U15493 (N_15493,N_11944,N_12870);
nor U15494 (N_15494,N_11275,N_10548);
or U15495 (N_15495,N_14959,N_14804);
nor U15496 (N_15496,N_11638,N_14794);
or U15497 (N_15497,N_10670,N_14616);
and U15498 (N_15498,N_10035,N_11757);
nand U15499 (N_15499,N_12792,N_10219);
or U15500 (N_15500,N_14312,N_12353);
nor U15501 (N_15501,N_10545,N_13402);
nor U15502 (N_15502,N_14906,N_10859);
and U15503 (N_15503,N_14135,N_12267);
or U15504 (N_15504,N_10843,N_11191);
nand U15505 (N_15505,N_13887,N_14281);
nand U15506 (N_15506,N_10623,N_14886);
nand U15507 (N_15507,N_13477,N_10620);
nand U15508 (N_15508,N_13184,N_13762);
or U15509 (N_15509,N_10585,N_12796);
nand U15510 (N_15510,N_10725,N_14182);
xnor U15511 (N_15511,N_12457,N_14174);
and U15512 (N_15512,N_12985,N_12797);
or U15513 (N_15513,N_14691,N_10003);
and U15514 (N_15514,N_10325,N_10466);
or U15515 (N_15515,N_13366,N_13462);
or U15516 (N_15516,N_12420,N_13170);
xnor U15517 (N_15517,N_14113,N_13458);
nor U15518 (N_15518,N_10244,N_12182);
and U15519 (N_15519,N_12238,N_12203);
or U15520 (N_15520,N_12396,N_11378);
nand U15521 (N_15521,N_14795,N_10930);
and U15522 (N_15522,N_13898,N_13648);
or U15523 (N_15523,N_13928,N_11533);
nand U15524 (N_15524,N_14404,N_12869);
or U15525 (N_15525,N_12791,N_12825);
or U15526 (N_15526,N_10657,N_14318);
and U15527 (N_15527,N_12598,N_13368);
and U15528 (N_15528,N_11207,N_11883);
and U15529 (N_15529,N_10688,N_14151);
nor U15530 (N_15530,N_13370,N_14783);
nor U15531 (N_15531,N_10812,N_14342);
and U15532 (N_15532,N_14095,N_13065);
and U15533 (N_15533,N_10563,N_10191);
or U15534 (N_15534,N_10519,N_12359);
nand U15535 (N_15535,N_14681,N_11904);
nand U15536 (N_15536,N_12005,N_14405);
and U15537 (N_15537,N_13088,N_14949);
nor U15538 (N_15538,N_12201,N_14111);
nand U15539 (N_15539,N_11173,N_11853);
xnor U15540 (N_15540,N_10682,N_11720);
nor U15541 (N_15541,N_14400,N_13859);
nor U15542 (N_15542,N_10064,N_13858);
nand U15543 (N_15543,N_13577,N_10551);
nand U15544 (N_15544,N_13830,N_12400);
or U15545 (N_15545,N_14943,N_13530);
or U15546 (N_15546,N_14044,N_14164);
nor U15547 (N_15547,N_12648,N_13304);
nand U15548 (N_15548,N_14277,N_13588);
nand U15549 (N_15549,N_12220,N_11370);
and U15550 (N_15550,N_13014,N_10355);
and U15551 (N_15551,N_10965,N_13337);
nor U15552 (N_15552,N_14460,N_13470);
nor U15553 (N_15553,N_11484,N_12607);
nand U15554 (N_15554,N_10847,N_13624);
nor U15555 (N_15555,N_10572,N_10374);
nand U15556 (N_15556,N_11225,N_10065);
nand U15557 (N_15557,N_11927,N_12567);
nor U15558 (N_15558,N_14597,N_12442);
nand U15559 (N_15559,N_14373,N_10618);
nor U15560 (N_15560,N_12086,N_11421);
or U15561 (N_15561,N_13452,N_12510);
and U15562 (N_15562,N_11582,N_10341);
or U15563 (N_15563,N_11740,N_11056);
and U15564 (N_15564,N_13908,N_11021);
or U15565 (N_15565,N_14868,N_12564);
nand U15566 (N_15566,N_14390,N_10184);
and U15567 (N_15567,N_12502,N_13531);
nor U15568 (N_15568,N_13970,N_14703);
nor U15569 (N_15569,N_13384,N_10696);
or U15570 (N_15570,N_13242,N_10894);
nor U15571 (N_15571,N_11898,N_13164);
or U15572 (N_15572,N_14625,N_14825);
or U15573 (N_15573,N_12892,N_11862);
and U15574 (N_15574,N_10352,N_13824);
nand U15575 (N_15575,N_14409,N_10308);
nand U15576 (N_15576,N_14708,N_14433);
nand U15577 (N_15577,N_14006,N_14439);
or U15578 (N_15578,N_14707,N_13834);
nand U15579 (N_15579,N_12454,N_13580);
nor U15580 (N_15580,N_11003,N_11881);
or U15581 (N_15581,N_13015,N_13334);
or U15582 (N_15582,N_14988,N_12046);
or U15583 (N_15583,N_11201,N_13193);
nor U15584 (N_15584,N_13619,N_12914);
nor U15585 (N_15585,N_10216,N_13962);
nor U15586 (N_15586,N_11017,N_14117);
nand U15587 (N_15587,N_14677,N_12265);
or U15588 (N_15588,N_14986,N_13268);
nor U15589 (N_15589,N_13712,N_12449);
nor U15590 (N_15590,N_14237,N_11594);
or U15591 (N_15591,N_12489,N_13092);
nand U15592 (N_15592,N_10433,N_12130);
or U15593 (N_15593,N_14421,N_10617);
nor U15594 (N_15594,N_11072,N_10635);
or U15595 (N_15595,N_11450,N_13396);
nor U15596 (N_15596,N_12889,N_13292);
and U15597 (N_15597,N_11156,N_10646);
and U15598 (N_15598,N_13175,N_11184);
nand U15599 (N_15599,N_12805,N_11492);
nor U15600 (N_15600,N_12894,N_10923);
nand U15601 (N_15601,N_11246,N_10287);
nand U15602 (N_15602,N_11057,N_14455);
nor U15603 (N_15603,N_12803,N_12240);
xnor U15604 (N_15604,N_12612,N_13070);
nand U15605 (N_15605,N_11300,N_12067);
nor U15606 (N_15606,N_14297,N_11040);
or U15607 (N_15607,N_10515,N_13983);
nand U15608 (N_15608,N_13307,N_14376);
nand U15609 (N_15609,N_10260,N_11229);
and U15610 (N_15610,N_10097,N_12838);
nor U15611 (N_15611,N_10322,N_12346);
nand U15612 (N_15612,N_12377,N_11042);
or U15613 (N_15613,N_11373,N_13353);
and U15614 (N_15614,N_10109,N_12365);
nor U15615 (N_15615,N_10608,N_12908);
and U15616 (N_15616,N_13741,N_11120);
nor U15617 (N_15617,N_13517,N_10409);
nand U15618 (N_15618,N_11045,N_13395);
or U15619 (N_15619,N_13024,N_14434);
nand U15620 (N_15620,N_11882,N_13294);
nor U15621 (N_15621,N_12701,N_10018);
nor U15622 (N_15622,N_12503,N_11457);
nand U15623 (N_15623,N_13213,N_10424);
nor U15624 (N_15624,N_11126,N_14660);
and U15625 (N_15625,N_13285,N_13997);
nand U15626 (N_15626,N_11493,N_13545);
or U15627 (N_15627,N_11458,N_10641);
nor U15628 (N_15628,N_14282,N_10735);
nor U15629 (N_15629,N_11169,N_10467);
or U15630 (N_15630,N_13778,N_10911);
nand U15631 (N_15631,N_12526,N_13625);
nand U15632 (N_15632,N_10423,N_13091);
nand U15633 (N_15633,N_12000,N_13074);
or U15634 (N_15634,N_14598,N_14658);
nand U15635 (N_15635,N_14235,N_12073);
or U15636 (N_15636,N_14447,N_12684);
nand U15637 (N_15637,N_10402,N_10256);
nand U15638 (N_15638,N_11698,N_12071);
and U15639 (N_15639,N_13922,N_10746);
and U15640 (N_15640,N_13207,N_11055);
nor U15641 (N_15641,N_12755,N_11892);
and U15642 (N_15642,N_12720,N_14679);
or U15643 (N_15643,N_12589,N_12679);
or U15644 (N_15644,N_10273,N_13176);
or U15645 (N_15645,N_10517,N_10387);
or U15646 (N_15646,N_13838,N_14005);
nor U15647 (N_15647,N_14722,N_10010);
or U15648 (N_15648,N_13479,N_11890);
nor U15649 (N_15649,N_14491,N_12758);
and U15650 (N_15650,N_12208,N_10416);
nor U15651 (N_15651,N_10280,N_12922);
nor U15652 (N_15652,N_14498,N_14700);
or U15653 (N_15653,N_10916,N_13939);
and U15654 (N_15654,N_14379,N_14454);
and U15655 (N_15655,N_13934,N_11875);
or U15656 (N_15656,N_10110,N_10626);
nand U15657 (N_15657,N_12298,N_10811);
or U15658 (N_15658,N_13821,N_13635);
nor U15659 (N_15659,N_13355,N_11347);
and U15660 (N_15660,N_11706,N_12749);
or U15661 (N_15661,N_13115,N_12305);
nand U15662 (N_15662,N_13114,N_11663);
and U15663 (N_15663,N_10228,N_10801);
nand U15664 (N_15664,N_12219,N_13212);
and U15665 (N_15665,N_11955,N_10518);
and U15666 (N_15666,N_10292,N_10481);
nor U15667 (N_15667,N_13668,N_13409);
and U15668 (N_15668,N_11342,N_10428);
or U15669 (N_15669,N_12910,N_10562);
nand U15670 (N_15670,N_12516,N_14966);
nand U15671 (N_15671,N_13151,N_14513);
and U15672 (N_15672,N_14760,N_13284);
nor U15673 (N_15673,N_12014,N_11285);
and U15674 (N_15674,N_13492,N_14110);
nand U15675 (N_15675,N_11058,N_11715);
and U15676 (N_15676,N_11085,N_10113);
and U15677 (N_15677,N_11241,N_12167);
and U15678 (N_15678,N_10510,N_14852);
or U15679 (N_15679,N_11541,N_10289);
xnor U15680 (N_15680,N_10323,N_11943);
and U15681 (N_15681,N_11335,N_13875);
nor U15682 (N_15682,N_10302,N_11522);
nor U15683 (N_15683,N_14377,N_10330);
nand U15684 (N_15684,N_10829,N_12136);
nor U15685 (N_15685,N_10381,N_12428);
nand U15686 (N_15686,N_10012,N_12006);
or U15687 (N_15687,N_11133,N_11404);
or U15688 (N_15688,N_10647,N_10961);
or U15689 (N_15689,N_14800,N_12254);
nor U15690 (N_15690,N_14313,N_14995);
or U15691 (N_15691,N_10861,N_13519);
nor U15692 (N_15692,N_12297,N_12829);
nand U15693 (N_15693,N_12592,N_10942);
or U15694 (N_15694,N_14353,N_12967);
nor U15695 (N_15695,N_11481,N_14850);
and U15696 (N_15696,N_11135,N_12854);
xnor U15697 (N_15697,N_13581,N_12763);
or U15698 (N_15698,N_14781,N_10760);
nor U15699 (N_15699,N_12157,N_10614);
or U15700 (N_15700,N_14029,N_12898);
nand U15701 (N_15701,N_11902,N_10233);
and U15702 (N_15702,N_10363,N_12711);
nor U15703 (N_15703,N_14997,N_10223);
nand U15704 (N_15704,N_12639,N_12655);
xnor U15705 (N_15705,N_13658,N_10753);
and U15706 (N_15706,N_11730,N_12374);
nor U15707 (N_15707,N_12277,N_12291);
nor U15708 (N_15708,N_13744,N_13801);
nor U15709 (N_15709,N_12843,N_10303);
or U15710 (N_15710,N_10777,N_12674);
nor U15711 (N_15711,N_10241,N_13953);
nand U15712 (N_15712,N_10021,N_10063);
and U15713 (N_15713,N_12602,N_13263);
nor U15714 (N_15714,N_12042,N_14228);
and U15715 (N_15715,N_11159,N_10705);
nor U15716 (N_15716,N_11817,N_10200);
or U15717 (N_15717,N_13631,N_12392);
or U15718 (N_15718,N_14127,N_12080);
and U15719 (N_15719,N_12129,N_10586);
or U15720 (N_15720,N_10913,N_14650);
nand U15721 (N_15721,N_13759,N_13799);
and U15722 (N_15722,N_13499,N_14566);
nand U15723 (N_15723,N_10591,N_10203);
nor U15724 (N_15724,N_14951,N_14375);
nor U15725 (N_15725,N_10880,N_12872);
nor U15726 (N_15726,N_14797,N_10908);
and U15727 (N_15727,N_11873,N_12625);
or U15728 (N_15728,N_11295,N_12362);
or U15729 (N_15729,N_14530,N_12239);
nand U15730 (N_15730,N_12741,N_10581);
nor U15731 (N_15731,N_13999,N_12117);
and U15732 (N_15732,N_12765,N_10174);
or U15733 (N_15733,N_10275,N_12477);
nor U15734 (N_15734,N_13613,N_14413);
and U15735 (N_15735,N_13984,N_13754);
or U15736 (N_15736,N_13445,N_12261);
or U15737 (N_15737,N_10043,N_11977);
or U15738 (N_15738,N_10603,N_13792);
nand U15739 (N_15739,N_11784,N_10578);
xnor U15740 (N_15740,N_14291,N_13463);
nor U15741 (N_15741,N_11960,N_11433);
and U15742 (N_15742,N_14283,N_13264);
or U15743 (N_15743,N_14240,N_11301);
nand U15744 (N_15744,N_11033,N_14251);
nor U15745 (N_15745,N_12308,N_13427);
and U15746 (N_15746,N_11833,N_12287);
nor U15747 (N_15747,N_10261,N_13585);
or U15748 (N_15748,N_13281,N_13551);
nand U15749 (N_15749,N_11561,N_12681);
and U15750 (N_15750,N_14941,N_14126);
nor U15751 (N_15751,N_14730,N_11068);
nor U15752 (N_15752,N_14626,N_10660);
and U15753 (N_15753,N_11138,N_13440);
or U15754 (N_15754,N_10159,N_13177);
and U15755 (N_15755,N_13782,N_11741);
nor U15756 (N_15756,N_14897,N_11736);
nor U15757 (N_15757,N_13256,N_14035);
or U15758 (N_15758,N_10195,N_10905);
nor U15759 (N_15759,N_10312,N_13132);
or U15760 (N_15760,N_14623,N_14406);
or U15761 (N_15761,N_10827,N_10900);
nand U15762 (N_15762,N_10500,N_12895);
or U15763 (N_15763,N_14961,N_12924);
or U15764 (N_15764,N_10815,N_13544);
and U15765 (N_15765,N_10513,N_13753);
and U15766 (N_15766,N_10619,N_14330);
nor U15767 (N_15767,N_12804,N_12806);
or U15768 (N_15768,N_13633,N_10277);
or U15769 (N_15769,N_14422,N_11070);
and U15770 (N_15770,N_12070,N_12222);
or U15771 (N_15771,N_10814,N_10080);
and U15772 (N_15772,N_11473,N_13681);
nand U15773 (N_15773,N_12360,N_12429);
nor U15774 (N_15774,N_12296,N_12166);
and U15775 (N_15775,N_12206,N_13878);
and U15776 (N_15776,N_14930,N_10582);
nor U15777 (N_15777,N_11654,N_10448);
nand U15778 (N_15778,N_14982,N_12369);
nor U15779 (N_15779,N_13220,N_13764);
or U15780 (N_15780,N_10687,N_11915);
and U15781 (N_15781,N_10403,N_14099);
nor U15782 (N_15782,N_11818,N_11323);
and U15783 (N_15783,N_10307,N_12976);
nand U15784 (N_15784,N_14223,N_14162);
and U15785 (N_15785,N_14101,N_13543);
and U15786 (N_15786,N_14065,N_14642);
or U15787 (N_15787,N_10884,N_13453);
or U15788 (N_15788,N_10810,N_12911);
and U15789 (N_15789,N_12560,N_12386);
or U15790 (N_15790,N_14067,N_13936);
nand U15791 (N_15791,N_12727,N_11962);
or U15792 (N_15792,N_14842,N_11310);
nor U15793 (N_15793,N_10396,N_11205);
and U15794 (N_15794,N_13052,N_12745);
nand U15795 (N_15795,N_14579,N_11773);
nor U15796 (N_15796,N_13795,N_14158);
nand U15797 (N_15797,N_12537,N_14839);
nor U15798 (N_15798,N_14201,N_10625);
nor U15799 (N_15799,N_14074,N_11793);
nand U15800 (N_15800,N_11891,N_13397);
or U15801 (N_15801,N_11116,N_14619);
nor U15802 (N_15802,N_10721,N_10494);
nor U15803 (N_15803,N_12022,N_10918);
nand U15804 (N_15804,N_10938,N_14233);
and U15805 (N_15805,N_12987,N_13938);
nand U15806 (N_15806,N_10132,N_13467);
and U15807 (N_15807,N_13952,N_14560);
and U15808 (N_15808,N_14261,N_12867);
nor U15809 (N_15809,N_12101,N_14572);
nand U15810 (N_15810,N_12658,N_13202);
nor U15811 (N_15811,N_14860,N_12430);
nor U15812 (N_15812,N_11778,N_10734);
or U15813 (N_15813,N_11107,N_12863);
and U15814 (N_15814,N_12488,N_11780);
nand U15815 (N_15815,N_12035,N_13387);
nand U15816 (N_15816,N_14519,N_11239);
and U15817 (N_15817,N_12977,N_12713);
and U15818 (N_15818,N_13682,N_14310);
nor U15819 (N_15819,N_12543,N_11947);
or U15820 (N_15820,N_14262,N_13166);
and U15821 (N_15821,N_14829,N_11361);
nand U15822 (N_15822,N_13260,N_13236);
nor U15823 (N_15823,N_10771,N_11384);
or U15824 (N_15824,N_11446,N_12776);
and U15825 (N_15825,N_12139,N_10211);
nand U15826 (N_15826,N_11969,N_10852);
or U15827 (N_15827,N_10689,N_12295);
and U15828 (N_15828,N_11506,N_12693);
and U15829 (N_15829,N_12041,N_14157);
xor U15830 (N_15830,N_14919,N_12371);
and U15831 (N_15831,N_14060,N_13038);
xnor U15832 (N_15832,N_10589,N_12092);
and U15833 (N_15833,N_14289,N_11733);
xnor U15834 (N_15834,N_14140,N_11671);
nand U15835 (N_15835,N_11750,N_11799);
nand U15836 (N_15836,N_10783,N_14200);
and U15837 (N_15837,N_14003,N_13805);
and U15838 (N_15838,N_14929,N_13894);
nor U15839 (N_15839,N_12285,N_14765);
and U15840 (N_15840,N_13388,N_13975);
and U15841 (N_15841,N_13827,N_14514);
or U15842 (N_15842,N_11075,N_12675);
or U15843 (N_15843,N_10521,N_11998);
nand U15844 (N_15844,N_12065,N_13902);
nor U15845 (N_15845,N_11928,N_10975);
xor U15846 (N_15846,N_14286,N_14905);
or U15847 (N_15847,N_11052,N_12998);
nor U15848 (N_15848,N_12256,N_11512);
and U15849 (N_15849,N_14191,N_12834);
nand U15850 (N_15850,N_10046,N_14721);
nor U15851 (N_15851,N_11726,N_12330);
nor U15852 (N_15852,N_11217,N_10039);
nor U15853 (N_15853,N_13086,N_13518);
nor U15854 (N_15854,N_14475,N_10390);
xor U15855 (N_15855,N_11914,N_14901);
nor U15856 (N_15856,N_13675,N_12259);
nor U15857 (N_15857,N_13129,N_10769);
or U15858 (N_15858,N_11376,N_10004);
nand U15859 (N_15859,N_13627,N_12289);
nand U15860 (N_15860,N_14994,N_11922);
or U15861 (N_15861,N_10702,N_12840);
nand U15862 (N_15862,N_10955,N_10885);
nor U15863 (N_15863,N_14116,N_13111);
and U15864 (N_15864,N_14629,N_10839);
or U15865 (N_15865,N_13568,N_11106);
xor U15866 (N_15866,N_14690,N_11146);
or U15867 (N_15867,N_12968,N_12334);
and U15868 (N_15868,N_12226,N_10663);
or U15869 (N_15869,N_14232,N_10613);
or U15870 (N_15870,N_10675,N_13800);
nor U15871 (N_15871,N_10347,N_11372);
or U15872 (N_15872,N_13901,N_11496);
and U15873 (N_15873,N_11354,N_12345);
xor U15874 (N_15874,N_10082,N_12339);
and U15875 (N_15875,N_14775,N_10557);
nor U15876 (N_15876,N_14090,N_10145);
or U15877 (N_15877,N_14841,N_12160);
nor U15878 (N_15878,N_12282,N_14528);
xnor U15879 (N_15879,N_10294,N_13900);
nor U15880 (N_15880,N_10826,N_13608);
and U15881 (N_15881,N_13640,N_11803);
or U15882 (N_15882,N_12098,N_11157);
nor U15883 (N_15883,N_11329,N_13715);
and U15884 (N_15884,N_10817,N_14399);
nor U15885 (N_15885,N_14788,N_14504);
and U15886 (N_15886,N_11713,N_11062);
nand U15887 (N_15887,N_14030,N_12415);
or U15888 (N_15888,N_13669,N_11470);
nand U15889 (N_15889,N_12197,N_11824);
nor U15890 (N_15890,N_12083,N_12984);
nor U15891 (N_15891,N_12004,N_10946);
nand U15892 (N_15892,N_14302,N_12164);
and U15893 (N_15893,N_14903,N_12148);
and U15894 (N_15894,N_12821,N_11826);
nand U15895 (N_15895,N_13378,N_11979);
and U15896 (N_15896,N_10800,N_14354);
nor U15897 (N_15897,N_12134,N_10270);
xor U15898 (N_15898,N_14676,N_12520);
xnor U15899 (N_15899,N_14877,N_14202);
and U15900 (N_15900,N_12153,N_12225);
or U15901 (N_15901,N_13977,N_11460);
and U15902 (N_15902,N_10161,N_10217);
nand U15903 (N_15903,N_13249,N_11327);
and U15904 (N_15904,N_10272,N_14939);
nand U15905 (N_15905,N_12513,N_11624);
or U15906 (N_15906,N_11356,N_13541);
or U15907 (N_15907,N_10209,N_14149);
nand U15908 (N_15908,N_14462,N_13230);
or U15909 (N_15909,N_13575,N_11455);
nor U15910 (N_15910,N_10634,N_10430);
and U15911 (N_15911,N_11290,N_12737);
nor U15912 (N_15912,N_12644,N_12514);
or U15913 (N_15913,N_11982,N_12191);
or U15914 (N_15914,N_12397,N_12996);
xnor U15915 (N_15915,N_10227,N_10225);
nand U15916 (N_15916,N_14457,N_13891);
nand U15917 (N_15917,N_12284,N_11102);
and U15918 (N_15918,N_13219,N_12169);
nand U15919 (N_15919,N_13618,N_14602);
nand U15920 (N_15920,N_10830,N_10824);
nand U15921 (N_15921,N_14503,N_14050);
and U15922 (N_15922,N_12764,N_10786);
nand U15923 (N_15923,N_11630,N_14608);
and U15924 (N_15924,N_11461,N_13287);
nor U15925 (N_15925,N_10086,N_13172);
nand U15926 (N_15926,N_13763,N_11729);
nor U15927 (N_15927,N_11260,N_14978);
and U15928 (N_15928,N_14141,N_13590);
nor U15929 (N_15929,N_11504,N_10989);
or U15930 (N_15930,N_12581,N_11214);
nand U15931 (N_15931,N_13837,N_14792);
nor U15932 (N_15932,N_10306,N_14640);
nor U15933 (N_15933,N_14426,N_13101);
and U15934 (N_15934,N_11908,N_10169);
or U15935 (N_15935,N_13234,N_12568);
or U15936 (N_15936,N_10296,N_10963);
nand U15937 (N_15937,N_13059,N_11264);
nor U15938 (N_15938,N_13250,N_12072);
or U15939 (N_15939,N_14264,N_13706);
nand U15940 (N_15940,N_12657,N_13182);
nand U15941 (N_15941,N_11734,N_12104);
nand U15942 (N_15942,N_10742,N_13216);
or U15943 (N_15943,N_10271,N_11893);
nor U15944 (N_15944,N_14716,N_13095);
nand U15945 (N_15945,N_13747,N_10378);
or U15946 (N_15946,N_12556,N_10005);
nor U15947 (N_15947,N_10936,N_11247);
nand U15948 (N_15948,N_13783,N_14858);
or U15949 (N_15949,N_13072,N_14244);
and U15950 (N_15950,N_13273,N_13930);
nand U15951 (N_15951,N_11478,N_13688);
nand U15952 (N_15952,N_12007,N_14520);
and U15953 (N_15953,N_11871,N_12927);
xnor U15954 (N_15954,N_13010,N_13863);
nand U15955 (N_15955,N_12331,N_10279);
nand U15956 (N_15956,N_14510,N_13087);
nand U15957 (N_15957,N_10532,N_12962);
nor U15958 (N_15958,N_14070,N_11129);
nand U15959 (N_15959,N_11447,N_11165);
and U15960 (N_15960,N_10094,N_13138);
and U15961 (N_15961,N_12554,N_13586);
or U15962 (N_15962,N_11035,N_11995);
and U15963 (N_15963,N_10120,N_10422);
or U15964 (N_15964,N_10796,N_13865);
nand U15965 (N_15965,N_14827,N_13344);
nand U15966 (N_15966,N_13168,N_12832);
nor U15967 (N_15967,N_13697,N_14219);
and U15968 (N_15968,N_12109,N_14024);
nand U15969 (N_15969,N_11574,N_10367);
nand U15970 (N_15970,N_11835,N_10208);
nand U15971 (N_15971,N_11718,N_10570);
and U15972 (N_15972,N_14361,N_14380);
and U15973 (N_15973,N_10020,N_10445);
or U15974 (N_15974,N_12828,N_11851);
xor U15975 (N_15975,N_11432,N_14296);
nand U15976 (N_15976,N_10985,N_11786);
nand U15977 (N_15977,N_13143,N_11349);
or U15978 (N_15978,N_11712,N_12161);
nand U15979 (N_15979,N_12793,N_11863);
xor U15980 (N_15980,N_10264,N_12668);
nand U15981 (N_15981,N_12257,N_11800);
and U15982 (N_15982,N_13836,N_14207);
and U15983 (N_15983,N_10098,N_13761);
or U15984 (N_15984,N_11695,N_11089);
nor U15985 (N_15985,N_13709,N_14324);
nand U15986 (N_15986,N_14134,N_14845);
nand U15987 (N_15987,N_10804,N_14702);
nor U15988 (N_15988,N_10050,N_10939);
nand U15989 (N_15989,N_14896,N_13696);
xor U15990 (N_15990,N_11791,N_13982);
nor U15991 (N_15991,N_10944,N_13360);
nor U15992 (N_15992,N_12817,N_13060);
nor U15993 (N_15993,N_13311,N_11554);
or U15994 (N_15994,N_14107,N_12944);
and U15995 (N_15995,N_12686,N_12733);
or U15996 (N_15996,N_10924,N_13639);
or U15997 (N_15997,N_13146,N_14639);
or U15998 (N_15998,N_14059,N_14785);
or U15999 (N_15999,N_10484,N_10164);
or U16000 (N_16000,N_13299,N_12954);
nand U16001 (N_16001,N_12087,N_14371);
and U16002 (N_16002,N_11105,N_12055);
nor U16003 (N_16003,N_12263,N_10840);
nor U16004 (N_16004,N_14588,N_14813);
nor U16005 (N_16005,N_14774,N_10757);
or U16006 (N_16006,N_14280,N_12855);
nand U16007 (N_16007,N_14571,N_10348);
nand U16008 (N_16008,N_12881,N_13325);
nand U16009 (N_16009,N_11375,N_11854);
and U16010 (N_16010,N_10000,N_10281);
nand U16011 (N_16011,N_13948,N_12907);
nor U16012 (N_16012,N_13896,N_11785);
or U16013 (N_16013,N_13520,N_10075);
and U16014 (N_16014,N_12294,N_12642);
nand U16015 (N_16015,N_12058,N_13828);
nor U16016 (N_16016,N_11865,N_14414);
or U16017 (N_16017,N_13662,N_14968);
nand U16018 (N_16018,N_10909,N_10040);
or U16019 (N_16019,N_13149,N_11683);
or U16020 (N_16020,N_11249,N_12919);
or U16021 (N_16021,N_13854,N_14488);
and U16022 (N_16022,N_11200,N_14355);
or U16023 (N_16023,N_13379,N_13235);
nor U16024 (N_16024,N_13459,N_11684);
xor U16025 (N_16025,N_13286,N_11145);
nor U16026 (N_16026,N_11294,N_13536);
and U16027 (N_16027,N_12786,N_10971);
nor U16028 (N_16028,N_10222,N_12629);
and U16029 (N_16029,N_12586,N_11658);
nand U16030 (N_16030,N_10081,N_14651);
and U16031 (N_16031,N_13700,N_14876);
and U16032 (N_16032,N_14934,N_14867);
nand U16033 (N_16033,N_11846,N_13113);
nand U16034 (N_16034,N_11359,N_11764);
nand U16035 (N_16035,N_10701,N_11272);
nor U16036 (N_16036,N_10512,N_12757);
or U16037 (N_16037,N_11777,N_12490);
or U16038 (N_16038,N_11187,N_11238);
nand U16039 (N_16039,N_11253,N_14438);
nand U16040 (N_16040,N_13003,N_14958);
or U16041 (N_16041,N_11215,N_10105);
or U16042 (N_16042,N_11385,N_10121);
nor U16043 (N_16043,N_10514,N_10720);
nand U16044 (N_16044,N_14386,N_13691);
nor U16045 (N_16045,N_11985,N_14287);
and U16046 (N_16046,N_11289,N_11188);
nand U16047 (N_16047,N_11336,N_13210);
or U16048 (N_16048,N_12694,N_14864);
and U16049 (N_16049,N_14348,N_11830);
and U16050 (N_16050,N_13390,N_12125);
nand U16051 (N_16051,N_12012,N_11179);
and U16052 (N_16052,N_11591,N_11725);
nand U16053 (N_16053,N_10436,N_14446);
and U16054 (N_16054,N_11383,N_11091);
nor U16055 (N_16055,N_14124,N_11847);
and U16056 (N_16056,N_13076,N_12692);
nor U16057 (N_16057,N_14000,N_13443);
nor U16058 (N_16058,N_12632,N_11006);
or U16059 (N_16059,N_12499,N_13737);
nand U16060 (N_16060,N_12948,N_10928);
and U16061 (N_16061,N_10616,N_12443);
and U16062 (N_16062,N_10717,N_13864);
nand U16063 (N_16063,N_10326,N_10158);
nor U16064 (N_16064,N_13475,N_14544);
nor U16065 (N_16065,N_14518,N_11983);
and U16066 (N_16066,N_14309,N_13428);
nor U16067 (N_16067,N_11237,N_10160);
xor U16068 (N_16068,N_14187,N_10419);
and U16069 (N_16069,N_11659,N_13162);
or U16070 (N_16070,N_12383,N_11939);
nand U16071 (N_16071,N_11297,N_12486);
nor U16072 (N_16072,N_13342,N_13811);
xor U16073 (N_16073,N_13317,N_11277);
and U16074 (N_16074,N_13671,N_12617);
or U16075 (N_16075,N_13912,N_14317);
or U16076 (N_16076,N_14875,N_14088);
nand U16077 (N_16077,N_14757,N_10991);
nand U16078 (N_16078,N_10051,N_11023);
or U16079 (N_16079,N_11117,N_14960);
and U16080 (N_16080,N_12472,N_10499);
or U16081 (N_16081,N_12857,N_13259);
and U16082 (N_16082,N_13039,N_10196);
or U16083 (N_16083,N_10288,N_10245);
and U16084 (N_16084,N_10201,N_13472);
and U16085 (N_16085,N_13380,N_14288);
xor U16086 (N_16086,N_11223,N_13558);
and U16087 (N_16087,N_10386,N_13924);
and U16088 (N_16088,N_11653,N_11344);
and U16089 (N_16089,N_12901,N_12349);
and U16090 (N_16090,N_12237,N_12483);
nor U16091 (N_16091,N_14278,N_10333);
or U16092 (N_16092,N_14383,N_12703);
or U16093 (N_16093,N_14601,N_10183);
nand U16094 (N_16094,N_13075,N_14773);
or U16095 (N_16095,N_12601,N_11772);
and U16096 (N_16096,N_12135,N_11679);
nor U16097 (N_16097,N_14384,N_13159);
nand U16098 (N_16098,N_13150,N_13290);
nor U16099 (N_16099,N_12521,N_13825);
and U16100 (N_16100,N_14305,N_11907);
nor U16101 (N_16101,N_10568,N_12389);
or U16102 (N_16102,N_12227,N_14587);
nor U16103 (N_16103,N_13322,N_11050);
or U16104 (N_16104,N_14473,N_14055);
nand U16105 (N_16105,N_13529,N_10779);
nand U16106 (N_16106,N_14345,N_12699);
or U16107 (N_16107,N_13215,N_12856);
nor U16108 (N_16108,N_10544,N_12528);
nor U16109 (N_16109,N_11941,N_14777);
nand U16110 (N_16110,N_11583,N_10748);
nand U16111 (N_16111,N_11548,N_12103);
nor U16112 (N_16112,N_10360,N_14469);
nor U16113 (N_16113,N_12982,N_10969);
or U16114 (N_16114,N_12509,N_14670);
and U16115 (N_16115,N_13133,N_11924);
and U16116 (N_16116,N_14753,N_14411);
nand U16117 (N_16117,N_10072,N_11868);
and U16118 (N_16118,N_13238,N_10253);
or U16119 (N_16119,N_10152,N_10215);
or U16120 (N_16120,N_12039,N_11054);
nor U16121 (N_16121,N_13909,N_13352);
or U16122 (N_16122,N_13062,N_12525);
xor U16123 (N_16123,N_13016,N_11000);
nor U16124 (N_16124,N_11255,N_13027);
nand U16125 (N_16125,N_13243,N_11270);
or U16126 (N_16126,N_13701,N_14523);
xnor U16127 (N_16127,N_11758,N_12333);
nor U16128 (N_16128,N_10737,N_11417);
nand U16129 (N_16129,N_14382,N_14225);
or U16130 (N_16130,N_11689,N_11407);
or U16131 (N_16131,N_14293,N_13813);
nand U16132 (N_16132,N_12057,N_14072);
nand U16133 (N_16133,N_12966,N_12303);
and U16134 (N_16134,N_12364,N_10667);
xor U16135 (N_16135,N_14590,N_10903);
or U16136 (N_16136,N_14335,N_13710);
or U16137 (N_16137,N_11507,N_11124);
nor U16138 (N_16138,N_10248,N_12384);
nor U16139 (N_16139,N_10738,N_14334);
and U16140 (N_16140,N_14043,N_11010);
and U16141 (N_16141,N_13947,N_11025);
and U16142 (N_16142,N_10536,N_13594);
nor U16143 (N_16143,N_13267,N_11080);
or U16144 (N_16144,N_12969,N_14304);
or U16145 (N_16145,N_12916,N_13118);
and U16146 (N_16146,N_13913,N_12344);
or U16147 (N_16147,N_13797,N_14256);
or U16148 (N_16148,N_11196,N_13121);
and U16149 (N_16149,N_11234,N_11940);
or U16150 (N_16150,N_10310,N_12549);
nor U16151 (N_16151,N_14333,N_14495);
and U16152 (N_16152,N_11749,N_12761);
nor U16153 (N_16153,N_10175,N_11011);
nor U16154 (N_16154,N_13415,N_13152);
nand U16155 (N_16155,N_14805,N_11618);
or U16156 (N_16156,N_13186,N_10685);
or U16157 (N_16157,N_11155,N_10033);
and U16158 (N_16158,N_13622,N_11899);
nand U16159 (N_16159,N_10026,N_10412);
xnor U16160 (N_16160,N_13677,N_11008);
or U16161 (N_16161,N_10805,N_13694);
nor U16162 (N_16162,N_13572,N_14385);
nor U16163 (N_16163,N_11319,N_13626);
nor U16164 (N_16164,N_10282,N_14271);
nor U16165 (N_16165,N_12229,N_12214);
and U16166 (N_16166,N_13989,N_11071);
or U16167 (N_16167,N_10014,N_10855);
or U16168 (N_16168,N_14977,N_13742);
and U16169 (N_16169,N_11242,N_10030);
nor U16170 (N_16170,N_11534,N_11401);
or U16171 (N_16171,N_11434,N_11048);
or U16172 (N_16172,N_14089,N_13389);
or U16173 (N_16173,N_12112,N_10768);
nand U16174 (N_16174,N_13093,N_12932);
or U16175 (N_16175,N_10560,N_14594);
nor U16176 (N_16176,N_14444,N_14086);
and U16177 (N_16177,N_14511,N_11440);
and U16178 (N_16178,N_10115,N_14066);
nor U16179 (N_16179,N_11377,N_10340);
nor U16180 (N_16180,N_11787,N_14480);
or U16181 (N_16181,N_14779,N_10899);
or U16182 (N_16182,N_14179,N_14592);
xor U16183 (N_16183,N_13599,N_12874);
or U16184 (N_16184,N_13611,N_10607);
nand U16185 (N_16185,N_14249,N_10042);
and U16186 (N_16186,N_13579,N_14203);
or U16187 (N_16187,N_12107,N_12913);
nor U16188 (N_16188,N_14894,N_12995);
nand U16189 (N_16189,N_14284,N_10605);
or U16190 (N_16190,N_12013,N_13363);
or U16191 (N_16191,N_14880,N_10508);
nand U16192 (N_16192,N_13538,N_12312);
and U16193 (N_16193,N_11328,N_13136);
nand U16194 (N_16194,N_14300,N_10954);
or U16195 (N_16195,N_14236,N_12474);
or U16196 (N_16196,N_10321,N_13140);
nand U16197 (N_16197,N_14908,N_11919);
nor U16198 (N_16198,N_13232,N_12479);
nor U16199 (N_16199,N_10236,N_13593);
or U16200 (N_16200,N_10632,N_11759);
nand U16201 (N_16201,N_14553,N_11466);
nand U16202 (N_16202,N_14073,N_14145);
or U16203 (N_16203,N_11622,N_13491);
nand U16204 (N_16204,N_14809,N_12484);
nor U16205 (N_16205,N_13269,N_13911);
and U16206 (N_16206,N_12879,N_12446);
nor U16207 (N_16207,N_10949,N_13408);
nor U16208 (N_16208,N_11331,N_12853);
or U16209 (N_16209,N_10335,N_10463);
xor U16210 (N_16210,N_13021,N_11692);
xor U16211 (N_16211,N_13630,N_13686);
and U16212 (N_16212,N_13768,N_14595);
nor U16213 (N_16213,N_12099,N_12049);
or U16214 (N_16214,N_13487,N_14082);
nor U16215 (N_16215,N_12636,N_10637);
nand U16216 (N_16216,N_12159,N_14984);
nand U16217 (N_16217,N_12044,N_11840);
nand U16218 (N_16218,N_14206,N_14136);
or U16219 (N_16219,N_14265,N_11889);
nand U16220 (N_16220,N_12678,N_13985);
and U16221 (N_16221,N_10994,N_11271);
nand U16222 (N_16222,N_14417,N_14993);
nor U16223 (N_16223,N_14168,N_10866);
nand U16224 (N_16224,N_11885,N_10128);
nand U16225 (N_16225,N_12780,N_13254);
or U16226 (N_16226,N_12010,N_11104);
nand U16227 (N_16227,N_11802,N_11655);
and U16228 (N_16228,N_14613,N_12350);
nand U16229 (N_16229,N_11073,N_14883);
or U16230 (N_16230,N_13450,N_11454);
and U16231 (N_16231,N_10230,N_11330);
nor U16232 (N_16232,N_14754,N_11657);
and U16233 (N_16233,N_10892,N_10027);
or U16234 (N_16234,N_11218,N_13548);
nand U16235 (N_16235,N_13231,N_11974);
nor U16236 (N_16236,N_12189,N_11364);
and U16237 (N_16237,N_13343,N_10472);
nand U16238 (N_16238,N_13326,N_11748);
nor U16239 (N_16239,N_12414,N_11476);
and U16240 (N_16240,N_11127,N_12274);
and U16241 (N_16241,N_14152,N_14326);
and U16242 (N_16242,N_14540,N_14505);
and U16243 (N_16243,N_11613,N_13142);
nor U16244 (N_16244,N_13449,N_12955);
nor U16245 (N_16245,N_14253,N_14863);
nor U16246 (N_16246,N_12611,N_10413);
nand U16247 (N_16247,N_12628,N_14755);
and U16248 (N_16248,N_14577,N_10883);
nand U16249 (N_16249,N_10262,N_12762);
nand U16250 (N_16250,N_13597,N_10224);
or U16251 (N_16251,N_11267,N_10019);
and U16252 (N_16252,N_10788,N_14295);
nor U16253 (N_16253,N_13237,N_12517);
nor U16254 (N_16254,N_12590,N_14299);
nor U16255 (N_16255,N_13509,N_11020);
nand U16256 (N_16256,N_12772,N_13471);
and U16257 (N_16257,N_11586,N_11084);
nand U16258 (N_16258,N_13498,N_12871);
nor U16259 (N_16259,N_13291,N_10068);
nand U16260 (N_16260,N_13106,N_14893);
and U16261 (N_16261,N_11430,N_12950);
and U16262 (N_16262,N_14554,N_12595);
nor U16263 (N_16263,N_10061,N_13354);
and U16264 (N_16264,N_10334,N_14097);
nor U16265 (N_16265,N_11170,N_13437);
and U16266 (N_16266,N_14900,N_13289);
or U16267 (N_16267,N_12034,N_14857);
nor U16268 (N_16268,N_11281,N_13659);
or U16269 (N_16269,N_13044,N_14555);
and U16270 (N_16270,N_11456,N_12994);
or U16271 (N_16271,N_10555,N_14393);
nor U16272 (N_16272,N_11216,N_14212);
nor U16273 (N_16273,N_11966,N_14799);
or U16274 (N_16274,N_13784,N_14238);
nand U16275 (N_16275,N_10709,N_13277);
nand U16276 (N_16276,N_14272,N_14976);
or U16277 (N_16277,N_13766,N_11014);
nor U16278 (N_16278,N_10567,N_12120);
xor U16279 (N_16279,N_11321,N_13399);
nor U16280 (N_16280,N_13218,N_11299);
nor U16281 (N_16281,N_11641,N_10762);
and U16282 (N_16282,N_13940,N_12773);
or U16283 (N_16283,N_13007,N_11427);
xor U16284 (N_16284,N_13693,N_11282);
nand U16285 (N_16285,N_12152,N_13746);
and U16286 (N_16286,N_12026,N_14843);
nand U16287 (N_16287,N_10633,N_13461);
nor U16288 (N_16288,N_13990,N_13650);
or U16289 (N_16289,N_12858,N_10665);
xor U16290 (N_16290,N_13807,N_13228);
nor U16291 (N_16291,N_10857,N_10338);
nor U16292 (N_16292,N_10851,N_10600);
or U16293 (N_16293,N_12200,N_12800);
nand U16294 (N_16294,N_14147,N_10298);
nand U16295 (N_16295,N_12538,N_10754);
or U16296 (N_16296,N_14657,N_12802);
nand U16297 (N_16297,N_10761,N_11426);
nand U16298 (N_16298,N_12961,N_12826);
nand U16299 (N_16299,N_11431,N_11886);
nor U16300 (N_16300,N_10628,N_10462);
and U16301 (N_16301,N_10699,N_11876);
and U16302 (N_16302,N_11380,N_12036);
or U16303 (N_16303,N_10141,N_14865);
nor U16304 (N_16304,N_14665,N_14370);
nand U16305 (N_16305,N_13929,N_12940);
nor U16306 (N_16306,N_10022,N_11719);
nor U16307 (N_16307,N_14748,N_14586);
and U16308 (N_16308,N_11400,N_12505);
xnor U16309 (N_16309,N_12249,N_12467);
nor U16310 (N_16310,N_12110,N_10968);
and U16311 (N_16311,N_14193,N_13791);
nor U16312 (N_16312,N_14695,N_10137);
nor U16313 (N_16313,N_14109,N_12433);
xnor U16314 (N_16314,N_14128,N_10733);
nor U16315 (N_16315,N_12476,N_12613);
and U16316 (N_16316,N_14911,N_14084);
nor U16317 (N_16317,N_13623,N_11527);
or U16318 (N_16318,N_11015,N_11123);
and U16319 (N_16319,N_13297,N_10221);
nor U16320 (N_16320,N_11307,N_14561);
nand U16321 (N_16321,N_11751,N_13967);
or U16322 (N_16322,N_13573,N_12723);
nor U16323 (N_16323,N_10553,N_10452);
nand U16324 (N_16324,N_10006,N_12957);
and U16325 (N_16325,N_13552,N_10154);
or U16326 (N_16326,N_10179,N_10770);
xor U16327 (N_16327,N_14487,N_14408);
or U16328 (N_16328,N_13582,N_10251);
nor U16329 (N_16329,N_11024,N_11002);
or U16330 (N_16330,N_12577,N_12188);
and U16331 (N_16331,N_11867,N_10099);
and U16332 (N_16332,N_14464,N_11643);
or U16333 (N_16333,N_14453,N_11108);
xor U16334 (N_16334,N_14653,N_14840);
xnor U16335 (N_16335,N_13576,N_10238);
or U16336 (N_16336,N_11809,N_12837);
nand U16337 (N_16337,N_10747,N_14636);
or U16338 (N_16338,N_14729,N_13312);
and U16339 (N_16339,N_14666,N_12541);
nor U16340 (N_16340,N_14173,N_10016);
and U16341 (N_16341,N_12293,N_13767);
nand U16342 (N_16342,N_14924,N_12145);
or U16343 (N_16343,N_11192,N_13058);
and U16344 (N_16344,N_11485,N_11499);
nand U16345 (N_16345,N_13739,N_10405);
and U16346 (N_16346,N_11697,N_13899);
nor U16347 (N_16347,N_10542,N_14969);
and U16348 (N_16348,N_13189,N_14822);
or U16349 (N_16349,N_11060,N_12903);
or U16350 (N_16350,N_13873,N_10443);
and U16351 (N_16351,N_13931,N_11444);
nand U16352 (N_16352,N_13723,N_10186);
nand U16353 (N_16353,N_13444,N_13460);
or U16354 (N_16354,N_14075,N_14125);
and U16355 (N_16355,N_14578,N_11483);
and U16356 (N_16356,N_14521,N_14545);
or U16357 (N_16357,N_13199,N_11452);
or U16358 (N_16358,N_13144,N_10872);
nand U16359 (N_16359,N_10429,N_11395);
and U16360 (N_16360,N_10631,N_11302);
nor U16361 (N_16361,N_14163,N_12937);
nand U16362 (N_16362,N_12697,N_13278);
nand U16363 (N_16363,N_14485,N_11905);
nand U16364 (N_16364,N_11705,N_13211);
and U16365 (N_16365,N_11109,N_13079);
and U16366 (N_16366,N_14196,N_10170);
nand U16367 (N_16367,N_11537,N_14907);
or U16368 (N_16368,N_12271,N_10877);
and U16369 (N_16369,N_14667,N_13988);
or U16370 (N_16370,N_14153,N_10118);
or U16371 (N_16371,N_10540,N_13078);
nand U16372 (N_16372,N_14257,N_12064);
or U16373 (N_16373,N_13431,N_12888);
nand U16374 (N_16374,N_13067,N_10952);
and U16375 (N_16375,N_13951,N_11776);
and U16376 (N_16376,N_11814,N_13158);
nand U16377 (N_16377,N_12583,N_12393);
nor U16378 (N_16378,N_11788,N_12122);
xnor U16379 (N_16379,N_13481,N_12340);
nor U16380 (N_16380,N_14425,N_10459);
nor U16381 (N_16381,N_11148,N_11727);
or U16382 (N_16382,N_11137,N_13465);
and U16383 (N_16383,N_10621,N_12909);
and U16384 (N_16384,N_14638,N_12001);
and U16385 (N_16385,N_14684,N_13280);
and U16386 (N_16386,N_11304,N_12481);
and U16387 (N_16387,N_14918,N_12212);
xor U16388 (N_16388,N_11110,N_10523);
and U16389 (N_16389,N_11910,N_12902);
or U16390 (N_16390,N_11714,N_10106);
or U16391 (N_16391,N_13732,N_12174);
nor U16392 (N_16392,N_10671,N_13134);
and U16393 (N_16393,N_10674,N_10136);
or U16394 (N_16394,N_14909,N_12965);
nor U16395 (N_16395,N_10807,N_12054);
and U16396 (N_16396,N_13657,N_10242);
nand U16397 (N_16397,N_13125,N_10780);
nand U16398 (N_16398,N_10541,N_14654);
nor U16399 (N_16399,N_14663,N_12432);
xnor U16400 (N_16400,N_11337,N_11254);
and U16401 (N_16401,N_14706,N_12498);
nand U16402 (N_16402,N_11182,N_11122);
nor U16403 (N_16403,N_13446,N_13422);
and U16404 (N_16404,N_13602,N_11082);
and U16405 (N_16405,N_13609,N_10879);
or U16406 (N_16406,N_12653,N_14862);
or U16407 (N_16407,N_11843,N_11901);
nand U16408 (N_16408,N_14252,N_11822);
and U16409 (N_16409,N_11959,N_10606);
nand U16410 (N_16410,N_11190,N_11590);
nand U16411 (N_16411,N_11837,N_13321);
and U16412 (N_16412,N_14209,N_12126);
or U16413 (N_16413,N_13776,N_10656);
nor U16414 (N_16414,N_12672,N_13174);
or U16415 (N_16415,N_13826,N_11681);
and U16416 (N_16416,N_12747,N_11665);
xnor U16417 (N_16417,N_10718,N_11436);
and U16418 (N_16418,N_11703,N_12132);
nand U16419 (N_16419,N_14169,N_12591);
and U16420 (N_16420,N_11250,N_14301);
nand U16421 (N_16421,N_10048,N_10434);
or U16422 (N_16422,N_13248,N_11018);
nor U16423 (N_16423,N_13906,N_12963);
nor U16424 (N_16424,N_10820,N_13525);
or U16425 (N_16425,N_12945,N_13314);
and U16426 (N_16426,N_11374,N_13381);
and U16427 (N_16427,N_10373,N_13394);
or U16428 (N_16428,N_11406,N_12716);
nand U16429 (N_16429,N_12767,N_11278);
nand U16430 (N_16430,N_13524,N_14688);
xnor U16431 (N_16431,N_13810,N_13335);
and U16432 (N_16432,N_11811,N_10404);
nor U16433 (N_16433,N_13004,N_13698);
nor U16434 (N_16434,N_13829,N_14745);
nand U16435 (N_16435,N_10828,N_12971);
and U16436 (N_16436,N_14053,N_12466);
or U16437 (N_16437,N_13407,N_12440);
nand U16438 (N_16438,N_12268,N_12193);
and U16439 (N_16439,N_13972,N_12865);
xor U16440 (N_16440,N_10691,N_12492);
nor U16441 (N_16441,N_13598,N_10569);
or U16442 (N_16442,N_10379,N_10678);
or U16443 (N_16443,N_13644,N_10888);
nand U16444 (N_16444,N_13084,N_13019);
or U16445 (N_16445,N_14802,N_12530);
nor U16446 (N_16446,N_11397,N_10962);
nor U16447 (N_16447,N_13654,N_11968);
and U16448 (N_16448,N_13853,N_13606);
nor U16449 (N_16449,N_14810,N_12512);
or U16450 (N_16450,N_14526,N_11381);
nor U16451 (N_16451,N_12388,N_11790);
nand U16452 (N_16452,N_14807,N_13247);
nand U16453 (N_16453,N_11858,N_11220);
xor U16454 (N_16454,N_12162,N_11607);
nand U16455 (N_16455,N_10654,N_11967);
nand U16456 (N_16456,N_14516,N_10394);
and U16457 (N_16457,N_12958,N_12272);
nor U16458 (N_16458,N_11767,N_13098);
or U16459 (N_16459,N_13816,N_12401);
nand U16460 (N_16460,N_13504,N_10364);
nor U16461 (N_16461,N_14989,N_13110);
or U16462 (N_16462,N_12736,N_11462);
and U16463 (N_16463,N_14508,N_11298);
nand U16464 (N_16464,N_12376,N_14210);
nand U16465 (N_16465,N_14801,N_12290);
or U16466 (N_16466,N_11445,N_10058);
xor U16467 (N_16467,N_11569,N_10870);
and U16468 (N_16468,N_12947,N_10111);
and U16469 (N_16469,N_12833,N_13991);
or U16470 (N_16470,N_11142,N_11222);
xor U16471 (N_16471,N_10291,N_14532);
nor U16472 (N_16472,N_11988,N_10882);
and U16473 (N_16473,N_13840,N_10795);
and U16474 (N_16474,N_11360,N_14294);
or U16475 (N_16475,N_11615,N_10477);
nor U16476 (N_16476,N_10353,N_10102);
and U16477 (N_16477,N_10491,N_14423);
or U16478 (N_16478,N_12728,N_12391);
or U16479 (N_16479,N_13903,N_14402);
or U16480 (N_16480,N_14103,N_14786);
nand U16481 (N_16481,N_12131,N_10915);
or U16482 (N_16482,N_10008,N_12445);
nand U16483 (N_16483,N_11861,N_11739);
nand U16484 (N_16484,N_14938,N_14879);
and U16485 (N_16485,N_14471,N_11596);
nand U16486 (N_16486,N_12179,N_14445);
or U16487 (N_16487,N_10697,N_13028);
nand U16488 (N_16488,N_12523,N_12610);
or U16489 (N_16489,N_14395,N_10661);
nand U16490 (N_16490,N_13758,N_11236);
or U16491 (N_16491,N_11486,N_12138);
or U16492 (N_16492,N_14759,N_10919);
nand U16493 (N_16493,N_14685,N_10947);
nand U16494 (N_16494,N_13486,N_13601);
nand U16495 (N_16495,N_12619,N_13812);
or U16496 (N_16496,N_10290,N_11690);
nand U16497 (N_16497,N_13073,N_12536);
nand U16498 (N_16498,N_12421,N_14811);
or U16499 (N_16499,N_14359,N_10447);
nand U16500 (N_16500,N_12886,N_13532);
and U16501 (N_16501,N_13950,N_12700);
or U16502 (N_16502,N_10446,N_12774);
nor U16503 (N_16503,N_14338,N_10686);
and U16504 (N_16504,N_10846,N_11419);
nor U16505 (N_16505,N_11030,N_13780);
or U16506 (N_16506,N_13029,N_11980);
nand U16507 (N_16507,N_12676,N_11946);
or U16508 (N_16508,N_10156,N_10552);
and U16509 (N_16509,N_12557,N_10690);
and U16510 (N_16510,N_12320,N_12452);
nor U16511 (N_16511,N_13521,N_13351);
nor U16512 (N_16512,N_12210,N_12258);
and U16513 (N_16513,N_12704,N_11677);
or U16514 (N_16514,N_14105,N_10549);
and U16515 (N_16515,N_11408,N_14955);
nor U16516 (N_16516,N_11292,N_14243);
or U16517 (N_16517,N_11161,N_13956);
or U16518 (N_16518,N_13927,N_10649);
nand U16519 (N_16519,N_11832,N_13882);
nor U16520 (N_16520,N_14250,N_13651);
or U16521 (N_16521,N_12419,N_13769);
nor U16522 (N_16522,N_13457,N_12814);
and U16523 (N_16523,N_10104,N_11369);
nor U16524 (N_16524,N_11171,N_13208);
xor U16525 (N_16525,N_13089,N_12100);
and U16526 (N_16526,N_11629,N_13944);
nor U16527 (N_16527,N_10031,N_10509);
or U16528 (N_16528,N_12300,N_11756);
and U16529 (N_16529,N_11553,N_13757);
nor U16530 (N_16530,N_10887,N_11115);
nand U16531 (N_16531,N_13224,N_12074);
nand U16532 (N_16532,N_13629,N_10502);
and U16533 (N_16533,N_10874,N_10309);
nand U16534 (N_16534,N_10254,N_12730);
and U16535 (N_16535,N_14419,N_12063);
or U16536 (N_16536,N_10148,N_13774);
nand U16537 (N_16537,N_10808,N_10729);
and U16538 (N_16538,N_12060,N_13405);
and U16539 (N_16539,N_10139,N_11845);
or U16540 (N_16540,N_11935,N_10377);
nand U16541 (N_16541,N_10976,N_13540);
or U16542 (N_16542,N_10527,N_12032);
nor U16543 (N_16543,N_10305,N_13844);
and U16544 (N_16544,N_14652,N_11459);
or U16545 (N_16545,N_12273,N_13755);
and U16546 (N_16546,N_12051,N_11087);
and U16547 (N_16547,N_10007,N_12495);
nor U16548 (N_16548,N_14435,N_13333);
nand U16549 (N_16549,N_14749,N_12204);
and U16550 (N_16550,N_10782,N_12952);
nand U16551 (N_16551,N_12096,N_10803);
and U16552 (N_16552,N_14175,N_13116);
nor U16553 (N_16553,N_13564,N_14895);
nor U16554 (N_16554,N_11810,N_13842);
nand U16555 (N_16555,N_14668,N_12559);
nand U16556 (N_16556,N_12224,N_11244);
and U16557 (N_16557,N_14583,N_12077);
and U16558 (N_16558,N_13661,N_12173);
or U16559 (N_16559,N_14183,N_14039);
nor U16560 (N_16560,N_14248,N_14673);
nor U16561 (N_16561,N_14549,N_12778);
or U16562 (N_16562,N_13187,N_11921);
and U16563 (N_16563,N_13037,N_11412);
and U16564 (N_16564,N_12302,N_13957);
or U16565 (N_16565,N_14620,N_14156);
nand U16566 (N_16566,N_11177,N_14967);
or U16567 (N_16567,N_12053,N_14964);
nand U16568 (N_16568,N_13591,N_11012);
nor U16569 (N_16569,N_12405,N_13533);
nor U16570 (N_16570,N_10346,N_12553);
nand U16571 (N_16571,N_11367,N_12614);
and U16572 (N_16572,N_14009,N_13958);
nor U16573 (N_16573,N_12236,N_14023);
nand U16574 (N_16574,N_10601,N_13017);
nor U16575 (N_16575,N_12015,N_13303);
or U16576 (N_16576,N_10604,N_11570);
nor U16577 (N_16577,N_12280,N_13786);
or U16578 (N_16578,N_14478,N_13403);
nor U16579 (N_16579,N_14068,N_10460);
nor U16580 (N_16580,N_14327,N_10397);
and U16581 (N_16581,N_14790,N_10833);
and U16582 (N_16582,N_11528,N_10679);
and U16583 (N_16583,N_12760,N_10162);
nand U16584 (N_16584,N_13566,N_13429);
nor U16585 (N_16585,N_14432,N_13494);
and U16586 (N_16586,N_10398,N_14987);
xor U16587 (N_16587,N_12794,N_12608);
or U16588 (N_16588,N_14953,N_14170);
and U16589 (N_16589,N_13288,N_11005);
or U16590 (N_16590,N_12574,N_11368);
and U16591 (N_16591,N_12753,N_11438);
or U16592 (N_16592,N_10593,N_10792);
and U16593 (N_16593,N_13729,N_12981);
nor U16594 (N_16594,N_10664,N_13386);
and U16595 (N_16595,N_12600,N_11978);
xor U16596 (N_16596,N_14723,N_13188);
nor U16597 (N_16597,N_10266,N_11128);
nor U16598 (N_16598,N_12677,N_12045);
or U16599 (N_16599,N_11632,N_14167);
or U16600 (N_16600,N_14835,N_13454);
or U16601 (N_16601,N_14017,N_12094);
nand U16602 (N_16602,N_14245,N_11952);
nand U16603 (N_16603,N_11971,N_10138);
xor U16604 (N_16604,N_14247,N_14004);
nand U16605 (N_16605,N_13806,N_14509);
nand U16606 (N_16606,N_11640,N_10715);
nor U16607 (N_16607,N_13935,N_10257);
nand U16608 (N_16608,N_10475,N_14367);
nor U16609 (N_16609,N_12335,N_11930);
nor U16610 (N_16610,N_14412,N_14712);
nor U16611 (N_16611,N_13664,N_13738);
and U16612 (N_16612,N_12518,N_11598);
nand U16613 (N_16613,N_12037,N_14217);
and U16614 (N_16614,N_14443,N_13203);
or U16615 (N_16615,N_13305,N_12093);
and U16616 (N_16616,N_10028,N_12009);
nand U16617 (N_16617,N_12529,N_13064);
nand U16618 (N_16618,N_11595,N_11194);
nand U16619 (N_16619,N_11451,N_14186);
nand U16620 (N_16620,N_13293,N_13255);
and U16621 (N_16621,N_11311,N_11162);
and U16622 (N_16622,N_10009,N_11699);
or U16623 (N_16623,N_10126,N_14607);
nand U16624 (N_16624,N_14551,N_14787);
and U16625 (N_16625,N_10898,N_12899);
nand U16626 (N_16626,N_13614,N_13849);
or U16627 (N_16627,N_12534,N_11549);
and U16628 (N_16628,N_12640,N_14427);
or U16629 (N_16629,N_11219,N_14032);
or U16630 (N_16630,N_13647,N_10147);
or U16631 (N_16631,N_10455,N_10743);
or U16632 (N_16632,N_10559,N_12275);
or U16633 (N_16633,N_12321,N_14682);
or U16634 (N_16634,N_10258,N_12493);
or U16635 (N_16635,N_13672,N_12234);
and U16636 (N_16636,N_14092,N_11662);
nor U16637 (N_16637,N_14621,N_12689);
and U16638 (N_16638,N_13862,N_14889);
nor U16639 (N_16639,N_10062,N_13549);
or U16640 (N_16640,N_11338,N_13733);
and U16641 (N_16641,N_14466,N_10468);
or U16642 (N_16642,N_10240,N_10561);
and U16643 (N_16643,N_10736,N_11870);
or U16644 (N_16644,N_10787,N_11864);
nor U16645 (N_16645,N_11286,N_13173);
and U16646 (N_16646,N_14719,N_12066);
nor U16647 (N_16647,N_10395,N_11923);
nand U16648 (N_16648,N_10937,N_11816);
nor U16649 (N_16649,N_14565,N_11064);
nor U16650 (N_16650,N_10327,N_13976);
nand U16651 (N_16651,N_14693,N_11031);
and U16652 (N_16652,N_10206,N_13978);
nor U16653 (N_16653,N_12319,N_14761);
nor U16654 (N_16654,N_10789,N_11158);
xnor U16655 (N_16655,N_10318,N_14323);
and U16656 (N_16656,N_14837,N_11118);
nor U16657 (N_16657,N_13434,N_13506);
and U16658 (N_16658,N_14627,N_12147);
nor U16659 (N_16659,N_10311,N_11672);
or U16660 (N_16660,N_14034,N_10794);
and U16661 (N_16661,N_10778,N_11505);
or U16662 (N_16662,N_12456,N_13171);
and U16663 (N_16663,N_12385,N_11423);
nor U16664 (N_16664,N_12635,N_14947);
nor U16665 (N_16665,N_12959,N_13373);
nand U16666 (N_16666,N_10550,N_12599);
or U16667 (N_16667,N_10652,N_12852);
nor U16668 (N_16668,N_14331,N_14564);
and U16669 (N_16669,N_12544,N_13722);
and U16670 (N_16670,N_14585,N_11513);
or U16671 (N_16671,N_10594,N_14780);
nand U16672 (N_16672,N_12382,N_12949);
or U16673 (N_16673,N_12552,N_12408);
or U16674 (N_16674,N_14077,N_11515);
or U16675 (N_16675,N_13295,N_11490);
or U16676 (N_16676,N_13923,N_14506);
and U16677 (N_16677,N_10592,N_11121);
nand U16678 (N_16678,N_11240,N_13217);
nor U16679 (N_16679,N_10252,N_12508);
or U16680 (N_16680,N_13245,N_10528);
and U16681 (N_16681,N_11611,N_14734);
or U16682 (N_16682,N_14216,N_12637);
or U16683 (N_16683,N_10056,N_14328);
nor U16684 (N_16684,N_12785,N_14100);
nand U16685 (N_16685,N_14692,N_10538);
or U16686 (N_16686,N_14161,N_10122);
nor U16687 (N_16687,N_11547,N_11317);
nor U16688 (N_16688,N_14007,N_13547);
xor U16689 (N_16689,N_13419,N_12260);
nor U16690 (N_16690,N_11520,N_14885);
and U16691 (N_16691,N_10023,N_10868);
nand U16692 (N_16692,N_14750,N_13775);
nor U16693 (N_16693,N_13516,N_12878);
nand U16694 (N_16694,N_13500,N_14752);
nor U16695 (N_16695,N_14770,N_14308);
and U16696 (N_16696,N_13327,N_10032);
nand U16697 (N_16697,N_11670,N_10818);
nor U16698 (N_16698,N_12724,N_11094);
or U16699 (N_16699,N_10365,N_11771);
or U16700 (N_16700,N_13596,N_13359);
nand U16701 (N_16701,N_10950,N_10992);
nand U16702 (N_16702,N_14922,N_14683);
or U16703 (N_16703,N_10752,N_10790);
or U16704 (N_16704,N_13559,N_13617);
or U16705 (N_16705,N_12789,N_10193);
or U16706 (N_16706,N_12059,N_11227);
and U16707 (N_16707,N_13539,N_10074);
nor U16708 (N_16708,N_13080,N_13699);
and U16709 (N_16709,N_13822,N_12496);
and U16710 (N_16710,N_12402,N_12928);
nor U16711 (N_16711,N_12782,N_10440);
and U16712 (N_16712,N_14866,N_12170);
nand U16713 (N_16713,N_13066,N_14048);
or U16714 (N_16714,N_12606,N_14063);
nor U16715 (N_16715,N_12980,N_14689);
or U16716 (N_16716,N_11707,N_11183);
and U16717 (N_16717,N_14704,N_13391);
nand U16718 (N_16718,N_13108,N_10998);
nand U16719 (N_16719,N_13861,N_12183);
nand U16720 (N_16720,N_13393,N_10401);
nor U16721 (N_16721,N_14854,N_13469);
nand U16722 (N_16722,N_10902,N_12115);
and U16723 (N_16723,N_14710,N_11836);
nand U16724 (N_16724,N_12008,N_10285);
nor U16725 (N_16725,N_11920,N_11825);
nand U16726 (N_16726,N_12154,N_13430);
or U16727 (N_16727,N_11578,N_12081);
and U16728 (N_16728,N_14823,N_12199);
nand U16729 (N_16729,N_12603,N_12367);
nor U16730 (N_16730,N_11546,N_13135);
nor U16731 (N_16731,N_13258,N_10400);
and U16732 (N_16732,N_14891,N_10385);
xor U16733 (N_16733,N_13603,N_14803);
nor U16734 (N_16734,N_14859,N_12939);
nand U16735 (N_16735,N_10130,N_13716);
or U16736 (N_16736,N_13346,N_14448);
or U16737 (N_16737,N_12799,N_14499);
nand U16738 (N_16738,N_10146,N_10988);
nor U16739 (N_16739,N_14001,N_10610);
or U16740 (N_16740,N_14631,N_14461);
nand U16741 (N_16741,N_13945,N_10658);
and U16742 (N_16742,N_12571,N_12168);
nor U16743 (N_16743,N_12507,N_13049);
nand U16744 (N_16744,N_13690,N_10001);
nor U16745 (N_16745,N_10076,N_11389);
or U16746 (N_16746,N_12561,N_11053);
nor U16747 (N_16747,N_10907,N_11167);
nor U16748 (N_16748,N_12095,N_14027);
nor U16749 (N_16749,N_11954,N_12646);
nor U16750 (N_16750,N_11208,N_10093);
or U16751 (N_16751,N_14332,N_11975);
nand U16752 (N_16752,N_11437,N_12448);
or U16753 (N_16753,N_13147,N_13274);
nor U16754 (N_16754,N_10474,N_11806);
nand U16755 (N_16755,N_14465,N_11334);
and U16756 (N_16756,N_12622,N_10194);
nor U16757 (N_16757,N_11602,N_11204);
or U16758 (N_16758,N_10831,N_13107);
nand U16759 (N_16759,N_10837,N_11545);
nand U16760 (N_16760,N_14102,N_10226);
or U16761 (N_16761,N_10449,N_10229);
and U16762 (N_16762,N_13226,N_12410);
or U16763 (N_16763,N_13365,N_14180);
nor U16764 (N_16764,N_10951,N_13013);
and U16765 (N_16765,N_11807,N_14533);
nor U16766 (N_16766,N_14612,N_14197);
or U16767 (N_16767,N_13752,N_14040);
nor U16768 (N_16768,N_13347,N_12084);
and U16769 (N_16769,N_14542,N_13137);
nand U16770 (N_16770,N_14933,N_10842);
nand U16771 (N_16771,N_10891,N_12578);
nand U16772 (N_16772,N_11467,N_12379);
and U16773 (N_16773,N_11666,N_12620);
or U16774 (N_16774,N_12085,N_12424);
nor U16775 (N_16775,N_12841,N_12989);
nand U16776 (N_16776,N_11379,N_14697);
nor U16777 (N_16777,N_11721,N_11132);
and U16778 (N_16778,N_14019,N_11065);
xnor U16779 (N_16779,N_10210,N_12111);
nand U16780 (N_16780,N_11044,N_11931);
xnor U16781 (N_16781,N_12630,N_11735);
nor U16782 (N_16782,N_10117,N_11099);
and U16783 (N_16783,N_14012,N_13534);
xor U16784 (N_16784,N_10207,N_10408);
and U16785 (N_16785,N_14946,N_14699);
xor U16786 (N_16786,N_11346,N_12223);
or U16787 (N_16787,N_12144,N_12336);
nand U16788 (N_16788,N_11779,N_10953);
nor U16789 (N_16789,N_11168,N_14724);
and U16790 (N_16790,N_11147,N_11674);
nand U16791 (N_16791,N_10836,N_10958);
nand U16792 (N_16792,N_12241,N_12244);
or U16793 (N_16793,N_11737,N_10844);
xor U16794 (N_16794,N_11069,N_12491);
nor U16795 (N_16795,N_10906,N_14087);
and U16796 (N_16796,N_10237,N_11948);
and U16797 (N_16797,N_10295,N_12205);
and U16798 (N_16798,N_13847,N_13653);
or U16799 (N_16799,N_14615,N_11051);
nand U16800 (N_16800,N_10630,N_12056);
nor U16801 (N_16801,N_12931,N_11972);
or U16802 (N_16802,N_14458,N_10441);
nand U16803 (N_16803,N_13703,N_12846);
or U16804 (N_16804,N_13324,N_12021);
nor U16805 (N_16805,N_12770,N_11494);
or U16806 (N_16806,N_14192,N_10566);
and U16807 (N_16807,N_10437,N_12215);
or U16808 (N_16808,N_10489,N_13832);
and U16809 (N_16809,N_13507,N_14921);
nor U16810 (N_16810,N_13665,N_12566);
nor U16811 (N_16811,N_12951,N_10232);
nor U16812 (N_16812,N_11313,N_11872);
nor U16813 (N_16813,N_14872,N_10362);
or U16814 (N_16814,N_14483,N_14818);
or U16815 (N_16815,N_13123,N_10044);
nor U16816 (N_16816,N_11556,N_13809);
or U16817 (N_16817,N_13426,N_11414);
nand U16818 (N_16818,N_11700,N_10149);
nor U16819 (N_16819,N_11532,N_13907);
and U16820 (N_16820,N_12461,N_12378);
and U16821 (N_16821,N_14118,N_14166);
and U16822 (N_16822,N_11754,N_12002);
and U16823 (N_16823,N_10415,N_12079);
and U16824 (N_16824,N_14701,N_11197);
or U16825 (N_16825,N_14270,N_10473);
nand U16826 (N_16826,N_11617,N_13179);
and U16827 (N_16827,N_10669,N_13006);
or U16828 (N_16828,N_12746,N_13570);
or U16829 (N_16829,N_11046,N_11993);
nor U16830 (N_16830,N_11114,N_12876);
or U16831 (N_16831,N_12450,N_11839);
or U16832 (N_16832,N_13018,N_14630);
or U16833 (N_16833,N_14368,N_11688);
nor U16834 (N_16834,N_14940,N_14782);
or U16835 (N_16835,N_13881,N_11283);
or U16836 (N_16836,N_12885,N_11860);
and U16837 (N_16837,N_13942,N_11382);
and U16838 (N_16838,N_12974,N_14643);
and U16839 (N_16839,N_14472,N_13320);
and U16840 (N_16840,N_13411,N_10214);
nor U16841 (N_16841,N_12250,N_14350);
or U16842 (N_16842,N_14831,N_10871);
and U16843 (N_16843,N_12807,N_14669);
nand U16844 (N_16844,N_13251,N_12156);
nor U16845 (N_16845,N_12146,N_10931);
nand U16846 (N_16846,N_13206,N_10293);
nor U16847 (N_16847,N_12306,N_11424);
or U16848 (N_16848,N_12917,N_14844);
or U16849 (N_16849,N_12102,N_10964);
and U16850 (N_16850,N_12209,N_14705);
nand U16851 (N_16851,N_12739,N_10929);
and U16852 (N_16852,N_13423,N_10766);
nor U16853 (N_16853,N_12387,N_13937);
xor U16854 (N_16854,N_13730,N_14830);
and U16855 (N_16855,N_11747,N_10345);
nand U16856 (N_16856,N_14424,N_11951);
nor U16857 (N_16857,N_14112,N_13870);
nand U16858 (N_16858,N_10957,N_12262);
nor U16859 (N_16859,N_14008,N_12314);
nand U16860 (N_16860,N_12172,N_10342);
or U16861 (N_16861,N_12482,N_12251);
nand U16862 (N_16862,N_12823,N_13356);
nand U16863 (N_16863,N_11022,N_13845);
and U16864 (N_16864,N_14847,N_13933);
and U16865 (N_16865,N_10349,N_10383);
nand U16866 (N_16866,N_13501,N_10218);
nor U16867 (N_16867,N_10580,N_10700);
and U16868 (N_16868,N_12106,N_10172);
nand U16869 (N_16869,N_12725,N_11623);
nand U16870 (N_16870,N_13302,N_14833);
and U16871 (N_16871,N_12501,N_13719);
nor U16872 (N_16872,N_12451,N_12787);
nand U16873 (N_16873,N_12088,N_13895);
nand U16874 (N_16874,N_13798,N_11691);
and U16875 (N_16875,N_13313,N_11027);
and U16876 (N_16876,N_10442,N_14227);
or U16877 (N_16877,N_14176,N_10643);
or U16878 (N_16878,N_10739,N_11399);
and U16879 (N_16879,N_12151,N_11392);
nand U16880 (N_16880,N_12788,N_14389);
nor U16881 (N_16881,N_12504,N_13371);
nand U16882 (N_16882,N_11724,N_13282);
or U16883 (N_16883,N_13667,N_10692);
and U16884 (N_16884,N_10220,N_14014);
nor U16885 (N_16885,N_13993,N_14819);
and U16886 (N_16886,N_14184,N_10758);
nor U16887 (N_16887,N_13683,N_14747);
and U16888 (N_16888,N_12926,N_12744);
nand U16889 (N_16889,N_10435,N_12003);
and U16890 (N_16890,N_14246,N_14796);
or U16891 (N_16891,N_14912,N_11897);
and U16892 (N_16892,N_11113,N_14824);
or U16893 (N_16893,N_11259,N_11770);
nand U16894 (N_16894,N_14154,N_11535);
nand U16895 (N_16895,N_10516,N_14974);
and U16896 (N_16896,N_11795,N_11398);
and U16897 (N_16897,N_10773,N_12669);
or U16898 (N_16898,N_10015,N_10470);
nor U16899 (N_16899,N_11918,N_11856);
nand U16900 (N_16900,N_14656,N_13046);
nor U16901 (N_16901,N_14481,N_14437);
or U16902 (N_16902,N_11957,N_10945);
nor U16903 (N_16903,N_11016,N_12999);
xor U16904 (N_16904,N_11965,N_13096);
and U16905 (N_16905,N_14878,N_14568);
nand U16906 (N_16906,N_10694,N_11350);
and U16907 (N_16907,N_14133,N_14696);
and U16908 (N_16908,N_14932,N_12524);
nand U16909 (N_16909,N_11668,N_13077);
or U16910 (N_16910,N_12176,N_13919);
or U16911 (N_16911,N_14887,N_12020);
nand U16912 (N_16912,N_10974,N_10157);
nor U16913 (N_16913,N_14990,N_14812);
or U16914 (N_16914,N_13261,N_12142);
and U16915 (N_16915,N_10506,N_13330);
nor U16916 (N_16916,N_13221,N_12394);
nor U16917 (N_16917,N_11332,N_11732);
nand U16918 (N_16918,N_13270,N_10640);
and U16919 (N_16919,N_10802,N_10198);
and U16920 (N_16920,N_12866,N_13604);
nand U16921 (N_16921,N_12352,N_12435);
or U16922 (N_16922,N_13750,N_13884);
nor U16923 (N_16923,N_14372,N_14998);
and U16924 (N_16924,N_11949,N_13949);
or U16925 (N_16925,N_11588,N_12181);
and U16926 (N_16926,N_13705,N_13214);
or U16927 (N_16927,N_14381,N_10060);
nand U16928 (N_16928,N_12605,N_12338);
and U16929 (N_16929,N_13310,N_12411);
or U16930 (N_16930,N_10243,N_13262);
or U16931 (N_16931,N_10055,N_14486);
or U16932 (N_16932,N_11343,N_10498);
or U16933 (N_16933,N_11620,N_12890);
nand U16934 (N_16934,N_13161,N_11029);
nand U16935 (N_16935,N_12417,N_10940);
or U16936 (N_16936,N_12801,N_10259);
nor U16937 (N_16937,N_10182,N_11443);
or U16938 (N_16938,N_14591,N_10791);
nand U16939 (N_16939,N_11680,N_10977);
or U16940 (N_16940,N_11801,N_14732);
nand U16941 (N_16941,N_12017,N_12883);
or U16942 (N_16942,N_14649,N_13833);
nor U16943 (N_16943,N_13592,N_14647);
and U16944 (N_16944,N_11678,N_11351);
or U16945 (N_16945,N_11047,N_12366);
or U16946 (N_16946,N_14122,N_13309);
nor U16947 (N_16947,N_11371,N_11206);
and U16948 (N_16948,N_14945,N_14507);
and U16949 (N_16949,N_14016,N_12690);
nor U16950 (N_16950,N_11849,N_13578);
nand U16951 (N_16951,N_14094,N_12325);
nor U16952 (N_16952,N_10704,N_13702);
nand U16953 (N_16953,N_13272,N_14515);
and U16954 (N_16954,N_14576,N_13002);
and U16955 (N_16955,N_13926,N_12202);
and U16956 (N_16956,N_10376,N_13846);
and U16957 (N_16957,N_11610,N_13466);
nand U16958 (N_16958,N_10698,N_10772);
and U16959 (N_16959,N_11435,N_11585);
and U16960 (N_16960,N_11111,N_10680);
and U16961 (N_16961,N_14815,N_10078);
nand U16962 (N_16962,N_10192,N_10083);
nor U16963 (N_16963,N_10317,N_11614);
nor U16964 (N_16964,N_13515,N_10986);
or U16965 (N_16965,N_11001,N_10865);
nand U16966 (N_16966,N_12754,N_10816);
nor U16967 (N_16967,N_11762,N_13793);
and U16968 (N_16968,N_13257,N_10651);
or U16969 (N_16969,N_11049,N_11312);
and U16970 (N_16970,N_14534,N_13374);
nor U16971 (N_16971,N_14468,N_10368);
and U16972 (N_16972,N_12090,N_13048);
or U16973 (N_16973,N_10529,N_14013);
nor U16974 (N_16974,N_10713,N_14268);
nand U16975 (N_16975,N_12233,N_12447);
nor U16976 (N_16976,N_12973,N_13726);
nor U16977 (N_16977,N_14388,N_13760);
nor U16978 (N_16978,N_11288,N_11039);
or U16979 (N_16979,N_13879,N_13513);
or U16980 (N_16980,N_14347,N_10925);
and U16981 (N_16981,N_11403,N_12470);
or U16982 (N_16982,N_14452,N_11429);
or U16983 (N_16983,N_12315,N_11675);
and U16984 (N_16984,N_14645,N_14403);
or U16985 (N_16985,N_12859,N_13679);
nand U16986 (N_16986,N_11626,N_10822);
or U16987 (N_16987,N_13777,N_12587);
nand U16988 (N_16988,N_12163,N_12638);
and U16989 (N_16989,N_12150,N_10653);
or U16990 (N_16990,N_10370,N_14962);
nand U16991 (N_16991,N_14098,N_10079);
or U16992 (N_16992,N_10503,N_11765);
and U16993 (N_16993,N_12069,N_14557);
nor U16994 (N_16994,N_14139,N_10269);
or U16995 (N_16995,N_14362,N_14904);
and U16996 (N_16996,N_12715,N_13704);
nor U16997 (N_16997,N_10283,N_14208);
or U16998 (N_16998,N_14479,N_14160);
xnor U16999 (N_16999,N_14956,N_11925);
nor U17000 (N_17000,N_11340,N_14848);
or U17001 (N_17001,N_12633,N_13663);
nand U17002 (N_17002,N_13893,N_14285);
or U17003 (N_17003,N_10869,N_10714);
or U17004 (N_17004,N_12721,N_12455);
nor U17005 (N_17005,N_13674,N_10983);
nor U17006 (N_17006,N_11095,N_14771);
or U17007 (N_17007,N_12582,N_14398);
or U17008 (N_17008,N_14343,N_12288);
nand U17009 (N_17009,N_11305,N_11468);
nand U17010 (N_17010,N_12027,N_13960);
and U17011 (N_17011,N_13892,N_13523);
or U17012 (N_17012,N_11953,N_14624);
nor U17013 (N_17013,N_13265,N_11296);
nor U17014 (N_17014,N_10759,N_13508);
nor U17015 (N_17015,N_13418,N_11544);
or U17016 (N_17016,N_13885,N_13099);
and U17017 (N_17017,N_11339,N_13495);
nand U17018 (N_17018,N_13673,N_12075);
or U17019 (N_17019,N_10564,N_14646);
nand U17020 (N_17020,N_11542,N_14364);
nor U17021 (N_17021,N_10255,N_13605);
and U17022 (N_17022,N_13535,N_13684);
and U17023 (N_17023,N_14314,N_10598);
and U17024 (N_17024,N_13910,N_10505);
nor U17025 (N_17025,N_14965,N_11728);
nand U17026 (N_17026,N_11263,N_10037);
nor U17027 (N_17027,N_11753,N_14648);
nand U17028 (N_17028,N_13649,N_12942);
and U17029 (N_17029,N_12812,N_13398);
and U17030 (N_17030,N_13823,N_13331);
nand U17031 (N_17031,N_10712,N_12750);
nor U17032 (N_17032,N_12279,N_14428);
nand U17033 (N_17033,N_11074,N_12356);
and U17034 (N_17034,N_10756,N_10234);
and U17035 (N_17035,N_14580,N_11038);
nand U17036 (N_17036,N_14996,N_12245);
nor U17037 (N_17037,N_14659,N_14559);
xor U17038 (N_17038,N_13319,N_10444);
and U17039 (N_17039,N_10823,N_11903);
nand U17040 (N_17040,N_11519,N_14497);
nand U17041 (N_17041,N_10531,N_12558);
and U17042 (N_17042,N_13348,N_11511);
or U17043 (N_17043,N_14851,N_12722);
and U17044 (N_17044,N_11098,N_14224);
or U17045 (N_17045,N_10764,N_13271);
nor U17046 (N_17046,N_11503,N_14550);
and U17047 (N_17047,N_13200,N_14146);
nand U17048 (N_17048,N_11130,N_11500);
nor U17049 (N_17049,N_10612,N_10645);
or U17050 (N_17050,N_10873,N_10406);
nand U17051 (N_17051,N_14589,N_13889);
nor U17052 (N_17052,N_12695,N_11439);
or U17053 (N_17053,N_11410,N_12593);
nand U17054 (N_17054,N_12718,N_13435);
or U17055 (N_17055,N_14341,N_11526);
or U17056 (N_17056,N_13740,N_10749);
nor U17057 (N_17057,N_12824,N_10284);
or U17058 (N_17058,N_12934,N_10574);
nor U17059 (N_17059,N_12688,N_14010);
or U17060 (N_17060,N_11441,N_11119);
nor U17061 (N_17061,N_11393,N_12896);
or U17062 (N_17062,N_10862,N_10995);
or U17063 (N_17063,N_14392,N_10711);
or U17064 (N_17064,N_14874,N_12211);
or U17065 (N_17065,N_14610,N_14744);
and U17066 (N_17066,N_13223,N_11276);
nand U17067 (N_17067,N_14143,N_11820);
and U17068 (N_17068,N_14064,N_10205);
nand U17069 (N_17069,N_12656,N_13773);
and U17070 (N_17070,N_13932,N_13537);
and U17071 (N_17071,N_11992,N_10250);
or U17072 (N_17072,N_13112,N_14952);
xnor U17073 (N_17073,N_12016,N_14211);
and U17074 (N_17074,N_10485,N_13369);
or U17075 (N_17075,N_14531,N_14057);
and U17076 (N_17076,N_13043,N_13473);
or U17077 (N_17077,N_10681,N_11252);
nand U17078 (N_17078,N_13961,N_12616);
nand U17079 (N_17079,N_10025,N_12475);
and U17080 (N_17080,N_10002,N_13480);
or U17081 (N_17081,N_12565,N_11081);
nor U17082 (N_17082,N_11981,N_11090);
xor U17083 (N_17083,N_14541,N_12993);
and U17084 (N_17084,N_10987,N_13340);
nor U17085 (N_17085,N_11769,N_12861);
or U17086 (N_17086,N_10315,N_10615);
or U17087 (N_17087,N_10356,N_10776);
nand U17088 (N_17088,N_11841,N_11472);
and U17089 (N_17089,N_13666,N_11529);
and U17090 (N_17090,N_10890,N_13542);
nand U17091 (N_17091,N_10703,N_10453);
and U17092 (N_17092,N_12230,N_10722);
nor U17093 (N_17093,N_10119,N_10101);
nand U17094 (N_17094,N_11913,N_13616);
and U17095 (N_17095,N_13318,N_11273);
nand U17096 (N_17096,N_13734,N_12186);
nor U17097 (N_17097,N_12862,N_13124);
nor U17098 (N_17098,N_10371,N_10546);
and U17099 (N_17099,N_11819,N_12710);
nand U17100 (N_17100,N_12783,N_13621);
and U17101 (N_17101,N_13790,N_13482);
or U17102 (N_17102,N_11551,N_12918);
nand U17103 (N_17103,N_12991,N_12194);
or U17104 (N_17104,N_14662,N_10867);
nor U17105 (N_17105,N_11320,N_11471);
nand U17106 (N_17106,N_12025,N_11287);
nor U17107 (N_17107,N_13130,N_13127);
or U17108 (N_17108,N_13341,N_10648);
or U17109 (N_17109,N_10013,N_12624);
or U17110 (N_17110,N_13852,N_14420);
xnor U17111 (N_17111,N_13628,N_14076);
nor U17112 (N_17112,N_13748,N_10624);
nand U17113 (N_17113,N_10393,N_14980);
or U17114 (N_17114,N_12621,N_12427);
and U17115 (N_17115,N_10199,N_10212);
nor U17116 (N_17116,N_13718,N_12464);
or U17117 (N_17117,N_13167,N_11938);
nand U17118 (N_17118,N_13328,N_13451);
or U17119 (N_17119,N_13771,N_10848);
nand U17120 (N_17120,N_12596,N_12028);
nor U17121 (N_17121,N_11880,N_12822);
or U17122 (N_17122,N_10525,N_13600);
and U17123 (N_17123,N_14546,N_11501);
nand U17124 (N_17124,N_12680,N_13765);
nand U17125 (N_17125,N_11314,N_10644);
or U17126 (N_17126,N_14709,N_14181);
nand U17127 (N_17127,N_12108,N_11996);
xnor U17128 (N_17128,N_11396,N_11413);
or U17129 (N_17129,N_14266,N_12771);
nand U17130 (N_17130,N_14021,N_10960);
or U17131 (N_17131,N_12114,N_11745);
nand U17132 (N_17132,N_10189,N_10980);
or U17133 (N_17133,N_11879,N_14374);
or U17134 (N_17134,N_10045,N_10595);
and U17135 (N_17135,N_12562,N_11929);
xor U17136 (N_17136,N_11850,N_14429);
nand U17137 (N_17137,N_11813,N_11160);
nor U17138 (N_17138,N_11782,N_13905);
nor U17139 (N_17139,N_10041,N_14178);
and U17140 (N_17140,N_14054,N_11318);
and U17141 (N_17141,N_11648,N_10609);
nand U17142 (N_17142,N_13584,N_13031);
nor U17143 (N_17143,N_14431,N_11597);
and U17144 (N_17144,N_12597,N_13205);
and U17145 (N_17145,N_11203,N_12473);
or U17146 (N_17146,N_10417,N_11013);
nor U17147 (N_17147,N_11604,N_11763);
and U17148 (N_17148,N_14834,N_14558);
nand U17149 (N_17149,N_11633,N_14339);
xor U17150 (N_17150,N_11804,N_10239);
nand U17151 (N_17151,N_13183,N_12217);
or U17152 (N_17152,N_12685,N_11482);
and U17153 (N_17153,N_11387,N_11884);
nand U17154 (N_17154,N_11256,N_13180);
and U17155 (N_17155,N_11584,N_13160);
or U17156 (N_17156,N_12540,N_11673);
and U17157 (N_17157,N_13069,N_11577);
or U17158 (N_17158,N_11357,N_13856);
nand U17159 (N_17159,N_12292,N_10069);
and U17160 (N_17160,N_14766,N_11589);
and U17161 (N_17161,N_11134,N_14042);
or U17162 (N_17162,N_11650,N_10084);
nor U17163 (N_17163,N_14185,N_12390);
and U17164 (N_17164,N_11409,N_12255);
and U17165 (N_17165,N_11694,N_12546);
nor U17166 (N_17166,N_12304,N_12113);
or U17167 (N_17167,N_13850,N_14336);
nor U17168 (N_17168,N_10366,N_10114);
xnor U17169 (N_17169,N_12714,N_13421);
or U17170 (N_17170,N_13497,N_14527);
xnor U17171 (N_17171,N_14459,N_10501);
and U17172 (N_17172,N_12375,N_12497);
and U17173 (N_17173,N_11226,N_13382);
or U17174 (N_17174,N_13655,N_11209);
and U17175 (N_17175,N_10935,N_14622);
nand U17176 (N_17176,N_10059,N_10231);
or U17177 (N_17177,N_11874,N_11152);
and U17178 (N_17178,N_12311,N_10666);
and U17179 (N_17179,N_11815,N_12124);
or U17180 (N_17180,N_13736,N_12759);
nor U17181 (N_17181,N_11258,N_12195);
or U17182 (N_17182,N_13456,N_10392);
or U17183 (N_17183,N_12316,N_12815);
and U17184 (N_17184,N_14563,N_10476);
and U17185 (N_17185,N_10052,N_14713);
or U17186 (N_17186,N_10357,N_10835);
nor U17187 (N_17187,N_10793,N_11711);
and U17188 (N_17188,N_13831,N_14279);
or U17189 (N_17189,N_12018,N_10984);
nor U17190 (N_17190,N_10927,N_10627);
nor U17191 (N_17191,N_12133,N_13687);
nor U17192 (N_17192,N_13817,N_14159);
or U17193 (N_17193,N_12453,N_14242);
and U17194 (N_17194,N_12575,N_11274);
nor U17195 (N_17195,N_11601,N_14743);
or U17196 (N_17196,N_11646,N_12137);
nor U17197 (N_17197,N_11141,N_14215);
or U17198 (N_17198,N_13120,N_13610);
or U17199 (N_17199,N_11621,N_14768);
nor U17200 (N_17200,N_12500,N_11808);
nand U17201 (N_17201,N_14121,N_10304);
or U17202 (N_17202,N_14356,N_13225);
nor U17203 (N_17203,N_10577,N_10278);
and U17204 (N_17204,N_14687,N_14360);
nand U17205 (N_17205,N_14694,N_14931);
nand U17206 (N_17206,N_13412,N_12180);
or U17207 (N_17207,N_10107,N_12407);
or U17208 (N_17208,N_14655,N_12243);
nand U17209 (N_17209,N_10999,N_11906);
nor U17210 (N_17210,N_13660,N_10858);
or U17211 (N_17211,N_10372,N_14902);
and U17212 (N_17212,N_13839,N_12627);
nand U17213 (N_17213,N_11896,N_10727);
or U17214 (N_17214,N_14150,N_13196);
nand U17215 (N_17215,N_11442,N_14387);
nor U17216 (N_17216,N_14740,N_12766);
nand U17217 (N_17217,N_12930,N_12547);
nand U17218 (N_17218,N_13857,N_12877);
nor U17219 (N_17219,N_14449,N_11612);
nor U17220 (N_17220,N_12462,N_13721);
xor U17221 (N_17221,N_11262,N_12253);
nor U17222 (N_17222,N_14171,N_11178);
or U17223 (N_17223,N_14441,N_12395);
nor U17224 (N_17224,N_14269,N_14142);
nor U17225 (N_17225,N_13185,N_12682);
nor U17226 (N_17226,N_12933,N_13448);
or U17227 (N_17227,N_10716,N_12023);
nand U17228 (N_17228,N_10017,N_10100);
nor U17229 (N_17229,N_10602,N_10176);
nor U17230 (N_17230,N_12732,N_13986);
or U17231 (N_17231,N_11516,N_14606);
nand U17232 (N_17232,N_11266,N_11151);
nor U17233 (N_17233,N_14593,N_14026);
nor U17234 (N_17234,N_11525,N_13711);
or U17235 (N_17235,N_12105,N_11063);
nor U17236 (N_17236,N_13981,N_12850);
and U17237 (N_17237,N_14316,N_12119);
and U17238 (N_17238,N_12662,N_13036);
nor U17239 (N_17239,N_12836,N_14052);
or U17240 (N_17240,N_13361,N_10096);
nand U17241 (N_17241,N_11315,N_13442);
nor U17242 (N_17242,N_14254,N_12235);
nor U17243 (N_17243,N_11509,N_13802);
or U17244 (N_17244,N_14798,N_10763);
or U17245 (N_17245,N_11704,N_11508);
nand U17246 (N_17246,N_11390,N_13583);
and U17247 (N_17247,N_11257,N_12667);
and U17248 (N_17248,N_11562,N_11495);
nand U17249 (N_17249,N_14970,N_12860);
nand U17250 (N_17250,N_14450,N_12604);
and U17251 (N_17251,N_10832,N_12661);
nand U17252 (N_17252,N_11391,N_10629);
nor U17253 (N_17253,N_14720,N_13122);
and U17254 (N_17254,N_10047,N_14575);
nor U17255 (N_17255,N_10854,N_10571);
nand U17256 (N_17256,N_11738,N_11568);
and U17257 (N_17257,N_11997,N_10369);
or U17258 (N_17258,N_11565,N_14617);
or U17259 (N_17259,N_14011,N_11631);
nand U17260 (N_17260,N_12756,N_12048);
nor U17261 (N_17261,N_10838,N_10537);
or U17262 (N_17262,N_13085,N_13796);
xnor U17263 (N_17263,N_11316,N_10344);
or U17264 (N_17264,N_14091,N_12436);
nand U17265 (N_17265,N_14547,N_12897);
nor U17266 (N_17266,N_13632,N_13819);
and U17267 (N_17267,N_12647,N_13338);
and U17268 (N_17268,N_10487,N_13119);
nand U17269 (N_17269,N_13787,N_14599);
and U17270 (N_17270,N_13897,N_12444);
or U17271 (N_17271,N_11248,N_10108);
and U17272 (N_17272,N_11352,N_14267);
or U17273 (N_17273,N_13692,N_14973);
and U17274 (N_17274,N_13493,N_14873);
and U17275 (N_17275,N_13866,N_11269);
or U17276 (N_17276,N_10190,N_13082);
and U17277 (N_17277,N_13637,N_14574);
and U17278 (N_17278,N_14512,N_12029);
or U17279 (N_17279,N_11175,N_14132);
nor U17280 (N_17280,N_13522,N_14552);
or U17281 (N_17281,N_13000,N_10982);
or U17282 (N_17282,N_13483,N_10728);
or U17283 (N_17283,N_13001,N_13571);
nand U17284 (N_17284,N_10163,N_11766);
xnor U17285 (N_17285,N_12221,N_11887);
nand U17286 (N_17286,N_11362,N_12031);
or U17287 (N_17287,N_13503,N_10784);
nor U17288 (N_17288,N_13045,N_14155);
nor U17289 (N_17289,N_11077,N_10057);
nor U17290 (N_17290,N_13053,N_12618);
or U17291 (N_17291,N_11580,N_14213);
nand U17292 (N_17292,N_10490,N_10495);
nand U17293 (N_17293,N_13022,N_11153);
and U17294 (N_17294,N_14363,N_12351);
or U17295 (N_17295,N_10576,N_11322);
nor U17296 (N_17296,N_12673,N_13026);
and U17297 (N_17297,N_11566,N_11221);
nand U17298 (N_17298,N_12905,N_11144);
or U17299 (N_17299,N_13438,N_10432);
or U17300 (N_17300,N_14104,N_10482);
or U17301 (N_17301,N_12143,N_14581);
nand U17302 (N_17302,N_14979,N_10343);
or U17303 (N_17303,N_13804,N_10095);
nor U17304 (N_17304,N_11693,N_13410);
and U17305 (N_17305,N_12127,N_12177);
nand U17306 (N_17306,N_10853,N_11199);
nand U17307 (N_17307,N_14051,N_14584);
or U17308 (N_17308,N_14855,N_13612);
and U17309 (N_17309,N_14106,N_13023);
or U17310 (N_17310,N_10590,N_12645);
nor U17311 (N_17311,N_10493,N_14239);
nand U17312 (N_17312,N_13920,N_13553);
or U17313 (N_17313,N_13496,N_13420);
nand U17314 (N_17314,N_13735,N_11990);
and U17315 (N_17315,N_12313,N_11682);
or U17316 (N_17316,N_10775,N_10774);
or U17317 (N_17317,N_12936,N_11415);
and U17318 (N_17318,N_13883,N_11649);
and U17319 (N_17319,N_14325,N_10781);
nand U17320 (N_17320,N_13485,N_13012);
and U17321 (N_17321,N_14678,N_11768);
or U17322 (N_17322,N_10579,N_11911);
and U17323 (N_17323,N_11563,N_10054);
nor U17324 (N_17324,N_13413,N_14537);
nor U17325 (N_17325,N_11284,N_12047);
or U17326 (N_17326,N_13994,N_11637);
and U17327 (N_17327,N_10087,N_11394);
xor U17328 (N_17328,N_12580,N_12691);
or U17329 (N_17329,N_12584,N_10922);
and U17330 (N_17330,N_10533,N_14407);
or U17331 (N_17331,N_12839,N_14189);
nand U17332 (N_17332,N_11365,N_14733);
and U17333 (N_17333,N_14828,N_10611);
or U17334 (N_17334,N_11213,N_14188);
and U17335 (N_17335,N_12373,N_12731);
nand U17336 (N_17336,N_11755,N_13565);
nand U17337 (N_17337,N_11041,N_12712);
and U17338 (N_17338,N_13383,N_14442);
and U17339 (N_17339,N_10668,N_12709);
nor U17340 (N_17340,N_13646,N_14698);
and U17341 (N_17341,N_13436,N_11855);
nor U17342 (N_17342,N_14985,N_10450);
and U17343 (N_17343,N_13954,N_10535);
nand U17344 (N_17344,N_12659,N_13005);
xor U17345 (N_17345,N_11280,N_12997);
and U17346 (N_17346,N_12923,N_11702);
or U17347 (N_17347,N_12409,N_12276);
nand U17348 (N_17348,N_13569,N_12539);
or U17349 (N_17349,N_10135,N_12165);
nand U17350 (N_17350,N_14637,N_13980);
nor U17351 (N_17351,N_13574,N_14861);
and U17352 (N_17352,N_11101,N_12555);
and U17353 (N_17353,N_12269,N_13835);
and U17354 (N_17354,N_13139,N_14899);
and U17355 (N_17355,N_12665,N_12748);
and U17356 (N_17356,N_13779,N_12398);
and U17357 (N_17357,N_13468,N_14231);
or U17358 (N_17358,N_11230,N_14069);
or U17359 (N_17359,N_14205,N_13998);
nor U17360 (N_17360,N_12458,N_11067);
nor U17361 (N_17361,N_13855,N_13851);
or U17362 (N_17362,N_10496,N_13917);
and U17363 (N_17363,N_11950,N_14817);
and U17364 (N_17364,N_13974,N_12348);
nor U17365 (N_17365,N_10337,N_13401);
nor U17366 (N_17366,N_10901,N_11961);
nor U17367 (N_17367,N_13589,N_13678);
or U17368 (N_17368,N_14916,N_11869);
nor U17369 (N_17369,N_11934,N_10134);
and U17370 (N_17370,N_13642,N_12779);
nand U17371 (N_17371,N_10286,N_10683);
nor U17372 (N_17372,N_10133,N_13874);
or U17373 (N_17373,N_11083,N_11139);
and U17374 (N_17374,N_12149,N_11405);
nor U17375 (N_17375,N_13557,N_10123);
nand U17376 (N_17376,N_11593,N_10534);
nor U17377 (N_17377,N_11805,N_14735);
or U17378 (N_17378,N_13489,N_14303);
and U17379 (N_17379,N_10246,N_11717);
nor U17380 (N_17380,N_14418,N_10677);
nor U17381 (N_17381,N_10411,N_14758);
or U17382 (N_17382,N_13240,N_12213);
nor U17383 (N_17383,N_12769,N_14915);
and U17384 (N_17384,N_13433,N_10597);
nand U17385 (N_17385,N_14273,N_11552);
and U17386 (N_17386,N_14218,N_13918);
or U17387 (N_17387,N_14814,N_12515);
nor U17388 (N_17388,N_12043,N_14711);
nor U17389 (N_17389,N_13946,N_12278);
and U17390 (N_17390,N_10185,N_12827);
nor U17391 (N_17391,N_13514,N_10173);
nand U17392 (N_17392,N_11086,N_11539);
nor U17393 (N_17393,N_11355,N_13197);
nand U17394 (N_17394,N_13556,N_10316);
nor U17395 (N_17395,N_13502,N_12847);
or U17396 (N_17396,N_11716,N_13756);
nor U17397 (N_17397,N_14826,N_12038);
nand U17398 (N_17398,N_14047,N_13155);
and U17399 (N_17399,N_11235,N_10956);
or U17400 (N_17400,N_13914,N_10741);
nor U17401 (N_17401,N_12426,N_14477);
and U17402 (N_17402,N_10825,N_12752);
nor U17403 (N_17403,N_12880,N_14820);
and U17404 (N_17404,N_14731,N_10167);
and U17405 (N_17405,N_12938,N_13414);
or U17406 (N_17406,N_12912,N_13560);
and U17407 (N_17407,N_12956,N_10202);
nor U17408 (N_17408,N_13336,N_13102);
xor U17409 (N_17409,N_11722,N_11112);
and U17410 (N_17410,N_11647,N_14871);
or U17411 (N_17411,N_14772,N_14686);
or U17412 (N_17412,N_14603,N_14633);
or U17413 (N_17413,N_10171,N_13362);
and U17414 (N_17414,N_13279,N_10492);
nand U17415 (N_17415,N_14494,N_12323);
nand U17416 (N_17416,N_13634,N_13877);
nand U17417 (N_17417,N_12743,N_11333);
xnor U17418 (N_17418,N_11878,N_14536);
nand U17419 (N_17419,N_14890,N_13030);
and U17420 (N_17420,N_13432,N_11202);
nand U17421 (N_17421,N_12468,N_13720);
and U17422 (N_17422,N_14806,N_12687);
nor U17423 (N_17423,N_14258,N_14836);
nand U17424 (N_17424,N_10067,N_10706);
xor U17425 (N_17425,N_11243,N_11917);
nor U17426 (N_17426,N_13229,N_10695);
nor U17427 (N_17427,N_12198,N_12196);
or U17428 (N_17428,N_11709,N_12511);
nand U17429 (N_17429,N_11970,N_12030);
nor U17430 (N_17430,N_11231,N_10914);
nand U17431 (N_17431,N_14717,N_14078);
nor U17432 (N_17432,N_10912,N_10993);
nand U17433 (N_17433,N_13198,N_12851);
nor U17434 (N_17434,N_13392,N_11937);
nor U17435 (N_17435,N_12651,N_14177);
nor U17436 (N_17436,N_11783,N_14451);
nor U17437 (N_17437,N_13222,N_12355);
and U17438 (N_17438,N_14319,N_12576);
nor U17439 (N_17439,N_11792,N_10358);
nand U17440 (N_17440,N_11303,N_10204);
nand U17441 (N_17441,N_12816,N_14582);
xnor U17442 (N_17442,N_12187,N_11660);
nand U17443 (N_17443,N_14923,N_12434);
and U17444 (N_17444,N_13169,N_10036);
and U17445 (N_17445,N_12128,N_14517);
and U17446 (N_17446,N_11233,N_12019);
and U17447 (N_17447,N_14736,N_14489);
and U17448 (N_17448,N_14320,N_14728);
and U17449 (N_17449,N_11140,N_12706);
or U17450 (N_17450,N_13992,N_12953);
nor U17451 (N_17451,N_10878,N_10077);
nand U17452 (N_17452,N_14071,N_10875);
and U17453 (N_17453,N_14349,N_10389);
nor U17454 (N_17454,N_11842,N_14311);
and U17455 (N_17455,N_11402,N_10268);
and U17456 (N_17456,N_14397,N_11245);
or U17457 (N_17457,N_10168,N_14882);
nand U17458 (N_17458,N_11821,N_13455);
and U17459 (N_17459,N_10767,N_10089);
and U17460 (N_17460,N_13636,N_12875);
nor U17461 (N_17461,N_13848,N_10997);
nand U17462 (N_17462,N_10038,N_14762);
and U17463 (N_17463,N_11211,N_10034);
and U17464 (N_17464,N_10247,N_12283);
and U17465 (N_17465,N_11576,N_11502);
nor U17466 (N_17466,N_10740,N_10943);
and U17467 (N_17467,N_13941,N_10391);
nand U17468 (N_17468,N_14369,N_11645);
nand U17469 (N_17469,N_10662,N_13439);
nand U17470 (N_17470,N_14715,N_12810);
or U17471 (N_17471,N_11686,N_11958);
nor U17472 (N_17472,N_13904,N_10049);
nor U17473 (N_17473,N_12683,N_14190);
nor U17474 (N_17474,N_13676,N_10655);
or U17475 (N_17475,N_10765,N_11341);
or U17476 (N_17476,N_14130,N_11164);
nor U17477 (N_17477,N_10144,N_11150);
and U17478 (N_17478,N_10933,N_13156);
or U17479 (N_17479,N_12726,N_14138);
nor U17480 (N_17480,N_12207,N_10910);
and U17481 (N_17481,N_11798,N_12399);
or U17482 (N_17482,N_14926,N_13157);
or U17483 (N_17483,N_14971,N_11619);
and U17484 (N_17484,N_11976,N_14045);
and U17485 (N_17485,N_12707,N_13276);
and U17486 (N_17486,N_14975,N_14856);
or U17487 (N_17487,N_11416,N_11848);
and U17488 (N_17488,N_13727,N_11195);
nand U17489 (N_17489,N_11497,N_10140);
and U17490 (N_17490,N_11986,N_11096);
nor U17491 (N_17491,N_12808,N_14037);
nor U17492 (N_17492,N_11353,N_13165);
or U17493 (N_17493,N_10329,N_13871);
nand U17494 (N_17494,N_10380,N_11829);
nand U17495 (N_17495,N_10970,N_14522);
nor U17496 (N_17496,N_14137,N_14644);
nand U17497 (N_17497,N_12341,N_13329);
and U17498 (N_17498,N_14935,N_14080);
and U17499 (N_17499,N_13890,N_12900);
nand U17500 (N_17500,N_13703,N_11410);
and U17501 (N_17501,N_14000,N_13346);
nor U17502 (N_17502,N_12400,N_14872);
and U17503 (N_17503,N_12044,N_10294);
or U17504 (N_17504,N_10187,N_11827);
nand U17505 (N_17505,N_12757,N_10295);
nor U17506 (N_17506,N_12375,N_10551);
nand U17507 (N_17507,N_14751,N_12929);
nor U17508 (N_17508,N_12319,N_11613);
nand U17509 (N_17509,N_13739,N_12193);
nand U17510 (N_17510,N_14730,N_12181);
or U17511 (N_17511,N_12756,N_11507);
and U17512 (N_17512,N_14345,N_13389);
nand U17513 (N_17513,N_10757,N_13018);
or U17514 (N_17514,N_10693,N_12270);
and U17515 (N_17515,N_10654,N_13277);
or U17516 (N_17516,N_11810,N_12920);
and U17517 (N_17517,N_11910,N_10775);
or U17518 (N_17518,N_10503,N_12038);
nand U17519 (N_17519,N_14683,N_10897);
and U17520 (N_17520,N_14407,N_10449);
and U17521 (N_17521,N_13062,N_11991);
or U17522 (N_17522,N_10091,N_14193);
or U17523 (N_17523,N_14194,N_13189);
nor U17524 (N_17524,N_12052,N_12075);
or U17525 (N_17525,N_11870,N_10855);
nor U17526 (N_17526,N_14550,N_11247);
and U17527 (N_17527,N_11236,N_14706);
xor U17528 (N_17528,N_11357,N_14327);
and U17529 (N_17529,N_11184,N_11879);
nor U17530 (N_17530,N_10591,N_14055);
nand U17531 (N_17531,N_12777,N_14217);
and U17532 (N_17532,N_12437,N_12136);
nor U17533 (N_17533,N_10857,N_11096);
or U17534 (N_17534,N_10930,N_11941);
or U17535 (N_17535,N_13023,N_11987);
nor U17536 (N_17536,N_14175,N_10008);
or U17537 (N_17537,N_13627,N_10055);
nor U17538 (N_17538,N_12064,N_13544);
nor U17539 (N_17539,N_11882,N_10070);
nand U17540 (N_17540,N_12218,N_13741);
and U17541 (N_17541,N_10438,N_13091);
and U17542 (N_17542,N_13282,N_13962);
or U17543 (N_17543,N_11680,N_13929);
nor U17544 (N_17544,N_12854,N_11559);
and U17545 (N_17545,N_14588,N_13315);
nand U17546 (N_17546,N_10864,N_14522);
and U17547 (N_17547,N_14105,N_13088);
or U17548 (N_17548,N_14962,N_14563);
or U17549 (N_17549,N_13131,N_10978);
nand U17550 (N_17550,N_10504,N_10758);
nand U17551 (N_17551,N_12012,N_10122);
and U17552 (N_17552,N_12954,N_11451);
nand U17553 (N_17553,N_12514,N_11875);
and U17554 (N_17554,N_10348,N_10113);
nand U17555 (N_17555,N_12007,N_14822);
and U17556 (N_17556,N_10899,N_12745);
and U17557 (N_17557,N_13133,N_11947);
and U17558 (N_17558,N_14639,N_12995);
or U17559 (N_17559,N_12260,N_10501);
or U17560 (N_17560,N_14407,N_13820);
or U17561 (N_17561,N_10807,N_12997);
nand U17562 (N_17562,N_14979,N_13223);
nand U17563 (N_17563,N_12463,N_13430);
and U17564 (N_17564,N_12147,N_12277);
nor U17565 (N_17565,N_14940,N_13731);
nand U17566 (N_17566,N_10669,N_11603);
and U17567 (N_17567,N_12638,N_14614);
and U17568 (N_17568,N_12538,N_12554);
nand U17569 (N_17569,N_10136,N_11612);
nand U17570 (N_17570,N_12965,N_12343);
or U17571 (N_17571,N_13524,N_13519);
or U17572 (N_17572,N_11317,N_12346);
and U17573 (N_17573,N_11424,N_12090);
or U17574 (N_17574,N_11885,N_12531);
nor U17575 (N_17575,N_13956,N_14586);
nor U17576 (N_17576,N_14558,N_12392);
nor U17577 (N_17577,N_12949,N_10064);
nand U17578 (N_17578,N_12152,N_14530);
or U17579 (N_17579,N_12041,N_13423);
or U17580 (N_17580,N_12085,N_14080);
or U17581 (N_17581,N_10226,N_12647);
and U17582 (N_17582,N_13799,N_12476);
nand U17583 (N_17583,N_12149,N_13982);
nor U17584 (N_17584,N_11720,N_14305);
nor U17585 (N_17585,N_14816,N_11078);
nand U17586 (N_17586,N_14513,N_10943);
nand U17587 (N_17587,N_10061,N_14177);
or U17588 (N_17588,N_12280,N_13624);
nand U17589 (N_17589,N_10052,N_14926);
xnor U17590 (N_17590,N_13864,N_14427);
nand U17591 (N_17591,N_12903,N_11746);
and U17592 (N_17592,N_10683,N_12944);
nor U17593 (N_17593,N_14637,N_14922);
nor U17594 (N_17594,N_14880,N_11267);
nand U17595 (N_17595,N_14521,N_12880);
nor U17596 (N_17596,N_10239,N_12196);
nand U17597 (N_17597,N_12557,N_11274);
nor U17598 (N_17598,N_12498,N_14527);
nand U17599 (N_17599,N_12710,N_13297);
or U17600 (N_17600,N_12947,N_11190);
xnor U17601 (N_17601,N_12658,N_10898);
or U17602 (N_17602,N_11864,N_10795);
nor U17603 (N_17603,N_10950,N_10289);
nor U17604 (N_17604,N_14176,N_13238);
or U17605 (N_17605,N_11027,N_12126);
nand U17606 (N_17606,N_14089,N_11587);
nor U17607 (N_17607,N_13218,N_13581);
xnor U17608 (N_17608,N_11317,N_13435);
and U17609 (N_17609,N_14327,N_14363);
nor U17610 (N_17610,N_12633,N_12877);
or U17611 (N_17611,N_13111,N_11160);
nor U17612 (N_17612,N_13250,N_12388);
and U17613 (N_17613,N_11281,N_14576);
nor U17614 (N_17614,N_12242,N_10053);
nand U17615 (N_17615,N_14941,N_12867);
xor U17616 (N_17616,N_13716,N_13837);
nand U17617 (N_17617,N_13436,N_14023);
nand U17618 (N_17618,N_14024,N_11585);
nand U17619 (N_17619,N_10773,N_13607);
or U17620 (N_17620,N_12566,N_12958);
and U17621 (N_17621,N_12325,N_14883);
or U17622 (N_17622,N_10982,N_14626);
xor U17623 (N_17623,N_10512,N_12477);
or U17624 (N_17624,N_12096,N_10122);
nor U17625 (N_17625,N_14641,N_10264);
nor U17626 (N_17626,N_12099,N_13959);
nor U17627 (N_17627,N_13347,N_13100);
nand U17628 (N_17628,N_12015,N_13041);
or U17629 (N_17629,N_11862,N_12585);
or U17630 (N_17630,N_14145,N_10143);
and U17631 (N_17631,N_14571,N_10816);
nand U17632 (N_17632,N_10460,N_14230);
nand U17633 (N_17633,N_10216,N_13472);
nor U17634 (N_17634,N_10159,N_11045);
or U17635 (N_17635,N_13123,N_10196);
and U17636 (N_17636,N_12841,N_13270);
and U17637 (N_17637,N_12316,N_14264);
nand U17638 (N_17638,N_12504,N_11982);
or U17639 (N_17639,N_14777,N_10672);
and U17640 (N_17640,N_12803,N_11535);
or U17641 (N_17641,N_10679,N_12243);
or U17642 (N_17642,N_13163,N_12187);
nor U17643 (N_17643,N_11974,N_13320);
and U17644 (N_17644,N_12993,N_10630);
or U17645 (N_17645,N_11059,N_13353);
nand U17646 (N_17646,N_14930,N_11381);
or U17647 (N_17647,N_12679,N_14343);
nand U17648 (N_17648,N_13265,N_12776);
or U17649 (N_17649,N_10612,N_13001);
xor U17650 (N_17650,N_11221,N_11368);
nand U17651 (N_17651,N_12424,N_13267);
nand U17652 (N_17652,N_12045,N_12697);
nor U17653 (N_17653,N_14939,N_11393);
and U17654 (N_17654,N_13745,N_10608);
and U17655 (N_17655,N_12152,N_13122);
nor U17656 (N_17656,N_10407,N_12641);
nor U17657 (N_17657,N_12371,N_14716);
or U17658 (N_17658,N_12204,N_14207);
nor U17659 (N_17659,N_10937,N_10496);
nor U17660 (N_17660,N_14867,N_10326);
and U17661 (N_17661,N_11475,N_14410);
and U17662 (N_17662,N_14083,N_13205);
nand U17663 (N_17663,N_11654,N_11496);
and U17664 (N_17664,N_12855,N_13068);
nor U17665 (N_17665,N_14598,N_13436);
xor U17666 (N_17666,N_13526,N_12390);
nand U17667 (N_17667,N_11871,N_13717);
nand U17668 (N_17668,N_13096,N_11442);
nor U17669 (N_17669,N_10902,N_11171);
and U17670 (N_17670,N_12610,N_12456);
nor U17671 (N_17671,N_10348,N_10218);
nor U17672 (N_17672,N_14772,N_11342);
and U17673 (N_17673,N_14266,N_12945);
and U17674 (N_17674,N_12856,N_10655);
or U17675 (N_17675,N_12303,N_11623);
nor U17676 (N_17676,N_12503,N_11726);
nor U17677 (N_17677,N_14065,N_11672);
nand U17678 (N_17678,N_13993,N_12692);
nor U17679 (N_17679,N_12496,N_11460);
and U17680 (N_17680,N_11334,N_12541);
nor U17681 (N_17681,N_11419,N_14097);
or U17682 (N_17682,N_13508,N_10516);
or U17683 (N_17683,N_12738,N_14583);
nor U17684 (N_17684,N_10972,N_12351);
nand U17685 (N_17685,N_10919,N_12408);
nand U17686 (N_17686,N_13907,N_12289);
nand U17687 (N_17687,N_10597,N_10778);
nand U17688 (N_17688,N_11564,N_10119);
and U17689 (N_17689,N_12145,N_14385);
nand U17690 (N_17690,N_11748,N_12967);
and U17691 (N_17691,N_13979,N_11465);
or U17692 (N_17692,N_14342,N_13846);
and U17693 (N_17693,N_10630,N_13483);
nor U17694 (N_17694,N_11037,N_12841);
nand U17695 (N_17695,N_13614,N_10657);
nand U17696 (N_17696,N_12650,N_13449);
and U17697 (N_17697,N_13407,N_12295);
and U17698 (N_17698,N_10331,N_10994);
nand U17699 (N_17699,N_14892,N_11214);
nor U17700 (N_17700,N_10811,N_13662);
and U17701 (N_17701,N_13572,N_12322);
nor U17702 (N_17702,N_14746,N_13935);
or U17703 (N_17703,N_11530,N_13714);
nor U17704 (N_17704,N_10501,N_11698);
and U17705 (N_17705,N_14312,N_13390);
nand U17706 (N_17706,N_14005,N_12703);
nand U17707 (N_17707,N_11500,N_14503);
nand U17708 (N_17708,N_14471,N_14032);
nand U17709 (N_17709,N_12431,N_14761);
or U17710 (N_17710,N_13661,N_14814);
and U17711 (N_17711,N_13300,N_13569);
or U17712 (N_17712,N_10803,N_13862);
nor U17713 (N_17713,N_14503,N_11508);
nor U17714 (N_17714,N_14441,N_12964);
nor U17715 (N_17715,N_10441,N_12278);
or U17716 (N_17716,N_11774,N_12626);
xnor U17717 (N_17717,N_11912,N_10380);
nand U17718 (N_17718,N_14505,N_10432);
and U17719 (N_17719,N_11848,N_11771);
nor U17720 (N_17720,N_12731,N_13326);
and U17721 (N_17721,N_14207,N_13876);
and U17722 (N_17722,N_11592,N_13691);
and U17723 (N_17723,N_10750,N_11561);
and U17724 (N_17724,N_13224,N_14618);
and U17725 (N_17725,N_12393,N_14279);
or U17726 (N_17726,N_13569,N_14357);
nor U17727 (N_17727,N_14754,N_14712);
nor U17728 (N_17728,N_11144,N_14540);
nand U17729 (N_17729,N_11153,N_13684);
nand U17730 (N_17730,N_14971,N_10565);
nand U17731 (N_17731,N_10922,N_11384);
or U17732 (N_17732,N_10489,N_13912);
nor U17733 (N_17733,N_11770,N_12952);
or U17734 (N_17734,N_14610,N_14517);
nand U17735 (N_17735,N_11203,N_11589);
nand U17736 (N_17736,N_14307,N_10487);
nand U17737 (N_17737,N_13573,N_14012);
nor U17738 (N_17738,N_10683,N_12384);
nor U17739 (N_17739,N_12470,N_12313);
and U17740 (N_17740,N_11597,N_11571);
nand U17741 (N_17741,N_11424,N_11887);
and U17742 (N_17742,N_14769,N_12555);
and U17743 (N_17743,N_13969,N_13957);
or U17744 (N_17744,N_14659,N_14697);
nor U17745 (N_17745,N_10317,N_13257);
or U17746 (N_17746,N_14069,N_10363);
and U17747 (N_17747,N_10524,N_12629);
nor U17748 (N_17748,N_10958,N_13127);
xor U17749 (N_17749,N_11345,N_11969);
nor U17750 (N_17750,N_14123,N_12701);
or U17751 (N_17751,N_13997,N_11783);
and U17752 (N_17752,N_14167,N_13730);
nor U17753 (N_17753,N_12037,N_12872);
or U17754 (N_17754,N_14263,N_12578);
or U17755 (N_17755,N_14261,N_13194);
nor U17756 (N_17756,N_11192,N_13691);
nand U17757 (N_17757,N_12237,N_13320);
nor U17758 (N_17758,N_13897,N_14847);
nand U17759 (N_17759,N_11387,N_13851);
or U17760 (N_17760,N_12715,N_13324);
nor U17761 (N_17761,N_10416,N_10177);
or U17762 (N_17762,N_12838,N_10144);
nand U17763 (N_17763,N_12354,N_13081);
or U17764 (N_17764,N_11658,N_14820);
nor U17765 (N_17765,N_14755,N_14021);
or U17766 (N_17766,N_10254,N_14455);
nand U17767 (N_17767,N_14203,N_10594);
and U17768 (N_17768,N_11988,N_14312);
nor U17769 (N_17769,N_13000,N_10617);
nand U17770 (N_17770,N_11448,N_14720);
nor U17771 (N_17771,N_12083,N_13622);
or U17772 (N_17772,N_12474,N_14937);
nor U17773 (N_17773,N_10362,N_13307);
nor U17774 (N_17774,N_12503,N_11632);
xnor U17775 (N_17775,N_12849,N_14536);
nand U17776 (N_17776,N_10037,N_10288);
and U17777 (N_17777,N_13897,N_13472);
nor U17778 (N_17778,N_14790,N_11074);
and U17779 (N_17779,N_13919,N_11207);
nor U17780 (N_17780,N_12915,N_12295);
and U17781 (N_17781,N_10990,N_12217);
nor U17782 (N_17782,N_10373,N_10752);
nand U17783 (N_17783,N_14421,N_12468);
or U17784 (N_17784,N_13349,N_10853);
nand U17785 (N_17785,N_13539,N_10718);
xnor U17786 (N_17786,N_13388,N_10874);
or U17787 (N_17787,N_13432,N_10793);
or U17788 (N_17788,N_12116,N_13396);
and U17789 (N_17789,N_13455,N_11344);
and U17790 (N_17790,N_13485,N_11998);
nor U17791 (N_17791,N_13807,N_13084);
nor U17792 (N_17792,N_14620,N_13465);
nor U17793 (N_17793,N_13547,N_11045);
and U17794 (N_17794,N_14355,N_11850);
nor U17795 (N_17795,N_11346,N_13279);
and U17796 (N_17796,N_12609,N_10054);
nand U17797 (N_17797,N_13554,N_13645);
nor U17798 (N_17798,N_12449,N_13568);
or U17799 (N_17799,N_13140,N_14440);
nand U17800 (N_17800,N_11935,N_12027);
nor U17801 (N_17801,N_10443,N_10584);
and U17802 (N_17802,N_13975,N_14776);
and U17803 (N_17803,N_11470,N_13179);
or U17804 (N_17804,N_11779,N_13215);
nor U17805 (N_17805,N_11779,N_12107);
or U17806 (N_17806,N_13359,N_14577);
nand U17807 (N_17807,N_12241,N_10201);
and U17808 (N_17808,N_11995,N_13190);
or U17809 (N_17809,N_12649,N_14324);
or U17810 (N_17810,N_10592,N_10328);
nor U17811 (N_17811,N_13432,N_13712);
or U17812 (N_17812,N_13664,N_10829);
and U17813 (N_17813,N_14580,N_13605);
and U17814 (N_17814,N_13308,N_12951);
and U17815 (N_17815,N_10290,N_11517);
or U17816 (N_17816,N_12225,N_13416);
nor U17817 (N_17817,N_13803,N_14101);
and U17818 (N_17818,N_14295,N_12326);
nand U17819 (N_17819,N_10129,N_13060);
xor U17820 (N_17820,N_10732,N_12535);
or U17821 (N_17821,N_11850,N_12844);
or U17822 (N_17822,N_14551,N_14304);
nor U17823 (N_17823,N_12193,N_13204);
and U17824 (N_17824,N_11681,N_11731);
and U17825 (N_17825,N_12588,N_10962);
or U17826 (N_17826,N_12376,N_14376);
or U17827 (N_17827,N_14571,N_11475);
xor U17828 (N_17828,N_12646,N_12794);
nor U17829 (N_17829,N_10251,N_14258);
nand U17830 (N_17830,N_10325,N_10163);
nor U17831 (N_17831,N_10936,N_14843);
nand U17832 (N_17832,N_10396,N_14577);
nor U17833 (N_17833,N_12921,N_14493);
or U17834 (N_17834,N_11097,N_11945);
or U17835 (N_17835,N_10098,N_13243);
and U17836 (N_17836,N_11338,N_13800);
nand U17837 (N_17837,N_10009,N_13000);
xor U17838 (N_17838,N_12788,N_14127);
nand U17839 (N_17839,N_11138,N_11871);
and U17840 (N_17840,N_11695,N_10500);
and U17841 (N_17841,N_13714,N_12842);
or U17842 (N_17842,N_12640,N_12590);
or U17843 (N_17843,N_11797,N_11567);
or U17844 (N_17844,N_12154,N_14348);
nor U17845 (N_17845,N_14376,N_11946);
nand U17846 (N_17846,N_10995,N_10057);
or U17847 (N_17847,N_14890,N_10734);
and U17848 (N_17848,N_11668,N_13522);
and U17849 (N_17849,N_11417,N_12177);
nand U17850 (N_17850,N_12671,N_11428);
xor U17851 (N_17851,N_13304,N_13313);
nor U17852 (N_17852,N_11593,N_10883);
nand U17853 (N_17853,N_11105,N_12918);
nor U17854 (N_17854,N_11393,N_11146);
nand U17855 (N_17855,N_13806,N_12140);
nor U17856 (N_17856,N_11206,N_14536);
and U17857 (N_17857,N_10693,N_12826);
nand U17858 (N_17858,N_10509,N_12723);
nand U17859 (N_17859,N_11953,N_13770);
or U17860 (N_17860,N_13816,N_12323);
or U17861 (N_17861,N_14482,N_14650);
xnor U17862 (N_17862,N_11996,N_14863);
or U17863 (N_17863,N_11131,N_13775);
and U17864 (N_17864,N_10955,N_14885);
nand U17865 (N_17865,N_13111,N_12735);
and U17866 (N_17866,N_14835,N_11836);
or U17867 (N_17867,N_10601,N_14875);
nor U17868 (N_17868,N_14362,N_12280);
and U17869 (N_17869,N_11610,N_14848);
or U17870 (N_17870,N_11077,N_11885);
nand U17871 (N_17871,N_11673,N_13696);
or U17872 (N_17872,N_12581,N_14326);
or U17873 (N_17873,N_13338,N_14149);
or U17874 (N_17874,N_13008,N_10613);
and U17875 (N_17875,N_13997,N_10563);
or U17876 (N_17876,N_13708,N_13201);
nor U17877 (N_17877,N_14019,N_12688);
or U17878 (N_17878,N_13435,N_11150);
nand U17879 (N_17879,N_14719,N_14866);
and U17880 (N_17880,N_11776,N_14638);
or U17881 (N_17881,N_13559,N_12209);
and U17882 (N_17882,N_11381,N_11667);
or U17883 (N_17883,N_12493,N_11468);
and U17884 (N_17884,N_11113,N_12172);
or U17885 (N_17885,N_11251,N_12627);
nand U17886 (N_17886,N_10012,N_12578);
or U17887 (N_17887,N_11578,N_12055);
nand U17888 (N_17888,N_13680,N_12820);
nor U17889 (N_17889,N_14937,N_10180);
nor U17890 (N_17890,N_10278,N_10668);
nor U17891 (N_17891,N_14750,N_13403);
nand U17892 (N_17892,N_11514,N_13175);
nand U17893 (N_17893,N_12757,N_13710);
or U17894 (N_17894,N_14572,N_14347);
and U17895 (N_17895,N_13602,N_11940);
nand U17896 (N_17896,N_13920,N_11678);
and U17897 (N_17897,N_12575,N_10493);
nor U17898 (N_17898,N_14041,N_11078);
or U17899 (N_17899,N_13976,N_11225);
nand U17900 (N_17900,N_12866,N_14162);
and U17901 (N_17901,N_14225,N_11017);
nand U17902 (N_17902,N_11452,N_11539);
nand U17903 (N_17903,N_13599,N_14373);
nor U17904 (N_17904,N_13389,N_14945);
nor U17905 (N_17905,N_10187,N_11764);
nor U17906 (N_17906,N_12351,N_12129);
xnor U17907 (N_17907,N_12630,N_11883);
nand U17908 (N_17908,N_11236,N_10724);
nor U17909 (N_17909,N_13679,N_12608);
or U17910 (N_17910,N_13905,N_11128);
nand U17911 (N_17911,N_11537,N_12818);
nand U17912 (N_17912,N_12513,N_14157);
and U17913 (N_17913,N_14220,N_10141);
nand U17914 (N_17914,N_11492,N_14323);
nor U17915 (N_17915,N_13236,N_10130);
nand U17916 (N_17916,N_11508,N_13045);
nor U17917 (N_17917,N_10145,N_14676);
nor U17918 (N_17918,N_11353,N_14683);
and U17919 (N_17919,N_14574,N_11794);
nor U17920 (N_17920,N_12563,N_11868);
nor U17921 (N_17921,N_13004,N_12157);
and U17922 (N_17922,N_10596,N_12551);
and U17923 (N_17923,N_14194,N_12863);
or U17924 (N_17924,N_13666,N_14500);
or U17925 (N_17925,N_14674,N_12506);
and U17926 (N_17926,N_11711,N_13480);
xnor U17927 (N_17927,N_11077,N_10073);
xor U17928 (N_17928,N_13335,N_13232);
nand U17929 (N_17929,N_13741,N_13860);
nor U17930 (N_17930,N_12857,N_10849);
or U17931 (N_17931,N_12504,N_14396);
and U17932 (N_17932,N_10483,N_11419);
nand U17933 (N_17933,N_12937,N_11767);
or U17934 (N_17934,N_14340,N_11027);
or U17935 (N_17935,N_14780,N_13097);
nand U17936 (N_17936,N_10978,N_10847);
nand U17937 (N_17937,N_14054,N_10548);
nor U17938 (N_17938,N_12614,N_12478);
nand U17939 (N_17939,N_14584,N_10858);
nor U17940 (N_17940,N_11414,N_14619);
and U17941 (N_17941,N_10294,N_13004);
and U17942 (N_17942,N_11370,N_12283);
and U17943 (N_17943,N_13925,N_11084);
xor U17944 (N_17944,N_10106,N_12773);
or U17945 (N_17945,N_10740,N_10587);
nand U17946 (N_17946,N_13568,N_13536);
nor U17947 (N_17947,N_10735,N_10284);
nand U17948 (N_17948,N_12496,N_10658);
nor U17949 (N_17949,N_13937,N_14200);
or U17950 (N_17950,N_13672,N_12785);
nor U17951 (N_17951,N_11445,N_13522);
and U17952 (N_17952,N_13400,N_12215);
and U17953 (N_17953,N_11543,N_13010);
or U17954 (N_17954,N_12436,N_10299);
nand U17955 (N_17955,N_10963,N_11021);
or U17956 (N_17956,N_12388,N_11249);
and U17957 (N_17957,N_14764,N_10222);
nand U17958 (N_17958,N_12613,N_10166);
or U17959 (N_17959,N_11639,N_14674);
or U17960 (N_17960,N_10288,N_10668);
or U17961 (N_17961,N_10434,N_12251);
nor U17962 (N_17962,N_11674,N_12181);
nor U17963 (N_17963,N_13928,N_14407);
or U17964 (N_17964,N_10743,N_14731);
or U17965 (N_17965,N_11022,N_10598);
and U17966 (N_17966,N_14366,N_13963);
and U17967 (N_17967,N_12253,N_13689);
or U17968 (N_17968,N_13795,N_12006);
and U17969 (N_17969,N_10780,N_10173);
nand U17970 (N_17970,N_13086,N_11539);
nand U17971 (N_17971,N_10722,N_14076);
nand U17972 (N_17972,N_14030,N_10049);
nor U17973 (N_17973,N_11511,N_12285);
or U17974 (N_17974,N_11193,N_13600);
and U17975 (N_17975,N_14165,N_10355);
nor U17976 (N_17976,N_11608,N_13802);
nand U17977 (N_17977,N_12534,N_12806);
or U17978 (N_17978,N_10740,N_11262);
nand U17979 (N_17979,N_11585,N_13831);
nand U17980 (N_17980,N_11101,N_10093);
nor U17981 (N_17981,N_10825,N_11103);
or U17982 (N_17982,N_14346,N_14561);
nand U17983 (N_17983,N_10488,N_11750);
and U17984 (N_17984,N_12654,N_11551);
nand U17985 (N_17985,N_10593,N_12319);
or U17986 (N_17986,N_10344,N_12218);
and U17987 (N_17987,N_10954,N_10793);
or U17988 (N_17988,N_12958,N_12501);
and U17989 (N_17989,N_11648,N_11728);
nor U17990 (N_17990,N_13996,N_11320);
and U17991 (N_17991,N_11344,N_12979);
nand U17992 (N_17992,N_13626,N_10194);
or U17993 (N_17993,N_13682,N_14423);
nand U17994 (N_17994,N_13502,N_13444);
or U17995 (N_17995,N_12565,N_10941);
and U17996 (N_17996,N_11156,N_13966);
and U17997 (N_17997,N_12414,N_10680);
or U17998 (N_17998,N_13342,N_12821);
nor U17999 (N_17999,N_10881,N_14039);
xor U18000 (N_18000,N_14357,N_12425);
and U18001 (N_18001,N_13925,N_12837);
nor U18002 (N_18002,N_12477,N_14290);
or U18003 (N_18003,N_14387,N_13873);
nand U18004 (N_18004,N_11654,N_12303);
nand U18005 (N_18005,N_13947,N_11973);
nor U18006 (N_18006,N_11194,N_12826);
or U18007 (N_18007,N_13500,N_11403);
nand U18008 (N_18008,N_12691,N_10305);
or U18009 (N_18009,N_12876,N_14787);
nand U18010 (N_18010,N_12148,N_10087);
and U18011 (N_18011,N_13425,N_13445);
nand U18012 (N_18012,N_10475,N_14843);
nand U18013 (N_18013,N_10051,N_13406);
nor U18014 (N_18014,N_13689,N_11292);
nor U18015 (N_18015,N_10709,N_14759);
or U18016 (N_18016,N_12938,N_14984);
and U18017 (N_18017,N_10484,N_11863);
nor U18018 (N_18018,N_13678,N_14344);
and U18019 (N_18019,N_12149,N_14463);
nor U18020 (N_18020,N_13251,N_12640);
nand U18021 (N_18021,N_13287,N_10536);
and U18022 (N_18022,N_14640,N_12204);
or U18023 (N_18023,N_10545,N_14308);
nor U18024 (N_18024,N_12516,N_12032);
nand U18025 (N_18025,N_11327,N_13008);
or U18026 (N_18026,N_11338,N_13135);
nand U18027 (N_18027,N_12898,N_10205);
or U18028 (N_18028,N_14269,N_10039);
nand U18029 (N_18029,N_14626,N_13604);
nand U18030 (N_18030,N_13424,N_10138);
and U18031 (N_18031,N_12963,N_10671);
and U18032 (N_18032,N_10374,N_13487);
nand U18033 (N_18033,N_13160,N_13351);
nand U18034 (N_18034,N_14474,N_10607);
nor U18035 (N_18035,N_12202,N_10377);
nor U18036 (N_18036,N_11576,N_14031);
or U18037 (N_18037,N_13650,N_12910);
nor U18038 (N_18038,N_12959,N_10263);
nand U18039 (N_18039,N_12339,N_13940);
nand U18040 (N_18040,N_11160,N_14123);
nor U18041 (N_18041,N_11770,N_11358);
nand U18042 (N_18042,N_13800,N_14500);
and U18043 (N_18043,N_10202,N_10222);
nor U18044 (N_18044,N_10931,N_11677);
and U18045 (N_18045,N_10174,N_11421);
and U18046 (N_18046,N_14834,N_10230);
or U18047 (N_18047,N_13682,N_10217);
and U18048 (N_18048,N_13779,N_12656);
or U18049 (N_18049,N_10472,N_10413);
nand U18050 (N_18050,N_14566,N_11413);
nor U18051 (N_18051,N_12340,N_10316);
and U18052 (N_18052,N_13284,N_14109);
or U18053 (N_18053,N_11264,N_12764);
and U18054 (N_18054,N_14115,N_10013);
nor U18055 (N_18055,N_10329,N_11886);
and U18056 (N_18056,N_12027,N_12162);
nand U18057 (N_18057,N_12131,N_11067);
and U18058 (N_18058,N_11230,N_14637);
nor U18059 (N_18059,N_12817,N_13886);
or U18060 (N_18060,N_11783,N_13543);
nand U18061 (N_18061,N_13361,N_12837);
and U18062 (N_18062,N_12323,N_12204);
or U18063 (N_18063,N_11290,N_14307);
nand U18064 (N_18064,N_12919,N_11788);
and U18065 (N_18065,N_11870,N_14825);
nor U18066 (N_18066,N_13331,N_11256);
nor U18067 (N_18067,N_12840,N_13350);
and U18068 (N_18068,N_14983,N_13217);
nor U18069 (N_18069,N_10316,N_11341);
and U18070 (N_18070,N_12422,N_13872);
nor U18071 (N_18071,N_12986,N_11074);
nor U18072 (N_18072,N_12957,N_13422);
nand U18073 (N_18073,N_12019,N_11591);
nand U18074 (N_18074,N_12545,N_10738);
xnor U18075 (N_18075,N_12790,N_10649);
nand U18076 (N_18076,N_11709,N_11727);
or U18077 (N_18077,N_13437,N_14209);
and U18078 (N_18078,N_11086,N_12857);
or U18079 (N_18079,N_14697,N_11606);
nor U18080 (N_18080,N_13035,N_10134);
nor U18081 (N_18081,N_13301,N_13601);
nand U18082 (N_18082,N_11357,N_12190);
or U18083 (N_18083,N_11463,N_11330);
nor U18084 (N_18084,N_14987,N_12243);
nor U18085 (N_18085,N_14703,N_13450);
or U18086 (N_18086,N_12266,N_11529);
and U18087 (N_18087,N_13128,N_13489);
or U18088 (N_18088,N_14311,N_11287);
and U18089 (N_18089,N_10422,N_11410);
and U18090 (N_18090,N_10163,N_12572);
or U18091 (N_18091,N_10994,N_13654);
nand U18092 (N_18092,N_14827,N_13913);
nor U18093 (N_18093,N_13577,N_14549);
and U18094 (N_18094,N_12889,N_14853);
nand U18095 (N_18095,N_13423,N_13637);
and U18096 (N_18096,N_13700,N_10502);
or U18097 (N_18097,N_13522,N_11591);
nand U18098 (N_18098,N_11328,N_10745);
and U18099 (N_18099,N_13284,N_10380);
and U18100 (N_18100,N_10852,N_13224);
or U18101 (N_18101,N_10148,N_10600);
nand U18102 (N_18102,N_10890,N_11410);
or U18103 (N_18103,N_10197,N_11257);
and U18104 (N_18104,N_11575,N_12128);
nor U18105 (N_18105,N_14356,N_14774);
and U18106 (N_18106,N_10342,N_10629);
and U18107 (N_18107,N_11457,N_10230);
xnor U18108 (N_18108,N_14655,N_13877);
nand U18109 (N_18109,N_11774,N_13936);
or U18110 (N_18110,N_11480,N_14103);
or U18111 (N_18111,N_14153,N_14801);
and U18112 (N_18112,N_11362,N_13999);
nor U18113 (N_18113,N_14366,N_12397);
nor U18114 (N_18114,N_11723,N_12527);
nand U18115 (N_18115,N_10077,N_10464);
or U18116 (N_18116,N_10568,N_11563);
nor U18117 (N_18117,N_10186,N_11862);
nand U18118 (N_18118,N_11189,N_13495);
nand U18119 (N_18119,N_14500,N_10177);
and U18120 (N_18120,N_10844,N_12849);
nand U18121 (N_18121,N_11797,N_13868);
nor U18122 (N_18122,N_11470,N_14836);
and U18123 (N_18123,N_11039,N_12102);
nor U18124 (N_18124,N_10808,N_13514);
or U18125 (N_18125,N_11578,N_11094);
nor U18126 (N_18126,N_12080,N_13380);
nor U18127 (N_18127,N_10008,N_13245);
nand U18128 (N_18128,N_14673,N_10735);
nor U18129 (N_18129,N_12205,N_14008);
and U18130 (N_18130,N_10287,N_14731);
nand U18131 (N_18131,N_10638,N_14615);
nor U18132 (N_18132,N_13954,N_11146);
nor U18133 (N_18133,N_12345,N_12137);
and U18134 (N_18134,N_12741,N_12131);
nand U18135 (N_18135,N_10106,N_10437);
xor U18136 (N_18136,N_13465,N_14833);
and U18137 (N_18137,N_13490,N_13730);
or U18138 (N_18138,N_12290,N_10800);
nand U18139 (N_18139,N_11760,N_12992);
nand U18140 (N_18140,N_10280,N_12022);
xnor U18141 (N_18141,N_13919,N_14533);
or U18142 (N_18142,N_13274,N_11229);
nand U18143 (N_18143,N_14621,N_11442);
nor U18144 (N_18144,N_11070,N_10431);
nand U18145 (N_18145,N_11265,N_12666);
and U18146 (N_18146,N_14711,N_13267);
and U18147 (N_18147,N_13524,N_11380);
or U18148 (N_18148,N_12237,N_10355);
nor U18149 (N_18149,N_13130,N_14631);
nor U18150 (N_18150,N_12688,N_14359);
or U18151 (N_18151,N_12298,N_13796);
nor U18152 (N_18152,N_12062,N_10593);
and U18153 (N_18153,N_14368,N_11536);
or U18154 (N_18154,N_13868,N_12122);
nand U18155 (N_18155,N_14896,N_13336);
xor U18156 (N_18156,N_11641,N_10695);
nand U18157 (N_18157,N_14710,N_10820);
and U18158 (N_18158,N_12535,N_11037);
or U18159 (N_18159,N_12251,N_14502);
and U18160 (N_18160,N_14402,N_12518);
and U18161 (N_18161,N_12213,N_11042);
and U18162 (N_18162,N_13921,N_14788);
and U18163 (N_18163,N_10324,N_11705);
nor U18164 (N_18164,N_13668,N_13988);
nor U18165 (N_18165,N_10911,N_12398);
xor U18166 (N_18166,N_14575,N_10646);
and U18167 (N_18167,N_13068,N_13747);
or U18168 (N_18168,N_14597,N_12348);
or U18169 (N_18169,N_11460,N_12102);
or U18170 (N_18170,N_10182,N_14273);
or U18171 (N_18171,N_10243,N_13087);
nand U18172 (N_18172,N_12061,N_10471);
nor U18173 (N_18173,N_14471,N_13879);
nor U18174 (N_18174,N_13790,N_11366);
and U18175 (N_18175,N_14893,N_11380);
or U18176 (N_18176,N_13799,N_11067);
nor U18177 (N_18177,N_12114,N_10730);
or U18178 (N_18178,N_12636,N_13263);
and U18179 (N_18179,N_11993,N_12699);
and U18180 (N_18180,N_11975,N_11355);
nand U18181 (N_18181,N_14936,N_12760);
and U18182 (N_18182,N_13143,N_10043);
and U18183 (N_18183,N_13942,N_12073);
nor U18184 (N_18184,N_14232,N_11884);
or U18185 (N_18185,N_13256,N_12457);
or U18186 (N_18186,N_11149,N_10199);
nor U18187 (N_18187,N_13403,N_12042);
or U18188 (N_18188,N_12549,N_14635);
or U18189 (N_18189,N_10843,N_12552);
nor U18190 (N_18190,N_13948,N_10145);
or U18191 (N_18191,N_14661,N_12858);
and U18192 (N_18192,N_13671,N_13148);
nor U18193 (N_18193,N_10095,N_13180);
and U18194 (N_18194,N_13372,N_10185);
or U18195 (N_18195,N_14348,N_13185);
or U18196 (N_18196,N_13601,N_10670);
nor U18197 (N_18197,N_14055,N_14488);
nand U18198 (N_18198,N_11590,N_14810);
or U18199 (N_18199,N_14619,N_11650);
or U18200 (N_18200,N_14291,N_11665);
nor U18201 (N_18201,N_11862,N_12367);
or U18202 (N_18202,N_13623,N_12223);
nand U18203 (N_18203,N_11817,N_11929);
or U18204 (N_18204,N_11965,N_14519);
nand U18205 (N_18205,N_11736,N_10267);
or U18206 (N_18206,N_12072,N_10828);
nor U18207 (N_18207,N_11461,N_11863);
or U18208 (N_18208,N_13641,N_12633);
nand U18209 (N_18209,N_11379,N_13644);
nor U18210 (N_18210,N_12206,N_14757);
and U18211 (N_18211,N_14356,N_14618);
or U18212 (N_18212,N_13475,N_14009);
or U18213 (N_18213,N_10168,N_14177);
and U18214 (N_18214,N_13022,N_12197);
nor U18215 (N_18215,N_12556,N_11998);
or U18216 (N_18216,N_10583,N_13750);
nor U18217 (N_18217,N_11341,N_11115);
and U18218 (N_18218,N_12402,N_11762);
and U18219 (N_18219,N_11609,N_13448);
nor U18220 (N_18220,N_12253,N_13638);
nor U18221 (N_18221,N_13471,N_13682);
nor U18222 (N_18222,N_12863,N_13799);
nor U18223 (N_18223,N_10338,N_11484);
or U18224 (N_18224,N_12420,N_14567);
nand U18225 (N_18225,N_12669,N_11542);
or U18226 (N_18226,N_11962,N_12320);
nand U18227 (N_18227,N_14707,N_10641);
or U18228 (N_18228,N_12632,N_13335);
or U18229 (N_18229,N_11500,N_11292);
nor U18230 (N_18230,N_10985,N_12481);
nor U18231 (N_18231,N_10231,N_14491);
and U18232 (N_18232,N_13243,N_11125);
or U18233 (N_18233,N_10990,N_11755);
nor U18234 (N_18234,N_13675,N_14932);
or U18235 (N_18235,N_13635,N_10723);
nor U18236 (N_18236,N_11069,N_13966);
or U18237 (N_18237,N_13630,N_10570);
nor U18238 (N_18238,N_11620,N_11164);
nand U18239 (N_18239,N_12018,N_14212);
and U18240 (N_18240,N_11078,N_11776);
or U18241 (N_18241,N_13845,N_13859);
nor U18242 (N_18242,N_14162,N_14259);
or U18243 (N_18243,N_10634,N_10949);
nand U18244 (N_18244,N_12840,N_14637);
or U18245 (N_18245,N_11630,N_10120);
or U18246 (N_18246,N_13381,N_12953);
or U18247 (N_18247,N_10189,N_10337);
and U18248 (N_18248,N_10786,N_12857);
nand U18249 (N_18249,N_11178,N_14602);
or U18250 (N_18250,N_11485,N_12413);
and U18251 (N_18251,N_11189,N_13662);
nor U18252 (N_18252,N_13848,N_10668);
nand U18253 (N_18253,N_10275,N_13481);
xor U18254 (N_18254,N_14551,N_14438);
or U18255 (N_18255,N_14766,N_13705);
or U18256 (N_18256,N_10776,N_13603);
nand U18257 (N_18257,N_11397,N_14287);
nor U18258 (N_18258,N_13836,N_11759);
xor U18259 (N_18259,N_11831,N_14787);
and U18260 (N_18260,N_13188,N_12371);
nand U18261 (N_18261,N_12791,N_12880);
nand U18262 (N_18262,N_11882,N_12526);
or U18263 (N_18263,N_12580,N_11873);
nand U18264 (N_18264,N_10758,N_14883);
nor U18265 (N_18265,N_14105,N_14585);
and U18266 (N_18266,N_12415,N_11931);
and U18267 (N_18267,N_10158,N_11002);
and U18268 (N_18268,N_14017,N_11518);
nand U18269 (N_18269,N_11473,N_11748);
and U18270 (N_18270,N_10090,N_11360);
nand U18271 (N_18271,N_12618,N_12776);
nor U18272 (N_18272,N_14578,N_11561);
nor U18273 (N_18273,N_10136,N_12088);
and U18274 (N_18274,N_11596,N_10820);
nor U18275 (N_18275,N_12615,N_14860);
or U18276 (N_18276,N_14524,N_14604);
and U18277 (N_18277,N_14136,N_10647);
xnor U18278 (N_18278,N_13199,N_11062);
and U18279 (N_18279,N_13414,N_12601);
nor U18280 (N_18280,N_11678,N_14782);
xnor U18281 (N_18281,N_13758,N_11664);
nor U18282 (N_18282,N_11603,N_13329);
nor U18283 (N_18283,N_11443,N_13165);
or U18284 (N_18284,N_14636,N_12581);
or U18285 (N_18285,N_13151,N_10742);
and U18286 (N_18286,N_11065,N_14494);
nor U18287 (N_18287,N_13168,N_10126);
or U18288 (N_18288,N_11521,N_13796);
nand U18289 (N_18289,N_11422,N_10942);
or U18290 (N_18290,N_11687,N_10220);
xnor U18291 (N_18291,N_10602,N_10035);
or U18292 (N_18292,N_12466,N_13897);
nand U18293 (N_18293,N_14386,N_13297);
nand U18294 (N_18294,N_11792,N_12402);
nor U18295 (N_18295,N_12450,N_10266);
and U18296 (N_18296,N_14711,N_11696);
nor U18297 (N_18297,N_10582,N_14576);
nor U18298 (N_18298,N_14009,N_14732);
nor U18299 (N_18299,N_14588,N_14482);
nand U18300 (N_18300,N_12602,N_10794);
nor U18301 (N_18301,N_10504,N_11020);
nor U18302 (N_18302,N_13962,N_10133);
nand U18303 (N_18303,N_11048,N_13331);
nor U18304 (N_18304,N_13999,N_13981);
nand U18305 (N_18305,N_12938,N_11664);
and U18306 (N_18306,N_12322,N_11255);
nand U18307 (N_18307,N_11618,N_12627);
xnor U18308 (N_18308,N_10216,N_11520);
nand U18309 (N_18309,N_10814,N_12905);
nor U18310 (N_18310,N_10884,N_12432);
nor U18311 (N_18311,N_12337,N_11528);
xnor U18312 (N_18312,N_13729,N_12867);
nand U18313 (N_18313,N_13663,N_12588);
nand U18314 (N_18314,N_11949,N_10456);
nand U18315 (N_18315,N_10076,N_11152);
nor U18316 (N_18316,N_11260,N_11615);
or U18317 (N_18317,N_10526,N_12659);
and U18318 (N_18318,N_13967,N_12472);
nor U18319 (N_18319,N_11375,N_12418);
and U18320 (N_18320,N_10385,N_10996);
nor U18321 (N_18321,N_12026,N_11947);
or U18322 (N_18322,N_10281,N_13905);
and U18323 (N_18323,N_14336,N_12335);
nand U18324 (N_18324,N_11260,N_11203);
or U18325 (N_18325,N_12798,N_12070);
nand U18326 (N_18326,N_10288,N_11832);
nor U18327 (N_18327,N_13216,N_14903);
or U18328 (N_18328,N_14231,N_12738);
nand U18329 (N_18329,N_14310,N_13237);
or U18330 (N_18330,N_11895,N_14271);
and U18331 (N_18331,N_13437,N_14264);
nand U18332 (N_18332,N_10352,N_11620);
or U18333 (N_18333,N_13689,N_11760);
nand U18334 (N_18334,N_13209,N_11586);
or U18335 (N_18335,N_10377,N_13614);
and U18336 (N_18336,N_12143,N_14908);
nor U18337 (N_18337,N_12538,N_13089);
nor U18338 (N_18338,N_14963,N_13599);
and U18339 (N_18339,N_14574,N_11473);
or U18340 (N_18340,N_14600,N_11305);
nand U18341 (N_18341,N_11806,N_12483);
or U18342 (N_18342,N_11795,N_10935);
nor U18343 (N_18343,N_14808,N_11177);
and U18344 (N_18344,N_10891,N_13079);
nand U18345 (N_18345,N_11501,N_11062);
nor U18346 (N_18346,N_13269,N_10173);
or U18347 (N_18347,N_12689,N_10663);
nand U18348 (N_18348,N_11657,N_10283);
nor U18349 (N_18349,N_10519,N_14212);
or U18350 (N_18350,N_13528,N_12210);
nand U18351 (N_18351,N_12484,N_13274);
nor U18352 (N_18352,N_14443,N_13188);
and U18353 (N_18353,N_11987,N_10554);
nor U18354 (N_18354,N_14787,N_14564);
nor U18355 (N_18355,N_13608,N_11351);
nor U18356 (N_18356,N_11016,N_12243);
or U18357 (N_18357,N_10703,N_10031);
nand U18358 (N_18358,N_13723,N_11604);
or U18359 (N_18359,N_11732,N_12480);
nand U18360 (N_18360,N_11431,N_12849);
or U18361 (N_18361,N_11185,N_12033);
and U18362 (N_18362,N_11588,N_10729);
nand U18363 (N_18363,N_14147,N_11226);
nor U18364 (N_18364,N_12903,N_11411);
or U18365 (N_18365,N_10236,N_11858);
and U18366 (N_18366,N_13233,N_10728);
and U18367 (N_18367,N_13185,N_12580);
or U18368 (N_18368,N_12468,N_10081);
nor U18369 (N_18369,N_10465,N_13052);
nor U18370 (N_18370,N_14271,N_11011);
and U18371 (N_18371,N_14233,N_12792);
nor U18372 (N_18372,N_12199,N_14424);
nand U18373 (N_18373,N_11554,N_14562);
or U18374 (N_18374,N_10403,N_13803);
nand U18375 (N_18375,N_14714,N_10260);
or U18376 (N_18376,N_11595,N_14647);
and U18377 (N_18377,N_13352,N_12517);
and U18378 (N_18378,N_13276,N_14082);
nand U18379 (N_18379,N_13760,N_13547);
nor U18380 (N_18380,N_13050,N_14308);
or U18381 (N_18381,N_12837,N_12688);
and U18382 (N_18382,N_14904,N_12623);
or U18383 (N_18383,N_10398,N_11569);
nor U18384 (N_18384,N_11051,N_10515);
nor U18385 (N_18385,N_11315,N_10884);
or U18386 (N_18386,N_13103,N_11472);
or U18387 (N_18387,N_12509,N_10040);
and U18388 (N_18388,N_12122,N_10114);
or U18389 (N_18389,N_10543,N_13273);
nor U18390 (N_18390,N_14044,N_10500);
nand U18391 (N_18391,N_13865,N_12339);
nand U18392 (N_18392,N_10172,N_10707);
or U18393 (N_18393,N_14276,N_13981);
and U18394 (N_18394,N_13904,N_10652);
nor U18395 (N_18395,N_12215,N_11087);
nand U18396 (N_18396,N_11199,N_11779);
nor U18397 (N_18397,N_12224,N_12943);
nand U18398 (N_18398,N_12753,N_12730);
nor U18399 (N_18399,N_10847,N_11451);
or U18400 (N_18400,N_14500,N_14698);
nor U18401 (N_18401,N_13840,N_10103);
and U18402 (N_18402,N_12546,N_14944);
nand U18403 (N_18403,N_10291,N_14035);
and U18404 (N_18404,N_13748,N_14496);
nand U18405 (N_18405,N_10112,N_12155);
and U18406 (N_18406,N_14487,N_10500);
or U18407 (N_18407,N_14297,N_10841);
nor U18408 (N_18408,N_12270,N_10090);
and U18409 (N_18409,N_10421,N_10866);
or U18410 (N_18410,N_11140,N_12671);
and U18411 (N_18411,N_13518,N_13764);
nand U18412 (N_18412,N_12319,N_14295);
or U18413 (N_18413,N_14054,N_11374);
and U18414 (N_18414,N_12420,N_11661);
or U18415 (N_18415,N_12470,N_12243);
or U18416 (N_18416,N_11885,N_12087);
nand U18417 (N_18417,N_12169,N_12046);
nor U18418 (N_18418,N_14142,N_11914);
and U18419 (N_18419,N_10438,N_12814);
nor U18420 (N_18420,N_10602,N_11190);
or U18421 (N_18421,N_10819,N_14967);
and U18422 (N_18422,N_13715,N_14065);
or U18423 (N_18423,N_10995,N_12536);
nor U18424 (N_18424,N_13396,N_13934);
nand U18425 (N_18425,N_10575,N_12366);
and U18426 (N_18426,N_14455,N_14647);
nand U18427 (N_18427,N_12332,N_13538);
nand U18428 (N_18428,N_12862,N_13046);
or U18429 (N_18429,N_12463,N_12710);
and U18430 (N_18430,N_13432,N_14091);
nand U18431 (N_18431,N_11944,N_14571);
nor U18432 (N_18432,N_13610,N_10585);
nand U18433 (N_18433,N_10514,N_10806);
or U18434 (N_18434,N_13694,N_13331);
or U18435 (N_18435,N_13980,N_14880);
or U18436 (N_18436,N_14870,N_10336);
or U18437 (N_18437,N_11648,N_12090);
or U18438 (N_18438,N_14753,N_10258);
or U18439 (N_18439,N_13939,N_10969);
nor U18440 (N_18440,N_13000,N_13910);
and U18441 (N_18441,N_11671,N_14856);
and U18442 (N_18442,N_12744,N_13729);
nor U18443 (N_18443,N_13444,N_10799);
nand U18444 (N_18444,N_12595,N_11876);
and U18445 (N_18445,N_13006,N_10437);
nor U18446 (N_18446,N_11678,N_14742);
nand U18447 (N_18447,N_13131,N_11608);
and U18448 (N_18448,N_12140,N_14859);
nand U18449 (N_18449,N_11966,N_13698);
nand U18450 (N_18450,N_14104,N_11726);
xnor U18451 (N_18451,N_14093,N_13394);
and U18452 (N_18452,N_11574,N_13981);
nand U18453 (N_18453,N_14829,N_10710);
nand U18454 (N_18454,N_11127,N_11383);
and U18455 (N_18455,N_10065,N_13221);
and U18456 (N_18456,N_10916,N_10301);
and U18457 (N_18457,N_13635,N_11924);
or U18458 (N_18458,N_13252,N_10601);
nand U18459 (N_18459,N_14790,N_11531);
or U18460 (N_18460,N_13760,N_13743);
nor U18461 (N_18461,N_11856,N_10465);
and U18462 (N_18462,N_13290,N_12553);
or U18463 (N_18463,N_14089,N_12823);
xor U18464 (N_18464,N_11498,N_11415);
nand U18465 (N_18465,N_13412,N_14170);
nor U18466 (N_18466,N_11158,N_13594);
nor U18467 (N_18467,N_11728,N_13507);
nand U18468 (N_18468,N_13113,N_11985);
nor U18469 (N_18469,N_13489,N_14317);
nand U18470 (N_18470,N_11518,N_13241);
xor U18471 (N_18471,N_11312,N_11757);
and U18472 (N_18472,N_12702,N_12761);
and U18473 (N_18473,N_13359,N_10368);
or U18474 (N_18474,N_12235,N_13198);
or U18475 (N_18475,N_13828,N_14190);
and U18476 (N_18476,N_10114,N_12120);
nor U18477 (N_18477,N_10794,N_11777);
nand U18478 (N_18478,N_14941,N_13940);
or U18479 (N_18479,N_11270,N_11151);
xnor U18480 (N_18480,N_12757,N_11969);
nand U18481 (N_18481,N_14416,N_10441);
and U18482 (N_18482,N_10157,N_10956);
or U18483 (N_18483,N_13682,N_10314);
or U18484 (N_18484,N_13419,N_10364);
or U18485 (N_18485,N_14524,N_13847);
and U18486 (N_18486,N_14628,N_14273);
xor U18487 (N_18487,N_10137,N_10315);
or U18488 (N_18488,N_14596,N_12512);
xnor U18489 (N_18489,N_13534,N_13775);
or U18490 (N_18490,N_14914,N_13179);
and U18491 (N_18491,N_11483,N_12080);
nand U18492 (N_18492,N_10320,N_14334);
and U18493 (N_18493,N_13678,N_13707);
nand U18494 (N_18494,N_12975,N_11657);
nand U18495 (N_18495,N_12596,N_10656);
nand U18496 (N_18496,N_13578,N_12715);
and U18497 (N_18497,N_12952,N_14256);
and U18498 (N_18498,N_10283,N_12470);
or U18499 (N_18499,N_11161,N_12843);
and U18500 (N_18500,N_11114,N_12994);
or U18501 (N_18501,N_11630,N_12509);
xor U18502 (N_18502,N_11780,N_11721);
or U18503 (N_18503,N_12662,N_10084);
xnor U18504 (N_18504,N_11999,N_10873);
nor U18505 (N_18505,N_12175,N_14211);
nand U18506 (N_18506,N_11615,N_11324);
and U18507 (N_18507,N_11748,N_12314);
or U18508 (N_18508,N_11693,N_13054);
and U18509 (N_18509,N_12679,N_10520);
or U18510 (N_18510,N_13433,N_14586);
nor U18511 (N_18511,N_10230,N_14416);
nor U18512 (N_18512,N_12489,N_11448);
nand U18513 (N_18513,N_14334,N_12796);
and U18514 (N_18514,N_13137,N_11073);
or U18515 (N_18515,N_10869,N_12690);
and U18516 (N_18516,N_12583,N_14364);
nor U18517 (N_18517,N_12919,N_10325);
nand U18518 (N_18518,N_13753,N_13717);
nand U18519 (N_18519,N_11545,N_13526);
nand U18520 (N_18520,N_10019,N_10608);
or U18521 (N_18521,N_12267,N_13072);
and U18522 (N_18522,N_12980,N_12921);
nor U18523 (N_18523,N_14587,N_13932);
or U18524 (N_18524,N_11456,N_10802);
and U18525 (N_18525,N_14957,N_11723);
or U18526 (N_18526,N_10197,N_13018);
and U18527 (N_18527,N_10473,N_11141);
nand U18528 (N_18528,N_10920,N_12499);
or U18529 (N_18529,N_10540,N_12715);
or U18530 (N_18530,N_10966,N_13625);
nand U18531 (N_18531,N_12033,N_10619);
and U18532 (N_18532,N_12061,N_13917);
or U18533 (N_18533,N_13811,N_11148);
nor U18534 (N_18534,N_13698,N_13225);
or U18535 (N_18535,N_12753,N_13837);
and U18536 (N_18536,N_12373,N_12214);
nand U18537 (N_18537,N_13238,N_11633);
and U18538 (N_18538,N_10627,N_14675);
nor U18539 (N_18539,N_13324,N_13138);
xor U18540 (N_18540,N_12227,N_10787);
or U18541 (N_18541,N_14077,N_13891);
or U18542 (N_18542,N_13210,N_13719);
nand U18543 (N_18543,N_11680,N_13129);
and U18544 (N_18544,N_13918,N_12744);
and U18545 (N_18545,N_11099,N_12550);
and U18546 (N_18546,N_13914,N_10566);
or U18547 (N_18547,N_12302,N_12844);
and U18548 (N_18548,N_11962,N_12909);
nand U18549 (N_18549,N_10726,N_13235);
nor U18550 (N_18550,N_11408,N_12599);
nand U18551 (N_18551,N_14268,N_10612);
nand U18552 (N_18552,N_11349,N_12040);
xor U18553 (N_18553,N_14254,N_14522);
nor U18554 (N_18554,N_14049,N_12297);
and U18555 (N_18555,N_10561,N_14627);
and U18556 (N_18556,N_12568,N_11593);
nor U18557 (N_18557,N_13079,N_14847);
and U18558 (N_18558,N_11673,N_13216);
and U18559 (N_18559,N_12806,N_13507);
nand U18560 (N_18560,N_12351,N_10452);
or U18561 (N_18561,N_13869,N_14950);
nor U18562 (N_18562,N_13234,N_13192);
or U18563 (N_18563,N_12107,N_11912);
and U18564 (N_18564,N_10179,N_14474);
nand U18565 (N_18565,N_11270,N_10729);
and U18566 (N_18566,N_13544,N_11226);
and U18567 (N_18567,N_14953,N_11349);
and U18568 (N_18568,N_13930,N_12714);
and U18569 (N_18569,N_13331,N_12998);
or U18570 (N_18570,N_12127,N_14585);
or U18571 (N_18571,N_10953,N_12715);
or U18572 (N_18572,N_14754,N_12050);
or U18573 (N_18573,N_11962,N_12265);
or U18574 (N_18574,N_10966,N_14918);
or U18575 (N_18575,N_12718,N_12693);
or U18576 (N_18576,N_14001,N_14889);
or U18577 (N_18577,N_13608,N_12294);
or U18578 (N_18578,N_14283,N_12845);
and U18579 (N_18579,N_10119,N_13595);
or U18580 (N_18580,N_14201,N_13572);
nor U18581 (N_18581,N_11960,N_11797);
or U18582 (N_18582,N_14150,N_12010);
or U18583 (N_18583,N_12876,N_12277);
nor U18584 (N_18584,N_11988,N_12112);
and U18585 (N_18585,N_14976,N_10844);
nor U18586 (N_18586,N_14991,N_11955);
nor U18587 (N_18587,N_14059,N_13157);
nor U18588 (N_18588,N_12776,N_12539);
nor U18589 (N_18589,N_12664,N_13504);
xor U18590 (N_18590,N_13248,N_12565);
and U18591 (N_18591,N_13098,N_14877);
nand U18592 (N_18592,N_10034,N_14977);
nor U18593 (N_18593,N_13326,N_12791);
nor U18594 (N_18594,N_12893,N_10266);
or U18595 (N_18595,N_10906,N_14520);
nor U18596 (N_18596,N_12967,N_10952);
or U18597 (N_18597,N_14424,N_10636);
nor U18598 (N_18598,N_11566,N_14014);
and U18599 (N_18599,N_11868,N_10924);
xor U18600 (N_18600,N_10529,N_10546);
or U18601 (N_18601,N_10435,N_14676);
nor U18602 (N_18602,N_11692,N_10358);
nand U18603 (N_18603,N_14733,N_11894);
nor U18604 (N_18604,N_11786,N_14561);
and U18605 (N_18605,N_13291,N_12249);
and U18606 (N_18606,N_12462,N_14922);
and U18607 (N_18607,N_13748,N_10399);
or U18608 (N_18608,N_11146,N_13570);
nand U18609 (N_18609,N_12259,N_10305);
and U18610 (N_18610,N_14421,N_11710);
nand U18611 (N_18611,N_14617,N_12944);
nor U18612 (N_18612,N_10308,N_14896);
or U18613 (N_18613,N_13368,N_13587);
xor U18614 (N_18614,N_10214,N_10196);
or U18615 (N_18615,N_10902,N_10813);
and U18616 (N_18616,N_11712,N_12727);
and U18617 (N_18617,N_12493,N_12321);
nor U18618 (N_18618,N_12689,N_13684);
and U18619 (N_18619,N_13679,N_12198);
nor U18620 (N_18620,N_12704,N_12743);
and U18621 (N_18621,N_11773,N_12807);
nor U18622 (N_18622,N_10200,N_12794);
nand U18623 (N_18623,N_13229,N_12637);
and U18624 (N_18624,N_14795,N_12142);
nand U18625 (N_18625,N_11006,N_14677);
and U18626 (N_18626,N_13541,N_10806);
nor U18627 (N_18627,N_13042,N_10394);
or U18628 (N_18628,N_14727,N_14753);
and U18629 (N_18629,N_13856,N_13646);
nor U18630 (N_18630,N_14656,N_13348);
xor U18631 (N_18631,N_11340,N_14291);
or U18632 (N_18632,N_14255,N_10500);
nor U18633 (N_18633,N_14219,N_11270);
or U18634 (N_18634,N_10867,N_12381);
or U18635 (N_18635,N_11882,N_14237);
nand U18636 (N_18636,N_13053,N_10366);
nand U18637 (N_18637,N_13231,N_10128);
or U18638 (N_18638,N_14545,N_13636);
or U18639 (N_18639,N_11956,N_11614);
or U18640 (N_18640,N_13610,N_14190);
or U18641 (N_18641,N_14067,N_12850);
nor U18642 (N_18642,N_10540,N_11132);
nand U18643 (N_18643,N_10467,N_14246);
and U18644 (N_18644,N_11201,N_14568);
xor U18645 (N_18645,N_12317,N_13404);
xor U18646 (N_18646,N_12349,N_10125);
and U18647 (N_18647,N_14152,N_10491);
or U18648 (N_18648,N_13177,N_12859);
or U18649 (N_18649,N_12506,N_13232);
or U18650 (N_18650,N_12622,N_10892);
nand U18651 (N_18651,N_11720,N_14210);
and U18652 (N_18652,N_13151,N_10732);
nor U18653 (N_18653,N_12762,N_10499);
nor U18654 (N_18654,N_13115,N_12039);
nor U18655 (N_18655,N_13781,N_10455);
nor U18656 (N_18656,N_10336,N_14667);
or U18657 (N_18657,N_11260,N_12382);
nor U18658 (N_18658,N_11641,N_11640);
or U18659 (N_18659,N_12985,N_14256);
or U18660 (N_18660,N_10343,N_14777);
xor U18661 (N_18661,N_14968,N_13026);
nor U18662 (N_18662,N_11095,N_10709);
and U18663 (N_18663,N_12056,N_11601);
nand U18664 (N_18664,N_14964,N_13437);
and U18665 (N_18665,N_12678,N_13922);
xor U18666 (N_18666,N_11935,N_12979);
and U18667 (N_18667,N_10624,N_12870);
nand U18668 (N_18668,N_10532,N_13564);
nor U18669 (N_18669,N_14678,N_10146);
xor U18670 (N_18670,N_11588,N_10487);
or U18671 (N_18671,N_14488,N_10173);
and U18672 (N_18672,N_12180,N_10887);
nand U18673 (N_18673,N_14707,N_14570);
and U18674 (N_18674,N_10128,N_14855);
or U18675 (N_18675,N_13522,N_11305);
nor U18676 (N_18676,N_11189,N_13027);
nand U18677 (N_18677,N_11759,N_10108);
nand U18678 (N_18678,N_11143,N_11961);
nor U18679 (N_18679,N_14321,N_11673);
nand U18680 (N_18680,N_10448,N_10717);
nand U18681 (N_18681,N_13689,N_14439);
nand U18682 (N_18682,N_13782,N_11110);
nand U18683 (N_18683,N_10615,N_10376);
and U18684 (N_18684,N_13740,N_13470);
nand U18685 (N_18685,N_12833,N_10672);
or U18686 (N_18686,N_14165,N_14576);
nor U18687 (N_18687,N_11097,N_11155);
and U18688 (N_18688,N_12555,N_14505);
and U18689 (N_18689,N_12381,N_10634);
and U18690 (N_18690,N_14259,N_12614);
nor U18691 (N_18691,N_12401,N_11008);
nor U18692 (N_18692,N_13034,N_13627);
and U18693 (N_18693,N_12595,N_11621);
and U18694 (N_18694,N_12275,N_10316);
nor U18695 (N_18695,N_13411,N_11563);
or U18696 (N_18696,N_13621,N_13409);
and U18697 (N_18697,N_14918,N_13244);
and U18698 (N_18698,N_13797,N_13684);
or U18699 (N_18699,N_11887,N_10751);
or U18700 (N_18700,N_10818,N_14109);
nor U18701 (N_18701,N_12894,N_14004);
and U18702 (N_18702,N_10706,N_14501);
or U18703 (N_18703,N_14990,N_13028);
nor U18704 (N_18704,N_12689,N_14319);
and U18705 (N_18705,N_14211,N_10365);
or U18706 (N_18706,N_11194,N_12264);
nor U18707 (N_18707,N_13708,N_12628);
nand U18708 (N_18708,N_10382,N_12016);
or U18709 (N_18709,N_11688,N_10140);
nand U18710 (N_18710,N_11790,N_10463);
or U18711 (N_18711,N_11356,N_10351);
nand U18712 (N_18712,N_12618,N_14267);
and U18713 (N_18713,N_13149,N_14683);
nand U18714 (N_18714,N_10983,N_11929);
or U18715 (N_18715,N_13799,N_12252);
nand U18716 (N_18716,N_14965,N_14691);
nand U18717 (N_18717,N_10392,N_10634);
nand U18718 (N_18718,N_13194,N_11688);
nor U18719 (N_18719,N_13189,N_13481);
nor U18720 (N_18720,N_12629,N_13287);
and U18721 (N_18721,N_12169,N_12508);
nor U18722 (N_18722,N_12226,N_13034);
nand U18723 (N_18723,N_14949,N_11162);
and U18724 (N_18724,N_14708,N_10854);
or U18725 (N_18725,N_13543,N_10184);
and U18726 (N_18726,N_14920,N_12374);
nor U18727 (N_18727,N_10709,N_10401);
nand U18728 (N_18728,N_14622,N_13481);
and U18729 (N_18729,N_10764,N_12979);
nand U18730 (N_18730,N_10578,N_12028);
nor U18731 (N_18731,N_10302,N_12707);
or U18732 (N_18732,N_11864,N_13683);
nor U18733 (N_18733,N_14447,N_14814);
nor U18734 (N_18734,N_11716,N_11527);
or U18735 (N_18735,N_14399,N_11701);
and U18736 (N_18736,N_11467,N_13963);
nand U18737 (N_18737,N_13006,N_12759);
xnor U18738 (N_18738,N_14986,N_10065);
and U18739 (N_18739,N_12103,N_14298);
nand U18740 (N_18740,N_12131,N_10762);
and U18741 (N_18741,N_13338,N_13455);
and U18742 (N_18742,N_11872,N_11570);
nand U18743 (N_18743,N_14154,N_11958);
or U18744 (N_18744,N_12725,N_14408);
nand U18745 (N_18745,N_10920,N_12297);
and U18746 (N_18746,N_11935,N_14028);
nand U18747 (N_18747,N_10203,N_12372);
and U18748 (N_18748,N_10680,N_11580);
or U18749 (N_18749,N_10190,N_12631);
and U18750 (N_18750,N_10834,N_14066);
or U18751 (N_18751,N_14244,N_13434);
nor U18752 (N_18752,N_13486,N_13380);
and U18753 (N_18753,N_10961,N_12290);
nor U18754 (N_18754,N_10512,N_10227);
and U18755 (N_18755,N_13405,N_10725);
nand U18756 (N_18756,N_12535,N_13766);
nand U18757 (N_18757,N_14851,N_11834);
and U18758 (N_18758,N_11995,N_11443);
nor U18759 (N_18759,N_11028,N_12361);
nand U18760 (N_18760,N_11566,N_11084);
nand U18761 (N_18761,N_14928,N_11438);
nor U18762 (N_18762,N_11568,N_14456);
and U18763 (N_18763,N_11362,N_11014);
nand U18764 (N_18764,N_11559,N_13650);
and U18765 (N_18765,N_14544,N_13127);
nor U18766 (N_18766,N_11016,N_10020);
nand U18767 (N_18767,N_14831,N_10238);
or U18768 (N_18768,N_12478,N_12421);
or U18769 (N_18769,N_14724,N_11550);
or U18770 (N_18770,N_14960,N_12457);
nand U18771 (N_18771,N_12388,N_11633);
nor U18772 (N_18772,N_11315,N_13019);
or U18773 (N_18773,N_11591,N_11874);
nor U18774 (N_18774,N_11055,N_14559);
nand U18775 (N_18775,N_10899,N_12794);
xnor U18776 (N_18776,N_14848,N_11849);
or U18777 (N_18777,N_11240,N_11605);
or U18778 (N_18778,N_14750,N_14328);
nor U18779 (N_18779,N_10070,N_11479);
and U18780 (N_18780,N_12042,N_12739);
and U18781 (N_18781,N_14074,N_12015);
and U18782 (N_18782,N_12719,N_10560);
nand U18783 (N_18783,N_13649,N_14841);
nor U18784 (N_18784,N_10487,N_10635);
and U18785 (N_18785,N_13771,N_10575);
or U18786 (N_18786,N_10897,N_13036);
nor U18787 (N_18787,N_10773,N_12102);
nor U18788 (N_18788,N_11320,N_14313);
and U18789 (N_18789,N_12289,N_11761);
or U18790 (N_18790,N_14868,N_12385);
or U18791 (N_18791,N_14394,N_10223);
or U18792 (N_18792,N_10877,N_11180);
or U18793 (N_18793,N_12736,N_10465);
nor U18794 (N_18794,N_14958,N_14669);
nor U18795 (N_18795,N_11249,N_13261);
or U18796 (N_18796,N_13816,N_10986);
nor U18797 (N_18797,N_12943,N_12250);
and U18798 (N_18798,N_12168,N_12067);
and U18799 (N_18799,N_13036,N_10850);
or U18800 (N_18800,N_10870,N_10684);
nand U18801 (N_18801,N_10579,N_12590);
and U18802 (N_18802,N_14883,N_14056);
and U18803 (N_18803,N_13932,N_11747);
nor U18804 (N_18804,N_13964,N_10761);
or U18805 (N_18805,N_11488,N_13186);
and U18806 (N_18806,N_12158,N_14601);
nor U18807 (N_18807,N_14331,N_14629);
nand U18808 (N_18808,N_10231,N_11864);
and U18809 (N_18809,N_11020,N_13331);
or U18810 (N_18810,N_12635,N_14750);
and U18811 (N_18811,N_11891,N_10192);
nor U18812 (N_18812,N_10150,N_10907);
nor U18813 (N_18813,N_10881,N_14619);
nand U18814 (N_18814,N_11973,N_11509);
and U18815 (N_18815,N_10702,N_13120);
and U18816 (N_18816,N_13167,N_11102);
nand U18817 (N_18817,N_12257,N_13255);
and U18818 (N_18818,N_14411,N_10130);
nand U18819 (N_18819,N_10805,N_10889);
and U18820 (N_18820,N_11424,N_13285);
nor U18821 (N_18821,N_13399,N_13208);
and U18822 (N_18822,N_13604,N_11730);
nand U18823 (N_18823,N_10757,N_14706);
and U18824 (N_18824,N_10554,N_11564);
nand U18825 (N_18825,N_13102,N_12085);
and U18826 (N_18826,N_12242,N_10050);
nor U18827 (N_18827,N_11209,N_14925);
nor U18828 (N_18828,N_14953,N_14195);
nand U18829 (N_18829,N_13258,N_10577);
or U18830 (N_18830,N_10666,N_10682);
nor U18831 (N_18831,N_13201,N_13761);
nand U18832 (N_18832,N_10741,N_10883);
and U18833 (N_18833,N_12395,N_10453);
and U18834 (N_18834,N_11168,N_13020);
nand U18835 (N_18835,N_10326,N_12024);
nor U18836 (N_18836,N_10161,N_11274);
xor U18837 (N_18837,N_10791,N_11276);
or U18838 (N_18838,N_11693,N_14224);
xnor U18839 (N_18839,N_11320,N_14728);
nor U18840 (N_18840,N_11447,N_10867);
nand U18841 (N_18841,N_10648,N_12622);
and U18842 (N_18842,N_10297,N_13094);
and U18843 (N_18843,N_13869,N_12701);
nor U18844 (N_18844,N_13094,N_11872);
nand U18845 (N_18845,N_11773,N_11521);
nor U18846 (N_18846,N_11091,N_11117);
or U18847 (N_18847,N_10639,N_14394);
nand U18848 (N_18848,N_10138,N_13254);
nand U18849 (N_18849,N_13120,N_10921);
nand U18850 (N_18850,N_13087,N_14962);
nor U18851 (N_18851,N_13537,N_10548);
nor U18852 (N_18852,N_12118,N_12852);
and U18853 (N_18853,N_13101,N_13797);
nand U18854 (N_18854,N_12304,N_11793);
nand U18855 (N_18855,N_12516,N_11021);
nor U18856 (N_18856,N_13358,N_14102);
or U18857 (N_18857,N_12913,N_14205);
nor U18858 (N_18858,N_14273,N_10041);
or U18859 (N_18859,N_12581,N_10376);
nor U18860 (N_18860,N_12956,N_13445);
or U18861 (N_18861,N_14331,N_11605);
and U18862 (N_18862,N_14295,N_13180);
nor U18863 (N_18863,N_10755,N_12091);
or U18864 (N_18864,N_14741,N_13349);
or U18865 (N_18865,N_12199,N_13413);
nand U18866 (N_18866,N_11022,N_12534);
nand U18867 (N_18867,N_14995,N_10778);
nor U18868 (N_18868,N_14966,N_13858);
or U18869 (N_18869,N_12307,N_12255);
nor U18870 (N_18870,N_14923,N_11369);
or U18871 (N_18871,N_10472,N_11402);
nor U18872 (N_18872,N_14949,N_12934);
and U18873 (N_18873,N_14493,N_14657);
nand U18874 (N_18874,N_10121,N_13581);
nor U18875 (N_18875,N_10993,N_10624);
nand U18876 (N_18876,N_14485,N_12409);
xor U18877 (N_18877,N_14024,N_12557);
and U18878 (N_18878,N_10585,N_14438);
nand U18879 (N_18879,N_10415,N_14029);
nor U18880 (N_18880,N_14487,N_10832);
and U18881 (N_18881,N_13531,N_11234);
nand U18882 (N_18882,N_12902,N_11173);
nand U18883 (N_18883,N_13818,N_14649);
and U18884 (N_18884,N_13481,N_11732);
nor U18885 (N_18885,N_12395,N_13325);
and U18886 (N_18886,N_11273,N_12280);
or U18887 (N_18887,N_13373,N_11757);
and U18888 (N_18888,N_12088,N_13244);
and U18889 (N_18889,N_12941,N_10528);
nor U18890 (N_18890,N_13821,N_13418);
nand U18891 (N_18891,N_11241,N_12569);
nand U18892 (N_18892,N_14430,N_12463);
nand U18893 (N_18893,N_13066,N_13124);
and U18894 (N_18894,N_11517,N_11354);
or U18895 (N_18895,N_10199,N_10123);
and U18896 (N_18896,N_13671,N_14108);
or U18897 (N_18897,N_13567,N_13706);
and U18898 (N_18898,N_10300,N_12351);
nand U18899 (N_18899,N_14747,N_13804);
and U18900 (N_18900,N_10895,N_13141);
nor U18901 (N_18901,N_12397,N_10243);
nand U18902 (N_18902,N_11014,N_12614);
and U18903 (N_18903,N_12048,N_14908);
or U18904 (N_18904,N_11186,N_11516);
or U18905 (N_18905,N_13443,N_11263);
and U18906 (N_18906,N_10430,N_13871);
or U18907 (N_18907,N_11528,N_13930);
nor U18908 (N_18908,N_12343,N_10867);
or U18909 (N_18909,N_12780,N_13240);
and U18910 (N_18910,N_11195,N_10272);
and U18911 (N_18911,N_12040,N_14051);
nand U18912 (N_18912,N_11695,N_12435);
and U18913 (N_18913,N_11522,N_12551);
or U18914 (N_18914,N_12133,N_10209);
nor U18915 (N_18915,N_12456,N_13224);
or U18916 (N_18916,N_13554,N_11334);
nand U18917 (N_18917,N_12269,N_13099);
nor U18918 (N_18918,N_10588,N_14627);
or U18919 (N_18919,N_12421,N_14306);
nand U18920 (N_18920,N_12851,N_14312);
nor U18921 (N_18921,N_10613,N_13378);
or U18922 (N_18922,N_11529,N_13496);
and U18923 (N_18923,N_13803,N_13126);
nand U18924 (N_18924,N_13135,N_13724);
or U18925 (N_18925,N_14479,N_11831);
nand U18926 (N_18926,N_11222,N_11539);
and U18927 (N_18927,N_13191,N_14960);
and U18928 (N_18928,N_13078,N_13481);
nor U18929 (N_18929,N_12019,N_13736);
nor U18930 (N_18930,N_10667,N_10000);
xnor U18931 (N_18931,N_11381,N_12944);
or U18932 (N_18932,N_12197,N_14800);
or U18933 (N_18933,N_11344,N_12308);
or U18934 (N_18934,N_13455,N_12855);
nand U18935 (N_18935,N_13187,N_10610);
nor U18936 (N_18936,N_14448,N_12188);
nor U18937 (N_18937,N_14947,N_14375);
and U18938 (N_18938,N_12394,N_12229);
or U18939 (N_18939,N_11383,N_12330);
and U18940 (N_18940,N_13152,N_11381);
nand U18941 (N_18941,N_10484,N_13279);
nor U18942 (N_18942,N_14184,N_12165);
or U18943 (N_18943,N_11232,N_14714);
nand U18944 (N_18944,N_12769,N_10122);
nand U18945 (N_18945,N_14504,N_11087);
or U18946 (N_18946,N_14944,N_10770);
or U18947 (N_18947,N_11806,N_12801);
or U18948 (N_18948,N_11271,N_12586);
and U18949 (N_18949,N_11506,N_10990);
nand U18950 (N_18950,N_13015,N_10225);
nor U18951 (N_18951,N_10185,N_14790);
and U18952 (N_18952,N_13735,N_10232);
nor U18953 (N_18953,N_12338,N_11779);
and U18954 (N_18954,N_10039,N_10874);
and U18955 (N_18955,N_10315,N_12655);
or U18956 (N_18956,N_12791,N_10374);
nand U18957 (N_18957,N_13438,N_10861);
nand U18958 (N_18958,N_10261,N_11556);
nor U18959 (N_18959,N_13587,N_11694);
nor U18960 (N_18960,N_12442,N_14639);
or U18961 (N_18961,N_11733,N_13047);
nand U18962 (N_18962,N_13899,N_10180);
or U18963 (N_18963,N_13456,N_13362);
or U18964 (N_18964,N_14858,N_14946);
nand U18965 (N_18965,N_10846,N_14240);
nand U18966 (N_18966,N_14823,N_10205);
nor U18967 (N_18967,N_13857,N_10532);
nand U18968 (N_18968,N_11254,N_14389);
or U18969 (N_18969,N_10973,N_11425);
and U18970 (N_18970,N_12187,N_10268);
nand U18971 (N_18971,N_11145,N_12178);
nor U18972 (N_18972,N_13808,N_13778);
nor U18973 (N_18973,N_13109,N_10457);
or U18974 (N_18974,N_13561,N_10204);
or U18975 (N_18975,N_10697,N_10941);
nand U18976 (N_18976,N_10231,N_14053);
or U18977 (N_18977,N_13727,N_11332);
nand U18978 (N_18978,N_11673,N_14389);
or U18979 (N_18979,N_11121,N_10296);
or U18980 (N_18980,N_12260,N_13438);
or U18981 (N_18981,N_13153,N_13193);
nand U18982 (N_18982,N_14975,N_11136);
or U18983 (N_18983,N_11199,N_13953);
nor U18984 (N_18984,N_13807,N_12707);
nand U18985 (N_18985,N_10260,N_11961);
nand U18986 (N_18986,N_13785,N_12619);
and U18987 (N_18987,N_10625,N_14640);
nor U18988 (N_18988,N_11647,N_14817);
and U18989 (N_18989,N_10853,N_12109);
nand U18990 (N_18990,N_10555,N_12991);
or U18991 (N_18991,N_10692,N_10462);
nand U18992 (N_18992,N_11499,N_14804);
and U18993 (N_18993,N_11133,N_13980);
nor U18994 (N_18994,N_11558,N_14926);
nor U18995 (N_18995,N_11566,N_14303);
nor U18996 (N_18996,N_13527,N_12967);
and U18997 (N_18997,N_12188,N_12325);
nor U18998 (N_18998,N_14236,N_13445);
and U18999 (N_18999,N_11064,N_14058);
and U19000 (N_19000,N_10666,N_10129);
and U19001 (N_19001,N_14043,N_14210);
nand U19002 (N_19002,N_10544,N_14703);
and U19003 (N_19003,N_10384,N_11619);
nand U19004 (N_19004,N_12275,N_10056);
or U19005 (N_19005,N_14348,N_14526);
nor U19006 (N_19006,N_11904,N_11983);
and U19007 (N_19007,N_12229,N_10256);
and U19008 (N_19008,N_14889,N_14670);
xnor U19009 (N_19009,N_14488,N_10192);
and U19010 (N_19010,N_11164,N_12814);
and U19011 (N_19011,N_13011,N_14765);
xnor U19012 (N_19012,N_14319,N_14304);
and U19013 (N_19013,N_10214,N_11441);
and U19014 (N_19014,N_11154,N_13177);
nand U19015 (N_19015,N_11062,N_11363);
nor U19016 (N_19016,N_11120,N_14235);
nand U19017 (N_19017,N_14417,N_10069);
nand U19018 (N_19018,N_13540,N_10675);
and U19019 (N_19019,N_12908,N_13436);
nand U19020 (N_19020,N_13577,N_10067);
and U19021 (N_19021,N_13642,N_14585);
or U19022 (N_19022,N_13439,N_12423);
nor U19023 (N_19023,N_12711,N_11874);
and U19024 (N_19024,N_11352,N_10921);
or U19025 (N_19025,N_14446,N_12834);
and U19026 (N_19026,N_12377,N_10539);
and U19027 (N_19027,N_14489,N_13716);
nand U19028 (N_19028,N_13534,N_11054);
nand U19029 (N_19029,N_10551,N_11863);
or U19030 (N_19030,N_11526,N_13349);
nor U19031 (N_19031,N_11277,N_12661);
or U19032 (N_19032,N_12007,N_14620);
nor U19033 (N_19033,N_11479,N_13635);
or U19034 (N_19034,N_12261,N_14019);
nand U19035 (N_19035,N_12673,N_10598);
and U19036 (N_19036,N_11724,N_13899);
and U19037 (N_19037,N_14343,N_12542);
or U19038 (N_19038,N_10517,N_13890);
or U19039 (N_19039,N_12956,N_14636);
or U19040 (N_19040,N_14142,N_12085);
and U19041 (N_19041,N_11471,N_11727);
nand U19042 (N_19042,N_14811,N_10760);
nand U19043 (N_19043,N_10260,N_12284);
nor U19044 (N_19044,N_11858,N_10373);
nand U19045 (N_19045,N_12224,N_13460);
nor U19046 (N_19046,N_10044,N_13666);
nor U19047 (N_19047,N_14103,N_10241);
or U19048 (N_19048,N_14623,N_13990);
nand U19049 (N_19049,N_14139,N_12463);
and U19050 (N_19050,N_13314,N_13248);
nor U19051 (N_19051,N_10865,N_11372);
or U19052 (N_19052,N_11907,N_10548);
nand U19053 (N_19053,N_13721,N_13767);
and U19054 (N_19054,N_10977,N_11027);
and U19055 (N_19055,N_13915,N_12198);
and U19056 (N_19056,N_12438,N_13947);
or U19057 (N_19057,N_11728,N_11797);
nand U19058 (N_19058,N_14607,N_13959);
nand U19059 (N_19059,N_14710,N_11041);
nor U19060 (N_19060,N_13179,N_12608);
or U19061 (N_19061,N_13375,N_14461);
or U19062 (N_19062,N_14648,N_12033);
xor U19063 (N_19063,N_12706,N_13089);
and U19064 (N_19064,N_14326,N_13192);
nand U19065 (N_19065,N_11390,N_10036);
xnor U19066 (N_19066,N_14617,N_13453);
nand U19067 (N_19067,N_12088,N_13379);
and U19068 (N_19068,N_13214,N_14723);
and U19069 (N_19069,N_14783,N_12691);
nand U19070 (N_19070,N_12272,N_13405);
nor U19071 (N_19071,N_14352,N_14572);
and U19072 (N_19072,N_13117,N_10231);
nand U19073 (N_19073,N_10024,N_11722);
or U19074 (N_19074,N_14153,N_10549);
xor U19075 (N_19075,N_12740,N_12541);
or U19076 (N_19076,N_14845,N_14997);
nor U19077 (N_19077,N_10907,N_11211);
nor U19078 (N_19078,N_11209,N_10512);
and U19079 (N_19079,N_14570,N_14360);
and U19080 (N_19080,N_10412,N_14414);
nand U19081 (N_19081,N_12236,N_10080);
nand U19082 (N_19082,N_10398,N_13422);
and U19083 (N_19083,N_10843,N_12991);
and U19084 (N_19084,N_14976,N_11701);
nand U19085 (N_19085,N_10925,N_14506);
and U19086 (N_19086,N_14321,N_12153);
nand U19087 (N_19087,N_14073,N_12585);
nand U19088 (N_19088,N_11785,N_11528);
or U19089 (N_19089,N_12624,N_13751);
nor U19090 (N_19090,N_11523,N_13151);
nor U19091 (N_19091,N_11686,N_14681);
or U19092 (N_19092,N_10061,N_14576);
or U19093 (N_19093,N_12432,N_12978);
or U19094 (N_19094,N_14759,N_14008);
or U19095 (N_19095,N_12121,N_10385);
or U19096 (N_19096,N_13819,N_10699);
and U19097 (N_19097,N_14024,N_14815);
and U19098 (N_19098,N_12209,N_14036);
nor U19099 (N_19099,N_11729,N_10444);
nor U19100 (N_19100,N_10683,N_11702);
nor U19101 (N_19101,N_12335,N_13613);
or U19102 (N_19102,N_10913,N_12919);
and U19103 (N_19103,N_13681,N_10038);
or U19104 (N_19104,N_13133,N_12290);
or U19105 (N_19105,N_11670,N_11922);
nor U19106 (N_19106,N_11513,N_12236);
or U19107 (N_19107,N_12653,N_13031);
nor U19108 (N_19108,N_14455,N_13526);
and U19109 (N_19109,N_10726,N_14754);
or U19110 (N_19110,N_12626,N_12255);
and U19111 (N_19111,N_10138,N_14631);
and U19112 (N_19112,N_12004,N_10316);
or U19113 (N_19113,N_14098,N_10874);
nor U19114 (N_19114,N_10141,N_12476);
nand U19115 (N_19115,N_10259,N_12762);
nand U19116 (N_19116,N_12846,N_14719);
xor U19117 (N_19117,N_12183,N_13188);
nand U19118 (N_19118,N_10866,N_14647);
nand U19119 (N_19119,N_11086,N_13374);
nor U19120 (N_19120,N_13460,N_14958);
nand U19121 (N_19121,N_11588,N_12168);
and U19122 (N_19122,N_11292,N_13412);
nand U19123 (N_19123,N_14414,N_11482);
and U19124 (N_19124,N_14401,N_10260);
and U19125 (N_19125,N_12321,N_13098);
or U19126 (N_19126,N_13141,N_11541);
or U19127 (N_19127,N_12295,N_12380);
nor U19128 (N_19128,N_12003,N_10521);
and U19129 (N_19129,N_14655,N_14899);
and U19130 (N_19130,N_10961,N_11702);
nand U19131 (N_19131,N_10049,N_13788);
or U19132 (N_19132,N_13276,N_12427);
or U19133 (N_19133,N_10119,N_10443);
nand U19134 (N_19134,N_13405,N_13773);
nand U19135 (N_19135,N_12208,N_12324);
and U19136 (N_19136,N_14979,N_10256);
and U19137 (N_19137,N_14117,N_12621);
or U19138 (N_19138,N_10315,N_13976);
nand U19139 (N_19139,N_12453,N_13245);
nor U19140 (N_19140,N_10254,N_14052);
or U19141 (N_19141,N_11747,N_13786);
nand U19142 (N_19142,N_10758,N_12566);
and U19143 (N_19143,N_10702,N_12132);
nand U19144 (N_19144,N_10644,N_10256);
nor U19145 (N_19145,N_11811,N_14410);
nor U19146 (N_19146,N_13645,N_10696);
or U19147 (N_19147,N_12802,N_10477);
nor U19148 (N_19148,N_14085,N_11494);
or U19149 (N_19149,N_11966,N_10663);
nand U19150 (N_19150,N_14549,N_11080);
or U19151 (N_19151,N_12173,N_10531);
and U19152 (N_19152,N_13289,N_12338);
or U19153 (N_19153,N_10229,N_10413);
and U19154 (N_19154,N_12877,N_13983);
nor U19155 (N_19155,N_12379,N_12197);
nor U19156 (N_19156,N_13120,N_14987);
or U19157 (N_19157,N_11639,N_13049);
nand U19158 (N_19158,N_12415,N_11525);
nand U19159 (N_19159,N_11979,N_14486);
nand U19160 (N_19160,N_11851,N_10073);
or U19161 (N_19161,N_12288,N_12931);
or U19162 (N_19162,N_10220,N_12804);
xor U19163 (N_19163,N_12368,N_10770);
and U19164 (N_19164,N_10634,N_12796);
and U19165 (N_19165,N_10243,N_11816);
nand U19166 (N_19166,N_12311,N_10987);
xnor U19167 (N_19167,N_14515,N_12993);
and U19168 (N_19168,N_12196,N_11260);
and U19169 (N_19169,N_10748,N_11490);
nor U19170 (N_19170,N_13162,N_14781);
nand U19171 (N_19171,N_13641,N_10164);
nor U19172 (N_19172,N_13973,N_12988);
nand U19173 (N_19173,N_10516,N_11748);
nand U19174 (N_19174,N_13347,N_12115);
xnor U19175 (N_19175,N_12509,N_14437);
nand U19176 (N_19176,N_14653,N_12883);
and U19177 (N_19177,N_10294,N_14977);
nand U19178 (N_19178,N_10449,N_11634);
nand U19179 (N_19179,N_13184,N_12266);
and U19180 (N_19180,N_12860,N_12270);
and U19181 (N_19181,N_14554,N_12434);
nand U19182 (N_19182,N_13268,N_12971);
and U19183 (N_19183,N_13468,N_12990);
and U19184 (N_19184,N_13223,N_14868);
nand U19185 (N_19185,N_12027,N_11158);
xnor U19186 (N_19186,N_14441,N_14213);
and U19187 (N_19187,N_10196,N_12576);
or U19188 (N_19188,N_11247,N_14716);
nand U19189 (N_19189,N_10859,N_14342);
or U19190 (N_19190,N_12229,N_12507);
nor U19191 (N_19191,N_10172,N_13338);
and U19192 (N_19192,N_13396,N_11466);
or U19193 (N_19193,N_13392,N_11642);
nand U19194 (N_19194,N_12988,N_14675);
nor U19195 (N_19195,N_14841,N_12951);
or U19196 (N_19196,N_10626,N_14148);
nor U19197 (N_19197,N_12680,N_14400);
nor U19198 (N_19198,N_12465,N_14949);
nor U19199 (N_19199,N_11367,N_14468);
nand U19200 (N_19200,N_11626,N_13838);
and U19201 (N_19201,N_14184,N_10144);
nor U19202 (N_19202,N_12540,N_11079);
nand U19203 (N_19203,N_10174,N_12645);
nand U19204 (N_19204,N_14568,N_10786);
nor U19205 (N_19205,N_10113,N_10364);
nor U19206 (N_19206,N_13841,N_13383);
xor U19207 (N_19207,N_10047,N_10714);
and U19208 (N_19208,N_11952,N_10463);
and U19209 (N_19209,N_10192,N_10788);
nand U19210 (N_19210,N_13283,N_13432);
nor U19211 (N_19211,N_13942,N_13766);
nand U19212 (N_19212,N_13246,N_14113);
and U19213 (N_19213,N_14334,N_10498);
nor U19214 (N_19214,N_13197,N_14626);
or U19215 (N_19215,N_13824,N_11781);
nor U19216 (N_19216,N_13628,N_10444);
or U19217 (N_19217,N_11136,N_14639);
nand U19218 (N_19218,N_12972,N_13456);
and U19219 (N_19219,N_11877,N_11872);
nand U19220 (N_19220,N_14374,N_11922);
nor U19221 (N_19221,N_12408,N_11978);
nor U19222 (N_19222,N_11364,N_13470);
nor U19223 (N_19223,N_12356,N_13439);
nand U19224 (N_19224,N_13557,N_11033);
nand U19225 (N_19225,N_12199,N_11360);
and U19226 (N_19226,N_11809,N_12967);
nand U19227 (N_19227,N_12524,N_13535);
nand U19228 (N_19228,N_10402,N_12730);
or U19229 (N_19229,N_13740,N_14397);
and U19230 (N_19230,N_10035,N_14481);
nand U19231 (N_19231,N_13973,N_11339);
and U19232 (N_19232,N_14108,N_11781);
or U19233 (N_19233,N_11621,N_11267);
and U19234 (N_19234,N_13631,N_14696);
or U19235 (N_19235,N_13610,N_12934);
nor U19236 (N_19236,N_14672,N_10961);
nor U19237 (N_19237,N_12129,N_12204);
nand U19238 (N_19238,N_12083,N_14984);
xor U19239 (N_19239,N_14161,N_12719);
or U19240 (N_19240,N_14399,N_10859);
nor U19241 (N_19241,N_12236,N_14122);
xor U19242 (N_19242,N_11684,N_10565);
or U19243 (N_19243,N_13187,N_13396);
or U19244 (N_19244,N_13677,N_13706);
or U19245 (N_19245,N_14459,N_13610);
or U19246 (N_19246,N_11797,N_13718);
nand U19247 (N_19247,N_11791,N_13681);
nor U19248 (N_19248,N_12859,N_10884);
nand U19249 (N_19249,N_12109,N_14125);
nand U19250 (N_19250,N_11958,N_12317);
nor U19251 (N_19251,N_13834,N_10032);
nor U19252 (N_19252,N_11996,N_14374);
nand U19253 (N_19253,N_13236,N_12581);
nor U19254 (N_19254,N_12085,N_13911);
nand U19255 (N_19255,N_11460,N_11217);
or U19256 (N_19256,N_10717,N_11260);
nand U19257 (N_19257,N_10235,N_11048);
nand U19258 (N_19258,N_12131,N_10532);
or U19259 (N_19259,N_13080,N_12614);
nand U19260 (N_19260,N_11342,N_13034);
nor U19261 (N_19261,N_10290,N_11933);
and U19262 (N_19262,N_13927,N_10286);
nand U19263 (N_19263,N_10271,N_12737);
nor U19264 (N_19264,N_11359,N_10721);
nand U19265 (N_19265,N_12592,N_12907);
or U19266 (N_19266,N_12676,N_11502);
nor U19267 (N_19267,N_10342,N_13547);
and U19268 (N_19268,N_11661,N_11316);
and U19269 (N_19269,N_10093,N_11471);
and U19270 (N_19270,N_14991,N_12529);
and U19271 (N_19271,N_14842,N_13333);
and U19272 (N_19272,N_11362,N_12373);
and U19273 (N_19273,N_13444,N_12893);
and U19274 (N_19274,N_11877,N_12928);
nand U19275 (N_19275,N_10177,N_12263);
and U19276 (N_19276,N_14977,N_13597);
nor U19277 (N_19277,N_13600,N_10724);
nor U19278 (N_19278,N_14230,N_12345);
xnor U19279 (N_19279,N_10418,N_12639);
and U19280 (N_19280,N_11019,N_11853);
nor U19281 (N_19281,N_11932,N_13183);
or U19282 (N_19282,N_10365,N_13806);
or U19283 (N_19283,N_10538,N_12080);
and U19284 (N_19284,N_14664,N_11358);
and U19285 (N_19285,N_10155,N_11342);
xnor U19286 (N_19286,N_14846,N_14969);
nand U19287 (N_19287,N_13448,N_14217);
nor U19288 (N_19288,N_10092,N_10980);
nand U19289 (N_19289,N_11139,N_13814);
and U19290 (N_19290,N_13875,N_14069);
or U19291 (N_19291,N_13441,N_14588);
nor U19292 (N_19292,N_10871,N_11586);
xor U19293 (N_19293,N_14009,N_14422);
nor U19294 (N_19294,N_11769,N_13463);
or U19295 (N_19295,N_13583,N_14774);
nand U19296 (N_19296,N_14711,N_12439);
or U19297 (N_19297,N_10529,N_14003);
nand U19298 (N_19298,N_10065,N_14045);
or U19299 (N_19299,N_10810,N_13160);
nor U19300 (N_19300,N_13443,N_14231);
and U19301 (N_19301,N_10492,N_14677);
nor U19302 (N_19302,N_14230,N_14384);
and U19303 (N_19303,N_10641,N_14411);
and U19304 (N_19304,N_11088,N_13548);
nor U19305 (N_19305,N_11154,N_14331);
nand U19306 (N_19306,N_14244,N_12274);
or U19307 (N_19307,N_11844,N_11790);
nand U19308 (N_19308,N_14560,N_11188);
and U19309 (N_19309,N_12820,N_14674);
or U19310 (N_19310,N_13853,N_10540);
nor U19311 (N_19311,N_13361,N_13614);
or U19312 (N_19312,N_11307,N_11397);
nand U19313 (N_19313,N_12050,N_14636);
and U19314 (N_19314,N_14450,N_14180);
or U19315 (N_19315,N_12232,N_11760);
nor U19316 (N_19316,N_14290,N_11897);
or U19317 (N_19317,N_11737,N_14008);
or U19318 (N_19318,N_12168,N_14712);
and U19319 (N_19319,N_13042,N_14123);
nor U19320 (N_19320,N_14607,N_10387);
nand U19321 (N_19321,N_11691,N_13950);
nand U19322 (N_19322,N_10701,N_13809);
and U19323 (N_19323,N_10139,N_12562);
nand U19324 (N_19324,N_13272,N_10911);
nand U19325 (N_19325,N_14625,N_11641);
or U19326 (N_19326,N_12370,N_14072);
xor U19327 (N_19327,N_13759,N_10015);
or U19328 (N_19328,N_13912,N_10669);
nor U19329 (N_19329,N_14538,N_13233);
or U19330 (N_19330,N_10227,N_12947);
nor U19331 (N_19331,N_12955,N_12316);
nor U19332 (N_19332,N_12408,N_13145);
and U19333 (N_19333,N_11086,N_14719);
and U19334 (N_19334,N_10882,N_10301);
or U19335 (N_19335,N_10590,N_11523);
and U19336 (N_19336,N_11552,N_14982);
nand U19337 (N_19337,N_11099,N_11882);
or U19338 (N_19338,N_13261,N_12269);
nor U19339 (N_19339,N_12998,N_11565);
nand U19340 (N_19340,N_12531,N_11884);
and U19341 (N_19341,N_10707,N_11940);
and U19342 (N_19342,N_10139,N_12842);
nor U19343 (N_19343,N_12324,N_14597);
or U19344 (N_19344,N_10703,N_10420);
or U19345 (N_19345,N_11015,N_14665);
nand U19346 (N_19346,N_12278,N_14296);
nand U19347 (N_19347,N_13586,N_14236);
nand U19348 (N_19348,N_10458,N_10069);
nand U19349 (N_19349,N_13844,N_10445);
nand U19350 (N_19350,N_14202,N_12077);
nand U19351 (N_19351,N_11664,N_10331);
or U19352 (N_19352,N_11058,N_12969);
nor U19353 (N_19353,N_12274,N_11159);
nor U19354 (N_19354,N_12912,N_10126);
nor U19355 (N_19355,N_14166,N_10092);
nor U19356 (N_19356,N_11126,N_10823);
or U19357 (N_19357,N_10202,N_11157);
nor U19358 (N_19358,N_10818,N_10582);
nor U19359 (N_19359,N_14749,N_13503);
nand U19360 (N_19360,N_14927,N_12869);
or U19361 (N_19361,N_10573,N_10084);
nor U19362 (N_19362,N_11817,N_13417);
nor U19363 (N_19363,N_14336,N_11913);
and U19364 (N_19364,N_10039,N_10000);
and U19365 (N_19365,N_13215,N_12103);
and U19366 (N_19366,N_12071,N_14959);
or U19367 (N_19367,N_14791,N_10546);
and U19368 (N_19368,N_13308,N_14706);
nand U19369 (N_19369,N_14250,N_10981);
or U19370 (N_19370,N_12486,N_14091);
nand U19371 (N_19371,N_13565,N_12815);
and U19372 (N_19372,N_10946,N_10963);
and U19373 (N_19373,N_13094,N_14589);
and U19374 (N_19374,N_13869,N_14308);
and U19375 (N_19375,N_14375,N_13140);
nor U19376 (N_19376,N_11199,N_14939);
xor U19377 (N_19377,N_14476,N_12047);
or U19378 (N_19378,N_11871,N_11791);
and U19379 (N_19379,N_14542,N_11076);
or U19380 (N_19380,N_11535,N_14876);
nor U19381 (N_19381,N_13066,N_12936);
nand U19382 (N_19382,N_11295,N_10186);
or U19383 (N_19383,N_14577,N_14538);
and U19384 (N_19384,N_12712,N_11350);
and U19385 (N_19385,N_11644,N_11415);
or U19386 (N_19386,N_11727,N_12609);
and U19387 (N_19387,N_10976,N_14392);
nand U19388 (N_19388,N_13624,N_13284);
nand U19389 (N_19389,N_10830,N_11772);
or U19390 (N_19390,N_11602,N_12873);
or U19391 (N_19391,N_10171,N_12520);
nor U19392 (N_19392,N_12967,N_14213);
and U19393 (N_19393,N_10280,N_11623);
or U19394 (N_19394,N_12544,N_11076);
xnor U19395 (N_19395,N_13178,N_12850);
or U19396 (N_19396,N_14866,N_13714);
nor U19397 (N_19397,N_13842,N_10679);
nor U19398 (N_19398,N_11767,N_14559);
nand U19399 (N_19399,N_12805,N_11601);
and U19400 (N_19400,N_14649,N_13878);
nor U19401 (N_19401,N_14817,N_11361);
or U19402 (N_19402,N_12886,N_13811);
nor U19403 (N_19403,N_12624,N_14470);
nor U19404 (N_19404,N_14945,N_13419);
or U19405 (N_19405,N_10990,N_14566);
or U19406 (N_19406,N_10969,N_13770);
nor U19407 (N_19407,N_13125,N_14334);
and U19408 (N_19408,N_13526,N_14355);
or U19409 (N_19409,N_12903,N_13896);
and U19410 (N_19410,N_14622,N_14090);
nand U19411 (N_19411,N_14413,N_13591);
and U19412 (N_19412,N_13854,N_12211);
or U19413 (N_19413,N_12195,N_12235);
nand U19414 (N_19414,N_14636,N_11679);
nor U19415 (N_19415,N_14326,N_11431);
nand U19416 (N_19416,N_11849,N_14861);
nor U19417 (N_19417,N_10698,N_10560);
and U19418 (N_19418,N_11138,N_10814);
or U19419 (N_19419,N_12027,N_11120);
nand U19420 (N_19420,N_13130,N_10240);
and U19421 (N_19421,N_13468,N_10270);
nor U19422 (N_19422,N_10131,N_10395);
or U19423 (N_19423,N_14830,N_13556);
nor U19424 (N_19424,N_10520,N_14748);
or U19425 (N_19425,N_14754,N_13972);
or U19426 (N_19426,N_14973,N_13195);
or U19427 (N_19427,N_14475,N_12723);
nand U19428 (N_19428,N_10680,N_13391);
and U19429 (N_19429,N_11033,N_12145);
and U19430 (N_19430,N_13360,N_10014);
nor U19431 (N_19431,N_13052,N_11277);
nor U19432 (N_19432,N_14357,N_10789);
or U19433 (N_19433,N_14586,N_12235);
and U19434 (N_19434,N_10948,N_13204);
nand U19435 (N_19435,N_13439,N_14361);
or U19436 (N_19436,N_14970,N_12252);
and U19437 (N_19437,N_11938,N_14221);
and U19438 (N_19438,N_13148,N_14040);
or U19439 (N_19439,N_14086,N_10143);
nand U19440 (N_19440,N_14250,N_10177);
or U19441 (N_19441,N_14346,N_14418);
or U19442 (N_19442,N_10940,N_13066);
xor U19443 (N_19443,N_13786,N_13572);
nor U19444 (N_19444,N_12742,N_11225);
and U19445 (N_19445,N_14934,N_11469);
and U19446 (N_19446,N_11960,N_13233);
or U19447 (N_19447,N_10082,N_10413);
or U19448 (N_19448,N_14441,N_12409);
nor U19449 (N_19449,N_13594,N_13079);
and U19450 (N_19450,N_10000,N_12567);
and U19451 (N_19451,N_10957,N_14236);
or U19452 (N_19452,N_11918,N_12845);
nand U19453 (N_19453,N_11432,N_12185);
nand U19454 (N_19454,N_13624,N_13388);
or U19455 (N_19455,N_14652,N_13942);
and U19456 (N_19456,N_12430,N_14730);
and U19457 (N_19457,N_14788,N_12092);
xor U19458 (N_19458,N_12371,N_12580);
or U19459 (N_19459,N_14946,N_14509);
and U19460 (N_19460,N_10851,N_10503);
nor U19461 (N_19461,N_11180,N_11059);
or U19462 (N_19462,N_12897,N_13990);
or U19463 (N_19463,N_13712,N_11504);
nand U19464 (N_19464,N_10105,N_14772);
xor U19465 (N_19465,N_12451,N_13071);
and U19466 (N_19466,N_13116,N_14628);
nand U19467 (N_19467,N_13103,N_11178);
and U19468 (N_19468,N_14545,N_10321);
nor U19469 (N_19469,N_13575,N_12158);
nand U19470 (N_19470,N_10584,N_10990);
nor U19471 (N_19471,N_14625,N_10781);
or U19472 (N_19472,N_13278,N_13084);
and U19473 (N_19473,N_11602,N_11389);
or U19474 (N_19474,N_11095,N_13401);
nor U19475 (N_19475,N_12380,N_10380);
and U19476 (N_19476,N_11309,N_11440);
and U19477 (N_19477,N_12493,N_13357);
nor U19478 (N_19478,N_11190,N_10183);
or U19479 (N_19479,N_12630,N_13680);
nor U19480 (N_19480,N_11696,N_12615);
nor U19481 (N_19481,N_11530,N_13352);
and U19482 (N_19482,N_11156,N_11090);
and U19483 (N_19483,N_13304,N_14478);
or U19484 (N_19484,N_12461,N_13808);
and U19485 (N_19485,N_11530,N_10194);
and U19486 (N_19486,N_12308,N_13966);
nor U19487 (N_19487,N_14198,N_13213);
nor U19488 (N_19488,N_12222,N_14749);
or U19489 (N_19489,N_14241,N_13472);
and U19490 (N_19490,N_13222,N_13143);
nand U19491 (N_19491,N_10409,N_12586);
and U19492 (N_19492,N_14957,N_13106);
and U19493 (N_19493,N_12039,N_11563);
nor U19494 (N_19494,N_12909,N_13771);
nand U19495 (N_19495,N_12259,N_10299);
nand U19496 (N_19496,N_12168,N_14438);
or U19497 (N_19497,N_11916,N_10084);
and U19498 (N_19498,N_12785,N_14634);
and U19499 (N_19499,N_12372,N_11195);
and U19500 (N_19500,N_13676,N_10019);
or U19501 (N_19501,N_12964,N_12745);
and U19502 (N_19502,N_11867,N_10786);
nor U19503 (N_19503,N_13564,N_12702);
or U19504 (N_19504,N_14775,N_12959);
nor U19505 (N_19505,N_11135,N_12006);
nor U19506 (N_19506,N_11082,N_14270);
nor U19507 (N_19507,N_11154,N_12577);
nor U19508 (N_19508,N_10406,N_10888);
or U19509 (N_19509,N_14119,N_13448);
and U19510 (N_19510,N_13019,N_11586);
or U19511 (N_19511,N_13275,N_13438);
nand U19512 (N_19512,N_11601,N_14651);
nand U19513 (N_19513,N_11145,N_10108);
and U19514 (N_19514,N_14173,N_14599);
nor U19515 (N_19515,N_10143,N_14969);
nor U19516 (N_19516,N_11981,N_12824);
nor U19517 (N_19517,N_10846,N_13999);
and U19518 (N_19518,N_10254,N_14532);
or U19519 (N_19519,N_10190,N_13221);
nand U19520 (N_19520,N_11672,N_10738);
or U19521 (N_19521,N_14815,N_13549);
nand U19522 (N_19522,N_13366,N_11897);
and U19523 (N_19523,N_13553,N_13882);
and U19524 (N_19524,N_10151,N_13783);
nor U19525 (N_19525,N_10737,N_13959);
nor U19526 (N_19526,N_11081,N_13661);
nor U19527 (N_19527,N_12000,N_14899);
nand U19528 (N_19528,N_10006,N_10940);
nor U19529 (N_19529,N_10667,N_13142);
or U19530 (N_19530,N_11187,N_10084);
and U19531 (N_19531,N_11137,N_14033);
and U19532 (N_19532,N_10795,N_11907);
nand U19533 (N_19533,N_13882,N_10637);
nand U19534 (N_19534,N_11501,N_11181);
or U19535 (N_19535,N_11374,N_10893);
nor U19536 (N_19536,N_12410,N_13928);
xor U19537 (N_19537,N_13965,N_11538);
xor U19538 (N_19538,N_10866,N_10414);
nand U19539 (N_19539,N_12072,N_10804);
nor U19540 (N_19540,N_12434,N_11721);
xor U19541 (N_19541,N_13712,N_13379);
nand U19542 (N_19542,N_11517,N_10563);
and U19543 (N_19543,N_11158,N_10323);
and U19544 (N_19544,N_12701,N_10798);
or U19545 (N_19545,N_13494,N_14819);
and U19546 (N_19546,N_12167,N_11085);
and U19547 (N_19547,N_13098,N_11068);
nor U19548 (N_19548,N_10603,N_11249);
nor U19549 (N_19549,N_11447,N_10363);
nor U19550 (N_19550,N_12288,N_12201);
nor U19551 (N_19551,N_13769,N_13995);
and U19552 (N_19552,N_10892,N_14109);
nor U19553 (N_19553,N_12427,N_13332);
nand U19554 (N_19554,N_12785,N_13276);
nand U19555 (N_19555,N_12915,N_10610);
nor U19556 (N_19556,N_12059,N_12074);
xor U19557 (N_19557,N_10220,N_13703);
nand U19558 (N_19558,N_14212,N_10613);
or U19559 (N_19559,N_10115,N_11646);
nand U19560 (N_19560,N_13523,N_10263);
nor U19561 (N_19561,N_11782,N_10697);
and U19562 (N_19562,N_13726,N_11710);
or U19563 (N_19563,N_13628,N_13900);
nor U19564 (N_19564,N_14865,N_10050);
and U19565 (N_19565,N_11979,N_10130);
and U19566 (N_19566,N_10874,N_13120);
nor U19567 (N_19567,N_14409,N_13346);
nor U19568 (N_19568,N_11668,N_14042);
or U19569 (N_19569,N_13215,N_13076);
nand U19570 (N_19570,N_11891,N_13658);
and U19571 (N_19571,N_13669,N_12705);
nand U19572 (N_19572,N_10413,N_14624);
or U19573 (N_19573,N_12681,N_12428);
nor U19574 (N_19574,N_12718,N_11124);
or U19575 (N_19575,N_11434,N_14743);
nand U19576 (N_19576,N_12293,N_11525);
nor U19577 (N_19577,N_10316,N_14032);
and U19578 (N_19578,N_13318,N_11635);
or U19579 (N_19579,N_12716,N_14678);
nor U19580 (N_19580,N_11850,N_14934);
nor U19581 (N_19581,N_10602,N_10012);
and U19582 (N_19582,N_11630,N_10737);
nor U19583 (N_19583,N_14847,N_14888);
nand U19584 (N_19584,N_12193,N_10872);
nand U19585 (N_19585,N_11560,N_10090);
nand U19586 (N_19586,N_13432,N_13784);
nand U19587 (N_19587,N_12935,N_13827);
nor U19588 (N_19588,N_12275,N_14566);
and U19589 (N_19589,N_12321,N_10597);
or U19590 (N_19590,N_10291,N_12867);
nor U19591 (N_19591,N_14078,N_13570);
and U19592 (N_19592,N_11883,N_11719);
nand U19593 (N_19593,N_12579,N_11347);
nor U19594 (N_19594,N_12651,N_12726);
and U19595 (N_19595,N_10246,N_14064);
nor U19596 (N_19596,N_11395,N_14178);
and U19597 (N_19597,N_10413,N_12802);
or U19598 (N_19598,N_11447,N_14634);
and U19599 (N_19599,N_14075,N_11883);
or U19600 (N_19600,N_13599,N_13038);
or U19601 (N_19601,N_14361,N_10309);
nand U19602 (N_19602,N_10917,N_14611);
xor U19603 (N_19603,N_12819,N_12502);
xnor U19604 (N_19604,N_10180,N_14509);
and U19605 (N_19605,N_10574,N_14430);
nand U19606 (N_19606,N_14778,N_12988);
and U19607 (N_19607,N_12118,N_11270);
and U19608 (N_19608,N_12499,N_13720);
nand U19609 (N_19609,N_14836,N_13827);
and U19610 (N_19610,N_10854,N_10797);
and U19611 (N_19611,N_11378,N_13084);
and U19612 (N_19612,N_14986,N_12101);
or U19613 (N_19613,N_13144,N_14039);
and U19614 (N_19614,N_12402,N_14533);
or U19615 (N_19615,N_14632,N_12225);
nand U19616 (N_19616,N_13462,N_14509);
nand U19617 (N_19617,N_12889,N_10441);
nor U19618 (N_19618,N_12739,N_13531);
or U19619 (N_19619,N_14660,N_11926);
or U19620 (N_19620,N_13066,N_14625);
nand U19621 (N_19621,N_10123,N_12040);
nor U19622 (N_19622,N_12278,N_12879);
or U19623 (N_19623,N_12287,N_11894);
and U19624 (N_19624,N_14056,N_10664);
or U19625 (N_19625,N_12674,N_10095);
and U19626 (N_19626,N_14312,N_10742);
nor U19627 (N_19627,N_14070,N_11683);
and U19628 (N_19628,N_13448,N_10263);
nor U19629 (N_19629,N_13933,N_12403);
nand U19630 (N_19630,N_10083,N_13445);
nor U19631 (N_19631,N_13094,N_14763);
nor U19632 (N_19632,N_11054,N_10188);
nand U19633 (N_19633,N_13811,N_14376);
nor U19634 (N_19634,N_12195,N_14801);
nand U19635 (N_19635,N_10389,N_10058);
nor U19636 (N_19636,N_11915,N_10524);
nand U19637 (N_19637,N_10842,N_14278);
nand U19638 (N_19638,N_11886,N_11087);
or U19639 (N_19639,N_12726,N_12657);
and U19640 (N_19640,N_10232,N_10017);
or U19641 (N_19641,N_11741,N_12099);
or U19642 (N_19642,N_14565,N_10100);
nand U19643 (N_19643,N_12296,N_10821);
nor U19644 (N_19644,N_13443,N_12324);
nand U19645 (N_19645,N_14202,N_14490);
nand U19646 (N_19646,N_14562,N_10206);
nand U19647 (N_19647,N_13498,N_14064);
or U19648 (N_19648,N_11458,N_12623);
or U19649 (N_19649,N_11113,N_12872);
or U19650 (N_19650,N_13672,N_13396);
nand U19651 (N_19651,N_11513,N_10604);
and U19652 (N_19652,N_12419,N_10382);
or U19653 (N_19653,N_10662,N_14520);
or U19654 (N_19654,N_10468,N_13922);
and U19655 (N_19655,N_10563,N_13970);
nand U19656 (N_19656,N_11333,N_11484);
or U19657 (N_19657,N_11990,N_11333);
and U19658 (N_19658,N_14873,N_12745);
nand U19659 (N_19659,N_11887,N_12460);
nor U19660 (N_19660,N_13460,N_14014);
nand U19661 (N_19661,N_13246,N_14440);
and U19662 (N_19662,N_12501,N_11723);
and U19663 (N_19663,N_13636,N_13694);
and U19664 (N_19664,N_11324,N_12138);
or U19665 (N_19665,N_10095,N_14107);
and U19666 (N_19666,N_11817,N_13146);
and U19667 (N_19667,N_14547,N_10169);
or U19668 (N_19668,N_10799,N_13104);
or U19669 (N_19669,N_13264,N_12611);
xor U19670 (N_19670,N_11222,N_13936);
or U19671 (N_19671,N_11011,N_13836);
nor U19672 (N_19672,N_11245,N_13327);
nand U19673 (N_19673,N_10612,N_14105);
nor U19674 (N_19674,N_14593,N_14942);
or U19675 (N_19675,N_12520,N_13300);
or U19676 (N_19676,N_11093,N_10785);
and U19677 (N_19677,N_12292,N_12553);
and U19678 (N_19678,N_14030,N_13630);
xor U19679 (N_19679,N_13912,N_14230);
or U19680 (N_19680,N_12633,N_11631);
and U19681 (N_19681,N_10683,N_14166);
or U19682 (N_19682,N_13397,N_12647);
or U19683 (N_19683,N_14280,N_13277);
nand U19684 (N_19684,N_11334,N_14520);
nor U19685 (N_19685,N_12017,N_12757);
nand U19686 (N_19686,N_12570,N_11139);
and U19687 (N_19687,N_13909,N_13782);
nand U19688 (N_19688,N_12974,N_11271);
and U19689 (N_19689,N_11456,N_13123);
nand U19690 (N_19690,N_10081,N_10098);
and U19691 (N_19691,N_14270,N_14246);
and U19692 (N_19692,N_11767,N_11970);
nor U19693 (N_19693,N_14929,N_12500);
nor U19694 (N_19694,N_12143,N_11937);
or U19695 (N_19695,N_10361,N_10481);
and U19696 (N_19696,N_11919,N_12754);
and U19697 (N_19697,N_10789,N_12460);
nor U19698 (N_19698,N_10205,N_11001);
or U19699 (N_19699,N_14514,N_13867);
nand U19700 (N_19700,N_11285,N_11831);
or U19701 (N_19701,N_13769,N_11517);
nor U19702 (N_19702,N_12789,N_11599);
nand U19703 (N_19703,N_11716,N_14283);
and U19704 (N_19704,N_14740,N_14622);
and U19705 (N_19705,N_13945,N_13256);
nand U19706 (N_19706,N_12379,N_11021);
or U19707 (N_19707,N_12395,N_11901);
or U19708 (N_19708,N_14965,N_10461);
nor U19709 (N_19709,N_14281,N_11765);
or U19710 (N_19710,N_10286,N_12355);
nor U19711 (N_19711,N_14936,N_10835);
xnor U19712 (N_19712,N_14607,N_10055);
xnor U19713 (N_19713,N_14510,N_10293);
nand U19714 (N_19714,N_12770,N_13014);
nand U19715 (N_19715,N_12225,N_13798);
nand U19716 (N_19716,N_10495,N_13565);
nor U19717 (N_19717,N_14314,N_13067);
nand U19718 (N_19718,N_11952,N_14606);
xor U19719 (N_19719,N_13160,N_14376);
nor U19720 (N_19720,N_11181,N_11324);
nor U19721 (N_19721,N_10297,N_14917);
nor U19722 (N_19722,N_13050,N_11738);
and U19723 (N_19723,N_13058,N_12234);
or U19724 (N_19724,N_10511,N_11716);
nor U19725 (N_19725,N_10400,N_14373);
or U19726 (N_19726,N_10388,N_12821);
or U19727 (N_19727,N_12905,N_10081);
nand U19728 (N_19728,N_10184,N_11129);
and U19729 (N_19729,N_10408,N_14825);
nor U19730 (N_19730,N_11803,N_10115);
nor U19731 (N_19731,N_12532,N_10413);
and U19732 (N_19732,N_12023,N_13205);
nand U19733 (N_19733,N_11961,N_12017);
nor U19734 (N_19734,N_13135,N_10203);
and U19735 (N_19735,N_11571,N_11714);
nand U19736 (N_19736,N_12248,N_12387);
nand U19737 (N_19737,N_14027,N_12970);
or U19738 (N_19738,N_12761,N_12099);
nand U19739 (N_19739,N_11931,N_11765);
and U19740 (N_19740,N_10875,N_13827);
nand U19741 (N_19741,N_14651,N_10726);
nand U19742 (N_19742,N_13792,N_14995);
and U19743 (N_19743,N_11575,N_13198);
nand U19744 (N_19744,N_14981,N_12176);
and U19745 (N_19745,N_10150,N_10243);
and U19746 (N_19746,N_14611,N_10011);
and U19747 (N_19747,N_14661,N_13970);
and U19748 (N_19748,N_10620,N_10863);
nor U19749 (N_19749,N_13810,N_10260);
nand U19750 (N_19750,N_11678,N_13572);
and U19751 (N_19751,N_14591,N_11524);
and U19752 (N_19752,N_10736,N_13221);
nor U19753 (N_19753,N_10345,N_13685);
or U19754 (N_19754,N_14441,N_11238);
nand U19755 (N_19755,N_13826,N_10640);
nand U19756 (N_19756,N_14691,N_14087);
or U19757 (N_19757,N_13820,N_12538);
nor U19758 (N_19758,N_10646,N_12420);
and U19759 (N_19759,N_11604,N_11551);
nor U19760 (N_19760,N_10421,N_14074);
xor U19761 (N_19761,N_12592,N_13386);
nor U19762 (N_19762,N_13145,N_13166);
and U19763 (N_19763,N_10046,N_10592);
or U19764 (N_19764,N_10095,N_14389);
nor U19765 (N_19765,N_10763,N_13399);
nor U19766 (N_19766,N_10909,N_11177);
xnor U19767 (N_19767,N_11386,N_14697);
and U19768 (N_19768,N_10695,N_11378);
nand U19769 (N_19769,N_13955,N_14195);
nor U19770 (N_19770,N_12130,N_12122);
nor U19771 (N_19771,N_11344,N_10838);
or U19772 (N_19772,N_14422,N_10023);
and U19773 (N_19773,N_10684,N_11216);
and U19774 (N_19774,N_12882,N_10536);
nand U19775 (N_19775,N_12048,N_11610);
nand U19776 (N_19776,N_12636,N_10949);
or U19777 (N_19777,N_10276,N_10707);
and U19778 (N_19778,N_10823,N_10435);
nor U19779 (N_19779,N_11652,N_12821);
and U19780 (N_19780,N_11672,N_10217);
nand U19781 (N_19781,N_12004,N_11812);
and U19782 (N_19782,N_13677,N_11283);
or U19783 (N_19783,N_11001,N_12996);
nand U19784 (N_19784,N_13713,N_11441);
and U19785 (N_19785,N_10679,N_13877);
and U19786 (N_19786,N_11701,N_10258);
nand U19787 (N_19787,N_12234,N_12189);
nand U19788 (N_19788,N_14181,N_14089);
or U19789 (N_19789,N_14510,N_13900);
or U19790 (N_19790,N_11306,N_14570);
nand U19791 (N_19791,N_10696,N_14114);
and U19792 (N_19792,N_13107,N_11277);
and U19793 (N_19793,N_14913,N_11392);
nor U19794 (N_19794,N_13190,N_10708);
nor U19795 (N_19795,N_14601,N_14908);
or U19796 (N_19796,N_10472,N_12821);
and U19797 (N_19797,N_12684,N_12714);
nand U19798 (N_19798,N_14255,N_10497);
or U19799 (N_19799,N_10427,N_13705);
or U19800 (N_19800,N_13950,N_14002);
or U19801 (N_19801,N_11564,N_10890);
and U19802 (N_19802,N_10301,N_12084);
and U19803 (N_19803,N_11647,N_10460);
and U19804 (N_19804,N_13966,N_11129);
nand U19805 (N_19805,N_14818,N_14388);
nor U19806 (N_19806,N_11533,N_13676);
nor U19807 (N_19807,N_11687,N_12807);
nand U19808 (N_19808,N_11577,N_12277);
nand U19809 (N_19809,N_11708,N_12696);
and U19810 (N_19810,N_12339,N_14404);
and U19811 (N_19811,N_14430,N_11889);
nand U19812 (N_19812,N_12341,N_10458);
nand U19813 (N_19813,N_14710,N_11639);
nand U19814 (N_19814,N_10764,N_13452);
and U19815 (N_19815,N_12042,N_10357);
nor U19816 (N_19816,N_10329,N_13416);
or U19817 (N_19817,N_10847,N_14684);
and U19818 (N_19818,N_12301,N_11826);
nor U19819 (N_19819,N_12129,N_11028);
and U19820 (N_19820,N_13158,N_12919);
and U19821 (N_19821,N_12353,N_11948);
and U19822 (N_19822,N_12640,N_11824);
nand U19823 (N_19823,N_12050,N_12049);
nand U19824 (N_19824,N_10556,N_12116);
and U19825 (N_19825,N_12089,N_12845);
or U19826 (N_19826,N_13080,N_10201);
nor U19827 (N_19827,N_13787,N_14614);
nand U19828 (N_19828,N_12949,N_11871);
xnor U19829 (N_19829,N_10608,N_13194);
nor U19830 (N_19830,N_12475,N_10348);
nand U19831 (N_19831,N_13954,N_13810);
xor U19832 (N_19832,N_11736,N_11367);
nand U19833 (N_19833,N_12593,N_14410);
or U19834 (N_19834,N_14905,N_10891);
and U19835 (N_19835,N_11231,N_11723);
nand U19836 (N_19836,N_14084,N_12828);
nand U19837 (N_19837,N_14041,N_13757);
nor U19838 (N_19838,N_14965,N_13185);
and U19839 (N_19839,N_12153,N_12704);
and U19840 (N_19840,N_10499,N_14787);
nand U19841 (N_19841,N_12790,N_14346);
nand U19842 (N_19842,N_14256,N_12439);
nor U19843 (N_19843,N_10099,N_11607);
or U19844 (N_19844,N_13529,N_12145);
nand U19845 (N_19845,N_12655,N_11372);
nor U19846 (N_19846,N_10258,N_11021);
and U19847 (N_19847,N_14307,N_10161);
and U19848 (N_19848,N_14212,N_12191);
and U19849 (N_19849,N_11503,N_12576);
nand U19850 (N_19850,N_12755,N_10716);
nor U19851 (N_19851,N_11143,N_13542);
nand U19852 (N_19852,N_12162,N_12458);
nand U19853 (N_19853,N_10867,N_10821);
nand U19854 (N_19854,N_10915,N_13671);
nand U19855 (N_19855,N_12782,N_13551);
nand U19856 (N_19856,N_10605,N_10892);
nand U19857 (N_19857,N_14903,N_10446);
nor U19858 (N_19858,N_14967,N_12417);
nor U19859 (N_19859,N_11900,N_14257);
or U19860 (N_19860,N_12775,N_10402);
or U19861 (N_19861,N_13539,N_14973);
or U19862 (N_19862,N_12956,N_10439);
and U19863 (N_19863,N_10783,N_11673);
and U19864 (N_19864,N_12811,N_10541);
or U19865 (N_19865,N_12303,N_10827);
and U19866 (N_19866,N_11327,N_13386);
nor U19867 (N_19867,N_12069,N_12073);
nand U19868 (N_19868,N_12790,N_13027);
or U19869 (N_19869,N_10302,N_10636);
nand U19870 (N_19870,N_14841,N_12301);
or U19871 (N_19871,N_14881,N_13254);
nand U19872 (N_19872,N_14725,N_11892);
or U19873 (N_19873,N_11033,N_12251);
and U19874 (N_19874,N_10843,N_10102);
or U19875 (N_19875,N_11833,N_10596);
or U19876 (N_19876,N_10681,N_10303);
and U19877 (N_19877,N_12913,N_14465);
nor U19878 (N_19878,N_13951,N_13499);
nor U19879 (N_19879,N_10323,N_13592);
and U19880 (N_19880,N_14469,N_14347);
nor U19881 (N_19881,N_10184,N_10797);
nand U19882 (N_19882,N_14344,N_12185);
nor U19883 (N_19883,N_11735,N_12626);
and U19884 (N_19884,N_13631,N_10629);
or U19885 (N_19885,N_14774,N_10685);
and U19886 (N_19886,N_10391,N_12369);
nor U19887 (N_19887,N_12162,N_14088);
and U19888 (N_19888,N_14320,N_10746);
nand U19889 (N_19889,N_10120,N_12822);
and U19890 (N_19890,N_10521,N_12094);
or U19891 (N_19891,N_12325,N_14142);
or U19892 (N_19892,N_14788,N_12669);
or U19893 (N_19893,N_12417,N_14612);
and U19894 (N_19894,N_10807,N_13573);
or U19895 (N_19895,N_10851,N_10265);
and U19896 (N_19896,N_10682,N_10236);
or U19897 (N_19897,N_13313,N_14576);
and U19898 (N_19898,N_14535,N_14252);
and U19899 (N_19899,N_10039,N_14837);
and U19900 (N_19900,N_14889,N_10397);
or U19901 (N_19901,N_13747,N_11758);
xor U19902 (N_19902,N_10661,N_14183);
nand U19903 (N_19903,N_12695,N_14224);
nor U19904 (N_19904,N_11916,N_11784);
nand U19905 (N_19905,N_14062,N_11407);
or U19906 (N_19906,N_13324,N_11538);
nand U19907 (N_19907,N_10095,N_10449);
nand U19908 (N_19908,N_10103,N_10919);
or U19909 (N_19909,N_13387,N_14623);
and U19910 (N_19910,N_13993,N_13638);
and U19911 (N_19911,N_11214,N_13722);
and U19912 (N_19912,N_10292,N_12989);
and U19913 (N_19913,N_10863,N_12628);
nand U19914 (N_19914,N_10921,N_11470);
nor U19915 (N_19915,N_14763,N_12234);
nand U19916 (N_19916,N_14675,N_13921);
or U19917 (N_19917,N_12200,N_12791);
nand U19918 (N_19918,N_14023,N_11212);
nor U19919 (N_19919,N_10982,N_10510);
and U19920 (N_19920,N_14538,N_11157);
nand U19921 (N_19921,N_14480,N_11034);
or U19922 (N_19922,N_11244,N_12671);
and U19923 (N_19923,N_14714,N_14406);
or U19924 (N_19924,N_13536,N_13444);
nor U19925 (N_19925,N_11926,N_11657);
nor U19926 (N_19926,N_10625,N_11293);
nor U19927 (N_19927,N_10536,N_14791);
nand U19928 (N_19928,N_14626,N_14247);
nand U19929 (N_19929,N_14439,N_14328);
nor U19930 (N_19930,N_14666,N_13785);
nand U19931 (N_19931,N_10736,N_12761);
nand U19932 (N_19932,N_12399,N_11926);
nand U19933 (N_19933,N_12865,N_10659);
or U19934 (N_19934,N_12206,N_13992);
and U19935 (N_19935,N_13558,N_12842);
or U19936 (N_19936,N_13870,N_12928);
and U19937 (N_19937,N_12611,N_13227);
nand U19938 (N_19938,N_13400,N_14261);
nor U19939 (N_19939,N_10811,N_14260);
nand U19940 (N_19940,N_14089,N_14879);
and U19941 (N_19941,N_12973,N_14020);
and U19942 (N_19942,N_10493,N_10510);
xnor U19943 (N_19943,N_13687,N_13274);
and U19944 (N_19944,N_10685,N_10301);
and U19945 (N_19945,N_12326,N_14012);
nand U19946 (N_19946,N_12235,N_14858);
nor U19947 (N_19947,N_12774,N_14298);
or U19948 (N_19948,N_11235,N_10612);
or U19949 (N_19949,N_11085,N_10917);
nand U19950 (N_19950,N_14795,N_13521);
nor U19951 (N_19951,N_14141,N_11662);
or U19952 (N_19952,N_10305,N_13163);
or U19953 (N_19953,N_11307,N_12710);
nor U19954 (N_19954,N_13126,N_10275);
or U19955 (N_19955,N_11382,N_14555);
nor U19956 (N_19956,N_10723,N_12830);
nor U19957 (N_19957,N_13014,N_12197);
or U19958 (N_19958,N_12889,N_14037);
nor U19959 (N_19959,N_13307,N_11799);
nor U19960 (N_19960,N_14647,N_10202);
xor U19961 (N_19961,N_12580,N_13811);
nand U19962 (N_19962,N_10403,N_13739);
nor U19963 (N_19963,N_10959,N_14309);
nor U19964 (N_19964,N_10159,N_10090);
nor U19965 (N_19965,N_14854,N_13351);
and U19966 (N_19966,N_10700,N_13423);
nor U19967 (N_19967,N_12410,N_14043);
nand U19968 (N_19968,N_12396,N_11274);
and U19969 (N_19969,N_11625,N_10034);
nor U19970 (N_19970,N_10461,N_12184);
nor U19971 (N_19971,N_12722,N_10707);
and U19972 (N_19972,N_11443,N_13065);
nor U19973 (N_19973,N_11209,N_13053);
and U19974 (N_19974,N_11241,N_10262);
and U19975 (N_19975,N_13271,N_11778);
nor U19976 (N_19976,N_11050,N_11973);
or U19977 (N_19977,N_12235,N_13385);
nand U19978 (N_19978,N_13206,N_14728);
xnor U19979 (N_19979,N_14872,N_14867);
nand U19980 (N_19980,N_14279,N_13394);
and U19981 (N_19981,N_10889,N_14464);
or U19982 (N_19982,N_10307,N_10962);
or U19983 (N_19983,N_13883,N_14185);
and U19984 (N_19984,N_14312,N_12483);
nand U19985 (N_19985,N_10560,N_12490);
nand U19986 (N_19986,N_13197,N_14352);
or U19987 (N_19987,N_12137,N_11786);
nor U19988 (N_19988,N_13634,N_11404);
nor U19989 (N_19989,N_13808,N_10602);
nand U19990 (N_19990,N_14759,N_14693);
nor U19991 (N_19991,N_10780,N_13713);
or U19992 (N_19992,N_13557,N_10350);
nor U19993 (N_19993,N_14450,N_12104);
nand U19994 (N_19994,N_12785,N_14729);
nor U19995 (N_19995,N_10322,N_13279);
or U19996 (N_19996,N_11951,N_12411);
and U19997 (N_19997,N_13394,N_10511);
nand U19998 (N_19998,N_14992,N_11531);
nand U19999 (N_19999,N_10471,N_10878);
and U20000 (N_20000,N_19424,N_17206);
and U20001 (N_20001,N_17720,N_16391);
nor U20002 (N_20002,N_17901,N_15753);
nor U20003 (N_20003,N_19568,N_17135);
nor U20004 (N_20004,N_15086,N_16570);
nand U20005 (N_20005,N_16525,N_18963);
or U20006 (N_20006,N_16464,N_18526);
nand U20007 (N_20007,N_17384,N_19198);
nor U20008 (N_20008,N_19323,N_15449);
nor U20009 (N_20009,N_18075,N_15723);
nand U20010 (N_20010,N_16226,N_19681);
and U20011 (N_20011,N_19754,N_18096);
and U20012 (N_20012,N_19661,N_15480);
and U20013 (N_20013,N_16383,N_18218);
nor U20014 (N_20014,N_17685,N_17528);
or U20015 (N_20015,N_15100,N_19548);
nand U20016 (N_20016,N_16136,N_16129);
or U20017 (N_20017,N_17480,N_17498);
or U20018 (N_20018,N_15616,N_16470);
nor U20019 (N_20019,N_15475,N_18694);
nand U20020 (N_20020,N_17549,N_15857);
and U20021 (N_20021,N_16177,N_19648);
and U20022 (N_20022,N_15305,N_15945);
nor U20023 (N_20023,N_17648,N_15702);
or U20024 (N_20024,N_18232,N_15694);
nand U20025 (N_20025,N_15301,N_15924);
nor U20026 (N_20026,N_18444,N_19854);
or U20027 (N_20027,N_17620,N_16825);
nor U20028 (N_20028,N_19387,N_15370);
and U20029 (N_20029,N_16860,N_19928);
and U20030 (N_20030,N_17764,N_16764);
nand U20031 (N_20031,N_17338,N_15745);
or U20032 (N_20032,N_15153,N_18280);
or U20033 (N_20033,N_16432,N_19709);
and U20034 (N_20034,N_15986,N_15633);
and U20035 (N_20035,N_17533,N_15018);
nor U20036 (N_20036,N_15619,N_18046);
nor U20037 (N_20037,N_18691,N_15428);
and U20038 (N_20038,N_19159,N_17262);
or U20039 (N_20039,N_18071,N_15941);
nand U20040 (N_20040,N_17220,N_17725);
nand U20041 (N_20041,N_18577,N_15258);
or U20042 (N_20042,N_18150,N_16424);
and U20043 (N_20043,N_19690,N_16593);
nand U20044 (N_20044,N_15617,N_15991);
or U20045 (N_20045,N_18297,N_16133);
nor U20046 (N_20046,N_15295,N_16793);
nand U20047 (N_20047,N_17547,N_18567);
and U20048 (N_20048,N_18951,N_17825);
nand U20049 (N_20049,N_19589,N_17164);
nand U20050 (N_20050,N_15909,N_18665);
nor U20051 (N_20051,N_15858,N_18580);
and U20052 (N_20052,N_15185,N_19465);
nand U20053 (N_20053,N_15077,N_17509);
nor U20054 (N_20054,N_18401,N_16152);
nand U20055 (N_20055,N_18138,N_16228);
and U20056 (N_20056,N_17370,N_16818);
nand U20057 (N_20057,N_15877,N_18782);
nand U20058 (N_20058,N_17123,N_15459);
or U20059 (N_20059,N_18326,N_16655);
or U20060 (N_20060,N_19268,N_18576);
nand U20061 (N_20061,N_19591,N_16477);
xnor U20062 (N_20062,N_17689,N_18914);
nand U20063 (N_20063,N_16043,N_17834);
and U20064 (N_20064,N_16947,N_19535);
and U20065 (N_20065,N_15040,N_15341);
nor U20066 (N_20066,N_18373,N_16552);
nand U20067 (N_20067,N_15698,N_18304);
and U20068 (N_20068,N_15285,N_19992);
or U20069 (N_20069,N_17558,N_15188);
nand U20070 (N_20070,N_18099,N_18014);
or U20071 (N_20071,N_18797,N_18349);
nand U20072 (N_20072,N_17969,N_19788);
nand U20073 (N_20073,N_16255,N_16234);
nand U20074 (N_20074,N_18796,N_17639);
nor U20075 (N_20075,N_17881,N_17068);
and U20076 (N_20076,N_17622,N_15764);
nor U20077 (N_20077,N_17083,N_16911);
nor U20078 (N_20078,N_18406,N_15397);
nor U20079 (N_20079,N_19861,N_18186);
or U20080 (N_20080,N_19726,N_15066);
or U20081 (N_20081,N_17497,N_18662);
nand U20082 (N_20082,N_15042,N_15297);
xor U20083 (N_20083,N_18722,N_15555);
nor U20084 (N_20084,N_15932,N_15596);
nor U20085 (N_20085,N_19066,N_19893);
and U20086 (N_20086,N_17112,N_19354);
nand U20087 (N_20087,N_15179,N_19973);
nor U20088 (N_20088,N_16538,N_15422);
nor U20089 (N_20089,N_19679,N_16758);
and U20090 (N_20090,N_18231,N_15187);
and U20091 (N_20091,N_17682,N_17499);
and U20092 (N_20092,N_17636,N_19881);
and U20093 (N_20093,N_16375,N_15056);
and U20094 (N_20094,N_16091,N_15410);
nor U20095 (N_20095,N_17299,N_18953);
and U20096 (N_20096,N_19674,N_17264);
nor U20097 (N_20097,N_17275,N_18487);
nor U20098 (N_20098,N_17148,N_19031);
nor U20099 (N_20099,N_17715,N_17102);
nor U20100 (N_20100,N_19121,N_15947);
nand U20101 (N_20101,N_17230,N_18791);
or U20102 (N_20102,N_17159,N_18434);
and U20103 (N_20103,N_17623,N_16931);
nor U20104 (N_20104,N_16119,N_16224);
xnor U20105 (N_20105,N_19575,N_15504);
or U20106 (N_20106,N_18975,N_16263);
or U20107 (N_20107,N_16379,N_15780);
xor U20108 (N_20108,N_18435,N_15168);
nor U20109 (N_20109,N_16347,N_19801);
nand U20110 (N_20110,N_15256,N_18621);
and U20111 (N_20111,N_18678,N_19576);
nor U20112 (N_20112,N_16637,N_16123);
nand U20113 (N_20113,N_15752,N_16493);
nand U20114 (N_20114,N_15071,N_19489);
or U20115 (N_20115,N_16985,N_16285);
nor U20116 (N_20116,N_18421,N_18093);
or U20117 (N_20117,N_15980,N_17696);
or U20118 (N_20118,N_15244,N_19889);
and U20119 (N_20119,N_17386,N_17035);
xnor U20120 (N_20120,N_19014,N_16395);
and U20121 (N_20121,N_19175,N_18635);
or U20122 (N_20122,N_15070,N_18419);
xnor U20123 (N_20123,N_15224,N_15750);
nor U20124 (N_20124,N_19902,N_19839);
nand U20125 (N_20125,N_19696,N_16015);
nor U20126 (N_20126,N_18300,N_16067);
nand U20127 (N_20127,N_19356,N_19860);
nor U20128 (N_20128,N_16856,N_19852);
nor U20129 (N_20129,N_15448,N_18536);
nor U20130 (N_20130,N_19638,N_15695);
or U20131 (N_20131,N_17291,N_15242);
nor U20132 (N_20132,N_15769,N_16438);
or U20133 (N_20133,N_17144,N_16559);
nand U20134 (N_20134,N_16926,N_16474);
or U20135 (N_20135,N_15704,N_15593);
nand U20136 (N_20136,N_15240,N_16631);
nand U20137 (N_20137,N_18780,N_19780);
or U20138 (N_20138,N_15574,N_18115);
nand U20139 (N_20139,N_15349,N_17310);
or U20140 (N_20140,N_15784,N_19764);
nor U20141 (N_20141,N_18196,N_18831);
nand U20142 (N_20142,N_17548,N_15110);
or U20143 (N_20143,N_19233,N_18517);
nor U20144 (N_20144,N_16394,N_18820);
nand U20145 (N_20145,N_16299,N_18067);
or U20146 (N_20146,N_17566,N_16690);
or U20147 (N_20147,N_18396,N_15530);
or U20148 (N_20148,N_16699,N_17846);
nor U20149 (N_20149,N_16501,N_19436);
nand U20150 (N_20150,N_15966,N_15908);
and U20151 (N_20151,N_19484,N_18054);
or U20152 (N_20152,N_18399,N_15145);
and U20153 (N_20153,N_15847,N_18497);
or U20154 (N_20154,N_17772,N_16960);
and U20155 (N_20155,N_18660,N_17941);
nand U20156 (N_20156,N_18763,N_16280);
nand U20157 (N_20157,N_15853,N_16336);
nand U20158 (N_20158,N_17302,N_19834);
nor U20159 (N_20159,N_18141,N_19459);
and U20160 (N_20160,N_19285,N_19182);
and U20161 (N_20161,N_19110,N_15737);
nand U20162 (N_20162,N_16420,N_18769);
and U20163 (N_20163,N_15304,N_15231);
and U20164 (N_20164,N_17329,N_17245);
and U20165 (N_20165,N_18155,N_15293);
nor U20166 (N_20166,N_18704,N_17002);
or U20167 (N_20167,N_16198,N_17237);
and U20168 (N_20168,N_19993,N_15507);
nand U20169 (N_20169,N_17782,N_16784);
nor U20170 (N_20170,N_16385,N_18184);
nand U20171 (N_20171,N_16717,N_15629);
nor U20172 (N_20172,N_16109,N_16589);
and U20173 (N_20173,N_18047,N_17292);
nor U20174 (N_20174,N_17960,N_18857);
nor U20175 (N_20175,N_17356,N_19400);
nand U20176 (N_20176,N_16791,N_15717);
nand U20177 (N_20177,N_15866,N_17057);
nand U20178 (N_20178,N_16542,N_18625);
nand U20179 (N_20179,N_19539,N_19134);
and U20180 (N_20180,N_15862,N_18659);
and U20181 (N_20181,N_19294,N_16075);
or U20182 (N_20182,N_19776,N_17693);
or U20183 (N_20183,N_19064,N_16135);
nand U20184 (N_20184,N_15691,N_19030);
nand U20185 (N_20185,N_16756,N_17223);
or U20186 (N_20186,N_18516,N_15097);
or U20187 (N_20187,N_18412,N_16881);
nor U20188 (N_20188,N_18031,N_19440);
nand U20189 (N_20189,N_18732,N_18420);
nand U20190 (N_20190,N_16629,N_16688);
and U20191 (N_20191,N_19841,N_18139);
nor U20192 (N_20192,N_17698,N_16889);
and U20193 (N_20193,N_18165,N_15204);
and U20194 (N_20194,N_18018,N_17400);
nand U20195 (N_20195,N_15514,N_16610);
and U20196 (N_20196,N_16476,N_17633);
nor U20197 (N_20197,N_18823,N_16130);
and U20198 (N_20198,N_16310,N_17768);
and U20199 (N_20199,N_18927,N_17086);
nor U20200 (N_20200,N_16929,N_15130);
nor U20201 (N_20201,N_19366,N_18249);
and U20202 (N_20202,N_18631,N_18573);
and U20203 (N_20203,N_19847,N_19891);
nor U20204 (N_20204,N_19451,N_15521);
nand U20205 (N_20205,N_17081,N_15103);
or U20206 (N_20206,N_17402,N_19107);
and U20207 (N_20207,N_15218,N_19678);
nor U20208 (N_20208,N_15848,N_18575);
or U20209 (N_20209,N_16617,N_16058);
nand U20210 (N_20210,N_16846,N_19136);
or U20211 (N_20211,N_19078,N_17465);
or U20212 (N_20212,N_15815,N_18158);
xnor U20213 (N_20213,N_19099,N_17198);
or U20214 (N_20214,N_17712,N_15518);
nand U20215 (N_20215,N_15875,N_18239);
or U20216 (N_20216,N_17185,N_18889);
or U20217 (N_20217,N_16319,N_18759);
nor U20218 (N_20218,N_19607,N_15373);
and U20219 (N_20219,N_19037,N_18008);
or U20220 (N_20220,N_17048,N_17030);
nor U20221 (N_20221,N_15257,N_15113);
and U20222 (N_20222,N_18070,N_16718);
nand U20223 (N_20223,N_15385,N_19765);
and U20224 (N_20224,N_19925,N_19739);
or U20225 (N_20225,N_16528,N_16536);
or U20226 (N_20226,N_18990,N_17239);
and U20227 (N_20227,N_17004,N_18157);
or U20228 (N_20228,N_17663,N_18793);
or U20229 (N_20229,N_16546,N_19132);
and U20230 (N_20230,N_16526,N_19442);
and U20231 (N_20231,N_16887,N_18730);
or U20232 (N_20232,N_15824,N_19097);
xor U20233 (N_20233,N_16606,N_15687);
and U20234 (N_20234,N_16973,N_19142);
xor U20235 (N_20235,N_18287,N_18336);
nor U20236 (N_20236,N_16763,N_16754);
and U20237 (N_20237,N_16357,N_17607);
nand U20238 (N_20238,N_17171,N_15332);
or U20239 (N_20239,N_17094,N_18431);
or U20240 (N_20240,N_18168,N_17982);
or U20241 (N_20241,N_15429,N_15860);
and U20242 (N_20242,N_18933,N_18605);
nor U20243 (N_20243,N_16068,N_18306);
or U20244 (N_20244,N_16961,N_18537);
xnor U20245 (N_20245,N_16866,N_19602);
or U20246 (N_20246,N_16706,N_19297);
and U20247 (N_20247,N_17121,N_18883);
and U20248 (N_20248,N_19131,N_16298);
or U20249 (N_20249,N_16668,N_19305);
or U20250 (N_20250,N_17388,N_16425);
nand U20251 (N_20251,N_19370,N_19334);
nand U20252 (N_20252,N_18266,N_16583);
nand U20253 (N_20253,N_19426,N_17863);
or U20254 (N_20254,N_18610,N_15600);
and U20255 (N_20255,N_16809,N_15928);
or U20256 (N_20256,N_19831,N_15522);
and U20257 (N_20257,N_18827,N_15176);
and U20258 (N_20258,N_18807,N_16799);
or U20259 (N_20259,N_19206,N_19051);
nor U20260 (N_20260,N_15300,N_16861);
or U20261 (N_20261,N_19228,N_17426);
nand U20262 (N_20262,N_18585,N_15586);
nand U20263 (N_20263,N_19139,N_16323);
nand U20264 (N_20264,N_16288,N_18522);
nor U20265 (N_20265,N_18225,N_19315);
or U20266 (N_20266,N_15568,N_19542);
nor U20267 (N_20267,N_17677,N_18560);
nand U20268 (N_20268,N_15227,N_15200);
nand U20269 (N_20269,N_18983,N_16871);
nor U20270 (N_20270,N_18657,N_17732);
and U20271 (N_20271,N_19878,N_19406);
or U20272 (N_20272,N_17878,N_18729);
and U20273 (N_20273,N_17832,N_15724);
and U20274 (N_20274,N_17404,N_18481);
and U20275 (N_20275,N_18207,N_15251);
xor U20276 (N_20276,N_15566,N_17563);
nor U20277 (N_20277,N_19615,N_16806);
and U20278 (N_20278,N_15817,N_19324);
nand U20279 (N_20279,N_16019,N_15778);
nor U20280 (N_20280,N_15026,N_16732);
nand U20281 (N_20281,N_17635,N_16267);
nand U20282 (N_20282,N_16485,N_16553);
nand U20283 (N_20283,N_18140,N_18019);
nor U20284 (N_20284,N_18030,N_18501);
or U20285 (N_20285,N_19558,N_19380);
nand U20286 (N_20286,N_19526,N_17103);
or U20287 (N_20287,N_15790,N_16588);
nor U20288 (N_20288,N_16838,N_19649);
and U20289 (N_20289,N_17105,N_18620);
or U20290 (N_20290,N_18252,N_15747);
and U20291 (N_20291,N_15962,N_16697);
or U20292 (N_20292,N_15392,N_18463);
and U20293 (N_20293,N_16657,N_18709);
or U20294 (N_20294,N_15509,N_15033);
or U20295 (N_20295,N_15235,N_15961);
or U20296 (N_20296,N_19572,N_18460);
or U20297 (N_20297,N_19209,N_19769);
or U20298 (N_20298,N_19787,N_16164);
or U20299 (N_20299,N_18080,N_16500);
and U20300 (N_20300,N_15995,N_19812);
or U20301 (N_20301,N_15874,N_19579);
and U20302 (N_20302,N_15431,N_16450);
or U20303 (N_20303,N_18918,N_17947);
or U20304 (N_20304,N_16026,N_19583);
or U20305 (N_20305,N_19501,N_15317);
nor U20306 (N_20306,N_15641,N_18328);
nor U20307 (N_20307,N_17487,N_15309);
and U20308 (N_20308,N_16434,N_19061);
nand U20309 (N_20309,N_17532,N_16498);
or U20310 (N_20310,N_15842,N_17373);
xor U20311 (N_20311,N_15589,N_16696);
and U20312 (N_20312,N_19267,N_17007);
nor U20313 (N_20313,N_19219,N_18959);
nand U20314 (N_20314,N_17330,N_19417);
and U20315 (N_20315,N_19316,N_18826);
or U20316 (N_20316,N_19537,N_19570);
and U20317 (N_20317,N_15579,N_16550);
nand U20318 (N_20318,N_15833,N_15748);
nor U20319 (N_20319,N_19123,N_15976);
and U20320 (N_20320,N_17496,N_18394);
nand U20321 (N_20321,N_18125,N_17080);
nor U20322 (N_20322,N_19389,N_19864);
nand U20323 (N_20323,N_16486,N_15280);
nand U20324 (N_20324,N_16864,N_19924);
nor U20325 (N_20325,N_18204,N_19164);
nor U20326 (N_20326,N_19035,N_16977);
nor U20327 (N_20327,N_18962,N_16539);
or U20328 (N_20328,N_18583,N_16286);
nand U20329 (N_20329,N_16948,N_19898);
and U20330 (N_20330,N_16940,N_18205);
and U20331 (N_20331,N_15794,N_18809);
or U20332 (N_20332,N_19269,N_17321);
nor U20333 (N_20333,N_15831,N_19706);
or U20334 (N_20334,N_19786,N_15358);
or U20335 (N_20335,N_15742,N_19517);
or U20336 (N_20336,N_16331,N_16408);
nand U20337 (N_20337,N_18818,N_19205);
nor U20338 (N_20338,N_16449,N_16895);
nand U20339 (N_20339,N_16236,N_16257);
nand U20340 (N_20340,N_17506,N_16480);
or U20341 (N_20341,N_16937,N_19819);
or U20342 (N_20342,N_18525,N_19922);
nor U20343 (N_20343,N_16175,N_18092);
nand U20344 (N_20344,N_17043,N_19138);
and U20345 (N_20345,N_15744,N_16715);
nor U20346 (N_20346,N_18867,N_16975);
nand U20347 (N_20347,N_15660,N_15163);
nand U20348 (N_20348,N_15871,N_15832);
nand U20349 (N_20349,N_15000,N_18840);
or U20350 (N_20350,N_17414,N_18923);
nand U20351 (N_20351,N_19434,N_15271);
or U20352 (N_20352,N_19995,N_16780);
or U20353 (N_20353,N_16007,N_17805);
or U20354 (N_20354,N_17456,N_15693);
or U20355 (N_20355,N_17613,N_16609);
or U20356 (N_20356,N_18436,N_17348);
or U20357 (N_20357,N_19065,N_19493);
xnor U20358 (N_20358,N_19803,N_15148);
or U20359 (N_20359,N_19951,N_17054);
nor U20360 (N_20360,N_19813,N_15653);
nand U20361 (N_20361,N_19200,N_16191);
or U20362 (N_20362,N_18873,N_18222);
nor U20363 (N_20363,N_16905,N_16436);
or U20364 (N_20364,N_18454,N_18085);
nor U20365 (N_20365,N_16746,N_16206);
nand U20366 (N_20366,N_16906,N_16457);
or U20367 (N_20367,N_18779,N_16579);
and U20368 (N_20368,N_18428,N_18344);
or U20369 (N_20369,N_16810,N_15802);
or U20370 (N_20370,N_15972,N_16046);
or U20371 (N_20371,N_18395,N_16390);
nand U20372 (N_20372,N_15345,N_16030);
nand U20373 (N_20373,N_19608,N_17812);
or U20374 (N_20374,N_16057,N_15846);
nand U20375 (N_20375,N_15347,N_18016);
nor U20376 (N_20376,N_18377,N_17170);
nor U20377 (N_20377,N_16185,N_16915);
nand U20378 (N_20378,N_18050,N_16796);
or U20379 (N_20379,N_17405,N_15914);
nor U20380 (N_20380,N_18183,N_18323);
or U20381 (N_20381,N_18926,N_17576);
or U20382 (N_20382,N_19204,N_15570);
or U20383 (N_20383,N_18281,N_16146);
and U20384 (N_20384,N_18663,N_15039);
nand U20385 (N_20385,N_17991,N_18871);
nor U20386 (N_20386,N_17151,N_17042);
nand U20387 (N_20387,N_17705,N_17443);
or U20388 (N_20388,N_18708,N_15222);
and U20389 (N_20389,N_18864,N_18540);
xor U20390 (N_20390,N_18726,N_16761);
and U20391 (N_20391,N_19859,N_17913);
or U20392 (N_20392,N_19835,N_15709);
nand U20393 (N_20393,N_18211,N_16287);
and U20394 (N_20394,N_15627,N_19603);
and U20395 (N_20395,N_15164,N_19226);
or U20396 (N_20396,N_19309,N_16983);
nand U20397 (N_20397,N_19277,N_18682);
or U20398 (N_20398,N_16909,N_18408);
and U20399 (N_20399,N_19077,N_16828);
xor U20400 (N_20400,N_16956,N_15850);
nor U20401 (N_20401,N_16454,N_19873);
or U20402 (N_20402,N_16523,N_17630);
nand U20403 (N_20403,N_18720,N_17598);
and U20404 (N_20404,N_16644,N_19842);
nand U20405 (N_20405,N_15840,N_15116);
nor U20406 (N_20406,N_16264,N_19740);
nand U20407 (N_20407,N_16031,N_15472);
nand U20408 (N_20408,N_17179,N_15795);
nor U20409 (N_20409,N_18701,N_19783);
nor U20410 (N_20410,N_15444,N_15869);
nor U20411 (N_20411,N_17201,N_15706);
nand U20412 (N_20412,N_16202,N_19668);
or U20413 (N_20413,N_17557,N_15282);
nand U20414 (N_20414,N_17312,N_18478);
and U20415 (N_20415,N_18033,N_18679);
or U20416 (N_20416,N_17126,N_16568);
xnor U20417 (N_20417,N_16064,N_18764);
nor U20418 (N_20418,N_19985,N_18307);
nand U20419 (N_20419,N_16767,N_15361);
nor U20420 (N_20420,N_16775,N_18371);
nor U20421 (N_20421,N_15245,N_16632);
nand U20422 (N_20422,N_17175,N_19704);
nand U20423 (N_20423,N_17062,N_17501);
or U20424 (N_20424,N_17228,N_15788);
nor U20425 (N_20425,N_18044,N_17536);
nor U20426 (N_20426,N_18221,N_15538);
xor U20427 (N_20427,N_15830,N_19251);
nand U20428 (N_20428,N_17606,N_15314);
or U20429 (N_20429,N_17922,N_16343);
nor U20430 (N_20430,N_17395,N_17739);
and U20431 (N_20431,N_19943,N_19724);
nand U20432 (N_20432,N_16330,N_17744);
or U20433 (N_20433,N_18804,N_18579);
nand U20434 (N_20434,N_18913,N_17483);
or U20435 (N_20435,N_15664,N_16415);
nor U20436 (N_20436,N_17318,N_18152);
and U20437 (N_20437,N_17500,N_17104);
or U20438 (N_20438,N_16245,N_18861);
or U20439 (N_20439,N_19283,N_15837);
nor U20440 (N_20440,N_15284,N_15183);
and U20441 (N_20441,N_16088,N_15855);
nand U20442 (N_20442,N_18968,N_16456);
nand U20443 (N_20443,N_17824,N_19475);
nor U20444 (N_20444,N_16592,N_15474);
nand U20445 (N_20445,N_18856,N_16679);
nand U20446 (N_20446,N_19784,N_16188);
nor U20447 (N_20447,N_17628,N_15630);
nand U20448 (N_20448,N_18135,N_17195);
nor U20449 (N_20449,N_16886,N_19553);
nand U20450 (N_20450,N_15469,N_15208);
nor U20451 (N_20451,N_17357,N_16976);
nand U20452 (N_20452,N_16414,N_17671);
and U20453 (N_20453,N_15072,N_15159);
or U20454 (N_20454,N_18107,N_17806);
nor U20455 (N_20455,N_18034,N_18039);
nand U20456 (N_20456,N_19004,N_19116);
xnor U20457 (N_20457,N_15632,N_18228);
or U20458 (N_20458,N_15697,N_15019);
nand U20459 (N_20459,N_15528,N_19443);
or U20460 (N_20460,N_17521,N_17281);
nand U20461 (N_20461,N_16665,N_17013);
or U20462 (N_20462,N_18322,N_15220);
and U20463 (N_20463,N_15733,N_18250);
and U20464 (N_20464,N_19430,N_19849);
nand U20465 (N_20465,N_17000,N_17323);
nand U20466 (N_20466,N_19643,N_17450);
and U20467 (N_20467,N_16630,N_19347);
or U20468 (N_20468,N_16704,N_17877);
nor U20469 (N_20469,N_17778,N_15675);
nand U20470 (N_20470,N_15771,N_19083);
or U20471 (N_20471,N_18242,N_17934);
nand U20472 (N_20472,N_16624,N_18775);
nor U20473 (N_20473,N_15175,N_15290);
nand U20474 (N_20474,N_17714,N_18374);
and U20475 (N_20475,N_18269,N_16356);
and U20476 (N_20476,N_19033,N_15090);
nor U20477 (N_20477,N_18645,N_18234);
nand U20478 (N_20478,N_18197,N_15131);
nand U20479 (N_20479,N_16667,N_17334);
or U20480 (N_20480,N_18619,N_15551);
and U20481 (N_20481,N_18865,N_15174);
or U20482 (N_20482,N_18439,N_16103);
nand U20483 (N_20483,N_16197,N_16124);
or U20484 (N_20484,N_19896,N_17711);
nor U20485 (N_20485,N_16281,N_16824);
or U20486 (N_20486,N_19041,N_19557);
nor U20487 (N_20487,N_17781,N_18899);
nand U20488 (N_20488,N_15982,N_16882);
or U20489 (N_20489,N_18132,N_19223);
or U20490 (N_20490,N_19203,N_16229);
and U20491 (N_20491,N_19516,N_17362);
nand U20492 (N_20492,N_16178,N_19075);
and U20493 (N_20493,N_17853,N_15180);
and U20494 (N_20494,N_19279,N_16673);
and U20495 (N_20495,N_15759,N_17896);
or U20496 (N_20496,N_19897,N_18061);
nand U20497 (N_20497,N_19923,N_17385);
nor U20498 (N_20498,N_16814,N_15648);
nor U20499 (N_20499,N_18987,N_15930);
and U20500 (N_20500,N_17279,N_19042);
or U20501 (N_20501,N_16110,N_15402);
nand U20502 (N_20502,N_16195,N_18145);
nand U20503 (N_20503,N_18052,N_15396);
nor U20504 (N_20504,N_15191,N_16072);
or U20505 (N_20505,N_19773,N_19564);
or U20506 (N_20506,N_16529,N_17192);
nand U20507 (N_20507,N_17784,N_19750);
nor U20508 (N_20508,N_19628,N_17061);
and U20509 (N_20509,N_15523,N_19670);
xnor U20510 (N_20510,N_19730,N_16958);
and U20511 (N_20511,N_16170,N_18534);
nand U20512 (N_20512,N_16627,N_19053);
or U20513 (N_20513,N_16847,N_16974);
nor U20514 (N_20514,N_19733,N_15513);
or U20515 (N_20515,N_15901,N_17326);
or U20516 (N_20516,N_18166,N_17700);
or U20517 (N_20517,N_17572,N_17430);
xnor U20518 (N_20518,N_18542,N_16853);
and U20519 (N_20519,N_15313,N_16509);
nor U20520 (N_20520,N_16218,N_16174);
nor U20521 (N_20521,N_16325,N_19533);
and U20522 (N_20522,N_15192,N_18602);
and U20523 (N_20523,N_16618,N_15956);
nand U20524 (N_20524,N_17656,N_18120);
and U20525 (N_20525,N_17090,N_16795);
nor U20526 (N_20526,N_15059,N_17347);
nand U20527 (N_20527,N_19917,N_17591);
nand U20528 (N_20528,N_16324,N_16180);
and U20529 (N_20529,N_16512,N_18247);
xnor U20530 (N_20530,N_19531,N_15010);
or U20531 (N_20531,N_18649,N_15193);
and U20532 (N_20532,N_18658,N_16510);
and U20533 (N_20533,N_15984,N_18450);
and U20534 (N_20534,N_19016,N_17319);
and U20535 (N_20535,N_17023,N_19474);
and U20536 (N_20536,N_19697,N_18376);
nand U20537 (N_20537,N_18251,N_15604);
and U20538 (N_20538,N_15162,N_19609);
nand U20539 (N_20539,N_19068,N_19098);
or U20540 (N_20540,N_18697,N_18043);
nand U20541 (N_20541,N_17755,N_19384);
and U20542 (N_20542,N_18427,N_15957);
or U20543 (N_20543,N_18528,N_19450);
or U20544 (N_20544,N_15057,N_17133);
nand U20545 (N_20545,N_18193,N_16765);
or U20546 (N_20546,N_19906,N_16161);
nor U20547 (N_20547,N_16837,N_15466);
and U20548 (N_20548,N_16467,N_19000);
and U20549 (N_20549,N_19437,N_18226);
nand U20550 (N_20550,N_17021,N_18206);
nand U20551 (N_20551,N_16942,N_17051);
or U20552 (N_20552,N_17095,N_19463);
nor U20553 (N_20553,N_19676,N_15854);
or U20554 (N_20554,N_16591,N_19409);
nand U20555 (N_20555,N_17939,N_18170);
and U20556 (N_20556,N_18609,N_15092);
nand U20557 (N_20557,N_17132,N_17736);
nand U20558 (N_20558,N_16078,N_16261);
or U20559 (N_20559,N_17336,N_18904);
and U20560 (N_20560,N_19689,N_18646);
or U20561 (N_20561,N_19351,N_19227);
nand U20562 (N_20562,N_16201,N_16563);
nor U20563 (N_20563,N_19371,N_17787);
nand U20564 (N_20564,N_15940,N_19006);
or U20565 (N_20565,N_17452,N_16115);
nor U20566 (N_20566,N_18049,N_16018);
nand U20567 (N_20567,N_19723,N_18341);
nand U20568 (N_20568,N_15864,N_16710);
nand U20569 (N_20569,N_17688,N_18384);
nor U20570 (N_20570,N_18090,N_17129);
nor U20571 (N_20571,N_15563,N_16716);
or U20572 (N_20572,N_19342,N_18130);
nor U20573 (N_20573,N_16469,N_17644);
nand U20574 (N_20574,N_18693,N_17225);
xor U20575 (N_20575,N_19682,N_15420);
nand U20576 (N_20576,N_17217,N_17672);
nand U20577 (N_20577,N_17097,N_15031);
and U20578 (N_20578,N_18946,N_19369);
or U20579 (N_20579,N_18862,N_19588);
xor U20580 (N_20580,N_15997,N_17134);
nor U20581 (N_20581,N_18134,N_19241);
and U20582 (N_20582,N_17332,N_16276);
or U20583 (N_20583,N_15025,N_17811);
and U20584 (N_20584,N_15834,N_15624);
nand U20585 (N_20585,N_16471,N_16647);
and U20586 (N_20586,N_16044,N_19937);
nor U20587 (N_20587,N_15649,N_16441);
nor U20588 (N_20588,N_19288,N_16040);
and U20589 (N_20589,N_19256,N_17455);
nand U20590 (N_20590,N_19632,N_18305);
nor U20591 (N_20591,N_16227,N_16413);
or U20592 (N_20592,N_18642,N_17462);
and U20593 (N_20593,N_18551,N_17482);
and U20594 (N_20594,N_19867,N_15421);
and U20595 (N_20595,N_15254,N_15124);
and U20596 (N_20596,N_17907,N_16640);
or U20597 (N_20597,N_16156,N_18364);
and U20598 (N_20598,N_18668,N_19187);
xor U20599 (N_20599,N_15166,N_17588);
nor U20600 (N_20600,N_18386,N_18562);
xnor U20601 (N_20601,N_16719,N_19795);
nor U20602 (N_20602,N_16004,N_16894);
and U20603 (N_20603,N_17885,N_19524);
and U20604 (N_20604,N_18816,N_15582);
or U20605 (N_20605,N_19817,N_16694);
nor U20606 (N_20606,N_19981,N_16393);
nand U20607 (N_20607,N_19382,N_15094);
and U20608 (N_20608,N_19665,N_16334);
and U20609 (N_20609,N_19652,N_19621);
nor U20610 (N_20610,N_15136,N_19024);
nor U20611 (N_20611,N_15981,N_19586);
and U20612 (N_20612,N_17603,N_19495);
and U20613 (N_20613,N_16590,N_15246);
and U20614 (N_20614,N_16282,N_19892);
nand U20615 (N_20615,N_19270,N_15348);
or U20616 (N_20616,N_15964,N_15949);
nor U20617 (N_20617,N_18728,N_15277);
or U20618 (N_20618,N_17205,N_16835);
nor U20619 (N_20619,N_17382,N_17227);
or U20620 (N_20620,N_19163,N_18843);
or U20621 (N_20621,N_17797,N_16167);
xor U20622 (N_20622,N_15490,N_17944);
nand U20623 (N_20623,N_15440,N_17735);
and U20624 (N_20624,N_19308,N_19433);
nor U20625 (N_20625,N_19341,N_15493);
nand U20626 (N_20626,N_18629,N_18808);
and U20627 (N_20627,N_18948,N_18738);
and U20628 (N_20628,N_15430,N_15414);
and U20629 (N_20629,N_18064,N_18437);
nand U20630 (N_20630,N_16516,N_17921);
or U20631 (N_20631,N_19169,N_15205);
nor U20632 (N_20632,N_15963,N_17261);
and U20633 (N_20633,N_19504,N_17376);
nor U20634 (N_20634,N_18190,N_16333);
nor U20635 (N_20635,N_16405,N_17260);
nand U20636 (N_20636,N_15710,N_16928);
nor U20637 (N_20637,N_17818,N_19503);
nor U20638 (N_20638,N_16896,N_16095);
nor U20639 (N_20639,N_18550,N_17854);
or U20640 (N_20640,N_16358,N_16404);
nor U20641 (N_20641,N_17124,N_19230);
or U20642 (N_20642,N_15950,N_16634);
and U20643 (N_20643,N_18219,N_19688);
nand U20644 (N_20644,N_19193,N_15915);
or U20645 (N_20645,N_15768,N_19569);
or U20646 (N_20646,N_19386,N_17970);
nand U20647 (N_20647,N_19528,N_18961);
nor U20648 (N_20648,N_19153,N_15128);
nand U20649 (N_20649,N_19001,N_18667);
and U20650 (N_20650,N_17244,N_15152);
and U20651 (N_20651,N_18453,N_18153);
nor U20652 (N_20652,N_16237,N_16747);
and U20653 (N_20653,N_18638,N_16789);
or U20654 (N_20654,N_15371,N_18805);
nor U20655 (N_20655,N_17277,N_19545);
nand U20656 (N_20656,N_15366,N_18753);
xnor U20657 (N_20657,N_16619,N_18502);
nor U20658 (N_20658,N_19177,N_19253);
or U20659 (N_20659,N_18757,N_16573);
nor U20660 (N_20660,N_17641,N_18278);
and U20661 (N_20661,N_19980,N_15170);
nor U20662 (N_20662,N_19278,N_19863);
nand U20663 (N_20663,N_16893,N_17754);
nand U20664 (N_20664,N_19320,N_16023);
and U20665 (N_20665,N_18590,N_17392);
nor U20666 (N_20666,N_15828,N_15810);
nand U20667 (N_20667,N_19630,N_19975);
and U20668 (N_20668,N_18964,N_15380);
xnor U20669 (N_20669,N_16844,N_15614);
or U20670 (N_20670,N_16781,N_15841);
nand U20671 (N_20671,N_17408,N_18591);
nand U20672 (N_20672,N_16971,N_16444);
and U20673 (N_20673,N_19388,N_19408);
nor U20674 (N_20674,N_17910,N_16725);
or U20675 (N_20675,N_18264,N_16969);
nand U20676 (N_20676,N_16492,N_17809);
nand U20677 (N_20677,N_15013,N_15236);
and U20678 (N_20678,N_18664,N_16041);
or U20679 (N_20679,N_16490,N_19254);
and U20680 (N_20680,N_19659,N_16777);
nand U20681 (N_20681,N_15307,N_17010);
or U20682 (N_20682,N_15143,N_18089);
nand U20683 (N_20683,N_16978,N_15722);
or U20684 (N_20684,N_19735,N_16684);
nand U20685 (N_20685,N_18509,N_17428);
nand U20686 (N_20686,N_19275,N_18429);
nand U20687 (N_20687,N_17579,N_19422);
nor U20688 (N_20688,N_18122,N_16112);
nor U20689 (N_20689,N_19809,N_15411);
nor U20690 (N_20690,N_19930,N_15409);
nor U20691 (N_20691,N_19664,N_16307);
and U20692 (N_20692,N_18712,N_18907);
and U20693 (N_20693,N_17977,N_15878);
or U20694 (N_20694,N_17139,N_15863);
xor U20695 (N_20695,N_16622,N_18992);
and U20696 (N_20696,N_16061,N_19590);
nand U20697 (N_20697,N_16440,N_17795);
and U20698 (N_20698,N_18599,N_16827);
nor U20699 (N_20699,N_15178,N_17364);
xor U20700 (N_20700,N_19108,N_16616);
nand U20701 (N_20701,N_16190,N_16337);
nor U20702 (N_20702,N_15519,N_17213);
or U20703 (N_20703,N_18267,N_18647);
and U20704 (N_20704,N_17599,N_19178);
nor U20705 (N_20705,N_15117,N_15926);
nor U20706 (N_20706,N_17964,N_19357);
nor U20707 (N_20707,N_17092,N_17514);
nand U20708 (N_20708,N_15439,N_15763);
nand U20709 (N_20709,N_17196,N_19161);
and U20710 (N_20710,N_19325,N_16731);
and U20711 (N_20711,N_17852,N_17962);
nor U20712 (N_20712,N_16412,N_18380);
nor U20713 (N_20713,N_15499,N_16691);
nand U20714 (N_20714,N_15658,N_19651);
nand U20715 (N_20715,N_17022,N_15413);
or U20716 (N_20716,N_19214,N_17339);
nand U20717 (N_20717,N_15372,N_18858);
and U20718 (N_20718,N_17494,N_19500);
xnor U20719 (N_20719,N_17507,N_17140);
and U20720 (N_20720,N_19396,N_18382);
or U20721 (N_20721,N_15147,N_17569);
and U20722 (N_20722,N_17138,N_19767);
or U20723 (N_20723,N_17773,N_19420);
and U20724 (N_20724,N_19953,N_18390);
nor U20725 (N_20725,N_19620,N_19983);
nand U20726 (N_20726,N_17657,N_16505);
nor U20727 (N_20727,N_15650,N_15442);
or U20728 (N_20728,N_15913,N_18527);
and U20729 (N_20729,N_16724,N_15655);
nor U20730 (N_20730,N_18814,N_15547);
nor U20731 (N_20731,N_18832,N_19768);
or U20732 (N_20732,N_15822,N_16650);
nand U20733 (N_20733,N_17908,N_16238);
or U20734 (N_20734,N_16317,N_15427);
and U20735 (N_20735,N_15028,N_17117);
nand U20736 (N_20736,N_16008,N_18777);
nand U20737 (N_20737,N_18896,N_15067);
nand U20738 (N_20738,N_16303,N_18655);
and U20739 (N_20739,N_17618,N_17088);
nand U20740 (N_20740,N_16150,N_15288);
or U20741 (N_20741,N_19184,N_17959);
nand U20742 (N_20742,N_18792,N_15318);
nor U20743 (N_20743,N_15731,N_17699);
nor U20744 (N_20744,N_17612,N_17573);
and U20745 (N_20745,N_19799,N_19958);
nor U20746 (N_20746,N_15789,N_15577);
nand U20747 (N_20747,N_17726,N_15921);
nor U20748 (N_20748,N_16290,N_17071);
nand U20749 (N_20749,N_19307,N_18467);
or U20750 (N_20750,N_16193,N_17238);
or U20751 (N_20751,N_19645,N_15760);
and U20752 (N_20752,N_18148,N_19120);
xor U20753 (N_20753,N_19731,N_15037);
and U20754 (N_20754,N_19904,N_16020);
and U20755 (N_20755,N_19040,N_19346);
nand U20756 (N_20756,N_16098,N_16001);
nor U20757 (N_20757,N_16292,N_19046);
nor U20758 (N_20758,N_18051,N_16502);
nand U20759 (N_20759,N_18048,N_15041);
or U20760 (N_20760,N_16805,N_19728);
and U20761 (N_20761,N_19757,N_15645);
or U20762 (N_20762,N_18829,N_15339);
and U20763 (N_20763,N_16342,N_18403);
or U20764 (N_20764,N_16762,N_17519);
nand U20765 (N_20765,N_17471,N_18564);
nor U20766 (N_20766,N_18461,N_19144);
and U20767 (N_20767,N_19122,N_15455);
and U20768 (N_20768,N_19439,N_15502);
or U20769 (N_20769,N_17538,N_16662);
and U20770 (N_20770,N_18622,N_15058);
nand U20771 (N_20771,N_16217,N_15584);
nor U20772 (N_20772,N_18325,N_16199);
nand U20773 (N_20773,N_19623,N_16384);
or U20774 (N_20774,N_19968,N_19372);
and U20775 (N_20775,N_18925,N_19870);
and U20776 (N_20776,N_17508,N_19280);
nand U20777 (N_20777,N_17857,N_16663);
nor U20778 (N_20778,N_19317,N_16851);
nand U20779 (N_20779,N_16143,N_19751);
or U20780 (N_20780,N_19126,N_19477);
and U20781 (N_20781,N_17187,N_15172);
or U20782 (N_20782,N_19600,N_19977);
nand U20783 (N_20783,N_15987,N_17686);
and U20784 (N_20784,N_17766,N_15725);
and U20785 (N_20785,N_15248,N_18653);
nor U20786 (N_20786,N_15524,N_18671);
and U20787 (N_20787,N_15644,N_18588);
and U20788 (N_20788,N_16468,N_17439);
and U20789 (N_20789,N_17413,N_19345);
and U20790 (N_20790,N_19079,N_17723);
or U20791 (N_20791,N_15274,N_19418);
nor U20792 (N_20792,N_18087,N_17110);
nor U20793 (N_20793,N_15023,N_17974);
nor U20794 (N_20794,N_18136,N_17984);
nor U20795 (N_20795,N_19089,N_16594);
or U20796 (N_20796,N_15106,N_16120);
or U20797 (N_20797,N_18494,N_15491);
nand U20798 (N_20798,N_18751,N_15252);
nand U20799 (N_20799,N_19225,N_15591);
or U20800 (N_20800,N_16934,N_15477);
and U20801 (N_20801,N_19470,N_17311);
and U20802 (N_20802,N_18785,N_18714);
nor U20803 (N_20803,N_19982,N_16034);
nor U20804 (N_20804,N_17769,N_15775);
nor U20805 (N_20805,N_19355,N_15900);
nor U20806 (N_20806,N_18950,N_18565);
and U20807 (N_20807,N_16025,N_19987);
nand U20808 (N_20808,N_19239,N_18137);
nor U20809 (N_20809,N_19662,N_18931);
nand U20810 (N_20810,N_15936,N_16740);
and U20811 (N_20811,N_16912,N_16965);
nand U20812 (N_20812,N_17272,N_19034);
or U20813 (N_20813,N_16738,N_17145);
and U20814 (N_20814,N_15108,N_15948);
nor U20815 (N_20815,N_18628,N_18783);
nand U20816 (N_20816,N_18253,N_19499);
nor U20817 (N_20817,N_18179,N_19263);
nand U20818 (N_20818,N_19912,N_16353);
and U20819 (N_20819,N_18492,N_15905);
nand U20820 (N_20820,N_15762,N_15558);
xnor U20821 (N_20821,N_16562,N_19429);
or U20822 (N_20822,N_18942,N_18936);
nor U20823 (N_20823,N_18582,N_19711);
and U20824 (N_20824,N_17638,N_17475);
nand U20825 (N_20825,N_15767,N_18472);
nor U20826 (N_20826,N_16370,N_16080);
and U20827 (N_20827,N_18812,N_15196);
or U20828 (N_20828,N_17307,N_19186);
or U20829 (N_20829,N_15622,N_19229);
nand U20830 (N_20830,N_18503,N_19592);
and U20831 (N_20831,N_15275,N_18294);
nor U20832 (N_20832,N_17203,N_19210);
nor U20833 (N_20833,N_16140,N_18194);
or U20834 (N_20834,N_15638,N_16116);
or U20835 (N_20835,N_19713,N_19687);
and U20836 (N_20836,N_18167,N_15728);
nand U20837 (N_20837,N_19816,N_18102);
and U20838 (N_20838,N_18365,N_15906);
and U20839 (N_20839,N_17971,N_18627);
and U20840 (N_20840,N_18510,N_19367);
nand U20841 (N_20841,N_16878,N_19353);
and U20842 (N_20842,N_19455,N_19258);
nor U20843 (N_20843,N_17582,N_17418);
nor U20844 (N_20844,N_18223,N_15215);
nor U20845 (N_20845,N_19582,N_19701);
or U20846 (N_20846,N_19446,N_19330);
and U20847 (N_20847,N_18880,N_16820);
nor U20848 (N_20848,N_19686,N_15340);
or U20849 (N_20849,N_18877,N_19287);
or U20850 (N_20850,N_17442,N_18333);
and U20851 (N_20851,N_18995,N_18471);
or U20852 (N_20852,N_17049,N_15211);
nor U20853 (N_20853,N_16409,N_16513);
nor U20854 (N_20854,N_17985,N_18847);
and U20855 (N_20855,N_15468,N_17869);
or U20856 (N_20856,N_15662,N_15177);
and U20857 (N_20857,N_16941,N_18477);
nor U20858 (N_20858,N_16659,N_19393);
and U20859 (N_20859,N_15554,N_16497);
nor U20860 (N_20860,N_15461,N_19669);
or U20861 (N_20861,N_19580,N_16613);
or U20862 (N_20862,N_19326,N_17721);
nand U20863 (N_20863,N_19112,N_15109);
or U20864 (N_20864,N_16774,N_16350);
nor U20865 (N_20865,N_17989,N_17879);
or U20866 (N_20866,N_19168,N_17082);
nand U20867 (N_20867,N_18817,N_15967);
nand U20868 (N_20868,N_15456,N_19311);
and U20869 (N_20869,N_19509,N_19466);
or U20870 (N_20870,N_17900,N_15457);
nand U20871 (N_20871,N_19299,N_15325);
or U20872 (N_20872,N_17314,N_17293);
or U20873 (N_20873,N_15515,N_16904);
and U20874 (N_20874,N_19063,N_18762);
nand U20875 (N_20875,N_17309,N_16314);
and U20876 (N_20876,N_15700,N_19172);
nor U20877 (N_20877,N_19821,N_18500);
and U20878 (N_20878,N_17350,N_18970);
or U20879 (N_20879,N_16870,N_18112);
nor U20880 (N_20880,N_15891,N_18312);
or U20881 (N_20881,N_16099,N_15095);
or U20882 (N_20882,N_16345,N_19617);
nand U20883 (N_20883,N_16021,N_16750);
nor U20884 (N_20884,N_19365,N_18988);
and U20885 (N_20885,N_15573,N_16359);
or U20886 (N_20886,N_15652,N_19486);
nor U20887 (N_20887,N_16305,N_16803);
nand U20888 (N_20888,N_17040,N_17271);
or U20889 (N_20889,N_19794,N_15434);
nand U20890 (N_20890,N_15990,N_15705);
and U20891 (N_20891,N_16154,N_15149);
nor U20892 (N_20892,N_18952,N_17923);
nor U20893 (N_20893,N_16875,N_15454);
or U20894 (N_20894,N_17835,N_15343);
or U20895 (N_20895,N_18029,N_16608);
nand U20896 (N_20896,N_18440,N_15261);
nand U20897 (N_20897,N_18062,N_16950);
or U20898 (N_20898,N_17551,N_16964);
nand U20899 (N_20899,N_16104,N_18596);
or U20900 (N_20900,N_17914,N_18744);
and U20901 (N_20901,N_17331,N_19410);
and U20902 (N_20902,N_17451,N_17830);
or U20903 (N_20903,N_17760,N_17836);
or U20904 (N_20904,N_15264,N_15939);
nor U20905 (N_20905,N_18844,N_17009);
nand U20906 (N_20906,N_17807,N_16620);
nor U20907 (N_20907,N_18905,N_18901);
or U20908 (N_20908,N_16070,N_15044);
nor U20909 (N_20909,N_16548,N_15433);
and U20910 (N_20910,N_18824,N_19394);
nand U20911 (N_20911,N_17851,N_18684);
nor U20912 (N_20912,N_15194,N_16782);
nand U20913 (N_20913,N_19848,N_17276);
and U20914 (N_20914,N_15816,N_18607);
nand U20915 (N_20915,N_17235,N_18418);
or U20916 (N_20916,N_15820,N_19606);
nand U20917 (N_20917,N_18273,N_19502);
and U20918 (N_20918,N_19675,N_17718);
or U20919 (N_20919,N_17643,N_16183);
and U20920 (N_20920,N_16128,N_15861);
and U20921 (N_20921,N_18128,N_17926);
or U20922 (N_20922,N_17745,N_16250);
nand U20923 (N_20923,N_18169,N_15053);
and U20924 (N_20924,N_17993,N_15329);
nor U20925 (N_20925,N_19838,N_17981);
nor U20926 (N_20926,N_19753,N_15151);
nor U20927 (N_20927,N_17074,N_18630);
xor U20928 (N_20928,N_16561,N_19047);
or U20929 (N_20929,N_17297,N_18566);
and U20930 (N_20930,N_19522,N_18109);
nor U20931 (N_20931,N_17180,N_16396);
and U20932 (N_20932,N_18240,N_17848);
nor U20933 (N_20933,N_18547,N_18956);
nor U20934 (N_20934,N_18648,N_15249);
and U20935 (N_20935,N_16522,N_16700);
xor U20936 (N_20936,N_19960,N_19415);
nor U20937 (N_20937,N_15907,N_18331);
nor U20938 (N_20938,N_18593,N_17575);
nand U20939 (N_20939,N_18745,N_19758);
and U20940 (N_20940,N_18587,N_16300);
or U20941 (N_20941,N_17448,N_17457);
nand U20942 (N_20942,N_19359,N_15403);
and U20943 (N_20943,N_19866,N_15543);
nand U20944 (N_20944,N_15383,N_18445);
nor U20945 (N_20945,N_19201,N_16231);
nor U20946 (N_20946,N_18220,N_19722);
or U20947 (N_20947,N_17113,N_17207);
or U20948 (N_20948,N_19827,N_17706);
nand U20949 (N_20949,N_17932,N_16855);
and U20950 (N_20950,N_19782,N_16661);
nand U20951 (N_20951,N_17390,N_16214);
or U20952 (N_20952,N_18081,N_18742);
or U20953 (N_20953,N_17353,N_18012);
nor U20954 (N_20954,N_17059,N_15585);
or U20955 (N_20955,N_15556,N_15173);
nor U20956 (N_20956,N_15024,N_15011);
nor U20957 (N_20957,N_18895,N_17979);
nor U20958 (N_20958,N_19360,N_18059);
nand U20959 (N_20959,N_15203,N_19496);
or U20960 (N_20960,N_19633,N_17282);
or U20961 (N_20961,N_18358,N_18514);
nor U20962 (N_20962,N_17802,N_15974);
nand U20963 (N_20963,N_19403,N_15531);
or U20964 (N_20964,N_19947,N_17427);
nand U20965 (N_20965,N_19133,N_17526);
nand U20966 (N_20966,N_17945,N_15501);
or U20967 (N_20967,N_17590,N_18215);
or U20968 (N_20968,N_16482,N_16625);
or U20969 (N_20969,N_19100,N_19021);
nand U20970 (N_20970,N_19836,N_19948);
nand U20971 (N_20971,N_15322,N_19901);
or U20972 (N_20972,N_18608,N_15388);
nor U20973 (N_20973,N_16981,N_16243);
or U20974 (N_20974,N_18392,N_16922);
or U20975 (N_20975,N_15545,N_15265);
nor U20976 (N_20976,N_17445,N_19019);
nand U20977 (N_20977,N_16959,N_18330);
and U20978 (N_20978,N_18886,N_19844);
nor U20979 (N_20979,N_15761,N_18634);
or U20980 (N_20980,N_15576,N_19349);
and U20981 (N_20981,N_15485,N_18214);
nand U20982 (N_20982,N_16783,N_17828);
or U20983 (N_20983,N_15273,N_18898);
nand U20984 (N_20984,N_18432,N_16635);
nand U20985 (N_20985,N_17681,N_17114);
and U20986 (N_20986,N_17990,N_17212);
nor U20987 (N_20987,N_19657,N_16943);
nor U20988 (N_20988,N_17295,N_19574);
nand U20989 (N_20989,N_18869,N_18446);
or U20990 (N_20990,N_17649,N_16368);
nand U20991 (N_20991,N_19899,N_17527);
and U20992 (N_20992,N_18520,N_15541);
and U20993 (N_20993,N_19216,N_17716);
nor U20994 (N_20994,N_19018,N_15473);
or U20995 (N_20995,N_18617,N_17241);
nor U20996 (N_20996,N_19823,N_16674);
and U20997 (N_20997,N_15452,N_18830);
nand U20998 (N_20998,N_15093,N_19352);
or U20999 (N_20999,N_17354,N_19003);
nand U21000 (N_21000,N_18613,N_17742);
and U21001 (N_21001,N_18375,N_19049);
nor U21002 (N_21002,N_19025,N_17669);
or U21003 (N_21003,N_19698,N_17172);
or U21004 (N_21004,N_17654,N_17136);
and U21005 (N_21005,N_19013,N_17785);
and U21006 (N_21006,N_17873,N_16504);
nor U21007 (N_21007,N_17800,N_17252);
nor U21008 (N_21008,N_15668,N_19846);
nor U21009 (N_21009,N_17804,N_19156);
nand U21010 (N_21010,N_18284,N_16885);
nand U21011 (N_21011,N_19479,N_16069);
nor U21012 (N_21012,N_18430,N_15663);
or U21013 (N_21013,N_16275,N_19379);
nand U21014 (N_21014,N_18848,N_16479);
and U21015 (N_21015,N_16316,N_17122);
and U21016 (N_21016,N_18770,N_15272);
and U21017 (N_21017,N_19865,N_15527);
nor U21018 (N_21018,N_17034,N_15333);
or U21019 (N_21019,N_16678,N_17668);
and U21020 (N_21020,N_18160,N_17491);
nor U21021 (N_21021,N_17069,N_18932);
nand U21022 (N_21022,N_17360,N_16801);
or U21023 (N_21023,N_18174,N_16551);
and U21024 (N_21024,N_18882,N_18669);
and U21025 (N_21025,N_19934,N_16984);
nand U21026 (N_21026,N_15281,N_15384);
or U21027 (N_21027,N_16711,N_16658);
and U21028 (N_21028,N_16623,N_16531);
nand U21029 (N_21029,N_15657,N_17704);
nor U21030 (N_21030,N_15150,N_18972);
nor U21031 (N_21031,N_16203,N_16830);
and U21032 (N_21032,N_17381,N_17433);
nand U21033 (N_21033,N_19057,N_18930);
or U21034 (N_21034,N_16223,N_15741);
and U21035 (N_21035,N_17515,N_16917);
or U21036 (N_21036,N_15843,N_15182);
and U21037 (N_21037,N_18977,N_19129);
or U21038 (N_21038,N_17966,N_19264);
nor U21039 (N_21039,N_15312,N_16351);
or U21040 (N_21040,N_16832,N_15575);
nand U21041 (N_21041,N_17577,N_18283);
nor U21042 (N_21042,N_15395,N_17709);
and U21043 (N_21043,N_17883,N_15757);
nor U21044 (N_21044,N_15919,N_17595);
nand U21045 (N_21045,N_15184,N_17253);
nor U21046 (N_21046,N_19054,N_15539);
nand U21047 (N_21047,N_18173,N_16683);
nor U21048 (N_21048,N_16776,N_16987);
and U21049 (N_21049,N_18835,N_18002);
nor U21050 (N_21050,N_19956,N_17897);
nor U21051 (N_21051,N_15020,N_17470);
nand U21052 (N_21052,N_15365,N_17488);
nor U21053 (N_21053,N_17884,N_19130);
nand U21054 (N_21054,N_19220,N_18229);
nand U21055 (N_21055,N_16785,N_19578);
nor U21056 (N_21056,N_16672,N_19658);
or U21057 (N_21057,N_16863,N_15350);
nor U21058 (N_21058,N_18296,N_15233);
and U21059 (N_21059,N_17796,N_16296);
nand U21060 (N_21060,N_15805,N_18626);
nand U21061 (N_21061,N_16794,N_18182);
nand U21062 (N_21062,N_17838,N_16423);
nand U21063 (N_21063,N_16643,N_16585);
nor U21064 (N_21064,N_16084,N_16100);
and U21065 (N_21065,N_16179,N_18201);
nand U21066 (N_21066,N_19584,N_17872);
and U21067 (N_21067,N_15262,N_16615);
xor U21068 (N_21068,N_15631,N_18397);
nor U21069 (N_21069,N_18518,N_15535);
nor U21070 (N_21070,N_19286,N_19999);
or U21071 (N_21071,N_17424,N_18754);
and U21072 (N_21072,N_15399,N_15207);
nand U21073 (N_21073,N_17368,N_17673);
or U21074 (N_21074,N_19111,N_15885);
or U21075 (N_21075,N_17667,N_17694);
or U21076 (N_21076,N_19124,N_15683);
nor U21077 (N_21077,N_17289,N_19375);
and U21078 (N_21078,N_16991,N_18944);
and U21079 (N_21079,N_19546,N_17058);
nor U21080 (N_21080,N_15785,N_17903);
and U21081 (N_21081,N_15595,N_19540);
and U21082 (N_21082,N_18837,N_18947);
nor U21083 (N_21083,N_15126,N_17867);
nand U21084 (N_21084,N_16421,N_16329);
and U21085 (N_21085,N_19038,N_17753);
nor U21086 (N_21086,N_16461,N_18719);
nor U21087 (N_21087,N_17387,N_15316);
nor U21088 (N_21088,N_19114,N_18001);
and U21089 (N_21089,N_18188,N_15003);
nand U21090 (N_21090,N_19337,N_17823);
or U21091 (N_21091,N_19454,N_16071);
nor U21092 (N_21092,N_16698,N_19084);
and U21093 (N_21093,N_19008,N_16426);
nand U21094 (N_21094,N_18557,N_16748);
or U21095 (N_21095,N_16074,N_16378);
nand U21096 (N_21096,N_18991,N_15578);
nor U21097 (N_21097,N_16813,N_17890);
and U21098 (N_21098,N_16918,N_19811);
and U21099 (N_21099,N_19321,N_15916);
or U21100 (N_21100,N_15618,N_17317);
and U21101 (N_21101,N_19348,N_16695);
and U21102 (N_21102,N_17814,N_18885);
and U21103 (N_21103,N_19514,N_19734);
nand U21104 (N_21104,N_16555,N_18960);
or U21105 (N_21105,N_17053,N_19343);
nand U21106 (N_21106,N_15014,N_19481);
and U21107 (N_21107,N_15508,N_19967);
nor U21108 (N_21108,N_17358,N_19272);
and U21109 (N_21109,N_19190,N_15155);
nor U21110 (N_21110,N_15336,N_16240);
and U21111 (N_21111,N_15302,N_18981);
nor U21112 (N_21112,N_16270,N_16289);
and U21113 (N_21113,N_16176,N_15276);
and U21114 (N_21114,N_18227,N_15352);
and U21115 (N_21115,N_17651,N_16189);
nor U21116 (N_21116,N_17248,N_19916);
nand U21117 (N_21117,N_19989,N_15793);
nand U21118 (N_21118,N_17813,N_19073);
nand U21119 (N_21119,N_17490,N_18041);
and U21120 (N_21120,N_16373,N_17670);
nand U21121 (N_21121,N_18363,N_16812);
nor U21122 (N_21122,N_18286,N_18295);
or U21123 (N_21123,N_18378,N_19525);
or U21124 (N_21124,N_16752,N_15946);
xnor U21125 (N_21125,N_19921,N_19797);
nand U21126 (N_21126,N_19173,N_18790);
and U21127 (N_21127,N_18891,N_18853);
nor U21128 (N_21128,N_18005,N_15996);
nand U21129 (N_21129,N_18262,N_19327);
nand U21130 (N_21130,N_19654,N_16519);
or U21131 (N_21131,N_18114,N_15054);
nand U21132 (N_21132,N_18037,N_17478);
or U21133 (N_21133,N_19248,N_17473);
or U21134 (N_21134,N_19986,N_16848);
or U21135 (N_21135,N_18178,N_16213);
and U21136 (N_21136,N_18700,N_19744);
or U21137 (N_21137,N_18498,N_19508);
or U21138 (N_21138,N_17378,N_17895);
or U21139 (N_21139,N_17799,N_17767);
nor U21140 (N_21140,N_19996,N_19276);
nand U21141 (N_21141,N_17539,N_19488);
and U21142 (N_21142,N_15216,N_15532);
nor U21143 (N_21143,N_15102,N_15890);
or U21144 (N_21144,N_16073,N_17406);
or U21145 (N_21145,N_18308,N_19610);
nand U21146 (N_21146,N_19165,N_15389);
nor U21147 (N_21147,N_15046,N_19456);
nand U21148 (N_21148,N_19862,N_15603);
or U21149 (N_21149,N_18616,N_17999);
nand U21150 (N_21150,N_17189,N_19742);
xor U21151 (N_21151,N_16352,N_18973);
nand U21152 (N_21152,N_18938,N_17287);
and U21153 (N_21153,N_17777,N_15882);
nor U21154 (N_21154,N_15096,N_16867);
nor U21155 (N_21155,N_18774,N_18939);
and U21156 (N_21156,N_19705,N_19720);
or U21157 (N_21157,N_15931,N_18084);
nand U21158 (N_21158,N_17308,N_15602);
and U21159 (N_21159,N_16660,N_18612);
nand U21160 (N_21160,N_19460,N_18643);
or U21161 (N_21161,N_15688,N_18765);
and U21162 (N_21162,N_15520,N_16518);
and U21163 (N_21163,N_18483,N_17288);
and U21164 (N_21164,N_19529,N_19166);
nor U21165 (N_21165,N_18641,N_17679);
nand U21166 (N_21166,N_19145,N_17425);
and U21167 (N_21167,N_16670,N_17469);
nor U21168 (N_21168,N_17936,N_16266);
xnor U21169 (N_21169,N_15553,N_18803);
nand U21170 (N_21170,N_17056,N_16295);
nor U21171 (N_21171,N_16995,N_19085);
and U21172 (N_21172,N_15529,N_17410);
nor U21173 (N_21173,N_18834,N_19691);
nor U21174 (N_21174,N_16192,N_17858);
nor U21175 (N_21175,N_19473,N_18236);
nor U21176 (N_21176,N_17477,N_19512);
nand U21177 (N_21177,N_17675,N_15696);
or U21178 (N_21178,N_15690,N_15417);
or U21179 (N_21179,N_17541,N_16297);
or U21180 (N_21180,N_17574,N_15715);
xor U21181 (N_21181,N_15391,N_16901);
or U21182 (N_21182,N_17933,N_16532);
and U21183 (N_21183,N_15922,N_17437);
xnor U21184 (N_21184,N_18595,N_16294);
and U21185 (N_21185,N_18718,N_15101);
nand U21186 (N_21186,N_19962,N_18057);
or U21187 (N_21187,N_17313,N_18291);
or U21188 (N_21188,N_17256,N_16726);
nand U21189 (N_21189,N_16398,N_15954);
or U21190 (N_21190,N_18470,N_17026);
nand U21191 (N_21191,N_19792,N_15640);
and U21192 (N_21192,N_19624,N_19938);
or U21193 (N_21193,N_16933,N_15779);
and U21194 (N_21194,N_18890,N_17407);
and U21195 (N_21195,N_16302,N_19703);
nand U21196 (N_21196,N_19082,N_18311);
nor U21197 (N_21197,N_15206,N_17965);
and U21198 (N_21198,N_17204,N_18656);
nor U21199 (N_21199,N_19876,N_15423);
nor U21200 (N_21200,N_16253,N_18479);
and U21201 (N_21201,N_18402,N_18776);
nor U21202 (N_21202,N_18293,N_18749);
nor U21203 (N_21203,N_18346,N_18941);
or U21204 (N_21204,N_18455,N_17817);
nand U21205 (N_21205,N_16826,N_19549);
nor U21206 (N_21206,N_15800,N_19453);
or U21207 (N_21207,N_15894,N_17916);
nor U21208 (N_21208,N_17243,N_16769);
and U21209 (N_21209,N_17419,N_17534);
nand U21210 (N_21210,N_16982,N_18841);
and U21211 (N_21211,N_18989,N_18416);
nand U21212 (N_21212,N_18465,N_18507);
and U21213 (N_21213,N_18175,N_17169);
and U21214 (N_21214,N_15083,N_17440);
and U21215 (N_21215,N_19260,N_17880);
or U21216 (N_21216,N_19472,N_15202);
and U21217 (N_21217,N_18292,N_15123);
and U21218 (N_21218,N_19694,N_15605);
and U21219 (N_21219,N_15979,N_19119);
nor U21220 (N_21220,N_18400,N_15354);
or U21221 (N_21221,N_18772,N_19629);
nor U21222 (N_21222,N_18187,N_17265);
or U21223 (N_21223,N_19497,N_16118);
and U21224 (N_21224,N_18747,N_17011);
nor U21225 (N_21225,N_19319,N_19826);
nand U21226 (N_21226,N_19966,N_17697);
and U21227 (N_21227,N_15253,N_16360);
and U21228 (N_21228,N_17738,N_18592);
and U21229 (N_21229,N_16642,N_17708);
nor U21230 (N_21230,N_17860,N_16145);
and U21231 (N_21231,N_16315,N_16134);
nor U21232 (N_21232,N_16727,N_16149);
nand U21233 (N_21233,N_16633,N_18066);
nand U21234 (N_21234,N_16681,N_15959);
or U21235 (N_21235,N_16196,N_15823);
nor U21236 (N_21236,N_15707,N_19715);
nor U21237 (N_21237,N_18673,N_17072);
or U21238 (N_21238,N_17174,N_18600);
or U21239 (N_21239,N_15685,N_18958);
nor U21240 (N_21240,N_16344,N_16923);
or U21241 (N_21241,N_16277,N_18108);
or U21242 (N_21242,N_16210,N_18559);
xnor U21243 (N_21243,N_19712,N_15673);
nand U21244 (N_21244,N_16371,N_17098);
and U21245 (N_21245,N_16957,N_16212);
nor U21246 (N_21246,N_17610,N_16751);
or U21247 (N_21247,N_16651,N_19074);
nand U21248 (N_21248,N_16366,N_15865);
or U21249 (N_21249,N_17161,N_16511);
or U21250 (N_21250,N_17928,N_16466);
nor U21251 (N_21251,N_18546,N_19685);
or U21252 (N_21252,N_15503,N_17759);
nand U21253 (N_21253,N_17660,N_16427);
nor U21254 (N_21254,N_16865,N_18024);
nand U21255 (N_21255,N_16038,N_18261);
nor U21256 (N_21256,N_15017,N_16654);
nor U21257 (N_21257,N_15321,N_15798);
and U21258 (N_21258,N_15588,N_18379);
nand U21259 (N_21259,N_18982,N_16052);
xnor U21260 (N_21260,N_16692,N_19045);
nand U21261 (N_21261,N_18452,N_17611);
nand U21262 (N_21262,N_18456,N_17815);
or U21263 (N_21263,N_15621,N_17918);
or U21264 (N_21264,N_18589,N_16132);
and U21265 (N_21265,N_15034,N_15471);
and U21266 (N_21266,N_16157,N_15880);
nand U21267 (N_21267,N_19458,N_16545);
nand U21268 (N_21268,N_16262,N_17052);
or U21269 (N_21269,N_18897,N_18356);
xor U21270 (N_21270,N_15975,N_15381);
nor U21271 (N_21271,N_15770,N_19961);
nand U21272 (N_21272,N_19515,N_16365);
nand U21273 (N_21273,N_16208,N_18504);
nor U21274 (N_21274,N_15988,N_16169);
nand U21275 (N_21275,N_17038,N_17153);
nor U21276 (N_21276,N_18315,N_18213);
nand U21277 (N_21277,N_18966,N_15628);
nor U21278 (N_21278,N_19137,N_17905);
and U21279 (N_21279,N_17046,N_18313);
or U21280 (N_21280,N_16246,N_17597);
or U21281 (N_21281,N_17737,N_19707);
nor U21282 (N_21282,N_19412,N_17303);
nand U21283 (N_21283,N_18574,N_17516);
nand U21284 (N_21284,N_16560,N_19759);
nand U21285 (N_21285,N_19259,N_15758);
nand U21286 (N_21286,N_18499,N_19749);
and U21287 (N_21287,N_17891,N_16077);
and U21288 (N_21288,N_15993,N_16338);
nor U21289 (N_21289,N_15849,N_16544);
and U21290 (N_21290,N_16162,N_18411);
nor U21291 (N_21291,N_16535,N_17060);
nor U21292 (N_21292,N_16773,N_18996);
or U21293 (N_21293,N_16576,N_17379);
or U21294 (N_21294,N_19012,N_15319);
or U21295 (N_21295,N_18027,N_18721);
nand U21296 (N_21296,N_18118,N_16335);
nor U21297 (N_21297,N_18784,N_17550);
and U21298 (N_21298,N_19552,N_16096);
and U21299 (N_21299,N_15809,N_17077);
and U21300 (N_21300,N_15716,N_19894);
nand U21301 (N_21301,N_19677,N_19005);
nand U21302 (N_21302,N_15500,N_18422);
nor U21303 (N_21303,N_17614,N_15776);
nor U21304 (N_21304,N_19738,N_19805);
or U21305 (N_21305,N_18451,N_15065);
nand U21306 (N_21306,N_17434,N_16636);
nand U21307 (N_21307,N_19140,N_16011);
nor U21308 (N_21308,N_17537,N_15405);
nor U21309 (N_21309,N_18893,N_17771);
and U21310 (N_21310,N_18928,N_17100);
and U21311 (N_21311,N_15133,N_19231);
and U21312 (N_21312,N_17091,N_15720);
nand U21313 (N_21313,N_19274,N_16311);
and U21314 (N_21314,N_19060,N_16113);
or U21315 (N_21315,N_17367,N_19562);
nor U21316 (N_21316,N_18598,N_19990);
and U21317 (N_21317,N_19853,N_16760);
and U21318 (N_21318,N_19868,N_18971);
nand U21319 (N_21319,N_17609,N_17294);
nor U21320 (N_21320,N_19883,N_19756);
or U21321 (N_21321,N_18650,N_16927);
or U21322 (N_21322,N_15165,N_19593);
nand U21323 (N_21323,N_19237,N_19224);
nand U21324 (N_21324,N_18314,N_18263);
nand U21325 (N_21325,N_18268,N_17019);
nand U21326 (N_21326,N_16986,N_17975);
and U21327 (N_21327,N_18200,N_18584);
nor U21328 (N_21328,N_15190,N_17950);
and U21329 (N_21329,N_19663,N_17027);
nand U21330 (N_21330,N_17585,N_16452);
nand U21331 (N_21331,N_19941,N_16899);
and U21332 (N_21332,N_17200,N_17458);
nor U21333 (N_21333,N_15807,N_17731);
or U21334 (N_21334,N_18706,N_17841);
xnor U21335 (N_21335,N_15238,N_16872);
nor U21336 (N_21336,N_16142,N_18110);
or U21337 (N_21337,N_18147,N_19087);
nand U21338 (N_21338,N_19577,N_19340);
or U21339 (N_21339,N_17513,N_19890);
or U21340 (N_21340,N_18285,N_18327);
nand U21341 (N_21341,N_18257,N_15870);
and U21342 (N_21342,N_17957,N_18345);
nor U21343 (N_21343,N_18998,N_15856);
nand U21344 (N_21344,N_18879,N_15536);
nor U21345 (N_21345,N_19978,N_18921);
nand U21346 (N_21346,N_19358,N_19653);
nor U21347 (N_21347,N_17359,N_19304);
and U21348 (N_21348,N_18810,N_16251);
nor U21349 (N_21349,N_16151,N_15038);
nor U21350 (N_21350,N_16341,N_15726);
nor U21351 (N_21351,N_16131,N_17954);
nand U21352 (N_21352,N_18833,N_17917);
nor U21353 (N_21353,N_16823,N_18768);
or U21354 (N_21354,N_18045,N_15099);
nand U21355 (N_21355,N_18368,N_17581);
nand U21356 (N_21356,N_17270,N_17625);
and U21357 (N_21357,N_17523,N_19151);
nor U21358 (N_21358,N_17727,N_17929);
nor U21359 (N_21359,N_16063,N_15844);
and U21360 (N_21360,N_15968,N_18210);
nor U21361 (N_21361,N_16547,N_17889);
or U21362 (N_21362,N_15416,N_18105);
nand U21363 (N_21363,N_17008,N_17728);
or U21364 (N_21364,N_17748,N_17467);
nand U21365 (N_21365,N_16873,N_18806);
nand U21366 (N_21366,N_17342,N_15089);
and U21367 (N_21367,N_16022,N_15969);
or U21368 (N_21368,N_16829,N_16419);
or U21369 (N_21369,N_17770,N_15879);
nand U21370 (N_21370,N_19959,N_15814);
and U21371 (N_21371,N_18851,N_16381);
nand U21372 (N_21372,N_19262,N_16859);
nor U21373 (N_21373,N_18329,N_19671);
nand U21374 (N_21374,N_15055,N_17249);
nand U21375 (N_21375,N_17182,N_19974);
nor U21376 (N_21376,N_15736,N_17567);
nand U21377 (N_21377,N_15154,N_17543);
nor U21378 (N_21378,N_19207,N_15406);
nor U21379 (N_21379,N_18674,N_17938);
nor U21380 (N_21380,N_17904,N_15432);
and U21381 (N_21381,N_16013,N_16759);
or U21382 (N_21382,N_18475,N_19743);
nand U21383 (N_21383,N_19850,N_18603);
and U21384 (N_21384,N_19541,N_16083);
nand U21385 (N_21385,N_16029,N_16556);
or U21386 (N_21386,N_18695,N_15898);
xor U21387 (N_21387,N_16407,N_19523);
nor U21388 (N_21388,N_16463,N_19807);
nor U21389 (N_21389,N_16076,N_18639);
or U21390 (N_21390,N_15888,N_16428);
or U21391 (N_21391,N_16990,N_15310);
or U21392 (N_21392,N_17931,N_19845);
and U21393 (N_21393,N_18009,N_15599);
and U21394 (N_21394,N_16055,N_17429);
and U21395 (N_21395,N_19413,N_16232);
nand U21396 (N_21396,N_15467,N_17017);
xor U21397 (N_21397,N_19291,N_15699);
nand U21398 (N_21398,N_17214,N_17849);
or U21399 (N_21399,N_15732,N_19747);
and U21400 (N_21400,N_17661,N_16137);
and U21401 (N_21401,N_16465,N_16920);
or U21402 (N_21402,N_15127,N_17847);
nand U21403 (N_21403,N_16766,N_15626);
nand U21404 (N_21404,N_17666,N_15897);
and U21405 (N_21405,N_17076,N_18324);
and U21406 (N_21406,N_15495,N_18533);
nand U21407 (N_21407,N_18581,N_15572);
or U21408 (N_21408,N_16897,N_17626);
and U21409 (N_21409,N_19513,N_18530);
and U21410 (N_21410,N_15918,N_15601);
nor U21411 (N_21411,N_19775,N_19421);
and U21412 (N_21412,N_16540,N_15884);
or U21413 (N_21413,N_16612,N_16952);
nor U21414 (N_21414,N_15571,N_16565);
nand U21415 (N_21415,N_15835,N_16439);
nor U21416 (N_21416,N_17202,N_18355);
or U21417 (N_21417,N_16259,N_19556);
or U21418 (N_21418,N_18318,N_17665);
and U21419 (N_21419,N_15201,N_17064);
or U21420 (N_21420,N_17535,N_15021);
nor U21421 (N_21421,N_17943,N_17504);
nor U21422 (N_21422,N_17919,N_16056);
and U21423 (N_21423,N_18870,N_17394);
xnor U21424 (N_21424,N_17029,N_17028);
nand U21425 (N_21425,N_17949,N_18023);
and U21426 (N_21426,N_15782,N_19245);
or U21427 (N_21427,N_15324,N_19314);
xnor U21428 (N_21428,N_16166,N_15078);
nor U21429 (N_21429,N_18614,N_16534);
and U21430 (N_21430,N_18156,N_17556);
and U21431 (N_21431,N_15328,N_19672);
and U21432 (N_21432,N_19748,N_19461);
nand U21433 (N_21433,N_17233,N_19457);
nor U21434 (N_21434,N_15787,N_19313);
xor U21435 (N_21435,N_16935,N_19235);
and U21436 (N_21436,N_19762,N_16309);
and U21437 (N_21437,N_16082,N_16702);
or U21438 (N_21438,N_16094,N_18342);
nand U21439 (N_21439,N_16857,N_16081);
and U21440 (N_21440,N_15247,N_19702);
or U21441 (N_21441,N_16107,N_15344);
nor U21442 (N_21442,N_15680,N_15498);
nand U21443 (N_21443,N_17154,N_18821);
nand U21444 (N_21444,N_15122,N_18473);
and U21445 (N_21445,N_18828,N_19218);
nand U21446 (N_21446,N_16821,N_18692);
nand U21447 (N_21447,N_18042,N_15952);
nor U21448 (N_21448,N_16819,N_19627);
nor U21449 (N_21449,N_19806,N_17653);
and U21450 (N_21450,N_15872,N_17152);
or U21451 (N_21451,N_15613,N_16656);
and U21452 (N_21452,N_19055,N_19790);
nor U21453 (N_21453,N_18801,N_19335);
or U21454 (N_21454,N_19716,N_18095);
nand U21455 (N_21455,N_19566,N_17887);
nand U21456 (N_21456,N_15886,N_16293);
and U21457 (N_21457,N_16999,N_17560);
nand U21458 (N_21458,N_16006,N_19076);
and U21459 (N_21459,N_16646,N_17266);
nand U21460 (N_21460,N_19127,N_15482);
nand U21461 (N_21461,N_18859,N_16730);
and U21462 (N_21462,N_19785,N_17642);
nor U21463 (N_21463,N_19563,N_19438);
nor U21464 (N_21464,N_16417,N_17351);
nand U21465 (N_21465,N_18515,N_19614);
nand U21466 (N_21466,N_15517,N_15876);
xnor U21467 (N_21467,N_19257,N_18748);
or U21468 (N_21468,N_16574,N_15971);
xnor U21469 (N_21469,N_15279,N_16114);
nor U21470 (N_21470,N_17365,N_19940);
and U21471 (N_21471,N_19914,N_16144);
and U21472 (N_21472,N_18496,N_15360);
or U21473 (N_21473,N_16032,N_17810);
or U21474 (N_21474,N_18929,N_15773);
and U21475 (N_21475,N_18563,N_16807);
or U21476 (N_21476,N_17645,N_19102);
or U21477 (N_21477,N_19128,N_17484);
or U21478 (N_21478,N_15873,N_18789);
and U21479 (N_21479,N_19872,N_17808);
nand U21480 (N_21480,N_15394,N_18387);
nor U21481 (N_21481,N_18073,N_15250);
xor U21482 (N_21482,N_18506,N_16172);
and U21483 (N_21483,N_16247,N_17955);
and U21484 (N_21484,N_17184,N_17875);
nor U21485 (N_21485,N_17794,N_18458);
nand U21486 (N_21486,N_15169,N_18854);
nand U21487 (N_21487,N_15460,N_15351);
nor U21488 (N_21488,N_19655,N_15651);
nand U21489 (N_21489,N_19103,N_18984);
and U21490 (N_21490,N_19900,N_17412);
and U21491 (N_21491,N_18026,N_18233);
nand U21492 (N_21492,N_16599,N_18800);
nand U21493 (N_21493,N_15646,N_15214);
xnor U21494 (N_21494,N_19174,N_16435);
xnor U21495 (N_21495,N_19777,N_16900);
xor U21496 (N_21496,N_15994,N_17664);
xnor U21497 (N_21497,N_15808,N_17018);
and U21498 (N_21498,N_19271,N_15867);
xor U21499 (N_21499,N_16376,N_19955);
or U21500 (N_21500,N_18922,N_18549);
nor U21501 (N_21501,N_16549,N_18980);
and U21502 (N_21502,N_19547,N_19395);
nand U21503 (N_21503,N_16967,N_16230);
nor U21504 (N_21504,N_15812,N_17719);
and U21505 (N_21505,N_16301,N_17829);
nor U21506 (N_21506,N_15654,N_19331);
and U21507 (N_21507,N_18716,N_19246);
xor U21508 (N_21508,N_18849,N_17325);
and U21509 (N_21509,N_15692,N_16962);
nor U21510 (N_21510,N_17646,N_15337);
and U21511 (N_21511,N_19929,N_17747);
nand U21512 (N_21512,N_18601,N_18548);
or U21513 (N_21513,N_18191,N_19289);
and U21514 (N_21514,N_15346,N_19222);
nor U21515 (N_21515,N_18969,N_18799);
and U21516 (N_21516,N_19007,N_16066);
and U21517 (N_21517,N_15419,N_16049);
nor U21518 (N_21518,N_15818,N_16354);
or U21519 (N_21519,N_19143,N_15665);
nand U21520 (N_21520,N_16597,N_15766);
or U21521 (N_21521,N_15268,N_17383);
nand U21522 (N_21522,N_16355,N_15721);
and U21523 (N_21523,N_17335,N_19935);
nand U21524 (N_21524,N_16778,N_16945);
or U21525 (N_21525,N_16012,N_16564);
nand U21526 (N_21526,N_19644,N_16382);
and U21527 (N_21527,N_15080,N_19613);
or U21528 (N_21528,N_17843,N_17305);
nand U21529 (N_21529,N_15464,N_19741);
nor U21530 (N_21530,N_19954,N_17986);
and U21531 (N_21531,N_18038,N_19766);
nand U21532 (N_21532,N_17423,N_18739);
or U21533 (N_21533,N_17571,N_17958);
nand U21534 (N_21534,N_18909,N_17631);
nor U21535 (N_21535,N_15634,N_16248);
nor U21536 (N_21536,N_19232,N_16735);
nand U21537 (N_21537,N_16533,N_18825);
or U21538 (N_21538,N_18069,N_19385);
or U21539 (N_21539,N_17988,N_17403);
nor U21540 (N_21540,N_15451,N_16186);
or U21541 (N_21541,N_19595,N_16604);
or U21542 (N_21542,N_15661,N_16148);
nor U21543 (N_21543,N_17333,N_18195);
nand U21544 (N_21544,N_19559,N_17632);
nor U21545 (N_21545,N_15609,N_17946);
nor U21546 (N_21546,N_17258,N_15002);
nor U21547 (N_21547,N_16804,N_18680);
and U21548 (N_21548,N_19988,N_15676);
and U21549 (N_21549,N_15114,N_19067);
nand U21550 (N_21550,N_16841,N_16483);
and U21551 (N_21551,N_18360,N_18056);
or U21552 (N_21552,N_19824,N_17158);
nor U21553 (N_21553,N_17449,N_15299);
nand U21554 (N_21554,N_17322,N_16086);
nand U21555 (N_21555,N_17047,N_16291);
or U21556 (N_21556,N_17231,N_17001);
and U21557 (N_21557,N_17037,N_17604);
nand U21558 (N_21558,N_18920,N_18511);
nand U21559 (N_21559,N_19036,N_15400);
nand U21560 (N_21560,N_18270,N_17454);
nor U21561 (N_21561,N_16024,N_17788);
or U21562 (N_21562,N_15315,N_17580);
and U21563 (N_21563,N_18523,N_17911);
nand U21564 (N_21564,N_18766,N_17393);
or U21565 (N_21565,N_18594,N_15084);
nand U21566 (N_21566,N_19915,N_17306);
or U21567 (N_21567,N_19043,N_16225);
nand U21568 (N_21568,N_16447,N_17106);
nor U21569 (N_21569,N_19945,N_15269);
nand U21570 (N_21570,N_17328,N_16207);
nor U21571 (N_21571,N_16200,N_18271);
nand U21572 (N_21572,N_16877,N_18532);
or U21573 (N_21573,N_17587,N_17396);
xor U21574 (N_21574,N_18260,N_15045);
nor U21575 (N_21575,N_18654,N_18543);
nor U21576 (N_21576,N_16506,N_16168);
nor U21577 (N_21577,N_19217,N_16085);
or U21578 (N_21578,N_19363,N_16489);
and U21579 (N_21579,N_15567,N_15141);
nand U21580 (N_21580,N_18036,N_15607);
nor U21581 (N_21581,N_16713,N_17283);
xnor U21582 (N_21582,N_18644,N_18976);
nor U21583 (N_21583,N_19160,N_17137);
and U21584 (N_21584,N_17790,N_15217);
and U21585 (N_21585,N_18724,N_16770);
nor U21586 (N_21586,N_18836,N_19791);
nand U21587 (N_21587,N_16187,N_17621);
nor U21588 (N_21588,N_15929,N_18245);
nand U21589 (N_21589,N_17920,N_17320);
nand U21590 (N_21590,N_17827,N_17850);
nor U21591 (N_21591,N_15625,N_15342);
or U21592 (N_21592,N_18082,N_16216);
and U21593 (N_21593,N_15047,N_19984);
nor U21594 (N_21594,N_18357,N_17822);
nand U21595 (N_21595,N_19462,N_17337);
and U21596 (N_21596,N_16884,N_18338);
nor U21597 (N_21597,N_16387,N_17789);
and U21598 (N_21598,N_17691,N_16400);
nand U21599 (N_21599,N_15983,N_17162);
and U21600 (N_21600,N_17522,N_16693);
nand U21601 (N_21601,N_17460,N_18063);
nand U21602 (N_21602,N_15356,N_19090);
nand U21603 (N_21603,N_19798,N_16854);
xor U21604 (N_21604,N_16537,N_16741);
and U21605 (N_21605,N_17066,N_15379);
or U21606 (N_21606,N_19976,N_18277);
nor U21607 (N_21607,N_19875,N_15755);
and U21608 (N_21608,N_17363,N_15542);
and U21609 (N_21609,N_19095,N_19377);
or U21610 (N_21610,N_18025,N_17375);
or U21611 (N_21611,N_17892,N_15404);
nand U21612 (N_21612,N_18426,N_15119);
or U21613 (N_21613,N_18301,N_17286);
and U21614 (N_21614,N_17493,N_15087);
nor U21615 (N_21615,N_17792,N_18343);
nand U21616 (N_21616,N_19871,N_15069);
nor U21617 (N_21617,N_15357,N_16779);
and U21618 (N_21618,N_15098,N_18370);
and U21619 (N_21619,N_19810,N_19510);
nor U21620 (N_21620,N_16499,N_19972);
nor U21621 (N_21621,N_15765,N_16790);
nand U21622 (N_21622,N_18079,N_18361);
and U21623 (N_21623,N_17925,N_16602);
or U21624 (N_21624,N_18672,N_17055);
nand U21625 (N_21625,N_15064,N_15443);
and U21626 (N_21626,N_16349,N_17909);
nor U21627 (N_21627,N_15107,N_17366);
nand U21628 (N_21628,N_19781,N_17399);
or U21629 (N_21629,N_17215,N_15937);
or U21630 (N_21630,N_15935,N_16429);
or U21631 (N_21631,N_17246,N_19480);
and U21632 (N_21632,N_16924,N_17762);
nor U21633 (N_21633,N_16734,N_19887);
or U21634 (N_21634,N_19903,N_15378);
and U21635 (N_21635,N_19195,N_17150);
or U21636 (N_21636,N_15637,N_16339);
nand U21637 (N_21637,N_17045,N_16914);
or U21638 (N_21638,N_16954,N_16603);
and U21639 (N_21639,N_16306,N_18065);
nand U21640 (N_21640,N_16416,N_17178);
and U21641 (N_21641,N_16953,N_16687);
nand U21642 (N_21642,N_16401,N_19056);
and U21643 (N_21643,N_18359,N_19815);
and U21644 (N_21644,N_17713,N_16580);
or U21645 (N_21645,N_19373,N_19118);
nand U21646 (N_21646,N_17695,N_19449);
nand U21647 (N_21647,N_19407,N_18908);
nand U21648 (N_21648,N_15210,N_17707);
xor U21649 (N_21649,N_16274,N_18852);
nand U21650 (N_21650,N_15426,N_16723);
nor U21651 (N_21651,N_18119,N_16092);
or U21652 (N_21652,N_15643,N_17316);
nand U21653 (N_21653,N_15458,N_17589);
or U21654 (N_21654,N_17758,N_19452);
xnor U21655 (N_21655,N_18151,N_19832);
nand U21656 (N_21656,N_16771,N_16811);
or U21657 (N_21657,N_15920,N_17776);
nand U21658 (N_21658,N_16980,N_18750);
and U21659 (N_21659,N_19431,N_17987);
or U21660 (N_21660,N_15689,N_19117);
nand U21661 (N_21661,N_18433,N_17479);
nor U21662 (N_21662,N_19856,N_17793);
nor U21663 (N_21663,N_16194,N_16402);
nor U21664 (N_21664,N_19284,N_19212);
nor U21665 (N_21665,N_16443,N_16481);
or U21666 (N_21666,N_16059,N_15134);
nand U21667 (N_21667,N_18198,N_19115);
or U21668 (N_21668,N_18615,N_15636);
xnor U21669 (N_21669,N_16002,N_16708);
nor U21670 (N_21670,N_16326,N_17044);
nor U21671 (N_21671,N_19918,N_19101);
nand U21672 (N_21672,N_18369,N_17520);
and U21673 (N_21673,N_17012,N_17107);
nor U21674 (N_21674,N_16628,N_15032);
nand U21675 (N_21675,N_17039,N_19939);
or U21676 (N_21676,N_18003,N_15899);
or U21677 (N_21677,N_19879,N_15803);
or U21678 (N_21678,N_18352,N_17377);
xor U21679 (N_21679,N_17352,N_18171);
nor U21680 (N_21680,N_17640,N_16089);
nand U21681 (N_21681,N_19544,N_16093);
nor U21682 (N_21682,N_16753,N_19238);
or U21683 (N_21683,N_17983,N_18258);
nand U21684 (N_21684,N_16097,N_18545);
or U21685 (N_21685,N_17826,N_18687);
and U21686 (N_21686,N_17995,N_15738);
nand U21687 (N_21687,N_19997,N_19800);
xnor U21688 (N_21688,N_19445,N_18335);
nor U21689 (N_21689,N_15903,N_19069);
nor U21690 (N_21690,N_19946,N_16822);
nand U21691 (N_21691,N_19998,N_18424);
and U21692 (N_21692,N_19435,N_15684);
and U21693 (N_21693,N_16913,N_16265);
nor U21694 (N_21694,N_18097,N_19598);
nor U21695 (N_21695,N_15635,N_15157);
nand U21696 (N_21696,N_16016,N_16664);
or U21697 (N_21697,N_17674,N_16005);
and U21698 (N_21698,N_16742,N_16621);
or U21699 (N_21699,N_18060,N_17505);
nand U21700 (N_21700,N_17973,N_15938);
or U21701 (N_21701,N_16003,N_15359);
nor U21702 (N_21702,N_19555,N_18040);
nor U21703 (N_21703,N_16979,N_16587);
and U21704 (N_21704,N_16925,N_17073);
or U21705 (N_21705,N_17131,N_16946);
or U21706 (N_21706,N_18337,N_18737);
xnor U21707 (N_21707,N_18385,N_16422);
nor U21708 (N_21708,N_17236,N_17592);
nand U21709 (N_21709,N_17324,N_17280);
or U21710 (N_21710,N_15291,N_17304);
nor U21711 (N_21711,N_16233,N_16966);
and U21712 (N_21712,N_19771,N_19913);
nor U21713 (N_21713,N_18866,N_17224);
or U21714 (N_21714,N_19157,N_18482);
nand U21715 (N_21715,N_19249,N_18022);
or U21716 (N_21716,N_17481,N_16524);
nand U21717 (N_21717,N_17740,N_17147);
nor U21718 (N_21718,N_16141,N_16241);
nand U21719 (N_21719,N_17820,N_15845);
and U21720 (N_21720,N_18255,N_18469);
or U21721 (N_21721,N_15232,N_17562);
nand U21722 (N_21722,N_19818,N_19383);
nor U21723 (N_21723,N_18558,N_15797);
or U21724 (N_21724,N_17078,N_19874);
or U21725 (N_21725,N_15749,N_17075);
nor U21726 (N_21726,N_18943,N_18710);
and U21727 (N_21727,N_15408,N_16530);
nor U21728 (N_21728,N_16963,N_15445);
or U21729 (N_21729,N_18887,N_19478);
nor U21730 (N_21730,N_16181,N_18438);
or U21731 (N_21731,N_19543,N_18309);
or U21732 (N_21732,N_18154,N_18781);
and U21733 (N_21733,N_16858,N_16418);
or U21734 (N_21734,N_19802,N_19882);
nor U21735 (N_21735,N_17994,N_17143);
nand U21736 (N_21736,N_17629,N_15186);
and U21737 (N_21737,N_17033,N_18670);
nand U21738 (N_21738,N_19050,N_16788);
and U21739 (N_21739,N_18123,N_17578);
nor U21740 (N_21740,N_15129,N_17186);
and U21741 (N_21741,N_19979,N_17255);
or U21742 (N_21742,N_18524,N_15362);
or U21743 (N_21743,N_18940,N_18410);
and U21744 (N_21744,N_19141,N_15813);
and U21745 (N_21745,N_17476,N_15012);
nor U21746 (N_21746,N_16768,N_19796);
or U21747 (N_21747,N_15992,N_18443);
nand U21748 (N_21748,N_16932,N_18334);
or U21749 (N_21749,N_17084,N_16272);
or U21750 (N_21750,N_15171,N_16062);
nor U21751 (N_21751,N_15132,N_18053);
xnor U21752 (N_21752,N_15999,N_17545);
or U21753 (N_21753,N_16736,N_19022);
nand U21754 (N_21754,N_17859,N_18488);
and U21755 (N_21755,N_15597,N_19464);
and U21756 (N_21756,N_19109,N_15829);
nand U21757 (N_21757,N_18254,N_16158);
or U21758 (N_21758,N_15016,N_17935);
nand U21759 (N_21759,N_19392,N_19858);
nand U21760 (N_21760,N_15610,N_17624);
or U21761 (N_21761,N_18495,N_19965);
and U21762 (N_21762,N_16397,N_17296);
or U21763 (N_21763,N_17655,N_19551);
or U21764 (N_21764,N_18661,N_17173);
nand U21765 (N_21765,N_15073,N_16090);
or U21766 (N_21766,N_18978,N_19532);
nand U21767 (N_21767,N_18243,N_15167);
nand U21768 (N_21768,N_17502,N_18860);
or U21769 (N_21769,N_15484,N_19789);
and U21770 (N_21770,N_19404,N_19911);
or U21771 (N_21771,N_19027,N_18391);
nor U21772 (N_21772,N_19909,N_19044);
or U21773 (N_21773,N_15076,N_15569);
and U21774 (N_21774,N_15483,N_19969);
nand U21775 (N_21775,N_16036,N_16850);
and U21776 (N_21776,N_16575,N_16204);
or U21777 (N_21777,N_17845,N_18815);
and U21778 (N_21778,N_16744,N_16520);
or U21779 (N_21779,N_16127,N_15137);
or U21780 (N_21780,N_16321,N_19908);
xnor U21781 (N_21781,N_16938,N_18974);
nor U21782 (N_21782,N_19105,N_16010);
nand U21783 (N_21783,N_15598,N_19511);
nor U21784 (N_21784,N_16163,N_16831);
and U21785 (N_21785,N_18162,N_15615);
nand U21786 (N_21786,N_17602,N_18457);
and U21787 (N_21787,N_19612,N_15594);
or U21788 (N_21788,N_19683,N_15298);
nand U21789 (N_21789,N_18350,N_17397);
and U21790 (N_21790,N_17953,N_19646);
or U21791 (N_21791,N_16125,N_19070);
and U21792 (N_21792,N_19530,N_17634);
nor U21793 (N_21793,N_18246,N_15868);
or U21794 (N_21794,N_17775,N_18491);
and U21795 (N_21795,N_17992,N_19176);
and U21796 (N_21796,N_17842,N_16737);
and U21797 (N_21797,N_17176,N_16808);
nand U21798 (N_21798,N_16939,N_16445);
or U21799 (N_21799,N_15353,N_17466);
nand U21800 (N_21800,N_16605,N_17888);
and U21801 (N_21801,N_17420,N_18756);
nand U21802 (N_21802,N_15719,N_15955);
nand U21803 (N_21803,N_18997,N_17269);
or U21804 (N_21804,N_16970,N_15006);
or U21805 (N_21805,N_18618,N_16254);
or U21806 (N_21806,N_19830,N_19444);
or U21807 (N_21807,N_17087,N_18303);
and U21808 (N_21808,N_18310,N_18633);
nor U21809 (N_21809,N_18935,N_16677);
or U21810 (N_21810,N_17099,N_15212);
or U21811 (N_21811,N_17531,N_19010);
or U21812 (N_21812,N_18683,N_15091);
or U21813 (N_21813,N_18916,N_19428);
nor U21814 (N_21814,N_15050,N_17020);
and U21815 (N_21815,N_19071,N_16720);
and U21816 (N_21816,N_16839,N_15367);
nor U21817 (N_21817,N_18794,N_19196);
or U21818 (N_21818,N_15181,N_16874);
nand U21819 (N_21819,N_16121,N_19708);
or U21820 (N_21820,N_18208,N_15550);
and U21821 (N_21821,N_19573,N_16101);
nand U21822 (N_21822,N_17191,N_15681);
nor U21823 (N_21823,N_19680,N_18275);
or U21824 (N_21824,N_18985,N_15792);
or U21825 (N_21825,N_16117,N_19673);
nor U21826 (N_21826,N_15374,N_17750);
and U21827 (N_21827,N_17474,N_19581);
xor U21828 (N_21828,N_18133,N_16998);
nand U21829 (N_21829,N_19194,N_17690);
nor U21830 (N_21830,N_16283,N_15060);
nor U21831 (N_21831,N_16184,N_19146);
and U21832 (N_21832,N_18554,N_17763);
xnor U21833 (N_21833,N_19188,N_16666);
nand U21834 (N_21834,N_19944,N_17156);
nor U21835 (N_21835,N_19329,N_15118);
nor U21836 (N_21836,N_16488,N_18485);
or U21837 (N_21837,N_16852,N_15989);
nand U21838 (N_21838,N_18241,N_18302);
and U21839 (N_21839,N_17461,N_15229);
or U21840 (N_21840,N_16638,N_18786);
nor U21841 (N_21841,N_15338,N_16802);
or U21842 (N_21842,N_15497,N_17005);
nor U21843 (N_21843,N_17882,N_16304);
nor U21844 (N_21844,N_17422,N_17564);
nand U21845 (N_21845,N_18480,N_18248);
nor U21846 (N_21846,N_16332,N_16968);
xor U21847 (N_21847,N_19828,N_19519);
and U21848 (N_21848,N_19888,N_15839);
or U21849 (N_21849,N_15398,N_18126);
nand U21850 (N_21850,N_15306,N_16728);
or U21851 (N_21851,N_15263,N_17952);
nor U21852 (N_21852,N_17050,N_18113);
or U21853 (N_21853,N_17031,N_17976);
and U21854 (N_21854,N_18367,N_17730);
nand U21855 (N_21855,N_19605,N_17149);
nand U21856 (N_21856,N_17209,N_15160);
nand U21857 (N_21857,N_19300,N_19684);
or U21858 (N_21858,N_18813,N_15209);
and U21859 (N_21859,N_18508,N_15549);
nor U21860 (N_21860,N_16155,N_15859);
and U21861 (N_21861,N_19152,N_19752);
nor U21862 (N_21862,N_17765,N_16988);
and U21863 (N_21863,N_18448,N_15973);
or U21864 (N_21864,N_17627,N_15363);
nand U21865 (N_21865,N_19482,N_18020);
nand U21866 (N_21866,N_18417,N_17014);
nor U21867 (N_21867,N_15424,N_17998);
nand U21868 (N_21868,N_19255,N_15447);
nor U21869 (N_21869,N_16671,N_15670);
or U21870 (N_21870,N_16028,N_16951);
nand U21871 (N_21871,N_17167,N_15958);
nor U21872 (N_21872,N_19667,N_15713);
or U21873 (N_21873,N_18741,N_17063);
and U21874 (N_21874,N_19717,N_15612);
nand U21875 (N_21875,N_17600,N_16543);
nand U21876 (N_21876,N_15492,N_15063);
nand U21877 (N_21877,N_16458,N_17746);
nand U21878 (N_21878,N_18404,N_17181);
or U21879 (N_21879,N_18521,N_17193);
nand U21880 (N_21880,N_19170,N_18512);
nor U21881 (N_21881,N_15904,N_19622);
and U21882 (N_21882,N_17724,N_17369);
or U21883 (N_21883,N_19567,N_15004);
nor U21884 (N_21884,N_15730,N_16930);
nor U21885 (N_21885,N_18142,N_17489);
and U21886 (N_21886,N_18317,N_16205);
nand U21887 (N_21887,N_18735,N_15494);
nor U21888 (N_21888,N_18224,N_15703);
nand U21889 (N_21889,N_15156,N_19837);
nor U21890 (N_21890,N_18320,N_15804);
and U21891 (N_21891,N_15791,N_18531);
and U21892 (N_21892,N_17868,N_18484);
nor U21893 (N_21893,N_16278,N_18715);
or U21894 (N_21894,N_18711,N_18121);
nand U21895 (N_21895,N_19244,N_19616);
and U21896 (N_21896,N_17065,N_17041);
nand U21897 (N_21897,N_17510,N_19213);
and U21898 (N_21898,N_16171,N_19487);
xor U21899 (N_21899,N_18381,N_16182);
and U21900 (N_21900,N_17924,N_19150);
or U21901 (N_21901,N_19640,N_19931);
nor U21902 (N_21902,N_18606,N_18372);
nor U21903 (N_21903,N_16714,N_16648);
nor U21904 (N_21904,N_19755,N_19350);
nand U21905 (N_21905,N_17111,N_17188);
nor U21906 (N_21906,N_18000,N_19699);
and U21907 (N_21907,N_17870,N_15453);
xor U21908 (N_21908,N_19647,N_15951);
nand U21909 (N_21909,N_16403,N_17530);
or U21910 (N_21910,N_19094,N_15985);
nor U21911 (N_21911,N_19197,N_19240);
nor U21912 (N_21912,N_18256,N_15476);
nand U21913 (N_21913,N_16755,N_16053);
nor U21914 (N_21914,N_15144,N_17586);
or U21915 (N_21915,N_18876,N_16411);
or U21916 (N_21916,N_18237,N_15111);
nand U21917 (N_21917,N_17798,N_16815);
or U21918 (N_21918,N_16892,N_18624);
nor U21919 (N_21919,N_15382,N_15009);
nand U21920 (N_21920,N_15677,N_19303);
or U21921 (N_21921,N_15125,N_16515);
and U21922 (N_21922,N_17512,N_19919);
nor U21923 (N_21923,N_19920,N_17016);
nor U21924 (N_21924,N_17032,N_19185);
nand U21925 (N_21925,N_15048,N_18366);
nor U21926 (N_21926,N_19660,N_18111);
or U21927 (N_21927,N_17980,N_17871);
nor U21928 (N_21928,N_15375,N_15355);
nor U21929 (N_21929,N_19091,N_15230);
or U21930 (N_21930,N_16027,N_17594);
or U21931 (N_21931,N_15260,N_18216);
nand U21932 (N_21932,N_18986,N_19641);
xnor U21933 (N_21933,N_18015,N_18078);
and U21934 (N_21934,N_18892,N_19154);
and U21935 (N_21935,N_18771,N_17226);
or U21936 (N_21936,N_17468,N_19779);
nand U21937 (N_21937,N_15623,N_15051);
or U21938 (N_21938,N_18875,N_19301);
or U21939 (N_21939,N_19601,N_19825);
or U21940 (N_21940,N_18468,N_19793);
nor U21941 (N_21941,N_19023,N_17864);
and U21942 (N_21942,N_15537,N_17861);
nand U21943 (N_21943,N_18459,N_18902);
and U21944 (N_21944,N_17257,N_17968);
nand U21945 (N_21945,N_16256,N_18007);
nor U21946 (N_21946,N_18189,N_18689);
nor U21947 (N_21947,N_16645,N_15580);
nand U21948 (N_21948,N_16517,N_17355);
and U21949 (N_21949,N_16453,N_19808);
or U21950 (N_21950,N_15139,N_16949);
and U21951 (N_21951,N_15323,N_18637);
xnor U21952 (N_21952,N_16308,N_15225);
and U21953 (N_21953,N_19059,N_15682);
nand U21954 (N_21954,N_18743,N_16327);
or U21955 (N_21955,N_19265,N_15756);
nand U21956 (N_21956,N_19963,N_18413);
nor U21957 (N_21957,N_15505,N_19425);
or U21958 (N_21958,N_17678,N_17659);
or U21959 (N_21959,N_19498,N_15927);
nor U21960 (N_21960,N_18117,N_17608);
and U21961 (N_21961,N_17568,N_17692);
and U21962 (N_21962,N_16669,N_18802);
nand U21963 (N_21963,N_18425,N_15801);
nor U21964 (N_21964,N_16462,N_18289);
nor U21965 (N_21965,N_16514,N_18571);
nand U21966 (N_21966,N_16689,N_18462);
nand U21967 (N_21967,N_15821,N_15043);
and U21968 (N_21968,N_18340,N_19135);
nor U21969 (N_21969,N_15583,N_18917);
and U21970 (N_21970,N_16997,N_19505);
nand U21971 (N_21971,N_17157,N_15889);
and U21972 (N_21972,N_16816,N_15239);
nand U21973 (N_21973,N_17967,N_16993);
and U21974 (N_21974,N_17701,N_19949);
and U21975 (N_21975,N_16484,N_19192);
or U21976 (N_21976,N_16527,N_15062);
xnor U21977 (N_21977,N_19447,N_15450);
and U21978 (N_21978,N_18415,N_15825);
and U21979 (N_21979,N_17101,N_18586);
or U21980 (N_21980,N_16843,N_17601);
nor U21981 (N_21981,N_17819,N_16503);
nor U21982 (N_21982,N_17229,N_17015);
or U21983 (N_21983,N_17349,N_17561);
nand U21984 (N_21984,N_15606,N_19002);
nand U21985 (N_21985,N_15393,N_16919);
and U21986 (N_21986,N_15559,N_18143);
and U21987 (N_21987,N_15977,N_17722);
nand U21988 (N_21988,N_19390,N_16126);
and U21989 (N_21989,N_15135,N_18632);
nor U21990 (N_21990,N_18819,N_16880);
nor U21991 (N_21991,N_17464,N_19700);
or U21992 (N_21992,N_17552,N_18955);
nand U21993 (N_21993,N_15146,N_18731);
nand U21994 (N_21994,N_16722,N_19772);
and U21995 (N_21995,N_18209,N_19507);
and U21996 (N_21996,N_17254,N_19666);
and U21997 (N_21997,N_18884,N_18529);
or U21998 (N_21998,N_19092,N_18076);
and U21999 (N_21999,N_19857,N_19527);
nor U22000 (N_22000,N_15895,N_17752);
nor U22001 (N_22001,N_17142,N_15386);
nand U22002 (N_22002,N_17915,N_17222);
or U22003 (N_22003,N_19361,N_17710);
xnor U22004 (N_22004,N_15608,N_17199);
nor U22005 (N_22005,N_16994,N_18159);
nand U22006 (N_22006,N_16313,N_15934);
or U22007 (N_22007,N_19148,N_18466);
xnor U22008 (N_22008,N_15533,N_16437);
and U22009 (N_22009,N_19167,N_17389);
and U22010 (N_22010,N_16105,N_17583);
nor U22011 (N_22011,N_15286,N_18541);
nand U22012 (N_22012,N_16139,N_15008);
nand U22013 (N_22013,N_18699,N_16252);
or U22014 (N_22014,N_19820,N_19211);
nand U22015 (N_22015,N_19714,N_16936);
nand U22016 (N_22016,N_18017,N_16279);
nand U22017 (N_22017,N_18288,N_17340);
nor U22018 (N_22018,N_18640,N_15436);
nand U22019 (N_22019,N_16992,N_15425);
xnor U22020 (N_22020,N_16037,N_16380);
or U22021 (N_22021,N_16410,N_15534);
and U22022 (N_22022,N_16685,N_16051);
nor U22023 (N_22023,N_16220,N_19242);
and U22024 (N_22024,N_17899,N_15679);
nand U22025 (N_22025,N_19905,N_18449);
nand U22026 (N_22026,N_19804,N_15052);
nor U22027 (N_22027,N_18734,N_16222);
and U22028 (N_22028,N_17274,N_19208);
or U22029 (N_22029,N_15965,N_18773);
nor U22030 (N_22030,N_16322,N_17855);
and U22031 (N_22031,N_15283,N_15796);
or U22032 (N_22032,N_15036,N_17940);
xor U22033 (N_22033,N_16614,N_17024);
and U22034 (N_22034,N_19877,N_16268);
nand U22035 (N_22035,N_18878,N_16372);
or U22036 (N_22036,N_18538,N_17109);
or U22037 (N_22037,N_18705,N_18685);
and U22038 (N_22038,N_15735,N_16431);
nor U22039 (N_22039,N_19729,N_18217);
nor U22040 (N_22040,N_19732,N_16916);
nand U22041 (N_22041,N_19058,N_16676);
nand U22042 (N_22042,N_15308,N_19416);
or U22043 (N_22043,N_18442,N_15590);
nand U22044 (N_22044,N_15925,N_17218);
or U22045 (N_22045,N_15671,N_15942);
or U22046 (N_22046,N_17300,N_16800);
and U22047 (N_22047,N_16890,N_18172);
nor U22048 (N_22048,N_15746,N_17268);
or U22049 (N_22049,N_16902,N_15923);
nor U22050 (N_22050,N_18192,N_17127);
nand U22051 (N_22051,N_16273,N_19236);
and U22052 (N_22052,N_16106,N_18348);
and U22053 (N_22053,N_18934,N_18993);
nand U22054 (N_22054,N_15112,N_17898);
nand U22055 (N_22055,N_15223,N_17662);
nor U22056 (N_22056,N_18937,N_16745);
or U22057 (N_22057,N_15806,N_17432);
or U22058 (N_22058,N_18103,N_15068);
nor U22059 (N_22059,N_17119,N_19088);
nor U22060 (N_22060,N_15320,N_15667);
and U22061 (N_22061,N_16675,N_18319);
nor U22062 (N_22062,N_16586,N_19374);
and U22063 (N_22063,N_15255,N_15401);
nand U22064 (N_22064,N_16743,N_15564);
or U22065 (N_22065,N_17733,N_19774);
and U22066 (N_22066,N_19180,N_17165);
nor U22067 (N_22067,N_15892,N_17894);
nor U22068 (N_22068,N_17415,N_17251);
and U22069 (N_22069,N_18703,N_16798);
or U22070 (N_22070,N_16242,N_15364);
nor U22071 (N_22071,N_17972,N_16786);
nand U22072 (N_22072,N_18409,N_17963);
and U22073 (N_22073,N_17559,N_17125);
nand U22074 (N_22074,N_18129,N_19282);
nand U22075 (N_22075,N_18074,N_18725);
and U22076 (N_22076,N_17542,N_19907);
nand U22077 (N_22077,N_15718,N_18476);
nand U22078 (N_22078,N_17327,N_17912);
nor U22079 (N_22079,N_15197,N_16433);
nand U22080 (N_22080,N_15819,N_15674);
nor U22081 (N_22081,N_18104,N_17211);
or U22082 (N_22082,N_15734,N_19310);
or U22083 (N_22083,N_19113,N_15330);
and U22084 (N_22084,N_16364,N_18265);
or U22085 (N_22085,N_19550,N_16160);
or U22086 (N_22086,N_19414,N_15142);
and U22087 (N_22087,N_15376,N_15540);
or U22088 (N_22088,N_15278,N_16102);
nand U22089 (N_22089,N_16014,N_16475);
nor U22090 (N_22090,N_15138,N_17371);
or U22091 (N_22091,N_19886,N_19957);
nand U22092 (N_22092,N_16340,N_15852);
nand U22093 (N_22093,N_18447,N_16472);
nor U22094 (N_22094,N_19932,N_19770);
nor U22095 (N_22095,N_17067,N_15827);
nand U22096 (N_22096,N_19381,N_15669);
nand U22097 (N_22097,N_15226,N_17250);
nor U22098 (N_22098,N_15902,N_15237);
and U22099 (N_22099,N_19778,N_18798);
nand U22100 (N_22100,N_17902,N_19761);
or U22101 (N_22101,N_19695,N_16033);
nand U22102 (N_22102,N_15488,N_15708);
xor U22103 (N_22103,N_17070,N_18513);
nand U22104 (N_22104,N_15243,N_15075);
nor U22105 (N_22105,N_15912,N_17652);
nor U22106 (N_22106,N_19339,N_15158);
nand U22107 (N_22107,N_18544,N_18464);
or U22108 (N_22108,N_19639,N_16399);
or U22109 (N_22109,N_15512,N_15270);
nand U22110 (N_22110,N_19936,N_17617);
or U22111 (N_22111,N_18290,N_19427);
nor U22112 (N_22112,N_17290,N_15221);
nor U22113 (N_22113,N_19039,N_16346);
nor U22114 (N_22114,N_16908,N_19448);
nand U22115 (N_22115,N_16772,N_19538);
or U22116 (N_22116,N_17128,N_19518);
and U22117 (N_22117,N_15296,N_19162);
or U22118 (N_22118,N_18881,N_19471);
or U22119 (N_22119,N_15407,N_15960);
and U22120 (N_22120,N_15587,N_19106);
nor U22121 (N_22121,N_19763,N_16460);
nor U22122 (N_22122,N_17194,N_19693);
and U22123 (N_22123,N_18752,N_15030);
and U22124 (N_22124,N_18690,N_18474);
nand U22125 (N_22125,N_15783,N_15121);
nand U22126 (N_22126,N_19104,N_15061);
and U22127 (N_22127,N_15751,N_19843);
xor U22128 (N_22128,N_18144,N_17441);
or U22129 (N_22129,N_15511,N_16541);
or U22130 (N_22130,N_19727,N_15287);
and U22131 (N_22131,N_15557,N_18101);
and U22132 (N_22132,N_15334,N_19364);
nand U22133 (N_22133,N_18957,N_18212);
nand U22134 (N_22134,N_15326,N_19093);
or U22135 (N_22135,N_18767,N_18623);
or U22136 (N_22136,N_19927,N_16601);
or U22137 (N_22137,N_18949,N_16682);
and U22138 (N_22138,N_15082,N_18299);
or U22139 (N_22139,N_17160,N_19332);
and U22140 (N_22140,N_17183,N_15561);
or U22141 (N_22141,N_15714,N_19181);
or U22142 (N_22142,N_16757,N_19432);
or U22143 (N_22143,N_16584,N_17862);
nor U22144 (N_22144,N_15666,N_18389);
and U22145 (N_22145,N_17130,N_15368);
or U22146 (N_22146,N_18230,N_16017);
and U22147 (N_22147,N_18611,N_17146);
nand U22148 (N_22148,N_16787,N_18717);
nand U22149 (N_22149,N_19822,N_17492);
and U22150 (N_22150,N_18321,N_18778);
nor U22151 (N_22151,N_19560,N_17438);
or U22152 (N_22152,N_18553,N_15085);
nor U22153 (N_22153,N_18713,N_16868);
or U22154 (N_22154,N_19534,N_19368);
nor U22155 (N_22155,N_16361,N_18106);
nand U22156 (N_22156,N_17540,N_15412);
nor U22157 (N_22157,N_17247,N_19411);
nand U22158 (N_22158,N_17115,N_15678);
or U22159 (N_22159,N_16239,N_19052);
nor U22160 (N_22160,N_15786,N_16739);
nor U22161 (N_22161,N_16571,N_15933);
or U22162 (N_22162,N_17345,N_17593);
and U22163 (N_22163,N_17341,N_18795);
nor U22164 (N_22164,N_19833,N_18185);
and U22165 (N_22165,N_17459,N_18572);
or U22166 (N_22166,N_18347,N_18244);
nor U22167 (N_22167,N_16165,N_17619);
or U22168 (N_22168,N_18011,N_17518);
nand U22169 (N_22169,N_17108,N_16367);
nor U22170 (N_22170,N_17886,N_19521);
and U22171 (N_22171,N_17436,N_17285);
nand U22172 (N_22172,N_17791,N_19266);
and U22173 (N_22173,N_15896,N_17079);
nand U22174 (N_22174,N_17546,N_18945);
or U22175 (N_22175,N_18569,N_18688);
nor U22176 (N_22176,N_19072,N_15435);
nand U22177 (N_22177,N_18354,N_19215);
or U22178 (N_22178,N_16582,N_15266);
and U22179 (N_22179,N_16888,N_15015);
or U22180 (N_22180,N_17284,N_16050);
and U22181 (N_22181,N_18021,N_19494);
or U22182 (N_22182,N_17463,N_16312);
nor U22183 (N_22183,N_19328,N_17409);
or U22184 (N_22184,N_17435,N_15289);
or U22185 (N_22185,N_18965,N_16883);
nand U22186 (N_22186,N_19252,N_16652);
or U22187 (N_22187,N_17190,N_17391);
nor U22188 (N_22188,N_17177,N_19011);
nand U22189 (N_22189,N_16596,N_15441);
or U22190 (N_22190,N_18083,N_16611);
nand U22191 (N_22191,N_18681,N_18383);
and U22192 (N_22192,N_15478,N_19250);
nand U22193 (N_22193,N_16558,N_18398);
or U22194 (N_22194,N_15754,N_19736);
or U22195 (N_22195,N_19490,N_16377);
and U22196 (N_22196,N_18423,N_19096);
or U22197 (N_22197,N_18912,N_19295);
nand U22198 (N_22198,N_17503,N_15620);
nor U22199 (N_22199,N_15437,N_17361);
nand U22200 (N_22200,N_17267,N_19469);
nor U22201 (N_22201,N_17472,N_19378);
nand U22202 (N_22202,N_19933,N_15446);
or U22203 (N_22203,N_18597,N_19293);
or U22204 (N_22204,N_18274,N_16836);
or U22205 (N_22205,N_17615,N_18100);
or U22206 (N_22206,N_18911,N_16639);
or U22207 (N_22207,N_18915,N_19710);
nand U22208 (N_22208,N_15079,N_16108);
or U22209 (N_22209,N_17343,N_17315);
and U22210 (N_22210,N_18272,N_15525);
or U22211 (N_22211,N_16159,N_17278);
and U22212 (N_22212,N_18164,N_19851);
and U22213 (N_22213,N_19261,N_15496);
or U22214 (N_22214,N_17118,N_15027);
or U22215 (N_22215,N_19296,N_15219);
and U22216 (N_22216,N_16607,N_18910);
nor U22217 (N_22217,N_19554,N_18388);
nand U22218 (N_22218,N_15327,N_18035);
and U22219 (N_22219,N_17948,N_16876);
nor U22220 (N_22220,N_15711,N_19737);
nor U22221 (N_22221,N_15772,N_17234);
and U22222 (N_22222,N_19492,N_18967);
or U22223 (N_22223,N_19441,N_19344);
and U22224 (N_22224,N_17485,N_17757);
nor U22225 (N_22225,N_15546,N_18199);
and U22226 (N_22226,N_16122,N_18838);
or U22227 (N_22227,N_19179,N_15489);
nand U22228 (N_22228,N_19650,N_16626);
nand U22229 (N_22229,N_15292,N_18316);
and U22230 (N_22230,N_16557,N_19191);
nor U22231 (N_22231,N_15387,N_18761);
nand U22232 (N_22232,N_19970,N_18839);
or U22233 (N_22233,N_19725,N_18539);
or U22234 (N_22234,N_19306,N_19081);
and U22235 (N_22235,N_18058,N_18696);
and U22236 (N_22236,N_17680,N_19333);
or U22237 (N_22237,N_17786,N_19637);
or U22238 (N_22238,N_18010,N_18279);
and U22239 (N_22239,N_15611,N_19009);
and U22240 (N_22240,N_16921,N_19234);
and U22241 (N_22241,N_15001,N_15506);
nor U22242 (N_22242,N_17937,N_18979);
and U22243 (N_22243,N_18202,N_15140);
nand U22244 (N_22244,N_17155,N_15712);
nor U22245 (N_22245,N_17263,N_15007);
or U22246 (N_22246,N_17840,N_19942);
nand U22247 (N_22247,N_19243,N_17221);
nor U22248 (N_22248,N_16862,N_15562);
and U22249 (N_22249,N_16507,N_15105);
nor U22250 (N_22250,N_17683,N_18489);
or U22251 (N_22251,N_17232,N_18146);
and U22252 (N_22252,N_17524,N_18131);
and U22253 (N_22253,N_15438,N_15642);
or U22254 (N_22254,N_16598,N_17743);
and U22255 (N_22255,N_15826,N_16649);
nor U22256 (N_22256,N_18676,N_18077);
nor U22257 (N_22257,N_16459,N_16712);
nand U22258 (N_22258,N_16578,N_16572);
nor U22259 (N_22259,N_17219,N_18850);
nand U22260 (N_22260,N_17416,N_18493);
nor U22261 (N_22261,N_19719,N_16035);
and U22262 (N_22262,N_16792,N_15189);
nor U22263 (N_22263,N_16491,N_19338);
or U22264 (N_22264,N_19994,N_15415);
nor U22265 (N_22265,N_15516,N_18124);
and U22266 (N_22266,N_19926,N_15267);
and U22267 (N_22267,N_19814,N_15799);
nand U22268 (N_22268,N_16271,N_19483);
nor U22269 (N_22269,N_17298,N_19565);
nor U22270 (N_22270,N_18351,N_17374);
or U22271 (N_22271,N_16989,N_16817);
or U22272 (N_22272,N_18636,N_16944);
or U22273 (N_22273,N_17036,N_16392);
and U22274 (N_22274,N_16211,N_19017);
nand U22275 (N_22275,N_19221,N_18698);
and U22276 (N_22276,N_15081,N_18755);
and U22277 (N_22277,N_16566,N_18176);
or U22278 (N_22278,N_18758,N_17447);
or U22279 (N_22279,N_18999,N_15195);
nand U22280 (N_22280,N_16320,N_19971);
and U22281 (N_22281,N_18855,N_19561);
nand U22282 (N_22282,N_15294,N_18490);
and U22283 (N_22283,N_15781,N_18652);
or U22284 (N_22284,N_17893,N_16000);
and U22285 (N_22285,N_16910,N_19336);
nand U22286 (N_22286,N_18552,N_19869);
or U22287 (N_22287,N_18604,N_16879);
nand U22288 (N_22288,N_18163,N_15998);
nor U22289 (N_22289,N_15701,N_15470);
nand U22290 (N_22290,N_16048,N_16042);
or U22291 (N_22291,N_17372,N_16258);
or U22292 (N_22292,N_16707,N_19467);
nand U22293 (N_22293,N_18086,N_19692);
nor U22294 (N_22294,N_18407,N_15029);
and U22295 (N_22295,N_19506,N_17208);
nor U22296 (N_22296,N_16709,N_18006);
nor U22297 (N_22297,N_16833,N_19401);
or U22298 (N_22298,N_15303,N_16374);
and U22299 (N_22299,N_16138,N_15978);
or U22300 (N_22300,N_18028,N_18362);
or U22301 (N_22301,N_17756,N_18736);
nor U22302 (N_22302,N_16348,N_16478);
nand U22303 (N_22303,N_17844,N_17240);
and U22304 (N_22304,N_15049,N_19015);
nand U22305 (N_22305,N_15022,N_15774);
and U22306 (N_22306,N_15565,N_17996);
nand U22307 (N_22307,N_18702,N_18276);
nand U22308 (N_22308,N_17529,N_19611);
and U22309 (N_22309,N_16907,N_17729);
or U22310 (N_22310,N_15836,N_15088);
and U22311 (N_22311,N_18055,N_18116);
or U22312 (N_22312,N_16215,N_17141);
nand U22313 (N_22313,N_19634,N_15035);
and U22314 (N_22314,N_16318,N_18094);
or U22315 (N_22315,N_17210,N_16442);
nand U22316 (N_22316,N_16521,N_17687);
xnor U22317 (N_22317,N_19631,N_19855);
or U22318 (N_22318,N_15479,N_19635);
or U22319 (N_22319,N_16955,N_19596);
nor U22320 (N_22320,N_16369,N_18788);
and U22321 (N_22321,N_16328,N_16680);
nand U22322 (N_22322,N_16733,N_16869);
or U22323 (N_22323,N_18906,N_19594);
nor U22324 (N_22324,N_17544,N_16903);
nor U22325 (N_22325,N_18894,N_19597);
or U22326 (N_22326,N_19656,N_16581);
nand U22327 (N_22327,N_15115,N_17417);
or U22328 (N_22328,N_19158,N_17637);
nor U22329 (N_22329,N_16834,N_15005);
and U22330 (N_22330,N_16686,N_17344);
and U22331 (N_22331,N_17273,N_19952);
nand U22332 (N_22332,N_16087,N_19376);
nand U22333 (N_22333,N_17259,N_19991);
nand U22334 (N_22334,N_19423,N_16705);
nand U22335 (N_22335,N_19312,N_15486);
or U22336 (N_22336,N_19485,N_18919);
or U22337 (N_22337,N_17703,N_17398);
nand U22338 (N_22338,N_16496,N_18414);
or U22339 (N_22339,N_15917,N_15953);
or U22340 (N_22340,N_19760,N_16047);
nand U22341 (N_22341,N_15883,N_19399);
and U22342 (N_22342,N_17089,N_18727);
nand U22343 (N_22343,N_15944,N_19273);
nand U22344 (N_22344,N_15465,N_16721);
or U22345 (N_22345,N_19625,N_18651);
nand U22346 (N_22346,N_18441,N_17565);
or U22347 (N_22347,N_19147,N_15228);
and U22348 (N_22348,N_17596,N_18561);
and U22349 (N_22349,N_16060,N_15811);
nand U22350 (N_22350,N_17684,N_18568);
or U22351 (N_22351,N_17942,N_17927);
nor U22352 (N_22352,N_15198,N_19964);
nand U22353 (N_22353,N_19322,N_15838);
nand U22354 (N_22354,N_17676,N_19476);
or U22355 (N_22355,N_18032,N_19536);
xnor U22356 (N_22356,N_18068,N_16039);
xnor U22357 (N_22357,N_18723,N_17168);
or U22358 (N_22358,N_17866,N_16219);
and U22359 (N_22359,N_16729,N_19746);
or U22360 (N_22360,N_17833,N_16569);
nor U22361 (N_22361,N_17166,N_19910);
and U22362 (N_22362,N_18666,N_19619);
nor U22363 (N_22363,N_19745,N_16235);
nand U22364 (N_22364,N_19884,N_18903);
and U22365 (N_22365,N_17554,N_19642);
and U22366 (N_22366,N_18733,N_16221);
nor U22367 (N_22367,N_19587,N_15777);
nand U22368 (N_22368,N_15234,N_16249);
nand U22369 (N_22369,N_17555,N_15970);
nand U22370 (N_22370,N_16845,N_15548);
nand U22371 (N_22371,N_17380,N_15074);
and U22372 (N_22372,N_19721,N_19026);
or U22373 (N_22373,N_15740,N_18677);
nor U22374 (N_22374,N_19032,N_15911);
and U22375 (N_22375,N_19840,N_15335);
nand U22376 (N_22376,N_18405,N_19398);
nand U22377 (N_22377,N_16209,N_19599);
nor U22378 (N_22378,N_18555,N_15656);
nand U22379 (N_22379,N_19171,N_17961);
and U22380 (N_22380,N_19125,N_16996);
nor U22381 (N_22381,N_15851,N_19618);
nand U22382 (N_22382,N_16363,N_17856);
nor U22383 (N_22383,N_15377,N_17876);
or U22384 (N_22384,N_18339,N_19183);
nand U22385 (N_22385,N_17444,N_18846);
nand U22386 (N_22386,N_15161,N_17421);
or U22387 (N_22387,N_16269,N_16045);
and U22388 (N_22388,N_17779,N_18149);
nor U22389 (N_22389,N_19491,N_18707);
or U22390 (N_22390,N_16430,N_18874);
or U22391 (N_22391,N_18842,N_18787);
nand U22392 (N_22392,N_19405,N_16898);
and U22393 (N_22393,N_16406,N_17446);
nand U22394 (N_22394,N_17495,N_17025);
or U22395 (N_22395,N_17163,N_17783);
or U22396 (N_22396,N_15560,N_18353);
and U22397 (N_22397,N_18088,N_15331);
nand U22398 (N_22398,N_19155,N_17120);
and U22399 (N_22399,N_15199,N_19149);
nand U22400 (N_22400,N_18235,N_15659);
or U22401 (N_22401,N_16891,N_15487);
nand U22402 (N_22402,N_18098,N_18863);
and U22403 (N_22403,N_17816,N_17930);
or U22404 (N_22404,N_16244,N_17242);
and U22405 (N_22405,N_18332,N_17997);
and U22406 (N_22406,N_19397,N_16153);
and U22407 (N_22407,N_16577,N_18924);
or U22408 (N_22408,N_16009,N_18180);
nand U22409 (N_22409,N_19950,N_18868);
or U22410 (N_22410,N_17096,N_16842);
nor U22411 (N_22411,N_19281,N_18535);
nor U22412 (N_22412,N_17605,N_18127);
or U22413 (N_22413,N_18298,N_18760);
nand U22414 (N_22414,N_17658,N_16849);
or U22415 (N_22415,N_16701,N_15104);
or U22416 (N_22416,N_17650,N_17216);
and U22417 (N_22417,N_18746,N_17821);
and U22418 (N_22418,N_16567,N_17717);
nand U22419 (N_22419,N_17801,N_18570);
nor U22420 (N_22420,N_18282,N_19520);
and U22421 (N_22421,N_18888,N_18556);
nand U22422 (N_22422,N_17839,N_16362);
or U22423 (N_22423,N_17411,N_16703);
nand U22424 (N_22424,N_15743,N_19247);
and U22425 (N_22425,N_17837,N_18900);
nand U22426 (N_22426,N_19585,N_18954);
or U22427 (N_22427,N_19636,N_16487);
or U22428 (N_22428,N_15120,N_15552);
nor U22429 (N_22429,N_16455,N_19391);
and U22430 (N_22430,N_16554,N_17956);
or U22431 (N_22431,N_17570,N_15739);
nand U22432 (N_22432,N_15727,N_16079);
or U22433 (N_22433,N_17511,N_17006);
or U22434 (N_22434,N_19302,N_19290);
and U22435 (N_22435,N_16448,N_17906);
and U22436 (N_22436,N_16173,N_18013);
nor U22437 (N_22437,N_16389,N_19626);
nor U22438 (N_22438,N_15510,N_17803);
nand U22439 (N_22439,N_15639,N_18072);
or U22440 (N_22440,N_18675,N_16446);
or U22441 (N_22441,N_15259,N_18177);
and U22442 (N_22442,N_17780,N_19468);
and U22443 (N_22443,N_16508,N_18238);
nor U22444 (N_22444,N_17702,N_15526);
or U22445 (N_22445,N_19571,N_18181);
nand U22446 (N_22446,N_18393,N_17486);
and U22447 (N_22447,N_16147,N_15592);
and U22448 (N_22448,N_17831,N_15241);
or U22449 (N_22449,N_19020,N_19880);
or U22450 (N_22450,N_16600,N_19402);
or U22451 (N_22451,N_17431,N_18811);
nand U22452 (N_22452,N_17453,N_17085);
and U22453 (N_22453,N_16641,N_17301);
or U22454 (N_22454,N_16111,N_15481);
nand U22455 (N_22455,N_15390,N_15893);
and U22456 (N_22456,N_17865,N_15581);
and U22457 (N_22457,N_15462,N_15647);
nor U22458 (N_22458,N_19080,N_17517);
nor U22459 (N_22459,N_17647,N_15910);
xor U22460 (N_22460,N_15311,N_16054);
nand U22461 (N_22461,N_18259,N_18486);
or U22462 (N_22462,N_18578,N_19199);
and U22463 (N_22463,N_15686,N_19604);
nor U22464 (N_22464,N_19895,N_18161);
xnor U22465 (N_22465,N_17616,N_15887);
nor U22466 (N_22466,N_15418,N_17774);
and U22467 (N_22467,N_16495,N_16260);
and U22468 (N_22468,N_19318,N_17525);
or U22469 (N_22469,N_17874,N_18740);
or U22470 (N_22470,N_17197,N_19419);
nand U22471 (N_22471,N_16284,N_19062);
nor U22472 (N_22472,N_19028,N_16494);
or U22473 (N_22473,N_17951,N_17584);
and U22474 (N_22474,N_16388,N_15213);
nand U22475 (N_22475,N_16972,N_15544);
and U22476 (N_22476,N_19885,N_17093);
and U22477 (N_22477,N_18686,N_19189);
nor U22478 (N_22478,N_17003,N_17116);
or U22479 (N_22479,N_15943,N_18004);
nor U22480 (N_22480,N_16386,N_19202);
or U22481 (N_22481,N_15672,N_19718);
and U22482 (N_22482,N_18519,N_19298);
nand U22483 (N_22483,N_18091,N_17741);
or U22484 (N_22484,N_18203,N_17749);
or U22485 (N_22485,N_16749,N_18505);
or U22486 (N_22486,N_17978,N_19029);
and U22487 (N_22487,N_16797,N_19086);
nand U22488 (N_22488,N_15881,N_17751);
nor U22489 (N_22489,N_17346,N_18845);
or U22490 (N_22490,N_17401,N_19362);
nand U22491 (N_22491,N_16473,N_17761);
nor U22492 (N_22492,N_17734,N_19292);
or U22493 (N_22493,N_18872,N_15463);
or U22494 (N_22494,N_19829,N_16451);
or U22495 (N_22495,N_17553,N_18994);
and U22496 (N_22496,N_16065,N_19048);
and U22497 (N_22497,N_16595,N_15729);
nor U22498 (N_22498,N_15369,N_16840);
nor U22499 (N_22499,N_18822,N_16653);
nand U22500 (N_22500,N_15430,N_18144);
or U22501 (N_22501,N_19640,N_16098);
nand U22502 (N_22502,N_19022,N_19338);
or U22503 (N_22503,N_16414,N_16216);
and U22504 (N_22504,N_19286,N_19043);
nand U22505 (N_22505,N_16821,N_17916);
nor U22506 (N_22506,N_17560,N_18495);
or U22507 (N_22507,N_16236,N_17621);
and U22508 (N_22508,N_18953,N_17046);
nand U22509 (N_22509,N_16918,N_17875);
and U22510 (N_22510,N_19752,N_17701);
and U22511 (N_22511,N_16219,N_17584);
and U22512 (N_22512,N_18992,N_17670);
nor U22513 (N_22513,N_18983,N_18825);
nand U22514 (N_22514,N_17755,N_19070);
or U22515 (N_22515,N_16801,N_18052);
or U22516 (N_22516,N_15215,N_16947);
and U22517 (N_22517,N_17595,N_15834);
or U22518 (N_22518,N_16778,N_19429);
nor U22519 (N_22519,N_19691,N_19704);
or U22520 (N_22520,N_15745,N_16035);
nand U22521 (N_22521,N_16393,N_15816);
nor U22522 (N_22522,N_16922,N_19481);
nand U22523 (N_22523,N_18724,N_19391);
or U22524 (N_22524,N_16548,N_16752);
nand U22525 (N_22525,N_19452,N_16474);
and U22526 (N_22526,N_18890,N_19592);
nor U22527 (N_22527,N_18030,N_15435);
and U22528 (N_22528,N_16101,N_16725);
nor U22529 (N_22529,N_15664,N_15213);
nand U22530 (N_22530,N_17710,N_15076);
nand U22531 (N_22531,N_17891,N_15016);
nand U22532 (N_22532,N_18211,N_18056);
nand U22533 (N_22533,N_18526,N_19180);
and U22534 (N_22534,N_15655,N_18164);
nor U22535 (N_22535,N_15306,N_17481);
and U22536 (N_22536,N_18850,N_17486);
nand U22537 (N_22537,N_16479,N_19929);
nand U22538 (N_22538,N_15124,N_16072);
nor U22539 (N_22539,N_18473,N_15852);
and U22540 (N_22540,N_19042,N_19739);
or U22541 (N_22541,N_17395,N_19700);
or U22542 (N_22542,N_18946,N_17105);
nor U22543 (N_22543,N_18435,N_16877);
nand U22544 (N_22544,N_16319,N_19636);
nor U22545 (N_22545,N_17841,N_17813);
nor U22546 (N_22546,N_16200,N_19454);
nor U22547 (N_22547,N_18231,N_15463);
nand U22548 (N_22548,N_15286,N_18289);
xnor U22549 (N_22549,N_19123,N_16976);
nor U22550 (N_22550,N_17180,N_18233);
nor U22551 (N_22551,N_18089,N_18999);
and U22552 (N_22552,N_16313,N_15367);
and U22553 (N_22553,N_16355,N_18166);
nand U22554 (N_22554,N_17602,N_19434);
nor U22555 (N_22555,N_16337,N_16621);
nor U22556 (N_22556,N_15953,N_18694);
nand U22557 (N_22557,N_19535,N_16494);
nor U22558 (N_22558,N_15821,N_17887);
nor U22559 (N_22559,N_18465,N_19276);
nand U22560 (N_22560,N_16039,N_15024);
nand U22561 (N_22561,N_16936,N_15946);
and U22562 (N_22562,N_18462,N_18886);
or U22563 (N_22563,N_17893,N_18156);
or U22564 (N_22564,N_19521,N_18283);
and U22565 (N_22565,N_15959,N_15756);
nand U22566 (N_22566,N_15573,N_17895);
nand U22567 (N_22567,N_19588,N_18275);
nand U22568 (N_22568,N_15421,N_18347);
nor U22569 (N_22569,N_17116,N_16822);
nand U22570 (N_22570,N_17376,N_19041);
or U22571 (N_22571,N_15006,N_19673);
nor U22572 (N_22572,N_16089,N_16728);
or U22573 (N_22573,N_17613,N_17229);
and U22574 (N_22574,N_16646,N_16550);
or U22575 (N_22575,N_16820,N_19306);
and U22576 (N_22576,N_19113,N_18384);
or U22577 (N_22577,N_16132,N_18298);
nand U22578 (N_22578,N_15266,N_16255);
and U22579 (N_22579,N_17355,N_18873);
nand U22580 (N_22580,N_18531,N_17072);
and U22581 (N_22581,N_16059,N_15371);
or U22582 (N_22582,N_15093,N_18698);
nand U22583 (N_22583,N_15449,N_17778);
or U22584 (N_22584,N_18956,N_16955);
or U22585 (N_22585,N_18680,N_16612);
and U22586 (N_22586,N_18010,N_17913);
nand U22587 (N_22587,N_16414,N_18466);
and U22588 (N_22588,N_17648,N_16275);
and U22589 (N_22589,N_15040,N_17659);
and U22590 (N_22590,N_19970,N_18699);
nand U22591 (N_22591,N_18590,N_18110);
nor U22592 (N_22592,N_15008,N_17222);
nor U22593 (N_22593,N_16082,N_16572);
nand U22594 (N_22594,N_18903,N_17977);
and U22595 (N_22595,N_15190,N_19903);
and U22596 (N_22596,N_19874,N_16871);
nor U22597 (N_22597,N_18726,N_19876);
and U22598 (N_22598,N_19560,N_18994);
nand U22599 (N_22599,N_15191,N_15245);
or U22600 (N_22600,N_18494,N_18679);
nand U22601 (N_22601,N_15131,N_18108);
nand U22602 (N_22602,N_19176,N_19281);
and U22603 (N_22603,N_16605,N_15957);
and U22604 (N_22604,N_19830,N_19358);
and U22605 (N_22605,N_17727,N_16624);
nor U22606 (N_22606,N_18426,N_15278);
and U22607 (N_22607,N_15248,N_15068);
or U22608 (N_22608,N_15710,N_15915);
nand U22609 (N_22609,N_16093,N_17431);
or U22610 (N_22610,N_17229,N_15427);
and U22611 (N_22611,N_18815,N_19816);
or U22612 (N_22612,N_16245,N_17893);
nor U22613 (N_22613,N_18431,N_15978);
and U22614 (N_22614,N_18241,N_18226);
nand U22615 (N_22615,N_17305,N_17119);
nand U22616 (N_22616,N_19572,N_16254);
nand U22617 (N_22617,N_15637,N_16084);
nor U22618 (N_22618,N_15823,N_19392);
nor U22619 (N_22619,N_19308,N_19972);
or U22620 (N_22620,N_18917,N_15269);
nor U22621 (N_22621,N_16951,N_19681);
or U22622 (N_22622,N_15675,N_17058);
and U22623 (N_22623,N_16925,N_15451);
nor U22624 (N_22624,N_17568,N_18776);
nor U22625 (N_22625,N_19659,N_18938);
or U22626 (N_22626,N_19125,N_16314);
or U22627 (N_22627,N_17443,N_15116);
nor U22628 (N_22628,N_17932,N_17380);
and U22629 (N_22629,N_17776,N_18419);
or U22630 (N_22630,N_16909,N_16480);
nand U22631 (N_22631,N_19180,N_15639);
xor U22632 (N_22632,N_19386,N_16710);
or U22633 (N_22633,N_18973,N_16828);
and U22634 (N_22634,N_19206,N_18669);
and U22635 (N_22635,N_16006,N_15006);
or U22636 (N_22636,N_18482,N_17204);
or U22637 (N_22637,N_15021,N_16397);
and U22638 (N_22638,N_16779,N_19485);
nand U22639 (N_22639,N_16742,N_15556);
nor U22640 (N_22640,N_16566,N_19644);
nand U22641 (N_22641,N_18566,N_18417);
and U22642 (N_22642,N_16584,N_17223);
nand U22643 (N_22643,N_18323,N_19517);
nand U22644 (N_22644,N_18540,N_19173);
xor U22645 (N_22645,N_18188,N_16289);
and U22646 (N_22646,N_16630,N_19536);
or U22647 (N_22647,N_18454,N_15464);
or U22648 (N_22648,N_18732,N_19107);
nand U22649 (N_22649,N_15274,N_19887);
and U22650 (N_22650,N_19232,N_19635);
or U22651 (N_22651,N_19469,N_15640);
and U22652 (N_22652,N_19023,N_18535);
and U22653 (N_22653,N_17526,N_16977);
xor U22654 (N_22654,N_16783,N_15705);
and U22655 (N_22655,N_18841,N_17844);
nand U22656 (N_22656,N_15657,N_17243);
nor U22657 (N_22657,N_18175,N_19552);
or U22658 (N_22658,N_15721,N_17952);
or U22659 (N_22659,N_19390,N_15067);
nand U22660 (N_22660,N_15837,N_18219);
nand U22661 (N_22661,N_15537,N_16575);
nand U22662 (N_22662,N_18747,N_15006);
and U22663 (N_22663,N_19181,N_18962);
nor U22664 (N_22664,N_19161,N_15508);
and U22665 (N_22665,N_15512,N_18179);
xnor U22666 (N_22666,N_17912,N_15446);
nand U22667 (N_22667,N_16672,N_17712);
or U22668 (N_22668,N_18757,N_15984);
or U22669 (N_22669,N_15993,N_17681);
and U22670 (N_22670,N_19431,N_16862);
and U22671 (N_22671,N_16210,N_19984);
nand U22672 (N_22672,N_19048,N_17263);
or U22673 (N_22673,N_18629,N_19632);
and U22674 (N_22674,N_16337,N_19426);
nand U22675 (N_22675,N_19746,N_16059);
nor U22676 (N_22676,N_19387,N_19833);
nor U22677 (N_22677,N_17492,N_16515);
and U22678 (N_22678,N_19742,N_16746);
and U22679 (N_22679,N_17224,N_18362);
and U22680 (N_22680,N_19463,N_18665);
or U22681 (N_22681,N_15951,N_19682);
and U22682 (N_22682,N_16435,N_16775);
and U22683 (N_22683,N_16717,N_15058);
or U22684 (N_22684,N_16841,N_19296);
and U22685 (N_22685,N_17559,N_16395);
nor U22686 (N_22686,N_19961,N_15535);
nor U22687 (N_22687,N_16639,N_15717);
and U22688 (N_22688,N_19686,N_16743);
nor U22689 (N_22689,N_19062,N_15608);
or U22690 (N_22690,N_18720,N_17736);
and U22691 (N_22691,N_19303,N_16757);
or U22692 (N_22692,N_16115,N_15805);
or U22693 (N_22693,N_16843,N_18436);
or U22694 (N_22694,N_19752,N_18763);
nand U22695 (N_22695,N_16678,N_15336);
and U22696 (N_22696,N_19653,N_19588);
or U22697 (N_22697,N_16652,N_18584);
or U22698 (N_22698,N_16726,N_15824);
and U22699 (N_22699,N_18659,N_19395);
xor U22700 (N_22700,N_17888,N_17042);
and U22701 (N_22701,N_17220,N_19276);
nor U22702 (N_22702,N_16114,N_17973);
or U22703 (N_22703,N_18592,N_16206);
or U22704 (N_22704,N_19259,N_15792);
nand U22705 (N_22705,N_18272,N_16742);
and U22706 (N_22706,N_19855,N_17878);
or U22707 (N_22707,N_16319,N_17759);
and U22708 (N_22708,N_17952,N_16257);
and U22709 (N_22709,N_18710,N_17728);
and U22710 (N_22710,N_19489,N_16807);
and U22711 (N_22711,N_19686,N_19671);
or U22712 (N_22712,N_17443,N_15624);
nand U22713 (N_22713,N_17438,N_19623);
nor U22714 (N_22714,N_16393,N_18866);
or U22715 (N_22715,N_18003,N_19289);
nor U22716 (N_22716,N_16092,N_15456);
or U22717 (N_22717,N_18696,N_19446);
nor U22718 (N_22718,N_17792,N_16890);
nand U22719 (N_22719,N_17656,N_16959);
or U22720 (N_22720,N_16925,N_15894);
nand U22721 (N_22721,N_15448,N_17541);
and U22722 (N_22722,N_18002,N_16670);
nand U22723 (N_22723,N_19366,N_17898);
nor U22724 (N_22724,N_19663,N_19451);
nand U22725 (N_22725,N_18592,N_18152);
or U22726 (N_22726,N_19193,N_19377);
nor U22727 (N_22727,N_16206,N_17976);
or U22728 (N_22728,N_18480,N_15740);
or U22729 (N_22729,N_18636,N_16161);
or U22730 (N_22730,N_16078,N_19152);
nand U22731 (N_22731,N_15140,N_18621);
nor U22732 (N_22732,N_18624,N_16301);
or U22733 (N_22733,N_15831,N_19428);
and U22734 (N_22734,N_19696,N_15028);
nand U22735 (N_22735,N_16623,N_16381);
xnor U22736 (N_22736,N_16716,N_15328);
nor U22737 (N_22737,N_19713,N_16131);
and U22738 (N_22738,N_16411,N_16856);
and U22739 (N_22739,N_16593,N_15533);
or U22740 (N_22740,N_15410,N_19820);
nand U22741 (N_22741,N_19967,N_16042);
nor U22742 (N_22742,N_15112,N_17094);
and U22743 (N_22743,N_15504,N_15048);
nor U22744 (N_22744,N_16968,N_17923);
nor U22745 (N_22745,N_15734,N_18797);
nor U22746 (N_22746,N_19125,N_19033);
nor U22747 (N_22747,N_19395,N_16704);
nand U22748 (N_22748,N_18467,N_15841);
nor U22749 (N_22749,N_16172,N_18423);
or U22750 (N_22750,N_16349,N_18054);
nand U22751 (N_22751,N_19364,N_16970);
or U22752 (N_22752,N_15120,N_19371);
or U22753 (N_22753,N_16629,N_15811);
or U22754 (N_22754,N_18462,N_15438);
or U22755 (N_22755,N_19213,N_16974);
and U22756 (N_22756,N_17889,N_15529);
and U22757 (N_22757,N_17441,N_16406);
and U22758 (N_22758,N_17652,N_19710);
and U22759 (N_22759,N_17470,N_15016);
and U22760 (N_22760,N_16250,N_19813);
and U22761 (N_22761,N_16598,N_18315);
or U22762 (N_22762,N_19997,N_16325);
nor U22763 (N_22763,N_15490,N_15235);
and U22764 (N_22764,N_18641,N_19735);
nor U22765 (N_22765,N_15459,N_19920);
or U22766 (N_22766,N_17538,N_15366);
nand U22767 (N_22767,N_19630,N_19146);
and U22768 (N_22768,N_16290,N_16741);
nand U22769 (N_22769,N_15090,N_16737);
nand U22770 (N_22770,N_17664,N_16011);
or U22771 (N_22771,N_16248,N_15647);
or U22772 (N_22772,N_18474,N_19471);
or U22773 (N_22773,N_17503,N_15921);
nor U22774 (N_22774,N_19624,N_17548);
nor U22775 (N_22775,N_16396,N_17846);
or U22776 (N_22776,N_15426,N_19775);
and U22777 (N_22777,N_17065,N_16398);
nor U22778 (N_22778,N_18970,N_17301);
and U22779 (N_22779,N_18460,N_18279);
or U22780 (N_22780,N_18685,N_19162);
and U22781 (N_22781,N_18385,N_15343);
or U22782 (N_22782,N_19773,N_15587);
nand U22783 (N_22783,N_18420,N_15159);
xnor U22784 (N_22784,N_18529,N_17259);
or U22785 (N_22785,N_15883,N_15688);
and U22786 (N_22786,N_17230,N_17715);
and U22787 (N_22787,N_18450,N_15997);
or U22788 (N_22788,N_19554,N_18296);
and U22789 (N_22789,N_18751,N_19601);
and U22790 (N_22790,N_17836,N_18535);
nor U22791 (N_22791,N_15537,N_18631);
nor U22792 (N_22792,N_15952,N_17433);
nand U22793 (N_22793,N_16767,N_18329);
xor U22794 (N_22794,N_17089,N_16047);
nor U22795 (N_22795,N_16922,N_18411);
nand U22796 (N_22796,N_18064,N_18366);
or U22797 (N_22797,N_17594,N_18188);
and U22798 (N_22798,N_19389,N_16275);
and U22799 (N_22799,N_17880,N_18905);
nand U22800 (N_22800,N_15413,N_19549);
nand U22801 (N_22801,N_18625,N_18736);
nand U22802 (N_22802,N_18004,N_18662);
nor U22803 (N_22803,N_19471,N_18131);
nand U22804 (N_22804,N_19984,N_17505);
and U22805 (N_22805,N_19784,N_18787);
and U22806 (N_22806,N_17328,N_19149);
nand U22807 (N_22807,N_17569,N_16765);
and U22808 (N_22808,N_17972,N_17302);
xor U22809 (N_22809,N_19169,N_17807);
or U22810 (N_22810,N_18790,N_18726);
or U22811 (N_22811,N_16480,N_19055);
or U22812 (N_22812,N_17233,N_18731);
or U22813 (N_22813,N_17165,N_15600);
nand U22814 (N_22814,N_19153,N_15836);
or U22815 (N_22815,N_18141,N_16670);
nor U22816 (N_22816,N_17182,N_16987);
nor U22817 (N_22817,N_15339,N_15974);
nor U22818 (N_22818,N_19811,N_19483);
nand U22819 (N_22819,N_19202,N_18796);
nand U22820 (N_22820,N_19769,N_15658);
nor U22821 (N_22821,N_17025,N_16376);
nor U22822 (N_22822,N_16789,N_19491);
nand U22823 (N_22823,N_18271,N_16688);
or U22824 (N_22824,N_15586,N_15582);
and U22825 (N_22825,N_19924,N_19000);
and U22826 (N_22826,N_17391,N_16171);
or U22827 (N_22827,N_17162,N_19226);
or U22828 (N_22828,N_17800,N_19983);
and U22829 (N_22829,N_16612,N_15804);
nor U22830 (N_22830,N_19952,N_17755);
and U22831 (N_22831,N_18062,N_17402);
nor U22832 (N_22832,N_17005,N_19506);
and U22833 (N_22833,N_17430,N_15826);
or U22834 (N_22834,N_15082,N_17077);
and U22835 (N_22835,N_16953,N_15022);
nor U22836 (N_22836,N_19681,N_19363);
nand U22837 (N_22837,N_17273,N_17528);
or U22838 (N_22838,N_16521,N_18679);
nor U22839 (N_22839,N_18402,N_17152);
and U22840 (N_22840,N_18905,N_17204);
or U22841 (N_22841,N_15476,N_15389);
nor U22842 (N_22842,N_17741,N_19542);
or U22843 (N_22843,N_15684,N_17281);
or U22844 (N_22844,N_16317,N_16627);
or U22845 (N_22845,N_19433,N_19732);
and U22846 (N_22846,N_17653,N_16313);
or U22847 (N_22847,N_15344,N_19093);
nor U22848 (N_22848,N_19065,N_19918);
or U22849 (N_22849,N_15049,N_19350);
nor U22850 (N_22850,N_18328,N_18506);
nor U22851 (N_22851,N_17051,N_16167);
nand U22852 (N_22852,N_17570,N_15401);
nand U22853 (N_22853,N_15238,N_16420);
and U22854 (N_22854,N_17356,N_18426);
or U22855 (N_22855,N_17756,N_15310);
xor U22856 (N_22856,N_19765,N_19754);
or U22857 (N_22857,N_19639,N_17344);
nand U22858 (N_22858,N_19586,N_15182);
and U22859 (N_22859,N_18880,N_16669);
nor U22860 (N_22860,N_15643,N_16383);
and U22861 (N_22861,N_17506,N_16315);
and U22862 (N_22862,N_18769,N_19081);
and U22863 (N_22863,N_19539,N_19323);
or U22864 (N_22864,N_15581,N_17615);
nand U22865 (N_22865,N_16859,N_19883);
nand U22866 (N_22866,N_18203,N_16920);
and U22867 (N_22867,N_15244,N_19140);
nand U22868 (N_22868,N_16843,N_19040);
nand U22869 (N_22869,N_17919,N_16883);
nor U22870 (N_22870,N_16171,N_17030);
or U22871 (N_22871,N_18920,N_15061);
and U22872 (N_22872,N_19133,N_16751);
and U22873 (N_22873,N_18002,N_16281);
nand U22874 (N_22874,N_15631,N_16305);
nand U22875 (N_22875,N_15001,N_16192);
and U22876 (N_22876,N_17060,N_19376);
and U22877 (N_22877,N_15570,N_15851);
and U22878 (N_22878,N_15946,N_18709);
and U22879 (N_22879,N_16904,N_18844);
or U22880 (N_22880,N_17853,N_15443);
and U22881 (N_22881,N_18794,N_17192);
or U22882 (N_22882,N_18522,N_19301);
xor U22883 (N_22883,N_16672,N_18164);
nand U22884 (N_22884,N_19509,N_16146);
and U22885 (N_22885,N_18958,N_17502);
nand U22886 (N_22886,N_15643,N_15773);
nand U22887 (N_22887,N_15951,N_15070);
and U22888 (N_22888,N_17061,N_16676);
nor U22889 (N_22889,N_18349,N_15404);
xnor U22890 (N_22890,N_16784,N_15778);
or U22891 (N_22891,N_16622,N_17619);
nor U22892 (N_22892,N_16181,N_16563);
nor U22893 (N_22893,N_15621,N_17751);
and U22894 (N_22894,N_17699,N_17106);
nand U22895 (N_22895,N_16090,N_17952);
xor U22896 (N_22896,N_18642,N_16575);
nand U22897 (N_22897,N_19364,N_18422);
xnor U22898 (N_22898,N_18108,N_16270);
nor U22899 (N_22899,N_18140,N_17923);
nand U22900 (N_22900,N_19195,N_15139);
nand U22901 (N_22901,N_15201,N_16749);
or U22902 (N_22902,N_16269,N_19082);
or U22903 (N_22903,N_17021,N_17540);
nor U22904 (N_22904,N_18677,N_15304);
and U22905 (N_22905,N_19219,N_15081);
nand U22906 (N_22906,N_17581,N_18241);
or U22907 (N_22907,N_17501,N_17134);
nand U22908 (N_22908,N_15962,N_15527);
or U22909 (N_22909,N_16474,N_16476);
and U22910 (N_22910,N_16995,N_19196);
nand U22911 (N_22911,N_17641,N_16645);
nand U22912 (N_22912,N_19719,N_18776);
nor U22913 (N_22913,N_18576,N_19414);
and U22914 (N_22914,N_16768,N_17327);
and U22915 (N_22915,N_16158,N_19420);
nand U22916 (N_22916,N_16409,N_18429);
nand U22917 (N_22917,N_19076,N_19420);
nand U22918 (N_22918,N_19672,N_17285);
nand U22919 (N_22919,N_18324,N_15732);
and U22920 (N_22920,N_16466,N_16876);
nand U22921 (N_22921,N_19040,N_16256);
nand U22922 (N_22922,N_19704,N_18570);
or U22923 (N_22923,N_17707,N_17643);
and U22924 (N_22924,N_18672,N_15765);
nand U22925 (N_22925,N_15575,N_19056);
nor U22926 (N_22926,N_18135,N_19216);
and U22927 (N_22927,N_15913,N_15201);
and U22928 (N_22928,N_19533,N_19082);
and U22929 (N_22929,N_15483,N_18867);
and U22930 (N_22930,N_17627,N_18953);
nor U22931 (N_22931,N_17960,N_19668);
nor U22932 (N_22932,N_19473,N_15898);
and U22933 (N_22933,N_15746,N_17161);
nor U22934 (N_22934,N_18447,N_16827);
nand U22935 (N_22935,N_18013,N_16295);
or U22936 (N_22936,N_17163,N_16762);
nand U22937 (N_22937,N_16344,N_18975);
nand U22938 (N_22938,N_16132,N_16084);
nand U22939 (N_22939,N_17040,N_15585);
or U22940 (N_22940,N_19159,N_19734);
and U22941 (N_22941,N_16956,N_19212);
nor U22942 (N_22942,N_15501,N_17417);
and U22943 (N_22943,N_16011,N_17234);
nor U22944 (N_22944,N_19216,N_15547);
and U22945 (N_22945,N_19516,N_19096);
or U22946 (N_22946,N_18148,N_19302);
nand U22947 (N_22947,N_15364,N_15964);
and U22948 (N_22948,N_17049,N_17578);
nand U22949 (N_22949,N_15802,N_19222);
nor U22950 (N_22950,N_18607,N_19070);
or U22951 (N_22951,N_17842,N_19438);
and U22952 (N_22952,N_16829,N_16489);
and U22953 (N_22953,N_17451,N_16450);
or U22954 (N_22954,N_17343,N_17632);
nor U22955 (N_22955,N_18189,N_19186);
nor U22956 (N_22956,N_16662,N_18190);
nand U22957 (N_22957,N_18749,N_18691);
or U22958 (N_22958,N_16483,N_18394);
and U22959 (N_22959,N_16099,N_15998);
and U22960 (N_22960,N_18854,N_16219);
and U22961 (N_22961,N_19230,N_19827);
and U22962 (N_22962,N_17653,N_15256);
nand U22963 (N_22963,N_15652,N_17084);
nand U22964 (N_22964,N_18520,N_18273);
nand U22965 (N_22965,N_19874,N_17447);
or U22966 (N_22966,N_18764,N_18864);
nand U22967 (N_22967,N_18012,N_17248);
nor U22968 (N_22968,N_16750,N_17829);
or U22969 (N_22969,N_18376,N_18387);
or U22970 (N_22970,N_17182,N_16523);
and U22971 (N_22971,N_18653,N_16472);
nand U22972 (N_22972,N_18023,N_19967);
and U22973 (N_22973,N_18758,N_16794);
or U22974 (N_22974,N_19203,N_19616);
and U22975 (N_22975,N_19871,N_19525);
or U22976 (N_22976,N_16499,N_19806);
nor U22977 (N_22977,N_16280,N_18313);
and U22978 (N_22978,N_17624,N_16105);
nand U22979 (N_22979,N_17337,N_15083);
and U22980 (N_22980,N_15426,N_17160);
or U22981 (N_22981,N_16128,N_19976);
or U22982 (N_22982,N_15607,N_18845);
and U22983 (N_22983,N_18856,N_16064);
and U22984 (N_22984,N_15146,N_16169);
or U22985 (N_22985,N_16325,N_19032);
nor U22986 (N_22986,N_19889,N_15515);
or U22987 (N_22987,N_16326,N_19936);
nor U22988 (N_22988,N_18164,N_16373);
nor U22989 (N_22989,N_15923,N_19490);
and U22990 (N_22990,N_19624,N_17680);
nor U22991 (N_22991,N_17805,N_18747);
nand U22992 (N_22992,N_16235,N_18383);
nand U22993 (N_22993,N_18644,N_15727);
or U22994 (N_22994,N_18475,N_17049);
or U22995 (N_22995,N_17989,N_15220);
or U22996 (N_22996,N_16284,N_18858);
and U22997 (N_22997,N_18012,N_16136);
nor U22998 (N_22998,N_16922,N_17863);
nor U22999 (N_22999,N_19440,N_19239);
and U23000 (N_23000,N_15387,N_15015);
xnor U23001 (N_23001,N_15759,N_17055);
nand U23002 (N_23002,N_19233,N_18949);
nor U23003 (N_23003,N_19001,N_17590);
nand U23004 (N_23004,N_17841,N_18178);
nand U23005 (N_23005,N_19455,N_15760);
nand U23006 (N_23006,N_18114,N_16806);
nand U23007 (N_23007,N_17984,N_19740);
nand U23008 (N_23008,N_17354,N_17044);
nor U23009 (N_23009,N_17314,N_16427);
nor U23010 (N_23010,N_15493,N_15014);
nand U23011 (N_23011,N_19228,N_16659);
nand U23012 (N_23012,N_15026,N_19368);
and U23013 (N_23013,N_17345,N_15243);
or U23014 (N_23014,N_19695,N_18869);
xor U23015 (N_23015,N_17548,N_18683);
and U23016 (N_23016,N_18503,N_16129);
and U23017 (N_23017,N_19728,N_16372);
nand U23018 (N_23018,N_18414,N_17257);
and U23019 (N_23019,N_19211,N_19296);
nand U23020 (N_23020,N_16403,N_17701);
or U23021 (N_23021,N_17015,N_18353);
nand U23022 (N_23022,N_17993,N_17061);
or U23023 (N_23023,N_16656,N_19373);
nand U23024 (N_23024,N_16266,N_19101);
nand U23025 (N_23025,N_15011,N_19807);
or U23026 (N_23026,N_18621,N_19986);
or U23027 (N_23027,N_18843,N_18215);
nor U23028 (N_23028,N_17684,N_18921);
nand U23029 (N_23029,N_19472,N_19571);
or U23030 (N_23030,N_19353,N_16337);
nor U23031 (N_23031,N_19470,N_18977);
nor U23032 (N_23032,N_15059,N_19599);
nand U23033 (N_23033,N_19697,N_18304);
or U23034 (N_23034,N_15286,N_16875);
or U23035 (N_23035,N_19721,N_19555);
nand U23036 (N_23036,N_18841,N_18877);
or U23037 (N_23037,N_16109,N_19317);
nor U23038 (N_23038,N_19979,N_18507);
nor U23039 (N_23039,N_16272,N_17719);
nor U23040 (N_23040,N_19066,N_15728);
nand U23041 (N_23041,N_16469,N_16566);
nor U23042 (N_23042,N_19274,N_19125);
or U23043 (N_23043,N_15275,N_17895);
nand U23044 (N_23044,N_15796,N_19385);
xor U23045 (N_23045,N_17135,N_17853);
xnor U23046 (N_23046,N_17916,N_18924);
or U23047 (N_23047,N_16856,N_19376);
and U23048 (N_23048,N_18983,N_17578);
and U23049 (N_23049,N_18015,N_15121);
or U23050 (N_23050,N_18698,N_19740);
and U23051 (N_23051,N_15153,N_17957);
or U23052 (N_23052,N_16356,N_16251);
or U23053 (N_23053,N_16184,N_15527);
nor U23054 (N_23054,N_17269,N_15570);
or U23055 (N_23055,N_18457,N_15549);
nand U23056 (N_23056,N_18873,N_15656);
nor U23057 (N_23057,N_15408,N_16815);
nor U23058 (N_23058,N_15626,N_16451);
nor U23059 (N_23059,N_19830,N_16748);
and U23060 (N_23060,N_17477,N_16541);
and U23061 (N_23061,N_16301,N_17648);
and U23062 (N_23062,N_17530,N_16510);
and U23063 (N_23063,N_17221,N_18627);
nand U23064 (N_23064,N_16345,N_17332);
and U23065 (N_23065,N_15079,N_15732);
nor U23066 (N_23066,N_18500,N_19396);
nor U23067 (N_23067,N_19770,N_16992);
and U23068 (N_23068,N_18861,N_15586);
or U23069 (N_23069,N_16346,N_17431);
nand U23070 (N_23070,N_19312,N_19499);
and U23071 (N_23071,N_17678,N_19453);
nor U23072 (N_23072,N_19646,N_17249);
and U23073 (N_23073,N_17191,N_17023);
nor U23074 (N_23074,N_15876,N_16951);
and U23075 (N_23075,N_18937,N_15167);
nor U23076 (N_23076,N_19146,N_15740);
or U23077 (N_23077,N_16008,N_18403);
nand U23078 (N_23078,N_18687,N_16588);
nand U23079 (N_23079,N_19873,N_16863);
nand U23080 (N_23080,N_18959,N_16577);
nor U23081 (N_23081,N_16704,N_18033);
xor U23082 (N_23082,N_17389,N_17978);
or U23083 (N_23083,N_16762,N_17968);
and U23084 (N_23084,N_18559,N_17934);
nand U23085 (N_23085,N_19549,N_15929);
nor U23086 (N_23086,N_18988,N_17250);
nor U23087 (N_23087,N_19218,N_17993);
or U23088 (N_23088,N_19980,N_18713);
or U23089 (N_23089,N_19801,N_15600);
nor U23090 (N_23090,N_18913,N_16778);
and U23091 (N_23091,N_18914,N_17657);
nand U23092 (N_23092,N_16880,N_16193);
nor U23093 (N_23093,N_16290,N_15671);
nand U23094 (N_23094,N_17261,N_15790);
nor U23095 (N_23095,N_17574,N_18315);
and U23096 (N_23096,N_15374,N_16606);
or U23097 (N_23097,N_19970,N_17146);
and U23098 (N_23098,N_15625,N_16129);
and U23099 (N_23099,N_15926,N_16140);
or U23100 (N_23100,N_19662,N_16929);
or U23101 (N_23101,N_16236,N_19601);
xnor U23102 (N_23102,N_17528,N_18037);
nor U23103 (N_23103,N_18844,N_17731);
nor U23104 (N_23104,N_15411,N_18940);
and U23105 (N_23105,N_16531,N_19905);
and U23106 (N_23106,N_17256,N_19307);
nand U23107 (N_23107,N_16469,N_16908);
nor U23108 (N_23108,N_15978,N_18264);
and U23109 (N_23109,N_16985,N_18318);
nand U23110 (N_23110,N_18069,N_15135);
and U23111 (N_23111,N_15267,N_17096);
xor U23112 (N_23112,N_19942,N_17985);
or U23113 (N_23113,N_19085,N_18541);
or U23114 (N_23114,N_15484,N_19059);
nor U23115 (N_23115,N_18870,N_16253);
and U23116 (N_23116,N_19482,N_16695);
nand U23117 (N_23117,N_16942,N_18476);
xor U23118 (N_23118,N_15947,N_18258);
or U23119 (N_23119,N_15833,N_18951);
or U23120 (N_23120,N_16939,N_17052);
nand U23121 (N_23121,N_18038,N_16347);
nor U23122 (N_23122,N_17809,N_16581);
nand U23123 (N_23123,N_16432,N_18923);
nor U23124 (N_23124,N_17620,N_16556);
or U23125 (N_23125,N_17319,N_16548);
nor U23126 (N_23126,N_17665,N_17669);
nand U23127 (N_23127,N_18836,N_15038);
or U23128 (N_23128,N_16655,N_16411);
nand U23129 (N_23129,N_18512,N_18736);
or U23130 (N_23130,N_15407,N_16849);
nand U23131 (N_23131,N_17241,N_19544);
or U23132 (N_23132,N_19230,N_15965);
or U23133 (N_23133,N_16976,N_17671);
nand U23134 (N_23134,N_18529,N_17162);
nor U23135 (N_23135,N_18037,N_16381);
or U23136 (N_23136,N_16213,N_18171);
nor U23137 (N_23137,N_17351,N_16735);
or U23138 (N_23138,N_16296,N_19615);
or U23139 (N_23139,N_16552,N_15815);
or U23140 (N_23140,N_17718,N_16449);
and U23141 (N_23141,N_19746,N_15340);
nand U23142 (N_23142,N_19088,N_17256);
nor U23143 (N_23143,N_17549,N_17804);
nand U23144 (N_23144,N_17515,N_18294);
xnor U23145 (N_23145,N_19764,N_15900);
xnor U23146 (N_23146,N_18926,N_18255);
nand U23147 (N_23147,N_15381,N_15304);
and U23148 (N_23148,N_15278,N_17416);
or U23149 (N_23149,N_19778,N_17534);
nand U23150 (N_23150,N_19196,N_18502);
or U23151 (N_23151,N_18237,N_16965);
nor U23152 (N_23152,N_17387,N_19521);
and U23153 (N_23153,N_15537,N_19754);
nor U23154 (N_23154,N_19474,N_15074);
and U23155 (N_23155,N_16494,N_15609);
or U23156 (N_23156,N_17993,N_16718);
or U23157 (N_23157,N_15081,N_18480);
nor U23158 (N_23158,N_16242,N_17270);
or U23159 (N_23159,N_18798,N_16761);
nand U23160 (N_23160,N_18265,N_19042);
nand U23161 (N_23161,N_18703,N_19024);
nand U23162 (N_23162,N_15501,N_17512);
and U23163 (N_23163,N_17345,N_17862);
xnor U23164 (N_23164,N_17146,N_15928);
and U23165 (N_23165,N_19712,N_18722);
or U23166 (N_23166,N_16845,N_15517);
nand U23167 (N_23167,N_17154,N_16695);
or U23168 (N_23168,N_16676,N_17369);
nand U23169 (N_23169,N_15608,N_19264);
nand U23170 (N_23170,N_19929,N_15373);
and U23171 (N_23171,N_18442,N_18846);
and U23172 (N_23172,N_17002,N_17186);
and U23173 (N_23173,N_15921,N_17588);
nand U23174 (N_23174,N_15976,N_18894);
or U23175 (N_23175,N_19719,N_18316);
nor U23176 (N_23176,N_19748,N_19777);
and U23177 (N_23177,N_16022,N_17863);
nand U23178 (N_23178,N_16335,N_18282);
and U23179 (N_23179,N_17764,N_15680);
and U23180 (N_23180,N_15520,N_19623);
nor U23181 (N_23181,N_18824,N_19765);
and U23182 (N_23182,N_15682,N_19418);
nor U23183 (N_23183,N_17169,N_15352);
nand U23184 (N_23184,N_15717,N_15530);
and U23185 (N_23185,N_17364,N_19869);
or U23186 (N_23186,N_17369,N_18950);
and U23187 (N_23187,N_16112,N_18327);
or U23188 (N_23188,N_19577,N_15022);
and U23189 (N_23189,N_18153,N_15242);
and U23190 (N_23190,N_16349,N_19200);
nor U23191 (N_23191,N_19046,N_15180);
or U23192 (N_23192,N_17417,N_17521);
nand U23193 (N_23193,N_16704,N_16495);
nand U23194 (N_23194,N_18398,N_15296);
nand U23195 (N_23195,N_16817,N_15125);
or U23196 (N_23196,N_15017,N_19270);
nor U23197 (N_23197,N_17143,N_16488);
nand U23198 (N_23198,N_18860,N_18862);
nor U23199 (N_23199,N_19167,N_17177);
and U23200 (N_23200,N_19804,N_17694);
or U23201 (N_23201,N_15159,N_15733);
and U23202 (N_23202,N_18299,N_15232);
or U23203 (N_23203,N_17578,N_16159);
or U23204 (N_23204,N_18633,N_18179);
nand U23205 (N_23205,N_18662,N_16345);
or U23206 (N_23206,N_18418,N_16083);
or U23207 (N_23207,N_16009,N_18997);
and U23208 (N_23208,N_19882,N_19586);
or U23209 (N_23209,N_15034,N_19266);
nor U23210 (N_23210,N_17394,N_17972);
nor U23211 (N_23211,N_15726,N_15848);
and U23212 (N_23212,N_19598,N_17353);
or U23213 (N_23213,N_15508,N_18135);
or U23214 (N_23214,N_18282,N_15722);
nor U23215 (N_23215,N_18125,N_17067);
and U23216 (N_23216,N_19637,N_19530);
and U23217 (N_23217,N_19190,N_19141);
nor U23218 (N_23218,N_17249,N_15424);
nand U23219 (N_23219,N_18855,N_17897);
nand U23220 (N_23220,N_19587,N_15625);
nor U23221 (N_23221,N_16915,N_19960);
nor U23222 (N_23222,N_18334,N_15440);
nor U23223 (N_23223,N_16330,N_17060);
or U23224 (N_23224,N_19744,N_18119);
and U23225 (N_23225,N_19670,N_19574);
and U23226 (N_23226,N_16295,N_16012);
and U23227 (N_23227,N_17637,N_17128);
or U23228 (N_23228,N_19796,N_19712);
and U23229 (N_23229,N_16273,N_18670);
nand U23230 (N_23230,N_16855,N_15375);
or U23231 (N_23231,N_16999,N_19726);
or U23232 (N_23232,N_18912,N_18541);
nand U23233 (N_23233,N_15669,N_17590);
or U23234 (N_23234,N_16020,N_15894);
or U23235 (N_23235,N_18301,N_18067);
nand U23236 (N_23236,N_16966,N_18762);
and U23237 (N_23237,N_19039,N_18237);
or U23238 (N_23238,N_15402,N_18077);
nand U23239 (N_23239,N_16409,N_15224);
and U23240 (N_23240,N_17967,N_17669);
nand U23241 (N_23241,N_16594,N_18760);
and U23242 (N_23242,N_15889,N_17798);
and U23243 (N_23243,N_15881,N_15423);
nand U23244 (N_23244,N_19422,N_15213);
or U23245 (N_23245,N_19316,N_15692);
nor U23246 (N_23246,N_15383,N_16227);
nand U23247 (N_23247,N_18781,N_16779);
nand U23248 (N_23248,N_17972,N_17365);
and U23249 (N_23249,N_15506,N_19845);
nand U23250 (N_23250,N_15112,N_15420);
nand U23251 (N_23251,N_15602,N_17216);
or U23252 (N_23252,N_19786,N_18507);
xor U23253 (N_23253,N_16180,N_15810);
nor U23254 (N_23254,N_19113,N_15169);
and U23255 (N_23255,N_15507,N_18767);
nand U23256 (N_23256,N_17079,N_18544);
or U23257 (N_23257,N_16461,N_15009);
and U23258 (N_23258,N_16971,N_16300);
and U23259 (N_23259,N_17146,N_16929);
nor U23260 (N_23260,N_15103,N_18729);
and U23261 (N_23261,N_19116,N_15021);
nand U23262 (N_23262,N_17624,N_15475);
nand U23263 (N_23263,N_16165,N_15013);
or U23264 (N_23264,N_17582,N_17208);
or U23265 (N_23265,N_15444,N_19959);
nor U23266 (N_23266,N_17445,N_17106);
or U23267 (N_23267,N_16927,N_18273);
or U23268 (N_23268,N_16262,N_16164);
nand U23269 (N_23269,N_16331,N_16673);
and U23270 (N_23270,N_15152,N_18162);
nand U23271 (N_23271,N_19645,N_18322);
xnor U23272 (N_23272,N_15793,N_18731);
nor U23273 (N_23273,N_16653,N_18705);
nand U23274 (N_23274,N_19001,N_15271);
nor U23275 (N_23275,N_17029,N_16481);
nand U23276 (N_23276,N_15281,N_15141);
and U23277 (N_23277,N_19780,N_15212);
or U23278 (N_23278,N_16950,N_18452);
nor U23279 (N_23279,N_16671,N_19505);
and U23280 (N_23280,N_15383,N_18816);
nor U23281 (N_23281,N_17301,N_15416);
nand U23282 (N_23282,N_16082,N_15735);
and U23283 (N_23283,N_18839,N_18593);
or U23284 (N_23284,N_19597,N_18149);
and U23285 (N_23285,N_17381,N_18687);
nor U23286 (N_23286,N_15442,N_15184);
and U23287 (N_23287,N_19047,N_16667);
nor U23288 (N_23288,N_15053,N_18039);
nor U23289 (N_23289,N_19461,N_17524);
nor U23290 (N_23290,N_15662,N_19608);
nand U23291 (N_23291,N_17756,N_17701);
or U23292 (N_23292,N_15835,N_19047);
nand U23293 (N_23293,N_16469,N_17407);
and U23294 (N_23294,N_18370,N_15199);
nor U23295 (N_23295,N_19500,N_17600);
or U23296 (N_23296,N_19044,N_19994);
or U23297 (N_23297,N_15790,N_19584);
or U23298 (N_23298,N_18594,N_18950);
nand U23299 (N_23299,N_19750,N_19956);
and U23300 (N_23300,N_16961,N_18751);
or U23301 (N_23301,N_18149,N_18019);
and U23302 (N_23302,N_15291,N_15874);
nand U23303 (N_23303,N_19465,N_16072);
and U23304 (N_23304,N_19782,N_16399);
or U23305 (N_23305,N_19724,N_15051);
or U23306 (N_23306,N_17499,N_19012);
and U23307 (N_23307,N_17769,N_18899);
nor U23308 (N_23308,N_18870,N_16898);
nand U23309 (N_23309,N_17387,N_15036);
nand U23310 (N_23310,N_15474,N_17600);
and U23311 (N_23311,N_18412,N_16127);
nand U23312 (N_23312,N_15358,N_16398);
nor U23313 (N_23313,N_17891,N_19140);
or U23314 (N_23314,N_15112,N_17478);
nor U23315 (N_23315,N_18940,N_16393);
or U23316 (N_23316,N_19741,N_18329);
and U23317 (N_23317,N_17464,N_16812);
nor U23318 (N_23318,N_18029,N_15053);
xor U23319 (N_23319,N_18856,N_18125);
nand U23320 (N_23320,N_19029,N_15968);
and U23321 (N_23321,N_17771,N_17642);
or U23322 (N_23322,N_18163,N_18858);
nor U23323 (N_23323,N_15389,N_17899);
nand U23324 (N_23324,N_19468,N_16670);
or U23325 (N_23325,N_15723,N_19067);
nor U23326 (N_23326,N_17965,N_16037);
nor U23327 (N_23327,N_18221,N_18883);
and U23328 (N_23328,N_18856,N_17889);
or U23329 (N_23329,N_17859,N_17120);
or U23330 (N_23330,N_18634,N_18371);
nand U23331 (N_23331,N_19936,N_16793);
and U23332 (N_23332,N_15414,N_19538);
nand U23333 (N_23333,N_16931,N_16824);
nand U23334 (N_23334,N_18485,N_19116);
nand U23335 (N_23335,N_19510,N_18617);
nor U23336 (N_23336,N_19036,N_17051);
nand U23337 (N_23337,N_19128,N_17205);
xnor U23338 (N_23338,N_16369,N_16207);
nor U23339 (N_23339,N_16509,N_16564);
and U23340 (N_23340,N_16678,N_17250);
or U23341 (N_23341,N_16330,N_17827);
nor U23342 (N_23342,N_16394,N_17355);
or U23343 (N_23343,N_18697,N_19358);
nor U23344 (N_23344,N_19803,N_19492);
nand U23345 (N_23345,N_18203,N_18835);
nand U23346 (N_23346,N_17264,N_18689);
and U23347 (N_23347,N_18447,N_18100);
or U23348 (N_23348,N_15453,N_16628);
xnor U23349 (N_23349,N_15058,N_15978);
or U23350 (N_23350,N_19134,N_15970);
or U23351 (N_23351,N_19966,N_18372);
nor U23352 (N_23352,N_19026,N_15121);
and U23353 (N_23353,N_17811,N_19493);
and U23354 (N_23354,N_17627,N_19509);
xnor U23355 (N_23355,N_17403,N_16265);
nand U23356 (N_23356,N_17186,N_15752);
or U23357 (N_23357,N_17624,N_16689);
and U23358 (N_23358,N_16155,N_18329);
and U23359 (N_23359,N_15738,N_18116);
nor U23360 (N_23360,N_18806,N_17001);
or U23361 (N_23361,N_15410,N_15678);
nand U23362 (N_23362,N_15447,N_18878);
nand U23363 (N_23363,N_18828,N_18248);
nor U23364 (N_23364,N_15898,N_19777);
nor U23365 (N_23365,N_15786,N_15410);
nor U23366 (N_23366,N_17853,N_17140);
nor U23367 (N_23367,N_17002,N_15097);
or U23368 (N_23368,N_17423,N_17084);
or U23369 (N_23369,N_18500,N_15915);
and U23370 (N_23370,N_15496,N_19971);
nor U23371 (N_23371,N_15789,N_16215);
nand U23372 (N_23372,N_16444,N_16047);
nor U23373 (N_23373,N_15192,N_19841);
nor U23374 (N_23374,N_19827,N_17567);
nand U23375 (N_23375,N_19427,N_17797);
or U23376 (N_23376,N_17826,N_17639);
nand U23377 (N_23377,N_17554,N_16983);
and U23378 (N_23378,N_19106,N_16014);
nor U23379 (N_23379,N_15619,N_16720);
nor U23380 (N_23380,N_15638,N_16943);
nand U23381 (N_23381,N_19318,N_18729);
nor U23382 (N_23382,N_17457,N_16225);
and U23383 (N_23383,N_19715,N_18997);
or U23384 (N_23384,N_16252,N_18382);
nand U23385 (N_23385,N_17296,N_16602);
and U23386 (N_23386,N_17384,N_16734);
and U23387 (N_23387,N_17590,N_17105);
nand U23388 (N_23388,N_16817,N_16642);
or U23389 (N_23389,N_18603,N_17305);
or U23390 (N_23390,N_17388,N_19500);
xor U23391 (N_23391,N_17965,N_19438);
xnor U23392 (N_23392,N_16912,N_15358);
and U23393 (N_23393,N_18457,N_16658);
xor U23394 (N_23394,N_16816,N_17232);
or U23395 (N_23395,N_19333,N_15461);
nand U23396 (N_23396,N_15039,N_17483);
nor U23397 (N_23397,N_15691,N_16590);
or U23398 (N_23398,N_16423,N_19619);
nor U23399 (N_23399,N_18639,N_19506);
nand U23400 (N_23400,N_15993,N_17566);
and U23401 (N_23401,N_17177,N_17456);
nand U23402 (N_23402,N_15593,N_18057);
nand U23403 (N_23403,N_19766,N_18359);
nand U23404 (N_23404,N_18830,N_17335);
and U23405 (N_23405,N_15444,N_19438);
and U23406 (N_23406,N_19833,N_17775);
nor U23407 (N_23407,N_15911,N_17625);
or U23408 (N_23408,N_18853,N_18326);
xnor U23409 (N_23409,N_16194,N_16225);
and U23410 (N_23410,N_19624,N_18836);
or U23411 (N_23411,N_17808,N_19994);
or U23412 (N_23412,N_16884,N_16730);
nor U23413 (N_23413,N_15309,N_15659);
nor U23414 (N_23414,N_18851,N_19004);
nand U23415 (N_23415,N_18749,N_15149);
nor U23416 (N_23416,N_15555,N_18775);
or U23417 (N_23417,N_19457,N_15449);
nor U23418 (N_23418,N_17438,N_15261);
nand U23419 (N_23419,N_17412,N_19044);
nor U23420 (N_23420,N_17225,N_17812);
nand U23421 (N_23421,N_15421,N_17540);
and U23422 (N_23422,N_18554,N_18639);
or U23423 (N_23423,N_17492,N_19581);
nor U23424 (N_23424,N_15774,N_15199);
and U23425 (N_23425,N_17843,N_15273);
nand U23426 (N_23426,N_19624,N_15605);
and U23427 (N_23427,N_15557,N_19747);
nor U23428 (N_23428,N_15925,N_19725);
or U23429 (N_23429,N_18867,N_15916);
nor U23430 (N_23430,N_17241,N_16400);
and U23431 (N_23431,N_17943,N_17769);
nand U23432 (N_23432,N_16321,N_19580);
and U23433 (N_23433,N_15029,N_17962);
xor U23434 (N_23434,N_16865,N_16974);
nor U23435 (N_23435,N_16880,N_19503);
and U23436 (N_23436,N_16873,N_16124);
nor U23437 (N_23437,N_17248,N_16777);
nand U23438 (N_23438,N_17057,N_17654);
or U23439 (N_23439,N_18577,N_15821);
nor U23440 (N_23440,N_17348,N_16871);
and U23441 (N_23441,N_16547,N_18541);
or U23442 (N_23442,N_16274,N_17080);
nand U23443 (N_23443,N_17931,N_15142);
nor U23444 (N_23444,N_19668,N_18793);
nand U23445 (N_23445,N_19865,N_15423);
and U23446 (N_23446,N_19269,N_19545);
and U23447 (N_23447,N_19881,N_17275);
nor U23448 (N_23448,N_17940,N_15636);
and U23449 (N_23449,N_19373,N_15863);
nand U23450 (N_23450,N_15945,N_19076);
and U23451 (N_23451,N_18693,N_17220);
or U23452 (N_23452,N_17550,N_16662);
nand U23453 (N_23453,N_17328,N_17230);
and U23454 (N_23454,N_15489,N_19988);
or U23455 (N_23455,N_15777,N_18501);
and U23456 (N_23456,N_16204,N_15125);
or U23457 (N_23457,N_19421,N_16309);
nand U23458 (N_23458,N_18827,N_15366);
and U23459 (N_23459,N_18031,N_16018);
nor U23460 (N_23460,N_15117,N_19080);
nand U23461 (N_23461,N_19418,N_16863);
nand U23462 (N_23462,N_16671,N_17457);
and U23463 (N_23463,N_18410,N_15047);
nor U23464 (N_23464,N_16891,N_16291);
nor U23465 (N_23465,N_16542,N_15736);
nand U23466 (N_23466,N_18679,N_18766);
nand U23467 (N_23467,N_15891,N_17372);
nor U23468 (N_23468,N_18638,N_18794);
and U23469 (N_23469,N_17889,N_18535);
nor U23470 (N_23470,N_17068,N_15794);
nor U23471 (N_23471,N_16242,N_16178);
and U23472 (N_23472,N_18122,N_16717);
nor U23473 (N_23473,N_19637,N_17190);
or U23474 (N_23474,N_16278,N_15787);
nor U23475 (N_23475,N_19506,N_18628);
nand U23476 (N_23476,N_15245,N_15107);
or U23477 (N_23477,N_19618,N_18375);
nand U23478 (N_23478,N_18596,N_15158);
or U23479 (N_23479,N_19751,N_19053);
nor U23480 (N_23480,N_16788,N_16523);
nor U23481 (N_23481,N_19181,N_19959);
and U23482 (N_23482,N_17734,N_18627);
nor U23483 (N_23483,N_17973,N_18992);
nor U23484 (N_23484,N_16689,N_16549);
or U23485 (N_23485,N_15466,N_15998);
nor U23486 (N_23486,N_17882,N_17910);
nand U23487 (N_23487,N_19628,N_17280);
nor U23488 (N_23488,N_19933,N_18812);
and U23489 (N_23489,N_16577,N_15941);
or U23490 (N_23490,N_17657,N_18595);
and U23491 (N_23491,N_18499,N_16129);
nor U23492 (N_23492,N_15490,N_17812);
or U23493 (N_23493,N_16009,N_19084);
or U23494 (N_23494,N_16648,N_16780);
nor U23495 (N_23495,N_16939,N_19528);
or U23496 (N_23496,N_18335,N_17117);
and U23497 (N_23497,N_19340,N_18906);
nor U23498 (N_23498,N_16758,N_18195);
and U23499 (N_23499,N_16430,N_15796);
or U23500 (N_23500,N_15100,N_15778);
or U23501 (N_23501,N_18213,N_17026);
or U23502 (N_23502,N_18763,N_18268);
nand U23503 (N_23503,N_18676,N_15088);
or U23504 (N_23504,N_15361,N_17934);
nor U23505 (N_23505,N_19218,N_15942);
or U23506 (N_23506,N_19924,N_18102);
and U23507 (N_23507,N_19136,N_19429);
or U23508 (N_23508,N_18107,N_16935);
or U23509 (N_23509,N_17238,N_17007);
or U23510 (N_23510,N_15054,N_17137);
nand U23511 (N_23511,N_18029,N_19689);
or U23512 (N_23512,N_17534,N_19116);
nand U23513 (N_23513,N_19138,N_17741);
nor U23514 (N_23514,N_16828,N_16849);
nor U23515 (N_23515,N_15451,N_19020);
nand U23516 (N_23516,N_18393,N_15377);
nand U23517 (N_23517,N_15201,N_17735);
or U23518 (N_23518,N_16220,N_16999);
or U23519 (N_23519,N_16262,N_16069);
or U23520 (N_23520,N_16940,N_17234);
or U23521 (N_23521,N_15475,N_17284);
xor U23522 (N_23522,N_19728,N_17854);
or U23523 (N_23523,N_18114,N_18735);
and U23524 (N_23524,N_19062,N_16359);
or U23525 (N_23525,N_19932,N_16584);
xor U23526 (N_23526,N_17020,N_17381);
or U23527 (N_23527,N_15177,N_16311);
nand U23528 (N_23528,N_15268,N_18639);
nor U23529 (N_23529,N_17907,N_16454);
or U23530 (N_23530,N_19332,N_18526);
nand U23531 (N_23531,N_15994,N_16676);
nand U23532 (N_23532,N_15419,N_19948);
or U23533 (N_23533,N_17917,N_19574);
xor U23534 (N_23534,N_15868,N_19663);
or U23535 (N_23535,N_17951,N_16437);
or U23536 (N_23536,N_19679,N_16893);
and U23537 (N_23537,N_17794,N_19409);
and U23538 (N_23538,N_15876,N_15130);
nand U23539 (N_23539,N_15388,N_19712);
nand U23540 (N_23540,N_16903,N_18244);
nand U23541 (N_23541,N_18872,N_17114);
nor U23542 (N_23542,N_16468,N_19007);
nand U23543 (N_23543,N_18392,N_18064);
nand U23544 (N_23544,N_15277,N_15679);
and U23545 (N_23545,N_16138,N_17810);
and U23546 (N_23546,N_18186,N_15904);
nand U23547 (N_23547,N_18617,N_17746);
nand U23548 (N_23548,N_16390,N_17859);
nand U23549 (N_23549,N_17369,N_16547);
or U23550 (N_23550,N_16445,N_15974);
nor U23551 (N_23551,N_18966,N_18779);
or U23552 (N_23552,N_19482,N_19881);
and U23553 (N_23553,N_19413,N_15248);
and U23554 (N_23554,N_15442,N_18473);
nor U23555 (N_23555,N_19346,N_19448);
and U23556 (N_23556,N_16700,N_16814);
and U23557 (N_23557,N_15988,N_16646);
and U23558 (N_23558,N_16544,N_15529);
nand U23559 (N_23559,N_18688,N_19214);
and U23560 (N_23560,N_19616,N_19592);
nor U23561 (N_23561,N_18664,N_16365);
nand U23562 (N_23562,N_16324,N_17074);
or U23563 (N_23563,N_19508,N_15738);
and U23564 (N_23564,N_18302,N_18055);
or U23565 (N_23565,N_16549,N_17655);
nor U23566 (N_23566,N_15132,N_15453);
and U23567 (N_23567,N_16908,N_15031);
and U23568 (N_23568,N_15135,N_16521);
and U23569 (N_23569,N_16195,N_18605);
or U23570 (N_23570,N_16089,N_15682);
or U23571 (N_23571,N_19993,N_17924);
nor U23572 (N_23572,N_19774,N_16306);
nor U23573 (N_23573,N_19260,N_19121);
and U23574 (N_23574,N_19938,N_19030);
or U23575 (N_23575,N_16395,N_15884);
or U23576 (N_23576,N_18890,N_17190);
nand U23577 (N_23577,N_18534,N_15179);
nand U23578 (N_23578,N_19579,N_19327);
or U23579 (N_23579,N_19987,N_17041);
and U23580 (N_23580,N_15960,N_19780);
or U23581 (N_23581,N_19549,N_17289);
and U23582 (N_23582,N_15297,N_19584);
and U23583 (N_23583,N_17795,N_19175);
or U23584 (N_23584,N_18552,N_15787);
nand U23585 (N_23585,N_15551,N_17205);
nor U23586 (N_23586,N_16726,N_19827);
and U23587 (N_23587,N_19834,N_19139);
or U23588 (N_23588,N_17030,N_15616);
and U23589 (N_23589,N_18470,N_19152);
nand U23590 (N_23590,N_16856,N_17459);
nand U23591 (N_23591,N_15629,N_16521);
nor U23592 (N_23592,N_15924,N_17330);
xor U23593 (N_23593,N_15724,N_16055);
nor U23594 (N_23594,N_19748,N_18367);
nand U23595 (N_23595,N_17642,N_16950);
and U23596 (N_23596,N_16922,N_18429);
nor U23597 (N_23597,N_15995,N_19116);
or U23598 (N_23598,N_17690,N_18039);
nand U23599 (N_23599,N_19243,N_19971);
nand U23600 (N_23600,N_19438,N_17252);
nor U23601 (N_23601,N_17629,N_16765);
or U23602 (N_23602,N_17254,N_17009);
nand U23603 (N_23603,N_15031,N_17824);
or U23604 (N_23604,N_17015,N_18788);
and U23605 (N_23605,N_17316,N_16787);
and U23606 (N_23606,N_18208,N_19002);
nor U23607 (N_23607,N_19599,N_15942);
nor U23608 (N_23608,N_15731,N_19704);
nand U23609 (N_23609,N_18727,N_15270);
nand U23610 (N_23610,N_15249,N_18135);
and U23611 (N_23611,N_15039,N_19104);
nor U23612 (N_23612,N_16137,N_16196);
nand U23613 (N_23613,N_19026,N_15117);
nor U23614 (N_23614,N_17033,N_16368);
or U23615 (N_23615,N_16797,N_18745);
nor U23616 (N_23616,N_18355,N_15778);
or U23617 (N_23617,N_19664,N_15544);
xnor U23618 (N_23618,N_19251,N_18118);
nand U23619 (N_23619,N_19205,N_15326);
or U23620 (N_23620,N_15431,N_16118);
and U23621 (N_23621,N_18123,N_19799);
nor U23622 (N_23622,N_15116,N_15640);
or U23623 (N_23623,N_19880,N_19184);
and U23624 (N_23624,N_15257,N_17522);
nor U23625 (N_23625,N_16899,N_16135);
xor U23626 (N_23626,N_16703,N_15752);
or U23627 (N_23627,N_15897,N_18967);
nor U23628 (N_23628,N_18233,N_18850);
nand U23629 (N_23629,N_18863,N_16432);
nor U23630 (N_23630,N_15478,N_17717);
nor U23631 (N_23631,N_15555,N_18353);
nor U23632 (N_23632,N_17143,N_19652);
or U23633 (N_23633,N_17157,N_17547);
and U23634 (N_23634,N_15429,N_17731);
nand U23635 (N_23635,N_15744,N_19487);
and U23636 (N_23636,N_16871,N_17582);
or U23637 (N_23637,N_15543,N_18781);
and U23638 (N_23638,N_18727,N_15381);
and U23639 (N_23639,N_16651,N_18676);
and U23640 (N_23640,N_17793,N_19682);
nor U23641 (N_23641,N_17958,N_18490);
or U23642 (N_23642,N_17238,N_15341);
or U23643 (N_23643,N_17716,N_15767);
xnor U23644 (N_23644,N_19665,N_16384);
nor U23645 (N_23645,N_18284,N_19242);
nand U23646 (N_23646,N_16577,N_15158);
nor U23647 (N_23647,N_18675,N_16602);
and U23648 (N_23648,N_19594,N_18897);
nor U23649 (N_23649,N_17182,N_17047);
and U23650 (N_23650,N_16791,N_16191);
nor U23651 (N_23651,N_15955,N_19443);
nand U23652 (N_23652,N_17286,N_18339);
nand U23653 (N_23653,N_16304,N_19440);
nand U23654 (N_23654,N_18242,N_16922);
nand U23655 (N_23655,N_18970,N_19697);
nand U23656 (N_23656,N_18584,N_16125);
or U23657 (N_23657,N_16423,N_17039);
and U23658 (N_23658,N_15473,N_18707);
or U23659 (N_23659,N_15106,N_15170);
and U23660 (N_23660,N_19294,N_18487);
nand U23661 (N_23661,N_19757,N_15089);
and U23662 (N_23662,N_19508,N_19241);
nor U23663 (N_23663,N_15232,N_19697);
nand U23664 (N_23664,N_19155,N_17664);
and U23665 (N_23665,N_16090,N_19870);
and U23666 (N_23666,N_16215,N_19393);
or U23667 (N_23667,N_17345,N_16617);
nand U23668 (N_23668,N_16992,N_17686);
and U23669 (N_23669,N_18333,N_15805);
nand U23670 (N_23670,N_19061,N_16776);
nand U23671 (N_23671,N_19664,N_16580);
and U23672 (N_23672,N_16433,N_15839);
or U23673 (N_23673,N_19351,N_17498);
nor U23674 (N_23674,N_19261,N_15719);
nor U23675 (N_23675,N_16233,N_16984);
nand U23676 (N_23676,N_17700,N_15664);
and U23677 (N_23677,N_16696,N_19850);
or U23678 (N_23678,N_17832,N_15579);
nand U23679 (N_23679,N_18868,N_18320);
nor U23680 (N_23680,N_19773,N_16617);
and U23681 (N_23681,N_15868,N_15446);
nor U23682 (N_23682,N_18636,N_19120);
xnor U23683 (N_23683,N_17363,N_18525);
or U23684 (N_23684,N_18732,N_19152);
nor U23685 (N_23685,N_19439,N_19707);
and U23686 (N_23686,N_17596,N_16851);
nand U23687 (N_23687,N_15356,N_15544);
or U23688 (N_23688,N_18930,N_17550);
nand U23689 (N_23689,N_16699,N_19629);
nand U23690 (N_23690,N_17868,N_19917);
nand U23691 (N_23691,N_16311,N_15321);
nor U23692 (N_23692,N_18189,N_18726);
and U23693 (N_23693,N_19382,N_18987);
and U23694 (N_23694,N_17082,N_15341);
nand U23695 (N_23695,N_18844,N_18163);
and U23696 (N_23696,N_15850,N_15995);
and U23697 (N_23697,N_18826,N_16727);
or U23698 (N_23698,N_16296,N_19149);
nand U23699 (N_23699,N_18522,N_15852);
nor U23700 (N_23700,N_17074,N_17180);
nand U23701 (N_23701,N_19797,N_16035);
or U23702 (N_23702,N_16844,N_17806);
nor U23703 (N_23703,N_15816,N_16131);
and U23704 (N_23704,N_19316,N_17585);
nand U23705 (N_23705,N_18895,N_15408);
nand U23706 (N_23706,N_18075,N_16878);
or U23707 (N_23707,N_16265,N_16679);
or U23708 (N_23708,N_16893,N_17001);
or U23709 (N_23709,N_18730,N_18624);
nand U23710 (N_23710,N_15695,N_15532);
or U23711 (N_23711,N_18692,N_18168);
and U23712 (N_23712,N_15802,N_15585);
nor U23713 (N_23713,N_18112,N_18376);
nor U23714 (N_23714,N_17573,N_17083);
and U23715 (N_23715,N_19489,N_15074);
nand U23716 (N_23716,N_16303,N_19346);
nand U23717 (N_23717,N_16534,N_18340);
nand U23718 (N_23718,N_19887,N_17280);
or U23719 (N_23719,N_16974,N_19526);
and U23720 (N_23720,N_17604,N_16350);
and U23721 (N_23721,N_16002,N_18883);
nand U23722 (N_23722,N_16964,N_17035);
xor U23723 (N_23723,N_15911,N_16357);
or U23724 (N_23724,N_18913,N_15451);
or U23725 (N_23725,N_18342,N_18833);
and U23726 (N_23726,N_18474,N_19533);
or U23727 (N_23727,N_17545,N_19739);
nor U23728 (N_23728,N_15396,N_18269);
nor U23729 (N_23729,N_17489,N_15563);
nor U23730 (N_23730,N_16366,N_17289);
nand U23731 (N_23731,N_18830,N_17927);
nand U23732 (N_23732,N_17267,N_19095);
or U23733 (N_23733,N_18188,N_19836);
or U23734 (N_23734,N_18174,N_16053);
nand U23735 (N_23735,N_17396,N_19898);
nor U23736 (N_23736,N_19385,N_17243);
and U23737 (N_23737,N_19393,N_15653);
and U23738 (N_23738,N_15507,N_18552);
or U23739 (N_23739,N_15821,N_16956);
nor U23740 (N_23740,N_18685,N_18671);
or U23741 (N_23741,N_16975,N_16553);
and U23742 (N_23742,N_17723,N_15464);
nor U23743 (N_23743,N_18934,N_17154);
nor U23744 (N_23744,N_15929,N_18642);
nor U23745 (N_23745,N_16014,N_17184);
nand U23746 (N_23746,N_18557,N_18628);
or U23747 (N_23747,N_17664,N_19367);
or U23748 (N_23748,N_19012,N_16645);
nor U23749 (N_23749,N_15839,N_17392);
nand U23750 (N_23750,N_18759,N_19415);
nor U23751 (N_23751,N_19345,N_17528);
or U23752 (N_23752,N_19686,N_16045);
and U23753 (N_23753,N_19453,N_17508);
and U23754 (N_23754,N_17923,N_18487);
or U23755 (N_23755,N_15867,N_17160);
nand U23756 (N_23756,N_19870,N_18384);
and U23757 (N_23757,N_18373,N_19284);
nand U23758 (N_23758,N_16149,N_18213);
nor U23759 (N_23759,N_15123,N_18017);
nand U23760 (N_23760,N_15752,N_15104);
nor U23761 (N_23761,N_18284,N_16760);
nand U23762 (N_23762,N_18362,N_15563);
or U23763 (N_23763,N_16964,N_15504);
nor U23764 (N_23764,N_18923,N_18571);
or U23765 (N_23765,N_19089,N_16962);
nand U23766 (N_23766,N_15486,N_17097);
nor U23767 (N_23767,N_15742,N_19012);
nor U23768 (N_23768,N_18684,N_15563);
nand U23769 (N_23769,N_18695,N_16833);
nor U23770 (N_23770,N_17368,N_16893);
or U23771 (N_23771,N_15921,N_19559);
nor U23772 (N_23772,N_17820,N_19657);
or U23773 (N_23773,N_19682,N_16133);
or U23774 (N_23774,N_15034,N_19077);
nand U23775 (N_23775,N_16805,N_18794);
or U23776 (N_23776,N_17314,N_15788);
nand U23777 (N_23777,N_18948,N_17979);
nand U23778 (N_23778,N_19776,N_15726);
or U23779 (N_23779,N_17453,N_19445);
nor U23780 (N_23780,N_17520,N_19279);
nand U23781 (N_23781,N_19160,N_19176);
or U23782 (N_23782,N_19746,N_19956);
nand U23783 (N_23783,N_15775,N_19688);
xnor U23784 (N_23784,N_15937,N_18334);
or U23785 (N_23785,N_18747,N_15963);
nand U23786 (N_23786,N_18418,N_15144);
nand U23787 (N_23787,N_19739,N_16888);
nand U23788 (N_23788,N_17356,N_19114);
nor U23789 (N_23789,N_15537,N_16420);
nand U23790 (N_23790,N_18071,N_18499);
nand U23791 (N_23791,N_15085,N_18542);
nand U23792 (N_23792,N_16926,N_16276);
nand U23793 (N_23793,N_19451,N_18904);
or U23794 (N_23794,N_17076,N_15967);
and U23795 (N_23795,N_18752,N_18262);
and U23796 (N_23796,N_16910,N_19472);
and U23797 (N_23797,N_16757,N_19562);
and U23798 (N_23798,N_19219,N_17127);
nor U23799 (N_23799,N_18270,N_18660);
nor U23800 (N_23800,N_16385,N_19933);
nand U23801 (N_23801,N_15102,N_15153);
or U23802 (N_23802,N_16643,N_16500);
or U23803 (N_23803,N_15197,N_15319);
nand U23804 (N_23804,N_19196,N_18488);
nor U23805 (N_23805,N_15623,N_15866);
and U23806 (N_23806,N_16165,N_16870);
nand U23807 (N_23807,N_15046,N_15958);
and U23808 (N_23808,N_19571,N_16003);
nor U23809 (N_23809,N_16002,N_18275);
or U23810 (N_23810,N_16802,N_19184);
or U23811 (N_23811,N_15580,N_16946);
and U23812 (N_23812,N_18767,N_18026);
and U23813 (N_23813,N_15708,N_16580);
and U23814 (N_23814,N_17198,N_16473);
nand U23815 (N_23815,N_15398,N_17597);
or U23816 (N_23816,N_19774,N_19519);
or U23817 (N_23817,N_17246,N_16623);
nor U23818 (N_23818,N_18752,N_19898);
or U23819 (N_23819,N_19827,N_17138);
or U23820 (N_23820,N_16912,N_17718);
and U23821 (N_23821,N_19967,N_15512);
nand U23822 (N_23822,N_15204,N_19760);
and U23823 (N_23823,N_18784,N_17456);
and U23824 (N_23824,N_15470,N_19203);
and U23825 (N_23825,N_16567,N_19438);
and U23826 (N_23826,N_18370,N_19289);
nor U23827 (N_23827,N_15783,N_19669);
and U23828 (N_23828,N_18256,N_18092);
and U23829 (N_23829,N_16345,N_15929);
nand U23830 (N_23830,N_19672,N_18240);
nor U23831 (N_23831,N_16840,N_18772);
and U23832 (N_23832,N_18588,N_17729);
nand U23833 (N_23833,N_16506,N_15440);
nand U23834 (N_23834,N_16328,N_16477);
nand U23835 (N_23835,N_18998,N_18813);
or U23836 (N_23836,N_17617,N_16764);
nand U23837 (N_23837,N_19567,N_18072);
or U23838 (N_23838,N_17492,N_16736);
and U23839 (N_23839,N_16714,N_19679);
or U23840 (N_23840,N_16407,N_19921);
nor U23841 (N_23841,N_18850,N_18126);
and U23842 (N_23842,N_15641,N_16743);
nand U23843 (N_23843,N_15216,N_17814);
nand U23844 (N_23844,N_15189,N_17064);
nor U23845 (N_23845,N_15117,N_16156);
nand U23846 (N_23846,N_16264,N_19861);
and U23847 (N_23847,N_19269,N_17473);
xor U23848 (N_23848,N_18644,N_16852);
nand U23849 (N_23849,N_16290,N_17645);
and U23850 (N_23850,N_18594,N_16405);
and U23851 (N_23851,N_16010,N_19014);
and U23852 (N_23852,N_17780,N_19528);
and U23853 (N_23853,N_18854,N_18409);
or U23854 (N_23854,N_17723,N_15675);
xor U23855 (N_23855,N_17262,N_19841);
nor U23856 (N_23856,N_18221,N_19149);
nand U23857 (N_23857,N_17686,N_16364);
nand U23858 (N_23858,N_16217,N_17046);
nor U23859 (N_23859,N_16997,N_19887);
nand U23860 (N_23860,N_16827,N_18498);
nand U23861 (N_23861,N_17347,N_18972);
and U23862 (N_23862,N_15141,N_19267);
or U23863 (N_23863,N_19659,N_18420);
nor U23864 (N_23864,N_17052,N_16127);
or U23865 (N_23865,N_18853,N_15914);
nor U23866 (N_23866,N_17948,N_19884);
and U23867 (N_23867,N_17246,N_19969);
and U23868 (N_23868,N_17818,N_19114);
or U23869 (N_23869,N_17751,N_17749);
nand U23870 (N_23870,N_16373,N_16175);
nor U23871 (N_23871,N_15339,N_17887);
and U23872 (N_23872,N_17661,N_18747);
and U23873 (N_23873,N_18927,N_15544);
xor U23874 (N_23874,N_17605,N_15275);
xnor U23875 (N_23875,N_15482,N_18768);
nand U23876 (N_23876,N_15179,N_18233);
nand U23877 (N_23877,N_15846,N_15908);
and U23878 (N_23878,N_18258,N_16536);
nand U23879 (N_23879,N_19359,N_15130);
nand U23880 (N_23880,N_15707,N_16959);
nor U23881 (N_23881,N_18910,N_19941);
or U23882 (N_23882,N_16463,N_15866);
or U23883 (N_23883,N_16314,N_18031);
nand U23884 (N_23884,N_19853,N_15170);
and U23885 (N_23885,N_17046,N_18323);
nand U23886 (N_23886,N_16951,N_17337);
or U23887 (N_23887,N_15925,N_16662);
nand U23888 (N_23888,N_17090,N_19415);
nand U23889 (N_23889,N_18913,N_18683);
and U23890 (N_23890,N_16295,N_15563);
and U23891 (N_23891,N_19632,N_17788);
xnor U23892 (N_23892,N_16799,N_15677);
or U23893 (N_23893,N_16595,N_16340);
and U23894 (N_23894,N_19026,N_16072);
nand U23895 (N_23895,N_16082,N_17966);
nor U23896 (N_23896,N_15151,N_15888);
nor U23897 (N_23897,N_17330,N_19754);
or U23898 (N_23898,N_19563,N_19839);
or U23899 (N_23899,N_15542,N_16907);
nor U23900 (N_23900,N_16806,N_16308);
nand U23901 (N_23901,N_18716,N_16850);
nor U23902 (N_23902,N_16426,N_15162);
or U23903 (N_23903,N_18220,N_19892);
nand U23904 (N_23904,N_16938,N_18692);
and U23905 (N_23905,N_18869,N_16293);
or U23906 (N_23906,N_16941,N_18563);
nand U23907 (N_23907,N_18443,N_19611);
nand U23908 (N_23908,N_19372,N_18664);
and U23909 (N_23909,N_17350,N_17361);
nor U23910 (N_23910,N_16167,N_17245);
nand U23911 (N_23911,N_18393,N_16771);
nand U23912 (N_23912,N_17782,N_16608);
or U23913 (N_23913,N_18888,N_16963);
nor U23914 (N_23914,N_15751,N_16484);
and U23915 (N_23915,N_19014,N_17034);
nand U23916 (N_23916,N_19711,N_18583);
nand U23917 (N_23917,N_18514,N_16508);
and U23918 (N_23918,N_16883,N_16501);
or U23919 (N_23919,N_19888,N_16096);
nand U23920 (N_23920,N_15435,N_19528);
nand U23921 (N_23921,N_19386,N_18880);
nor U23922 (N_23922,N_15854,N_15948);
or U23923 (N_23923,N_17693,N_16211);
nand U23924 (N_23924,N_19099,N_16255);
nand U23925 (N_23925,N_19166,N_17031);
nand U23926 (N_23926,N_19455,N_17802);
or U23927 (N_23927,N_17036,N_16271);
or U23928 (N_23928,N_15747,N_15278);
nand U23929 (N_23929,N_19621,N_17306);
xnor U23930 (N_23930,N_15897,N_17481);
nor U23931 (N_23931,N_15046,N_15936);
or U23932 (N_23932,N_18253,N_18325);
nand U23933 (N_23933,N_15874,N_17569);
and U23934 (N_23934,N_16508,N_15616);
nand U23935 (N_23935,N_18342,N_19729);
or U23936 (N_23936,N_19052,N_19047);
and U23937 (N_23937,N_17035,N_18669);
and U23938 (N_23938,N_18631,N_17872);
and U23939 (N_23939,N_18525,N_16799);
nand U23940 (N_23940,N_18498,N_16950);
and U23941 (N_23941,N_19601,N_19134);
nand U23942 (N_23942,N_17027,N_15942);
nand U23943 (N_23943,N_15663,N_19464);
nand U23944 (N_23944,N_17495,N_19583);
nand U23945 (N_23945,N_17787,N_15916);
and U23946 (N_23946,N_19423,N_17709);
and U23947 (N_23947,N_16324,N_17082);
nand U23948 (N_23948,N_16627,N_19790);
and U23949 (N_23949,N_18067,N_17424);
nor U23950 (N_23950,N_18597,N_15411);
and U23951 (N_23951,N_19105,N_19622);
and U23952 (N_23952,N_15645,N_19724);
or U23953 (N_23953,N_18692,N_17374);
nand U23954 (N_23954,N_16092,N_16225);
or U23955 (N_23955,N_16735,N_16162);
nand U23956 (N_23956,N_16853,N_17993);
nor U23957 (N_23957,N_19193,N_16530);
nor U23958 (N_23958,N_15591,N_17111);
or U23959 (N_23959,N_17274,N_15106);
or U23960 (N_23960,N_18737,N_17569);
nand U23961 (N_23961,N_16992,N_15290);
nor U23962 (N_23962,N_16508,N_15447);
nand U23963 (N_23963,N_18958,N_15507);
nand U23964 (N_23964,N_15571,N_18450);
or U23965 (N_23965,N_17723,N_19052);
or U23966 (N_23966,N_16727,N_18924);
and U23967 (N_23967,N_17091,N_17311);
or U23968 (N_23968,N_17796,N_19774);
nor U23969 (N_23969,N_15878,N_17513);
xor U23970 (N_23970,N_17679,N_19750);
nand U23971 (N_23971,N_15697,N_19690);
and U23972 (N_23972,N_18934,N_15266);
or U23973 (N_23973,N_18975,N_19532);
or U23974 (N_23974,N_18870,N_19079);
nand U23975 (N_23975,N_17765,N_17742);
and U23976 (N_23976,N_17367,N_19482);
nor U23977 (N_23977,N_16639,N_17107);
and U23978 (N_23978,N_18846,N_16286);
nand U23979 (N_23979,N_18124,N_16798);
or U23980 (N_23980,N_18904,N_18505);
nand U23981 (N_23981,N_16559,N_16878);
nor U23982 (N_23982,N_17021,N_18568);
or U23983 (N_23983,N_15288,N_17671);
or U23984 (N_23984,N_15292,N_16546);
and U23985 (N_23985,N_15022,N_15693);
and U23986 (N_23986,N_15763,N_15111);
and U23987 (N_23987,N_18446,N_19286);
or U23988 (N_23988,N_19401,N_18006);
or U23989 (N_23989,N_16424,N_15537);
nor U23990 (N_23990,N_18382,N_17350);
or U23991 (N_23991,N_16303,N_15383);
nor U23992 (N_23992,N_15034,N_19159);
or U23993 (N_23993,N_19585,N_16059);
nor U23994 (N_23994,N_16087,N_19492);
and U23995 (N_23995,N_19211,N_15457);
nand U23996 (N_23996,N_18504,N_18282);
nor U23997 (N_23997,N_17895,N_15797);
nand U23998 (N_23998,N_18223,N_18202);
nand U23999 (N_23999,N_19779,N_15364);
nand U24000 (N_24000,N_16931,N_17956);
and U24001 (N_24001,N_19123,N_19978);
nand U24002 (N_24002,N_15825,N_19061);
nor U24003 (N_24003,N_16309,N_19335);
or U24004 (N_24004,N_18505,N_17463);
nor U24005 (N_24005,N_17306,N_15058);
and U24006 (N_24006,N_19594,N_18082);
nor U24007 (N_24007,N_19791,N_17600);
nor U24008 (N_24008,N_16509,N_16109);
and U24009 (N_24009,N_16364,N_17145);
and U24010 (N_24010,N_18451,N_15662);
nor U24011 (N_24011,N_15109,N_19865);
nor U24012 (N_24012,N_16497,N_18100);
nor U24013 (N_24013,N_19108,N_18619);
or U24014 (N_24014,N_18793,N_15572);
nor U24015 (N_24015,N_19846,N_17154);
or U24016 (N_24016,N_16559,N_15711);
and U24017 (N_24017,N_17508,N_15143);
or U24018 (N_24018,N_15199,N_16966);
and U24019 (N_24019,N_16803,N_18277);
and U24020 (N_24020,N_16065,N_16907);
nor U24021 (N_24021,N_16371,N_16833);
or U24022 (N_24022,N_15103,N_18797);
or U24023 (N_24023,N_18922,N_18075);
or U24024 (N_24024,N_15401,N_17762);
nor U24025 (N_24025,N_18807,N_17125);
nand U24026 (N_24026,N_17307,N_17844);
and U24027 (N_24027,N_18152,N_15474);
nor U24028 (N_24028,N_16755,N_15447);
and U24029 (N_24029,N_19972,N_18574);
and U24030 (N_24030,N_16053,N_15566);
nor U24031 (N_24031,N_15558,N_15772);
nor U24032 (N_24032,N_19738,N_18561);
nand U24033 (N_24033,N_19239,N_18734);
nor U24034 (N_24034,N_18475,N_15062);
and U24035 (N_24035,N_17036,N_16852);
and U24036 (N_24036,N_16598,N_16001);
nor U24037 (N_24037,N_17468,N_16769);
or U24038 (N_24038,N_17654,N_18559);
or U24039 (N_24039,N_18921,N_17401);
or U24040 (N_24040,N_19093,N_16897);
nand U24041 (N_24041,N_18843,N_17351);
and U24042 (N_24042,N_17371,N_19166);
nand U24043 (N_24043,N_15940,N_19508);
and U24044 (N_24044,N_17619,N_15879);
nor U24045 (N_24045,N_16425,N_15327);
and U24046 (N_24046,N_18709,N_17132);
or U24047 (N_24047,N_16134,N_18682);
or U24048 (N_24048,N_16398,N_17265);
nor U24049 (N_24049,N_15135,N_17473);
nor U24050 (N_24050,N_19680,N_17599);
xor U24051 (N_24051,N_15013,N_18566);
and U24052 (N_24052,N_17730,N_18565);
and U24053 (N_24053,N_16541,N_15713);
nand U24054 (N_24054,N_15300,N_19810);
and U24055 (N_24055,N_18854,N_17689);
nand U24056 (N_24056,N_18904,N_18305);
nor U24057 (N_24057,N_16592,N_19372);
xor U24058 (N_24058,N_19277,N_19538);
nor U24059 (N_24059,N_17330,N_15810);
or U24060 (N_24060,N_17439,N_16923);
nor U24061 (N_24061,N_17783,N_17994);
nand U24062 (N_24062,N_18270,N_15448);
nor U24063 (N_24063,N_17651,N_15355);
nand U24064 (N_24064,N_16225,N_15538);
or U24065 (N_24065,N_15468,N_15180);
or U24066 (N_24066,N_16347,N_16838);
nand U24067 (N_24067,N_15043,N_17427);
nor U24068 (N_24068,N_16385,N_15190);
xor U24069 (N_24069,N_16306,N_15366);
or U24070 (N_24070,N_19788,N_18230);
and U24071 (N_24071,N_15514,N_16647);
or U24072 (N_24072,N_16821,N_17600);
and U24073 (N_24073,N_19194,N_19186);
and U24074 (N_24074,N_16767,N_16143);
or U24075 (N_24075,N_19651,N_16784);
and U24076 (N_24076,N_15257,N_17374);
nor U24077 (N_24077,N_18891,N_19471);
nor U24078 (N_24078,N_17711,N_18250);
and U24079 (N_24079,N_17545,N_18890);
and U24080 (N_24080,N_17473,N_15579);
and U24081 (N_24081,N_15340,N_19435);
nand U24082 (N_24082,N_17088,N_15880);
nor U24083 (N_24083,N_16439,N_15382);
or U24084 (N_24084,N_17798,N_19879);
nand U24085 (N_24085,N_17483,N_15506);
nor U24086 (N_24086,N_19407,N_18273);
xor U24087 (N_24087,N_19678,N_19412);
nor U24088 (N_24088,N_18515,N_17457);
and U24089 (N_24089,N_16557,N_19485);
and U24090 (N_24090,N_17032,N_15311);
or U24091 (N_24091,N_15695,N_18826);
or U24092 (N_24092,N_18632,N_19211);
and U24093 (N_24093,N_19148,N_19290);
nand U24094 (N_24094,N_19908,N_17674);
nand U24095 (N_24095,N_18024,N_19841);
or U24096 (N_24096,N_18949,N_18328);
and U24097 (N_24097,N_15352,N_16546);
and U24098 (N_24098,N_18642,N_15936);
and U24099 (N_24099,N_17267,N_17077);
or U24100 (N_24100,N_17893,N_16918);
and U24101 (N_24101,N_19675,N_16693);
or U24102 (N_24102,N_17801,N_17590);
or U24103 (N_24103,N_16052,N_17956);
and U24104 (N_24104,N_17675,N_18314);
and U24105 (N_24105,N_19929,N_15866);
or U24106 (N_24106,N_17582,N_17229);
nand U24107 (N_24107,N_15580,N_17722);
nand U24108 (N_24108,N_18022,N_15798);
or U24109 (N_24109,N_19148,N_17763);
nand U24110 (N_24110,N_16624,N_18698);
or U24111 (N_24111,N_16001,N_16082);
nand U24112 (N_24112,N_19178,N_15435);
nand U24113 (N_24113,N_16241,N_18489);
nand U24114 (N_24114,N_16794,N_18444);
nor U24115 (N_24115,N_15373,N_17200);
and U24116 (N_24116,N_19607,N_16527);
nand U24117 (N_24117,N_18963,N_18510);
nand U24118 (N_24118,N_17634,N_15428);
or U24119 (N_24119,N_19754,N_15110);
and U24120 (N_24120,N_18466,N_18616);
nor U24121 (N_24121,N_16157,N_18200);
xor U24122 (N_24122,N_17476,N_18611);
and U24123 (N_24123,N_17815,N_19455);
nor U24124 (N_24124,N_17605,N_18688);
nand U24125 (N_24125,N_16729,N_17004);
nor U24126 (N_24126,N_18359,N_16706);
nand U24127 (N_24127,N_19883,N_17356);
nor U24128 (N_24128,N_17553,N_18582);
nand U24129 (N_24129,N_15596,N_17101);
nand U24130 (N_24130,N_15309,N_15009);
and U24131 (N_24131,N_18580,N_19471);
or U24132 (N_24132,N_16724,N_19493);
and U24133 (N_24133,N_17407,N_15677);
nand U24134 (N_24134,N_19181,N_17972);
nor U24135 (N_24135,N_18261,N_16627);
or U24136 (N_24136,N_17100,N_15229);
and U24137 (N_24137,N_16317,N_19059);
and U24138 (N_24138,N_15028,N_18158);
nor U24139 (N_24139,N_19073,N_15427);
and U24140 (N_24140,N_16185,N_19382);
and U24141 (N_24141,N_17413,N_19244);
nor U24142 (N_24142,N_19519,N_17630);
nor U24143 (N_24143,N_18043,N_16363);
and U24144 (N_24144,N_18275,N_15415);
and U24145 (N_24145,N_16323,N_15234);
and U24146 (N_24146,N_19301,N_15017);
nor U24147 (N_24147,N_17477,N_16206);
nand U24148 (N_24148,N_19763,N_15555);
and U24149 (N_24149,N_17244,N_15970);
and U24150 (N_24150,N_17293,N_18561);
and U24151 (N_24151,N_16979,N_15875);
nor U24152 (N_24152,N_17311,N_15398);
or U24153 (N_24153,N_16941,N_16358);
nand U24154 (N_24154,N_18402,N_17227);
or U24155 (N_24155,N_17108,N_15280);
and U24156 (N_24156,N_17849,N_18321);
and U24157 (N_24157,N_19275,N_15787);
nand U24158 (N_24158,N_16750,N_18594);
and U24159 (N_24159,N_19717,N_18304);
nor U24160 (N_24160,N_18485,N_17831);
nor U24161 (N_24161,N_17417,N_18222);
nand U24162 (N_24162,N_17819,N_17765);
and U24163 (N_24163,N_19657,N_17506);
and U24164 (N_24164,N_19901,N_18929);
nor U24165 (N_24165,N_18316,N_15391);
nand U24166 (N_24166,N_16718,N_15073);
nor U24167 (N_24167,N_17029,N_15170);
nand U24168 (N_24168,N_16809,N_19460);
nor U24169 (N_24169,N_15923,N_19810);
nand U24170 (N_24170,N_15825,N_18152);
nor U24171 (N_24171,N_18771,N_15282);
xor U24172 (N_24172,N_16822,N_15108);
nand U24173 (N_24173,N_15162,N_18936);
nand U24174 (N_24174,N_18075,N_15037);
nand U24175 (N_24175,N_17542,N_15850);
nor U24176 (N_24176,N_16335,N_18241);
nand U24177 (N_24177,N_19156,N_16004);
nand U24178 (N_24178,N_19405,N_18832);
and U24179 (N_24179,N_17433,N_18441);
nor U24180 (N_24180,N_15397,N_17134);
xor U24181 (N_24181,N_18852,N_17679);
nor U24182 (N_24182,N_16653,N_19261);
nand U24183 (N_24183,N_15701,N_16720);
xnor U24184 (N_24184,N_17435,N_18123);
and U24185 (N_24185,N_15808,N_15663);
or U24186 (N_24186,N_16735,N_18151);
and U24187 (N_24187,N_16028,N_15796);
or U24188 (N_24188,N_18454,N_17997);
or U24189 (N_24189,N_16331,N_17158);
or U24190 (N_24190,N_17138,N_16670);
or U24191 (N_24191,N_16774,N_18007);
and U24192 (N_24192,N_19901,N_18611);
and U24193 (N_24193,N_15221,N_17730);
or U24194 (N_24194,N_18891,N_16450);
or U24195 (N_24195,N_15965,N_16586);
nor U24196 (N_24196,N_17196,N_16184);
or U24197 (N_24197,N_18735,N_17680);
nor U24198 (N_24198,N_16835,N_18266);
nor U24199 (N_24199,N_15962,N_19162);
and U24200 (N_24200,N_16818,N_17578);
and U24201 (N_24201,N_16871,N_16978);
xor U24202 (N_24202,N_15899,N_18763);
and U24203 (N_24203,N_15615,N_17750);
and U24204 (N_24204,N_15404,N_17307);
or U24205 (N_24205,N_15530,N_16460);
nor U24206 (N_24206,N_18564,N_17956);
nand U24207 (N_24207,N_16580,N_15205);
or U24208 (N_24208,N_17799,N_18970);
nor U24209 (N_24209,N_19808,N_17411);
nand U24210 (N_24210,N_16643,N_18415);
or U24211 (N_24211,N_19987,N_19351);
nand U24212 (N_24212,N_15996,N_16475);
nand U24213 (N_24213,N_19964,N_17267);
nand U24214 (N_24214,N_15069,N_16079);
xor U24215 (N_24215,N_18117,N_19993);
nand U24216 (N_24216,N_15219,N_16341);
and U24217 (N_24217,N_17384,N_15404);
or U24218 (N_24218,N_15685,N_16251);
nor U24219 (N_24219,N_16645,N_15172);
or U24220 (N_24220,N_19597,N_17381);
nand U24221 (N_24221,N_18767,N_15073);
and U24222 (N_24222,N_15593,N_16537);
and U24223 (N_24223,N_17797,N_17354);
nand U24224 (N_24224,N_19880,N_19253);
and U24225 (N_24225,N_15835,N_15049);
nand U24226 (N_24226,N_18707,N_18176);
nor U24227 (N_24227,N_18294,N_16264);
nor U24228 (N_24228,N_19998,N_15937);
or U24229 (N_24229,N_17753,N_17947);
or U24230 (N_24230,N_16361,N_19888);
or U24231 (N_24231,N_17554,N_19943);
and U24232 (N_24232,N_18619,N_17574);
and U24233 (N_24233,N_16046,N_15670);
nand U24234 (N_24234,N_15638,N_16308);
nor U24235 (N_24235,N_18023,N_17124);
xor U24236 (N_24236,N_15005,N_17810);
xor U24237 (N_24237,N_15982,N_17398);
nor U24238 (N_24238,N_18121,N_18054);
nor U24239 (N_24239,N_16174,N_17094);
and U24240 (N_24240,N_18293,N_17442);
and U24241 (N_24241,N_17970,N_17020);
nor U24242 (N_24242,N_17214,N_19281);
or U24243 (N_24243,N_15697,N_16014);
nor U24244 (N_24244,N_15104,N_16419);
nor U24245 (N_24245,N_17814,N_15220);
nor U24246 (N_24246,N_15494,N_19243);
or U24247 (N_24247,N_18294,N_17964);
and U24248 (N_24248,N_18125,N_16626);
nand U24249 (N_24249,N_18646,N_19278);
or U24250 (N_24250,N_15410,N_19509);
nand U24251 (N_24251,N_16114,N_19369);
or U24252 (N_24252,N_17260,N_15336);
xor U24253 (N_24253,N_15239,N_15166);
nor U24254 (N_24254,N_15295,N_19911);
or U24255 (N_24255,N_16393,N_18449);
nor U24256 (N_24256,N_16838,N_16092);
nor U24257 (N_24257,N_19794,N_15011);
and U24258 (N_24258,N_18527,N_18540);
and U24259 (N_24259,N_15648,N_16405);
or U24260 (N_24260,N_17226,N_18136);
nor U24261 (N_24261,N_18783,N_19622);
and U24262 (N_24262,N_17919,N_15230);
and U24263 (N_24263,N_19308,N_16353);
nor U24264 (N_24264,N_17471,N_16119);
nor U24265 (N_24265,N_15019,N_18698);
and U24266 (N_24266,N_18534,N_15393);
nor U24267 (N_24267,N_18788,N_16486);
and U24268 (N_24268,N_18519,N_15832);
nor U24269 (N_24269,N_16849,N_17058);
nor U24270 (N_24270,N_19805,N_16565);
or U24271 (N_24271,N_16766,N_16228);
xnor U24272 (N_24272,N_16815,N_16772);
xor U24273 (N_24273,N_16603,N_19660);
nand U24274 (N_24274,N_19108,N_17982);
nand U24275 (N_24275,N_19034,N_19610);
nand U24276 (N_24276,N_17258,N_19887);
nand U24277 (N_24277,N_19334,N_15086);
nand U24278 (N_24278,N_15494,N_19654);
and U24279 (N_24279,N_17299,N_15584);
and U24280 (N_24280,N_17278,N_15911);
nand U24281 (N_24281,N_17974,N_17723);
or U24282 (N_24282,N_16379,N_15033);
nor U24283 (N_24283,N_19568,N_18153);
nor U24284 (N_24284,N_19142,N_17795);
or U24285 (N_24285,N_17944,N_16211);
or U24286 (N_24286,N_18395,N_17572);
nand U24287 (N_24287,N_16199,N_16542);
or U24288 (N_24288,N_17093,N_17753);
and U24289 (N_24289,N_19358,N_18664);
nor U24290 (N_24290,N_16428,N_19801);
and U24291 (N_24291,N_19140,N_19721);
nor U24292 (N_24292,N_15489,N_16133);
nor U24293 (N_24293,N_17780,N_18000);
or U24294 (N_24294,N_16690,N_16030);
nor U24295 (N_24295,N_19702,N_16118);
or U24296 (N_24296,N_16848,N_17006);
nand U24297 (N_24297,N_15771,N_18436);
nand U24298 (N_24298,N_15142,N_16535);
nor U24299 (N_24299,N_17943,N_19289);
nor U24300 (N_24300,N_16391,N_16056);
or U24301 (N_24301,N_18321,N_19812);
or U24302 (N_24302,N_17370,N_15500);
nand U24303 (N_24303,N_15595,N_15343);
and U24304 (N_24304,N_16148,N_17089);
or U24305 (N_24305,N_19340,N_15269);
and U24306 (N_24306,N_18178,N_18699);
nand U24307 (N_24307,N_18302,N_15087);
nor U24308 (N_24308,N_17358,N_17377);
nand U24309 (N_24309,N_15912,N_18462);
nor U24310 (N_24310,N_17810,N_15361);
or U24311 (N_24311,N_17806,N_15078);
or U24312 (N_24312,N_17044,N_18452);
nor U24313 (N_24313,N_15209,N_15708);
or U24314 (N_24314,N_17115,N_16271);
nand U24315 (N_24315,N_17976,N_17924);
nand U24316 (N_24316,N_16305,N_16656);
nand U24317 (N_24317,N_19623,N_19776);
or U24318 (N_24318,N_16513,N_17242);
and U24319 (N_24319,N_18026,N_15372);
nand U24320 (N_24320,N_16278,N_16753);
xnor U24321 (N_24321,N_16454,N_19659);
xnor U24322 (N_24322,N_18245,N_16957);
nand U24323 (N_24323,N_19394,N_15720);
and U24324 (N_24324,N_17105,N_19280);
nor U24325 (N_24325,N_19964,N_16930);
nor U24326 (N_24326,N_17324,N_17623);
nand U24327 (N_24327,N_17192,N_16483);
nor U24328 (N_24328,N_16743,N_16735);
nand U24329 (N_24329,N_18639,N_18842);
and U24330 (N_24330,N_18315,N_17616);
nor U24331 (N_24331,N_17499,N_19314);
or U24332 (N_24332,N_16894,N_16292);
or U24333 (N_24333,N_15447,N_15762);
nor U24334 (N_24334,N_18167,N_18705);
nand U24335 (N_24335,N_15024,N_15935);
nor U24336 (N_24336,N_15966,N_19620);
or U24337 (N_24337,N_19594,N_15235);
nand U24338 (N_24338,N_19418,N_15453);
nor U24339 (N_24339,N_18058,N_15241);
and U24340 (N_24340,N_16006,N_15863);
and U24341 (N_24341,N_15502,N_19503);
nor U24342 (N_24342,N_15863,N_16966);
and U24343 (N_24343,N_15933,N_18857);
nor U24344 (N_24344,N_16028,N_17767);
or U24345 (N_24345,N_16363,N_15489);
nand U24346 (N_24346,N_16203,N_18560);
and U24347 (N_24347,N_16281,N_18596);
and U24348 (N_24348,N_16660,N_18114);
nor U24349 (N_24349,N_18025,N_15221);
nand U24350 (N_24350,N_16227,N_17900);
nand U24351 (N_24351,N_17062,N_15782);
xnor U24352 (N_24352,N_17425,N_17740);
nand U24353 (N_24353,N_15376,N_19805);
or U24354 (N_24354,N_19214,N_15276);
nand U24355 (N_24355,N_15883,N_19389);
or U24356 (N_24356,N_16629,N_18735);
or U24357 (N_24357,N_17676,N_15785);
or U24358 (N_24358,N_18176,N_16926);
nor U24359 (N_24359,N_19496,N_17174);
and U24360 (N_24360,N_16690,N_19868);
and U24361 (N_24361,N_19743,N_15140);
xor U24362 (N_24362,N_16304,N_15622);
and U24363 (N_24363,N_19171,N_17191);
nand U24364 (N_24364,N_16836,N_16635);
or U24365 (N_24365,N_16150,N_15992);
or U24366 (N_24366,N_15957,N_19009);
nor U24367 (N_24367,N_16826,N_16428);
or U24368 (N_24368,N_18295,N_17786);
or U24369 (N_24369,N_18872,N_17425);
and U24370 (N_24370,N_18186,N_16532);
nor U24371 (N_24371,N_18600,N_17145);
nor U24372 (N_24372,N_19336,N_18392);
nand U24373 (N_24373,N_16078,N_16270);
and U24374 (N_24374,N_16514,N_18256);
nand U24375 (N_24375,N_17089,N_16585);
and U24376 (N_24376,N_17294,N_16793);
and U24377 (N_24377,N_18230,N_16270);
nand U24378 (N_24378,N_19707,N_19530);
nor U24379 (N_24379,N_18557,N_16257);
or U24380 (N_24380,N_19768,N_17563);
or U24381 (N_24381,N_18679,N_18754);
and U24382 (N_24382,N_19668,N_18029);
nor U24383 (N_24383,N_15646,N_16474);
or U24384 (N_24384,N_19538,N_16113);
and U24385 (N_24385,N_19987,N_17909);
nand U24386 (N_24386,N_18809,N_17079);
or U24387 (N_24387,N_19649,N_16797);
and U24388 (N_24388,N_16832,N_16514);
nor U24389 (N_24389,N_18351,N_18747);
or U24390 (N_24390,N_16969,N_15167);
or U24391 (N_24391,N_18514,N_15498);
nor U24392 (N_24392,N_16441,N_16558);
xnor U24393 (N_24393,N_17144,N_19284);
or U24394 (N_24394,N_16935,N_18086);
or U24395 (N_24395,N_17532,N_17895);
nand U24396 (N_24396,N_19182,N_15538);
xnor U24397 (N_24397,N_16186,N_15309);
nor U24398 (N_24398,N_16646,N_19961);
and U24399 (N_24399,N_15492,N_16344);
nor U24400 (N_24400,N_18421,N_15954);
and U24401 (N_24401,N_15776,N_15265);
nand U24402 (N_24402,N_17619,N_15027);
nor U24403 (N_24403,N_15147,N_15064);
and U24404 (N_24404,N_18741,N_15276);
nand U24405 (N_24405,N_19120,N_19226);
and U24406 (N_24406,N_16667,N_16997);
and U24407 (N_24407,N_17733,N_19106);
or U24408 (N_24408,N_15015,N_16512);
nand U24409 (N_24409,N_17426,N_19916);
nor U24410 (N_24410,N_16272,N_19925);
nor U24411 (N_24411,N_19158,N_15986);
nor U24412 (N_24412,N_16416,N_19647);
or U24413 (N_24413,N_16532,N_18756);
nor U24414 (N_24414,N_17751,N_18047);
or U24415 (N_24415,N_17739,N_15403);
or U24416 (N_24416,N_16051,N_18290);
nand U24417 (N_24417,N_18952,N_15634);
xor U24418 (N_24418,N_17054,N_16005);
xnor U24419 (N_24419,N_15929,N_19632);
or U24420 (N_24420,N_16883,N_17193);
or U24421 (N_24421,N_19299,N_16949);
nor U24422 (N_24422,N_19012,N_17216);
and U24423 (N_24423,N_16221,N_18566);
xor U24424 (N_24424,N_19642,N_18185);
and U24425 (N_24425,N_19846,N_19594);
and U24426 (N_24426,N_18954,N_16852);
or U24427 (N_24427,N_16984,N_18436);
nor U24428 (N_24428,N_17676,N_15801);
or U24429 (N_24429,N_19026,N_16557);
nor U24430 (N_24430,N_16122,N_17371);
nor U24431 (N_24431,N_15051,N_16332);
nor U24432 (N_24432,N_15366,N_16765);
nand U24433 (N_24433,N_19229,N_16645);
xnor U24434 (N_24434,N_15432,N_16040);
and U24435 (N_24435,N_18541,N_19042);
or U24436 (N_24436,N_18910,N_18750);
or U24437 (N_24437,N_15992,N_15642);
and U24438 (N_24438,N_19987,N_18392);
and U24439 (N_24439,N_19022,N_15543);
or U24440 (N_24440,N_18958,N_19020);
nand U24441 (N_24441,N_19379,N_19851);
nor U24442 (N_24442,N_15272,N_17158);
and U24443 (N_24443,N_15461,N_19467);
nor U24444 (N_24444,N_18565,N_17189);
or U24445 (N_24445,N_18276,N_17415);
nor U24446 (N_24446,N_19451,N_17081);
nand U24447 (N_24447,N_18423,N_18649);
and U24448 (N_24448,N_18183,N_15642);
or U24449 (N_24449,N_18289,N_16391);
nand U24450 (N_24450,N_15952,N_17197);
and U24451 (N_24451,N_19807,N_18326);
and U24452 (N_24452,N_16833,N_18856);
and U24453 (N_24453,N_16380,N_16694);
and U24454 (N_24454,N_18264,N_19502);
and U24455 (N_24455,N_15210,N_15232);
nor U24456 (N_24456,N_19279,N_17956);
nor U24457 (N_24457,N_17209,N_15575);
nor U24458 (N_24458,N_16783,N_16527);
nor U24459 (N_24459,N_15854,N_18771);
and U24460 (N_24460,N_16380,N_15563);
or U24461 (N_24461,N_18244,N_18582);
xnor U24462 (N_24462,N_17099,N_17593);
and U24463 (N_24463,N_18132,N_18255);
nand U24464 (N_24464,N_15647,N_15567);
nand U24465 (N_24465,N_19359,N_18438);
and U24466 (N_24466,N_18811,N_19878);
or U24467 (N_24467,N_16207,N_19212);
or U24468 (N_24468,N_19047,N_19756);
nand U24469 (N_24469,N_16384,N_17446);
and U24470 (N_24470,N_18068,N_15272);
nor U24471 (N_24471,N_17344,N_19716);
or U24472 (N_24472,N_18186,N_19560);
nand U24473 (N_24473,N_15041,N_17255);
nor U24474 (N_24474,N_16226,N_19800);
nor U24475 (N_24475,N_18141,N_18284);
nor U24476 (N_24476,N_19470,N_18438);
nor U24477 (N_24477,N_19692,N_19634);
or U24478 (N_24478,N_19986,N_15617);
and U24479 (N_24479,N_17264,N_18154);
or U24480 (N_24480,N_16009,N_18703);
nand U24481 (N_24481,N_18162,N_19684);
nand U24482 (N_24482,N_18395,N_15209);
or U24483 (N_24483,N_16688,N_16720);
nor U24484 (N_24484,N_19987,N_17593);
nand U24485 (N_24485,N_19679,N_19738);
nor U24486 (N_24486,N_17872,N_15603);
and U24487 (N_24487,N_17280,N_19516);
or U24488 (N_24488,N_18937,N_16146);
or U24489 (N_24489,N_18890,N_16764);
nor U24490 (N_24490,N_15248,N_15655);
nor U24491 (N_24491,N_16039,N_17866);
xnor U24492 (N_24492,N_16639,N_17925);
nor U24493 (N_24493,N_18713,N_18138);
and U24494 (N_24494,N_16556,N_15392);
or U24495 (N_24495,N_17962,N_18327);
or U24496 (N_24496,N_16879,N_15829);
nand U24497 (N_24497,N_16108,N_17677);
nand U24498 (N_24498,N_15265,N_15083);
or U24499 (N_24499,N_15720,N_17116);
or U24500 (N_24500,N_15039,N_18492);
nor U24501 (N_24501,N_18698,N_16829);
nand U24502 (N_24502,N_18064,N_15273);
or U24503 (N_24503,N_19409,N_15580);
or U24504 (N_24504,N_16832,N_18406);
and U24505 (N_24505,N_17555,N_17975);
or U24506 (N_24506,N_18405,N_15715);
nor U24507 (N_24507,N_16950,N_16311);
nand U24508 (N_24508,N_19249,N_18507);
xnor U24509 (N_24509,N_18742,N_16001);
or U24510 (N_24510,N_18431,N_19492);
or U24511 (N_24511,N_15846,N_15420);
nor U24512 (N_24512,N_19883,N_18779);
nor U24513 (N_24513,N_15927,N_16873);
and U24514 (N_24514,N_15552,N_18638);
or U24515 (N_24515,N_18179,N_17179);
nand U24516 (N_24516,N_19627,N_18526);
or U24517 (N_24517,N_19058,N_18865);
or U24518 (N_24518,N_19290,N_16703);
nor U24519 (N_24519,N_17988,N_17048);
nor U24520 (N_24520,N_16183,N_17732);
and U24521 (N_24521,N_15762,N_16611);
or U24522 (N_24522,N_18178,N_18101);
xor U24523 (N_24523,N_18907,N_19245);
and U24524 (N_24524,N_16073,N_19964);
nor U24525 (N_24525,N_15215,N_19295);
nor U24526 (N_24526,N_17892,N_15570);
nor U24527 (N_24527,N_17893,N_18770);
nand U24528 (N_24528,N_16111,N_15516);
and U24529 (N_24529,N_18218,N_15698);
or U24530 (N_24530,N_18440,N_17896);
or U24531 (N_24531,N_17185,N_19725);
or U24532 (N_24532,N_18437,N_19963);
and U24533 (N_24533,N_15448,N_19864);
nor U24534 (N_24534,N_16107,N_16920);
nor U24535 (N_24535,N_18613,N_19727);
or U24536 (N_24536,N_18337,N_17477);
nand U24537 (N_24537,N_18081,N_15244);
xnor U24538 (N_24538,N_16638,N_16302);
or U24539 (N_24539,N_18938,N_16841);
nor U24540 (N_24540,N_18236,N_19629);
or U24541 (N_24541,N_19453,N_16909);
nand U24542 (N_24542,N_16262,N_17948);
or U24543 (N_24543,N_19154,N_15484);
nand U24544 (N_24544,N_18391,N_18494);
or U24545 (N_24545,N_17915,N_16618);
nor U24546 (N_24546,N_15777,N_18622);
nand U24547 (N_24547,N_19799,N_15110);
nor U24548 (N_24548,N_19001,N_18530);
and U24549 (N_24549,N_15327,N_15017);
nand U24550 (N_24550,N_19077,N_15472);
or U24551 (N_24551,N_15818,N_15117);
and U24552 (N_24552,N_19103,N_19427);
and U24553 (N_24553,N_19520,N_17395);
xor U24554 (N_24554,N_15105,N_16643);
nor U24555 (N_24555,N_18709,N_16590);
nor U24556 (N_24556,N_18396,N_18453);
nor U24557 (N_24557,N_16941,N_15147);
nand U24558 (N_24558,N_15266,N_17941);
nand U24559 (N_24559,N_17318,N_15754);
and U24560 (N_24560,N_17490,N_16892);
nand U24561 (N_24561,N_15140,N_15357);
nor U24562 (N_24562,N_16868,N_17750);
or U24563 (N_24563,N_19173,N_18859);
nand U24564 (N_24564,N_18117,N_16410);
nand U24565 (N_24565,N_15927,N_19382);
nand U24566 (N_24566,N_19588,N_18277);
nand U24567 (N_24567,N_16725,N_15887);
nand U24568 (N_24568,N_16097,N_17120);
nor U24569 (N_24569,N_16913,N_16131);
nor U24570 (N_24570,N_19052,N_16088);
and U24571 (N_24571,N_16631,N_19469);
nor U24572 (N_24572,N_18452,N_15042);
and U24573 (N_24573,N_17055,N_16589);
nand U24574 (N_24574,N_19557,N_19469);
or U24575 (N_24575,N_19334,N_16120);
nand U24576 (N_24576,N_19278,N_15572);
and U24577 (N_24577,N_17834,N_16424);
nand U24578 (N_24578,N_17587,N_17317);
and U24579 (N_24579,N_16076,N_17528);
or U24580 (N_24580,N_19010,N_18007);
nor U24581 (N_24581,N_16691,N_18524);
and U24582 (N_24582,N_19042,N_18695);
nand U24583 (N_24583,N_17529,N_18646);
and U24584 (N_24584,N_16786,N_18035);
nor U24585 (N_24585,N_17578,N_16897);
nand U24586 (N_24586,N_17876,N_17895);
nand U24587 (N_24587,N_19784,N_17105);
and U24588 (N_24588,N_17648,N_17333);
or U24589 (N_24589,N_19322,N_18697);
nand U24590 (N_24590,N_15186,N_19625);
or U24591 (N_24591,N_18529,N_18802);
and U24592 (N_24592,N_15677,N_19721);
or U24593 (N_24593,N_19589,N_18520);
and U24594 (N_24594,N_15689,N_16335);
nor U24595 (N_24595,N_15668,N_16680);
and U24596 (N_24596,N_15315,N_16067);
or U24597 (N_24597,N_15959,N_18432);
nand U24598 (N_24598,N_15005,N_16610);
nor U24599 (N_24599,N_18003,N_18125);
nand U24600 (N_24600,N_16455,N_15768);
and U24601 (N_24601,N_19070,N_17846);
or U24602 (N_24602,N_15198,N_17231);
and U24603 (N_24603,N_15055,N_15514);
or U24604 (N_24604,N_18538,N_16971);
and U24605 (N_24605,N_15101,N_19898);
or U24606 (N_24606,N_19995,N_15619);
nand U24607 (N_24607,N_15792,N_19489);
nand U24608 (N_24608,N_18543,N_15914);
or U24609 (N_24609,N_15954,N_16880);
or U24610 (N_24610,N_16798,N_17512);
or U24611 (N_24611,N_16617,N_17780);
or U24612 (N_24612,N_15463,N_18051);
nand U24613 (N_24613,N_17526,N_17826);
nand U24614 (N_24614,N_16524,N_15572);
or U24615 (N_24615,N_17759,N_15769);
nand U24616 (N_24616,N_15488,N_16750);
nand U24617 (N_24617,N_15464,N_17356);
and U24618 (N_24618,N_17464,N_18110);
nor U24619 (N_24619,N_19595,N_19519);
or U24620 (N_24620,N_15668,N_17731);
nor U24621 (N_24621,N_16361,N_18619);
and U24622 (N_24622,N_17424,N_19116);
nor U24623 (N_24623,N_18838,N_15930);
nor U24624 (N_24624,N_15534,N_15624);
or U24625 (N_24625,N_18468,N_16274);
nand U24626 (N_24626,N_18498,N_18242);
or U24627 (N_24627,N_15781,N_16015);
or U24628 (N_24628,N_18454,N_17650);
or U24629 (N_24629,N_15133,N_15237);
xnor U24630 (N_24630,N_17533,N_18102);
nand U24631 (N_24631,N_18722,N_15862);
nor U24632 (N_24632,N_15865,N_19368);
and U24633 (N_24633,N_19207,N_19277);
nor U24634 (N_24634,N_15219,N_18928);
or U24635 (N_24635,N_19190,N_18767);
nor U24636 (N_24636,N_19961,N_18788);
and U24637 (N_24637,N_15361,N_18415);
nor U24638 (N_24638,N_17196,N_19422);
nand U24639 (N_24639,N_16773,N_16858);
and U24640 (N_24640,N_19635,N_16536);
nand U24641 (N_24641,N_15690,N_15597);
xor U24642 (N_24642,N_17216,N_17068);
or U24643 (N_24643,N_16754,N_19811);
and U24644 (N_24644,N_16447,N_19939);
xnor U24645 (N_24645,N_15075,N_19877);
and U24646 (N_24646,N_15443,N_15902);
nor U24647 (N_24647,N_16645,N_17006);
and U24648 (N_24648,N_15139,N_18066);
nor U24649 (N_24649,N_17339,N_16607);
and U24650 (N_24650,N_15994,N_17988);
nand U24651 (N_24651,N_18463,N_16831);
nand U24652 (N_24652,N_15111,N_16625);
xnor U24653 (N_24653,N_19089,N_17824);
nand U24654 (N_24654,N_19830,N_19234);
and U24655 (N_24655,N_17376,N_16966);
nand U24656 (N_24656,N_17209,N_15425);
nand U24657 (N_24657,N_15804,N_19109);
nor U24658 (N_24658,N_17017,N_19092);
and U24659 (N_24659,N_19441,N_18180);
and U24660 (N_24660,N_16360,N_19031);
nor U24661 (N_24661,N_17307,N_15418);
and U24662 (N_24662,N_19979,N_17884);
nor U24663 (N_24663,N_19372,N_15333);
and U24664 (N_24664,N_18942,N_17466);
and U24665 (N_24665,N_17125,N_15803);
nor U24666 (N_24666,N_17625,N_15561);
and U24667 (N_24667,N_17111,N_17647);
or U24668 (N_24668,N_16477,N_15872);
or U24669 (N_24669,N_16104,N_19931);
nor U24670 (N_24670,N_18739,N_16400);
nand U24671 (N_24671,N_17311,N_16495);
and U24672 (N_24672,N_19858,N_19140);
and U24673 (N_24673,N_18820,N_16455);
nand U24674 (N_24674,N_17499,N_15388);
nor U24675 (N_24675,N_16836,N_17967);
nor U24676 (N_24676,N_17091,N_16813);
or U24677 (N_24677,N_18511,N_17020);
or U24678 (N_24678,N_17750,N_17345);
nand U24679 (N_24679,N_16680,N_16088);
or U24680 (N_24680,N_18969,N_19855);
and U24681 (N_24681,N_18275,N_16306);
nand U24682 (N_24682,N_18695,N_18732);
and U24683 (N_24683,N_17360,N_17140);
nand U24684 (N_24684,N_18201,N_19969);
or U24685 (N_24685,N_17619,N_16976);
or U24686 (N_24686,N_19342,N_16659);
nand U24687 (N_24687,N_18187,N_19864);
nand U24688 (N_24688,N_15823,N_18097);
nand U24689 (N_24689,N_16937,N_15644);
nand U24690 (N_24690,N_19354,N_15879);
or U24691 (N_24691,N_15029,N_17002);
nand U24692 (N_24692,N_15523,N_18843);
and U24693 (N_24693,N_18566,N_15805);
nor U24694 (N_24694,N_18809,N_18481);
nor U24695 (N_24695,N_19238,N_15141);
xnor U24696 (N_24696,N_19009,N_17960);
nor U24697 (N_24697,N_15160,N_17462);
nand U24698 (N_24698,N_19217,N_16581);
nor U24699 (N_24699,N_17804,N_19834);
nor U24700 (N_24700,N_17693,N_18770);
nor U24701 (N_24701,N_15512,N_15132);
nor U24702 (N_24702,N_16662,N_17962);
nand U24703 (N_24703,N_17307,N_15111);
or U24704 (N_24704,N_15963,N_15625);
and U24705 (N_24705,N_19712,N_15750);
or U24706 (N_24706,N_15104,N_17827);
nand U24707 (N_24707,N_16668,N_17108);
or U24708 (N_24708,N_15496,N_18434);
and U24709 (N_24709,N_17293,N_19650);
nor U24710 (N_24710,N_18746,N_19060);
nor U24711 (N_24711,N_17868,N_15751);
nand U24712 (N_24712,N_15625,N_19719);
or U24713 (N_24713,N_17032,N_19777);
or U24714 (N_24714,N_18807,N_18011);
and U24715 (N_24715,N_17529,N_18361);
or U24716 (N_24716,N_19038,N_16863);
nor U24717 (N_24717,N_15265,N_17435);
or U24718 (N_24718,N_16417,N_16646);
or U24719 (N_24719,N_17879,N_15246);
nor U24720 (N_24720,N_19707,N_19507);
or U24721 (N_24721,N_19220,N_16301);
and U24722 (N_24722,N_18101,N_16492);
or U24723 (N_24723,N_19312,N_19385);
and U24724 (N_24724,N_17637,N_17665);
nor U24725 (N_24725,N_18373,N_16826);
nor U24726 (N_24726,N_18170,N_15190);
or U24727 (N_24727,N_15272,N_19965);
or U24728 (N_24728,N_19447,N_17887);
nand U24729 (N_24729,N_18578,N_18417);
nor U24730 (N_24730,N_19740,N_15198);
nand U24731 (N_24731,N_16878,N_19454);
nor U24732 (N_24732,N_18028,N_15445);
and U24733 (N_24733,N_16945,N_19314);
nand U24734 (N_24734,N_18428,N_16033);
nand U24735 (N_24735,N_16681,N_16551);
and U24736 (N_24736,N_19657,N_17108);
nand U24737 (N_24737,N_16889,N_19593);
xor U24738 (N_24738,N_15012,N_18850);
and U24739 (N_24739,N_19300,N_19601);
and U24740 (N_24740,N_16337,N_15677);
nand U24741 (N_24741,N_15884,N_17477);
nor U24742 (N_24742,N_17485,N_19134);
nand U24743 (N_24743,N_15183,N_17543);
and U24744 (N_24744,N_17224,N_16685);
or U24745 (N_24745,N_17142,N_19179);
or U24746 (N_24746,N_18600,N_15726);
nand U24747 (N_24747,N_17546,N_15322);
nor U24748 (N_24748,N_15780,N_17400);
nor U24749 (N_24749,N_17457,N_18126);
and U24750 (N_24750,N_16612,N_18705);
nand U24751 (N_24751,N_16798,N_15346);
and U24752 (N_24752,N_17019,N_17686);
or U24753 (N_24753,N_15312,N_19498);
nand U24754 (N_24754,N_19603,N_18754);
nor U24755 (N_24755,N_19920,N_15634);
nand U24756 (N_24756,N_17052,N_18859);
nor U24757 (N_24757,N_15415,N_19973);
and U24758 (N_24758,N_16321,N_17463);
and U24759 (N_24759,N_18574,N_17937);
or U24760 (N_24760,N_17816,N_16832);
and U24761 (N_24761,N_15968,N_17429);
nor U24762 (N_24762,N_15748,N_16021);
nor U24763 (N_24763,N_15596,N_16328);
nand U24764 (N_24764,N_19043,N_18900);
and U24765 (N_24765,N_17616,N_19225);
and U24766 (N_24766,N_16655,N_18865);
nand U24767 (N_24767,N_17845,N_17812);
or U24768 (N_24768,N_16462,N_15941);
and U24769 (N_24769,N_15567,N_19764);
and U24770 (N_24770,N_18011,N_15582);
and U24771 (N_24771,N_18373,N_15115);
nand U24772 (N_24772,N_19102,N_16908);
or U24773 (N_24773,N_15819,N_16465);
nor U24774 (N_24774,N_18190,N_19888);
or U24775 (N_24775,N_18612,N_16506);
nand U24776 (N_24776,N_19826,N_16341);
nor U24777 (N_24777,N_17062,N_18176);
or U24778 (N_24778,N_19042,N_19320);
and U24779 (N_24779,N_18173,N_18920);
or U24780 (N_24780,N_15319,N_19576);
and U24781 (N_24781,N_15888,N_17336);
nand U24782 (N_24782,N_17402,N_17957);
nor U24783 (N_24783,N_15702,N_17732);
and U24784 (N_24784,N_19062,N_16406);
nor U24785 (N_24785,N_16142,N_18184);
or U24786 (N_24786,N_15958,N_15822);
and U24787 (N_24787,N_18920,N_19560);
nor U24788 (N_24788,N_18967,N_18830);
or U24789 (N_24789,N_19647,N_16160);
nor U24790 (N_24790,N_18194,N_18481);
nand U24791 (N_24791,N_18487,N_19656);
nand U24792 (N_24792,N_19501,N_16738);
nor U24793 (N_24793,N_19935,N_15948);
or U24794 (N_24794,N_18061,N_18243);
and U24795 (N_24795,N_17017,N_16932);
nor U24796 (N_24796,N_17654,N_18677);
nor U24797 (N_24797,N_19493,N_19894);
or U24798 (N_24798,N_16879,N_15122);
and U24799 (N_24799,N_18294,N_19165);
nand U24800 (N_24800,N_19349,N_17568);
nor U24801 (N_24801,N_16831,N_17717);
xnor U24802 (N_24802,N_16216,N_17164);
and U24803 (N_24803,N_16631,N_17691);
nand U24804 (N_24804,N_15869,N_16246);
and U24805 (N_24805,N_19612,N_19800);
nand U24806 (N_24806,N_15587,N_18691);
nor U24807 (N_24807,N_15696,N_16288);
and U24808 (N_24808,N_16228,N_17480);
nand U24809 (N_24809,N_19016,N_19925);
nand U24810 (N_24810,N_18558,N_16867);
and U24811 (N_24811,N_16136,N_18833);
nor U24812 (N_24812,N_19803,N_19445);
nor U24813 (N_24813,N_18128,N_18999);
nor U24814 (N_24814,N_15811,N_17319);
nand U24815 (N_24815,N_19444,N_18786);
nand U24816 (N_24816,N_19088,N_16437);
nand U24817 (N_24817,N_16506,N_15821);
and U24818 (N_24818,N_17810,N_18701);
nand U24819 (N_24819,N_16995,N_18361);
nand U24820 (N_24820,N_17388,N_16746);
nor U24821 (N_24821,N_19528,N_15352);
nor U24822 (N_24822,N_15356,N_19844);
and U24823 (N_24823,N_19505,N_19909);
or U24824 (N_24824,N_17996,N_16187);
or U24825 (N_24825,N_17987,N_18880);
nor U24826 (N_24826,N_15128,N_16967);
or U24827 (N_24827,N_16190,N_15377);
nor U24828 (N_24828,N_19506,N_15799);
nand U24829 (N_24829,N_16874,N_17835);
nand U24830 (N_24830,N_19173,N_18784);
and U24831 (N_24831,N_16884,N_17530);
nor U24832 (N_24832,N_18424,N_19433);
nor U24833 (N_24833,N_17041,N_15753);
nand U24834 (N_24834,N_15795,N_16921);
or U24835 (N_24835,N_16249,N_19109);
or U24836 (N_24836,N_18220,N_17185);
nand U24837 (N_24837,N_19417,N_16610);
nand U24838 (N_24838,N_17684,N_17382);
and U24839 (N_24839,N_15241,N_19933);
or U24840 (N_24840,N_16074,N_17770);
nor U24841 (N_24841,N_17776,N_16890);
or U24842 (N_24842,N_17196,N_19402);
or U24843 (N_24843,N_19956,N_15423);
and U24844 (N_24844,N_19243,N_15604);
and U24845 (N_24845,N_15932,N_17709);
nand U24846 (N_24846,N_16829,N_17121);
nor U24847 (N_24847,N_18361,N_15042);
or U24848 (N_24848,N_15254,N_16543);
nor U24849 (N_24849,N_19441,N_17172);
or U24850 (N_24850,N_19962,N_15213);
and U24851 (N_24851,N_15770,N_18736);
and U24852 (N_24852,N_16698,N_18238);
and U24853 (N_24853,N_19469,N_17507);
and U24854 (N_24854,N_17673,N_19231);
and U24855 (N_24855,N_18779,N_17270);
nand U24856 (N_24856,N_19077,N_15818);
nor U24857 (N_24857,N_19201,N_15911);
and U24858 (N_24858,N_16887,N_18252);
or U24859 (N_24859,N_15375,N_19268);
nand U24860 (N_24860,N_16464,N_16673);
nand U24861 (N_24861,N_15492,N_17506);
or U24862 (N_24862,N_19946,N_19209);
and U24863 (N_24863,N_17431,N_17021);
or U24864 (N_24864,N_18038,N_18389);
or U24865 (N_24865,N_18642,N_19684);
and U24866 (N_24866,N_19166,N_19450);
nand U24867 (N_24867,N_19600,N_17744);
and U24868 (N_24868,N_16112,N_19393);
or U24869 (N_24869,N_18204,N_18732);
and U24870 (N_24870,N_18970,N_15004);
nor U24871 (N_24871,N_16069,N_15700);
or U24872 (N_24872,N_19482,N_18942);
nor U24873 (N_24873,N_18111,N_18465);
nand U24874 (N_24874,N_16604,N_15293);
and U24875 (N_24875,N_16810,N_18278);
nor U24876 (N_24876,N_16197,N_17271);
nor U24877 (N_24877,N_19874,N_16248);
and U24878 (N_24878,N_18214,N_18331);
nand U24879 (N_24879,N_19806,N_17518);
nor U24880 (N_24880,N_18652,N_15682);
and U24881 (N_24881,N_15252,N_16659);
or U24882 (N_24882,N_19403,N_16526);
xnor U24883 (N_24883,N_17682,N_19539);
and U24884 (N_24884,N_19175,N_18795);
and U24885 (N_24885,N_17792,N_19251);
and U24886 (N_24886,N_19986,N_17172);
nand U24887 (N_24887,N_15831,N_18439);
nand U24888 (N_24888,N_18350,N_16249);
nand U24889 (N_24889,N_15828,N_18414);
and U24890 (N_24890,N_16660,N_18376);
nand U24891 (N_24891,N_18887,N_16208);
and U24892 (N_24892,N_19921,N_19968);
nand U24893 (N_24893,N_16750,N_15355);
and U24894 (N_24894,N_18404,N_19985);
and U24895 (N_24895,N_16530,N_17289);
nor U24896 (N_24896,N_17692,N_17712);
xnor U24897 (N_24897,N_18412,N_15324);
xor U24898 (N_24898,N_16809,N_16216);
or U24899 (N_24899,N_17290,N_17186);
or U24900 (N_24900,N_18393,N_15583);
or U24901 (N_24901,N_15189,N_18451);
nor U24902 (N_24902,N_16069,N_15307);
and U24903 (N_24903,N_16088,N_17845);
nor U24904 (N_24904,N_15640,N_15059);
and U24905 (N_24905,N_15622,N_17435);
nand U24906 (N_24906,N_17754,N_18374);
nor U24907 (N_24907,N_17099,N_16137);
or U24908 (N_24908,N_19596,N_18598);
and U24909 (N_24909,N_17706,N_17282);
nand U24910 (N_24910,N_18883,N_17456);
nor U24911 (N_24911,N_15999,N_16044);
nor U24912 (N_24912,N_18193,N_16549);
or U24913 (N_24913,N_17859,N_15920);
nor U24914 (N_24914,N_15855,N_19583);
or U24915 (N_24915,N_18154,N_17839);
or U24916 (N_24916,N_16242,N_18763);
xnor U24917 (N_24917,N_16020,N_17649);
nor U24918 (N_24918,N_18558,N_15957);
nand U24919 (N_24919,N_17014,N_16300);
nand U24920 (N_24920,N_19943,N_15079);
or U24921 (N_24921,N_16782,N_18670);
nor U24922 (N_24922,N_17038,N_19649);
or U24923 (N_24923,N_15616,N_15589);
and U24924 (N_24924,N_18736,N_15704);
nor U24925 (N_24925,N_19552,N_16689);
and U24926 (N_24926,N_15099,N_16786);
nor U24927 (N_24927,N_16142,N_15553);
nor U24928 (N_24928,N_19839,N_18641);
nor U24929 (N_24929,N_18264,N_17957);
or U24930 (N_24930,N_15740,N_15917);
and U24931 (N_24931,N_19675,N_18122);
or U24932 (N_24932,N_15153,N_19281);
nor U24933 (N_24933,N_16011,N_17298);
and U24934 (N_24934,N_17053,N_18047);
nand U24935 (N_24935,N_19505,N_15805);
nor U24936 (N_24936,N_15634,N_16564);
nor U24937 (N_24937,N_18203,N_19862);
nor U24938 (N_24938,N_16256,N_16833);
xor U24939 (N_24939,N_17158,N_18063);
or U24940 (N_24940,N_17993,N_18356);
or U24941 (N_24941,N_15024,N_15928);
and U24942 (N_24942,N_17321,N_17916);
or U24943 (N_24943,N_18437,N_15207);
or U24944 (N_24944,N_18903,N_17502);
and U24945 (N_24945,N_15106,N_17896);
or U24946 (N_24946,N_18547,N_17897);
nor U24947 (N_24947,N_15036,N_15837);
and U24948 (N_24948,N_15378,N_19994);
and U24949 (N_24949,N_17473,N_16401);
or U24950 (N_24950,N_17362,N_18432);
nand U24951 (N_24951,N_15989,N_18025);
nand U24952 (N_24952,N_15182,N_16963);
or U24953 (N_24953,N_17033,N_19010);
and U24954 (N_24954,N_17880,N_17761);
nor U24955 (N_24955,N_16140,N_16564);
nor U24956 (N_24956,N_15153,N_18231);
and U24957 (N_24957,N_16514,N_17649);
and U24958 (N_24958,N_18594,N_18117);
nor U24959 (N_24959,N_18574,N_18669);
or U24960 (N_24960,N_16030,N_18659);
and U24961 (N_24961,N_17372,N_19485);
and U24962 (N_24962,N_18599,N_17451);
nor U24963 (N_24963,N_16527,N_16026);
or U24964 (N_24964,N_15773,N_19745);
nor U24965 (N_24965,N_17729,N_15799);
nand U24966 (N_24966,N_15376,N_17901);
nand U24967 (N_24967,N_17346,N_18230);
or U24968 (N_24968,N_19644,N_19035);
nor U24969 (N_24969,N_17363,N_16005);
nand U24970 (N_24970,N_18527,N_19402);
or U24971 (N_24971,N_16864,N_18188);
or U24972 (N_24972,N_15313,N_15762);
nand U24973 (N_24973,N_15154,N_15324);
and U24974 (N_24974,N_18439,N_15897);
and U24975 (N_24975,N_19992,N_16984);
and U24976 (N_24976,N_15211,N_18212);
or U24977 (N_24977,N_18428,N_19425);
or U24978 (N_24978,N_18353,N_18651);
nand U24979 (N_24979,N_16960,N_17597);
and U24980 (N_24980,N_17348,N_16104);
nand U24981 (N_24981,N_18012,N_16044);
nor U24982 (N_24982,N_18228,N_17471);
nand U24983 (N_24983,N_19364,N_16845);
and U24984 (N_24984,N_18248,N_19127);
nand U24985 (N_24985,N_16813,N_17669);
nand U24986 (N_24986,N_17360,N_17794);
nand U24987 (N_24987,N_19361,N_19665);
or U24988 (N_24988,N_15439,N_17748);
nor U24989 (N_24989,N_17499,N_19383);
and U24990 (N_24990,N_15426,N_17354);
or U24991 (N_24991,N_17766,N_15117);
or U24992 (N_24992,N_19652,N_16050);
nor U24993 (N_24993,N_17993,N_17758);
or U24994 (N_24994,N_18983,N_19659);
and U24995 (N_24995,N_17952,N_19593);
xnor U24996 (N_24996,N_19095,N_17692);
nand U24997 (N_24997,N_19144,N_19760);
nand U24998 (N_24998,N_15305,N_15217);
nor U24999 (N_24999,N_15482,N_19604);
nand UO_0 (O_0,N_20525,N_20111);
nor UO_1 (O_1,N_20671,N_21585);
nand UO_2 (O_2,N_24928,N_21481);
and UO_3 (O_3,N_23057,N_24096);
or UO_4 (O_4,N_22686,N_22587);
nand UO_5 (O_5,N_23589,N_20184);
nor UO_6 (O_6,N_21403,N_23811);
or UO_7 (O_7,N_22068,N_21531);
nor UO_8 (O_8,N_20674,N_21970);
nor UO_9 (O_9,N_20363,N_20771);
nand UO_10 (O_10,N_21544,N_20832);
nand UO_11 (O_11,N_22949,N_22244);
or UO_12 (O_12,N_24056,N_23067);
and UO_13 (O_13,N_22185,N_21751);
and UO_14 (O_14,N_21573,N_24880);
or UO_15 (O_15,N_24514,N_22164);
or UO_16 (O_16,N_22798,N_21662);
nand UO_17 (O_17,N_21789,N_20926);
nand UO_18 (O_18,N_23689,N_20396);
nand UO_19 (O_19,N_20319,N_23395);
and UO_20 (O_20,N_22089,N_23341);
nor UO_21 (O_21,N_22825,N_20931);
or UO_22 (O_22,N_23820,N_22869);
nor UO_23 (O_23,N_23650,N_22778);
nor UO_24 (O_24,N_21809,N_24165);
nand UO_25 (O_25,N_20117,N_21724);
nand UO_26 (O_26,N_23005,N_20008);
nor UO_27 (O_27,N_23239,N_22521);
nor UO_28 (O_28,N_22732,N_22119);
or UO_29 (O_29,N_22104,N_21367);
and UO_30 (O_30,N_21607,N_21208);
nor UO_31 (O_31,N_24859,N_20633);
or UO_32 (O_32,N_22930,N_21060);
or UO_33 (O_33,N_20435,N_23045);
and UO_34 (O_34,N_20238,N_23946);
nand UO_35 (O_35,N_22787,N_23298);
nand UO_36 (O_36,N_20989,N_23289);
and UO_37 (O_37,N_20880,N_22613);
nand UO_38 (O_38,N_20245,N_22906);
and UO_39 (O_39,N_24682,N_22756);
and UO_40 (O_40,N_21292,N_24889);
and UO_41 (O_41,N_21828,N_23934);
xnor UO_42 (O_42,N_20826,N_24585);
xnor UO_43 (O_43,N_24438,N_20770);
nand UO_44 (O_44,N_20107,N_24727);
nor UO_45 (O_45,N_20146,N_22877);
or UO_46 (O_46,N_23106,N_20376);
nand UO_47 (O_47,N_21555,N_23714);
nor UO_48 (O_48,N_24753,N_23938);
nand UO_49 (O_49,N_23182,N_23889);
xnor UO_50 (O_50,N_22811,N_22920);
nand UO_51 (O_51,N_22602,N_21890);
xor UO_52 (O_52,N_20666,N_20683);
or UO_53 (O_53,N_21342,N_21779);
and UO_54 (O_54,N_23685,N_24846);
and UO_55 (O_55,N_22248,N_21407);
and UO_56 (O_56,N_24146,N_24273);
or UO_57 (O_57,N_24281,N_24788);
or UO_58 (O_58,N_23090,N_24308);
or UO_59 (O_59,N_20642,N_23129);
or UO_60 (O_60,N_22017,N_21543);
nand UO_61 (O_61,N_20461,N_21119);
and UO_62 (O_62,N_22132,N_22958);
or UO_63 (O_63,N_24492,N_24774);
or UO_64 (O_64,N_23133,N_24093);
and UO_65 (O_65,N_23291,N_22243);
nand UO_66 (O_66,N_23127,N_23603);
nor UO_67 (O_67,N_22036,N_21478);
nor UO_68 (O_68,N_22428,N_23764);
and UO_69 (O_69,N_24521,N_24245);
nand UO_70 (O_70,N_20788,N_22421);
and UO_71 (O_71,N_22166,N_22658);
and UO_72 (O_72,N_20263,N_24848);
and UO_73 (O_73,N_24470,N_20682);
or UO_74 (O_74,N_20240,N_23619);
and UO_75 (O_75,N_22504,N_22139);
nand UO_76 (O_76,N_23211,N_23237);
nand UO_77 (O_77,N_22968,N_22010);
or UO_78 (O_78,N_24478,N_22302);
or UO_79 (O_79,N_24431,N_23943);
nand UO_80 (O_80,N_22839,N_23741);
and UO_81 (O_81,N_22843,N_23085);
nor UO_82 (O_82,N_23215,N_21755);
or UO_83 (O_83,N_24795,N_24474);
nand UO_84 (O_84,N_23801,N_22537);
and UO_85 (O_85,N_21620,N_22256);
nor UO_86 (O_86,N_23302,N_22468);
nand UO_87 (O_87,N_22300,N_22404);
nand UO_88 (O_88,N_24396,N_20566);
nand UO_89 (O_89,N_23144,N_23868);
and UO_90 (O_90,N_22519,N_24124);
and UO_91 (O_91,N_20650,N_20852);
nand UO_92 (O_92,N_23773,N_22129);
nor UO_93 (O_93,N_24183,N_24824);
or UO_94 (O_94,N_20743,N_23558);
or UO_95 (O_95,N_21784,N_23951);
and UO_96 (O_96,N_24404,N_20944);
and UO_97 (O_97,N_20897,N_22650);
nand UO_98 (O_98,N_20795,N_22826);
xnor UO_99 (O_99,N_23489,N_23798);
or UO_100 (O_100,N_23678,N_23973);
and UO_101 (O_101,N_21732,N_21722);
nor UO_102 (O_102,N_22317,N_22853);
nand UO_103 (O_103,N_24525,N_21864);
and UO_104 (O_104,N_23337,N_23830);
nor UO_105 (O_105,N_20802,N_22518);
nor UO_106 (O_106,N_24809,N_21632);
nand UO_107 (O_107,N_24046,N_20908);
nor UO_108 (O_108,N_20651,N_20123);
and UO_109 (O_109,N_20491,N_23480);
nand UO_110 (O_110,N_23561,N_22861);
or UO_111 (O_111,N_22603,N_23340);
or UO_112 (O_112,N_21856,N_24511);
or UO_113 (O_113,N_23674,N_20206);
nand UO_114 (O_114,N_24131,N_21140);
or UO_115 (O_115,N_24054,N_20617);
nand UO_116 (O_116,N_20954,N_23931);
xor UO_117 (O_117,N_20344,N_21390);
and UO_118 (O_118,N_20096,N_22580);
nor UO_119 (O_119,N_20160,N_24415);
nor UO_120 (O_120,N_22402,N_22560);
and UO_121 (O_121,N_21595,N_21214);
or UO_122 (O_122,N_23383,N_22640);
nor UO_123 (O_123,N_21319,N_24696);
nor UO_124 (O_124,N_24224,N_24570);
nor UO_125 (O_125,N_24445,N_20723);
nand UO_126 (O_126,N_24121,N_21956);
nand UO_127 (O_127,N_24579,N_21947);
nor UO_128 (O_128,N_21736,N_22279);
nand UO_129 (O_129,N_22507,N_22005);
nand UO_130 (O_130,N_20892,N_22750);
or UO_131 (O_131,N_23673,N_22437);
or UO_132 (O_132,N_21758,N_23817);
xor UO_133 (O_133,N_22349,N_20275);
and UO_134 (O_134,N_23040,N_22733);
nand UO_135 (O_135,N_20993,N_23477);
nor UO_136 (O_136,N_23010,N_20505);
nor UO_137 (O_137,N_20321,N_21220);
nand UO_138 (O_138,N_23012,N_21217);
or UO_139 (O_139,N_24671,N_20133);
or UO_140 (O_140,N_23802,N_23424);
or UO_141 (O_141,N_23479,N_21527);
nand UO_142 (O_142,N_24296,N_24238);
nor UO_143 (O_143,N_21932,N_24412);
and UO_144 (O_144,N_20046,N_22143);
nand UO_145 (O_145,N_24625,N_23353);
nor UO_146 (O_146,N_21160,N_21347);
or UO_147 (O_147,N_22395,N_20974);
or UO_148 (O_148,N_21392,N_20937);
and UO_149 (O_149,N_20958,N_22035);
nand UO_150 (O_150,N_21584,N_22142);
nor UO_151 (O_151,N_21039,N_22335);
nor UO_152 (O_152,N_20867,N_24651);
nand UO_153 (O_153,N_20113,N_22022);
or UO_154 (O_154,N_24029,N_23908);
and UO_155 (O_155,N_23474,N_22873);
or UO_156 (O_156,N_20393,N_23055);
nand UO_157 (O_157,N_20627,N_24354);
or UO_158 (O_158,N_20398,N_24299);
or UO_159 (O_159,N_22378,N_22969);
or UO_160 (O_160,N_20138,N_22148);
or UO_161 (O_161,N_21993,N_21882);
and UO_162 (O_162,N_23398,N_22495);
or UO_163 (O_163,N_20475,N_22170);
nor UO_164 (O_164,N_21193,N_24644);
and UO_165 (O_165,N_23418,N_23739);
or UO_166 (O_166,N_20091,N_21631);
and UO_167 (O_167,N_20988,N_20140);
nand UO_168 (O_168,N_23945,N_24145);
nor UO_169 (O_169,N_24469,N_21763);
nand UO_170 (O_170,N_21453,N_20135);
nor UO_171 (O_171,N_20131,N_20220);
or UO_172 (O_172,N_23980,N_23692);
and UO_173 (O_173,N_23833,N_20065);
and UO_174 (O_174,N_22789,N_23156);
nor UO_175 (O_175,N_21258,N_21004);
nand UO_176 (O_176,N_24444,N_23781);
nor UO_177 (O_177,N_24855,N_21357);
nand UO_178 (O_178,N_21752,N_21984);
or UO_179 (O_179,N_23136,N_21023);
nand UO_180 (O_180,N_24003,N_22784);
nand UO_181 (O_181,N_21723,N_21615);
or UO_182 (O_182,N_20447,N_24302);
nor UO_183 (O_183,N_20241,N_20553);
or UO_184 (O_184,N_22541,N_21561);
or UO_185 (O_185,N_20576,N_22528);
xor UO_186 (O_186,N_22846,N_21647);
nand UO_187 (O_187,N_23132,N_24668);
nor UO_188 (O_188,N_20339,N_23111);
and UO_189 (O_189,N_20596,N_24256);
nor UO_190 (O_190,N_23548,N_20468);
or UO_191 (O_191,N_22590,N_21688);
and UO_192 (O_192,N_24242,N_20702);
or UO_193 (O_193,N_22701,N_22891);
nand UO_194 (O_194,N_21735,N_23009);
or UO_195 (O_195,N_22351,N_24631);
nand UO_196 (O_196,N_21548,N_22200);
or UO_197 (O_197,N_24058,N_23879);
or UO_198 (O_198,N_20521,N_23500);
nor UO_199 (O_199,N_21813,N_21151);
nand UO_200 (O_200,N_23385,N_22411);
or UO_201 (O_201,N_23568,N_23587);
and UO_202 (O_202,N_23691,N_23078);
nand UO_203 (O_203,N_23499,N_23876);
nand UO_204 (O_204,N_23197,N_21501);
or UO_205 (O_205,N_24297,N_22074);
or UO_206 (O_206,N_22190,N_23074);
or UO_207 (O_207,N_22172,N_24070);
nor UO_208 (O_208,N_24317,N_20610);
nand UO_209 (O_209,N_24214,N_20174);
nand UO_210 (O_210,N_24346,N_21457);
and UO_211 (O_211,N_24035,N_22994);
nand UO_212 (O_212,N_24999,N_22597);
nand UO_213 (O_213,N_20535,N_24883);
nand UO_214 (O_214,N_23485,N_21408);
or UO_215 (O_215,N_23458,N_21569);
nand UO_216 (O_216,N_21502,N_20038);
nor UO_217 (O_217,N_20394,N_22015);
nand UO_218 (O_218,N_20044,N_21931);
or UO_219 (O_219,N_21883,N_24202);
nor UO_220 (O_220,N_23483,N_24482);
nor UO_221 (O_221,N_21166,N_24887);
nand UO_222 (O_222,N_21795,N_21935);
nand UO_223 (O_223,N_21837,N_21154);
nor UO_224 (O_224,N_22236,N_22814);
nand UO_225 (O_225,N_20580,N_24698);
and UO_226 (O_226,N_23999,N_20865);
or UO_227 (O_227,N_20209,N_22183);
nor UO_228 (O_228,N_21134,N_23233);
nand UO_229 (O_229,N_22888,N_23170);
nand UO_230 (O_230,N_22088,N_24140);
nand UO_231 (O_231,N_23818,N_20463);
nor UO_232 (O_232,N_22283,N_24501);
or UO_233 (O_233,N_20712,N_24784);
or UO_234 (O_234,N_21974,N_22127);
or UO_235 (O_235,N_20512,N_22358);
or UO_236 (O_236,N_24462,N_20186);
nor UO_237 (O_237,N_24369,N_23601);
or UO_238 (O_238,N_22987,N_22517);
nand UO_239 (O_239,N_22707,N_23331);
or UO_240 (O_240,N_20243,N_22638);
or UO_241 (O_241,N_20656,N_22633);
and UO_242 (O_242,N_21575,N_24991);
or UO_243 (O_243,N_21441,N_21131);
xor UO_244 (O_244,N_20382,N_21097);
nor UO_245 (O_245,N_21719,N_22496);
nand UO_246 (O_246,N_23583,N_20458);
nor UO_247 (O_247,N_24742,N_20011);
xor UO_248 (O_248,N_23232,N_21395);
nor UO_249 (O_249,N_21650,N_20711);
nand UO_250 (O_250,N_24132,N_20102);
or UO_251 (O_251,N_21571,N_22165);
nand UO_252 (O_252,N_24418,N_23274);
nand UO_253 (O_253,N_24832,N_23244);
nand UO_254 (O_254,N_23723,N_21138);
nor UO_255 (O_255,N_23544,N_20957);
nand UO_256 (O_256,N_22914,N_24507);
nor UO_257 (O_257,N_24216,N_23588);
or UO_258 (O_258,N_24122,N_22693);
and UO_259 (O_259,N_23929,N_22585);
and UO_260 (O_260,N_21918,N_20717);
nor UO_261 (O_261,N_22531,N_24149);
nor UO_262 (O_262,N_23081,N_24437);
nand UO_263 (O_263,N_21877,N_21398);
and UO_264 (O_264,N_24884,N_20597);
and UO_265 (O_265,N_21876,N_23667);
or UO_266 (O_266,N_22217,N_21169);
or UO_267 (O_267,N_24375,N_21269);
and UO_268 (O_268,N_23018,N_21000);
nand UO_269 (O_269,N_21659,N_22651);
nand UO_270 (O_270,N_23837,N_22067);
nand UO_271 (O_271,N_23357,N_24882);
and UO_272 (O_272,N_20188,N_20381);
xor UO_273 (O_273,N_24152,N_24740);
and UO_274 (O_274,N_22957,N_21845);
nor UO_275 (O_275,N_24810,N_21272);
and UO_276 (O_276,N_23482,N_22940);
and UO_277 (O_277,N_22672,N_21605);
nor UO_278 (O_278,N_24173,N_22614);
nand UO_279 (O_279,N_22193,N_22373);
nand UO_280 (O_280,N_23853,N_24630);
nand UO_281 (O_281,N_22357,N_21898);
or UO_282 (O_282,N_23841,N_20121);
or UO_283 (O_283,N_24968,N_21149);
nand UO_284 (O_284,N_21144,N_23854);
nor UO_285 (O_285,N_21657,N_22099);
or UO_286 (O_286,N_23622,N_21400);
nand UO_287 (O_287,N_21069,N_24190);
nand UO_288 (O_288,N_20699,N_22607);
nand UO_289 (O_289,N_23644,N_23140);
nand UO_290 (O_290,N_20756,N_23697);
or UO_291 (O_291,N_22606,N_23034);
nand UO_292 (O_292,N_23276,N_23217);
nand UO_293 (O_293,N_23070,N_21838);
or UO_294 (O_294,N_21022,N_21293);
or UO_295 (O_295,N_21579,N_21165);
or UO_296 (O_296,N_22838,N_22400);
and UO_297 (O_297,N_24557,N_22716);
nand UO_298 (O_298,N_24687,N_23297);
nor UO_299 (O_299,N_24179,N_24863);
nor UO_300 (O_300,N_22092,N_20840);
nor UO_301 (O_301,N_21881,N_22026);
nor UO_302 (O_302,N_21903,N_21899);
and UO_303 (O_303,N_22550,N_20839);
or UO_304 (O_304,N_24076,N_21827);
and UO_305 (O_305,N_22128,N_23962);
and UO_306 (O_306,N_22458,N_21284);
or UO_307 (O_307,N_21373,N_23570);
nand UO_308 (O_308,N_21841,N_20436);
nor UO_309 (O_309,N_21093,N_22626);
or UO_310 (O_310,N_24372,N_23277);
nand UO_311 (O_311,N_20779,N_24107);
and UO_312 (O_312,N_24321,N_24272);
nand UO_313 (O_313,N_22616,N_24204);
and UO_314 (O_314,N_23584,N_24148);
nor UO_315 (O_315,N_21787,N_24294);
and UO_316 (O_316,N_20152,N_24429);
and UO_317 (O_317,N_22058,N_21674);
nand UO_318 (O_318,N_20498,N_20349);
nand UO_319 (O_319,N_24258,N_24324);
or UO_320 (O_320,N_20546,N_21721);
and UO_321 (O_321,N_20303,N_24397);
or UO_322 (O_322,N_21793,N_20324);
nor UO_323 (O_323,N_22231,N_23971);
nor UO_324 (O_324,N_22485,N_21744);
nor UO_325 (O_325,N_20595,N_24279);
and UO_326 (O_326,N_21690,N_20000);
xor UO_327 (O_327,N_22145,N_24754);
nand UO_328 (O_328,N_22513,N_21622);
or UO_329 (O_329,N_22600,N_23778);
or UO_330 (O_330,N_24471,N_24390);
nand UO_331 (O_331,N_20979,N_24508);
and UO_332 (O_332,N_24476,N_23271);
or UO_333 (O_333,N_24506,N_21334);
nand UO_334 (O_334,N_24971,N_23702);
nor UO_335 (O_335,N_22298,N_23826);
nor UO_336 (O_336,N_20945,N_20244);
nor UO_337 (O_337,N_24876,N_20934);
nand UO_338 (O_338,N_21546,N_23662);
or UO_339 (O_339,N_20385,N_22188);
and UO_340 (O_340,N_20713,N_24684);
or UO_341 (O_341,N_21172,N_21218);
nor UO_342 (O_342,N_24167,N_21849);
nor UO_343 (O_343,N_24974,N_21871);
and UO_344 (O_344,N_20611,N_21757);
or UO_345 (O_345,N_22316,N_24691);
and UO_346 (O_346,N_21901,N_24681);
nand UO_347 (O_347,N_24161,N_21461);
nor UO_348 (O_348,N_22117,N_22682);
or UO_349 (O_349,N_21912,N_20480);
and UO_350 (O_350,N_22448,N_20659);
nor UO_351 (O_351,N_24977,N_20169);
and UO_352 (O_352,N_23746,N_23659);
and UO_353 (O_353,N_24979,N_21568);
and UO_354 (O_354,N_24878,N_21627);
or UO_355 (O_355,N_24075,N_22084);
and UO_356 (O_356,N_24472,N_23449);
and UO_357 (O_357,N_23135,N_20478);
and UO_358 (O_358,N_20946,N_24268);
nor UO_359 (O_359,N_23310,N_23982);
nor UO_360 (O_360,N_23473,N_20959);
and UO_361 (O_361,N_20714,N_24356);
nand UO_362 (O_362,N_23615,N_20272);
nor UO_363 (O_363,N_24073,N_23661);
or UO_364 (O_364,N_24153,N_20759);
nand UO_365 (O_365,N_20833,N_24042);
nor UO_366 (O_366,N_21071,N_20088);
nand UO_367 (O_367,N_21102,N_23236);
nand UO_368 (O_368,N_23719,N_22628);
nor UO_369 (O_369,N_20502,N_21634);
nor UO_370 (O_370,N_23141,N_23896);
and UO_371 (O_371,N_20551,N_23911);
nand UO_372 (O_372,N_23953,N_24331);
or UO_373 (O_373,N_24722,N_22858);
or UO_374 (O_374,N_21368,N_21547);
nor UO_375 (O_375,N_21613,N_20312);
and UO_376 (O_376,N_22024,N_20027);
or UO_377 (O_377,N_21678,N_20780);
or UO_378 (O_378,N_24293,N_20718);
nand UO_379 (O_379,N_23947,N_23326);
or UO_380 (O_380,N_20401,N_24419);
or UO_381 (O_381,N_23162,N_22227);
and UO_382 (O_382,N_24959,N_21670);
or UO_383 (O_383,N_20686,N_23950);
nand UO_384 (O_384,N_23177,N_23635);
and UO_385 (O_385,N_24633,N_20001);
and UO_386 (O_386,N_24729,N_22163);
nor UO_387 (O_387,N_21243,N_22424);
and UO_388 (O_388,N_20690,N_21957);
nand UO_389 (O_389,N_23623,N_21337);
nor UO_390 (O_390,N_21636,N_20167);
nand UO_391 (O_391,N_21648,N_22834);
nor UO_392 (O_392,N_23776,N_23035);
nor UO_393 (O_393,N_22044,N_24209);
and UO_394 (O_394,N_24700,N_23373);
nand UO_395 (O_395,N_23142,N_21550);
nand UO_396 (O_396,N_21282,N_21851);
and UO_397 (O_397,N_23567,N_24637);
or UO_398 (O_398,N_24561,N_22340);
and UO_399 (O_399,N_23810,N_22352);
nor UO_400 (O_400,N_22294,N_22813);
and UO_401 (O_401,N_20757,N_23284);
nor UO_402 (O_402,N_23541,N_24674);
or UO_403 (O_403,N_24866,N_24617);
or UO_404 (O_404,N_22649,N_23419);
nor UO_405 (O_405,N_21391,N_21557);
nor UO_406 (O_406,N_23348,N_22123);
or UO_407 (O_407,N_22558,N_24718);
xnor UO_408 (O_408,N_24648,N_24213);
and UO_409 (O_409,N_24484,N_24624);
or UO_410 (O_410,N_21271,N_22624);
nor UO_411 (O_411,N_21366,N_23161);
or UO_412 (O_412,N_23105,N_21860);
and UO_413 (O_413,N_24931,N_22105);
or UO_414 (O_414,N_20609,N_24577);
or UO_415 (O_415,N_22187,N_23308);
or UO_416 (O_416,N_21741,N_24839);
or UO_417 (O_417,N_20293,N_22848);
and UO_418 (O_418,N_23439,N_20271);
nor UO_419 (O_419,N_20900,N_20256);
and UO_420 (O_420,N_20288,N_20752);
and UO_421 (O_421,N_21139,N_24353);
nor UO_422 (O_422,N_21645,N_21431);
or UO_423 (O_423,N_21742,N_22175);
or UO_424 (O_424,N_24379,N_24546);
nand UO_425 (O_425,N_20591,N_24384);
and UO_426 (O_426,N_20040,N_23607);
nor UO_427 (O_427,N_20786,N_21710);
nand UO_428 (O_428,N_23511,N_20308);
and UO_429 (O_429,N_20998,N_21812);
or UO_430 (O_430,N_20857,N_20986);
nand UO_431 (O_431,N_21188,N_23430);
nand UO_432 (O_432,N_23509,N_23434);
and UO_433 (O_433,N_21892,N_24914);
and UO_434 (O_434,N_23243,N_23145);
or UO_435 (O_435,N_20790,N_22039);
nand UO_436 (O_436,N_23375,N_20049);
nor UO_437 (O_437,N_21425,N_20261);
nor UO_438 (O_438,N_21536,N_24626);
or UO_439 (O_439,N_24694,N_21082);
nor UO_440 (O_440,N_23917,N_22765);
nor UO_441 (O_441,N_21798,N_21640);
and UO_442 (O_442,N_20493,N_22241);
and UO_443 (O_443,N_21232,N_22601);
nor UO_444 (O_444,N_22678,N_24589);
nand UO_445 (O_445,N_22636,N_21381);
nor UO_446 (O_446,N_21331,N_24237);
nor UO_447 (O_447,N_22896,N_22997);
nand UO_448 (O_448,N_21517,N_20687);
and UO_449 (O_449,N_22345,N_24735);
and UO_450 (O_450,N_21580,N_24995);
nand UO_451 (O_451,N_22492,N_23964);
and UO_452 (O_452,N_21668,N_20539);
or UO_453 (O_453,N_24360,N_21534);
or UO_454 (O_454,N_20175,N_20289);
or UO_455 (O_455,N_20421,N_22396);
nand UO_456 (O_456,N_21929,N_20368);
and UO_457 (O_457,N_22878,N_22330);
nor UO_458 (O_458,N_22618,N_22717);
or UO_459 (O_459,N_22456,N_24115);
nand UO_460 (O_460,N_20004,N_20537);
nor UO_461 (O_461,N_20388,N_23463);
or UO_462 (O_462,N_22368,N_20248);
and UO_463 (O_463,N_20487,N_24551);
or UO_464 (O_464,N_21709,N_24162);
or UO_465 (O_465,N_24678,N_24826);
or UO_466 (O_466,N_22274,N_21486);
nand UO_467 (O_467,N_23576,N_21158);
nand UO_468 (O_468,N_23013,N_24447);
xor UO_469 (O_469,N_21302,N_20700);
or UO_470 (O_470,N_22252,N_24013);
and UO_471 (O_471,N_24225,N_21551);
xnor UO_472 (O_472,N_21869,N_23775);
nand UO_473 (O_473,N_23175,N_22598);
and UO_474 (O_474,N_22939,N_21317);
or UO_475 (O_475,N_22648,N_22107);
and UO_476 (O_476,N_23272,N_23311);
nand UO_477 (O_477,N_20348,N_22427);
nor UO_478 (O_478,N_20522,N_21835);
and UO_479 (O_479,N_21926,N_23454);
and UO_480 (O_480,N_20777,N_20429);
nor UO_481 (O_481,N_21848,N_23201);
or UO_482 (O_482,N_23645,N_23977);
and UO_483 (O_483,N_24236,N_20587);
and UO_484 (O_484,N_24591,N_23362);
or UO_485 (O_485,N_23916,N_22786);
nor UO_486 (O_486,N_23796,N_23376);
or UO_487 (O_487,N_23414,N_21048);
and UO_488 (O_488,N_21987,N_21930);
nand UO_489 (O_489,N_20875,N_20103);
xor UO_490 (O_490,N_22309,N_23073);
nor UO_491 (O_491,N_20215,N_22670);
or UO_492 (O_492,N_20407,N_24038);
nor UO_493 (O_493,N_21663,N_24730);
and UO_494 (O_494,N_21072,N_22239);
nand UO_495 (O_495,N_22312,N_21906);
nor UO_496 (O_496,N_22741,N_21460);
nor UO_497 (O_497,N_20932,N_22720);
or UO_498 (O_498,N_23008,N_23562);
nand UO_499 (O_499,N_20819,N_23805);
or UO_500 (O_500,N_21846,N_22574);
nor UO_501 (O_501,N_20267,N_20056);
or UO_502 (O_502,N_21018,N_24203);
and UO_503 (O_503,N_21333,N_22703);
or UO_504 (O_504,N_22779,N_21730);
nand UO_505 (O_505,N_20701,N_21565);
or UO_506 (O_506,N_22277,N_24166);
or UO_507 (O_507,N_20063,N_24329);
nor UO_508 (O_508,N_21281,N_23523);
nand UO_509 (O_509,N_21937,N_20424);
nand UO_510 (O_510,N_23351,N_22833);
nor UO_511 (O_511,N_21513,N_24187);
nor UO_512 (O_512,N_22000,N_21896);
and UO_513 (O_513,N_21737,N_22904);
xnor UO_514 (O_514,N_20903,N_20622);
and UO_515 (O_515,N_21420,N_21372);
nor UO_516 (O_516,N_22802,N_24665);
or UO_517 (O_517,N_21163,N_20961);
or UO_518 (O_518,N_24271,N_23037);
nand UO_519 (O_519,N_24782,N_24583);
and UO_520 (O_520,N_23611,N_24207);
nor UO_521 (O_521,N_24374,N_23745);
nor UO_522 (O_522,N_22532,N_21982);
and UO_523 (O_523,N_21338,N_23188);
or UO_524 (O_524,N_21278,N_21429);
or UO_525 (O_525,N_21897,N_22118);
and UO_526 (O_526,N_22646,N_22069);
or UO_527 (O_527,N_23226,N_21191);
xnor UO_528 (O_528,N_23264,N_21637);
and UO_529 (O_529,N_22526,N_23168);
or UO_530 (O_530,N_20246,N_22662);
nor UO_531 (O_531,N_21181,N_24015);
xor UO_532 (O_532,N_23065,N_20799);
nand UO_533 (O_533,N_22898,N_21270);
xor UO_534 (O_534,N_21308,N_20097);
nand UO_535 (O_535,N_20637,N_20772);
or UO_536 (O_536,N_20078,N_23116);
nand UO_537 (O_537,N_23671,N_24840);
nand UO_538 (O_538,N_20859,N_22261);
and UO_539 (O_539,N_20952,N_22554);
or UO_540 (O_540,N_20895,N_20171);
xor UO_541 (O_541,N_24241,N_23800);
or UO_542 (O_542,N_21448,N_23604);
or UO_543 (O_543,N_20504,N_20406);
or UO_544 (O_544,N_21796,N_21008);
nand UO_545 (O_545,N_22182,N_23641);
and UO_546 (O_546,N_24661,N_22311);
nand UO_547 (O_547,N_23757,N_22296);
and UO_548 (O_548,N_24695,N_23718);
nand UO_549 (O_549,N_22643,N_24950);
nor UO_550 (O_550,N_22795,N_21245);
nor UO_551 (O_551,N_23287,N_24018);
or UO_552 (O_552,N_21424,N_20812);
and UO_553 (O_553,N_23543,N_22667);
and UO_554 (O_554,N_22520,N_23266);
nand UO_555 (O_555,N_24969,N_23052);
nand UO_556 (O_556,N_21287,N_23769);
nor UO_557 (O_557,N_24796,N_24504);
xnor UO_558 (O_558,N_21529,N_24697);
or UO_559 (O_559,N_22555,N_23557);
nor UO_560 (O_560,N_23748,N_24243);
nor UO_561 (O_561,N_22307,N_24389);
or UO_562 (O_562,N_20888,N_20231);
nand UO_563 (O_563,N_24806,N_24232);
nor UO_564 (O_564,N_21351,N_23921);
nor UO_565 (O_565,N_22933,N_20423);
nand UO_566 (O_566,N_24976,N_23501);
xnor UO_567 (O_567,N_20531,N_24543);
nand UO_568 (O_568,N_23762,N_21012);
nand UO_569 (O_569,N_20471,N_22131);
or UO_570 (O_570,N_21275,N_21981);
and UO_571 (O_571,N_24467,N_24021);
and UO_572 (O_572,N_23360,N_23265);
nor UO_573 (O_573,N_23026,N_20644);
or UO_574 (O_574,N_20939,N_21010);
nor UO_575 (O_575,N_20473,N_21764);
nor UO_576 (O_576,N_22505,N_21754);
nand UO_577 (O_577,N_21041,N_20544);
or UO_578 (O_578,N_23267,N_22057);
nand UO_579 (O_579,N_23679,N_23970);
or UO_580 (O_580,N_22559,N_23785);
nand UO_581 (O_581,N_23758,N_21156);
nand UO_582 (O_582,N_20066,N_20764);
and UO_583 (O_583,N_21038,N_23328);
nand UO_584 (O_584,N_21803,N_22223);
and UO_585 (O_585,N_23595,N_22950);
nand UO_586 (O_586,N_20100,N_23218);
and UO_587 (O_587,N_23147,N_21867);
nand UO_588 (O_588,N_24539,N_21174);
or UO_589 (O_589,N_23514,N_24160);
and UO_590 (O_590,N_21988,N_24526);
nor UO_591 (O_591,N_20161,N_24082);
nand UO_592 (O_592,N_22673,N_20698);
and UO_593 (O_593,N_20605,N_21248);
and UO_594 (O_594,N_21108,N_23639);
or UO_595 (O_595,N_22253,N_22557);
and UO_596 (O_596,N_21850,N_22674);
nand UO_597 (O_597,N_20549,N_23782);
nor UO_598 (O_598,N_22301,N_20028);
or UO_599 (O_599,N_21223,N_23436);
nand UO_600 (O_600,N_23209,N_22721);
nor UO_601 (O_601,N_23877,N_24803);
nor UO_602 (O_602,N_20125,N_22641);
nor UO_603 (O_603,N_23347,N_20373);
nor UO_604 (O_604,N_21405,N_20536);
or UO_605 (O_605,N_22919,N_23327);
nor UO_606 (O_606,N_22233,N_21944);
and UO_607 (O_607,N_24807,N_21055);
or UO_608 (O_608,N_23143,N_23028);
nand UO_609 (O_609,N_20709,N_24421);
and UO_610 (O_610,N_20176,N_20089);
or UO_611 (O_611,N_23149,N_22791);
and UO_612 (O_612,N_24049,N_20681);
or UO_613 (O_613,N_24911,N_21578);
and UO_614 (O_614,N_21066,N_21076);
nand UO_615 (O_615,N_20408,N_22540);
or UO_616 (O_616,N_23521,N_20559);
nor UO_617 (O_617,N_24065,N_24494);
or UO_618 (O_618,N_20798,N_23126);
and UO_619 (O_619,N_23752,N_21075);
or UO_620 (O_620,N_23952,N_22016);
or UO_621 (O_621,N_23858,N_21115);
and UO_622 (O_622,N_24201,N_23616);
or UO_623 (O_623,N_20070,N_21888);
nor UO_624 (O_624,N_22893,N_22006);
or UO_625 (O_625,N_22880,N_24240);
nor UO_626 (O_626,N_22377,N_20023);
nand UO_627 (O_627,N_21748,N_21350);
nor UO_628 (O_628,N_21002,N_24770);
nand UO_629 (O_629,N_24143,N_22281);
nand UO_630 (O_630,N_21747,N_24408);
nand UO_631 (O_631,N_24420,N_21179);
nor UO_632 (O_632,N_20302,N_22980);
or UO_633 (O_633,N_24292,N_24212);
and UO_634 (O_634,N_23356,N_24712);
nand UO_635 (O_635,N_24274,N_21475);
nor UO_636 (O_636,N_23246,N_21161);
xnor UO_637 (O_637,N_23756,N_22125);
nor UO_638 (O_638,N_21304,N_24123);
nor UO_639 (O_639,N_21697,N_24027);
and UO_640 (O_640,N_22868,N_24886);
nor UO_641 (O_641,N_23680,N_23316);
nor UO_642 (O_642,N_20459,N_21263);
or UO_643 (O_643,N_20470,N_24517);
nand UO_644 (O_644,N_23415,N_24983);
or UO_645 (O_645,N_23221,N_21325);
nor UO_646 (O_646,N_23153,N_21875);
nand UO_647 (O_647,N_23549,N_24210);
or UO_648 (O_648,N_23783,N_24023);
xor UO_649 (O_649,N_24776,N_20565);
or UO_650 (O_650,N_20846,N_23432);
nand UO_651 (O_651,N_21518,N_22870);
nor UO_652 (O_652,N_20911,N_22455);
nor UO_653 (O_653,N_23472,N_20262);
nor UO_654 (O_654,N_20389,N_24529);
nand UO_655 (O_655,N_20987,N_21094);
and UO_656 (O_656,N_22909,N_21153);
nor UO_657 (O_657,N_21683,N_21194);
and UO_658 (O_658,N_21745,N_23918);
nor UO_659 (O_659,N_24595,N_23402);
nor UO_660 (O_660,N_24218,N_21505);
and UO_661 (O_661,N_24091,N_23260);
and UO_662 (O_662,N_24614,N_24351);
nor UO_663 (O_663,N_22629,N_24597);
nor UO_664 (O_664,N_21718,N_22757);
nor UO_665 (O_665,N_23608,N_24406);
or UO_666 (O_666,N_21049,N_24000);
nor UO_667 (O_667,N_22726,N_21265);
nor UO_668 (O_668,N_23553,N_24157);
nand UO_669 (O_669,N_23355,N_23652);
nor UO_670 (O_670,N_20018,N_22293);
or UO_671 (O_671,N_21058,N_23959);
nor UO_672 (O_672,N_22792,N_21354);
and UO_673 (O_673,N_23940,N_23176);
or UO_674 (O_674,N_23643,N_23379);
or UO_675 (O_675,N_23528,N_20518);
nand UO_676 (O_676,N_20894,N_22992);
and UO_677 (O_677,N_22394,N_22608);
nor UO_678 (O_678,N_24117,N_20604);
xor UO_679 (O_679,N_21708,N_21738);
nand UO_680 (O_680,N_24894,N_21426);
nor UO_681 (O_681,N_23229,N_22438);
nor UO_682 (O_682,N_20746,N_22596);
or UO_683 (O_683,N_24099,N_22079);
and UO_684 (O_684,N_21230,N_24175);
nand UO_685 (O_685,N_20168,N_23255);
nor UO_686 (O_686,N_20727,N_23507);
nand UO_687 (O_687,N_23349,N_20141);
nand UO_688 (O_688,N_22205,N_21766);
nand UO_689 (O_689,N_22581,N_20646);
and UO_690 (O_690,N_21387,N_21089);
and UO_691 (O_691,N_22710,N_21612);
or UO_692 (O_692,N_22196,N_24772);
and UO_693 (O_693,N_21576,N_21315);
nor UO_694 (O_694,N_20441,N_24276);
nor UO_695 (O_695,N_23069,N_24533);
or UO_696 (O_696,N_22974,N_24663);
nand UO_697 (O_697,N_20234,N_21423);
nor UO_698 (O_698,N_24303,N_23725);
xor UO_699 (O_699,N_22946,N_20200);
xnor UO_700 (O_700,N_23011,N_24679);
or UO_701 (O_701,N_20562,N_23535);
and UO_702 (O_702,N_23113,N_20890);
nand UO_703 (O_703,N_20838,N_21389);
nand UO_704 (O_704,N_22691,N_24677);
or UO_705 (O_705,N_23979,N_24495);
or UO_706 (O_706,N_23749,N_22611);
nand UO_707 (O_707,N_24086,N_24913);
nor UO_708 (O_708,N_20228,N_24189);
or UO_709 (O_709,N_22947,N_21206);
nor UO_710 (O_710,N_23231,N_20127);
nor UO_711 (O_711,N_24582,N_24620);
nand UO_712 (O_712,N_24955,N_21609);
or UO_713 (O_713,N_24632,N_23315);
nand UO_714 (O_714,N_21276,N_23440);
nand UO_715 (O_715,N_22287,N_24490);
or UO_716 (O_716,N_21286,N_22110);
xnor UO_717 (O_717,N_21309,N_24163);
or UO_718 (O_718,N_20377,N_23581);
or UO_719 (O_719,N_22491,N_20773);
nand UO_720 (O_720,N_24915,N_23322);
and UO_721 (O_721,N_24552,N_20881);
nor UO_722 (O_722,N_20219,N_24051);
nor UO_723 (O_723,N_22822,N_23064);
nand UO_724 (O_724,N_21189,N_24711);
and UO_725 (O_725,N_23377,N_23806);
nand UO_726 (O_726,N_22990,N_21133);
or UO_727 (O_727,N_21808,N_24330);
nor UO_728 (O_728,N_22593,N_24499);
and UO_729 (O_729,N_23210,N_20858);
nor UO_730 (O_730,N_20645,N_22775);
and UO_731 (O_731,N_23448,N_23437);
nor UO_732 (O_732,N_22925,N_23299);
and UO_733 (O_733,N_22383,N_22697);
or UO_734 (O_734,N_23913,N_23621);
nor UO_735 (O_735,N_22347,N_23152);
and UO_736 (O_736,N_23318,N_24151);
and UO_737 (O_737,N_24319,N_21530);
or UO_738 (O_738,N_22565,N_24628);
nor UO_739 (O_739,N_20296,N_20529);
and UO_740 (O_740,N_22014,N_20830);
nand UO_741 (O_741,N_20902,N_22288);
nand UO_742 (O_742,N_21991,N_22772);
nand UO_743 (O_743,N_22746,N_24970);
nand UO_744 (O_744,N_24048,N_20350);
and UO_745 (O_745,N_21202,N_24818);
nand UO_746 (O_746,N_21026,N_21227);
nor UO_747 (O_747,N_20236,N_20067);
nand UO_748 (O_748,N_20170,N_23048);
nand UO_749 (O_749,N_22154,N_24835);
and UO_750 (O_750,N_20912,N_24416);
or UO_751 (O_751,N_20577,N_21800);
or UO_752 (O_752,N_23654,N_22136);
and UO_753 (O_753,N_23203,N_20033);
and UO_754 (O_754,N_24310,N_21252);
or UO_755 (O_755,N_20982,N_24900);
nand UO_756 (O_756,N_20437,N_24298);
and UO_757 (O_757,N_22027,N_23932);
and UO_758 (O_758,N_22500,N_20673);
nor UO_759 (O_759,N_22998,N_21030);
or UO_760 (O_760,N_20785,N_22417);
and UO_761 (O_761,N_20705,N_20405);
nor UO_762 (O_762,N_22690,N_22114);
nand UO_763 (O_763,N_22954,N_22388);
or UO_764 (O_764,N_21829,N_23906);
or UO_765 (O_765,N_22856,N_23296);
or UO_766 (O_766,N_24466,N_24394);
and UO_767 (O_767,N_24972,N_24436);
nor UO_768 (O_768,N_23846,N_23948);
nor UO_769 (O_769,N_21237,N_23313);
or UO_770 (O_770,N_20374,N_20295);
nor UO_771 (O_771,N_21330,N_20101);
nand UO_772 (O_772,N_24799,N_21020);
and UO_773 (O_773,N_24221,N_22197);
nor UO_774 (O_774,N_21729,N_23883);
and UO_775 (O_775,N_22763,N_23828);
or UO_776 (O_776,N_21682,N_22482);
nor UO_777 (O_777,N_22681,N_22937);
nand UO_778 (O_778,N_21215,N_21825);
nand UO_779 (O_779,N_21535,N_21507);
or UO_780 (O_780,N_22081,N_20692);
and UO_781 (O_781,N_24425,N_21603);
nor UO_782 (O_782,N_21629,N_20554);
nand UO_783 (O_783,N_24112,N_23520);
and UO_784 (O_784,N_21854,N_21318);
and UO_785 (O_785,N_24831,N_22382);
nor UO_786 (O_786,N_22038,N_20367);
xnor UO_787 (O_787,N_22420,N_23022);
nor UO_788 (O_788,N_22752,N_21540);
or UO_789 (O_789,N_22653,N_23545);
nand UO_790 (O_790,N_21788,N_21079);
nor UO_791 (O_791,N_23092,N_20208);
and UO_792 (O_792,N_21972,N_23519);
xor UO_793 (O_793,N_22353,N_21815);
and UO_794 (O_794,N_24566,N_20805);
nor UO_795 (O_795,N_24041,N_22860);
nor UO_796 (O_796,N_22434,N_23824);
nor UO_797 (O_797,N_22331,N_21099);
nor UO_798 (O_798,N_24721,N_24786);
and UO_799 (O_799,N_23098,N_20026);
or UO_800 (O_800,N_24477,N_23875);
xor UO_801 (O_801,N_24726,N_20179);
nand UO_802 (O_802,N_22116,N_24755);
and UO_803 (O_803,N_20420,N_22028);
nand UO_804 (O_804,N_22286,N_24917);
nor UO_805 (O_805,N_22264,N_22093);
or UO_806 (O_806,N_23335,N_23850);
and UO_807 (O_807,N_22433,N_21195);
nand UO_808 (O_808,N_20149,N_22876);
and UO_809 (O_809,N_22452,N_20556);
nand UO_810 (O_810,N_24265,N_23121);
and UO_811 (O_811,N_23930,N_22471);
nand UO_812 (O_812,N_22314,N_23386);
nor UO_813 (O_813,N_23625,N_21844);
or UO_814 (O_814,N_24736,N_21979);
nor UO_815 (O_815,N_21560,N_22403);
and UO_816 (O_816,N_24935,N_22186);
nor UO_817 (O_817,N_21047,N_23086);
nor UO_818 (O_818,N_24284,N_22048);
nor UO_819 (O_819,N_23793,N_24002);
or UO_820 (O_820,N_21990,N_20218);
and UO_821 (O_821,N_23339,N_21822);
nor UO_822 (O_822,N_24461,N_21488);
and UO_823 (O_823,N_23204,N_20793);
and UO_824 (O_824,N_24364,N_22828);
nand UO_825 (O_825,N_22612,N_22416);
or UO_826 (O_826,N_21785,N_22435);
nand UO_827 (O_827,N_23772,N_23655);
or UO_828 (O_828,N_20064,N_21698);
nor UO_829 (O_829,N_21031,N_24649);
and UO_830 (O_830,N_24936,N_22334);
nor UO_831 (O_831,N_24098,N_21482);
and UO_832 (O_832,N_20885,N_24670);
or UO_833 (O_833,N_22589,N_24660);
and UO_834 (O_834,N_21437,N_23984);
and UO_835 (O_835,N_20889,N_20162);
nand UO_836 (O_836,N_21977,N_24822);
nor UO_837 (O_837,N_24813,N_21469);
and UO_838 (O_838,N_23563,N_24074);
or UO_839 (O_839,N_22282,N_24879);
and UO_840 (O_840,N_20628,N_23744);
and UO_841 (O_841,N_23066,N_24798);
and UO_842 (O_842,N_24830,N_23372);
nand UO_843 (O_843,N_22639,N_24575);
or UO_844 (O_844,N_20935,N_23780);
xnor UO_845 (O_845,N_23050,N_23513);
nand UO_846 (O_846,N_20837,N_20528);
nand UO_847 (O_847,N_20625,N_24101);
xnor UO_848 (O_848,N_23320,N_24881);
or UO_849 (O_849,N_23821,N_23598);
nor UO_850 (O_850,N_23476,N_24949);
nor UO_851 (O_851,N_21581,N_24910);
nor UO_852 (O_852,N_23468,N_24844);
and UO_853 (O_853,N_21592,N_21842);
and UO_854 (O_854,N_24277,N_20620);
or UO_855 (O_855,N_21147,N_21628);
nand UO_856 (O_856,N_20136,N_23036);
xnor UO_857 (O_857,N_22874,N_20909);
nor UO_858 (O_858,N_23974,N_24907);
nand UO_859 (O_859,N_23186,N_20438);
and UO_860 (O_860,N_24613,N_20371);
nor UO_861 (O_861,N_20265,N_23365);
and UO_862 (O_862,N_21159,N_22178);
and UO_863 (O_863,N_22790,N_23891);
nor UO_864 (O_864,N_21415,N_20317);
or UO_865 (O_865,N_22229,N_22836);
or UO_866 (O_866,N_21388,N_20728);
nor UO_867 (O_867,N_24605,N_24519);
nand UO_868 (O_868,N_21256,N_24340);
and UO_869 (O_869,N_20572,N_21652);
nor UO_870 (O_870,N_21073,N_23831);
nand UO_871 (O_871,N_23860,N_20260);
or UO_872 (O_872,N_22446,N_24434);
nor UO_873 (O_873,N_20327,N_23874);
nand UO_874 (O_874,N_24055,N_21226);
and UO_875 (O_875,N_22945,N_20851);
nand UO_876 (O_876,N_24990,N_22412);
and UO_877 (O_877,N_21943,N_20948);
and UO_878 (O_878,N_22539,N_22736);
and UO_879 (O_879,N_20269,N_21355);
nor UO_880 (O_880,N_22126,N_22729);
or UO_881 (O_881,N_21995,N_21413);
nand UO_882 (O_882,N_20370,N_22506);
and UO_883 (O_883,N_21335,N_20781);
nor UO_884 (O_884,N_21063,N_21121);
or UO_885 (O_885,N_23433,N_22897);
xor UO_886 (O_886,N_20210,N_23760);
nor UO_887 (O_887,N_20762,N_23578);
or UO_888 (O_888,N_22928,N_24641);
nand UO_889 (O_889,N_24386,N_23408);
and UO_890 (O_890,N_23208,N_22664);
or UO_891 (O_891,N_21125,N_22002);
nor UO_892 (O_892,N_23863,N_24382);
or UO_893 (O_893,N_20915,N_20928);
and UO_894 (O_894,N_20969,N_22177);
nand UO_895 (O_895,N_20981,N_20297);
and UO_896 (O_896,N_21919,N_23222);
and UO_897 (O_897,N_22857,N_24282);
and UO_898 (O_898,N_20164,N_24701);
nand UO_899 (O_899,N_23958,N_20629);
and UO_900 (O_900,N_21462,N_23114);
xor UO_901 (O_901,N_21520,N_24888);
and UO_902 (O_902,N_20083,N_21564);
and UO_903 (O_903,N_22620,N_22361);
nand UO_904 (O_904,N_22767,N_23809);
nand UO_905 (O_905,N_23967,N_22001);
nor UO_906 (O_906,N_20415,N_23957);
nand UO_907 (O_907,N_23382,N_24790);
or UO_908 (O_908,N_21007,N_23936);
or UO_909 (O_909,N_24985,N_23515);
nand UO_910 (O_910,N_24875,N_20287);
or UO_911 (O_911,N_23750,N_22490);
nor UO_912 (O_912,N_23389,N_23560);
or UO_913 (O_913,N_23404,N_21885);
nand UO_914 (O_914,N_23164,N_22106);
and UO_915 (O_915,N_21145,N_23822);
or UO_916 (O_916,N_23024,N_24805);
or UO_917 (O_917,N_22548,N_21832);
and UO_918 (O_918,N_20081,N_24920);
nand UO_919 (O_919,N_23792,N_23317);
and UO_920 (O_920,N_22271,N_22101);
and UO_921 (O_921,N_23118,N_22935);
and UO_922 (O_922,N_21653,N_21103);
or UO_923 (O_923,N_20791,N_24872);
nand UO_924 (O_924,N_22062,N_21411);
or UO_925 (O_925,N_24304,N_20828);
nor UO_926 (O_926,N_23453,N_24025);
nand UO_927 (O_927,N_23189,N_23722);
or UO_928 (O_928,N_22583,N_21135);
nor UO_929 (O_929,N_22885,N_20601);
nor UO_930 (O_930,N_23949,N_24709);
nand UO_931 (O_931,N_24253,N_23084);
nor UO_932 (O_932,N_22380,N_24196);
and UO_933 (O_933,N_24992,N_22680);
and UO_934 (O_934,N_21454,N_21068);
and UO_935 (O_935,N_20654,N_24930);
or UO_936 (O_936,N_23823,N_24797);
or UO_937 (O_937,N_20036,N_21510);
nor UO_938 (O_938,N_20333,N_22886);
nor UO_939 (O_939,N_24186,N_23735);
nand UO_940 (O_940,N_23677,N_20561);
xor UO_941 (O_941,N_22097,N_21604);
nor UO_942 (O_942,N_21199,N_20801);
and UO_943 (O_943,N_24373,N_22225);
nor UO_944 (O_944,N_20541,N_22902);
nand UO_945 (O_945,N_24853,N_22892);
or UO_946 (O_946,N_23390,N_24496);
and UO_947 (O_947,N_23062,N_22823);
nand UO_948 (O_948,N_22413,N_21013);
nor UO_949 (O_949,N_20284,N_21283);
nand UO_950 (O_950,N_24654,N_20019);
nor UO_951 (O_951,N_20803,N_22463);
nand UO_952 (O_952,N_21184,N_23456);
or UO_953 (O_953,N_23767,N_20082);
and UO_954 (O_954,N_20907,N_23687);
nand UO_955 (O_955,N_22564,N_24749);
or UO_956 (O_956,N_21294,N_21177);
or UO_957 (O_957,N_24540,N_22755);
or UO_958 (O_958,N_21033,N_24285);
nor UO_959 (O_959,N_21374,N_22268);
or UO_960 (O_960,N_21321,N_22374);
and UO_961 (O_961,N_22502,N_21633);
or UO_962 (O_962,N_20670,N_22617);
nand UO_963 (O_963,N_22121,N_22161);
nor UO_964 (O_964,N_22071,N_20950);
and UO_965 (O_965,N_21361,N_23816);
and UO_966 (O_966,N_21247,N_22389);
and UO_967 (O_967,N_21463,N_24426);
nor UO_968 (O_968,N_21332,N_23167);
nand UO_969 (O_969,N_22901,N_23346);
nand UO_970 (O_970,N_22883,N_20247);
and UO_971 (O_971,N_21915,N_24738);
and UO_972 (O_972,N_22372,N_20868);
or UO_973 (O_973,N_20087,N_24856);
xor UO_974 (O_974,N_20434,N_24489);
nor UO_975 (O_975,N_23710,N_22398);
nor UO_976 (O_976,N_21574,N_23646);
nand UO_977 (O_977,N_22305,N_22688);
nand UO_978 (O_978,N_20006,N_23788);
nor UO_979 (O_979,N_24081,N_22013);
nand UO_980 (O_980,N_21608,N_22604);
nand UO_981 (O_981,N_21777,N_24622);
nand UO_982 (O_982,N_20843,N_20489);
or UO_983 (O_983,N_20636,N_22173);
and UO_984 (O_984,N_24752,N_24505);
nor UO_985 (O_985,N_22797,N_21623);
or UO_986 (O_986,N_23159,N_24686);
nor UO_987 (O_987,N_23227,N_21235);
and UO_988 (O_988,N_20455,N_22844);
nand UO_989 (O_989,N_24759,N_21464);
or UO_990 (O_990,N_21840,N_21053);
or UO_991 (O_991,N_21665,N_24683);
or UO_992 (O_992,N_20351,N_21451);
nand UO_993 (O_993,N_20227,N_22410);
nor UO_994 (O_994,N_23629,N_21360);
nor UO_995 (O_995,N_23422,N_21820);
nand UO_996 (O_996,N_24414,N_21830);
nand UO_997 (O_997,N_20488,N_23994);
nor UO_998 (O_998,N_23252,N_22207);
or UO_999 (O_999,N_23878,N_21759);
and UO_1000 (O_1000,N_24653,N_24816);
or UO_1001 (O_1001,N_22498,N_23465);
and UO_1002 (O_1002,N_21950,N_22322);
and UO_1003 (O_1003,N_22759,N_24026);
or UO_1004 (O_1004,N_21422,N_23494);
nor UO_1005 (O_1005,N_23516,N_21111);
nor UO_1006 (O_1006,N_20873,N_22310);
and UO_1007 (O_1007,N_24007,N_20242);
nor UO_1008 (O_1008,N_20924,N_24001);
or UO_1009 (O_1009,N_20155,N_24634);
nor UO_1010 (O_1010,N_21532,N_23522);
or UO_1011 (O_1011,N_24246,N_23199);
nand UO_1012 (O_1012,N_23672,N_23235);
or UO_1013 (O_1013,N_24314,N_23965);
nor UO_1014 (O_1014,N_23481,N_24825);
nand UO_1015 (O_1015,N_20194,N_20119);
or UO_1016 (O_1016,N_24892,N_20495);
and UO_1017 (O_1017,N_24692,N_22511);
xor UO_1018 (O_1018,N_20352,N_20041);
nand UO_1019 (O_1019,N_24328,N_21288);
nand UO_1020 (O_1020,N_21602,N_24596);
or UO_1021 (O_1021,N_24217,N_24446);
nor UO_1022 (O_1022,N_23148,N_22444);
and UO_1023 (O_1023,N_20624,N_24147);
and UO_1024 (O_1024,N_22472,N_20126);
nand UO_1025 (O_1025,N_22475,N_24693);
nor UO_1026 (O_1026,N_24453,N_20910);
or UO_1027 (O_1027,N_20118,N_22854);
nor UO_1028 (O_1028,N_22921,N_24417);
and UO_1029 (O_1029,N_21802,N_24361);
or UO_1030 (O_1030,N_23881,N_24424);
or UO_1031 (O_1031,N_20300,N_23137);
or UO_1032 (O_1032,N_24771,N_24155);
nand UO_1033 (O_1033,N_24667,N_23469);
nor UO_1034 (O_1034,N_24144,N_23196);
nor UO_1035 (O_1035,N_23397,N_23928);
nand UO_1036 (O_1036,N_21015,N_23471);
nand UO_1037 (O_1037,N_24758,N_24126);
and UO_1038 (O_1038,N_21586,N_20213);
and UO_1039 (O_1039,N_24069,N_24043);
nor UO_1040 (O_1040,N_20972,N_23909);
nand UO_1041 (O_1041,N_20021,N_21567);
and UO_1042 (O_1042,N_24441,N_24728);
or UO_1043 (O_1043,N_21322,N_24989);
or UO_1044 (O_1044,N_21257,N_22112);
nor UO_1045 (O_1045,N_23288,N_20484);
nor UO_1046 (O_1046,N_21566,N_21807);
nand UO_1047 (O_1047,N_24548,N_24779);
nor UO_1048 (O_1048,N_22991,N_22768);
or UO_1049 (O_1049,N_21363,N_23676);
or UO_1050 (O_1050,N_24430,N_24248);
and UO_1051 (O_1051,N_22292,N_22489);
or UO_1052 (O_1052,N_20515,N_22375);
and UO_1053 (O_1053,N_24231,N_23505);
nor UO_1054 (O_1054,N_21404,N_24669);
nor UO_1055 (O_1055,N_23551,N_21909);
xnor UO_1056 (O_1056,N_20157,N_20479);
nor UO_1057 (O_1057,N_23484,N_24576);
nor UO_1058 (O_1058,N_20304,N_23076);
nand UO_1059 (O_1059,N_22508,N_20025);
and UO_1060 (O_1060,N_22955,N_20305);
nor UO_1061 (O_1061,N_24741,N_24957);
or UO_1062 (O_1062,N_21826,N_23179);
nand UO_1063 (O_1063,N_21489,N_24778);
or UO_1064 (O_1064,N_24400,N_23815);
nand UO_1065 (O_1065,N_22250,N_21521);
nor UO_1066 (O_1066,N_21259,N_21476);
nand UO_1067 (O_1067,N_21955,N_22276);
or UO_1068 (O_1068,N_22346,N_20929);
and UO_1069 (O_1069,N_22656,N_20640);
nor UO_1070 (O_1070,N_24269,N_22887);
and UO_1071 (O_1071,N_24680,N_23192);
nor UO_1072 (O_1072,N_20778,N_23790);
and UO_1073 (O_1073,N_23704,N_21428);
xnor UO_1074 (O_1074,N_23620,N_23431);
and UO_1075 (O_1075,N_24932,N_20426);
and UO_1076 (O_1076,N_23213,N_23983);
or UO_1077 (O_1077,N_20896,N_20999);
nor UO_1078 (O_1078,N_24792,N_23104);
nor UO_1079 (O_1079,N_22219,N_24647);
and UO_1080 (O_1080,N_24652,N_24777);
nand UO_1081 (O_1081,N_21821,N_22499);
nand UO_1082 (O_1082,N_20499,N_23715);
and UO_1083 (O_1083,N_21083,N_21976);
nand UO_1084 (O_1084,N_21003,N_21468);
nor UO_1085 (O_1085,N_22551,N_23565);
nor UO_1086 (O_1086,N_20338,N_21861);
nand UO_1087 (O_1087,N_22043,N_21493);
nand UO_1088 (O_1088,N_24040,N_21916);
or UO_1089 (O_1089,N_23915,N_20172);
nand UO_1090 (O_1090,N_24702,N_20996);
nand UO_1091 (O_1091,N_23131,N_22644);
nor UO_1092 (O_1092,N_23593,N_22535);
and UO_1093 (O_1093,N_23867,N_21700);
nor UO_1094 (O_1094,N_23648,N_23882);
and UO_1095 (O_1095,N_21880,N_23720);
nand UO_1096 (O_1096,N_24706,N_23912);
or UO_1097 (O_1097,N_21443,N_23825);
nor UO_1098 (O_1098,N_21681,N_23003);
and UO_1099 (O_1099,N_23381,N_20075);
or UO_1100 (O_1100,N_20574,N_20402);
nand UO_1101 (O_1101,N_22632,N_22480);
nand UO_1102 (O_1102,N_24357,N_21105);
nand UO_1103 (O_1103,N_21701,N_21780);
or UO_1104 (O_1104,N_23571,N_23089);
and UO_1105 (O_1105,N_21646,N_23134);
and UO_1106 (O_1106,N_20211,N_24071);
and UO_1107 (O_1107,N_23435,N_21162);
and UO_1108 (O_1108,N_23171,N_20453);
nand UO_1109 (O_1109,N_20608,N_22942);
and UO_1110 (O_1110,N_21277,N_22012);
nand UO_1111 (O_1111,N_24945,N_24463);
and UO_1112 (O_1112,N_22522,N_24405);
nor UO_1113 (O_1113,N_22051,N_20482);
nor UO_1114 (O_1114,N_21706,N_23307);
or UO_1115 (O_1115,N_22972,N_21006);
nor UO_1116 (O_1116,N_23658,N_20827);
nor UO_1117 (O_1117,N_21219,N_23443);
nand UO_1118 (O_1118,N_24088,N_21393);
xor UO_1119 (O_1119,N_21492,N_21183);
and UO_1120 (O_1120,N_22407,N_20588);
xor UO_1121 (O_1121,N_20431,N_23849);
and UO_1122 (O_1122,N_23636,N_22210);
and UO_1123 (O_1123,N_20331,N_24812);
or UO_1124 (O_1124,N_22959,N_23043);
nor UO_1125 (O_1125,N_24858,N_22466);
or UO_1126 (O_1126,N_20571,N_23058);
and UO_1127 (O_1127,N_21925,N_24536);
xor UO_1128 (O_1128,N_24594,N_24399);
and UO_1129 (O_1129,N_23717,N_22135);
nor UO_1130 (O_1130,N_23223,N_23508);
nand UO_1131 (O_1131,N_24523,N_24448);
or UO_1132 (O_1132,N_24781,N_24077);
nor UO_1133 (O_1133,N_21365,N_22760);
nand UO_1134 (O_1134,N_22422,N_21155);
and UO_1135 (O_1135,N_20369,N_20163);
nor UO_1136 (O_1136,N_23020,N_23993);
or UO_1137 (O_1137,N_22842,N_23151);
nor UO_1138 (O_1138,N_22711,N_22037);
or UO_1139 (O_1139,N_21019,N_20992);
nand UO_1140 (O_1140,N_20330,N_23096);
nand UO_1141 (O_1141,N_20301,N_24336);
nand UO_1142 (O_1142,N_20185,N_23688);
nand UO_1143 (O_1143,N_24191,N_22321);
nor UO_1144 (O_1144,N_24938,N_24449);
nand UO_1145 (O_1145,N_20630,N_24854);
nand UO_1146 (O_1146,N_22158,N_20276);
or UO_1147 (O_1147,N_20031,N_20343);
and UO_1148 (O_1148,N_23428,N_24345);
and UO_1149 (O_1149,N_21001,N_23510);
nor UO_1150 (O_1150,N_21928,N_24500);
and UO_1151 (O_1151,N_23871,N_22931);
and UO_1152 (O_1152,N_20448,N_20575);
and UO_1153 (O_1153,N_20193,N_20855);
and UO_1154 (O_1154,N_24488,N_24087);
or UO_1155 (O_1155,N_21998,N_21983);
nand UO_1156 (O_1156,N_20783,N_23200);
or UO_1157 (O_1157,N_24349,N_21465);
nand UO_1158 (O_1158,N_23391,N_23207);
or UO_1159 (O_1159,N_22588,N_21320);
nand UO_1160 (O_1160,N_24642,N_21642);
and UO_1161 (O_1161,N_21253,N_20158);
nand UO_1162 (O_1162,N_21516,N_20411);
nor UO_1163 (O_1163,N_21297,N_21792);
and UO_1164 (O_1164,N_22080,N_23550);
and UO_1165 (O_1165,N_24610,N_20722);
or UO_1166 (O_1166,N_21684,N_21433);
nand UO_1167 (O_1167,N_24906,N_22465);
nor UO_1168 (O_1168,N_21525,N_21035);
or UO_1169 (O_1169,N_21945,N_24852);
nor UO_1170 (O_1170,N_22149,N_20156);
or UO_1171 (O_1171,N_24403,N_24584);
nor UO_1172 (O_1172,N_20196,N_24905);
and UO_1173 (O_1173,N_24763,N_21037);
nor UO_1174 (O_1174,N_20810,N_20416);
or UO_1175 (O_1175,N_22344,N_21559);
or UO_1176 (O_1176,N_20730,N_24944);
or UO_1177 (O_1177,N_22151,N_23245);
xor UO_1178 (O_1178,N_24233,N_20866);
nor UO_1179 (O_1179,N_21671,N_23794);
nand UO_1180 (O_1180,N_22285,N_22781);
nand UO_1181 (O_1181,N_22181,N_24116);
nor UO_1182 (O_1182,N_21027,N_21279);
or UO_1183 (O_1183,N_21717,N_20632);
nor UO_1184 (O_1184,N_22579,N_24094);
and UO_1185 (O_1185,N_22875,N_21267);
nand UO_1186 (O_1186,N_22852,N_23518);
nand UO_1187 (O_1187,N_21606,N_21353);
nand UO_1188 (O_1188,N_22543,N_23963);
and UO_1189 (O_1189,N_20145,N_23734);
or UO_1190 (O_1190,N_20129,N_20901);
nor UO_1191 (O_1191,N_23706,N_23108);
nand UO_1192 (O_1192,N_20603,N_21975);
and UO_1193 (O_1193,N_20570,N_23602);
nand UO_1194 (O_1194,N_22975,N_22788);
nor UO_1195 (O_1195,N_21207,N_24264);
nand UO_1196 (O_1196,N_20538,N_22061);
nor UO_1197 (O_1197,N_21920,N_21817);
nand UO_1198 (O_1198,N_22408,N_21176);
nor UO_1199 (O_1199,N_23248,N_23082);
or UO_1200 (O_1200,N_21298,N_22666);
or UO_1201 (O_1201,N_23532,N_24761);
or UO_1202 (O_1202,N_20697,N_21948);
nand UO_1203 (O_1203,N_23388,N_21014);
and UO_1204 (O_1204,N_21669,N_20906);
or UO_1205 (O_1205,N_20543,N_22926);
and UO_1206 (O_1206,N_22676,N_23759);
nor UO_1207 (O_1207,N_24586,N_23343);
nor UO_1208 (O_1208,N_23942,N_23536);
and UO_1209 (O_1209,N_23187,N_22609);
and UO_1210 (O_1210,N_23797,N_22049);
or UO_1211 (O_1211,N_20964,N_20849);
or UO_1212 (O_1212,N_21806,N_22754);
nor UO_1213 (O_1213,N_22748,N_21100);
or UO_1214 (O_1214,N_23665,N_23063);
and UO_1215 (O_1215,N_21098,N_21971);
or UO_1216 (O_1216,N_24174,N_20863);
and UO_1217 (O_1217,N_24291,N_22426);
nand UO_1218 (O_1218,N_22066,N_21078);
nor UO_1219 (O_1219,N_23190,N_21661);
xor UO_1220 (O_1220,N_24988,N_24598);
nand UO_1221 (O_1221,N_22141,N_21810);
nand UO_1222 (O_1222,N_24006,N_22004);
nand UO_1223 (O_1223,N_23072,N_22983);
nand UO_1224 (O_1224,N_20792,N_20794);
or UO_1225 (O_1225,N_24211,N_24766);
nor UO_1226 (O_1226,N_24593,N_23573);
or UO_1227 (O_1227,N_24199,N_23743);
nor UO_1228 (O_1228,N_24278,N_24398);
nor UO_1229 (O_1229,N_24608,N_22153);
or UO_1230 (O_1230,N_20053,N_21610);
nand UO_1231 (O_1231,N_22397,N_20811);
nand UO_1232 (O_1232,N_22727,N_24857);
nor UO_1233 (O_1233,N_23091,N_21050);
nand UO_1234 (O_1234,N_20221,N_20254);
nor UO_1235 (O_1235,N_24312,N_24411);
nor UO_1236 (O_1236,N_23552,N_22007);
or UO_1237 (O_1237,N_24503,N_21556);
nand UO_1238 (O_1238,N_24739,N_24659);
and UO_1239 (O_1239,N_20995,N_24313);
or UO_1240 (O_1240,N_22663,N_21923);
or UO_1241 (O_1241,N_22365,N_20845);
and UO_1242 (O_1242,N_20569,N_21689);
nor UO_1243 (O_1243,N_20335,N_21057);
nor UO_1244 (O_1244,N_23933,N_20057);
nand UO_1245 (O_1245,N_23273,N_24865);
nor UO_1246 (O_1246,N_21801,N_23195);
nor UO_1247 (O_1247,N_21599,N_20024);
or UO_1248 (O_1248,N_21675,N_21847);
nor UO_1249 (O_1249,N_24047,N_20887);
or UO_1250 (O_1250,N_20606,N_22970);
and UO_1251 (O_1251,N_22159,N_21539);
and UO_1252 (O_1252,N_24502,N_23575);
nor UO_1253 (O_1253,N_23059,N_20511);
and UO_1254 (O_1254,N_22515,N_21563);
nor UO_1255 (O_1255,N_22090,N_20623);
and UO_1256 (O_1256,N_21933,N_22359);
nor UO_1257 (O_1257,N_23728,N_24169);
nor UO_1258 (O_1258,N_20069,N_20015);
nand UO_1259 (O_1259,N_24180,N_22327);
xor UO_1260 (O_1260,N_23990,N_22484);
or UO_1261 (O_1261,N_21514,N_21839);
or UO_1262 (O_1262,N_21554,N_22850);
or UO_1263 (O_1263,N_23281,N_20695);
or UO_1264 (O_1264,N_24987,N_21625);
nor UO_1265 (O_1265,N_22770,N_22783);
and UO_1266 (O_1266,N_20725,N_20427);
nand UO_1267 (O_1267,N_24897,N_20853);
or UO_1268 (O_1268,N_20251,N_22793);
and UO_1269 (O_1269,N_20978,N_21205);
nand UO_1270 (O_1270,N_23712,N_24344);
and UO_1271 (O_1271,N_22211,N_24128);
or UO_1272 (O_1272,N_22999,N_24079);
nor UO_1273 (O_1273,N_20497,N_24842);
nand UO_1274 (O_1274,N_20813,N_22806);
or UO_1275 (O_1275,N_21978,N_22423);
or UO_1276 (O_1276,N_20310,N_22029);
or UO_1277 (O_1277,N_22336,N_21936);
nand UO_1278 (O_1278,N_22150,N_22030);
and UO_1279 (O_1279,N_20467,N_20379);
nand UO_1280 (O_1280,N_23721,N_23559);
nor UO_1281 (O_1281,N_20259,N_20956);
nor UO_1282 (O_1282,N_22837,N_20675);
nand UO_1283 (O_1283,N_21900,N_21954);
or UO_1284 (O_1284,N_23812,N_20454);
nor UO_1285 (O_1285,N_20442,N_20669);
nor UO_1286 (O_1286,N_23101,N_21141);
or UO_1287 (O_1287,N_22619,N_20917);
nand UO_1288 (O_1288,N_23077,N_20706);
or UO_1289 (O_1289,N_23606,N_22445);
nand UO_1290 (O_1290,N_23290,N_20223);
and UO_1291 (O_1291,N_24109,N_20496);
or UO_1292 (O_1292,N_20257,N_20797);
or UO_1293 (O_1293,N_22687,N_23413);
or UO_1294 (O_1294,N_21328,N_20253);
nand UO_1295 (O_1295,N_21182,N_21251);
nand UO_1296 (O_1296,N_23495,N_24541);
nor UO_1297 (O_1297,N_22228,N_20573);
nand UO_1298 (O_1298,N_24440,N_21084);
nor UO_1299 (O_1299,N_20621,N_23122);
nand UO_1300 (O_1300,N_23083,N_20862);
nand UO_1301 (O_1301,N_24141,N_23184);
xnor UO_1302 (O_1302,N_24032,N_21124);
or UO_1303 (O_1303,N_21485,N_23944);
nand UO_1304 (O_1304,N_23294,N_21266);
nor UO_1305 (O_1305,N_21997,N_20962);
and UO_1306 (O_1306,N_21130,N_23627);
nor UO_1307 (O_1307,N_23663,N_20112);
and UO_1308 (O_1308,N_21962,N_22723);
nor UO_1309 (O_1309,N_20120,N_20104);
or UO_1310 (O_1310,N_21110,N_20592);
or UO_1311 (O_1311,N_20716,N_22431);
nand UO_1312 (O_1312,N_22415,N_24639);
or UO_1313 (O_1313,N_24325,N_24720);
nor UO_1314 (O_1314,N_21852,N_21344);
nand UO_1315 (O_1315,N_20599,N_20590);
or UO_1316 (O_1316,N_22742,N_22758);
nor UO_1317 (O_1317,N_20751,N_20970);
or UO_1318 (O_1318,N_22390,N_20122);
nor UO_1319 (O_1319,N_23533,N_20462);
and UO_1320 (O_1320,N_24600,N_23403);
nor UO_1321 (O_1321,N_23110,N_22464);
or UO_1322 (O_1322,N_20412,N_20898);
and UO_1323 (O_1323,N_24306,N_23956);
nand UO_1324 (O_1324,N_21641,N_23885);
and UO_1325 (O_1325,N_20404,N_24555);
and UO_1326 (O_1326,N_21291,N_24532);
or UO_1327 (O_1327,N_20032,N_22459);
and UO_1328 (O_1328,N_23007,N_23899);
and UO_1329 (O_1329,N_22406,N_20061);
nand UO_1330 (O_1330,N_23701,N_22391);
nand UO_1331 (O_1331,N_24367,N_22198);
or UO_1332 (O_1332,N_20106,N_20355);
nand UO_1333 (O_1333,N_20059,N_24464);
and UO_1334 (O_1334,N_22923,N_24022);
and UO_1335 (O_1335,N_20050,N_22724);
and UO_1336 (O_1336,N_24690,N_22546);
and UO_1337 (O_1337,N_24363,N_22738);
xor UO_1338 (O_1338,N_20139,N_21771);
nand UO_1339 (O_1339,N_24229,N_23030);
or UO_1340 (O_1340,N_20226,N_21436);
nand UO_1341 (O_1341,N_21907,N_21262);
nor UO_1342 (O_1342,N_22371,N_21471);
nor UO_1343 (O_1343,N_24085,N_21570);
nor UO_1344 (O_1344,N_21143,N_22708);
or UO_1345 (O_1345,N_23364,N_21804);
or UO_1346 (O_1346,N_23051,N_21702);
and UO_1347 (O_1347,N_23093,N_22647);
nor UO_1348 (O_1348,N_22936,N_23300);
and UO_1349 (O_1349,N_22524,N_20517);
nand UO_1350 (O_1350,N_21834,N_20967);
nor UO_1351 (O_1351,N_20748,N_22052);
or UO_1352 (O_1352,N_23421,N_20744);
nand UO_1353 (O_1353,N_20177,N_20685);
and UO_1354 (O_1354,N_20419,N_21196);
or UO_1355 (O_1355,N_24037,N_20860);
nand UO_1356 (O_1356,N_21203,N_22213);
nand UO_1357 (O_1357,N_23981,N_20923);
nand UO_1358 (O_1358,N_23814,N_23283);
and UO_1359 (O_1359,N_22668,N_23732);
nor UO_1360 (O_1360,N_20003,N_22487);
nand UO_1361 (O_1361,N_21490,N_20189);
nor UO_1362 (O_1362,N_24480,N_21450);
and UO_1363 (O_1363,N_24062,N_21965);
xnor UO_1364 (O_1364,N_23181,N_23324);
and UO_1365 (O_1365,N_21406,N_24618);
nand UO_1366 (O_1366,N_23280,N_24301);
nor UO_1367 (O_1367,N_23193,N_20761);
nor UO_1368 (O_1368,N_20361,N_20820);
nand UO_1369 (O_1369,N_21417,N_23095);
nand UO_1370 (O_1370,N_23021,N_22297);
nand UO_1371 (O_1371,N_21660,N_23504);
nor UO_1372 (O_1372,N_24756,N_23779);
nor UO_1373 (O_1373,N_22232,N_23000);
nand UO_1374 (O_1374,N_22108,N_23466);
nor UO_1375 (O_1375,N_22922,N_21397);
or UO_1376 (O_1376,N_23987,N_24993);
nand UO_1377 (O_1377,N_20094,N_22094);
nor UO_1378 (O_1378,N_21583,N_22761);
nand UO_1379 (O_1379,N_23503,N_23525);
or UO_1380 (O_1380,N_24612,N_23703);
and UO_1381 (O_1381,N_21713,N_24409);
and UO_1382 (O_1382,N_24862,N_23425);
nand UO_1383 (O_1383,N_22819,N_23638);
nand UO_1384 (O_1384,N_21816,N_20508);
nand UO_1385 (O_1385,N_24966,N_20178);
nor UO_1386 (O_1386,N_22194,N_21378);
or UO_1387 (O_1387,N_20775,N_22827);
or UO_1388 (O_1388,N_22130,N_20372);
nand UO_1389 (O_1389,N_23895,N_20619);
and UO_1390 (O_1390,N_20474,N_22944);
nand UO_1391 (O_1391,N_22985,N_22803);
or UO_1392 (O_1392,N_20012,N_24125);
and UO_1393 (O_1393,N_24228,N_23709);
nor UO_1394 (O_1394,N_20760,N_23367);
and UO_1395 (O_1395,N_20456,N_21326);
nor UO_1396 (O_1396,N_23789,N_20647);
nor UO_1397 (O_1397,N_20913,N_22376);
or UO_1398 (O_1398,N_22275,N_24901);
nor UO_1399 (O_1399,N_24097,N_24827);
nor UO_1400 (O_1400,N_21961,N_24747);
or UO_1401 (O_1401,N_22669,N_20309);
nand UO_1402 (O_1402,N_20109,N_23502);
or UO_1403 (O_1403,N_20816,N_24980);
and UO_1404 (O_1404,N_22785,N_24615);
and UO_1405 (O_1405,N_20594,N_21452);
nor UO_1406 (O_1406,N_23907,N_20433);
and UO_1407 (O_1407,N_22549,N_20252);
nand UO_1408 (O_1408,N_22730,N_21712);
and UO_1409 (O_1409,N_20567,N_24289);
nor UO_1410 (O_1410,N_22623,N_22167);
nand UO_1411 (O_1411,N_21244,N_20076);
nor UO_1412 (O_1412,N_20279,N_20661);
nand UO_1413 (O_1413,N_20649,N_20658);
or UO_1414 (O_1414,N_23730,N_23955);
nand UO_1415 (O_1415,N_20446,N_20918);
nand UO_1416 (O_1416,N_24954,N_20990);
and UO_1417 (O_1417,N_22544,N_24996);
nand UO_1418 (O_1418,N_24635,N_24347);
nand UO_1419 (O_1419,N_20380,N_23617);
or UO_1420 (O_1420,N_24601,N_22501);
nand UO_1421 (O_1421,N_22516,N_24197);
and UO_1422 (O_1422,N_24359,N_24982);
or UO_1423 (O_1423,N_24100,N_24725);
and UO_1424 (O_1424,N_21412,N_20689);
and UO_1425 (O_1425,N_20821,N_20836);
nand UO_1426 (O_1426,N_23653,N_23001);
nand UO_1427 (O_1427,N_20366,N_21446);
nand UO_1428 (O_1428,N_23890,N_21994);
nand UO_1429 (O_1429,N_21009,N_23726);
nand UO_1430 (O_1430,N_20501,N_21934);
or UO_1431 (O_1431,N_20510,N_24962);
or UO_1432 (O_1432,N_23851,N_23387);
and UO_1433 (O_1433,N_24688,N_24481);
nor UO_1434 (O_1434,N_24378,N_24609);
nor UO_1435 (O_1435,N_22805,N_20921);
or UO_1436 (O_1436,N_22989,N_21734);
or UO_1437 (O_1437,N_23427,N_21091);
nand UO_1438 (O_1438,N_24019,N_22102);
nand UO_1439 (O_1439,N_23194,N_20652);
or UO_1440 (O_1440,N_23605,N_21358);
or UO_1441 (O_1441,N_22553,N_24787);
nand UO_1442 (O_1442,N_22457,N_21951);
and UO_1443 (O_1443,N_20274,N_21508);
and UO_1444 (O_1444,N_24588,N_22355);
xor UO_1445 (O_1445,N_21200,N_21197);
or UO_1446 (O_1446,N_23609,N_23046);
and UO_1447 (O_1447,N_21855,N_21410);
or UO_1448 (O_1448,N_23540,N_22369);
or UO_1449 (O_1449,N_24114,N_20191);
or UO_1450 (O_1450,N_20691,N_21024);
or UO_1451 (O_1451,N_21096,N_20318);
and UO_1452 (O_1452,N_22155,N_21228);
nand UO_1453 (O_1453,N_22986,N_22745);
nor UO_1454 (O_1454,N_21692,N_24780);
and UO_1455 (O_1455,N_21434,N_24623);
nor UO_1456 (O_1456,N_20768,N_24515);
nand UO_1457 (O_1457,N_22685,N_24845);
and UO_1458 (O_1458,N_22393,N_22962);
and UO_1459 (O_1459,N_20796,N_24978);
nand UO_1460 (O_1460,N_20130,N_22009);
or UO_1461 (O_1461,N_22386,N_23124);
or UO_1462 (O_1462,N_22083,N_23847);
nor UO_1463 (O_1463,N_23359,N_22184);
nor UO_1464 (O_1464,N_20190,N_20953);
or UO_1465 (O_1465,N_20358,N_20273);
and UO_1466 (O_1466,N_22399,N_21192);
and UO_1467 (O_1467,N_20266,N_22086);
and UO_1468 (O_1468,N_20250,N_22267);
or UO_1469 (O_1469,N_20916,N_23107);
nor UO_1470 (O_1470,N_23384,N_21600);
and UO_1471 (O_1471,N_21819,N_21770);
or UO_1472 (O_1472,N_20469,N_22960);
or UO_1473 (O_1473,N_22719,N_22801);
nand UO_1474 (O_1474,N_20154,N_24323);
and UO_1475 (O_1475,N_22621,N_22692);
nand UO_1476 (O_1476,N_24638,N_23693);
or UO_1477 (O_1477,N_20766,N_24560);
nor UO_1478 (O_1478,N_21693,N_23396);
nand UO_1479 (O_1479,N_24643,N_21917);
nor UO_1480 (O_1480,N_21587,N_23827);
nor UO_1481 (O_1481,N_23309,N_21241);
nand UO_1482 (O_1482,N_24524,N_22782);
and UO_1483 (O_1483,N_21239,N_20357);
nor UO_1484 (O_1484,N_20893,N_22260);
and UO_1485 (O_1485,N_20583,N_20615);
nand UO_1486 (O_1486,N_22645,N_22440);
nor UO_1487 (O_1487,N_24733,N_20150);
nor UO_1488 (O_1488,N_24102,N_21062);
nand UO_1489 (O_1489,N_20410,N_22820);
nand UO_1490 (O_1490,N_23015,N_22180);
nor UO_1491 (O_1491,N_20114,N_23380);
or UO_1492 (O_1492,N_23618,N_23901);
nor UO_1493 (O_1493,N_21913,N_23412);
or UO_1494 (O_1494,N_20137,N_24286);
or UO_1495 (O_1495,N_23784,N_24817);
or UO_1496 (O_1496,N_20983,N_23099);
and UO_1497 (O_1497,N_24005,N_23325);
nor UO_1498 (O_1498,N_24864,N_22461);
and UO_1499 (O_1499,N_22572,N_20207);
and UO_1500 (O_1500,N_20737,N_22714);
nand UO_1501 (O_1501,N_20976,N_22363);
or UO_1502 (O_1502,N_23498,N_20831);
nor UO_1503 (O_1503,N_23736,N_23370);
nor UO_1504 (O_1504,N_21051,N_23242);
nor UO_1505 (O_1505,N_24748,N_23656);
or UO_1506 (O_1506,N_24902,N_21170);
or UO_1507 (O_1507,N_22098,N_24413);
or UO_1508 (O_1508,N_21487,N_20861);
and UO_1509 (O_1509,N_20693,N_20724);
nor UO_1510 (O_1510,N_22047,N_20527);
or UO_1511 (O_1511,N_24924,N_24808);
nand UO_1512 (O_1512,N_22847,N_21442);
nand UO_1513 (O_1513,N_24380,N_22060);
nand UO_1514 (O_1514,N_21240,N_22809);
or UO_1515 (O_1515,N_21427,N_23888);
xor UO_1516 (O_1516,N_22224,N_23637);
and UO_1517 (O_1517,N_24899,N_23138);
nor UO_1518 (O_1518,N_23526,N_24849);
or UO_1519 (O_1519,N_22753,N_20365);
and UO_1520 (O_1520,N_21761,N_21480);
nor UO_1521 (O_1521,N_24219,N_22884);
nand UO_1522 (O_1522,N_24965,N_21999);
or UO_1523 (O_1523,N_21506,N_20264);
or UO_1524 (O_1524,N_22342,N_21626);
nand UO_1525 (O_1525,N_22900,N_24828);
and UO_1526 (O_1526,N_20936,N_22077);
and UO_1527 (O_1527,N_24008,N_20052);
nor UO_1528 (O_1528,N_22615,N_21699);
nor UO_1529 (O_1529,N_21743,N_23305);
and UO_1530 (O_1530,N_20825,N_22414);
nor UO_1531 (O_1531,N_23442,N_20183);
nor UO_1532 (O_1532,N_22932,N_20217);
and UO_1533 (O_1533,N_20258,N_20663);
nand UO_1534 (O_1534,N_20079,N_22981);
xnor UO_1535 (O_1535,N_20822,N_23506);
nand UO_1536 (O_1536,N_22354,N_22831);
or UO_1537 (O_1537,N_21178,N_24024);
xor UO_1538 (O_1538,N_23670,N_20871);
nand UO_1539 (O_1539,N_21034,N_22815);
nand UO_1540 (O_1540,N_22095,N_21760);
nor UO_1541 (O_1541,N_21762,N_20235);
nand UO_1542 (O_1542,N_22995,N_22563);
nand UO_1543 (O_1543,N_24089,N_24860);
nor UO_1544 (O_1544,N_21113,N_20391);
nand UO_1545 (O_1545,N_24893,N_24129);
or UO_1546 (O_1546,N_21254,N_24621);
or UO_1547 (O_1547,N_22582,N_20378);
nor UO_1548 (O_1548,N_20492,N_20099);
and UO_1549 (O_1549,N_22769,N_20951);
nor UO_1550 (O_1550,N_21479,N_20030);
nand UO_1551 (O_1551,N_20919,N_20618);
nand UO_1552 (O_1552,N_20884,N_22206);
nor UO_1553 (O_1553,N_23991,N_22113);
nand UO_1554 (O_1554,N_22295,N_24707);
nor UO_1555 (O_1555,N_23628,N_23241);
or UO_1556 (O_1556,N_23954,N_20579);
or UO_1557 (O_1557,N_24050,N_24133);
xnor UO_1558 (O_1558,N_24571,N_22033);
and UO_1559 (O_1559,N_20360,N_24307);
or UO_1560 (O_1560,N_23155,N_22053);
nor UO_1561 (O_1561,N_23857,N_20187);
and UO_1562 (O_1562,N_21118,N_23633);
or UO_1563 (O_1563,N_21889,N_22290);
nor UO_1564 (O_1564,N_24497,N_22993);
or UO_1565 (O_1565,N_24012,N_20383);
and UO_1566 (O_1566,N_23060,N_23119);
and UO_1567 (O_1567,N_24388,N_24578);
xor UO_1568 (O_1568,N_23214,N_24030);
or UO_1569 (O_1569,N_23198,N_24366);
xor UO_1570 (O_1570,N_23594,N_22050);
nor UO_1571 (O_1571,N_23569,N_23682);
nor UO_1572 (O_1572,N_24986,N_20151);
or UO_1573 (O_1573,N_21299,N_23278);
nand UO_1574 (O_1574,N_24861,N_20758);
and UO_1575 (O_1575,N_23705,N_21863);
and UO_1576 (O_1576,N_20824,N_21704);
nand UO_1577 (O_1577,N_21772,N_22216);
nor UO_1578 (O_1578,N_22220,N_23270);
nor UO_1579 (O_1579,N_23880,N_24335);
and UO_1580 (O_1580,N_22392,N_24565);
nand UO_1581 (O_1581,N_22045,N_21445);
nor UO_1582 (O_1582,N_20413,N_24459);
and UO_1583 (O_1583,N_24941,N_23978);
nor UO_1584 (O_1584,N_21515,N_21768);
and UO_1585 (O_1585,N_22910,N_24457);
nand UO_1586 (O_1586,N_22679,N_20581);
nor UO_1587 (O_1587,N_24053,N_20182);
nand UO_1588 (O_1588,N_21687,N_20542);
or UO_1589 (O_1589,N_21168,N_23247);
nand UO_1590 (O_1590,N_21986,N_22091);
or UO_1591 (O_1591,N_20613,N_21753);
nand UO_1592 (O_1592,N_21477,N_21077);
nor UO_1593 (O_1593,N_20071,N_22956);
and UO_1594 (O_1594,N_20922,N_20774);
and UO_1595 (O_1595,N_23939,N_22927);
nand UO_1596 (O_1596,N_20255,N_20507);
nor UO_1597 (O_1597,N_22536,N_24689);
nand UO_1598 (O_1598,N_21129,N_20481);
or UO_1599 (O_1599,N_22362,N_23492);
and UO_1600 (O_1600,N_24869,N_23925);
nor UO_1601 (O_1601,N_21677,N_24833);
nor UO_1602 (O_1602,N_23624,N_20639);
or UO_1603 (O_1603,N_22169,N_20035);
or UO_1604 (O_1604,N_23240,N_23898);
or UO_1605 (O_1605,N_20678,N_22654);
or UO_1606 (O_1606,N_23669,N_23345);
and UO_1607 (O_1607,N_24836,N_20817);
nand UO_1608 (O_1608,N_20612,N_20332);
xnor UO_1609 (O_1609,N_21658,N_20707);
nor UO_1610 (O_1610,N_21107,N_21497);
nand UO_1611 (O_1611,N_20949,N_23049);
nand UO_1612 (O_1612,N_24762,N_23681);
nand UO_1613 (O_1613,N_24558,N_21966);
or UO_1614 (O_1614,N_24554,N_21229);
and UO_1615 (O_1615,N_24034,N_23539);
nor UO_1616 (O_1616,N_22214,N_24550);
or UO_1617 (O_1617,N_20733,N_21087);
and UO_1618 (O_1618,N_22706,N_20809);
and UO_1619 (O_1619,N_23600,N_23071);
nor UO_1620 (O_1620,N_24746,N_23897);
nand UO_1621 (O_1621,N_24934,N_23097);
or UO_1622 (O_1622,N_24912,N_21382);
or UO_1623 (O_1623,N_24656,N_22405);
nand UO_1624 (O_1624,N_22899,N_24535);
and UO_1625 (O_1625,N_21261,N_22367);
and UO_1626 (O_1626,N_23464,N_20329);
nand UO_1627 (O_1627,N_22238,N_22675);
nand UO_1628 (O_1628,N_24254,N_23795);
or UO_1629 (O_1629,N_20202,N_23251);
and UO_1630 (O_1630,N_23699,N_23657);
or UO_1631 (O_1631,N_23554,N_23451);
or UO_1632 (O_1632,N_21946,N_21064);
nand UO_1633 (O_1633,N_22963,N_22299);
or UO_1634 (O_1634,N_22103,N_21316);
nand UO_1635 (O_1635,N_22191,N_21211);
and UO_1636 (O_1636,N_20763,N_24198);
nand UO_1637 (O_1637,N_22064,N_21927);
and UO_1638 (O_1638,N_22821,N_20153);
nand UO_1639 (O_1639,N_20165,N_24890);
or UO_1640 (O_1640,N_22085,N_20334);
nand UO_1641 (O_1641,N_21377,N_20600);
nand UO_1642 (O_1642,N_22140,N_23989);
and UO_1643 (O_1643,N_20086,N_21043);
and UO_1644 (O_1644,N_21638,N_23572);
nor UO_1645 (O_1645,N_24095,N_22634);
nor UO_1646 (O_1646,N_20680,N_21250);
or UO_1647 (O_1647,N_20784,N_24090);
and UO_1648 (O_1648,N_24479,N_23191);
nor UO_1649 (O_1649,N_22907,N_22503);
nand UO_1650 (O_1650,N_20144,N_22642);
or UO_1651 (O_1651,N_20124,N_22943);
xor UO_1652 (O_1652,N_20930,N_21150);
nand UO_1653 (O_1653,N_21348,N_20029);
or UO_1654 (O_1654,N_24923,N_22556);
and UO_1655 (O_1655,N_20326,N_21095);
nor UO_1656 (O_1656,N_24106,N_22764);
or UO_1657 (O_1657,N_21385,N_21911);
or UO_1658 (O_1658,N_24537,N_22453);
and UO_1659 (O_1659,N_23068,N_21794);
nand UO_1660 (O_1660,N_22192,N_23361);
nor UO_1661 (O_1661,N_22657,N_22677);
and UO_1662 (O_1662,N_20043,N_21432);
or UO_1663 (O_1663,N_23582,N_20337);
or UO_1664 (O_1664,N_21831,N_24337);
nand UO_1665 (O_1665,N_22996,N_23174);
nor UO_1666 (O_1666,N_21767,N_20315);
nor UO_1667 (O_1667,N_21526,N_24587);
nor UO_1668 (O_1668,N_23004,N_20249);
and UO_1669 (O_1669,N_22915,N_20985);
nor UO_1670 (O_1670,N_24334,N_20037);
or UO_1671 (O_1671,N_23976,N_23859);
nand UO_1672 (O_1672,N_22031,N_21685);
and UO_1673 (O_1673,N_24057,N_23708);
and UO_1674 (O_1674,N_21589,N_23547);
and UO_1675 (O_1675,N_21370,N_21369);
xnor UO_1676 (O_1676,N_22478,N_20285);
and UO_1677 (O_1677,N_22168,N_20115);
and UO_1678 (O_1678,N_21879,N_21891);
and UO_1679 (O_1679,N_24017,N_23766);
and UO_1680 (O_1680,N_22204,N_24563);
nor UO_1681 (O_1681,N_20390,N_24815);
nor UO_1682 (O_1682,N_24300,N_23263);
and UO_1683 (O_1683,N_23564,N_23128);
nor UO_1684 (O_1684,N_23163,N_20239);
and UO_1685 (O_1685,N_22718,N_24432);
or UO_1686 (O_1686,N_20500,N_23444);
xor UO_1687 (O_1687,N_24220,N_22794);
or UO_1688 (O_1688,N_24564,N_23765);
or UO_1689 (O_1689,N_24765,N_22289);
and UO_1690 (O_1690,N_21384,N_24714);
nand UO_1691 (O_1691,N_22370,N_20641);
nand UO_1692 (O_1692,N_22917,N_20732);
or UO_1693 (O_1693,N_23591,N_20904);
or UO_1694 (O_1694,N_21289,N_23884);
and UO_1695 (O_1695,N_22460,N_23358);
or UO_1696 (O_1696,N_24998,N_20991);
and UO_1697 (O_1697,N_23920,N_24009);
and UO_1698 (O_1698,N_24574,N_24841);
nand UO_1699 (O_1699,N_24850,N_22523);
nor UO_1700 (O_1700,N_20116,N_23960);
xor UO_1701 (O_1701,N_21887,N_24393);
or UO_1702 (O_1702,N_21922,N_20450);
nor UO_1703 (O_1703,N_24569,N_23426);
and UO_1704 (O_1704,N_24401,N_22226);
or UO_1705 (O_1705,N_20347,N_24263);
or UO_1706 (O_1706,N_24768,N_22234);
nand UO_1707 (O_1707,N_24170,N_23306);
or UO_1708 (O_1708,N_20568,N_21455);
nor UO_1709 (O_1709,N_24518,N_21017);
nor UO_1710 (O_1710,N_23042,N_20443);
nand UO_1711 (O_1711,N_20311,N_24895);
or UO_1712 (O_1712,N_22303,N_24270);
or UO_1713 (O_1713,N_23724,N_23632);
or UO_1714 (O_1714,N_20616,N_23112);
or UO_1715 (O_1715,N_20353,N_24092);
and UO_1716 (O_1716,N_22889,N_21090);
nor UO_1717 (O_1717,N_21577,N_22189);
or UO_1718 (O_1718,N_21379,N_24156);
and UO_1719 (O_1719,N_23631,N_23642);
or UO_1720 (O_1720,N_21895,N_23029);
nand UO_1721 (O_1721,N_21824,N_22483);
nor UO_1722 (O_1722,N_21597,N_23988);
and UO_1723 (O_1723,N_23053,N_23462);
or UO_1724 (O_1724,N_20444,N_23250);
and UO_1725 (O_1725,N_22425,N_23033);
nor UO_1726 (O_1726,N_21122,N_23172);
and UO_1727 (O_1727,N_22527,N_22576);
nor UO_1728 (O_1728,N_24341,N_21246);
and UO_1729 (O_1729,N_20212,N_22263);
nand UO_1730 (O_1730,N_21324,N_20268);
nor UO_1731 (O_1731,N_22245,N_21204);
nand UO_1732 (O_1732,N_23301,N_24370);
and UO_1733 (O_1733,N_24568,N_23394);
xor UO_1734 (O_1734,N_21345,N_21952);
nor UO_1735 (O_1735,N_21870,N_24528);
or UO_1736 (O_1736,N_20872,N_22594);
and UO_1737 (O_1737,N_24487,N_21783);
nand UO_1738 (O_1738,N_22817,N_23922);
nor UO_1739 (O_1739,N_23027,N_22087);
and UO_1740 (O_1740,N_24664,N_21619);
nand UO_1741 (O_1741,N_23887,N_22240);
nor UO_1742 (O_1742,N_23892,N_21782);
nand UO_1743 (O_1743,N_23864,N_20524);
and UO_1744 (O_1744,N_20425,N_23845);
nand UO_1745 (O_1745,N_24737,N_20147);
or UO_1746 (O_1746,N_24320,N_22439);
or UO_1747 (O_1747,N_24943,N_21643);
and UO_1748 (O_1748,N_20808,N_20320);
or UO_1749 (O_1749,N_21942,N_22470);
nand UO_1750 (O_1750,N_21552,N_22971);
or UO_1751 (O_1751,N_20933,N_20439);
nand UO_1752 (O_1752,N_24940,N_24428);
nand UO_1753 (O_1753,N_23056,N_20963);
nor UO_1754 (O_1754,N_22924,N_24685);
or UO_1755 (O_1755,N_23333,N_24699);
and UO_1756 (O_1756,N_20316,N_20323);
nor UO_1757 (O_1757,N_22203,N_24194);
nor UO_1758 (O_1758,N_23855,N_22179);
and UO_1759 (O_1759,N_22586,N_20092);
and UO_1760 (O_1760,N_24111,N_23178);
nor UO_1761 (O_1761,N_24800,N_24309);
and UO_1762 (O_1762,N_24456,N_24158);
xor UO_1763 (O_1763,N_20662,N_22605);
nand UO_1764 (O_1764,N_20294,N_21558);
nand UO_1765 (O_1765,N_21499,N_22235);
nand UO_1766 (O_1766,N_24205,N_24105);
nor UO_1767 (O_1767,N_20054,N_23647);
nor UO_1768 (O_1768,N_23253,N_24847);
or UO_1769 (O_1769,N_21383,N_23512);
nand UO_1770 (O_1770,N_20980,N_22257);
nor UO_1771 (O_1771,N_20055,N_22222);
nor UO_1772 (O_1772,N_24483,N_21790);
nor UO_1773 (O_1773,N_22162,N_21352);
xor UO_1774 (O_1774,N_24775,N_20719);
or UO_1775 (O_1775,N_23399,N_24392);
nand UO_1776 (O_1776,N_21430,N_24251);
and UO_1777 (O_1777,N_21419,N_24138);
nor UO_1778 (O_1778,N_20940,N_24455);
or UO_1779 (O_1779,N_23038,N_20422);
nand UO_1780 (O_1780,N_20965,N_20905);
or UO_1781 (O_1781,N_21052,N_24376);
nand UO_1782 (O_1782,N_21511,N_20199);
or UO_1783 (O_1783,N_24458,N_22637);
or UO_1784 (O_1784,N_21740,N_21992);
nand UO_1785 (O_1785,N_22652,N_24377);
or UO_1786 (O_1786,N_22510,N_21989);
and UO_1787 (O_1787,N_24327,N_22731);
nand UO_1788 (O_1788,N_22911,N_20708);
nor UO_1789 (O_1789,N_24120,N_20017);
nand UO_1790 (O_1790,N_20879,N_21797);
or UO_1791 (O_1791,N_22529,N_20105);
and UO_1792 (O_1792,N_24195,N_22447);
or UO_1793 (O_1793,N_21329,N_22988);
xor UO_1794 (O_1794,N_21528,N_21672);
nand UO_1795 (O_1795,N_23755,N_23371);
or UO_1796 (O_1796,N_22242,N_22739);
nand UO_1797 (O_1797,N_23079,N_20346);
or UO_1798 (O_1798,N_23596,N_22712);
or UO_1799 (O_1799,N_21545,N_23352);
and UO_1800 (O_1800,N_24223,N_20850);
and UO_1801 (O_1801,N_20943,N_23768);
or UO_1802 (O_1802,N_23924,N_21601);
nand UO_1803 (O_1803,N_21814,N_20545);
nand UO_1804 (O_1804,N_24208,N_22266);
or UO_1805 (O_1805,N_24402,N_21040);
nor UO_1806 (O_1806,N_23409,N_21588);
nor UO_1807 (O_1807,N_21703,N_22630);
nand UO_1808 (O_1808,N_22477,N_22577);
and UO_1809 (O_1809,N_20298,N_20229);
nor UO_1810 (O_1810,N_22744,N_23968);
and UO_1811 (O_1811,N_21562,N_21886);
nor UO_1812 (O_1812,N_24903,N_23216);
nor UO_1813 (O_1813,N_20648,N_22728);
or UO_1814 (O_1814,N_23538,N_21630);
or UO_1815 (O_1815,N_24636,N_24339);
nor UO_1816 (O_1816,N_20841,N_20749);
nand UO_1817 (O_1817,N_23017,N_21114);
or UO_1818 (O_1818,N_22318,N_20657);
nand UO_1819 (O_1819,N_20564,N_20532);
and UO_1820 (O_1820,N_21418,N_21301);
nand UO_1821 (O_1821,N_20815,N_22665);
nor UO_1822 (O_1822,N_21904,N_21654);
and UO_1823 (O_1823,N_21336,N_23286);
nand UO_1824 (O_1824,N_22735,N_20585);
nor UO_1825 (O_1825,N_21117,N_23803);
nand UO_1826 (O_1826,N_24261,N_20842);
nor UO_1827 (O_1827,N_24333,N_24358);
nor UO_1828 (O_1828,N_22951,N_22122);
or UO_1829 (O_1829,N_24465,N_24255);
nand UO_1830 (O_1830,N_23293,N_20735);
nand UO_1831 (O_1831,N_20607,N_21306);
nand UO_1832 (O_1832,N_21594,N_24350);
and UO_1833 (O_1833,N_22247,N_23258);
nor UO_1834 (O_1834,N_23304,N_21884);
nor UO_1835 (O_1835,N_21985,N_24127);
xor UO_1836 (O_1836,N_21029,N_21691);
or UO_1837 (O_1837,N_23613,N_20856);
or UO_1838 (O_1838,N_20550,N_22032);
nand UO_1839 (O_1839,N_22137,N_22631);
or UO_1840 (O_1840,N_20563,N_24820);
and UO_1841 (O_1841,N_22350,N_21496);
or UO_1842 (O_1842,N_22743,N_21680);
nor UO_1843 (O_1843,N_21371,N_21314);
nor UO_1844 (O_1844,N_20014,N_21996);
nand UO_1845 (O_1845,N_20010,N_20237);
or UO_1846 (O_1846,N_24338,N_22313);
nor UO_1847 (O_1847,N_20513,N_20098);
or UO_1848 (O_1848,N_20134,N_21823);
nor UO_1849 (O_1849,N_21074,N_24724);
nor UO_1850 (O_1850,N_20891,N_23686);
or UO_1851 (O_1851,N_23626,N_23577);
nor UO_1852 (O_1852,N_23354,N_21963);
nand UO_1853 (O_1853,N_20428,N_24104);
nand UO_1854 (O_1854,N_21964,N_23392);
and UO_1855 (O_1855,N_23941,N_20280);
nor UO_1856 (O_1856,N_24371,N_22859);
nor UO_1857 (O_1857,N_23711,N_22829);
or UO_1858 (O_1858,N_23491,N_21778);
and UO_1859 (O_1859,N_24110,N_22046);
nor UO_1860 (O_1860,N_21843,N_23487);
and UO_1861 (O_1861,N_24929,N_21312);
nor UO_1862 (O_1862,N_21435,N_22320);
nor UO_1863 (O_1863,N_24801,N_23747);
nor UO_1864 (O_1864,N_22807,N_22567);
nand UO_1865 (O_1865,N_23819,N_23423);
nand UO_1866 (O_1866,N_23651,N_20181);
nor UO_1867 (O_1867,N_22134,N_21061);
and UO_1868 (O_1868,N_21474,N_22454);
or UO_1869 (O_1869,N_23180,N_24004);
or UO_1870 (O_1870,N_23457,N_20870);
nor UO_1871 (O_1871,N_24531,N_21152);
or UO_1872 (O_1872,N_21167,N_23634);
nand UO_1873 (O_1873,N_20938,N_23517);
and UO_1874 (O_1874,N_20672,N_20204);
nand UO_1875 (O_1875,N_24066,N_24137);
or UO_1876 (O_1876,N_21042,N_21231);
nand UO_1877 (O_1877,N_21967,N_21538);
or UO_1878 (O_1878,N_23002,N_22591);
or UO_1879 (O_1879,N_20721,N_21679);
nand UO_1880 (O_1880,N_22722,N_20677);
and UO_1881 (O_1881,N_22696,N_22251);
and UO_1882 (O_1882,N_21859,N_22280);
nand UO_1883 (O_1883,N_20039,N_20664);
or UO_1884 (O_1884,N_24509,N_23225);
nand UO_1885 (O_1885,N_22040,N_22124);
nor UO_1886 (O_1886,N_20375,N_24951);
and UO_1887 (O_1887,N_24871,N_23224);
nand UO_1888 (O_1888,N_21958,N_23054);
or UO_1889 (O_1889,N_21142,N_22542);
and UO_1890 (O_1890,N_22255,N_21495);
nand UO_1891 (O_1891,N_24750,N_22890);
or UO_1892 (O_1892,N_21614,N_24580);
and UO_1893 (O_1893,N_21296,N_21359);
nor UO_1894 (O_1894,N_22737,N_22929);
nor UO_1895 (O_1895,N_21549,N_20660);
nor UO_1896 (O_1896,N_23401,N_22908);
or UO_1897 (O_1897,N_20807,N_23684);
nand UO_1898 (O_1898,N_20582,N_22341);
and UO_1899 (O_1899,N_24318,N_21409);
or UO_1900 (O_1900,N_20578,N_23870);
nand UO_1901 (O_1901,N_20638,N_22777);
nand UO_1902 (O_1902,N_20753,N_20313);
or UO_1903 (O_1903,N_21221,N_21503);
and UO_1904 (O_1904,N_22063,N_20430);
or UO_1905 (O_1905,N_24134,N_22882);
or UO_1906 (O_1906,N_22176,N_21067);
nor UO_1907 (O_1907,N_24926,N_24769);
xnor UO_1908 (O_1908,N_21439,N_22713);
nor UO_1909 (O_1909,N_22430,N_21088);
or UO_1910 (O_1910,N_23169,N_22704);
and UO_1911 (O_1911,N_22934,N_21639);
nand UO_1912 (O_1912,N_22109,N_20847);
or UO_1913 (O_1913,N_24234,N_22366);
and UO_1914 (O_1914,N_22018,N_23450);
or UO_1915 (O_1915,N_21136,N_22237);
and UO_1916 (O_1916,N_22830,N_23405);
and UO_1917 (O_1917,N_23165,N_23023);
nand UO_1918 (O_1918,N_21127,N_24355);
and UO_1919 (O_1919,N_21104,N_24039);
and UO_1920 (O_1920,N_20016,N_21340);
nand UO_1921 (O_1921,N_23838,N_21865);
and UO_1922 (O_1922,N_24592,N_21696);
nor UO_1923 (O_1923,N_20072,N_21635);
nand UO_1924 (O_1924,N_22913,N_22146);
xor UO_1925 (O_1925,N_23914,N_24553);
or UO_1926 (O_1926,N_22218,N_23872);
nand UO_1927 (O_1927,N_24305,N_20899);
nand UO_1928 (O_1928,N_22894,N_20356);
nand UO_1929 (O_1929,N_24676,N_21541);
xor UO_1930 (O_1930,N_23524,N_24802);
and UO_1931 (O_1931,N_20731,N_23751);
and UO_1932 (O_1932,N_22966,N_24646);
and UO_1933 (O_1933,N_20975,N_24743);
and UO_1934 (O_1934,N_22324,N_23763);
and UO_1935 (O_1935,N_21028,N_21667);
xor UO_1936 (O_1936,N_23411,N_20128);
or UO_1937 (O_1937,N_20283,N_20457);
or UO_1938 (O_1938,N_22326,N_21394);
and UO_1939 (O_1939,N_24804,N_24168);
and UO_1940 (O_1940,N_21862,N_24814);
nand UO_1941 (O_1941,N_24226,N_22481);
and UO_1942 (O_1942,N_22766,N_24599);
nor UO_1943 (O_1943,N_22436,N_23338);
or UO_1944 (O_1944,N_24206,N_21524);
or UO_1945 (O_1945,N_23275,N_23937);
or UO_1946 (O_1946,N_20876,N_21739);
nand UO_1947 (O_1947,N_23220,N_24063);
nand UO_1948 (O_1948,N_20736,N_22494);
or UO_1949 (O_1949,N_23986,N_21212);
nand UO_1950 (O_1950,N_24192,N_22291);
and UO_1951 (O_1951,N_21664,N_20464);
nand UO_1952 (O_1952,N_22333,N_23445);
or UO_1953 (O_1953,N_23087,N_20058);
nand UO_1954 (O_1954,N_21264,N_21401);
or UO_1955 (O_1955,N_21458,N_24606);
and UO_1956 (O_1956,N_22384,N_20994);
and UO_1957 (O_1957,N_22488,N_23590);
and UO_1958 (O_1958,N_24491,N_20593);
xnor UO_1959 (O_1959,N_21467,N_22973);
nor UO_1960 (O_1960,N_24387,N_21731);
or UO_1961 (O_1961,N_20509,N_20090);
nand UO_1962 (O_1962,N_20095,N_21438);
nand UO_1963 (O_1963,N_24981,N_20173);
nor UO_1964 (O_1964,N_24439,N_24672);
and UO_1965 (O_1965,N_24142,N_22364);
nand UO_1966 (O_1966,N_24362,N_24315);
nand UO_1967 (O_1967,N_22441,N_21364);
xor UO_1968 (O_1968,N_21327,N_24952);
nor UO_1969 (O_1969,N_21776,N_20051);
nor UO_1970 (O_1970,N_21185,N_20667);
or UO_1971 (O_1971,N_24964,N_22660);
or UO_1972 (O_1972,N_23212,N_24556);
and UO_1973 (O_1973,N_23690,N_23580);
or UO_1974 (O_1974,N_22578,N_23486);
nand UO_1975 (O_1975,N_23886,N_22401);
and UO_1976 (O_1976,N_24433,N_24937);
nand UO_1977 (O_1977,N_24450,N_23566);
and UO_1978 (O_1978,N_24326,N_23319);
nand UO_1979 (O_1979,N_20108,N_21733);
or UO_1980 (O_1980,N_20740,N_20403);
nand UO_1981 (O_1981,N_22115,N_20814);
nand UO_1982 (O_1982,N_20715,N_22011);
nand UO_1983 (O_1983,N_22493,N_21715);
and UO_1984 (O_1984,N_24391,N_23630);
nand UO_1985 (O_1985,N_20080,N_21749);
nand UO_1986 (O_1986,N_23998,N_20483);
or UO_1987 (O_1987,N_23400,N_22512);
and UO_1988 (O_1988,N_22054,N_24783);
nand UO_1989 (O_1989,N_21290,N_22249);
nor UO_1990 (O_1990,N_23675,N_21456);
nand UO_1991 (O_1991,N_22800,N_20684);
nand UO_1992 (O_1992,N_20776,N_22337);
or UO_1993 (O_1993,N_24352,N_23205);
nand UO_1994 (O_1994,N_24640,N_24534);
and UO_1995 (O_1995,N_23902,N_23640);
and UO_1996 (O_1996,N_22751,N_23061);
nor UO_1997 (O_1997,N_20110,N_20704);
or UO_1998 (O_1998,N_23995,N_22545);
nor UO_1999 (O_1999,N_20914,N_24422);
nand UO_2000 (O_2000,N_24410,N_24177);
nand UO_2001 (O_2001,N_20703,N_21310);
nand UO_2002 (O_2002,N_24527,N_23694);
nand UO_2003 (O_2003,N_23754,N_23599);
nor UO_2004 (O_2004,N_23696,N_23323);
nor UO_2005 (O_2005,N_22818,N_24068);
and UO_2006 (O_2006,N_23972,N_24961);
xor UO_2007 (O_2007,N_22698,N_23185);
or UO_2008 (O_2008,N_23334,N_20997);
nor UO_2009 (O_2009,N_21313,N_21339);
and UO_2010 (O_2010,N_23285,N_23530);
nand UO_2011 (O_2011,N_24154,N_24877);
nor UO_2012 (O_2012,N_24581,N_23031);
and UO_2013 (O_2013,N_23006,N_20418);
and UO_2014 (O_2014,N_24821,N_24267);
or UO_2015 (O_2015,N_21611,N_22315);
or UO_2016 (O_2016,N_20676,N_24185);
nand UO_2017 (O_2017,N_20864,N_23856);
and UO_2018 (O_2018,N_24925,N_22530);
or UO_2019 (O_2019,N_24164,N_20314);
nand UO_2020 (O_2020,N_21059,N_23202);
nor UO_2021 (O_2021,N_21553,N_24072);
and UO_2022 (O_2022,N_22571,N_23461);
and UO_2023 (O_2023,N_21305,N_23829);
nor UO_2024 (O_2024,N_21746,N_20354);
xnor UO_2025 (O_2025,N_23716,N_20854);
or UO_2026 (O_2026,N_24590,N_20476);
or UO_2027 (O_2027,N_21380,N_21032);
xor UO_2028 (O_2028,N_23862,N_20552);
nand UO_2029 (O_2029,N_24288,N_21187);
xor UO_2030 (O_2030,N_22419,N_23125);
or UO_2031 (O_2031,N_20009,N_24171);
nand UO_2032 (O_2032,N_24922,N_23919);
nor UO_2033 (O_2033,N_22967,N_20955);
xor UO_2034 (O_2034,N_24657,N_22568);
xor UO_2035 (O_2035,N_20602,N_24997);
or UO_2036 (O_2036,N_22070,N_20883);
nand UO_2037 (O_2037,N_22304,N_21346);
nand UO_2038 (O_2038,N_20034,N_24715);
nor UO_2039 (O_2039,N_22538,N_20586);
or UO_2040 (O_2040,N_22065,N_21980);
nand UO_2041 (O_2041,N_20634,N_22689);
xor UO_2042 (O_2042,N_24732,N_21086);
and UO_2043 (O_2043,N_21853,N_20614);
nand UO_2044 (O_2044,N_23044,N_21137);
nor UO_2045 (O_2045,N_23910,N_22265);
nand UO_2046 (O_2046,N_24283,N_22072);
and UO_2047 (O_2047,N_20451,N_21225);
or UO_2048 (O_2048,N_24031,N_22473);
nand UO_2049 (O_2049,N_22023,N_24819);
or UO_2050 (O_2050,N_22476,N_24603);
or UO_2051 (O_2051,N_20635,N_20340);
and UO_2052 (O_2052,N_20520,N_24342);
nand UO_2053 (O_2053,N_24767,N_21473);
nor UO_2054 (O_2054,N_22734,N_23527);
or UO_2055 (O_2055,N_21858,N_21655);
nor UO_2056 (O_2056,N_20397,N_24452);
or UO_2057 (O_2057,N_24011,N_20787);
and UO_2058 (O_2058,N_22702,N_21673);
nand UO_2059 (O_2059,N_21833,N_21349);
and UO_2060 (O_2060,N_24545,N_24673);
and UO_2061 (O_2061,N_21011,N_24522);
nor UO_2062 (O_2062,N_23497,N_22111);
and UO_2063 (O_2063,N_24785,N_24627);
nor UO_2064 (O_2064,N_23117,N_22008);
and UO_2065 (O_2065,N_20741,N_20526);
nand UO_2066 (O_2066,N_23966,N_20005);
and UO_2067 (O_2067,N_23707,N_24200);
or UO_2068 (O_2068,N_22100,N_24262);
nor UO_2069 (O_2069,N_21421,N_20589);
or UO_2070 (O_2070,N_24407,N_22443);
nor UO_2071 (O_2071,N_21300,N_21582);
or UO_2072 (O_2072,N_22610,N_22202);
nand UO_2073 (O_2073,N_24919,N_22835);
or UO_2074 (O_2074,N_20767,N_22840);
or UO_2075 (O_2075,N_20560,N_24383);
nand UO_2076 (O_2076,N_24562,N_21112);
or UO_2077 (O_2077,N_23731,N_24250);
or UO_2078 (O_2078,N_22020,N_24530);
or UO_2079 (O_2079,N_21132,N_21233);
and UO_2080 (O_2080,N_21101,N_21222);
or UO_2081 (O_2081,N_21447,N_23852);
or UO_2082 (O_2082,N_22961,N_23614);
and UO_2083 (O_2083,N_24249,N_24460);
nand UO_2084 (O_2084,N_21081,N_24365);
nand UO_2085 (O_2085,N_20306,N_20060);
or UO_2086 (O_2086,N_24984,N_23873);
nand UO_2087 (O_2087,N_23279,N_22845);
or UO_2088 (O_2088,N_24078,N_24963);
and UO_2089 (O_2089,N_23905,N_20506);
or UO_2090 (O_2090,N_24247,N_23866);
nor UO_2091 (O_2091,N_21044,N_22003);
nand UO_2092 (O_2092,N_21973,N_20364);
nor UO_2093 (O_2093,N_24918,N_23592);
and UO_2094 (O_2094,N_23753,N_22258);
or UO_2095 (O_2095,N_22514,N_22700);
and UO_2096 (O_2096,N_20927,N_23869);
nor UO_2097 (O_2097,N_24036,N_23698);
or UO_2098 (O_2098,N_24933,N_21449);
nor UO_2099 (O_2099,N_23123,N_24222);
nand UO_2100 (O_2100,N_21593,N_21459);
or UO_2101 (O_2101,N_20307,N_23103);
nor UO_2102 (O_2102,N_20045,N_21224);
nor UO_2103 (O_2103,N_22865,N_20345);
nor UO_2104 (O_2104,N_23586,N_22019);
nor UO_2105 (O_2105,N_23668,N_23160);
nand UO_2106 (O_2106,N_23844,N_23926);
nor UO_2107 (O_2107,N_20490,N_23417);
nor UO_2108 (O_2108,N_22360,N_20806);
and UO_2109 (O_2109,N_23447,N_21375);
nor UO_2110 (O_2110,N_20754,N_22160);
or UO_2111 (O_2111,N_24794,N_21171);
nor UO_2112 (O_2112,N_23865,N_21509);
nand UO_2113 (O_2113,N_23047,N_20225);
and UO_2114 (O_2114,N_21045,N_21968);
nand UO_2115 (O_2115,N_22864,N_22867);
nand UO_2116 (O_2116,N_21921,N_22905);
nor UO_2117 (O_2117,N_24662,N_22409);
nor UO_2118 (O_2118,N_21190,N_23556);
nand UO_2119 (O_2119,N_23032,N_23996);
xor UO_2120 (O_2120,N_24119,N_20205);
or UO_2121 (O_2121,N_23597,N_23771);
and UO_2122 (O_2122,N_23534,N_23259);
or UO_2123 (O_2123,N_20281,N_24381);
and UO_2124 (O_2124,N_20047,N_24956);
and UO_2125 (O_2125,N_24719,N_22387);
or UO_2126 (O_2126,N_24395,N_22547);
and UO_2127 (O_2127,N_21750,N_23843);
or UO_2128 (O_2128,N_23368,N_24645);
nand UO_2129 (O_2129,N_22762,N_24061);
xor UO_2130 (O_2130,N_20738,N_21175);
nor UO_2131 (O_2131,N_24867,N_23039);
nand UO_2132 (O_2132,N_20533,N_20584);
nand UO_2133 (O_2133,N_24385,N_22552);
and UO_2134 (O_2134,N_22916,N_22862);
nor UO_2135 (O_2135,N_22442,N_20392);
or UO_2136 (O_2136,N_22284,N_21756);
nor UO_2137 (O_2137,N_21260,N_20514);
and UO_2138 (O_2138,N_22575,N_24368);
or UO_2139 (O_2139,N_20414,N_21116);
or UO_2140 (O_2140,N_20278,N_23312);
or UO_2141 (O_2141,N_23791,N_20598);
xnor UO_2142 (O_2142,N_20417,N_21080);
and UO_2143 (O_2143,N_24275,N_20073);
nor UO_2144 (O_2144,N_22338,N_22771);
and UO_2145 (O_2145,N_24703,N_22812);
or UO_2146 (O_2146,N_24083,N_20460);
nor UO_2147 (O_2147,N_22799,N_22796);
nor UO_2148 (O_2148,N_21341,N_23014);
and UO_2149 (O_2149,N_21707,N_23219);
nand UO_2150 (O_2150,N_24520,N_23146);
or UO_2151 (O_2151,N_21440,N_21591);
or UO_2152 (O_2152,N_22982,N_21295);
nor UO_2153 (O_2153,N_21617,N_23733);
nor UO_2154 (O_2154,N_22671,N_20270);
nand UO_2155 (O_2155,N_23115,N_24322);
or UO_2156 (O_2156,N_22059,N_22343);
nor UO_2157 (O_2157,N_20643,N_23904);
or UO_2158 (O_2158,N_20485,N_23903);
and UO_2159 (O_2159,N_24512,N_21236);
nand UO_2160 (O_2160,N_22903,N_24823);
and UO_2161 (O_2161,N_21651,N_21941);
and UO_2162 (O_2162,N_22144,N_21893);
and UO_2163 (O_2163,N_23555,N_23861);
nand UO_2164 (O_2164,N_21598,N_20002);
or UO_2165 (O_2165,N_23446,N_21726);
and UO_2166 (O_2166,N_20341,N_24193);
and UO_2167 (O_2167,N_24713,N_20984);
or UO_2168 (O_2168,N_21148,N_23256);
nor UO_2169 (O_2169,N_22979,N_23332);
nor UO_2170 (O_2170,N_21126,N_21765);
or UO_2171 (O_2171,N_23808,N_23542);
and UO_2172 (O_2172,N_22041,N_23438);
nor UO_2173 (O_2173,N_23102,N_23839);
nor UO_2174 (O_2174,N_23420,N_20745);
or UO_2175 (O_2175,N_24033,N_24760);
nor UO_2176 (O_2176,N_22323,N_23985);
nand UO_2177 (O_2177,N_21323,N_21590);
nor UO_2178 (O_2178,N_23019,N_20882);
nor UO_2179 (O_2179,N_20626,N_22627);
nand UO_2180 (O_2180,N_22246,N_20074);
and UO_2181 (O_2181,N_24028,N_20159);
or UO_2182 (O_2182,N_21938,N_24118);
nor UO_2183 (O_2183,N_22866,N_20679);
or UO_2184 (O_2184,N_21836,N_21273);
nand UO_2185 (O_2185,N_22078,N_23158);
and UO_2186 (O_2186,N_24731,N_21872);
nor UO_2187 (O_2187,N_20068,N_23664);
and UO_2188 (O_2188,N_24067,N_20290);
nor UO_2189 (O_2189,N_24150,N_21905);
nor UO_2190 (O_2190,N_23330,N_21494);
or UO_2191 (O_2191,N_23969,N_22699);
or UO_2192 (O_2192,N_24960,N_23292);
and UO_2193 (O_2193,N_20558,N_24629);
nand UO_2194 (O_2194,N_21873,N_24059);
nand UO_2195 (O_2195,N_23329,N_20800);
nand UO_2196 (O_2196,N_23088,N_21128);
or UO_2197 (O_2197,N_22174,N_20631);
and UO_2198 (O_2198,N_20233,N_23807);
nand UO_2199 (O_2199,N_20013,N_23262);
nor UO_2200 (O_2200,N_23894,N_20325);
nand UO_2201 (O_2201,N_22138,N_24084);
nor UO_2202 (O_2202,N_24443,N_20818);
nor UO_2203 (O_2203,N_22479,N_22816);
or UO_2204 (O_2204,N_22964,N_21728);
or UO_2205 (O_2205,N_20874,N_21466);
or UO_2206 (O_2206,N_24939,N_20198);
nand UO_2207 (O_2207,N_22780,N_21774);
nor UO_2208 (O_2208,N_23075,N_23206);
nand UO_2209 (O_2209,N_23840,N_21307);
and UO_2210 (O_2210,N_22871,N_23393);
and UO_2211 (O_2211,N_24650,N_22467);
or UO_2212 (O_2212,N_21444,N_24454);
nor UO_2213 (O_2213,N_20547,N_24870);
nand UO_2214 (O_2214,N_20747,N_20494);
or UO_2215 (O_2215,N_24516,N_22881);
nor UO_2216 (O_2216,N_20534,N_21676);
or UO_2217 (O_2217,N_22308,N_24764);
or UO_2218 (O_2218,N_24475,N_24973);
and UO_2219 (O_2219,N_22938,N_22171);
or UO_2220 (O_2220,N_24130,N_22278);
and UO_2221 (O_2221,N_20530,N_22262);
nor UO_2222 (O_2222,N_21399,N_23238);
or UO_2223 (O_2223,N_22034,N_22215);
and UO_2224 (O_2224,N_21868,N_22449);
nand UO_2225 (O_2225,N_20203,N_22776);
nand UO_2226 (O_2226,N_20742,N_20282);
or UO_2227 (O_2227,N_22810,N_22209);
or UO_2228 (O_2228,N_20328,N_22566);
and UO_2229 (O_2229,N_23490,N_20755);
nor UO_2230 (O_2230,N_21213,N_24604);
nand UO_2231 (O_2231,N_23835,N_20062);
nand UO_2232 (O_2232,N_22509,N_23467);
xor UO_2233 (O_2233,N_20835,N_21542);
nor UO_2234 (O_2234,N_22635,N_24045);
nor UO_2235 (O_2235,N_23366,N_22272);
and UO_2236 (O_2236,N_20077,N_23832);
nand UO_2237 (O_2237,N_20286,N_20399);
and UO_2238 (O_2238,N_23700,N_24010);
and UO_2239 (O_2239,N_22339,N_24287);
nand UO_2240 (O_2240,N_21249,N_20769);
or UO_2241 (O_2241,N_21874,N_23770);
nor UO_2242 (O_2242,N_24904,N_23268);
and UO_2243 (O_2243,N_22157,N_21781);
nand UO_2244 (O_2244,N_23363,N_21969);
nand UO_2245 (O_2245,N_23406,N_21960);
and UO_2246 (O_2246,N_20804,N_23834);
nand UO_2247 (O_2247,N_20516,N_23761);
nand UO_2248 (O_2248,N_22659,N_22385);
nand UO_2249 (O_2249,N_21878,N_23350);
and UO_2250 (O_2250,N_22705,N_24773);
nor UO_2251 (O_2251,N_22082,N_20523);
nand UO_2252 (O_2252,N_22977,N_21686);
or UO_2253 (O_2253,N_22863,N_22195);
or UO_2254 (O_2254,N_20947,N_22429);
or UO_2255 (O_2255,N_21572,N_21902);
nand UO_2256 (O_2256,N_24708,N_21106);
nand UO_2257 (O_2257,N_20503,N_20299);
nor UO_2258 (O_2258,N_21484,N_20216);
nand UO_2259 (O_2259,N_24244,N_21714);
nand UO_2260 (O_2260,N_20555,N_22254);
or UO_2261 (O_2261,N_22774,N_20232);
and UO_2262 (O_2262,N_20359,N_24442);
and UO_2263 (O_2263,N_22462,N_24942);
or UO_2264 (O_2264,N_24016,N_20093);
nand UO_2265 (O_2265,N_24958,N_24259);
nor UO_2266 (O_2266,N_24544,N_22073);
and UO_2267 (O_2267,N_22851,N_24139);
and UO_2268 (O_2268,N_20195,N_20941);
nand UO_2269 (O_2269,N_23848,N_23923);
and UO_2270 (O_2270,N_23139,N_24745);
or UO_2271 (O_2271,N_21376,N_24791);
and UO_2272 (O_2272,N_23612,N_24946);
nor UO_2273 (O_2273,N_24898,N_24975);
or UO_2274 (O_2274,N_24052,N_23257);
and UO_2275 (O_2275,N_23927,N_23786);
nor UO_2276 (O_2276,N_21537,N_21694);
nand UO_2277 (O_2277,N_21775,N_24616);
and UO_2278 (O_2278,N_22147,N_21805);
nand UO_2279 (O_2279,N_24188,N_22432);
or UO_2280 (O_2280,N_24172,N_24611);
or UO_2281 (O_2281,N_20869,N_24295);
nor UO_2282 (O_2282,N_21157,N_24908);
nand UO_2283 (O_2283,N_22976,N_23713);
or UO_2284 (O_2284,N_24834,N_20734);
and UO_2285 (O_2285,N_23429,N_24885);
nor UO_2286 (O_2286,N_23961,N_24675);
and UO_2287 (O_2287,N_21036,N_22773);
nor UO_2288 (O_2288,N_24716,N_20142);
and UO_2289 (O_2289,N_20192,N_22133);
nand UO_2290 (O_2290,N_20765,N_24184);
nor UO_2291 (O_2291,N_20720,N_24573);
nor UO_2292 (O_2292,N_21186,N_20400);
and UO_2293 (O_2293,N_24493,N_24547);
or UO_2294 (O_2294,N_21799,N_23488);
and UO_2295 (O_2295,N_22055,N_23460);
xor UO_2296 (O_2296,N_24549,N_22025);
nand UO_2297 (O_2297,N_20694,N_23774);
nand UO_2298 (O_2298,N_20848,N_21210);
nor UO_2299 (O_2299,N_20782,N_22325);
nor UO_2300 (O_2300,N_24994,N_20291);
and UO_2301 (O_2301,N_24567,N_20224);
or UO_2302 (O_2302,N_20085,N_23740);
or UO_2303 (O_2303,N_21949,N_22075);
nand UO_2304 (O_2304,N_22120,N_21695);
and UO_2305 (O_2305,N_23683,N_24602);
nor UO_2306 (O_2306,N_20387,N_21268);
nor UO_2307 (O_2307,N_21649,N_23893);
nor UO_2308 (O_2308,N_20844,N_24014);
and UO_2309 (O_2309,N_23230,N_23228);
and UO_2310 (O_2310,N_24159,N_23254);
and UO_2311 (O_2311,N_21504,N_22348);
and UO_2312 (O_2312,N_22533,N_24468);
nand UO_2313 (O_2313,N_21180,N_21522);
or UO_2314 (O_2314,N_23249,N_20440);
nor UO_2315 (O_2315,N_22562,N_24227);
nand UO_2316 (O_2316,N_23295,N_20449);
or UO_2317 (O_2317,N_21109,N_22212);
nand UO_2318 (O_2318,N_22941,N_20971);
nand UO_2319 (O_2319,N_21356,N_20977);
nor UO_2320 (O_2320,N_22683,N_20466);
or UO_2321 (O_2321,N_20432,N_20750);
nor UO_2322 (O_2322,N_20007,N_21285);
and UO_2323 (O_2323,N_20180,N_21666);
or UO_2324 (O_2324,N_24789,N_22201);
nand UO_2325 (O_2325,N_20277,N_21866);
or UO_2326 (O_2326,N_24607,N_23025);
or UO_2327 (O_2327,N_23496,N_23154);
and UO_2328 (O_2328,N_22269,N_20519);
nor UO_2329 (O_2329,N_21085,N_21939);
and UO_2330 (O_2330,N_21716,N_23344);
nand UO_2331 (O_2331,N_23975,N_24020);
nand UO_2332 (O_2332,N_22474,N_23261);
nor UO_2333 (O_2333,N_21216,N_21120);
nor UO_2334 (O_2334,N_24451,N_21914);
and UO_2335 (O_2335,N_23579,N_24953);
nand UO_2336 (O_2336,N_21959,N_22569);
nand UO_2337 (O_2337,N_21786,N_20653);
or UO_2338 (O_2338,N_21720,N_20668);
or UO_2339 (O_2339,N_22715,N_21054);
nand UO_2340 (O_2340,N_23537,N_24215);
nand UO_2341 (O_2341,N_21512,N_22879);
and UO_2342 (O_2342,N_20342,N_24723);
and UO_2343 (O_2343,N_23100,N_21123);
nand UO_2344 (O_2344,N_23166,N_20739);
nor UO_2345 (O_2345,N_22273,N_21953);
nor UO_2346 (O_2346,N_23737,N_24717);
nand UO_2347 (O_2347,N_20362,N_23804);
nor UO_2348 (O_2348,N_22259,N_24473);
nand UO_2349 (O_2349,N_21280,N_20834);
nor UO_2350 (O_2350,N_22356,N_20960);
nand UO_2351 (O_2351,N_24235,N_21773);
nor UO_2352 (O_2352,N_22306,N_22740);
nand UO_2353 (O_2353,N_20322,N_23455);
nand UO_2354 (O_2354,N_22855,N_22328);
and UO_2355 (O_2355,N_22709,N_23080);
nand UO_2356 (O_2356,N_23374,N_22208);
or UO_2357 (O_2357,N_23282,N_22486);
or UO_2358 (O_2358,N_20042,N_21894);
nor UO_2359 (O_2359,N_21343,N_22592);
nand UO_2360 (O_2360,N_24751,N_22948);
and UO_2361 (O_2361,N_22599,N_22570);
nand UO_2362 (O_2362,N_21056,N_22156);
nand UO_2363 (O_2363,N_22076,N_20925);
and UO_2364 (O_2364,N_20214,N_21791);
and UO_2365 (O_2365,N_21618,N_22661);
or UO_2366 (O_2366,N_23314,N_24182);
and UO_2367 (O_2367,N_24113,N_23321);
nor UO_2368 (O_2368,N_24843,N_24705);
and UO_2369 (O_2369,N_23777,N_23407);
or UO_2370 (O_2370,N_23459,N_22622);
nand UO_2371 (O_2371,N_22319,N_22804);
nand UO_2372 (O_2372,N_24542,N_23787);
nand UO_2373 (O_2373,N_20409,N_22625);
nor UO_2374 (O_2374,N_23183,N_23997);
nor UO_2375 (O_2375,N_23738,N_24485);
or UO_2376 (O_2376,N_21005,N_21491);
and UO_2377 (O_2377,N_20886,N_20968);
nand UO_2378 (O_2378,N_23531,N_22042);
nor UO_2379 (O_2379,N_24891,N_20201);
nor UO_2380 (O_2380,N_21727,N_22230);
nor UO_2381 (O_2381,N_20148,N_21483);
nor UO_2382 (O_2382,N_23729,N_21164);
nand UO_2383 (O_2383,N_21311,N_22595);
nor UO_2384 (O_2384,N_24135,N_24921);
and UO_2385 (O_2385,N_23150,N_23742);
and UO_2386 (O_2386,N_21857,N_21303);
nor UO_2387 (O_2387,N_23130,N_21705);
and UO_2388 (O_2388,N_20197,N_22329);
and UO_2389 (O_2389,N_23529,N_22912);
nand UO_2390 (O_2390,N_22824,N_23900);
nor UO_2391 (O_2391,N_24572,N_24793);
and UO_2392 (O_2392,N_20143,N_20729);
nor UO_2393 (O_2393,N_24510,N_23660);
nand UO_2394 (O_2394,N_23441,N_23478);
nand UO_2395 (O_2395,N_20132,N_24252);
nor UO_2396 (O_2396,N_20696,N_24064);
or UO_2397 (O_2397,N_21065,N_21416);
and UO_2398 (O_2398,N_24343,N_21414);
nor UO_2399 (O_2399,N_24868,N_20548);
nand UO_2400 (O_2400,N_20452,N_23836);
nor UO_2401 (O_2401,N_24332,N_22381);
or UO_2402 (O_2402,N_21198,N_24060);
nor UO_2403 (O_2403,N_23695,N_21472);
nand UO_2404 (O_2404,N_21818,N_24486);
nand UO_2405 (O_2405,N_23173,N_24290);
nor UO_2406 (O_2406,N_24948,N_23342);
nor UO_2407 (O_2407,N_21386,N_22534);
and UO_2408 (O_2408,N_22221,N_21209);
or UO_2409 (O_2409,N_23094,N_22849);
nor UO_2410 (O_2410,N_24874,N_23493);
nand UO_2411 (O_2411,N_21940,N_23369);
nand UO_2412 (O_2412,N_22418,N_24178);
nor UO_2413 (O_2413,N_22584,N_24239);
nand UO_2414 (O_2414,N_23727,N_20395);
and UO_2415 (O_2415,N_21046,N_23610);
nand UO_2416 (O_2416,N_23813,N_21242);
nand UO_2417 (O_2417,N_24181,N_20973);
or UO_2418 (O_2418,N_21910,N_22965);
nor UO_2419 (O_2419,N_20384,N_24513);
or UO_2420 (O_2420,N_24710,N_21711);
nand UO_2421 (O_2421,N_22895,N_22694);
or UO_2422 (O_2422,N_24967,N_22695);
or UO_2423 (O_2423,N_21924,N_24108);
and UO_2424 (O_2424,N_23336,N_21908);
nor UO_2425 (O_2425,N_24619,N_22978);
or UO_2426 (O_2426,N_23649,N_22379);
and UO_2427 (O_2427,N_21396,N_22497);
nor UO_2428 (O_2428,N_21523,N_23234);
or UO_2429 (O_2429,N_24080,N_24044);
or UO_2430 (O_2430,N_22525,N_21498);
nor UO_2431 (O_2431,N_24744,N_24260);
and UO_2432 (O_2432,N_20557,N_22152);
nand UO_2433 (O_2433,N_24829,N_24837);
or UO_2434 (O_2434,N_22918,N_23041);
and UO_2435 (O_2435,N_23546,N_21234);
or UO_2436 (O_2436,N_24427,N_23992);
nor UO_2437 (O_2437,N_23016,N_24538);
nand UO_2438 (O_2438,N_24658,N_22684);
nand UO_2439 (O_2439,N_24103,N_21470);
nand UO_2440 (O_2440,N_24498,N_23574);
nor UO_2441 (O_2441,N_22749,N_21769);
or UO_2442 (O_2442,N_21362,N_20230);
nand UO_2443 (O_2443,N_23303,N_20048);
or UO_2444 (O_2444,N_21070,N_20222);
and UO_2445 (O_2445,N_20477,N_24666);
nor UO_2446 (O_2446,N_24916,N_24316);
or UO_2447 (O_2447,N_22561,N_21500);
nor UO_2448 (O_2448,N_21656,N_22725);
and UO_2449 (O_2449,N_22199,N_22872);
or UO_2450 (O_2450,N_24435,N_21519);
nor UO_2451 (O_2451,N_24136,N_20920);
or UO_2452 (O_2452,N_22450,N_21402);
or UO_2453 (O_2453,N_24655,N_20166);
nand UO_2454 (O_2454,N_23378,N_21644);
or UO_2455 (O_2455,N_22451,N_23666);
xor UO_2456 (O_2456,N_22841,N_21146);
nor UO_2457 (O_2457,N_20292,N_24757);
and UO_2458 (O_2458,N_21092,N_20445);
nand UO_2459 (O_2459,N_22056,N_20878);
and UO_2460 (O_2460,N_24734,N_21621);
nand UO_2461 (O_2461,N_21616,N_21201);
and UO_2462 (O_2462,N_24927,N_22984);
nand UO_2463 (O_2463,N_20829,N_20022);
nor UO_2464 (O_2464,N_22808,N_22332);
or UO_2465 (O_2465,N_20386,N_21016);
xor UO_2466 (O_2466,N_23475,N_24811);
xnor UO_2467 (O_2467,N_20336,N_22953);
and UO_2468 (O_2468,N_21021,N_24559);
nand UO_2469 (O_2469,N_23410,N_23416);
nor UO_2470 (O_2470,N_24266,N_21624);
nand UO_2471 (O_2471,N_24230,N_22952);
nor UO_2472 (O_2472,N_20966,N_21725);
or UO_2473 (O_2473,N_20084,N_22096);
nor UO_2474 (O_2474,N_20020,N_24873);
and UO_2475 (O_2475,N_23585,N_24838);
nand UO_2476 (O_2476,N_22747,N_20823);
or UO_2477 (O_2477,N_23452,N_23157);
nor UO_2478 (O_2478,N_24851,N_24348);
or UO_2479 (O_2479,N_23109,N_21238);
nor UO_2480 (O_2480,N_24280,N_20789);
nand UO_2481 (O_2481,N_21274,N_20655);
and UO_2482 (O_2482,N_20688,N_20540);
or UO_2483 (O_2483,N_24257,N_20942);
and UO_2484 (O_2484,N_24176,N_23799);
and UO_2485 (O_2485,N_22270,N_23269);
or UO_2486 (O_2486,N_24423,N_23470);
nor UO_2487 (O_2487,N_23120,N_24909);
nor UO_2488 (O_2488,N_21533,N_21255);
or UO_2489 (O_2489,N_20465,N_22021);
nand UO_2490 (O_2490,N_24311,N_21173);
and UO_2491 (O_2491,N_24947,N_24896);
and UO_2492 (O_2492,N_21596,N_21025);
or UO_2493 (O_2493,N_21811,N_20472);
and UO_2494 (O_2494,N_22655,N_22832);
or UO_2495 (O_2495,N_22573,N_23842);
xor UO_2496 (O_2496,N_20665,N_20877);
or UO_2497 (O_2497,N_22469,N_23935);
nand UO_2498 (O_2498,N_20486,N_20710);
nand UO_2499 (O_2499,N_20726,N_24704);
and UO_2500 (O_2500,N_20672,N_24472);
nor UO_2501 (O_2501,N_24908,N_20310);
nor UO_2502 (O_2502,N_24053,N_23086);
and UO_2503 (O_2503,N_20587,N_21746);
nor UO_2504 (O_2504,N_23478,N_22309);
nor UO_2505 (O_2505,N_22385,N_23030);
and UO_2506 (O_2506,N_22107,N_23980);
xor UO_2507 (O_2507,N_23710,N_22809);
nand UO_2508 (O_2508,N_24844,N_24803);
and UO_2509 (O_2509,N_23833,N_22928);
nand UO_2510 (O_2510,N_23046,N_22615);
nor UO_2511 (O_2511,N_21308,N_24139);
and UO_2512 (O_2512,N_23543,N_21433);
nor UO_2513 (O_2513,N_22825,N_22575);
or UO_2514 (O_2514,N_23226,N_20307);
nand UO_2515 (O_2515,N_23590,N_24583);
or UO_2516 (O_2516,N_20933,N_23880);
nand UO_2517 (O_2517,N_24787,N_23028);
and UO_2518 (O_2518,N_20593,N_23436);
nand UO_2519 (O_2519,N_24475,N_22112);
or UO_2520 (O_2520,N_21385,N_21087);
and UO_2521 (O_2521,N_22320,N_22101);
nor UO_2522 (O_2522,N_20538,N_20520);
nand UO_2523 (O_2523,N_23819,N_22817);
and UO_2524 (O_2524,N_22147,N_23007);
nand UO_2525 (O_2525,N_24336,N_22252);
nand UO_2526 (O_2526,N_21051,N_24725);
and UO_2527 (O_2527,N_24509,N_22959);
or UO_2528 (O_2528,N_23903,N_22405);
and UO_2529 (O_2529,N_20551,N_20201);
and UO_2530 (O_2530,N_22505,N_21012);
nand UO_2531 (O_2531,N_23829,N_22793);
and UO_2532 (O_2532,N_21005,N_21740);
nand UO_2533 (O_2533,N_24506,N_21196);
nor UO_2534 (O_2534,N_21530,N_24550);
nand UO_2535 (O_2535,N_22934,N_23633);
nor UO_2536 (O_2536,N_22758,N_24401);
nor UO_2537 (O_2537,N_21711,N_24981);
or UO_2538 (O_2538,N_24126,N_22475);
nand UO_2539 (O_2539,N_24034,N_24225);
nor UO_2540 (O_2540,N_23715,N_22660);
or UO_2541 (O_2541,N_22447,N_23596);
and UO_2542 (O_2542,N_20133,N_20412);
nand UO_2543 (O_2543,N_21583,N_24445);
nor UO_2544 (O_2544,N_23464,N_23633);
or UO_2545 (O_2545,N_23631,N_23465);
nand UO_2546 (O_2546,N_20333,N_24100);
and UO_2547 (O_2547,N_20296,N_22738);
and UO_2548 (O_2548,N_21794,N_22556);
nor UO_2549 (O_2549,N_24696,N_22998);
or UO_2550 (O_2550,N_23468,N_20882);
nor UO_2551 (O_2551,N_20873,N_24327);
nand UO_2552 (O_2552,N_20424,N_20173);
nand UO_2553 (O_2553,N_24677,N_23222);
and UO_2554 (O_2554,N_22323,N_20412);
or UO_2555 (O_2555,N_22908,N_24432);
and UO_2556 (O_2556,N_24367,N_21665);
nand UO_2557 (O_2557,N_24643,N_22639);
and UO_2558 (O_2558,N_22877,N_23785);
and UO_2559 (O_2559,N_20774,N_23784);
nor UO_2560 (O_2560,N_23832,N_24817);
and UO_2561 (O_2561,N_23146,N_21125);
nand UO_2562 (O_2562,N_22208,N_21192);
nand UO_2563 (O_2563,N_22607,N_20714);
or UO_2564 (O_2564,N_23437,N_22295);
nand UO_2565 (O_2565,N_24820,N_20539);
xor UO_2566 (O_2566,N_24854,N_22715);
nor UO_2567 (O_2567,N_22848,N_23635);
nor UO_2568 (O_2568,N_23922,N_23691);
nor UO_2569 (O_2569,N_22667,N_23629);
nand UO_2570 (O_2570,N_22031,N_21622);
nor UO_2571 (O_2571,N_22144,N_23773);
nand UO_2572 (O_2572,N_22352,N_21408);
and UO_2573 (O_2573,N_21615,N_21542);
and UO_2574 (O_2574,N_23418,N_24561);
nor UO_2575 (O_2575,N_24693,N_21444);
or UO_2576 (O_2576,N_20226,N_21575);
or UO_2577 (O_2577,N_22646,N_24020);
nand UO_2578 (O_2578,N_21626,N_22782);
nand UO_2579 (O_2579,N_24184,N_22337);
nor UO_2580 (O_2580,N_22144,N_24357);
or UO_2581 (O_2581,N_23702,N_23497);
nor UO_2582 (O_2582,N_21160,N_22376);
nor UO_2583 (O_2583,N_24713,N_24160);
nand UO_2584 (O_2584,N_20077,N_20100);
nor UO_2585 (O_2585,N_21549,N_20673);
nand UO_2586 (O_2586,N_24812,N_21349);
nor UO_2587 (O_2587,N_21897,N_23748);
and UO_2588 (O_2588,N_24189,N_24399);
or UO_2589 (O_2589,N_22113,N_23709);
xor UO_2590 (O_2590,N_20056,N_24871);
nor UO_2591 (O_2591,N_24884,N_24180);
nand UO_2592 (O_2592,N_20678,N_23247);
or UO_2593 (O_2593,N_21861,N_23067);
and UO_2594 (O_2594,N_21425,N_22223);
or UO_2595 (O_2595,N_20001,N_20767);
nor UO_2596 (O_2596,N_22744,N_22787);
nand UO_2597 (O_2597,N_21652,N_22148);
and UO_2598 (O_2598,N_21954,N_23409);
nor UO_2599 (O_2599,N_23261,N_21631);
or UO_2600 (O_2600,N_24875,N_20505);
nor UO_2601 (O_2601,N_24347,N_22876);
nor UO_2602 (O_2602,N_24579,N_21936);
nand UO_2603 (O_2603,N_23773,N_24006);
nand UO_2604 (O_2604,N_20347,N_20054);
and UO_2605 (O_2605,N_21922,N_24920);
nand UO_2606 (O_2606,N_24603,N_20913);
nand UO_2607 (O_2607,N_21103,N_24488);
nor UO_2608 (O_2608,N_20842,N_22386);
nand UO_2609 (O_2609,N_20498,N_21743);
and UO_2610 (O_2610,N_24268,N_21236);
nor UO_2611 (O_2611,N_20050,N_21113);
nor UO_2612 (O_2612,N_22564,N_24323);
nand UO_2613 (O_2613,N_22878,N_24251);
and UO_2614 (O_2614,N_22091,N_22083);
and UO_2615 (O_2615,N_21325,N_21079);
nor UO_2616 (O_2616,N_22452,N_20061);
nor UO_2617 (O_2617,N_24708,N_23065);
or UO_2618 (O_2618,N_23023,N_23507);
or UO_2619 (O_2619,N_22483,N_21427);
and UO_2620 (O_2620,N_22275,N_23300);
or UO_2621 (O_2621,N_23203,N_23707);
or UO_2622 (O_2622,N_24942,N_24069);
or UO_2623 (O_2623,N_24983,N_21809);
and UO_2624 (O_2624,N_23045,N_24725);
nor UO_2625 (O_2625,N_20787,N_23536);
or UO_2626 (O_2626,N_23868,N_24602);
nor UO_2627 (O_2627,N_23698,N_24963);
nand UO_2628 (O_2628,N_24606,N_22302);
or UO_2629 (O_2629,N_24890,N_22351);
and UO_2630 (O_2630,N_24913,N_23892);
and UO_2631 (O_2631,N_20552,N_20076);
and UO_2632 (O_2632,N_24914,N_24259);
nand UO_2633 (O_2633,N_21566,N_21620);
or UO_2634 (O_2634,N_20209,N_20916);
nor UO_2635 (O_2635,N_22736,N_20704);
nand UO_2636 (O_2636,N_24872,N_24453);
or UO_2637 (O_2637,N_24493,N_20258);
and UO_2638 (O_2638,N_22052,N_21293);
nor UO_2639 (O_2639,N_24095,N_22692);
nand UO_2640 (O_2640,N_21671,N_23752);
or UO_2641 (O_2641,N_23217,N_24194);
and UO_2642 (O_2642,N_22035,N_23283);
or UO_2643 (O_2643,N_21392,N_21971);
or UO_2644 (O_2644,N_22182,N_23163);
and UO_2645 (O_2645,N_21329,N_23434);
nand UO_2646 (O_2646,N_20752,N_23148);
and UO_2647 (O_2647,N_21627,N_20389);
or UO_2648 (O_2648,N_21674,N_22134);
or UO_2649 (O_2649,N_20616,N_21724);
nand UO_2650 (O_2650,N_23294,N_20155);
or UO_2651 (O_2651,N_23396,N_22392);
and UO_2652 (O_2652,N_21593,N_24416);
nand UO_2653 (O_2653,N_23716,N_24382);
and UO_2654 (O_2654,N_22549,N_23359);
nor UO_2655 (O_2655,N_21764,N_21873);
nand UO_2656 (O_2656,N_24055,N_22217);
and UO_2657 (O_2657,N_24922,N_24855);
and UO_2658 (O_2658,N_21582,N_21434);
or UO_2659 (O_2659,N_23258,N_21500);
nand UO_2660 (O_2660,N_24777,N_20414);
or UO_2661 (O_2661,N_24436,N_22972);
nor UO_2662 (O_2662,N_21103,N_23264);
nand UO_2663 (O_2663,N_20928,N_21309);
nand UO_2664 (O_2664,N_20364,N_23930);
or UO_2665 (O_2665,N_20028,N_24708);
nand UO_2666 (O_2666,N_20597,N_23426);
nor UO_2667 (O_2667,N_24202,N_21423);
and UO_2668 (O_2668,N_21572,N_24581);
nand UO_2669 (O_2669,N_21958,N_21965);
and UO_2670 (O_2670,N_23836,N_22155);
nand UO_2671 (O_2671,N_23324,N_23856);
nand UO_2672 (O_2672,N_23340,N_24108);
nand UO_2673 (O_2673,N_20905,N_23954);
nor UO_2674 (O_2674,N_21588,N_24349);
nand UO_2675 (O_2675,N_20051,N_23536);
nand UO_2676 (O_2676,N_22061,N_24315);
nor UO_2677 (O_2677,N_23922,N_20979);
nor UO_2678 (O_2678,N_22718,N_22750);
nor UO_2679 (O_2679,N_24821,N_21334);
nand UO_2680 (O_2680,N_21522,N_24472);
nor UO_2681 (O_2681,N_20227,N_24102);
nand UO_2682 (O_2682,N_21701,N_23000);
or UO_2683 (O_2683,N_24956,N_24540);
and UO_2684 (O_2684,N_21809,N_22135);
nand UO_2685 (O_2685,N_22325,N_24795);
and UO_2686 (O_2686,N_20490,N_24484);
or UO_2687 (O_2687,N_21491,N_22298);
or UO_2688 (O_2688,N_21829,N_22745);
nor UO_2689 (O_2689,N_23818,N_20619);
or UO_2690 (O_2690,N_21255,N_24776);
or UO_2691 (O_2691,N_22034,N_24467);
and UO_2692 (O_2692,N_20235,N_20877);
nor UO_2693 (O_2693,N_23866,N_20439);
and UO_2694 (O_2694,N_24565,N_22610);
nand UO_2695 (O_2695,N_23887,N_22370);
or UO_2696 (O_2696,N_20948,N_21068);
nand UO_2697 (O_2697,N_24064,N_22198);
or UO_2698 (O_2698,N_22738,N_20230);
and UO_2699 (O_2699,N_20496,N_20388);
nand UO_2700 (O_2700,N_22259,N_21217);
and UO_2701 (O_2701,N_21451,N_20755);
or UO_2702 (O_2702,N_22729,N_21821);
or UO_2703 (O_2703,N_21200,N_23649);
or UO_2704 (O_2704,N_22647,N_24181);
nand UO_2705 (O_2705,N_20714,N_23520);
nand UO_2706 (O_2706,N_22305,N_24048);
xor UO_2707 (O_2707,N_21269,N_22888);
and UO_2708 (O_2708,N_22560,N_23941);
or UO_2709 (O_2709,N_22817,N_22941);
or UO_2710 (O_2710,N_22969,N_21776);
or UO_2711 (O_2711,N_21642,N_22305);
nor UO_2712 (O_2712,N_24204,N_23998);
and UO_2713 (O_2713,N_23503,N_22247);
or UO_2714 (O_2714,N_21982,N_21531);
nand UO_2715 (O_2715,N_24452,N_23420);
nand UO_2716 (O_2716,N_20569,N_22088);
and UO_2717 (O_2717,N_21974,N_24068);
nor UO_2718 (O_2718,N_23117,N_21835);
or UO_2719 (O_2719,N_21959,N_21940);
and UO_2720 (O_2720,N_20663,N_22228);
nor UO_2721 (O_2721,N_20671,N_20638);
and UO_2722 (O_2722,N_24368,N_20576);
nor UO_2723 (O_2723,N_24139,N_24009);
nor UO_2724 (O_2724,N_24315,N_24741);
or UO_2725 (O_2725,N_24842,N_22839);
nor UO_2726 (O_2726,N_24198,N_20811);
or UO_2727 (O_2727,N_20406,N_20740);
nor UO_2728 (O_2728,N_20892,N_21608);
and UO_2729 (O_2729,N_20210,N_20165);
nand UO_2730 (O_2730,N_22695,N_24820);
nand UO_2731 (O_2731,N_20290,N_21473);
or UO_2732 (O_2732,N_21606,N_21965);
and UO_2733 (O_2733,N_23533,N_24139);
and UO_2734 (O_2734,N_22391,N_22375);
or UO_2735 (O_2735,N_22153,N_21833);
nand UO_2736 (O_2736,N_24432,N_21966);
or UO_2737 (O_2737,N_22198,N_23118);
nand UO_2738 (O_2738,N_24122,N_24842);
or UO_2739 (O_2739,N_20018,N_20583);
nand UO_2740 (O_2740,N_23239,N_24127);
nor UO_2741 (O_2741,N_21623,N_23148);
nor UO_2742 (O_2742,N_24437,N_21729);
or UO_2743 (O_2743,N_22453,N_22020);
or UO_2744 (O_2744,N_23310,N_23606);
nand UO_2745 (O_2745,N_20112,N_21216);
nor UO_2746 (O_2746,N_22461,N_22614);
nand UO_2747 (O_2747,N_24290,N_20107);
nor UO_2748 (O_2748,N_24577,N_21557);
nor UO_2749 (O_2749,N_24956,N_22327);
or UO_2750 (O_2750,N_21117,N_21242);
or UO_2751 (O_2751,N_22165,N_22437);
or UO_2752 (O_2752,N_21612,N_24349);
xnor UO_2753 (O_2753,N_23545,N_24095);
nand UO_2754 (O_2754,N_20195,N_22641);
xor UO_2755 (O_2755,N_22969,N_22862);
nor UO_2756 (O_2756,N_21499,N_24182);
and UO_2757 (O_2757,N_22049,N_23267);
nor UO_2758 (O_2758,N_20305,N_24331);
nand UO_2759 (O_2759,N_23408,N_20946);
or UO_2760 (O_2760,N_22804,N_21067);
nor UO_2761 (O_2761,N_21583,N_23645);
or UO_2762 (O_2762,N_24399,N_24361);
nor UO_2763 (O_2763,N_23897,N_20981);
or UO_2764 (O_2764,N_20759,N_22439);
and UO_2765 (O_2765,N_20345,N_24444);
nor UO_2766 (O_2766,N_22145,N_22005);
nand UO_2767 (O_2767,N_21169,N_21246);
or UO_2768 (O_2768,N_21390,N_23697);
nand UO_2769 (O_2769,N_24022,N_24972);
nand UO_2770 (O_2770,N_21829,N_22198);
nand UO_2771 (O_2771,N_20034,N_20837);
nor UO_2772 (O_2772,N_20506,N_23451);
nand UO_2773 (O_2773,N_24297,N_23973);
and UO_2774 (O_2774,N_20472,N_22285);
or UO_2775 (O_2775,N_22754,N_22888);
nand UO_2776 (O_2776,N_20776,N_20941);
nand UO_2777 (O_2777,N_21218,N_20885);
or UO_2778 (O_2778,N_21379,N_22025);
nand UO_2779 (O_2779,N_20199,N_24481);
xor UO_2780 (O_2780,N_23517,N_22881);
nor UO_2781 (O_2781,N_21719,N_22730);
nand UO_2782 (O_2782,N_20668,N_23329);
nand UO_2783 (O_2783,N_22111,N_21071);
nand UO_2784 (O_2784,N_20810,N_23533);
nand UO_2785 (O_2785,N_21979,N_22374);
xor UO_2786 (O_2786,N_21164,N_24428);
nor UO_2787 (O_2787,N_24943,N_22974);
nand UO_2788 (O_2788,N_22160,N_22850);
or UO_2789 (O_2789,N_24896,N_23427);
or UO_2790 (O_2790,N_20318,N_21026);
nand UO_2791 (O_2791,N_23127,N_22734);
or UO_2792 (O_2792,N_21017,N_21266);
nor UO_2793 (O_2793,N_21724,N_24015);
nor UO_2794 (O_2794,N_22537,N_24318);
and UO_2795 (O_2795,N_22356,N_24303);
nor UO_2796 (O_2796,N_20574,N_21974);
nor UO_2797 (O_2797,N_22952,N_24034);
nor UO_2798 (O_2798,N_22288,N_23809);
nor UO_2799 (O_2799,N_21875,N_23128);
and UO_2800 (O_2800,N_23142,N_24978);
xor UO_2801 (O_2801,N_22032,N_23811);
xnor UO_2802 (O_2802,N_21037,N_21469);
and UO_2803 (O_2803,N_20352,N_24318);
nor UO_2804 (O_2804,N_21520,N_20256);
or UO_2805 (O_2805,N_23807,N_21954);
nor UO_2806 (O_2806,N_22534,N_21517);
xnor UO_2807 (O_2807,N_21746,N_22489);
nand UO_2808 (O_2808,N_22852,N_22022);
and UO_2809 (O_2809,N_21586,N_20370);
xnor UO_2810 (O_2810,N_21847,N_20950);
nand UO_2811 (O_2811,N_24771,N_23158);
or UO_2812 (O_2812,N_21267,N_23531);
and UO_2813 (O_2813,N_24527,N_22012);
or UO_2814 (O_2814,N_24925,N_23910);
and UO_2815 (O_2815,N_21903,N_22590);
nand UO_2816 (O_2816,N_21873,N_20156);
nand UO_2817 (O_2817,N_21336,N_20908);
or UO_2818 (O_2818,N_22073,N_20487);
or UO_2819 (O_2819,N_23226,N_24676);
and UO_2820 (O_2820,N_22469,N_23327);
nand UO_2821 (O_2821,N_23177,N_23323);
or UO_2822 (O_2822,N_20688,N_20908);
or UO_2823 (O_2823,N_24768,N_23434);
nand UO_2824 (O_2824,N_22406,N_23575);
and UO_2825 (O_2825,N_21759,N_21906);
nor UO_2826 (O_2826,N_20565,N_21027);
nand UO_2827 (O_2827,N_22500,N_24716);
nor UO_2828 (O_2828,N_24946,N_21752);
nand UO_2829 (O_2829,N_23105,N_20879);
nand UO_2830 (O_2830,N_22730,N_24369);
or UO_2831 (O_2831,N_21663,N_21530);
nand UO_2832 (O_2832,N_22063,N_22080);
or UO_2833 (O_2833,N_24139,N_23630);
nor UO_2834 (O_2834,N_24536,N_20507);
and UO_2835 (O_2835,N_23339,N_24240);
xor UO_2836 (O_2836,N_20562,N_20348);
or UO_2837 (O_2837,N_20905,N_20195);
nand UO_2838 (O_2838,N_21555,N_23891);
nand UO_2839 (O_2839,N_20251,N_20857);
nor UO_2840 (O_2840,N_20967,N_20829);
or UO_2841 (O_2841,N_22672,N_21274);
and UO_2842 (O_2842,N_21909,N_24274);
nor UO_2843 (O_2843,N_21137,N_22786);
and UO_2844 (O_2844,N_20345,N_23177);
nor UO_2845 (O_2845,N_23527,N_24826);
and UO_2846 (O_2846,N_23367,N_24728);
or UO_2847 (O_2847,N_24855,N_23482);
nand UO_2848 (O_2848,N_21604,N_24150);
or UO_2849 (O_2849,N_23150,N_21406);
nand UO_2850 (O_2850,N_22156,N_22455);
and UO_2851 (O_2851,N_22070,N_24283);
and UO_2852 (O_2852,N_21501,N_24216);
nor UO_2853 (O_2853,N_22166,N_24747);
or UO_2854 (O_2854,N_21840,N_23233);
and UO_2855 (O_2855,N_24298,N_22428);
nand UO_2856 (O_2856,N_21474,N_24433);
nor UO_2857 (O_2857,N_24093,N_23626);
or UO_2858 (O_2858,N_20486,N_21972);
nor UO_2859 (O_2859,N_21126,N_24907);
and UO_2860 (O_2860,N_20878,N_23444);
nand UO_2861 (O_2861,N_22741,N_20483);
nor UO_2862 (O_2862,N_22927,N_21033);
nor UO_2863 (O_2863,N_23235,N_21561);
nor UO_2864 (O_2864,N_23668,N_21005);
nand UO_2865 (O_2865,N_22125,N_20226);
and UO_2866 (O_2866,N_24409,N_22022);
or UO_2867 (O_2867,N_22297,N_20632);
or UO_2868 (O_2868,N_23331,N_22782);
and UO_2869 (O_2869,N_22171,N_20689);
nand UO_2870 (O_2870,N_23996,N_24709);
nor UO_2871 (O_2871,N_23673,N_24730);
nor UO_2872 (O_2872,N_21604,N_20260);
nand UO_2873 (O_2873,N_20182,N_24973);
or UO_2874 (O_2874,N_21908,N_21995);
and UO_2875 (O_2875,N_22045,N_23643);
nand UO_2876 (O_2876,N_21921,N_24656);
nor UO_2877 (O_2877,N_24816,N_23354);
and UO_2878 (O_2878,N_20458,N_22587);
and UO_2879 (O_2879,N_23410,N_22382);
nand UO_2880 (O_2880,N_22392,N_24427);
nand UO_2881 (O_2881,N_23225,N_23427);
nor UO_2882 (O_2882,N_21075,N_24636);
or UO_2883 (O_2883,N_23159,N_21602);
nand UO_2884 (O_2884,N_23750,N_22891);
and UO_2885 (O_2885,N_24332,N_22637);
nand UO_2886 (O_2886,N_20074,N_21018);
and UO_2887 (O_2887,N_23586,N_20210);
and UO_2888 (O_2888,N_20450,N_24040);
nand UO_2889 (O_2889,N_21166,N_20868);
and UO_2890 (O_2890,N_23882,N_22536);
nand UO_2891 (O_2891,N_24198,N_24244);
and UO_2892 (O_2892,N_20908,N_23122);
nand UO_2893 (O_2893,N_22499,N_22918);
xor UO_2894 (O_2894,N_22722,N_20808);
nand UO_2895 (O_2895,N_22814,N_24193);
or UO_2896 (O_2896,N_24389,N_22025);
nor UO_2897 (O_2897,N_21044,N_21506);
xor UO_2898 (O_2898,N_23082,N_21162);
nor UO_2899 (O_2899,N_23402,N_23892);
nor UO_2900 (O_2900,N_20084,N_24678);
nand UO_2901 (O_2901,N_21670,N_21916);
and UO_2902 (O_2902,N_21263,N_20900);
nand UO_2903 (O_2903,N_24567,N_24178);
nand UO_2904 (O_2904,N_23308,N_24830);
and UO_2905 (O_2905,N_24002,N_21531);
nor UO_2906 (O_2906,N_24490,N_24932);
and UO_2907 (O_2907,N_23588,N_21457);
or UO_2908 (O_2908,N_22861,N_21740);
and UO_2909 (O_2909,N_24531,N_23928);
or UO_2910 (O_2910,N_22967,N_23956);
and UO_2911 (O_2911,N_20435,N_23101);
or UO_2912 (O_2912,N_23271,N_21149);
nand UO_2913 (O_2913,N_20597,N_23350);
nor UO_2914 (O_2914,N_21645,N_23052);
nand UO_2915 (O_2915,N_21011,N_23526);
xnor UO_2916 (O_2916,N_20924,N_21971);
or UO_2917 (O_2917,N_22679,N_20436);
nor UO_2918 (O_2918,N_24242,N_22399);
and UO_2919 (O_2919,N_21815,N_20653);
and UO_2920 (O_2920,N_20910,N_24518);
xnor UO_2921 (O_2921,N_24756,N_20388);
and UO_2922 (O_2922,N_24255,N_22655);
or UO_2923 (O_2923,N_20854,N_22603);
and UO_2924 (O_2924,N_24901,N_20900);
and UO_2925 (O_2925,N_20827,N_20663);
nand UO_2926 (O_2926,N_22651,N_23043);
and UO_2927 (O_2927,N_24251,N_23113);
and UO_2928 (O_2928,N_21747,N_22017);
nor UO_2929 (O_2929,N_20009,N_20583);
nand UO_2930 (O_2930,N_20639,N_22173);
or UO_2931 (O_2931,N_22695,N_21537);
nor UO_2932 (O_2932,N_24634,N_24559);
nand UO_2933 (O_2933,N_21048,N_22043);
nor UO_2934 (O_2934,N_24054,N_23673);
or UO_2935 (O_2935,N_21093,N_21030);
nand UO_2936 (O_2936,N_20714,N_21173);
and UO_2937 (O_2937,N_21667,N_21047);
xor UO_2938 (O_2938,N_21264,N_24997);
and UO_2939 (O_2939,N_22181,N_21540);
nor UO_2940 (O_2940,N_21897,N_24016);
nor UO_2941 (O_2941,N_22128,N_23210);
nand UO_2942 (O_2942,N_20022,N_22209);
or UO_2943 (O_2943,N_20067,N_22470);
nand UO_2944 (O_2944,N_23833,N_21619);
xnor UO_2945 (O_2945,N_21410,N_20169);
nor UO_2946 (O_2946,N_20761,N_21329);
nor UO_2947 (O_2947,N_24764,N_21031);
nor UO_2948 (O_2948,N_20660,N_20680);
and UO_2949 (O_2949,N_24751,N_23492);
or UO_2950 (O_2950,N_22470,N_20153);
nor UO_2951 (O_2951,N_20796,N_21366);
and UO_2952 (O_2952,N_24986,N_22706);
and UO_2953 (O_2953,N_23517,N_23480);
nand UO_2954 (O_2954,N_24297,N_22952);
and UO_2955 (O_2955,N_22621,N_23444);
nand UO_2956 (O_2956,N_22989,N_24150);
nand UO_2957 (O_2957,N_21009,N_21420);
and UO_2958 (O_2958,N_21714,N_21017);
and UO_2959 (O_2959,N_20884,N_23278);
and UO_2960 (O_2960,N_21279,N_24624);
nor UO_2961 (O_2961,N_23673,N_20070);
and UO_2962 (O_2962,N_21465,N_24833);
or UO_2963 (O_2963,N_20034,N_22003);
nor UO_2964 (O_2964,N_24627,N_21136);
and UO_2965 (O_2965,N_20112,N_21668);
or UO_2966 (O_2966,N_23122,N_23028);
nor UO_2967 (O_2967,N_21443,N_21955);
and UO_2968 (O_2968,N_23598,N_23461);
nor UO_2969 (O_2969,N_22688,N_24156);
or UO_2970 (O_2970,N_23982,N_22329);
or UO_2971 (O_2971,N_24457,N_24809);
nand UO_2972 (O_2972,N_21187,N_21980);
nor UO_2973 (O_2973,N_22424,N_23243);
nor UO_2974 (O_2974,N_21120,N_23519);
nor UO_2975 (O_2975,N_23828,N_20524);
or UO_2976 (O_2976,N_20827,N_21803);
or UO_2977 (O_2977,N_21223,N_24159);
nand UO_2978 (O_2978,N_23034,N_20248);
or UO_2979 (O_2979,N_24070,N_23048);
or UO_2980 (O_2980,N_21628,N_20804);
nor UO_2981 (O_2981,N_23313,N_23607);
and UO_2982 (O_2982,N_23411,N_20989);
nand UO_2983 (O_2983,N_23101,N_21934);
xor UO_2984 (O_2984,N_23398,N_24279);
nand UO_2985 (O_2985,N_20569,N_23031);
xnor UO_2986 (O_2986,N_23381,N_22554);
and UO_2987 (O_2987,N_21869,N_22290);
and UO_2988 (O_2988,N_22135,N_22818);
nand UO_2989 (O_2989,N_24567,N_21144);
and UO_2990 (O_2990,N_24954,N_23395);
and UO_2991 (O_2991,N_24476,N_21026);
and UO_2992 (O_2992,N_23341,N_22829);
nor UO_2993 (O_2993,N_24209,N_21021);
and UO_2994 (O_2994,N_20935,N_24501);
xor UO_2995 (O_2995,N_22619,N_24381);
or UO_2996 (O_2996,N_23299,N_22137);
and UO_2997 (O_2997,N_20833,N_22748);
nor UO_2998 (O_2998,N_22381,N_23169);
nor UO_2999 (O_2999,N_22909,N_20804);
endmodule