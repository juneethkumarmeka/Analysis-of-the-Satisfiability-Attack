module basic_3000_30000_3500_25_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_434,In_639);
and U1 (N_1,In_86,In_2650);
nand U2 (N_2,In_2558,In_1457);
and U3 (N_3,In_657,In_2094);
and U4 (N_4,In_120,In_1323);
nor U5 (N_5,In_2127,In_502);
nor U6 (N_6,In_2122,In_167);
and U7 (N_7,In_2967,In_533);
xor U8 (N_8,In_364,In_209);
nand U9 (N_9,In_1612,In_1465);
nor U10 (N_10,In_2895,In_2853);
nor U11 (N_11,In_996,In_1657);
nor U12 (N_12,In_1091,In_340);
nand U13 (N_13,In_2433,In_741);
or U14 (N_14,In_1916,In_1039);
and U15 (N_15,In_1167,In_402);
and U16 (N_16,In_396,In_965);
nand U17 (N_17,In_1274,In_2364);
or U18 (N_18,In_1404,In_1893);
nand U19 (N_19,In_269,In_1829);
nor U20 (N_20,In_1576,In_174);
and U21 (N_21,In_688,In_2932);
nand U22 (N_22,In_1195,In_1765);
or U23 (N_23,In_1413,In_2004);
nor U24 (N_24,In_1368,In_2477);
nand U25 (N_25,In_419,In_2618);
nand U26 (N_26,In_2907,In_154);
nand U27 (N_27,In_2892,In_1611);
xnor U28 (N_28,In_2973,In_2472);
xor U29 (N_29,In_1444,In_2975);
and U30 (N_30,In_1494,In_1499);
and U31 (N_31,In_691,In_162);
or U32 (N_32,In_2214,In_1169);
or U33 (N_33,In_338,In_609);
nand U34 (N_34,In_508,In_2292);
nand U35 (N_35,In_816,In_481);
nand U36 (N_36,In_1172,In_1099);
nand U37 (N_37,In_1237,In_1985);
or U38 (N_38,In_760,In_2362);
or U39 (N_39,In_1939,In_2949);
nor U40 (N_40,In_1075,In_876);
nand U41 (N_41,In_1601,In_1745);
nand U42 (N_42,In_437,In_2185);
nand U43 (N_43,In_1786,In_737);
nor U44 (N_44,In_160,In_645);
nor U45 (N_45,In_904,In_1106);
xor U46 (N_46,In_656,In_539);
nor U47 (N_47,In_2116,In_1861);
or U48 (N_48,In_2587,In_266);
xnor U49 (N_49,In_715,In_2445);
nand U50 (N_50,In_1496,In_2675);
or U51 (N_51,In_834,In_2785);
or U52 (N_52,In_2888,In_673);
nand U53 (N_53,In_1770,In_1645);
nor U54 (N_54,In_633,In_1936);
nand U55 (N_55,In_545,In_998);
xor U56 (N_56,In_1729,In_1535);
and U57 (N_57,In_1986,In_446);
xnor U58 (N_58,In_18,In_8);
or U59 (N_59,In_333,In_662);
nor U60 (N_60,In_1026,In_2653);
and U61 (N_61,In_2134,In_507);
or U62 (N_62,In_1699,In_2673);
and U63 (N_63,In_1799,In_2055);
and U64 (N_64,In_1683,In_2464);
and U65 (N_65,In_1831,In_295);
and U66 (N_66,In_2099,In_125);
nor U67 (N_67,In_2304,In_359);
nor U68 (N_68,In_27,In_2542);
or U69 (N_69,In_2953,In_923);
xnor U70 (N_70,In_2746,In_1805);
or U71 (N_71,In_2103,In_2409);
nand U72 (N_72,In_2868,In_2818);
xor U73 (N_73,In_2490,In_58);
or U74 (N_74,In_1910,In_202);
nand U75 (N_75,In_2500,In_1079);
nor U76 (N_76,In_2148,In_728);
or U77 (N_77,In_1782,In_627);
nand U78 (N_78,In_726,In_2206);
nand U79 (N_79,In_98,In_2337);
or U80 (N_80,In_186,In_2905);
nor U81 (N_81,In_2549,In_2531);
nand U82 (N_82,In_599,In_2767);
nand U83 (N_83,In_577,In_999);
nor U84 (N_84,In_82,In_1084);
nand U85 (N_85,In_2093,In_2526);
or U86 (N_86,In_2072,In_879);
nor U87 (N_87,In_2832,In_1081);
nor U88 (N_88,In_2515,In_2312);
and U89 (N_89,In_1027,In_2846);
nand U90 (N_90,In_2488,In_1727);
nor U91 (N_91,In_1913,In_2585);
or U92 (N_92,In_714,In_975);
nand U93 (N_93,In_1788,In_518);
or U94 (N_94,In_2961,In_1955);
nand U95 (N_95,In_1684,In_808);
nor U96 (N_96,In_2437,In_795);
nor U97 (N_97,In_410,In_946);
nand U98 (N_98,In_2682,In_1073);
and U99 (N_99,In_1545,In_1232);
xnor U100 (N_100,In_399,In_1255);
xor U101 (N_101,In_487,In_351);
nor U102 (N_102,In_14,In_643);
xnor U103 (N_103,In_818,In_2513);
nor U104 (N_104,In_745,In_145);
and U105 (N_105,In_1031,In_2624);
xnor U106 (N_106,In_575,In_146);
and U107 (N_107,In_2229,In_981);
nor U108 (N_108,In_2797,In_43);
nand U109 (N_109,In_1108,In_2352);
nand U110 (N_110,In_2897,In_2271);
and U111 (N_111,In_1627,In_699);
nand U112 (N_112,In_1453,In_135);
xnor U113 (N_113,In_2788,In_2849);
nor U114 (N_114,In_1988,In_2984);
nand U115 (N_115,In_227,In_1762);
and U116 (N_116,In_2997,In_391);
nand U117 (N_117,In_225,In_592);
nor U118 (N_118,In_136,In_1262);
and U119 (N_119,In_2732,In_867);
xnor U120 (N_120,In_1514,In_2043);
nor U121 (N_121,In_652,In_881);
and U122 (N_122,In_1168,In_704);
nor U123 (N_123,In_980,In_2610);
or U124 (N_124,In_886,In_1830);
or U125 (N_125,In_1191,In_649);
and U126 (N_126,In_2783,In_378);
xnor U127 (N_127,In_1933,In_2728);
xnor U128 (N_128,In_233,In_2354);
nor U129 (N_129,In_598,In_2212);
nand U130 (N_130,In_460,In_1358);
nand U131 (N_131,In_1275,In_2082);
or U132 (N_132,In_189,In_2272);
nand U133 (N_133,In_517,In_1259);
xnor U134 (N_134,In_806,In_1973);
nor U135 (N_135,In_2369,In_2149);
and U136 (N_136,In_2405,In_170);
xnor U137 (N_137,In_1235,In_1481);
nand U138 (N_138,In_1726,In_1780);
or U139 (N_139,In_273,In_1490);
nor U140 (N_140,In_667,In_1510);
nand U141 (N_141,In_55,In_318);
xnor U142 (N_142,In_458,In_485);
nand U143 (N_143,In_612,In_566);
xor U144 (N_144,In_2224,In_1523);
nand U145 (N_145,In_1998,In_815);
or U146 (N_146,In_1568,In_81);
or U147 (N_147,In_2373,In_105);
xnor U148 (N_148,In_376,In_2681);
nor U149 (N_149,In_2139,In_917);
or U150 (N_150,In_89,In_2592);
or U151 (N_151,In_898,In_2484);
or U152 (N_152,In_2864,In_231);
or U153 (N_153,In_1258,In_2940);
nand U154 (N_154,In_187,In_672);
or U155 (N_155,In_634,In_4);
and U156 (N_156,In_83,In_1128);
xnor U157 (N_157,In_2883,In_1133);
or U158 (N_158,In_441,In_885);
nand U159 (N_159,In_669,In_2309);
xnor U160 (N_160,In_640,In_860);
xnor U161 (N_161,In_2316,In_552);
and U162 (N_162,In_1327,In_1375);
xor U163 (N_163,In_2138,In_2978);
and U164 (N_164,In_1739,In_2548);
nand U165 (N_165,In_286,In_2467);
and U166 (N_166,In_2482,In_2088);
nand U167 (N_167,In_2614,In_1025);
nor U168 (N_168,In_268,In_1418);
xnor U169 (N_169,In_254,In_2648);
xor U170 (N_170,In_1390,In_1000);
and U171 (N_171,In_1855,In_176);
xor U172 (N_172,In_1975,In_573);
or U173 (N_173,In_248,In_727);
nand U174 (N_174,In_931,In_793);
nand U175 (N_175,In_2249,In_1456);
or U176 (N_176,In_2104,In_2401);
nor U177 (N_177,In_2957,In_2635);
and U178 (N_178,In_2711,In_1342);
nor U179 (N_179,In_2047,In_2236);
or U180 (N_180,In_474,In_319);
xor U181 (N_181,In_814,In_2036);
or U182 (N_182,In_2399,In_1159);
nor U183 (N_183,In_758,In_2434);
and U184 (N_184,In_2349,In_828);
nand U185 (N_185,In_190,In_213);
and U186 (N_186,In_2486,In_2680);
nand U187 (N_187,In_973,In_1316);
and U188 (N_188,In_2903,In_1093);
xor U189 (N_189,In_514,In_2360);
and U190 (N_190,In_986,In_1953);
nor U191 (N_191,In_361,In_661);
or U192 (N_192,In_1595,In_2422);
xnor U193 (N_193,In_2649,In_1468);
xor U194 (N_194,In_2428,In_491);
nor U195 (N_195,In_835,In_2729);
and U196 (N_196,In_1277,In_2956);
nor U197 (N_197,In_1440,In_2756);
xnor U198 (N_198,In_1814,In_1567);
and U199 (N_199,In_2964,In_2935);
or U200 (N_200,In_841,In_937);
and U201 (N_201,In_2654,In_698);
nand U202 (N_202,In_2076,In_2306);
or U203 (N_203,In_520,In_1541);
nor U204 (N_204,In_2386,In_2628);
and U205 (N_205,In_450,In_1543);
and U206 (N_206,In_1615,In_984);
nand U207 (N_207,In_1878,In_2520);
nand U208 (N_208,In_1151,In_2987);
nand U209 (N_209,In_920,In_2252);
xnor U210 (N_210,In_2740,In_1113);
nor U211 (N_211,In_2462,In_1822);
nand U212 (N_212,In_194,In_321);
nor U213 (N_213,In_582,In_2198);
nor U214 (N_214,In_742,In_2992);
xor U215 (N_215,In_2166,In_792);
nor U216 (N_216,In_2847,In_433);
xnor U217 (N_217,In_2131,In_1532);
xor U218 (N_218,In_436,In_1055);
nand U219 (N_219,In_710,In_2263);
nor U220 (N_220,In_2000,In_1748);
or U221 (N_221,In_199,In_439);
or U222 (N_222,In_356,In_1386);
or U223 (N_223,In_2400,In_1944);
nor U224 (N_224,In_1226,In_1322);
nand U225 (N_225,In_2046,In_1520);
and U226 (N_226,In_991,In_944);
xnor U227 (N_227,In_2742,In_1420);
xor U228 (N_228,In_90,In_469);
nand U229 (N_229,In_1759,In_972);
xor U230 (N_230,In_2315,In_1573);
and U231 (N_231,In_1124,In_2516);
nand U232 (N_232,In_1890,In_1790);
and U233 (N_233,In_707,In_2078);
xor U234 (N_234,In_153,In_1847);
or U235 (N_235,In_1253,In_771);
xnor U236 (N_236,In_572,In_2473);
or U237 (N_237,In_671,In_1341);
nor U238 (N_238,In_137,In_994);
xor U239 (N_239,In_1455,In_467);
or U240 (N_240,In_1003,In_1330);
xor U241 (N_241,In_932,In_2596);
or U242 (N_242,In_322,In_493);
nor U243 (N_243,In_1302,In_635);
nor U244 (N_244,In_1584,In_49);
nand U245 (N_245,In_2511,In_1837);
and U246 (N_246,In_2408,In_1071);
xor U247 (N_247,In_964,In_1929);
and U248 (N_248,In_1451,In_790);
or U249 (N_249,In_264,In_2253);
or U250 (N_250,In_1834,In_1571);
and U251 (N_251,In_1065,In_1853);
or U252 (N_252,In_2660,In_1283);
and U253 (N_253,In_859,In_1845);
nand U254 (N_254,In_550,In_1279);
nor U255 (N_255,In_1742,In_234);
xnor U256 (N_256,In_345,In_2027);
or U257 (N_257,In_1648,In_463);
or U258 (N_258,In_2572,In_1044);
and U259 (N_259,In_1266,In_1981);
or U260 (N_260,In_509,In_1131);
nor U261 (N_261,In_247,In_2506);
nand U262 (N_262,In_1098,In_384);
nand U263 (N_263,In_2522,In_1807);
nor U264 (N_264,In_625,In_7);
and U265 (N_265,In_1697,In_2630);
nand U266 (N_266,In_259,In_2279);
and U267 (N_267,In_2418,In_1422);
or U268 (N_268,In_587,In_1392);
xnor U269 (N_269,In_1057,In_921);
nand U270 (N_270,In_2151,In_432);
and U271 (N_271,In_1558,In_59);
and U272 (N_272,In_2861,In_602);
xnor U273 (N_273,In_2189,In_60);
or U274 (N_274,In_1175,In_1459);
nor U275 (N_275,In_1118,In_1629);
nor U276 (N_276,In_1951,In_41);
nor U277 (N_277,In_855,In_72);
xor U278 (N_278,In_1467,In_2708);
xnor U279 (N_279,In_2208,In_342);
nand U280 (N_280,In_1889,In_1579);
nand U281 (N_281,In_918,In_2331);
and U282 (N_282,In_1556,In_1803);
nor U283 (N_283,In_2375,In_2085);
xnor U284 (N_284,In_2620,In_2750);
and U285 (N_285,In_2938,In_2102);
and U286 (N_286,In_1092,In_130);
nand U287 (N_287,In_2403,In_2246);
nor U288 (N_288,In_988,In_181);
nor U289 (N_289,In_486,In_119);
nand U290 (N_290,In_2398,In_772);
or U291 (N_291,In_2743,In_974);
nor U292 (N_292,In_71,In_896);
or U293 (N_293,In_1518,In_1512);
nand U294 (N_294,In_2985,In_2053);
xnor U295 (N_295,In_279,In_723);
xnor U296 (N_296,In_258,In_719);
nor U297 (N_297,In_884,In_1306);
xnor U298 (N_298,In_1136,In_1329);
nand U299 (N_299,In_2640,In_2901);
nand U300 (N_300,In_1557,In_736);
and U301 (N_301,In_1754,In_650);
or U302 (N_302,In_2319,In_2597);
nor U303 (N_303,In_2947,In_597);
and U304 (N_304,In_2095,In_2633);
xor U305 (N_305,In_1626,In_797);
or U306 (N_306,In_1117,In_159);
xor U307 (N_307,In_541,In_214);
nor U308 (N_308,In_516,In_1032);
nand U309 (N_309,In_20,In_1605);
and U310 (N_310,In_1993,In_2722);
nand U311 (N_311,In_1243,In_1236);
or U312 (N_312,In_217,In_725);
nand U313 (N_313,In_2251,In_2211);
nand U314 (N_314,In_1315,In_1711);
xnor U315 (N_315,In_1554,In_966);
xnor U316 (N_316,In_1529,In_561);
nand U317 (N_317,In_600,In_349);
or U318 (N_318,In_2824,In_524);
and U319 (N_319,In_1210,In_2672);
or U320 (N_320,In_1524,In_1408);
and U321 (N_321,In_1434,In_1307);
and U322 (N_322,In_761,In_1562);
and U323 (N_323,In_1876,In_1066);
xor U324 (N_324,In_1602,In_1013);
nand U325 (N_325,In_428,In_950);
nand U326 (N_326,In_1284,In_1298);
nor U327 (N_327,In_1694,In_2946);
or U328 (N_328,In_2790,In_2264);
nand U329 (N_329,In_2805,In_236);
or U330 (N_330,In_2782,In_1);
nor U331 (N_331,In_1990,In_2770);
or U332 (N_332,In_832,In_1396);
or U333 (N_333,In_499,In_894);
or U334 (N_334,In_1723,In_2871);
nor U335 (N_335,In_1129,In_1380);
and U336 (N_336,In_1812,In_132);
nand U337 (N_337,In_1549,In_1139);
xor U338 (N_338,In_2744,In_2210);
and U339 (N_339,In_440,In_74);
xnor U340 (N_340,In_564,In_2643);
or U341 (N_341,In_2730,In_2658);
nand U342 (N_342,In_1049,In_1426);
or U343 (N_343,In_1779,In_1692);
nand U344 (N_344,In_748,In_2110);
and U345 (N_345,In_2801,In_2071);
nand U346 (N_346,In_603,In_2245);
or U347 (N_347,In_2813,In_1351);
nor U348 (N_348,In_1888,In_2158);
or U349 (N_349,In_2645,In_1920);
nand U350 (N_350,In_1992,In_2809);
or U351 (N_351,In_2735,In_261);
xor U352 (N_352,In_2145,In_91);
and U353 (N_353,In_117,In_1760);
nand U354 (N_354,In_1511,In_489);
and U355 (N_355,In_2615,In_2923);
nor U356 (N_356,In_854,In_1379);
or U357 (N_357,In_680,In_2142);
and U358 (N_358,In_2005,In_352);
nor U359 (N_359,In_705,In_1968);
and U360 (N_360,In_1526,In_2494);
nand U361 (N_361,In_2980,In_2820);
xnor U362 (N_362,In_2642,In_940);
xnor U363 (N_363,In_2882,In_888);
nor U364 (N_364,In_1181,In_1371);
nand U365 (N_365,In_449,In_1116);
xor U366 (N_366,In_969,In_850);
nand U367 (N_367,In_822,In_15);
nand U368 (N_368,In_2705,In_2666);
nor U369 (N_369,In_2285,In_1718);
nand U370 (N_370,In_2350,In_1881);
xor U371 (N_371,In_873,In_17);
or U372 (N_372,In_2474,In_2411);
nor U373 (N_373,In_1634,In_1623);
xor U374 (N_374,In_1449,In_2108);
nand U375 (N_375,In_1078,In_1209);
nand U376 (N_376,In_185,In_1400);
xor U377 (N_377,In_694,In_1502);
nor U378 (N_378,In_2452,In_475);
xor U379 (N_379,In_968,In_911);
or U380 (N_380,In_1841,In_2583);
nand U381 (N_381,In_1197,In_1192);
nor U382 (N_382,In_37,In_2389);
nor U383 (N_383,In_1710,In_1072);
or U384 (N_384,In_954,In_1397);
nor U385 (N_385,In_274,In_1264);
or U386 (N_386,In_872,In_2217);
nand U387 (N_387,In_1208,In_2764);
nor U388 (N_388,In_2268,In_2812);
xnor U389 (N_389,In_293,In_2387);
xor U390 (N_390,In_2769,In_1163);
or U391 (N_391,In_2124,In_1184);
nand U392 (N_392,In_1970,In_2977);
or U393 (N_393,In_256,In_2966);
and U394 (N_394,In_1649,In_1646);
nand U395 (N_395,In_2107,In_2616);
xor U396 (N_396,In_1087,In_1176);
nor U397 (N_397,In_651,In_2427);
xor U398 (N_398,In_2365,In_1707);
xnor U399 (N_399,In_362,In_2657);
xnor U400 (N_400,In_2146,In_2848);
nor U401 (N_401,In_1155,In_1314);
and U402 (N_402,In_1771,In_2738);
nor U403 (N_403,In_1525,In_1503);
xor U404 (N_404,In_1317,In_2699);
nand U405 (N_405,In_2761,In_594);
nand U406 (N_406,In_2174,In_682);
nor U407 (N_407,In_2242,In_2412);
and U408 (N_408,In_1842,In_2248);
or U409 (N_409,In_1289,In_2070);
nor U410 (N_410,In_1187,In_1189);
xor U411 (N_411,In_1915,In_2567);
nor U412 (N_412,In_1714,In_1661);
nand U413 (N_413,In_265,In_512);
xor U414 (N_414,In_1585,In_2521);
nand U415 (N_415,In_501,In_1185);
or U416 (N_416,In_654,In_1958);
or U417 (N_417,In_2589,In_2033);
nand U418 (N_418,In_2209,In_1703);
and U419 (N_419,In_1717,In_607);
nor U420 (N_420,In_329,In_2836);
nor U421 (N_421,In_947,In_567);
nand U422 (N_422,In_2686,In_1002);
nand U423 (N_423,In_2752,In_1923);
xor U424 (N_424,In_906,In_608);
nor U425 (N_425,In_1040,In_1539);
and U426 (N_426,In_1828,In_1460);
and U427 (N_427,In_257,In_398);
nand U428 (N_428,In_2269,In_2918);
nand U429 (N_429,In_2425,In_2646);
or U430 (N_430,In_1464,In_942);
nor U431 (N_431,In_2188,In_341);
nand U432 (N_432,In_1276,In_833);
xnor U433 (N_433,In_1885,In_1220);
xnor U434 (N_434,In_1359,In_1416);
nand U435 (N_435,In_2243,In_1486);
or U436 (N_436,In_2493,In_1205);
nor U437 (N_437,In_2376,In_2822);
nand U438 (N_438,In_365,In_2974);
xor U439 (N_439,In_1731,In_1211);
nand U440 (N_440,In_2310,In_313);
and U441 (N_441,In_2579,In_2704);
or U442 (N_442,In_2419,In_2546);
or U443 (N_443,In_2540,In_2697);
xnor U444 (N_444,In_2969,In_716);
xor U445 (N_445,In_2713,In_1686);
and U446 (N_446,In_1493,In_2690);
nand U447 (N_447,In_1778,In_142);
xnor U448 (N_448,In_44,In_251);
and U449 (N_449,In_1665,In_5);
xor U450 (N_450,In_675,In_1100);
or U451 (N_451,In_683,In_1527);
or U452 (N_452,In_2225,In_1393);
xnor U453 (N_453,In_464,In_1917);
nand U454 (N_454,In_1569,In_2451);
and U455 (N_455,In_2431,In_735);
nor U456 (N_456,In_2678,In_1042);
xor U457 (N_457,In_1934,In_570);
and U458 (N_458,In_122,In_2265);
and U459 (N_459,In_1119,In_2458);
or U460 (N_460,In_646,In_381);
nor U461 (N_461,In_2695,In_2609);
and U462 (N_462,In_1685,In_1733);
xor U463 (N_463,In_579,In_591);
nand U464 (N_464,In_1469,In_1918);
and U465 (N_465,In_1265,In_1946);
or U466 (N_466,In_2677,In_2982);
nand U467 (N_467,In_1983,In_13);
nand U468 (N_468,In_112,In_703);
nor U469 (N_469,In_2867,In_1991);
xnor U470 (N_470,In_116,In_2361);
nand U471 (N_471,In_2016,In_2150);
nand U472 (N_472,In_2416,In_802);
or U473 (N_473,In_865,In_413);
nand U474 (N_474,In_35,In_1294);
or U475 (N_475,In_2731,In_1901);
or U476 (N_476,In_25,In_2232);
xnor U477 (N_477,In_2556,In_763);
and U478 (N_478,In_2012,In_337);
and U479 (N_479,In_1679,In_216);
and U480 (N_480,In_2886,In_2712);
or U481 (N_481,In_2578,In_1840);
xor U482 (N_482,In_1508,In_457);
or U483 (N_483,In_2636,In_708);
xnor U484 (N_484,In_853,In_168);
xnor U485 (N_485,In_220,In_1883);
nor U486 (N_486,In_1793,In_2955);
or U487 (N_487,In_2340,In_871);
nor U488 (N_488,In_526,In_2314);
and U489 (N_489,In_851,In_2240);
or U490 (N_490,In_848,In_1221);
nor U491 (N_491,In_2837,In_1482);
and U492 (N_492,In_241,In_803);
xnor U493 (N_493,In_644,In_1096);
or U494 (N_494,In_1326,In_1773);
or U495 (N_495,In_243,In_2167);
nand U496 (N_496,In_1001,In_2497);
and U497 (N_497,In_2739,In_431);
nand U498 (N_498,In_2890,In_2062);
xnor U499 (N_499,In_2880,In_369);
or U500 (N_500,In_47,In_200);
and U501 (N_501,In_239,In_201);
nor U502 (N_502,In_1257,In_1705);
or U503 (N_503,In_2178,In_197);
xor U504 (N_504,In_2835,In_204);
xor U505 (N_505,In_1154,In_1083);
nand U506 (N_506,In_12,In_1304);
and U507 (N_507,In_2988,In_1862);
nor U508 (N_508,In_863,In_1835);
nor U509 (N_509,In_2204,In_532);
xnor U510 (N_510,In_1170,In_180);
and U511 (N_511,In_2024,In_1141);
xnor U512 (N_512,In_2492,In_2057);
nor U513 (N_513,In_1349,In_2118);
nand U514 (N_514,In_2329,In_2569);
and U515 (N_515,In_2727,In_1688);
nor U516 (N_516,In_1638,In_1140);
xnor U517 (N_517,In_1162,In_770);
nor U518 (N_518,In_1412,In_93);
nor U519 (N_519,In_902,In_1147);
or U520 (N_520,In_796,In_2481);
xor U521 (N_521,In_2760,In_1942);
xnor U522 (N_522,In_355,In_2254);
nand U523 (N_523,In_595,In_179);
nor U524 (N_524,In_1012,In_1965);
nor U525 (N_525,In_729,In_1053);
xnor U526 (N_526,In_1409,In_1617);
or U527 (N_527,In_52,In_115);
and U528 (N_528,In_2220,In_2898);
and U529 (N_529,In_108,In_1407);
or U530 (N_530,In_1492,In_2367);
nor U531 (N_531,In_2745,In_470);
nor U532 (N_532,In_1473,In_2466);
nor U533 (N_533,In_2090,In_2165);
nor U534 (N_534,In_1063,In_1956);
xor U535 (N_535,In_1590,In_237);
xor U536 (N_536,In_2120,In_1364);
xnor U537 (N_537,In_306,In_1747);
nand U538 (N_538,In_2436,In_2470);
xnor U539 (N_539,In_2584,In_141);
nor U540 (N_540,In_1248,In_842);
xnor U541 (N_541,In_334,In_22);
nor U542 (N_542,In_270,In_1443);
nand U543 (N_543,In_971,In_2372);
or U544 (N_544,In_2344,In_331);
xor U545 (N_545,In_659,In_63);
or U546 (N_546,In_2152,In_1383);
or U547 (N_547,In_2018,In_647);
nor U548 (N_548,In_2504,In_1781);
nand U549 (N_549,In_2469,In_2663);
nor U550 (N_550,In_2202,In_372);
and U551 (N_551,In_2833,In_2244);
and U552 (N_552,In_2719,In_1600);
xor U553 (N_553,In_1452,In_2623);
nand U554 (N_554,In_2963,In_78);
and U555 (N_555,In_590,In_1662);
or U556 (N_556,In_2056,In_2595);
nor U557 (N_557,In_2830,In_1241);
or U558 (N_558,In_858,In_416);
nor U559 (N_559,In_547,In_2689);
and U560 (N_560,In_11,In_2662);
xnor U561 (N_561,In_2190,In_459);
xnor U562 (N_562,In_836,In_1997);
and U563 (N_563,In_1839,In_2562);
xor U564 (N_564,In_990,In_1150);
nand U565 (N_565,In_2866,In_549);
xor U566 (N_566,In_2064,In_303);
xor U567 (N_567,In_448,In_1219);
or U568 (N_568,In_963,In_676);
xor U569 (N_569,In_2280,In_150);
or U570 (N_570,In_2774,In_314);
or U571 (N_571,In_2748,In_987);
or U572 (N_572,In_2200,In_2463);
or U573 (N_573,In_212,In_2100);
nor U574 (N_574,In_619,In_128);
nor U575 (N_575,In_235,In_184);
and U576 (N_576,In_1332,In_42);
xnor U577 (N_577,In_1271,In_2395);
nand U578 (N_578,In_2561,In_2536);
xor U579 (N_579,In_505,In_1149);
nor U580 (N_580,In_2577,In_2336);
and U581 (N_581,In_2906,In_272);
nand U582 (N_582,In_110,In_1826);
and U583 (N_583,In_2996,In_468);
xor U584 (N_584,In_2889,In_2358);
nor U585 (N_585,In_2574,In_1033);
and U586 (N_586,In_1614,In_542);
nor U587 (N_587,In_995,In_1374);
nor U588 (N_588,In_2277,In_613);
and U589 (N_589,In_1869,In_928);
nor U590 (N_590,In_1706,In_1886);
nand U591 (N_591,In_1045,In_94);
xor U592 (N_592,In_218,In_1156);
and U593 (N_593,In_406,In_2363);
or U594 (N_594,In_2845,In_878);
nand U595 (N_595,In_936,In_377);
xor U596 (N_596,In_1994,In_2530);
xnor U597 (N_597,In_2951,In_2573);
and U598 (N_598,In_1547,In_260);
or U599 (N_599,In_350,In_23);
nor U600 (N_600,In_1308,In_1971);
or U601 (N_601,In_2478,In_2479);
nor U602 (N_602,In_1967,In_1125);
or U603 (N_603,In_1318,In_840);
nand U604 (N_604,In_2929,In_2551);
nor U605 (N_605,In_1378,In_1596);
nand U606 (N_606,In_1491,In_2241);
nand U607 (N_607,In_1566,In_1143);
or U608 (N_608,In_2130,In_1937);
nor U609 (N_609,In_1586,In_1103);
and U610 (N_610,In_305,In_171);
nand U611 (N_611,In_2667,In_623);
or U612 (N_612,In_638,In_483);
nor U613 (N_613,In_1836,In_862);
or U614 (N_614,In_755,In_1598);
nand U615 (N_615,In_1722,In_2215);
nor U616 (N_616,In_480,In_2817);
nand U617 (N_617,In_1043,In_2273);
nor U618 (N_618,In_941,In_2135);
and U619 (N_619,In_2112,In_1630);
and U620 (N_620,In_442,In_2948);
and U621 (N_621,In_788,In_371);
or U622 (N_622,In_1873,In_456);
or U623 (N_623,In_208,In_2570);
and U624 (N_624,In_1070,In_2958);
nand U625 (N_625,In_540,In_1670);
and U626 (N_626,In_2390,In_435);
xnor U627 (N_627,In_2096,In_812);
and U628 (N_628,In_961,In_2223);
nor U629 (N_629,In_2059,In_148);
xnor U630 (N_630,In_1682,In_9);
or U631 (N_631,In_712,In_2067);
nor U632 (N_632,In_1391,In_1769);
nor U633 (N_633,In_1047,In_2017);
xor U634 (N_634,In_1238,In_1776);
and U635 (N_635,In_1442,In_462);
or U636 (N_636,In_2588,In_1796);
nand U637 (N_637,In_1709,In_1216);
or U638 (N_638,In_2421,In_2457);
nand U639 (N_639,In_1182,In_632);
xnor U640 (N_640,In_2345,In_374);
nor U641 (N_641,In_622,In_1427);
nor U642 (N_642,In_1887,In_2776);
nand U643 (N_643,In_2916,In_1758);
nand U644 (N_644,In_776,In_2828);
xnor U645 (N_645,In_282,In_1107);
and U646 (N_646,In_717,In_2438);
nor U647 (N_647,In_1059,In_530);
and U648 (N_648,In_388,In_73);
and U649 (N_649,In_1144,In_1287);
nand U650 (N_650,In_2844,In_230);
xnor U651 (N_651,In_1009,In_821);
and U652 (N_652,In_2607,In_756);
nand U653 (N_653,In_2299,In_2608);
and U654 (N_654,In_1201,In_738);
nand U655 (N_655,In_2983,In_2839);
nand U656 (N_656,In_2850,In_2909);
nor U657 (N_657,In_1345,In_2454);
and U658 (N_658,In_2709,In_2625);
and U659 (N_659,In_1651,In_1179);
nand U660 (N_660,In_750,In_500);
nand U661 (N_661,In_686,In_407);
or U662 (N_662,In_1178,In_2307);
or U663 (N_663,In_2296,In_79);
or U664 (N_664,In_263,In_1112);
xnor U665 (N_665,In_1305,In_2525);
and U666 (N_666,In_2734,In_1218);
xnor U667 (N_667,In_2485,In_165);
or U668 (N_668,In_1787,In_2334);
and U669 (N_669,In_781,In_2619);
and U670 (N_670,In_1616,In_1884);
or U671 (N_671,In_1738,In_513);
nand U672 (N_672,In_1104,In_585);
nand U673 (N_673,In_1736,In_2971);
or U674 (N_674,In_2865,In_2159);
and U675 (N_675,In_2544,In_1454);
nand U676 (N_676,In_1363,In_198);
xor U677 (N_677,In_1852,In_1485);
nand U678 (N_678,In_1015,In_2054);
and U679 (N_679,In_629,In_2355);
or U680 (N_680,In_2718,In_553);
or U681 (N_681,In_967,In_1249);
and U682 (N_682,In_1680,In_267);
nor U683 (N_683,In_417,In_611);
or U684 (N_684,In_794,In_2388);
xor U685 (N_685,In_1746,In_2449);
and U686 (N_686,In_767,In_222);
xnor U687 (N_687,In_785,In_245);
nand U688 (N_688,In_2787,In_370);
nand U689 (N_689,In_1222,In_1476);
and U690 (N_690,In_1439,In_1328);
nand U691 (N_691,In_2972,In_2058);
xor U692 (N_692,In_2396,In_2203);
nand U693 (N_693,In_670,In_1406);
or U694 (N_694,In_1763,In_2133);
and U695 (N_695,In_2317,In_2301);
or U696 (N_696,In_1048,In_1982);
or U697 (N_697,In_825,In_1797);
nor U698 (N_698,In_2523,In_126);
and U699 (N_699,In_1522,In_2275);
or U700 (N_700,In_476,In_702);
nand U701 (N_701,In_1011,In_2930);
and U702 (N_702,In_67,In_1252);
or U703 (N_703,In_948,In_1980);
xnor U704 (N_704,In_461,In_856);
and U705 (N_705,In_1618,In_1902);
nor U706 (N_706,In_2392,In_138);
xor U707 (N_707,In_1344,In_477);
and U708 (N_708,In_1824,In_1200);
nor U709 (N_709,In_866,In_2305);
or U710 (N_710,In_621,In_1632);
or U711 (N_711,In_466,In_1542);
nor U712 (N_712,In_583,In_1435);
nand U713 (N_713,In_899,In_2637);
or U714 (N_714,In_1589,In_2656);
nor U715 (N_715,In_2716,In_300);
nand U716 (N_716,In_2063,In_2164);
nand U717 (N_717,In_1006,In_1483);
nand U718 (N_718,In_1250,In_1050);
xnor U719 (N_719,In_1817,In_1740);
and U720 (N_720,In_164,In_1984);
nand U721 (N_721,In_926,In_711);
and U722 (N_722,In_809,In_747);
or U723 (N_723,In_2563,In_54);
or U724 (N_724,In_1134,In_1534);
xnor U725 (N_725,In_2904,In_1863);
nor U726 (N_726,In_1681,In_2181);
and U727 (N_727,In_1766,In_443);
xnor U728 (N_728,In_111,In_2207);
and U729 (N_729,In_789,In_1952);
xor U730 (N_730,In_2586,In_1833);
or U731 (N_731,In_1676,In_1548);
nand U732 (N_732,In_1035,In_38);
or U733 (N_733,In_1577,In_891);
and U734 (N_734,In_957,In_2924);
and U735 (N_735,In_956,In_2233);
xnor U736 (N_736,In_1528,In_1702);
and U737 (N_737,In_2518,In_2311);
or U738 (N_738,In_2696,In_1978);
or U739 (N_739,In_2475,In_1171);
nor U740 (N_740,In_765,In_2338);
nor U741 (N_741,In_1735,In_1268);
nand U742 (N_742,In_2717,In_2976);
nand U743 (N_743,In_2723,In_1877);
or U744 (N_744,In_1749,In_496);
or U745 (N_745,In_1784,In_1521);
and U746 (N_746,In_617,In_2757);
nor U747 (N_747,In_1004,In_503);
nand U748 (N_748,In_454,In_2014);
nor U749 (N_749,In_2219,In_1867);
nor U750 (N_750,In_847,In_39);
nand U751 (N_751,In_69,In_1753);
nand U752 (N_752,In_2771,In_1285);
nor U753 (N_753,In_2075,In_1640);
or U754 (N_754,In_2276,In_2827);
and U755 (N_755,In_2979,In_1642);
nand U756 (N_756,In_2359,In_48);
nand U757 (N_757,In_2714,In_2749);
xor U758 (N_758,In_30,In_1637);
nor U759 (N_759,In_997,In_2028);
or U760 (N_760,In_2606,In_2507);
or U761 (N_761,In_424,In_1563);
xnor U762 (N_762,In_2920,In_2228);
or U763 (N_763,In_1114,In_978);
nand U764 (N_764,In_1935,In_1230);
nand U765 (N_765,In_528,In_1721);
and U766 (N_766,In_887,In_1014);
nand U767 (N_767,In_907,In_425);
or U768 (N_768,In_2747,In_1704);
xnor U769 (N_769,In_700,In_1868);
nor U770 (N_770,In_734,In_2460);
xor U771 (N_771,In_1450,In_1652);
nand U772 (N_772,In_344,In_2119);
or U773 (N_773,In_2706,In_2326);
nor U774 (N_774,In_535,In_2815);
nand U775 (N_775,In_2417,In_66);
nor U776 (N_776,In_210,In_864);
and U777 (N_777,In_2795,In_531);
or U778 (N_778,In_910,In_543);
and U779 (N_779,In_903,In_397);
and U780 (N_780,In_1094,In_515);
and U781 (N_781,In_1963,In_2519);
nor U782 (N_782,In_61,In_1300);
xor U783 (N_783,In_26,In_2187);
nor U784 (N_784,In_1606,In_1196);
nor U785 (N_785,In_718,In_277);
xnor U786 (N_786,In_2065,In_455);
and U787 (N_787,In_1666,In_140);
nor U788 (N_788,In_1969,In_2683);
nand U789 (N_789,In_1922,In_874);
xnor U790 (N_790,In_1639,In_2060);
or U791 (N_791,In_892,In_2079);
and U792 (N_792,In_1430,In_1938);
nor U793 (N_793,In_1856,In_1850);
and U794 (N_794,In_444,In_2140);
or U795 (N_795,In_1898,In_746);
xnor U796 (N_796,In_2591,In_1038);
nor U797 (N_797,In_408,In_2501);
xor U798 (N_798,In_778,In_335);
xor U799 (N_799,In_478,In_901);
xnor U800 (N_800,In_1540,In_289);
xor U801 (N_801,In_2862,In_1067);
nor U802 (N_802,In_2804,In_1123);
nand U803 (N_803,In_578,In_713);
nor U804 (N_804,In_1574,In_1689);
or U805 (N_805,In_733,In_510);
nor U806 (N_806,In_1925,In_50);
or U807 (N_807,In_730,In_2194);
xnor U808 (N_808,In_307,In_1555);
nand U809 (N_809,In_2039,In_2297);
nor U810 (N_810,In_240,In_1401);
nor U811 (N_811,In_1846,In_1858);
nor U812 (N_812,In_276,In_826);
and U813 (N_813,In_1537,In_2097);
or U814 (N_814,In_624,In_156);
nand U815 (N_815,In_2959,In_2191);
nand U816 (N_816,In_2598,In_390);
xor U817 (N_817,In_2934,In_2857);
and U818 (N_818,In_1414,In_1105);
nand U819 (N_819,In_2320,In_2391);
and U820 (N_820,In_2664,In_2626);
or U821 (N_821,In_1544,In_1489);
nand U822 (N_822,In_1239,In_1551);
nand U823 (N_823,In_905,In_1843);
nand U824 (N_824,In_1698,In_852);
or U825 (N_825,In_76,In_2255);
or U826 (N_826,In_3,In_2377);
xnor U827 (N_827,In_2081,In_1366);
xnor U828 (N_828,In_2881,In_211);
xnor U829 (N_829,In_330,In_2821);
xnor U830 (N_830,In_537,In_1478);
or U831 (N_831,In_422,In_889);
nor U832 (N_832,In_2814,In_2459);
nor U833 (N_833,In_472,In_1244);
nor U834 (N_834,In_1445,In_2565);
nor U835 (N_835,In_2221,In_2879);
nand U836 (N_836,In_805,In_2721);
or U837 (N_837,In_1487,In_1966);
and U838 (N_838,In_2294,In_506);
nor U839 (N_839,In_2002,In_2091);
or U840 (N_840,In_2442,In_1173);
xor U841 (N_841,In_1772,In_2509);
xnor U842 (N_842,In_77,In_869);
xor U843 (N_843,In_1854,In_762);
nor U844 (N_844,In_2019,In_2816);
and U845 (N_845,In_845,In_2851);
nand U846 (N_846,In_1206,In_1879);
and U847 (N_847,In_121,In_1774);
and U848 (N_848,In_1198,In_1767);
and U849 (N_849,In_1186,In_2256);
xor U850 (N_850,In_2286,In_2169);
or U851 (N_851,In_915,In_2084);
nand U852 (N_852,In_1020,In_2327);
nor U853 (N_853,In_922,In_1007);
nand U854 (N_854,In_34,In_51);
and U855 (N_855,In_775,In_684);
xnor U856 (N_856,In_70,In_2687);
xor U857 (N_857,In_1960,In_2455);
and U858 (N_858,In_2952,In_1570);
and U859 (N_859,In_977,In_1633);
xor U860 (N_860,In_246,In_2415);
or U861 (N_861,In_2670,In_379);
or U862 (N_862,In_2887,In_403);
xor U863 (N_863,In_2582,In_2917);
nor U864 (N_864,In_1909,In_830);
nand U865 (N_865,In_1687,In_1233);
xor U866 (N_866,In_1819,In_1437);
and U867 (N_867,In_1458,In_2199);
nand U868 (N_868,In_2856,In_571);
nor U869 (N_869,In_2308,In_2125);
xnor U870 (N_870,In_1756,In_309);
and U871 (N_871,In_2186,In_819);
or U872 (N_872,In_929,In_893);
and U873 (N_873,In_2318,In_1260);
xnor U874 (N_874,In_1463,In_2050);
nor U875 (N_875,In_2383,In_56);
xor U876 (N_876,In_605,In_1498);
or U877 (N_877,In_2503,In_238);
or U878 (N_878,In_301,In_1641);
xor U879 (N_879,In_935,In_2798);
nand U880 (N_880,In_1130,In_810);
or U881 (N_881,In_1800,In_1019);
or U882 (N_882,In_798,In_1311);
and U883 (N_883,In_1157,In_1572);
xor U884 (N_884,In_1603,In_87);
xor U885 (N_885,In_2724,In_521);
or U886 (N_886,In_1732,In_1372);
nor U887 (N_887,In_389,In_2810);
nand U888 (N_888,In_1907,In_799);
nor U889 (N_889,In_1823,In_1713);
nand U890 (N_890,In_2995,In_2679);
or U891 (N_891,In_2755,In_2925);
xnor U892 (N_892,In_400,In_253);
nand U893 (N_893,In_787,In_1926);
or U894 (N_894,In_1959,In_1387);
nor U895 (N_895,In_620,In_1872);
or U896 (N_896,In_2550,In_2632);
nand U897 (N_897,In_373,In_6);
nor U898 (N_898,In_1046,In_2290);
xor U899 (N_899,In_2179,In_2073);
xnor U900 (N_900,In_2962,In_495);
nor U901 (N_901,In_1354,In_1199);
nand U902 (N_902,In_2092,In_2176);
nor U903 (N_903,In_1504,In_2237);
or U904 (N_904,In_2231,In_2514);
nand U905 (N_905,In_244,In_366);
xnor U906 (N_906,In_2448,In_596);
and U907 (N_907,In_2576,In_1495);
and U908 (N_908,In_2325,In_1348);
xor U909 (N_909,In_658,In_2044);
xnor U910 (N_910,In_1190,In_2994);
and U911 (N_911,In_1999,In_430);
xnor U912 (N_912,In_631,In_813);
xnor U913 (N_913,In_801,In_753);
or U914 (N_914,In_2274,In_288);
and U915 (N_915,In_2032,In_2803);
xor U916 (N_916,In_877,In_1741);
and U917 (N_917,In_2111,In_2986);
or U918 (N_918,In_1160,In_554);
and U919 (N_919,In_630,In_1678);
nor U920 (N_920,In_1737,In_395);
nor U921 (N_921,In_2560,In_207);
xnor U922 (N_922,In_1871,In_2634);
nor U923 (N_923,In_2581,In_1398);
nor U924 (N_924,In_29,In_2566);
or U925 (N_925,In_1225,In_1575);
nor U926 (N_926,In_720,In_1058);
nor U927 (N_927,In_385,In_465);
and U928 (N_928,In_438,In_709);
nand U929 (N_929,In_2160,In_2291);
nand U930 (N_930,In_2736,In_177);
and U931 (N_931,In_1477,In_1362);
xor U932 (N_932,In_2227,In_2638);
and U933 (N_933,In_2568,In_1290);
nand U934 (N_934,In_1367,In_1578);
and U935 (N_935,In_749,In_1109);
and U936 (N_936,In_949,In_2792);
xor U937 (N_937,In_2852,In_2289);
xnor U938 (N_938,In_2098,In_2447);
nand U939 (N_939,In_2173,In_663);
nor U940 (N_940,In_2778,In_2424);
and U941 (N_941,In_1677,In_536);
nor U942 (N_942,In_1515,In_548);
and U943 (N_943,In_511,In_544);
xnor U944 (N_944,In_1355,In_2147);
or U945 (N_945,In_2247,In_383);
or U946 (N_946,In_909,In_2068);
or U947 (N_947,In_2685,In_2378);
or U948 (N_948,In_1278,In_2613);
and U949 (N_949,In_1950,In_2943);
and U950 (N_950,In_2393,In_163);
nor U951 (N_951,In_1610,In_1501);
xor U952 (N_952,In_1410,In_2238);
xnor U953 (N_953,In_1153,In_1794);
nand U954 (N_954,In_752,In_2617);
nor U955 (N_955,In_1775,In_1761);
or U956 (N_956,In_558,In_1813);
xor U957 (N_957,In_2604,In_2180);
xor U958 (N_958,In_453,In_2737);
and U959 (N_959,In_1750,In_1802);
and U960 (N_960,In_2132,In_426);
nor U961 (N_961,In_721,In_323);
nand U962 (N_962,In_2262,In_1764);
nand U963 (N_963,In_36,In_2235);
nand U964 (N_964,In_2944,In_1193);
xor U965 (N_965,In_409,In_2193);
xnor U966 (N_966,In_2733,In_317);
nand U967 (N_967,In_616,In_1622);
and U968 (N_968,In_2873,In_807);
nand U969 (N_969,In_1531,In_1132);
and U970 (N_970,In_846,In_1303);
nor U971 (N_971,In_2413,In_2671);
and U972 (N_972,In_1806,In_955);
xnor U973 (N_973,In_2491,In_1267);
nand U974 (N_974,In_1791,In_1030);
and U975 (N_975,In_1010,In_1338);
nor U976 (N_976,In_2779,In_989);
xor U977 (N_977,In_152,In_2332);
or U978 (N_978,In_2870,In_930);
or U979 (N_979,In_2177,In_2919);
and U980 (N_980,In_1479,In_1593);
nand U981 (N_981,In_2456,In_1866);
and U982 (N_982,In_2537,In_2205);
and U983 (N_983,In_327,In_1340);
nor U984 (N_984,In_525,In_560);
xnor U985 (N_985,In_2003,In_2950);
or U986 (N_986,In_1466,In_1940);
or U987 (N_987,In_2806,In_2791);
nor U988 (N_988,In_1536,In_706);
nor U989 (N_989,In_1976,In_2512);
and U990 (N_990,In_1301,In_302);
and U991 (N_991,In_519,In_2450);
or U992 (N_992,In_2293,In_1037);
xor U993 (N_993,In_2552,In_1783);
nor U994 (N_994,In_1720,In_2762);
nor U995 (N_995,In_290,In_1288);
nand U996 (N_996,In_2768,In_1860);
and U997 (N_997,In_2781,In_773);
or U998 (N_998,In_2498,In_2);
nor U999 (N_999,In_1008,In_2430);
nand U1000 (N_1000,In_2489,In_2216);
or U1001 (N_1001,In_2564,In_2402);
and U1002 (N_1002,In_925,In_2777);
nor U1003 (N_1003,In_1655,In_2011);
and U1004 (N_1004,In_332,In_1815);
or U1005 (N_1005,In_2644,In_1360);
xnor U1006 (N_1006,In_143,In_139);
or U1007 (N_1007,In_1419,In_1462);
or U1008 (N_1008,In_2545,In_2676);
or U1009 (N_1009,In_1339,In_677);
xnor U1010 (N_1010,In_584,In_1880);
nand U1011 (N_1011,In_2184,In_1251);
and U1012 (N_1012,In_2230,In_62);
xor U1013 (N_1013,In_346,In_2765);
xnor U1014 (N_1014,In_2921,In_664);
xor U1015 (N_1015,In_1472,In_1560);
xnor U1016 (N_1016,In_494,In_1894);
nand U1017 (N_1017,In_1353,In_824);
nor U1018 (N_1018,In_1795,In_1530);
nor U1019 (N_1019,In_1914,In_28);
xnor U1020 (N_1020,In_1875,In_2114);
or U1021 (N_1021,In_175,In_574);
and U1022 (N_1022,In_648,In_1947);
xnor U1023 (N_1023,In_1597,In_938);
or U1024 (N_1024,In_2811,In_232);
nor U1025 (N_1025,In_178,In_1734);
nand U1026 (N_1026,In_2432,In_559);
xor U1027 (N_1027,In_1158,In_1785);
or U1028 (N_1028,In_1552,In_2684);
or U1029 (N_1029,In_546,In_1954);
nand U1030 (N_1030,In_1183,In_2141);
or U1031 (N_1031,In_1701,In_2394);
or U1032 (N_1032,In_1644,In_1382);
xor U1033 (N_1033,In_1324,In_1757);
and U1034 (N_1034,In_2517,In_1448);
nand U1035 (N_1035,In_2858,In_46);
or U1036 (N_1036,In_2874,In_2911);
nor U1037 (N_1037,In_2622,In_193);
nor U1038 (N_1038,In_1900,In_2872);
xor U1039 (N_1039,In_2023,In_1282);
nor U1040 (N_1040,In_255,In_312);
and U1041 (N_1041,In_2049,In_569);
nand U1042 (N_1042,In_653,In_2555);
nor U1043 (N_1043,In_423,In_2353);
nor U1044 (N_1044,In_2668,In_897);
nor U1045 (N_1045,In_2960,In_2035);
and U1046 (N_1046,In_2692,In_2875);
xor U1047 (N_1047,In_1346,In_2900);
and U1048 (N_1048,In_2553,In_1565);
xor U1049 (N_1049,In_24,In_1921);
nor U1050 (N_1050,In_2066,In_1882);
nor U1051 (N_1051,In_2807,In_1928);
xnor U1052 (N_1052,In_610,In_2037);
nand U1053 (N_1053,In_2257,In_2527);
xor U1054 (N_1054,In_523,In_2117);
or U1055 (N_1055,In_529,In_2495);
nor U1056 (N_1056,In_1664,In_2908);
nor U1057 (N_1057,In_2006,In_829);
nand U1058 (N_1058,In_970,In_1979);
xor U1059 (N_1059,In_1897,In_637);
xnor U1060 (N_1060,In_2471,In_1507);
nand U1061 (N_1061,In_1809,In_1054);
and U1062 (N_1062,In_2789,In_952);
nor U1063 (N_1063,In_1165,In_45);
nand U1064 (N_1064,In_696,In_151);
nor U1065 (N_1065,In_1752,In_924);
xnor U1066 (N_1066,In_2183,In_2439);
nor U1067 (N_1067,In_1247,In_367);
nand U1068 (N_1068,In_421,In_983);
xor U1069 (N_1069,In_1357,In_1016);
or U1070 (N_1070,In_1844,In_249);
xor U1071 (N_1071,In_147,In_1337);
or U1072 (N_1072,In_2659,In_363);
and U1073 (N_1073,In_328,In_2590);
or U1074 (N_1074,In_1231,In_2627);
and U1075 (N_1075,In_2143,In_701);
or U1076 (N_1076,In_2300,In_1977);
or U1077 (N_1077,In_2758,In_568);
and U1078 (N_1078,In_451,In_1588);
xor U1079 (N_1079,In_2543,In_320);
xor U1080 (N_1080,In_2163,In_823);
nor U1081 (N_1081,In_57,In_2126);
xnor U1082 (N_1082,In_2854,In_1538);
nor U1083 (N_1083,In_538,In_1325);
xor U1084 (N_1084,In_1989,In_1653);
and U1085 (N_1085,In_919,In_2754);
xor U1086 (N_1086,In_641,In_1700);
xnor U1087 (N_1087,In_1509,In_2593);
and U1088 (N_1088,In_1148,In_870);
nand U1089 (N_1089,In_1365,In_1352);
and U1090 (N_1090,In_2499,In_2429);
and U1091 (N_1091,In_1591,In_2831);
nor U1092 (N_1092,In_1582,In_414);
nand U1093 (N_1093,In_1120,In_2420);
and U1094 (N_1094,In_951,In_993);
nand U1095 (N_1095,In_2083,In_2161);
or U1096 (N_1096,In_104,In_1825);
nor U1097 (N_1097,In_913,In_1777);
nand U1098 (N_1098,In_844,In_580);
nand U1099 (N_1099,In_2328,In_1017);
nor U1100 (N_1100,In_982,In_2669);
xor U1101 (N_1101,In_692,In_221);
nor U1102 (N_1102,In_182,In_2693);
and U1103 (N_1103,In_2534,In_2426);
nor U1104 (N_1104,In_1798,In_2213);
nand U1105 (N_1105,In_739,In_411);
and U1106 (N_1106,In_820,In_2153);
or U1107 (N_1107,In_166,In_1513);
and U1108 (N_1108,In_751,In_2025);
and U1109 (N_1109,In_2931,In_2295);
nand U1110 (N_1110,In_2772,In_2021);
nor U1111 (N_1111,In_1080,In_880);
nand U1112 (N_1112,In_144,In_1628);
or U1113 (N_1113,In_817,In_2197);
and U1114 (N_1114,In_1691,In_2611);
xor U1115 (N_1115,In_2406,In_96);
nor U1116 (N_1116,In_1090,In_2443);
and U1117 (N_1117,In_2342,In_2661);
and U1118 (N_1118,In_2218,In_368);
xor U1119 (N_1119,In_2998,In_2283);
nand U1120 (N_1120,In_2155,In_1319);
nor U1121 (N_1121,In_551,In_581);
or U1122 (N_1122,In_392,In_2571);
nor U1123 (N_1123,In_2838,In_2266);
and U1124 (N_1124,In_2086,In_2261);
xnor U1125 (N_1125,In_2123,In_2884);
and U1126 (N_1126,In_1436,In_380);
xor U1127 (N_1127,In_1669,In_1331);
or U1128 (N_1128,In_107,In_1930);
and U1129 (N_1129,In_1018,In_2502);
nand U1130 (N_1130,In_2258,In_1068);
nand U1131 (N_1131,In_1056,In_2524);
xor U1132 (N_1132,In_242,In_2259);
nor U1133 (N_1133,In_1293,In_1309);
or U1134 (N_1134,In_158,In_1273);
and U1135 (N_1135,In_497,In_2913);
nor U1136 (N_1136,In_2559,In_2182);
or U1137 (N_1137,In_1821,In_1943);
xnor U1138 (N_1138,In_1135,In_1580);
xnor U1139 (N_1139,In_895,In_2440);
nand U1140 (N_1140,In_2547,In_2535);
and U1141 (N_1141,In_2089,In_188);
or U1142 (N_1142,In_2860,In_1957);
nor U1143 (N_1143,In_412,In_113);
nor U1144 (N_1144,In_1996,In_2896);
xor U1145 (N_1145,In_1261,In_284);
nand U1146 (N_1146,In_1768,In_1376);
nor U1147 (N_1147,In_1074,In_1127);
xor U1148 (N_1148,In_161,In_2702);
nor U1149 (N_1149,In_2802,In_123);
nor U1150 (N_1150,In_2260,In_1062);
nand U1151 (N_1151,In_223,In_1668);
nor U1152 (N_1152,In_2453,In_2379);
xnor U1153 (N_1153,In_827,In_2168);
xor U1154 (N_1154,In_1696,In_1613);
and U1155 (N_1155,In_2694,In_53);
nor U1156 (N_1156,In_2157,In_1619);
or U1157 (N_1157,In_157,In_2902);
nor U1158 (N_1158,In_1021,In_1296);
nor U1159 (N_1159,In_283,In_628);
or U1160 (N_1160,In_1321,In_490);
nor U1161 (N_1161,In_2483,In_1384);
and U1162 (N_1162,In_1424,In_183);
xnor U1163 (N_1163,In_2385,In_393);
nand U1164 (N_1164,In_1517,In_666);
nor U1165 (N_1165,In_2435,In_784);
xnor U1166 (N_1166,In_985,In_1744);
or U1167 (N_1167,In_1654,In_2351);
or U1168 (N_1168,In_2031,In_2496);
nor U1169 (N_1169,In_1832,In_1423);
or U1170 (N_1170,In_2725,In_1270);
nor U1171 (N_1171,In_2446,In_278);
and U1172 (N_1172,In_2715,In_1228);
nor U1173 (N_1173,In_1431,In_1335);
nand U1174 (N_1174,In_1334,In_1660);
nor U1175 (N_1175,In_2339,In_2346);
or U1176 (N_1176,In_1256,In_2302);
or U1177 (N_1177,In_21,In_1415);
xnor U1178 (N_1178,In_1631,In_1269);
nor U1179 (N_1179,In_1932,In_1060);
nor U1180 (N_1180,In_2826,In_2808);
nand U1181 (N_1181,In_791,In_2928);
xor U1182 (N_1182,In_229,In_2476);
xnor U1183 (N_1183,In_1217,In_360);
or U1184 (N_1184,In_2370,In_2533);
or U1185 (N_1185,In_1246,In_1320);
nor U1186 (N_1186,In_693,In_1254);
and U1187 (N_1187,In_1077,In_2009);
nor U1188 (N_1188,In_1350,In_1428);
nand U1189 (N_1189,In_2368,In_2701);
nor U1190 (N_1190,In_1394,In_195);
xor U1191 (N_1191,In_1891,In_1370);
nand U1192 (N_1192,In_1719,In_1865);
nand U1193 (N_1193,In_484,In_2859);
xor U1194 (N_1194,In_219,In_2775);
xnor U1195 (N_1195,In_2773,In_1663);
and U1196 (N_1196,In_2698,In_1505);
nor U1197 (N_1197,In_2600,In_226);
nor U1198 (N_1198,In_2030,In_1421);
xor U1199 (N_1199,In_2468,In_2639);
xor U1200 (N_1200,In_429,N_601);
or U1201 (N_1201,N_1142,In_2045);
nor U1202 (N_1202,N_261,In_1667);
nor U1203 (N_1203,In_2371,In_2087);
and U1204 (N_1204,N_708,N_802);
nor U1205 (N_1205,N_963,N_271);
or U1206 (N_1206,N_304,N_496);
xor U1207 (N_1207,N_342,N_655);
and U1208 (N_1208,N_996,N_823);
nor U1209 (N_1209,N_108,In_1905);
xor U1210 (N_1210,In_1546,N_1026);
nor U1211 (N_1211,N_954,N_349);
and U1212 (N_1212,In_1292,N_375);
and U1213 (N_1213,In_2933,N_258);
nor U1214 (N_1214,In_415,In_1403);
nand U1215 (N_1215,In_2374,N_480);
nand U1216 (N_1216,N_1015,N_252);
nand U1217 (N_1217,N_448,N_967);
or U1218 (N_1218,N_900,N_285);
and U1219 (N_1219,In_1188,N_803);
xnor U1220 (N_1220,In_1399,N_1189);
nand U1221 (N_1221,N_378,N_113);
or U1222 (N_1222,N_1129,N_296);
and U1223 (N_1223,N_428,In_2322);
nor U1224 (N_1224,N_668,N_88);
xnor U1225 (N_1225,In_1089,N_644);
nand U1226 (N_1226,N_356,In_959);
nor U1227 (N_1227,In_2397,In_2381);
and U1228 (N_1228,N_563,N_365);
nand U1229 (N_1229,N_332,N_198);
or U1230 (N_1230,In_1851,N_976);
nor U1231 (N_1231,N_830,N_945);
or U1232 (N_1232,N_689,In_394);
or U1233 (N_1233,N_1162,N_466);
nand U1234 (N_1234,N_1075,N_598);
nor U1235 (N_1235,N_1041,N_594);
nand U1236 (N_1236,N_808,N_1097);
xor U1237 (N_1237,N_94,In_2162);
nor U1238 (N_1238,N_611,In_2407);
nor U1239 (N_1239,N_54,N_91);
or U1240 (N_1240,In_2282,N_732);
xnor U1241 (N_1241,N_132,N_926);
or U1242 (N_1242,N_959,N_694);
and U1243 (N_1243,In_2631,N_532);
nor U1244 (N_1244,In_33,N_44);
xor U1245 (N_1245,N_982,N_291);
xnor U1246 (N_1246,In_1161,In_2461);
xnor U1247 (N_1247,In_1122,N_487);
or U1248 (N_1248,N_255,N_506);
xnor U1249 (N_1249,N_66,N_1133);
and U1250 (N_1250,N_597,N_266);
nand U1251 (N_1251,N_141,N_595);
nand U1252 (N_1252,N_76,In_40);
nor U1253 (N_1253,In_2621,N_574);
xnor U1254 (N_1254,N_903,N_727);
and U1255 (N_1255,In_2926,N_118);
and U1256 (N_1256,N_1106,In_2899);
nand U1257 (N_1257,In_1234,N_1040);
xor U1258 (N_1258,N_476,N_393);
nand U1259 (N_1259,In_933,N_806);
and U1260 (N_1260,N_321,N_718);
or U1261 (N_1261,N_279,N_663);
or U1262 (N_1262,N_166,In_2020);
nor U1263 (N_1263,N_862,N_741);
nor U1264 (N_1264,In_1987,N_586);
and U1265 (N_1265,N_867,N_844);
or U1266 (N_1266,N_1172,N_204);
and U1267 (N_1267,N_866,N_951);
or U1268 (N_1268,N_878,N_922);
nand U1269 (N_1269,N_1063,N_210);
and U1270 (N_1270,In_1564,In_215);
and U1271 (N_1271,N_721,N_714);
xnor U1272 (N_1272,In_2751,N_1132);
nand U1273 (N_1273,N_914,N_283);
or U1274 (N_1274,In_1215,N_659);
nand U1275 (N_1275,N_560,In_2040);
nand U1276 (N_1276,In_1516,N_746);
xor U1277 (N_1277,N_67,N_173);
or U1278 (N_1278,N_429,N_119);
xor U1279 (N_1279,N_536,N_664);
nor U1280 (N_1280,N_392,N_1039);
nand U1281 (N_1281,N_992,In_1927);
or U1282 (N_1282,N_972,N_956);
nor U1283 (N_1283,N_339,N_1094);
or U1284 (N_1284,N_837,N_931);
nand U1285 (N_1285,In_196,N_768);
nor U1286 (N_1286,N_988,N_302);
and U1287 (N_1287,In_2077,N_220);
and U1288 (N_1288,In_1849,In_556);
xor U1289 (N_1289,In_1671,N_25);
and U1290 (N_1290,N_626,In_786);
xnor U1291 (N_1291,N_277,N_70);
nand U1292 (N_1292,N_1088,N_1111);
or U1293 (N_1293,N_705,In_294);
and U1294 (N_1294,N_348,In_1816);
nand U1295 (N_1295,In_2226,In_2196);
nor U1296 (N_1296,In_262,N_697);
and U1297 (N_1297,In_2234,N_1100);
nand U1298 (N_1298,In_1381,N_812);
xnor U1299 (N_1299,N_13,N_942);
nand U1300 (N_1300,In_743,N_894);
or U1301 (N_1301,N_971,In_2330);
or U1302 (N_1302,N_32,N_915);
xor U1303 (N_1303,N_522,N_278);
and U1304 (N_1304,In_774,In_2910);
xnor U1305 (N_1305,In_914,N_21);
and U1306 (N_1306,In_1755,N_670);
nand U1307 (N_1307,N_499,N_551);
xor U1308 (N_1308,N_540,N_1048);
and U1309 (N_1309,In_386,N_1161);
or U1310 (N_1310,In_1635,N_1177);
nand U1311 (N_1311,N_740,N_904);
xnor U1312 (N_1312,N_484,N_142);
or U1313 (N_1313,N_101,N_167);
and U1314 (N_1314,In_934,N_192);
nand U1315 (N_1315,N_759,N_1045);
xor U1316 (N_1316,In_636,N_1113);
or U1317 (N_1317,N_938,N_1058);
and U1318 (N_1318,N_274,N_691);
xor U1319 (N_1319,N_43,N_706);
nand U1320 (N_1320,In_304,N_92);
or U1321 (N_1321,N_1146,In_900);
or U1322 (N_1322,In_2999,N_337);
nand U1323 (N_1323,N_1053,In_2026);
xor U1324 (N_1324,N_315,In_292);
or U1325 (N_1325,In_780,N_99);
xor U1326 (N_1326,In_1690,In_1974);
and U1327 (N_1327,N_225,N_784);
xnor U1328 (N_1328,In_68,N_950);
xnor U1329 (N_1329,N_825,N_469);
or U1330 (N_1330,N_1150,In_1870);
nor U1331 (N_1331,N_405,In_2121);
nand U1332 (N_1332,N_890,N_1044);
or U1333 (N_1333,N_856,In_1429);
xor U1334 (N_1334,In_1028,In_1497);
and U1335 (N_1335,N_109,N_1152);
nor U1336 (N_1336,N_6,N_409);
and U1337 (N_1337,N_1153,N_213);
and U1338 (N_1338,In_2780,N_568);
nand U1339 (N_1339,N_769,In_2508);
and U1340 (N_1340,In_354,N_376);
or U1341 (N_1341,N_1085,N_916);
xor U1342 (N_1342,N_490,N_589);
and U1343 (N_1343,N_614,In_1811);
nor U1344 (N_1344,In_1180,In_1919);
and U1345 (N_1345,N_243,In_1389);
or U1346 (N_1346,N_548,In_1561);
xor U1347 (N_1347,N_1144,In_593);
nand U1348 (N_1348,In_2113,N_731);
xor U1349 (N_1349,N_48,N_1092);
and U1350 (N_1350,N_749,In_2357);
nor U1351 (N_1351,In_326,In_2794);
and U1352 (N_1352,In_482,N_911);
nor U1353 (N_1353,N_654,N_641);
nand U1354 (N_1354,N_1123,N_23);
and U1355 (N_1355,In_2539,N_236);
and U1356 (N_1356,In_1624,N_600);
nor U1357 (N_1357,N_368,In_296);
or U1358 (N_1358,N_455,In_75);
nand U1359 (N_1359,N_815,N_645);
and U1360 (N_1360,In_882,N_239);
or U1361 (N_1361,N_503,N_364);
nor U1362 (N_1362,In_1280,In_697);
or U1363 (N_1363,N_767,N_86);
and U1364 (N_1364,N_196,N_1003);
xor U1365 (N_1365,N_78,N_516);
nand U1366 (N_1366,N_460,N_703);
xor U1367 (N_1367,N_1021,In_285);
xor U1368 (N_1368,N_1110,N_845);
and U1369 (N_1369,N_89,N_573);
xnor U1370 (N_1370,In_2819,N_1055);
nor U1371 (N_1371,N_115,N_224);
nor U1372 (N_1372,In_642,In_1214);
and U1373 (N_1373,N_40,N_571);
or U1374 (N_1374,N_193,N_1147);
nand U1375 (N_1375,N_561,N_923);
and U1376 (N_1376,In_129,N_84);
or U1377 (N_1377,N_781,N_403);
xor U1378 (N_1378,N_724,N_1180);
nand U1379 (N_1379,In_2937,N_486);
and U1380 (N_1380,N_145,N_102);
or U1381 (N_1381,N_413,N_177);
xor U1382 (N_1382,In_1725,N_125);
nor U1383 (N_1383,In_2052,N_1156);
nand U1384 (N_1384,In_2487,In_101);
xnor U1385 (N_1385,In_1931,N_763);
nand U1386 (N_1386,In_754,N_1007);
and U1387 (N_1387,N_129,N_1182);
xnor U1388 (N_1388,In_1895,N_912);
nor U1389 (N_1389,N_228,In_16);
nand U1390 (N_1390,N_382,N_1072);
and U1391 (N_1391,N_287,In_2841);
nor U1392 (N_1392,N_515,N_424);
nor U1393 (N_1393,N_804,N_819);
nand U1394 (N_1394,In_2939,N_123);
xor U1395 (N_1395,N_700,N_504);
xnor U1396 (N_1396,N_465,In_764);
xor U1397 (N_1397,In_1519,In_1373);
xnor U1398 (N_1398,In_912,In_868);
nand U1399 (N_1399,N_523,N_776);
xor U1400 (N_1400,In_2015,N_260);
nand U1401 (N_1401,In_32,N_970);
xor U1402 (N_1402,In_420,N_895);
nor U1403 (N_1403,In_2382,N_305);
nor U1404 (N_1404,N_338,In_1608);
xnor U1405 (N_1405,N_229,In_2601);
xor U1406 (N_1406,N_68,N_1064);
or U1407 (N_1407,N_391,N_248);
xnor U1408 (N_1408,In_99,N_1199);
or U1409 (N_1409,In_1659,N_734);
and U1410 (N_1410,In_382,In_2172);
nor U1411 (N_1411,N_546,In_109);
or U1412 (N_1412,N_1087,N_1);
or U1413 (N_1413,N_816,N_352);
and U1414 (N_1414,N_233,In_2022);
nand U1415 (N_1415,In_2109,N_832);
nand U1416 (N_1416,N_169,N_328);
nor U1417 (N_1417,In_732,In_2799);
xor U1418 (N_1418,In_2741,N_957);
nor U1419 (N_1419,N_407,In_1177);
nor U1420 (N_1420,N_59,In_2128);
xnor U1421 (N_1421,N_1009,N_787);
nand U1422 (N_1422,N_467,In_1194);
xnor U1423 (N_1423,In_1592,N_160);
and U1424 (N_1424,In_1647,N_187);
or U1425 (N_1425,N_161,N_872);
nand U1426 (N_1426,N_853,N_650);
xnor U1427 (N_1427,N_122,N_358);
xor U1428 (N_1428,N_331,N_1096);
nand U1429 (N_1429,N_793,N_1069);
or U1430 (N_1430,N_754,N_998);
xor U1431 (N_1431,N_688,In_498);
nand U1432 (N_1432,In_2594,N_157);
nor U1433 (N_1433,In_2287,N_690);
nor U1434 (N_1434,In_252,In_1708);
and U1435 (N_1435,In_857,N_1174);
or U1436 (N_1436,N_1136,In_1949);
nand U1437 (N_1437,N_720,N_521);
xor U1438 (N_1438,N_936,In_1827);
xor U1439 (N_1439,N_286,N_453);
xnor U1440 (N_1440,N_692,In_1673);
nand U1441 (N_1441,N_120,N_292);
or U1442 (N_1442,In_308,N_75);
nor U1443 (N_1443,N_149,N_625);
or U1444 (N_1444,N_765,N_103);
xnor U1445 (N_1445,In_534,In_1166);
nor U1446 (N_1446,N_223,N_1022);
nor U1447 (N_1447,N_143,N_235);
nand U1448 (N_1448,N_762,N_404);
xnor U1449 (N_1449,In_401,N_334);
nand U1450 (N_1450,N_438,In_1297);
or U1451 (N_1451,N_442,In_172);
or U1452 (N_1452,In_604,N_535);
nor U1453 (N_1453,In_2707,N_1194);
and U1454 (N_1454,In_2324,In_1818);
nand U1455 (N_1455,In_2869,N_891);
or U1456 (N_1456,N_301,In_324);
nor U1457 (N_1457,In_722,In_1675);
nand U1458 (N_1458,N_478,N_319);
or U1459 (N_1459,N_18,N_146);
nand U1460 (N_1460,N_518,N_511);
nand U1461 (N_1461,In_1174,In_1213);
nand U1462 (N_1462,N_138,N_74);
xnor U1463 (N_1463,In_1604,In_1674);
nand U1464 (N_1464,N_753,N_609);
nand U1465 (N_1465,In_131,N_1043);
and U1466 (N_1466,In_118,N_502);
xnor U1467 (N_1467,In_2823,In_2599);
or U1468 (N_1468,In_916,N_1057);
and U1469 (N_1469,N_978,N_631);
nand U1470 (N_1470,N_683,N_362);
and U1471 (N_1471,N_905,N_698);
nand U1472 (N_1472,N_744,N_1066);
nand U1473 (N_1473,In_192,In_336);
nand U1474 (N_1474,In_768,N_1127);
and U1475 (N_1475,N_932,In_777);
xor U1476 (N_1476,N_826,In_1941);
xor U1477 (N_1477,In_1263,N_307);
or U1478 (N_1478,In_297,N_885);
nor U1479 (N_1479,In_206,In_1051);
and U1480 (N_1480,N_158,N_513);
nor U1481 (N_1481,N_795,In_1036);
or U1482 (N_1482,N_1124,N_716);
and U1483 (N_1483,In_2154,N_851);
nor U1484 (N_1484,N_1134,N_1001);
nor U1485 (N_1485,In_2554,In_861);
nor U1486 (N_1486,N_41,N_298);
nand U1487 (N_1487,N_807,In_404);
and U1488 (N_1488,N_237,In_2651);
or U1489 (N_1489,In_1005,N_71);
or U1490 (N_1490,In_2105,In_2029);
and U1491 (N_1491,N_294,In_1064);
xnor U1492 (N_1492,N_814,In_149);
xnor U1493 (N_1493,N_354,N_172);
xnor U1494 (N_1494,N_1109,In_2855);
and U1495 (N_1495,In_1446,N_1033);
nand U1496 (N_1496,In_2115,N_10);
or U1497 (N_1497,N_1115,In_133);
xor U1498 (N_1498,N_410,N_367);
nor U1499 (N_1499,N_877,N_1037);
nor U1500 (N_1500,In_2013,N_873);
nand U1501 (N_1501,In_2863,N_686);
or U1502 (N_1502,N_707,In_1599);
nor U1503 (N_1503,In_2356,In_85);
nand U1504 (N_1504,In_2968,N_676);
nor U1505 (N_1505,N_330,N_780);
or U1506 (N_1506,N_919,N_933);
or U1507 (N_1507,In_614,In_1432);
or U1508 (N_1508,N_1184,In_689);
nand U1509 (N_1509,In_1474,N_952);
xnor U1510 (N_1510,N_1195,In_2922);
or U1511 (N_1511,N_450,N_127);
or U1512 (N_1512,N_587,In_2575);
nor U1513 (N_1513,In_504,N_702);
or U1514 (N_1514,In_2894,N_30);
or U1515 (N_1515,In_2942,N_1070);
nor U1516 (N_1516,N_1159,N_105);
nand U1517 (N_1517,N_462,N_777);
and U1518 (N_1518,N_925,N_542);
nand U1519 (N_1519,In_2348,N_770);
xnor U1520 (N_1520,N_1187,In_224);
nand U1521 (N_1521,In_2893,N_419);
xor U1522 (N_1522,In_1607,N_289);
and U1523 (N_1523,N_195,N_530);
nor U1524 (N_1524,N_681,N_1131);
or U1525 (N_1525,N_893,In_1052);
nor U1526 (N_1526,N_987,N_33);
and U1527 (N_1527,In_1286,N_250);
xor U1528 (N_1528,In_291,N_1028);
nand U1529 (N_1529,N_756,N_558);
xnor U1530 (N_1530,In_155,In_2936);
and U1531 (N_1531,N_1196,In_1961);
nand U1532 (N_1532,N_345,N_569);
nor U1533 (N_1533,N_1186,N_1036);
or U1534 (N_1534,N_276,In_1583);
and U1535 (N_1535,N_1117,In_102);
and U1536 (N_1536,N_669,N_1032);
xnor U1537 (N_1537,In_1801,N_1082);
nor U1538 (N_1538,N_247,N_847);
or U1539 (N_1539,N_472,N_1171);
nor U1540 (N_1540,N_677,N_603);
or U1541 (N_1541,N_473,N_79);
or U1542 (N_1542,In_1310,In_97);
nand U1543 (N_1543,N_361,In_563);
or U1544 (N_1544,N_316,In_811);
nand U1545 (N_1545,N_990,N_788);
xnor U1546 (N_1546,N_343,N_549);
and U1547 (N_1547,In_939,In_2541);
xor U1548 (N_1548,N_355,N_11);
and U1549 (N_1549,In_281,In_838);
nand U1550 (N_1550,In_565,In_2720);
nor U1551 (N_1551,N_435,N_107);
nand U1552 (N_1552,N_805,N_621);
nor U1553 (N_1553,N_1017,In_1126);
xor U1554 (N_1554,N_840,N_1122);
xnor U1555 (N_1555,N_449,N_656);
nor U1556 (N_1556,In_1636,In_769);
or U1557 (N_1557,In_883,N_811);
nor U1558 (N_1558,N_865,N_612);
or U1559 (N_1559,N_318,N_1119);
or U1560 (N_1560,N_216,In_1291);
nand U1561 (N_1561,In_1411,N_1025);
nor U1562 (N_1562,N_322,N_596);
nor U1563 (N_1563,In_2222,N_444);
nor U1564 (N_1564,N_131,N_209);
nand U1565 (N_1565,N_607,N_350);
nor U1566 (N_1566,N_1103,N_46);
or U1567 (N_1567,N_1010,N_181);
xor U1568 (N_1568,N_100,N_1062);
and U1569 (N_1569,In_134,N_194);
or U1570 (N_1570,In_1227,N_185);
nor U1571 (N_1571,N_272,In_2323);
or U1572 (N_1572,N_57,In_1896);
and U1573 (N_1573,In_2528,N_81);
or U1574 (N_1574,N_344,In_2641);
or U1575 (N_1575,N_909,N_333);
xor U1576 (N_1576,N_1198,In_992);
and U1577 (N_1577,In_357,N_927);
nand U1578 (N_1578,In_2945,In_2423);
xor U1579 (N_1579,N_836,N_1011);
nand U1580 (N_1580,N_159,N_52);
xor U1581 (N_1581,N_72,In_1369);
or U1582 (N_1582,N_458,N_876);
nand U1583 (N_1583,N_726,N_649);
nand U1584 (N_1584,N_743,N_680);
or U1585 (N_1585,N_577,N_796);
xnor U1586 (N_1586,N_280,N_387);
nor U1587 (N_1587,N_208,In_1164);
nand U1588 (N_1588,N_979,N_779);
nand U1589 (N_1589,N_699,N_98);
or U1590 (N_1590,N_491,N_180);
and U1591 (N_1591,In_1804,In_1022);
or U1592 (N_1592,N_0,N_605);
or U1593 (N_1593,N_259,N_742);
or U1594 (N_1594,N_841,N_679);
or U1595 (N_1595,N_565,N_556);
xnor U1596 (N_1596,N_165,N_53);
xor U1597 (N_1597,N_827,In_2048);
nand U1598 (N_1598,N_417,N_541);
and U1599 (N_1599,N_562,In_418);
nor U1600 (N_1600,N_730,N_557);
xor U1601 (N_1601,In_945,N_1141);
nor U1602 (N_1602,In_1470,In_1550);
or U1603 (N_1603,N_953,In_2267);
nand U1604 (N_1604,N_634,N_1151);
nor U1605 (N_1605,N_1027,N_1126);
nor U1606 (N_1606,N_884,N_902);
nor U1607 (N_1607,N_218,N_682);
nor U1608 (N_1608,N_69,N_1107);
and U1609 (N_1609,N_673,N_31);
xnor U1610 (N_1610,In_1948,N_965);
and U1611 (N_1611,N_1114,In_2878);
nand U1612 (N_1612,N_396,In_655);
and U1613 (N_1613,N_590,N_1005);
nand U1614 (N_1614,N_222,In_2652);
and U1615 (N_1615,In_1343,N_369);
or U1616 (N_1616,In_2041,N_539);
or U1617 (N_1617,N_162,In_387);
and U1618 (N_1618,N_859,N_928);
nor U1619 (N_1619,N_997,N_789);
nand U1620 (N_1620,In_124,N_667);
nand U1621 (N_1621,N_717,N_745);
nand U1622 (N_1622,In_2281,In_127);
nor U1623 (N_1623,N_1067,N_402);
nand U1624 (N_1624,N_809,In_298);
xor U1625 (N_1625,N_580,N_564);
xor U1626 (N_1626,In_2603,N_163);
or U1627 (N_1627,N_95,N_879);
or U1628 (N_1628,N_50,In_2877);
or U1629 (N_1629,N_311,N_1038);
nand U1630 (N_1630,In_875,In_615);
xnor U1631 (N_1631,N_188,N_1188);
nand U1632 (N_1632,N_439,In_660);
nand U1633 (N_1633,N_899,N_251);
xor U1634 (N_1634,N_647,In_1904);
nor U1635 (N_1635,N_418,In_2106);
or U1636 (N_1636,In_205,N_269);
xnor U1637 (N_1637,N_456,N_863);
and U1638 (N_1638,In_2965,N_616);
nor U1639 (N_1639,N_12,N_148);
nand U1640 (N_1640,N_980,N_186);
nand U1641 (N_1641,N_665,In_2366);
xnor U1642 (N_1642,N_1020,In_1587);
nor U1643 (N_1643,In_843,In_2796);
nand U1644 (N_1644,N_973,In_2239);
nor U1645 (N_1645,In_1751,In_2532);
nand U1646 (N_1646,N_985,In_2786);
and U1647 (N_1647,In_2414,N_1019);
and U1648 (N_1648,N_327,In_782);
xnor U1649 (N_1649,N_1197,In_527);
nand U1650 (N_1650,N_999,N_1160);
nand U1651 (N_1651,N_299,N_918);
or U1652 (N_1652,In_1299,In_979);
xor U1653 (N_1653,In_311,N_817);
nor U1654 (N_1654,In_601,N_593);
and U1655 (N_1655,In_576,In_2993);
nor U1656 (N_1656,N_351,In_1029);
and U1657 (N_1657,In_626,In_2843);
xor U1658 (N_1658,N_520,In_2885);
nor U1659 (N_1659,N_268,In_316);
nand U1660 (N_1660,In_2876,N_871);
nand U1661 (N_1661,N_913,N_63);
nor U1662 (N_1662,In_1730,In_1145);
nor U1663 (N_1663,N_329,N_554);
or U1664 (N_1664,In_800,In_405);
nor U1665 (N_1665,N_678,N_388);
and U1666 (N_1666,In_287,N_529);
nor U1667 (N_1667,In_1224,N_930);
or U1668 (N_1668,N_1135,N_635);
nand U1669 (N_1669,N_1149,In_2703);
nand U1670 (N_1670,In_1041,N_1181);
nor U1671 (N_1671,N_408,In_1395);
nand U1672 (N_1672,N_643,N_1047);
nor U1673 (N_1673,In_1447,N_723);
nand U1674 (N_1674,In_1656,In_2074);
nor U1675 (N_1675,N_666,N_87);
xor U1676 (N_1676,N_443,In_1097);
nor U1677 (N_1677,N_1143,N_1068);
xnor U1678 (N_1678,N_591,N_295);
nand U1679 (N_1679,N_636,N_934);
or U1680 (N_1680,In_1838,N_948);
xor U1681 (N_1681,N_534,N_585);
nand U1682 (N_1682,N_842,N_93);
nor U1683 (N_1683,N_994,In_1672);
or U1684 (N_1684,N_618,N_901);
nor U1685 (N_1685,In_2612,In_1204);
and U1686 (N_1686,In_681,N_82);
nand U1687 (N_1687,N_323,N_713);
nor U1688 (N_1688,In_1728,N_949);
or U1689 (N_1689,N_671,In_2891);
or U1690 (N_1690,N_308,N_652);
nor U1691 (N_1691,N_341,N_615);
xor U1692 (N_1692,N_1091,In_2444);
xor U1693 (N_1693,N_488,N_481);
nand U1694 (N_1694,N_398,N_1175);
or U1695 (N_1695,N_599,N_920);
or U1696 (N_1696,N_60,N_137);
xor U1697 (N_1697,In_1695,N_974);
xor U1698 (N_1698,N_45,In_1082);
nand U1699 (N_1699,N_582,N_182);
or U1700 (N_1700,N_134,N_16);
nor U1701 (N_1701,In_2284,In_759);
nand U1702 (N_1702,In_618,N_1190);
and U1703 (N_1703,N_313,In_1272);
nor U1704 (N_1704,In_2038,N_130);
and U1705 (N_1705,In_1892,In_2629);
nand U1706 (N_1706,N_738,N_380);
or U1707 (N_1707,In_1034,In_1724);
xnor U1708 (N_1708,N_1155,N_501);
and U1709 (N_1709,In_2201,N_785);
xor U1710 (N_1710,N_267,N_207);
or U1711 (N_1711,N_1000,N_1077);
nand U1712 (N_1712,N_1098,N_1052);
xnor U1713 (N_1713,In_2674,In_169);
and U1714 (N_1714,N_461,In_1972);
nand U1715 (N_1715,N_1089,N_1059);
nor U1716 (N_1716,In_64,N_366);
or U1717 (N_1717,In_92,In_2602);
and U1718 (N_1718,In_2766,N_711);
or U1719 (N_1719,In_2288,N_800);
and U1720 (N_1720,In_2010,N_238);
and U1721 (N_1721,N_90,N_28);
xnor U1722 (N_1722,N_854,In_831);
or U1723 (N_1723,N_112,N_77);
or U1724 (N_1724,N_219,In_1336);
nand U1725 (N_1725,N_73,In_339);
nand U1726 (N_1726,N_494,N_29);
nand U1727 (N_1727,N_509,N_293);
and U1728 (N_1728,In_2171,N_921);
nor U1729 (N_1729,N_24,In_1240);
nand U1730 (N_1730,N_608,N_320);
nor U1731 (N_1731,In_943,N_775);
or U1732 (N_1732,N_1054,N_514);
nor U1733 (N_1733,In_1441,N_1154);
xnor U1734 (N_1734,N_191,N_774);
xnor U1735 (N_1735,In_1848,N_140);
xnor U1736 (N_1736,N_61,N_685);
nand U1737 (N_1737,N_898,N_1080);
xor U1738 (N_1738,N_373,N_833);
and U1739 (N_1739,In_1361,N_1118);
or U1740 (N_1740,In_1024,In_2970);
xor U1741 (N_1741,N_906,N_211);
or U1742 (N_1742,In_2990,N_80);
xor U1743 (N_1743,N_39,N_524);
nor U1744 (N_1744,N_1163,In_839);
xnor U1745 (N_1745,N_736,N_755);
nand U1746 (N_1746,N_772,In_1115);
nand U1747 (N_1747,N_543,In_837);
xnor U1748 (N_1748,N_324,In_2001);
xor U1749 (N_1749,In_783,N_846);
nand U1750 (N_1750,N_588,In_731);
or U1751 (N_1751,In_203,N_426);
or U1752 (N_1752,N_661,In_2954);
and U1753 (N_1753,N_124,N_111);
xor U1754 (N_1754,N_306,In_103);
nor U1755 (N_1755,In_1716,In_2410);
or U1756 (N_1756,N_526,In_1076);
xnor U1757 (N_1757,N_270,N_672);
xor U1758 (N_1758,In_1347,N_189);
and U1759 (N_1759,In_473,N_1112);
nor U1760 (N_1760,In_343,N_171);
xor U1761 (N_1761,N_416,In_2333);
nor U1762 (N_1762,In_1553,In_2580);
nor U1763 (N_1763,N_870,In_1295);
nor U1764 (N_1764,N_386,N_629);
nand U1765 (N_1765,N_857,In_2834);
xor U1766 (N_1766,N_1099,N_693);
or U1767 (N_1767,In_2665,In_2480);
and U1768 (N_1768,N_85,N_1138);
nor U1769 (N_1769,N_1139,N_758);
xnor U1770 (N_1770,In_1964,N_962);
nand U1771 (N_1771,N_452,N_750);
and U1772 (N_1772,N_135,In_2912);
xor U1773 (N_1773,N_431,In_2700);
or U1774 (N_1774,N_454,N_964);
or U1775 (N_1775,In_908,N_190);
or U1776 (N_1776,N_773,N_874);
or U1777 (N_1777,N_273,N_947);
nor U1778 (N_1778,N_710,N_147);
nand U1779 (N_1779,N_1191,In_1203);
nand U1780 (N_1780,In_1417,N_715);
nor U1781 (N_1781,N_425,N_550);
or U1782 (N_1782,N_966,N_483);
or U1783 (N_1783,N_657,N_935);
nor U1784 (N_1784,In_2007,N_421);
nand U1785 (N_1785,N_310,In_674);
and U1786 (N_1786,In_348,N_436);
nor U1787 (N_1787,In_1625,In_1621);
nand U1788 (N_1788,In_114,N_821);
nor U1789 (N_1789,In_0,N_786);
nor U1790 (N_1790,In_976,In_2941);
nor U1791 (N_1791,In_678,In_1962);
nor U1792 (N_1792,N_1178,In_315);
xor U1793 (N_1793,N_627,N_168);
and U1794 (N_1794,N_65,N_411);
or U1795 (N_1795,In_1388,In_679);
or U1796 (N_1796,In_2008,N_810);
xnor U1797 (N_1797,N_838,N_116);
nand U1798 (N_1798,N_1176,N_783);
nor U1799 (N_1799,In_1620,N_960);
xnor U1800 (N_1800,N_559,N_719);
nand U1801 (N_1801,In_65,In_740);
and U1802 (N_1802,In_1581,N_440);
xnor U1803 (N_1803,N_969,N_637);
nor U1804 (N_1804,N_981,N_164);
or U1805 (N_1805,N_1166,N_687);
nand U1806 (N_1806,N_771,N_62);
nand U1807 (N_1807,In_1789,N_638);
nor U1808 (N_1808,In_250,In_2759);
or U1809 (N_1809,N_1084,N_1013);
xor U1810 (N_1810,N_433,N_475);
nor U1811 (N_1811,N_430,In_562);
nand U1812 (N_1812,In_1121,N_538);
xnor U1813 (N_1813,N_374,N_946);
nor U1814 (N_1814,In_280,N_485);
and U1815 (N_1815,N_1008,N_4);
or U1816 (N_1816,N_56,In_1594);
xnor U1817 (N_1817,In_2042,N_422);
xnor U1818 (N_1818,N_1173,N_801);
and U1819 (N_1819,N_244,N_175);
nor U1820 (N_1820,N_648,N_883);
or U1821 (N_1821,N_1030,N_451);
xnor U1822 (N_1822,In_1995,In_100);
nand U1823 (N_1823,N_385,N_861);
xnor U1824 (N_1824,In_1069,In_2347);
nor U1825 (N_1825,N_1121,In_2175);
or U1826 (N_1826,N_1074,N_868);
xor U1827 (N_1827,In_766,In_1693);
nor U1828 (N_1828,In_1061,In_1377);
nand U1829 (N_1829,N_531,In_1152);
or U1830 (N_1830,In_588,In_1281);
nand U1831 (N_1831,In_2156,N_977);
or U1832 (N_1832,N_246,In_1874);
nor U1833 (N_1833,In_1207,N_1016);
and U1834 (N_1834,N_544,N_1128);
xor U1835 (N_1835,In_2404,In_2144);
xor U1836 (N_1836,N_1024,In_1658);
and U1837 (N_1837,In_2529,In_1810);
and U1838 (N_1838,In_2321,In_488);
nor U1839 (N_1839,N_1102,N_1073);
nor U1840 (N_1840,In_2195,In_2793);
or U1841 (N_1841,In_695,N_414);
or U1842 (N_1842,N_882,N_642);
nor U1843 (N_1843,N_212,N_199);
and U1844 (N_1844,N_1034,N_622);
nand U1845 (N_1845,N_371,N_1029);
or U1846 (N_1846,In_1912,N_17);
and U1847 (N_1847,N_1006,N_372);
nor U1848 (N_1848,N_1158,N_14);
xor U1849 (N_1849,N_848,In_1475);
or U1850 (N_1850,In_10,N_42);
xor U1851 (N_1851,In_2278,N_843);
or U1852 (N_1852,In_2137,N_824);
xnor U1853 (N_1853,N_479,In_1095);
nor U1854 (N_1854,In_557,N_1071);
nand U1855 (N_1855,In_1643,In_555);
nand U1856 (N_1856,N_508,In_2298);
nor U1857 (N_1857,N_1104,N_944);
xnor U1858 (N_1858,N_1049,N_1165);
xor U1859 (N_1859,In_2784,N_153);
nand U1860 (N_1860,In_1312,N_477);
and U1861 (N_1861,N_489,In_690);
or U1862 (N_1862,In_586,N_798);
or U1863 (N_1863,In_927,N_401);
or U1864 (N_1864,N_1179,In_1792);
and U1865 (N_1865,In_962,N_646);
and U1866 (N_1866,N_505,N_357);
or U1867 (N_1867,N_1169,N_892);
or U1868 (N_1868,N_864,N_1035);
and U1869 (N_1869,N_835,In_2915);
and U1870 (N_1870,In_2505,N_989);
nor U1871 (N_1871,In_106,N_151);
and U1872 (N_1872,N_126,In_1820);
and U1873 (N_1873,N_937,N_150);
xor U1874 (N_1874,In_1712,N_201);
or U1875 (N_1875,N_1023,In_2080);
xor U1876 (N_1876,N_1101,N_104);
or U1877 (N_1877,N_230,N_1046);
or U1878 (N_1878,In_606,N_1014);
xnor U1879 (N_1879,N_1065,In_1715);
nor U1880 (N_1880,N_200,N_752);
nor U1881 (N_1881,In_2710,N_47);
or U1882 (N_1882,In_2927,N_896);
and U1883 (N_1883,In_1023,N_986);
nor U1884 (N_1884,In_1859,N_828);
and U1885 (N_1885,N_993,N_660);
nand U1886 (N_1886,In_191,In_1650);
and U1887 (N_1887,In_1402,In_2647);
xnor U1888 (N_1888,In_1385,N_2);
nand U1889 (N_1889,N_1060,In_427);
or U1890 (N_1890,N_49,In_522);
or U1891 (N_1891,N_570,N_897);
and U1892 (N_1892,N_154,In_2341);
or U1893 (N_1893,In_1142,In_2061);
xor U1894 (N_1894,N_675,N_575);
or U1895 (N_1895,N_203,N_839);
or U1896 (N_1896,In_687,In_2343);
xnor U1897 (N_1897,N_1108,N_249);
or U1898 (N_1898,N_383,In_299);
and U1899 (N_1899,N_1076,In_1609);
nor U1900 (N_1900,N_347,N_395);
or U1901 (N_1901,In_19,N_377);
xnor U1902 (N_1902,N_790,N_696);
nor U1903 (N_1903,N_370,In_2129);
and U1904 (N_1904,N_470,N_492);
and U1905 (N_1905,In_1743,In_1484);
nand U1906 (N_1906,N_360,N_512);
nand U1907 (N_1907,N_566,N_1031);
xnor U1908 (N_1908,N_792,N_1079);
nand U1909 (N_1909,In_445,In_358);
or U1910 (N_1910,N_170,N_446);
nand U1911 (N_1911,N_178,N_254);
nor U1912 (N_1912,N_1170,In_2557);
xor U1913 (N_1913,N_924,In_2510);
nand U1914 (N_1914,N_434,N_764);
xnor U1915 (N_1915,N_1002,In_1202);
nand U1916 (N_1916,N_1167,N_83);
or U1917 (N_1917,In_2842,N_117);
xor U1918 (N_1918,N_240,N_447);
and U1919 (N_1919,N_139,N_1004);
xnor U1920 (N_1920,N_20,N_35);
or U1921 (N_1921,N_415,N_468);
nand U1922 (N_1922,N_257,In_2840);
and U1923 (N_1923,N_1168,In_1137);
nor U1924 (N_1924,In_2250,N_427);
xnor U1925 (N_1925,In_2069,In_2829);
and U1926 (N_1926,N_653,N_975);
xor U1927 (N_1927,N_445,N_381);
and U1928 (N_1928,N_340,N_281);
nor U1929 (N_1929,N_552,N_983);
nor U1930 (N_1930,N_1081,N_757);
and U1931 (N_1931,In_471,N_1116);
or U1932 (N_1932,N_474,N_1095);
or U1933 (N_1933,N_704,N_399);
and U1934 (N_1934,In_80,In_1857);
nor U1935 (N_1935,N_888,N_241);
xnor U1936 (N_1936,N_7,N_495);
and U1937 (N_1937,In_2101,N_533);
and U1938 (N_1938,In_2726,In_1506);
nand U1939 (N_1939,In_804,N_613);
xnor U1940 (N_1940,N_760,N_527);
or U1941 (N_1941,In_2136,In_2270);
nand U1942 (N_1942,N_858,In_88);
or U1943 (N_1943,In_1425,In_1906);
and U1944 (N_1944,N_303,N_640);
xor U1945 (N_1945,In_1461,In_228);
and U1946 (N_1946,N_1012,N_1090);
xor U1947 (N_1947,N_1148,In_2192);
and U1948 (N_1948,N_581,N_253);
nand U1949 (N_1949,In_1945,N_1185);
nand U1950 (N_1950,N_1018,N_359);
xnor U1951 (N_1951,In_375,In_31);
xor U1952 (N_1952,N_630,N_739);
nand U1953 (N_1953,N_733,In_1808);
xor U1954 (N_1954,In_2441,In_744);
and U1955 (N_1955,N_38,In_1533);
or U1956 (N_1956,N_179,N_961);
nor U1957 (N_1957,N_231,N_275);
nand U1958 (N_1958,In_2384,N_214);
nor U1959 (N_1959,N_849,N_282);
xor U1960 (N_1960,N_869,N_497);
nand U1961 (N_1961,N_227,In_95);
nand U1962 (N_1962,N_567,N_619);
xnor U1963 (N_1963,N_309,N_51);
or U1964 (N_1964,N_463,In_173);
nor U1965 (N_1965,In_2991,N_813);
nand U1966 (N_1966,N_1125,N_968);
nor U1967 (N_1967,In_1903,In_1924);
and U1968 (N_1968,N_394,In_310);
xor U1969 (N_1969,N_400,N_639);
nor U1970 (N_1970,In_1899,N_234);
xnor U1971 (N_1971,In_2753,N_886);
nand U1972 (N_1972,N_152,N_36);
or U1973 (N_1973,In_325,In_2763);
nand U1974 (N_1974,In_1313,N_1157);
nor U1975 (N_1975,N_729,In_1356);
nor U1976 (N_1976,N_799,N_1078);
or U1977 (N_1977,N_197,N_174);
nor U1978 (N_1978,N_984,In_665);
or U1979 (N_1979,In_2465,N_507);
or U1980 (N_1980,N_929,In_1405);
nand U1981 (N_1981,In_2605,N_317);
nor U1982 (N_1982,N_1145,N_326);
nor U1983 (N_1983,In_1086,N_632);
or U1984 (N_1984,N_471,In_2303);
nand U1985 (N_1985,In_2800,N_584);
or U1986 (N_1986,N_226,N_794);
nand U1987 (N_1987,N_658,N_406);
nor U1988 (N_1988,In_1245,In_2380);
nand U1989 (N_1989,N_881,N_880);
and U1990 (N_1990,N_288,N_156);
nand U1991 (N_1991,N_97,N_778);
nand U1992 (N_1992,In_2981,N_725);
nand U1993 (N_1993,N_34,N_875);
xor U1994 (N_1994,In_953,N_917);
nand U1995 (N_1995,N_547,N_761);
xor U1996 (N_1996,N_262,In_757);
xor U1997 (N_1997,N_290,N_457);
and U1998 (N_1998,In_589,N_420);
nand U1999 (N_1999,In_1146,N_15);
xnor U2000 (N_2000,N_384,N_37);
nor U2001 (N_2001,N_610,N_397);
and U2002 (N_2002,N_133,N_579);
nand U2003 (N_2003,N_300,N_202);
nand U2004 (N_2004,N_1056,N_389);
xor U2005 (N_2005,N_860,N_106);
xnor U2006 (N_2006,N_379,In_1138);
nand U2007 (N_2007,N_8,N_583);
or U2008 (N_2008,N_604,In_1433);
or U2009 (N_2009,N_624,N_184);
or U2010 (N_2010,N_850,N_709);
xnor U2011 (N_2011,N_592,In_685);
nand U2012 (N_2012,N_500,N_991);
nor U2013 (N_2013,In_1471,N_820);
nand U2014 (N_2014,N_1050,N_55);
nand U2015 (N_2015,N_958,N_390);
nor U2016 (N_2016,N_232,N_96);
nor U2017 (N_2017,N_205,In_724);
nand U2018 (N_2018,N_441,In_2688);
xnor U2019 (N_2019,In_1864,N_695);
or U2020 (N_2020,N_284,N_623);
nor U2021 (N_2021,In_1438,N_3);
or U2022 (N_2022,N_459,N_834);
and U2023 (N_2023,In_890,N_176);
nand U2024 (N_2024,N_432,N_19);
nand U2025 (N_2025,In_1911,N_245);
and U2026 (N_2026,N_701,N_628);
and U2027 (N_2027,N_22,N_737);
and U2028 (N_2028,N_263,N_1083);
and U2029 (N_2029,N_537,N_1061);
xor U2030 (N_2030,In_1223,N_748);
or U2031 (N_2031,N_855,N_155);
xnor U2032 (N_2032,N_940,N_183);
xnor U2033 (N_2033,N_545,In_1559);
xor U2034 (N_2034,N_423,N_831);
nand U2035 (N_2035,N_617,N_336);
or U2036 (N_2036,N_662,N_941);
nand U2037 (N_2037,N_528,N_1093);
xor U2038 (N_2038,N_674,N_576);
xnor U2039 (N_2039,In_1102,N_206);
and U2040 (N_2040,In_2825,In_2691);
nor U2041 (N_2041,N_221,In_849);
nor U2042 (N_2042,N_939,In_2914);
or U2043 (N_2043,N_265,N_633);
and U2044 (N_2044,N_1137,N_572);
and U2045 (N_2045,N_955,N_215);
or U2046 (N_2046,N_555,N_482);
or U2047 (N_2047,In_960,In_1333);
xnor U2048 (N_2048,N_908,N_910);
and U2049 (N_2049,N_314,N_1183);
xnor U2050 (N_2050,In_1242,N_110);
nand U2051 (N_2051,N_722,In_353);
nand U2052 (N_2052,N_1193,N_312);
xor U2053 (N_2053,N_852,N_517);
nor U2054 (N_2054,N_887,N_335);
and U2055 (N_2055,N_58,In_2051);
or U2056 (N_2056,N_510,In_958);
or U2057 (N_2057,In_1488,In_1212);
xor U2058 (N_2058,N_822,N_242);
nor U2059 (N_2059,N_735,N_498);
xor U2060 (N_2060,N_602,In_479);
and U2061 (N_2061,N_1042,In_1480);
and U2062 (N_2062,N_1130,In_2989);
xnor U2063 (N_2063,N_782,In_2313);
and U2064 (N_2064,N_907,N_728);
or U2065 (N_2065,In_452,N_1140);
nor U2066 (N_2066,N_26,In_2034);
or U2067 (N_2067,In_1085,N_829);
or U2068 (N_2068,N_1086,In_668);
nor U2069 (N_2069,In_275,N_578);
or U2070 (N_2070,N_493,N_712);
xor U2071 (N_2071,N_412,N_606);
nand U2072 (N_2072,N_766,In_1908);
nor U2073 (N_2073,N_1120,N_64);
xnor U2074 (N_2074,In_84,N_797);
nand U2075 (N_2075,N_264,N_363);
nor U2076 (N_2076,N_1192,In_779);
and U2077 (N_2077,In_2655,N_751);
nand U2078 (N_2078,N_791,N_136);
nor U2079 (N_2079,In_2538,N_325);
nor U2080 (N_2080,N_651,N_1164);
or U2081 (N_2081,N_5,In_447);
nand U2082 (N_2082,In_1088,N_818);
and U2083 (N_2083,In_1110,In_271);
xnor U2084 (N_2084,N_9,N_1051);
and U2085 (N_2085,N_144,In_492);
nor U2086 (N_2086,N_519,In_347);
xor U2087 (N_2087,N_114,N_256);
nand U2088 (N_2088,N_464,N_27);
xor U2089 (N_2089,N_525,In_1101);
nand U2090 (N_2090,In_1500,N_1105);
nor U2091 (N_2091,In_2170,N_889);
xor U2092 (N_2092,In_2335,N_747);
or U2093 (N_2093,N_121,N_995);
or U2094 (N_2094,N_437,In_1229);
nand U2095 (N_2095,N_553,N_620);
and U2096 (N_2096,N_684,N_128);
or U2097 (N_2097,N_943,N_353);
or U2098 (N_2098,N_297,In_1111);
nor U2099 (N_2099,N_217,N_346);
nand U2100 (N_2100,N_737,N_96);
and U2101 (N_2101,N_614,N_633);
and U2102 (N_2102,N_344,In_2936);
nor U2103 (N_2103,N_290,N_247);
and U2104 (N_2104,N_1152,In_1152);
xor U2105 (N_2105,In_1848,N_14);
xor U2106 (N_2106,N_1012,N_330);
or U2107 (N_2107,N_650,N_185);
and U2108 (N_2108,In_92,N_304);
xor U2109 (N_2109,N_1105,N_132);
nor U2110 (N_2110,N_1057,In_353);
nor U2111 (N_2111,N_535,N_473);
nand U2112 (N_2112,N_800,In_2074);
nor U2113 (N_2113,In_2647,In_2042);
or U2114 (N_2114,N_978,N_887);
and U2115 (N_2115,In_2010,N_257);
nand U2116 (N_2116,N_183,In_1892);
or U2117 (N_2117,N_966,N_362);
xor U2118 (N_2118,N_60,N_310);
nand U2119 (N_2119,N_582,In_674);
xor U2120 (N_2120,N_279,In_1804);
nand U2121 (N_2121,In_2109,In_1497);
nand U2122 (N_2122,In_2347,In_2532);
or U2123 (N_2123,N_597,In_2195);
xor U2124 (N_2124,In_2288,N_399);
nand U2125 (N_2125,In_2602,N_365);
nor U2126 (N_2126,In_339,N_117);
nor U2127 (N_2127,In_114,N_471);
or U2128 (N_2128,N_791,N_550);
and U2129 (N_2129,In_64,N_455);
nand U2130 (N_2130,In_2825,N_1087);
nor U2131 (N_2131,In_2759,In_2843);
or U2132 (N_2132,N_1185,N_990);
nand U2133 (N_2133,In_2080,N_536);
or U2134 (N_2134,In_192,N_808);
and U2135 (N_2135,N_1099,N_497);
nor U2136 (N_2136,In_1052,In_452);
nand U2137 (N_2137,N_1063,N_313);
and U2138 (N_2138,N_148,N_915);
or U2139 (N_2139,In_2109,N_1016);
or U2140 (N_2140,N_255,In_1945);
xor U2141 (N_2141,N_789,N_280);
nor U2142 (N_2142,N_884,N_467);
nand U2143 (N_2143,In_2799,In_1036);
xor U2144 (N_2144,In_1313,In_19);
nor U2145 (N_2145,N_514,In_129);
or U2146 (N_2146,N_403,N_1185);
and U2147 (N_2147,N_816,N_431);
nor U2148 (N_2148,In_118,In_2192);
xor U2149 (N_2149,In_588,In_1405);
nand U2150 (N_2150,N_962,N_920);
and U2151 (N_2151,In_1864,N_1085);
xnor U2152 (N_2152,In_838,N_374);
and U2153 (N_2153,N_81,In_2840);
nand U2154 (N_2154,In_1972,In_679);
nand U2155 (N_2155,N_1114,In_2843);
or U2156 (N_2156,N_664,N_565);
and U2157 (N_2157,N_1068,In_2162);
and U2158 (N_2158,In_1432,N_233);
nor U2159 (N_2159,N_915,N_36);
xor U2160 (N_2160,N_396,N_95);
nor U2161 (N_2161,N_870,In_2529);
xor U2162 (N_2162,In_1086,N_1049);
nor U2163 (N_2163,In_939,In_1446);
nand U2164 (N_2164,In_601,N_941);
and U2165 (N_2165,N_480,In_655);
nor U2166 (N_2166,N_576,N_908);
and U2167 (N_2167,N_1037,N_103);
and U2168 (N_2168,In_1672,In_1849);
nand U2169 (N_2169,N_94,In_1811);
and U2170 (N_2170,N_721,In_2282);
and U2171 (N_2171,N_669,N_1189);
nand U2172 (N_2172,In_339,In_2700);
or U2173 (N_2173,N_10,In_943);
nand U2174 (N_2174,In_1961,N_209);
nor U2175 (N_2175,In_849,In_2106);
xnor U2176 (N_2176,N_92,N_525);
or U2177 (N_2177,N_596,N_128);
and U2178 (N_2178,N_3,N_1154);
or U2179 (N_2179,N_45,N_473);
nand U2180 (N_2180,N_765,N_299);
and U2181 (N_2181,N_586,In_1962);
xnor U2182 (N_2182,In_294,In_149);
nand U2183 (N_2183,N_181,N_728);
nor U2184 (N_2184,In_129,In_2510);
nand U2185 (N_2185,In_1870,N_1195);
nor U2186 (N_2186,N_795,N_583);
or U2187 (N_2187,In_2990,In_1272);
nand U2188 (N_2188,In_291,N_138);
nand U2189 (N_2189,N_6,In_2594);
nor U2190 (N_2190,In_2201,N_499);
xnor U2191 (N_2191,In_1076,N_357);
nand U2192 (N_2192,In_1650,N_734);
nor U2193 (N_2193,In_1097,N_119);
nand U2194 (N_2194,N_943,N_875);
and U2195 (N_2195,N_1136,N_600);
nand U2196 (N_2196,N_1077,N_237);
xnor U2197 (N_2197,N_262,In_2020);
nand U2198 (N_2198,In_296,N_1182);
and U2199 (N_2199,N_334,N_584);
or U2200 (N_2200,N_577,In_1291);
nor U2201 (N_2201,N_914,N_610);
nand U2202 (N_2202,In_1433,N_379);
nor U2203 (N_2203,In_149,N_240);
or U2204 (N_2204,N_595,N_31);
nor U2205 (N_2205,N_756,In_2041);
xnor U2206 (N_2206,N_94,N_755);
nor U2207 (N_2207,N_666,N_975);
nor U2208 (N_2208,N_49,In_604);
or U2209 (N_2209,N_406,N_1161);
and U2210 (N_2210,N_924,N_258);
and U2211 (N_2211,N_811,N_46);
or U2212 (N_2212,In_1480,In_1177);
nand U2213 (N_2213,N_797,N_1116);
nand U2214 (N_2214,N_534,N_213);
nor U2215 (N_2215,In_84,In_1403);
nand U2216 (N_2216,N_989,N_986);
nor U2217 (N_2217,N_1192,In_1647);
nand U2218 (N_2218,In_2444,N_312);
and U2219 (N_2219,In_2505,N_311);
nand U2220 (N_2220,N_1191,In_2303);
nor U2221 (N_2221,N_823,N_611);
nand U2222 (N_2222,N_536,N_1146);
nand U2223 (N_2223,In_336,N_256);
xor U2224 (N_2224,In_325,N_710);
xor U2225 (N_2225,N_745,N_915);
and U2226 (N_2226,N_106,N_738);
nand U2227 (N_2227,N_1109,N_123);
nand U2228 (N_2228,In_1214,N_543);
nor U2229 (N_2229,In_1229,N_643);
or U2230 (N_2230,In_92,In_471);
nor U2231 (N_2231,In_2528,N_32);
and U2232 (N_2232,In_695,N_1045);
nor U2233 (N_2233,In_1229,N_883);
nor U2234 (N_2234,N_756,N_1114);
and U2235 (N_2235,In_215,N_257);
nor U2236 (N_2236,In_2441,N_639);
or U2237 (N_2237,In_1029,N_931);
nand U2238 (N_2238,In_169,In_1245);
nor U2239 (N_2239,N_1144,N_1114);
nor U2240 (N_2240,N_68,N_1196);
nor U2241 (N_2241,In_0,N_815);
nand U2242 (N_2242,In_665,In_1121);
xnor U2243 (N_2243,N_243,In_665);
nand U2244 (N_2244,In_191,In_2999);
nor U2245 (N_2245,N_1142,N_688);
or U2246 (N_2246,N_301,N_299);
nor U2247 (N_2247,N_724,In_722);
nand U2248 (N_2248,In_2298,N_699);
nand U2249 (N_2249,N_1028,In_311);
nand U2250 (N_2250,In_2322,In_1061);
or U2251 (N_2251,N_816,In_1089);
nor U2252 (N_2252,N_877,N_704);
nor U2253 (N_2253,N_540,In_1599);
nand U2254 (N_2254,N_536,N_612);
nand U2255 (N_2255,N_1009,N_183);
nand U2256 (N_2256,In_2759,N_965);
xnor U2257 (N_2257,N_238,In_252);
and U2258 (N_2258,N_844,In_618);
nor U2259 (N_2259,In_2763,N_332);
nand U2260 (N_2260,N_431,N_1162);
and U2261 (N_2261,N_57,N_74);
nor U2262 (N_2262,N_324,N_1006);
nand U2263 (N_2263,N_388,In_655);
and U2264 (N_2264,In_1674,N_1063);
xor U2265 (N_2265,In_1924,In_1069);
or U2266 (N_2266,In_2007,N_46);
or U2267 (N_2267,N_520,N_477);
and U2268 (N_2268,N_115,N_998);
nor U2269 (N_2269,N_565,N_651);
xnor U2270 (N_2270,In_292,N_451);
xor U2271 (N_2271,N_455,In_1810);
nor U2272 (N_2272,In_394,In_1559);
xnor U2273 (N_2273,N_299,In_2374);
or U2274 (N_2274,N_1193,N_1172);
and U2275 (N_2275,N_816,N_412);
and U2276 (N_2276,N_943,N_226);
nor U2277 (N_2277,N_928,N_740);
and U2278 (N_2278,N_1170,N_625);
xnor U2279 (N_2279,N_1136,N_928);
and U2280 (N_2280,N_8,In_2784);
or U2281 (N_2281,N_906,N_878);
and U2282 (N_2282,N_308,N_1053);
and U2283 (N_2283,N_379,N_653);
nor U2284 (N_2284,In_831,N_624);
nand U2285 (N_2285,N_1114,In_1110);
or U2286 (N_2286,In_1403,N_1172);
and U2287 (N_2287,In_2382,N_469);
and U2288 (N_2288,In_2007,N_953);
and U2289 (N_2289,N_451,In_1388);
and U2290 (N_2290,N_156,N_439);
and U2291 (N_2291,N_1003,N_691);
and U2292 (N_2292,N_306,N_975);
nand U2293 (N_2293,N_1147,In_2356);
nor U2294 (N_2294,N_1106,N_711);
nand U2295 (N_2295,In_868,N_998);
or U2296 (N_2296,In_2341,N_1157);
xnor U2297 (N_2297,N_735,In_2796);
nand U2298 (N_2298,In_2487,N_338);
nor U2299 (N_2299,N_835,N_762);
xor U2300 (N_2300,In_343,N_621);
nor U2301 (N_2301,N_107,N_1081);
xnor U2302 (N_2302,N_612,In_68);
or U2303 (N_2303,N_74,N_83);
nand U2304 (N_2304,In_934,In_1142);
and U2305 (N_2305,N_770,In_576);
and U2306 (N_2306,N_443,N_4);
or U2307 (N_2307,In_1475,In_1974);
xor U2308 (N_2308,In_786,N_100);
and U2309 (N_2309,In_2793,N_769);
or U2310 (N_2310,N_142,N_756);
or U2311 (N_2311,N_297,In_979);
nand U2312 (N_2312,N_866,N_439);
nor U2313 (N_2313,N_1085,In_1650);
nor U2314 (N_2314,N_1096,In_1712);
and U2315 (N_2315,N_2,N_488);
xor U2316 (N_2316,In_2284,N_135);
nand U2317 (N_2317,N_748,In_291);
nand U2318 (N_2318,N_891,N_353);
nand U2319 (N_2319,N_551,In_912);
or U2320 (N_2320,N_530,N_577);
xnor U2321 (N_2321,N_438,N_197);
xor U2322 (N_2322,N_604,N_207);
nand U2323 (N_2323,N_142,N_233);
nand U2324 (N_2324,N_802,N_69);
nor U2325 (N_2325,N_580,N_610);
and U2326 (N_2326,N_604,In_2842);
nand U2327 (N_2327,N_863,N_535);
nor U2328 (N_2328,N_247,N_22);
and U2329 (N_2329,N_382,In_2891);
nand U2330 (N_2330,N_793,N_262);
and U2331 (N_2331,N_877,In_2575);
or U2332 (N_2332,N_137,N_926);
nor U2333 (N_2333,In_690,N_905);
nor U2334 (N_2334,In_2878,N_312);
nand U2335 (N_2335,In_786,N_279);
and U2336 (N_2336,In_2914,N_13);
xor U2337 (N_2337,N_1026,N_1044);
or U2338 (N_2338,N_826,N_657);
xor U2339 (N_2339,N_397,N_15);
or U2340 (N_2340,N_860,N_219);
nor U2341 (N_2341,N_357,In_934);
and U2342 (N_2342,In_1607,In_2621);
nand U2343 (N_2343,N_732,In_1152);
xnor U2344 (N_2344,In_2869,In_1695);
or U2345 (N_2345,N_948,N_685);
or U2346 (N_2346,N_607,In_1962);
nor U2347 (N_2347,In_2601,In_1658);
and U2348 (N_2348,N_1137,In_2539);
and U2349 (N_2349,N_911,N_746);
nand U2350 (N_2350,N_335,In_1724);
xor U2351 (N_2351,N_1172,In_2910);
xor U2352 (N_2352,N_125,In_1659);
xor U2353 (N_2353,N_614,In_681);
and U2354 (N_2354,In_943,In_2154);
nand U2355 (N_2355,In_953,In_2575);
and U2356 (N_2356,In_1667,In_1110);
or U2357 (N_2357,In_1403,In_2641);
and U2358 (N_2358,N_156,N_963);
nor U2359 (N_2359,N_566,In_668);
xor U2360 (N_2360,In_958,N_577);
and U2361 (N_2361,In_934,N_308);
nand U2362 (N_2362,N_887,In_1101);
and U2363 (N_2363,In_804,N_34);
nand U2364 (N_2364,N_206,N_957);
nor U2365 (N_2365,N_1113,In_2993);
nor U2366 (N_2366,In_642,In_134);
nor U2367 (N_2367,N_943,N_916);
and U2368 (N_2368,N_585,N_381);
xnor U2369 (N_2369,N_191,N_469);
or U2370 (N_2370,N_718,In_64);
and U2371 (N_2371,N_1114,In_2397);
nand U2372 (N_2372,N_530,In_1607);
xor U2373 (N_2373,N_814,N_232);
xnor U2374 (N_2374,N_1174,N_330);
or U2375 (N_2375,N_679,In_2703);
xnor U2376 (N_2376,N_136,In_1052);
or U2377 (N_2377,In_743,N_998);
nor U2378 (N_2378,N_739,In_172);
or U2379 (N_2379,N_948,In_2647);
nand U2380 (N_2380,N_419,N_1044);
nor U2381 (N_2381,In_129,In_1730);
or U2382 (N_2382,In_262,N_753);
xor U2383 (N_2383,In_1024,In_2154);
or U2384 (N_2384,N_417,In_281);
nor U2385 (N_2385,N_168,In_2284);
or U2386 (N_2386,N_364,In_2843);
nand U2387 (N_2387,N_301,In_1082);
and U2388 (N_2388,N_1173,N_796);
and U2389 (N_2389,N_128,N_468);
and U2390 (N_2390,N_849,N_907);
or U2391 (N_2391,In_882,N_1162);
and U2392 (N_2392,In_1715,N_75);
or U2393 (N_2393,N_606,N_168);
and U2394 (N_2394,N_981,N_432);
nand U2395 (N_2395,N_122,N_879);
or U2396 (N_2396,N_22,N_481);
or U2397 (N_2397,N_262,N_997);
xor U2398 (N_2398,N_97,In_100);
and U2399 (N_2399,N_352,N_65);
nor U2400 (N_2400,N_1854,N_1525);
or U2401 (N_2401,N_1561,N_2181);
and U2402 (N_2402,N_2260,N_1536);
or U2403 (N_2403,N_1754,N_2092);
and U2404 (N_2404,N_2024,N_2118);
and U2405 (N_2405,N_2077,N_2262);
xnor U2406 (N_2406,N_1467,N_1821);
nand U2407 (N_2407,N_1229,N_2240);
xor U2408 (N_2408,N_1443,N_1303);
and U2409 (N_2409,N_2272,N_2352);
or U2410 (N_2410,N_1939,N_1394);
or U2411 (N_2411,N_2245,N_1699);
and U2412 (N_2412,N_1573,N_1970);
nor U2413 (N_2413,N_1825,N_2366);
nor U2414 (N_2414,N_1585,N_1709);
nand U2415 (N_2415,N_1982,N_2135);
xnor U2416 (N_2416,N_1484,N_2027);
and U2417 (N_2417,N_1824,N_1803);
or U2418 (N_2418,N_1514,N_1478);
xnor U2419 (N_2419,N_1398,N_1785);
and U2420 (N_2420,N_2259,N_1912);
xnor U2421 (N_2421,N_1847,N_1539);
nand U2422 (N_2422,N_1532,N_1203);
nand U2423 (N_2423,N_2398,N_2299);
or U2424 (N_2424,N_1527,N_1374);
nand U2425 (N_2425,N_2389,N_1746);
and U2426 (N_2426,N_1321,N_2195);
and U2427 (N_2427,N_2247,N_1818);
xnor U2428 (N_2428,N_2103,N_2007);
and U2429 (N_2429,N_1280,N_1548);
or U2430 (N_2430,N_1352,N_2186);
or U2431 (N_2431,N_1931,N_1545);
nand U2432 (N_2432,N_1780,N_1389);
nand U2433 (N_2433,N_1764,N_1950);
xor U2434 (N_2434,N_1210,N_1453);
nand U2435 (N_2435,N_1876,N_1397);
nand U2436 (N_2436,N_2091,N_1874);
xnor U2437 (N_2437,N_1889,N_1362);
and U2438 (N_2438,N_2095,N_2256);
nor U2439 (N_2439,N_1832,N_2392);
nand U2440 (N_2440,N_1762,N_2314);
nand U2441 (N_2441,N_1786,N_1700);
xnor U2442 (N_2442,N_1864,N_1972);
nor U2443 (N_2443,N_1396,N_2266);
nor U2444 (N_2444,N_1510,N_1259);
or U2445 (N_2445,N_2263,N_1835);
nand U2446 (N_2446,N_2222,N_2101);
nand U2447 (N_2447,N_1602,N_1424);
and U2448 (N_2448,N_1325,N_2242);
nand U2449 (N_2449,N_1610,N_1807);
xnor U2450 (N_2450,N_1621,N_1761);
nor U2451 (N_2451,N_1264,N_1569);
xor U2452 (N_2452,N_1246,N_1223);
xnor U2453 (N_2453,N_2133,N_2284);
nor U2454 (N_2454,N_1671,N_1468);
nor U2455 (N_2455,N_1712,N_1644);
and U2456 (N_2456,N_1693,N_1348);
nand U2457 (N_2457,N_1372,N_1523);
xor U2458 (N_2458,N_2105,N_2002);
or U2459 (N_2459,N_1886,N_2224);
and U2460 (N_2460,N_1645,N_2031);
xor U2461 (N_2461,N_1784,N_1639);
and U2462 (N_2462,N_1407,N_1216);
nor U2463 (N_2463,N_2173,N_2151);
nor U2464 (N_2464,N_1937,N_1568);
nand U2465 (N_2465,N_1476,N_1338);
xnor U2466 (N_2466,N_1625,N_1309);
nand U2467 (N_2467,N_2303,N_1350);
nand U2468 (N_2468,N_1479,N_1257);
or U2469 (N_2469,N_1885,N_1429);
xnor U2470 (N_2470,N_2042,N_1791);
nand U2471 (N_2471,N_2055,N_1675);
nor U2472 (N_2472,N_1236,N_1966);
or U2473 (N_2473,N_1243,N_1204);
and U2474 (N_2474,N_2276,N_1355);
xnor U2475 (N_2475,N_1540,N_1946);
nand U2476 (N_2476,N_1261,N_2280);
or U2477 (N_2477,N_2258,N_1595);
nor U2478 (N_2478,N_1522,N_1307);
xor U2479 (N_2479,N_2221,N_1969);
and U2480 (N_2480,N_1714,N_2023);
nor U2481 (N_2481,N_1924,N_1562);
xor U2482 (N_2482,N_2033,N_2124);
nor U2483 (N_2483,N_1418,N_2269);
nor U2484 (N_2484,N_1680,N_1575);
xnor U2485 (N_2485,N_1444,N_1715);
xor U2486 (N_2486,N_1778,N_2342);
nor U2487 (N_2487,N_1403,N_1883);
and U2488 (N_2488,N_2387,N_1538);
and U2489 (N_2489,N_1270,N_2008);
and U2490 (N_2490,N_1952,N_1341);
xor U2491 (N_2491,N_2134,N_1361);
or U2492 (N_2492,N_1357,N_2140);
nor U2493 (N_2493,N_2056,N_2312);
nor U2494 (N_2494,N_1853,N_2047);
or U2495 (N_2495,N_1892,N_2166);
xnor U2496 (N_2496,N_2097,N_2217);
nor U2497 (N_2497,N_1749,N_1209);
and U2498 (N_2498,N_2393,N_1776);
and U2499 (N_2499,N_1505,N_1301);
nor U2500 (N_2500,N_2106,N_1855);
xnor U2501 (N_2501,N_1928,N_1472);
or U2502 (N_2502,N_1897,N_1457);
nand U2503 (N_2503,N_1381,N_1419);
xnor U2504 (N_2504,N_2104,N_1801);
and U2505 (N_2505,N_1579,N_1686);
or U2506 (N_2506,N_2277,N_1289);
xor U2507 (N_2507,N_1668,N_2239);
nor U2508 (N_2508,N_1382,N_1617);
nor U2509 (N_2509,N_1238,N_1517);
and U2510 (N_2510,N_1490,N_1706);
nor U2511 (N_2511,N_1542,N_2063);
and U2512 (N_2512,N_1211,N_1449);
nand U2513 (N_2513,N_1475,N_1987);
xnor U2514 (N_2514,N_1239,N_1796);
or U2515 (N_2515,N_1446,N_1851);
and U2516 (N_2516,N_1566,N_2204);
xor U2517 (N_2517,N_1380,N_2309);
nor U2518 (N_2518,N_1705,N_2359);
nand U2519 (N_2519,N_1918,N_1624);
nand U2520 (N_2520,N_1438,N_1500);
and U2521 (N_2521,N_1554,N_2232);
and U2522 (N_2522,N_2174,N_1513);
nand U2523 (N_2523,N_2189,N_2330);
nand U2524 (N_2524,N_2334,N_1232);
or U2525 (N_2525,N_1976,N_1858);
or U2526 (N_2526,N_1465,N_1499);
nor U2527 (N_2527,N_1364,N_1590);
xor U2528 (N_2528,N_1725,N_1412);
and U2529 (N_2529,N_2046,N_2148);
and U2530 (N_2530,N_1531,N_2285);
nand U2531 (N_2531,N_2198,N_1423);
nor U2532 (N_2532,N_1766,N_2172);
xor U2533 (N_2533,N_1685,N_1681);
or U2534 (N_2534,N_1632,N_2053);
nor U2535 (N_2535,N_2257,N_1649);
or U2536 (N_2536,N_1451,N_1642);
or U2537 (N_2537,N_1752,N_1218);
or U2538 (N_2538,N_1616,N_1960);
nand U2539 (N_2539,N_1250,N_1284);
or U2540 (N_2540,N_2264,N_1529);
nor U2541 (N_2541,N_2391,N_1552);
and U2542 (N_2542,N_2094,N_1275);
nand U2543 (N_2543,N_2226,N_1676);
xor U2544 (N_2544,N_1589,N_2178);
or U2545 (N_2545,N_1417,N_1300);
nor U2546 (N_2546,N_1330,N_1359);
and U2547 (N_2547,N_1421,N_1975);
nand U2548 (N_2548,N_2337,N_1635);
xor U2549 (N_2549,N_1980,N_1323);
nand U2550 (N_2550,N_1800,N_1502);
and U2551 (N_2551,N_1326,N_1497);
nor U2552 (N_2552,N_1891,N_2233);
and U2553 (N_2553,N_1533,N_1650);
and U2554 (N_2554,N_1228,N_1739);
nand U2555 (N_2555,N_1290,N_2220);
nand U2556 (N_2556,N_1979,N_1599);
nand U2557 (N_2557,N_1734,N_2317);
or U2558 (N_2558,N_1881,N_1434);
nand U2559 (N_2559,N_2003,N_1385);
and U2560 (N_2560,N_2293,N_1692);
or U2561 (N_2561,N_2098,N_2193);
xnor U2562 (N_2562,N_1814,N_1276);
or U2563 (N_2563,N_2339,N_2304);
or U2564 (N_2564,N_1445,N_1311);
xor U2565 (N_2565,N_1859,N_2160);
nand U2566 (N_2566,N_2144,N_2397);
nor U2567 (N_2567,N_1313,N_1619);
nand U2568 (N_2568,N_1893,N_1741);
nand U2569 (N_2569,N_2292,N_1657);
and U2570 (N_2570,N_2017,N_2390);
nor U2571 (N_2571,N_2318,N_2347);
xor U2572 (N_2572,N_1331,N_2231);
xnor U2573 (N_2573,N_1557,N_1788);
nor U2574 (N_2574,N_2212,N_2321);
and U2575 (N_2575,N_1383,N_1318);
nor U2576 (N_2576,N_1875,N_1971);
nand U2577 (N_2577,N_2335,N_1600);
xor U2578 (N_2578,N_1750,N_2128);
xnor U2579 (N_2579,N_1528,N_1763);
or U2580 (N_2580,N_1813,N_1981);
and U2581 (N_2581,N_1420,N_1721);
and U2582 (N_2582,N_1314,N_1272);
nand U2583 (N_2583,N_1526,N_2332);
and U2584 (N_2584,N_2032,N_1368);
nand U2585 (N_2585,N_1636,N_1690);
xnor U2586 (N_2586,N_2227,N_1634);
and U2587 (N_2587,N_1217,N_1905);
nor U2588 (N_2588,N_1388,N_2274);
and U2589 (N_2589,N_2300,N_1578);
xnor U2590 (N_2590,N_1335,N_2307);
nor U2591 (N_2591,N_1392,N_2122);
or U2592 (N_2592,N_2080,N_2016);
or U2593 (N_2593,N_1244,N_1494);
or U2594 (N_2594,N_1425,N_1765);
nor U2595 (N_2595,N_2155,N_2015);
nor U2596 (N_2596,N_1833,N_2071);
nand U2597 (N_2597,N_2061,N_1406);
or U2598 (N_2598,N_1286,N_1748);
nor U2599 (N_2599,N_2371,N_1862);
nand U2600 (N_2600,N_2286,N_1456);
xor U2601 (N_2601,N_1201,N_1393);
and U2602 (N_2602,N_1867,N_1574);
nor U2603 (N_2603,N_1839,N_1996);
and U2604 (N_2604,N_1718,N_1790);
nand U2605 (N_2605,N_1520,N_1292);
xor U2606 (N_2606,N_2291,N_1304);
nor U2607 (N_2607,N_2281,N_1701);
nand U2608 (N_2608,N_2019,N_1684);
nor U2609 (N_2609,N_1435,N_1273);
and U2610 (N_2610,N_1237,N_1267);
xnor U2611 (N_2611,N_2325,N_1334);
and U2612 (N_2612,N_1911,N_1731);
nand U2613 (N_2613,N_1781,N_1998);
nor U2614 (N_2614,N_1751,N_1805);
or U2615 (N_2615,N_2111,N_1870);
xnor U2616 (N_2616,N_1955,N_2057);
and U2617 (N_2617,N_2184,N_1920);
and U2618 (N_2618,N_1951,N_2375);
xor U2619 (N_2619,N_1293,N_2253);
xnor U2620 (N_2620,N_2289,N_1852);
xor U2621 (N_2621,N_1450,N_2099);
or U2622 (N_2622,N_1391,N_1333);
and U2623 (N_2623,N_1985,N_1269);
xnor U2624 (N_2624,N_1507,N_1654);
nor U2625 (N_2625,N_1447,N_2038);
nand U2626 (N_2626,N_1935,N_1459);
and U2627 (N_2627,N_2117,N_2343);
nand U2628 (N_2628,N_1949,N_1667);
xor U2629 (N_2629,N_1506,N_1551);
xor U2630 (N_2630,N_2076,N_1241);
and U2631 (N_2631,N_2244,N_1227);
and U2632 (N_2632,N_1729,N_2197);
nor U2633 (N_2633,N_2176,N_1328);
and U2634 (N_2634,N_2320,N_1869);
nor U2635 (N_2635,N_1298,N_1519);
nor U2636 (N_2636,N_1547,N_1909);
or U2637 (N_2637,N_1512,N_2062);
and U2638 (N_2638,N_2014,N_1782);
nand U2639 (N_2639,N_1860,N_2145);
nor U2640 (N_2640,N_1888,N_1627);
xnor U2641 (N_2641,N_1698,N_1653);
nor U2642 (N_2642,N_1669,N_2079);
or U2643 (N_2643,N_1226,N_1959);
and U2644 (N_2644,N_1572,N_2183);
nor U2645 (N_2645,N_1903,N_1493);
nand U2646 (N_2646,N_1956,N_2029);
nor U2647 (N_2647,N_1367,N_1717);
and U2648 (N_2648,N_1295,N_1884);
nand U2649 (N_2649,N_1626,N_1342);
nor U2650 (N_2650,N_1622,N_1486);
and U2651 (N_2651,N_1454,N_1549);
xnor U2652 (N_2652,N_1999,N_2311);
nand U2653 (N_2653,N_2064,N_2261);
xnor U2654 (N_2654,N_1953,N_1466);
or U2655 (N_2655,N_2011,N_2030);
xor U2656 (N_2656,N_1936,N_2187);
nand U2657 (N_2657,N_1743,N_2351);
or U2658 (N_2658,N_2191,N_1377);
nor U2659 (N_2659,N_2288,N_1277);
and U2660 (N_2660,N_2157,N_1861);
and U2661 (N_2661,N_2296,N_1433);
nand U2662 (N_2662,N_2170,N_1254);
and U2663 (N_2663,N_2090,N_1887);
or U2664 (N_2664,N_1802,N_1260);
or U2665 (N_2665,N_2070,N_1319);
nand U2666 (N_2666,N_2177,N_2179);
xnor U2667 (N_2667,N_2346,N_2340);
nor U2668 (N_2668,N_1401,N_1722);
or U2669 (N_2669,N_2113,N_1395);
or U2670 (N_2670,N_2372,N_1612);
nor U2671 (N_2671,N_1212,N_2093);
nor U2672 (N_2672,N_1558,N_1735);
nor U2673 (N_2673,N_1808,N_1410);
nor U2674 (N_2674,N_1405,N_1591);
xor U2675 (N_2675,N_1643,N_1866);
and U2676 (N_2676,N_1235,N_2308);
nand U2677 (N_2677,N_1274,N_2035);
nand U2678 (N_2678,N_2089,N_1934);
and U2679 (N_2679,N_1683,N_1206);
nor U2680 (N_2680,N_1983,N_2147);
nand U2681 (N_2681,N_1580,N_2238);
and U2682 (N_2682,N_1581,N_1485);
nand U2683 (N_2683,N_1759,N_1598);
nor U2684 (N_2684,N_1637,N_1830);
or U2685 (N_2685,N_1663,N_2112);
and U2686 (N_2686,N_2230,N_1379);
and U2687 (N_2687,N_1899,N_1550);
xor U2688 (N_2688,N_1670,N_1365);
and U2689 (N_2689,N_2049,N_1770);
and U2690 (N_2690,N_2078,N_1305);
xnor U2691 (N_2691,N_2202,N_1332);
xor U2692 (N_2692,N_1339,N_2283);
nand U2693 (N_2693,N_2206,N_1652);
xor U2694 (N_2694,N_1521,N_1422);
xor U2695 (N_2695,N_1200,N_1838);
xnor U2696 (N_2696,N_1930,N_1471);
nor U2697 (N_2697,N_2158,N_2310);
and U2698 (N_2698,N_1409,N_1256);
or U2699 (N_2699,N_1224,N_2192);
nor U2700 (N_2700,N_1944,N_1702);
nor U2701 (N_2701,N_1515,N_1214);
nand U2702 (N_2702,N_1390,N_1358);
and U2703 (N_2703,N_1707,N_1263);
and U2704 (N_2704,N_2109,N_1288);
xor U2705 (N_2705,N_2378,N_1964);
nand U2706 (N_2706,N_1678,N_1340);
nand U2707 (N_2707,N_1504,N_1556);
nor U2708 (N_2708,N_2010,N_1315);
and U2709 (N_2709,N_1221,N_2004);
nor U2710 (N_2710,N_2246,N_1268);
or U2711 (N_2711,N_1695,N_2058);
xor U2712 (N_2712,N_1594,N_2126);
xor U2713 (N_2713,N_1220,N_1879);
or U2714 (N_2714,N_1414,N_1655);
or U2715 (N_2715,N_1961,N_1872);
and U2716 (N_2716,N_2075,N_2153);
and U2717 (N_2717,N_1795,N_1842);
nand U2718 (N_2718,N_1925,N_1817);
nor U2719 (N_2719,N_1916,N_1363);
and U2720 (N_2720,N_2306,N_1582);
or U2721 (N_2721,N_2249,N_2005);
nor U2722 (N_2722,N_2044,N_1845);
nor U2723 (N_2723,N_1296,N_1458);
xor U2724 (N_2724,N_1452,N_2265);
nor U2725 (N_2725,N_1461,N_1620);
xnor U2726 (N_2726,N_1809,N_2059);
nor U2727 (N_2727,N_2349,N_1386);
and U2728 (N_2728,N_2395,N_1738);
or U2729 (N_2729,N_2301,N_1427);
nor U2730 (N_2730,N_1587,N_2209);
xor U2731 (N_2731,N_1674,N_2255);
nand U2732 (N_2732,N_1601,N_1588);
xnor U2733 (N_2733,N_1481,N_2355);
xnor U2734 (N_2734,N_2287,N_1482);
nor U2735 (N_2735,N_1371,N_1828);
or U2736 (N_2736,N_1509,N_1400);
or U2737 (N_2737,N_1492,N_1753);
and U2738 (N_2738,N_1518,N_2013);
nand U2739 (N_2739,N_2386,N_2036);
or U2740 (N_2740,N_2048,N_2368);
nand U2741 (N_2741,N_2020,N_2107);
or U2742 (N_2742,N_1496,N_2074);
and U2743 (N_2743,N_2141,N_1844);
or U2744 (N_2744,N_1878,N_2188);
nand U2745 (N_2745,N_2248,N_1769);
and U2746 (N_2746,N_1963,N_2329);
xnor U2747 (N_2747,N_1720,N_1757);
xor U2748 (N_2748,N_1495,N_2116);
and U2749 (N_2749,N_1498,N_2072);
and U2750 (N_2750,N_1555,N_1399);
and U2751 (N_2751,N_2380,N_1863);
nand U2752 (N_2752,N_2379,N_2132);
nand U2753 (N_2753,N_2051,N_2367);
nand U2754 (N_2754,N_1902,N_1733);
or U2755 (N_2755,N_1648,N_1251);
nand U2756 (N_2756,N_2373,N_1322);
xnor U2757 (N_2757,N_1242,N_1213);
nand U2758 (N_2758,N_1689,N_1846);
or U2759 (N_2759,N_2073,N_2119);
xnor U2760 (N_2760,N_2376,N_2146);
and U2761 (N_2761,N_1868,N_1317);
and U2762 (N_2762,N_2382,N_1856);
xor U2763 (N_2763,N_1793,N_1724);
and U2764 (N_2764,N_1378,N_2383);
or U2765 (N_2765,N_2298,N_1834);
and U2766 (N_2766,N_1219,N_1615);
xor U2767 (N_2767,N_2137,N_1687);
xor U2768 (N_2768,N_2388,N_1345);
nor U2769 (N_2769,N_1907,N_2001);
xnor U2770 (N_2770,N_1503,N_2377);
or U2771 (N_2771,N_2028,N_1302);
nand U2772 (N_2772,N_2012,N_2052);
or U2773 (N_2773,N_1986,N_2254);
nand U2774 (N_2774,N_1815,N_2088);
nor U2775 (N_2775,N_1387,N_1660);
and U2776 (N_2776,N_2384,N_2152);
or U2777 (N_2777,N_1993,N_1994);
and U2778 (N_2778,N_1984,N_2194);
nand U2779 (N_2779,N_1437,N_1997);
nor U2780 (N_2780,N_1697,N_1758);
nand U2781 (N_2781,N_1898,N_1730);
or U2782 (N_2782,N_1583,N_1416);
or U2783 (N_2783,N_1929,N_1534);
and U2784 (N_2784,N_1408,N_1491);
nor U2785 (N_2785,N_2136,N_2305);
and U2786 (N_2786,N_1646,N_1265);
nor U2787 (N_2787,N_2139,N_1880);
xnor U2788 (N_2788,N_1932,N_2279);
nand U2789 (N_2789,N_2115,N_1941);
xnor U2790 (N_2790,N_1415,N_2009);
xnor U2791 (N_2791,N_1618,N_2295);
nor U2792 (N_2792,N_1316,N_1436);
nor U2793 (N_2793,N_1771,N_1320);
nand U2794 (N_2794,N_1366,N_1603);
and U2795 (N_2795,N_1560,N_2225);
nor U2796 (N_2796,N_1576,N_2114);
nor U2797 (N_2797,N_1727,N_1543);
nor U2798 (N_2798,N_1508,N_1823);
or U2799 (N_2799,N_1455,N_1673);
nor U2800 (N_2800,N_1567,N_1922);
nor U2801 (N_2801,N_1252,N_1713);
nand U2802 (N_2802,N_1662,N_1719);
nor U2803 (N_2803,N_1747,N_1439);
xor U2804 (N_2804,N_2338,N_1797);
nor U2805 (N_2805,N_2243,N_1370);
nand U2806 (N_2806,N_2370,N_1255);
xor U2807 (N_2807,N_1651,N_2081);
nand U2808 (N_2808,N_2327,N_2165);
or U2809 (N_2809,N_1404,N_2333);
or U2810 (N_2810,N_1816,N_1351);
xnor U2811 (N_2811,N_2237,N_2161);
and U2812 (N_2812,N_2026,N_1728);
nor U2813 (N_2813,N_2040,N_2069);
and U2814 (N_2814,N_2396,N_2313);
and U2815 (N_2815,N_2282,N_1544);
and U2816 (N_2816,N_2271,N_2235);
nor U2817 (N_2817,N_1977,N_2201);
and U2818 (N_2818,N_1921,N_2083);
nor U2819 (N_2819,N_2328,N_1462);
and U2820 (N_2820,N_1926,N_1877);
nand U2821 (N_2821,N_1894,N_1710);
xnor U2822 (N_2822,N_1756,N_1487);
xor U2823 (N_2823,N_1353,N_1957);
nand U2824 (N_2824,N_1248,N_2065);
and U2825 (N_2825,N_1948,N_1774);
and U2826 (N_2826,N_2360,N_2316);
nand U2827 (N_2827,N_1283,N_1895);
or U2828 (N_2828,N_2290,N_1772);
and U2829 (N_2829,N_2348,N_1850);
or U2830 (N_2830,N_1943,N_1773);
nand U2831 (N_2831,N_1777,N_1460);
and U2832 (N_2832,N_2207,N_2034);
nand U2833 (N_2833,N_1384,N_1967);
or U2834 (N_2834,N_1240,N_2068);
nand U2835 (N_2835,N_1822,N_2060);
or U2836 (N_2836,N_1463,N_2050);
or U2837 (N_2837,N_2143,N_1428);
xor U2838 (N_2838,N_1768,N_1278);
nor U2839 (N_2839,N_1740,N_1840);
nand U2840 (N_2840,N_2037,N_1890);
nor U2841 (N_2841,N_2341,N_2223);
nand U2842 (N_2842,N_2218,N_1604);
or U2843 (N_2843,N_2022,N_2219);
nand U2844 (N_2844,N_1611,N_1608);
or U2845 (N_2845,N_1630,N_2350);
xor U2846 (N_2846,N_1647,N_1716);
nor U2847 (N_2847,N_2067,N_1375);
xnor U2848 (N_2848,N_1470,N_1691);
nor U2849 (N_2849,N_1473,N_1836);
nor U2850 (N_2850,N_1792,N_1799);
nor U2851 (N_2851,N_1613,N_2154);
and U2852 (N_2852,N_2162,N_1837);
xnor U2853 (N_2853,N_1688,N_2381);
and U2854 (N_2854,N_1440,N_1933);
nand U2855 (N_2855,N_2267,N_1592);
xor U2856 (N_2856,N_2123,N_1411);
nand U2857 (N_2857,N_2125,N_1991);
nor U2858 (N_2858,N_2041,N_1990);
nor U2859 (N_2859,N_1742,N_1281);
nor U2860 (N_2860,N_2043,N_2211);
nor U2861 (N_2861,N_2210,N_2365);
nand U2862 (N_2862,N_2324,N_1570);
or U2863 (N_2863,N_1843,N_1628);
nor U2864 (N_2864,N_2163,N_2180);
or U2865 (N_2865,N_2039,N_1480);
nand U2866 (N_2866,N_1349,N_2363);
and U2867 (N_2867,N_1605,N_1992);
and U2868 (N_2868,N_1919,N_1344);
nand U2869 (N_2869,N_1343,N_1896);
xor U2870 (N_2870,N_2190,N_2294);
and U2871 (N_2871,N_1442,N_2167);
nor U2872 (N_2872,N_1483,N_1820);
or U2873 (N_2873,N_2086,N_2213);
xor U2874 (N_2874,N_1285,N_1917);
and U2875 (N_2875,N_2369,N_1658);
and U2876 (N_2876,N_2362,N_2268);
or U2877 (N_2877,N_2364,N_1641);
xor U2878 (N_2878,N_1369,N_1938);
xor U2879 (N_2879,N_1806,N_1559);
xor U2880 (N_2880,N_1553,N_1287);
nand U2881 (N_2881,N_1231,N_2149);
xnor U2882 (N_2882,N_1222,N_1535);
xnor U2883 (N_2883,N_1913,N_2121);
xnor U2884 (N_2884,N_2229,N_1811);
xnor U2885 (N_2885,N_2150,N_1910);
xor U2886 (N_2886,N_2045,N_2142);
and U2887 (N_2887,N_1789,N_2129);
or U2888 (N_2888,N_2021,N_2241);
xnor U2889 (N_2889,N_1312,N_1665);
and U2890 (N_2890,N_1812,N_1477);
or U2891 (N_2891,N_1848,N_1488);
or U2892 (N_2892,N_1631,N_1989);
or U2893 (N_2893,N_1965,N_2345);
nand U2894 (N_2894,N_2196,N_2385);
and U2895 (N_2895,N_2322,N_1623);
and U2896 (N_2896,N_1474,N_1373);
xnor U2897 (N_2897,N_2236,N_2171);
nand U2898 (N_2898,N_2358,N_2275);
and U2899 (N_2899,N_2159,N_1376);
and U2900 (N_2900,N_2326,N_2130);
and U2901 (N_2901,N_1464,N_1247);
nor U2902 (N_2902,N_2138,N_1233);
xnor U2903 (N_2903,N_2164,N_1208);
and U2904 (N_2904,N_2084,N_1230);
nand U2905 (N_2905,N_2234,N_1779);
nand U2906 (N_2906,N_1324,N_1974);
and U2907 (N_2907,N_1978,N_1565);
nand U2908 (N_2908,N_1968,N_1787);
and U2909 (N_2909,N_1694,N_1266);
nand U2910 (N_2910,N_2208,N_2100);
nand U2911 (N_2911,N_1873,N_1432);
nor U2912 (N_2912,N_2252,N_2315);
xor U2913 (N_2913,N_2302,N_1546);
nor U2914 (N_2914,N_1829,N_1672);
nor U2915 (N_2915,N_2025,N_2354);
nor U2916 (N_2916,N_2102,N_1633);
and U2917 (N_2917,N_2323,N_1947);
nor U2918 (N_2918,N_1299,N_1207);
xnor U2919 (N_2919,N_2006,N_1942);
nand U2920 (N_2920,N_1827,N_1819);
nor U2921 (N_2921,N_1901,N_1430);
xnor U2922 (N_2922,N_1291,N_2066);
nor U2923 (N_2923,N_2278,N_1656);
xnor U2924 (N_2924,N_2000,N_1988);
and U2925 (N_2925,N_1448,N_1597);
or U2926 (N_2926,N_1904,N_1489);
xnor U2927 (N_2927,N_1677,N_1614);
or U2928 (N_2928,N_2251,N_1962);
or U2929 (N_2929,N_1826,N_2374);
xor U2930 (N_2930,N_2096,N_2185);
and U2931 (N_2931,N_1234,N_1336);
or U2932 (N_2932,N_2131,N_2110);
xnor U2933 (N_2933,N_1571,N_1469);
nor U2934 (N_2934,N_1973,N_1958);
nor U2935 (N_2935,N_1882,N_2087);
nand U2936 (N_2936,N_2199,N_1664);
or U2937 (N_2937,N_2344,N_1607);
and U2938 (N_2938,N_1865,N_1541);
and U2939 (N_2939,N_1908,N_1659);
nand U2940 (N_2940,N_1783,N_1995);
or U2941 (N_2941,N_1945,N_1927);
nor U2942 (N_2942,N_1798,N_1745);
nand U2943 (N_2943,N_1329,N_2215);
or U2944 (N_2944,N_1794,N_2361);
xor U2945 (N_2945,N_1249,N_1732);
or U2946 (N_2946,N_2356,N_1584);
nand U2947 (N_2947,N_2082,N_1703);
nand U2948 (N_2948,N_1516,N_2127);
nand U2949 (N_2949,N_2169,N_2319);
nand U2950 (N_2950,N_1900,N_1327);
nand U2951 (N_2951,N_2200,N_1831);
nand U2952 (N_2952,N_1310,N_1441);
nor U2953 (N_2953,N_2205,N_2336);
xnor U2954 (N_2954,N_1723,N_2054);
and U2955 (N_2955,N_2156,N_2168);
xor U2956 (N_2956,N_1804,N_2120);
or U2957 (N_2957,N_1279,N_1354);
xor U2958 (N_2958,N_1696,N_1402);
xor U2959 (N_2959,N_2394,N_1225);
and U2960 (N_2960,N_1431,N_1245);
or U2961 (N_2961,N_1940,N_1501);
or U2962 (N_2962,N_1711,N_2175);
and U2963 (N_2963,N_1638,N_1426);
nor U2964 (N_2964,N_1294,N_1726);
xnor U2965 (N_2965,N_1857,N_1849);
and U2966 (N_2966,N_1704,N_1215);
nand U2967 (N_2967,N_1308,N_1760);
nor U2968 (N_2968,N_1271,N_2085);
nand U2969 (N_2969,N_1306,N_2353);
nand U2970 (N_2970,N_1914,N_1530);
nor U2971 (N_2971,N_1586,N_2216);
xor U2972 (N_2972,N_1346,N_1915);
xnor U2973 (N_2973,N_1347,N_2182);
xnor U2974 (N_2974,N_2273,N_2357);
xor U2975 (N_2975,N_1629,N_1810);
nand U2976 (N_2976,N_1841,N_1737);
nand U2977 (N_2977,N_1708,N_1954);
xor U2978 (N_2978,N_1923,N_1767);
or U2979 (N_2979,N_1609,N_1906);
or U2980 (N_2980,N_2018,N_1661);
nand U2981 (N_2981,N_2270,N_1258);
and U2982 (N_2982,N_1282,N_1679);
nand U2983 (N_2983,N_1413,N_2214);
and U2984 (N_2984,N_1593,N_1262);
nand U2985 (N_2985,N_1360,N_1755);
xor U2986 (N_2986,N_1577,N_1337);
xnor U2987 (N_2987,N_2228,N_1682);
xnor U2988 (N_2988,N_1205,N_2108);
and U2989 (N_2989,N_1666,N_1596);
or U2990 (N_2990,N_2250,N_1297);
nand U2991 (N_2991,N_1564,N_1356);
nor U2992 (N_2992,N_1736,N_1202);
or U2993 (N_2993,N_1775,N_1640);
nand U2994 (N_2994,N_2399,N_2203);
nor U2995 (N_2995,N_1253,N_1563);
or U2996 (N_2996,N_1744,N_1524);
nand U2997 (N_2997,N_1537,N_1606);
xnor U2998 (N_2998,N_2297,N_1511);
or U2999 (N_2999,N_1871,N_2331);
or U3000 (N_3000,N_2143,N_2384);
and U3001 (N_3001,N_1744,N_1251);
or U3002 (N_3002,N_1670,N_1926);
or U3003 (N_3003,N_1270,N_1839);
and U3004 (N_3004,N_1516,N_1490);
and U3005 (N_3005,N_2063,N_2072);
nor U3006 (N_3006,N_1800,N_2306);
nand U3007 (N_3007,N_2175,N_2229);
xnor U3008 (N_3008,N_2178,N_1952);
nor U3009 (N_3009,N_2158,N_2112);
nand U3010 (N_3010,N_1249,N_2206);
nor U3011 (N_3011,N_2016,N_2374);
nor U3012 (N_3012,N_1493,N_1833);
or U3013 (N_3013,N_1413,N_1672);
nand U3014 (N_3014,N_1241,N_2362);
xnor U3015 (N_3015,N_1429,N_1605);
or U3016 (N_3016,N_2086,N_1346);
and U3017 (N_3017,N_1298,N_1809);
nand U3018 (N_3018,N_1747,N_1560);
nand U3019 (N_3019,N_2210,N_2046);
xor U3020 (N_3020,N_2367,N_2285);
nand U3021 (N_3021,N_2122,N_1820);
nand U3022 (N_3022,N_1921,N_1431);
nand U3023 (N_3023,N_1903,N_1454);
xnor U3024 (N_3024,N_2189,N_2216);
xor U3025 (N_3025,N_1527,N_2114);
xnor U3026 (N_3026,N_1342,N_2128);
nand U3027 (N_3027,N_1568,N_1406);
or U3028 (N_3028,N_1611,N_2377);
nand U3029 (N_3029,N_2331,N_1422);
xnor U3030 (N_3030,N_1525,N_1289);
or U3031 (N_3031,N_1256,N_2176);
or U3032 (N_3032,N_1349,N_2142);
or U3033 (N_3033,N_1462,N_2080);
nand U3034 (N_3034,N_1346,N_1966);
and U3035 (N_3035,N_1441,N_2091);
xor U3036 (N_3036,N_1223,N_2042);
or U3037 (N_3037,N_1913,N_2265);
nor U3038 (N_3038,N_1384,N_1214);
nand U3039 (N_3039,N_2157,N_1668);
nor U3040 (N_3040,N_2001,N_1889);
nor U3041 (N_3041,N_1780,N_1442);
xnor U3042 (N_3042,N_1599,N_1881);
nand U3043 (N_3043,N_1788,N_1827);
or U3044 (N_3044,N_1436,N_1462);
and U3045 (N_3045,N_2323,N_2249);
nor U3046 (N_3046,N_1385,N_2284);
or U3047 (N_3047,N_1380,N_1389);
or U3048 (N_3048,N_1620,N_2219);
or U3049 (N_3049,N_2059,N_2349);
xor U3050 (N_3050,N_1334,N_1712);
and U3051 (N_3051,N_1936,N_2110);
and U3052 (N_3052,N_1232,N_2038);
or U3053 (N_3053,N_1501,N_2360);
or U3054 (N_3054,N_2214,N_1960);
or U3055 (N_3055,N_2050,N_2378);
nand U3056 (N_3056,N_2145,N_2076);
xnor U3057 (N_3057,N_1712,N_1382);
nand U3058 (N_3058,N_2018,N_1936);
xor U3059 (N_3059,N_2375,N_1496);
nor U3060 (N_3060,N_2115,N_1443);
and U3061 (N_3061,N_1846,N_1373);
or U3062 (N_3062,N_2119,N_1290);
xor U3063 (N_3063,N_1571,N_1735);
or U3064 (N_3064,N_2101,N_1619);
nand U3065 (N_3065,N_2026,N_1660);
or U3066 (N_3066,N_1573,N_1786);
nand U3067 (N_3067,N_1863,N_2339);
nor U3068 (N_3068,N_1669,N_2316);
nor U3069 (N_3069,N_2116,N_2109);
and U3070 (N_3070,N_2180,N_1613);
nand U3071 (N_3071,N_1325,N_1738);
and U3072 (N_3072,N_1479,N_1275);
nor U3073 (N_3073,N_1441,N_1949);
nand U3074 (N_3074,N_1867,N_1485);
and U3075 (N_3075,N_2187,N_1836);
xor U3076 (N_3076,N_1874,N_1483);
xor U3077 (N_3077,N_1810,N_1391);
and U3078 (N_3078,N_1405,N_1561);
and U3079 (N_3079,N_1248,N_2323);
or U3080 (N_3080,N_2228,N_1363);
and U3081 (N_3081,N_1632,N_1255);
nor U3082 (N_3082,N_2017,N_2148);
xnor U3083 (N_3083,N_1538,N_1327);
nor U3084 (N_3084,N_2350,N_2191);
and U3085 (N_3085,N_1514,N_1548);
or U3086 (N_3086,N_1878,N_1373);
nor U3087 (N_3087,N_1842,N_2291);
or U3088 (N_3088,N_2381,N_2073);
and U3089 (N_3089,N_1217,N_1496);
and U3090 (N_3090,N_2136,N_1495);
nand U3091 (N_3091,N_1266,N_2149);
nor U3092 (N_3092,N_1461,N_1238);
nand U3093 (N_3093,N_1319,N_2354);
and U3094 (N_3094,N_1718,N_1773);
or U3095 (N_3095,N_2269,N_1883);
nand U3096 (N_3096,N_2330,N_2155);
xnor U3097 (N_3097,N_2339,N_2320);
nand U3098 (N_3098,N_2130,N_1486);
xor U3099 (N_3099,N_1448,N_1523);
nor U3100 (N_3100,N_1217,N_2168);
or U3101 (N_3101,N_1959,N_1681);
and U3102 (N_3102,N_2106,N_1213);
or U3103 (N_3103,N_1880,N_1218);
xor U3104 (N_3104,N_2100,N_1915);
and U3105 (N_3105,N_1808,N_1771);
nand U3106 (N_3106,N_2027,N_1445);
nor U3107 (N_3107,N_2163,N_1762);
and U3108 (N_3108,N_1769,N_1577);
nand U3109 (N_3109,N_1842,N_1268);
nand U3110 (N_3110,N_1220,N_1636);
xnor U3111 (N_3111,N_1392,N_1722);
xor U3112 (N_3112,N_1722,N_1714);
and U3113 (N_3113,N_1945,N_2130);
nand U3114 (N_3114,N_1207,N_2083);
and U3115 (N_3115,N_2252,N_1931);
nor U3116 (N_3116,N_2194,N_1795);
xnor U3117 (N_3117,N_1546,N_2301);
nor U3118 (N_3118,N_1768,N_1900);
nand U3119 (N_3119,N_2293,N_1479);
xor U3120 (N_3120,N_2383,N_1733);
nor U3121 (N_3121,N_1756,N_2273);
xnor U3122 (N_3122,N_1868,N_2114);
nor U3123 (N_3123,N_2394,N_2183);
xor U3124 (N_3124,N_1339,N_2048);
xor U3125 (N_3125,N_2391,N_1435);
and U3126 (N_3126,N_1434,N_2021);
or U3127 (N_3127,N_1237,N_2315);
nand U3128 (N_3128,N_1698,N_2284);
and U3129 (N_3129,N_1902,N_1924);
nor U3130 (N_3130,N_1502,N_2192);
nand U3131 (N_3131,N_1742,N_2119);
and U3132 (N_3132,N_2222,N_2190);
nor U3133 (N_3133,N_1934,N_1569);
nand U3134 (N_3134,N_1507,N_2076);
or U3135 (N_3135,N_1691,N_1999);
or U3136 (N_3136,N_1632,N_1956);
or U3137 (N_3137,N_2368,N_2009);
and U3138 (N_3138,N_1382,N_1983);
and U3139 (N_3139,N_1942,N_2369);
xor U3140 (N_3140,N_1403,N_2271);
or U3141 (N_3141,N_1737,N_2393);
xnor U3142 (N_3142,N_1410,N_2062);
or U3143 (N_3143,N_1219,N_2149);
or U3144 (N_3144,N_1970,N_1499);
nand U3145 (N_3145,N_1411,N_2386);
nand U3146 (N_3146,N_1881,N_1552);
xnor U3147 (N_3147,N_1786,N_1693);
nand U3148 (N_3148,N_2285,N_1596);
nor U3149 (N_3149,N_1214,N_2019);
xnor U3150 (N_3150,N_2049,N_2248);
xnor U3151 (N_3151,N_2299,N_1946);
or U3152 (N_3152,N_1452,N_1213);
nor U3153 (N_3153,N_2311,N_1743);
xnor U3154 (N_3154,N_1914,N_1837);
and U3155 (N_3155,N_1843,N_1278);
nor U3156 (N_3156,N_1526,N_1250);
and U3157 (N_3157,N_2159,N_1355);
nor U3158 (N_3158,N_1885,N_2095);
or U3159 (N_3159,N_1441,N_1242);
nand U3160 (N_3160,N_2384,N_1406);
and U3161 (N_3161,N_2368,N_2381);
and U3162 (N_3162,N_1407,N_1885);
or U3163 (N_3163,N_2159,N_1461);
or U3164 (N_3164,N_1803,N_2218);
or U3165 (N_3165,N_1511,N_1677);
xor U3166 (N_3166,N_1512,N_1818);
and U3167 (N_3167,N_1893,N_2397);
or U3168 (N_3168,N_2108,N_2144);
nor U3169 (N_3169,N_1244,N_2301);
nor U3170 (N_3170,N_2101,N_2176);
and U3171 (N_3171,N_1924,N_1587);
or U3172 (N_3172,N_2015,N_1465);
or U3173 (N_3173,N_1770,N_1693);
nor U3174 (N_3174,N_2118,N_1622);
or U3175 (N_3175,N_1774,N_1819);
xnor U3176 (N_3176,N_1377,N_2208);
and U3177 (N_3177,N_2162,N_1378);
and U3178 (N_3178,N_1631,N_2095);
nor U3179 (N_3179,N_1651,N_1213);
xor U3180 (N_3180,N_2197,N_1710);
nor U3181 (N_3181,N_1513,N_1365);
nand U3182 (N_3182,N_1593,N_1417);
nor U3183 (N_3183,N_2130,N_2016);
xnor U3184 (N_3184,N_1589,N_1348);
or U3185 (N_3185,N_2093,N_1941);
and U3186 (N_3186,N_1318,N_1249);
or U3187 (N_3187,N_1654,N_1794);
xor U3188 (N_3188,N_2209,N_2070);
nor U3189 (N_3189,N_1596,N_2308);
and U3190 (N_3190,N_2015,N_1615);
and U3191 (N_3191,N_1425,N_1661);
nand U3192 (N_3192,N_2221,N_2193);
nand U3193 (N_3193,N_1223,N_2097);
nand U3194 (N_3194,N_2172,N_1950);
or U3195 (N_3195,N_2223,N_1381);
nand U3196 (N_3196,N_1421,N_1562);
or U3197 (N_3197,N_2127,N_1443);
nand U3198 (N_3198,N_1220,N_1310);
and U3199 (N_3199,N_1608,N_1255);
and U3200 (N_3200,N_1885,N_1463);
xnor U3201 (N_3201,N_1976,N_1819);
nand U3202 (N_3202,N_2123,N_1442);
and U3203 (N_3203,N_2076,N_1266);
xnor U3204 (N_3204,N_2312,N_1837);
and U3205 (N_3205,N_1683,N_1408);
and U3206 (N_3206,N_1666,N_2294);
nor U3207 (N_3207,N_1341,N_1642);
nand U3208 (N_3208,N_1888,N_1972);
nor U3209 (N_3209,N_2351,N_1845);
or U3210 (N_3210,N_1304,N_1672);
xor U3211 (N_3211,N_1666,N_2145);
xnor U3212 (N_3212,N_1614,N_2147);
xnor U3213 (N_3213,N_1597,N_2308);
xnor U3214 (N_3214,N_1421,N_2279);
nand U3215 (N_3215,N_1212,N_1671);
or U3216 (N_3216,N_2141,N_2250);
or U3217 (N_3217,N_2204,N_1772);
nor U3218 (N_3218,N_2126,N_2268);
or U3219 (N_3219,N_2199,N_1314);
nand U3220 (N_3220,N_1696,N_1445);
nor U3221 (N_3221,N_2293,N_1679);
nor U3222 (N_3222,N_2282,N_2342);
or U3223 (N_3223,N_2046,N_1792);
and U3224 (N_3224,N_2368,N_1455);
and U3225 (N_3225,N_1294,N_2059);
and U3226 (N_3226,N_1626,N_1478);
nand U3227 (N_3227,N_1664,N_1997);
nand U3228 (N_3228,N_2004,N_1281);
or U3229 (N_3229,N_1392,N_1849);
xor U3230 (N_3230,N_1211,N_1527);
or U3231 (N_3231,N_2090,N_2053);
or U3232 (N_3232,N_2237,N_1903);
xor U3233 (N_3233,N_2360,N_1857);
and U3234 (N_3234,N_1395,N_1482);
and U3235 (N_3235,N_1584,N_1340);
nand U3236 (N_3236,N_1667,N_1373);
nand U3237 (N_3237,N_2334,N_1819);
or U3238 (N_3238,N_2058,N_1954);
or U3239 (N_3239,N_1224,N_1411);
xor U3240 (N_3240,N_1566,N_2223);
nor U3241 (N_3241,N_1385,N_1550);
xnor U3242 (N_3242,N_1997,N_1418);
xor U3243 (N_3243,N_1498,N_2029);
nor U3244 (N_3244,N_1703,N_1866);
or U3245 (N_3245,N_1340,N_1987);
or U3246 (N_3246,N_1375,N_1233);
nand U3247 (N_3247,N_2067,N_1966);
and U3248 (N_3248,N_2308,N_1958);
nand U3249 (N_3249,N_1866,N_2363);
nor U3250 (N_3250,N_1330,N_1965);
or U3251 (N_3251,N_2191,N_1273);
xnor U3252 (N_3252,N_1512,N_1610);
xor U3253 (N_3253,N_1751,N_1415);
xnor U3254 (N_3254,N_1330,N_2122);
and U3255 (N_3255,N_1517,N_2210);
nor U3256 (N_3256,N_2164,N_1356);
nand U3257 (N_3257,N_2361,N_2299);
xor U3258 (N_3258,N_1418,N_1572);
nor U3259 (N_3259,N_2099,N_1434);
nor U3260 (N_3260,N_1204,N_1245);
nand U3261 (N_3261,N_1704,N_1668);
or U3262 (N_3262,N_1563,N_1652);
nand U3263 (N_3263,N_1982,N_2297);
nand U3264 (N_3264,N_1925,N_1377);
nand U3265 (N_3265,N_1985,N_1248);
or U3266 (N_3266,N_1367,N_1432);
and U3267 (N_3267,N_1450,N_2295);
xor U3268 (N_3268,N_1697,N_1391);
nand U3269 (N_3269,N_1739,N_2069);
or U3270 (N_3270,N_2094,N_1959);
or U3271 (N_3271,N_2215,N_2077);
xor U3272 (N_3272,N_1831,N_2311);
nor U3273 (N_3273,N_2356,N_1285);
or U3274 (N_3274,N_1975,N_1513);
nand U3275 (N_3275,N_1345,N_2004);
and U3276 (N_3276,N_2012,N_2077);
nand U3277 (N_3277,N_2336,N_1385);
nand U3278 (N_3278,N_1722,N_2270);
xnor U3279 (N_3279,N_2181,N_2388);
and U3280 (N_3280,N_1677,N_1691);
nand U3281 (N_3281,N_1896,N_1576);
nand U3282 (N_3282,N_1469,N_1597);
or U3283 (N_3283,N_1979,N_1666);
nor U3284 (N_3284,N_2122,N_2244);
nand U3285 (N_3285,N_1960,N_2093);
nand U3286 (N_3286,N_1472,N_2106);
and U3287 (N_3287,N_1895,N_1784);
or U3288 (N_3288,N_1405,N_1685);
xnor U3289 (N_3289,N_1519,N_1690);
nand U3290 (N_3290,N_1542,N_2074);
nor U3291 (N_3291,N_2373,N_1692);
nor U3292 (N_3292,N_2054,N_2070);
or U3293 (N_3293,N_1544,N_1963);
nand U3294 (N_3294,N_1995,N_2204);
xor U3295 (N_3295,N_1741,N_1887);
and U3296 (N_3296,N_2093,N_1937);
nand U3297 (N_3297,N_1930,N_1239);
and U3298 (N_3298,N_1494,N_1751);
nand U3299 (N_3299,N_1646,N_2359);
or U3300 (N_3300,N_1664,N_1632);
nand U3301 (N_3301,N_2258,N_1662);
and U3302 (N_3302,N_1372,N_1479);
xor U3303 (N_3303,N_1441,N_1231);
nand U3304 (N_3304,N_2235,N_1849);
and U3305 (N_3305,N_2167,N_1881);
nand U3306 (N_3306,N_1776,N_1557);
xor U3307 (N_3307,N_1702,N_1321);
nand U3308 (N_3308,N_2242,N_2148);
and U3309 (N_3309,N_1313,N_2151);
and U3310 (N_3310,N_2128,N_1771);
and U3311 (N_3311,N_2199,N_1590);
or U3312 (N_3312,N_1772,N_1536);
and U3313 (N_3313,N_1961,N_1627);
nand U3314 (N_3314,N_1594,N_1253);
nor U3315 (N_3315,N_1640,N_2200);
nand U3316 (N_3316,N_2373,N_2054);
nor U3317 (N_3317,N_2191,N_1956);
or U3318 (N_3318,N_1462,N_1781);
nor U3319 (N_3319,N_1855,N_1212);
xnor U3320 (N_3320,N_1314,N_2008);
xor U3321 (N_3321,N_1814,N_2034);
nor U3322 (N_3322,N_1595,N_1824);
or U3323 (N_3323,N_1746,N_1784);
nand U3324 (N_3324,N_1385,N_1663);
or U3325 (N_3325,N_1765,N_2141);
nor U3326 (N_3326,N_1537,N_1500);
nor U3327 (N_3327,N_1939,N_2020);
or U3328 (N_3328,N_2306,N_2292);
or U3329 (N_3329,N_1942,N_1450);
xor U3330 (N_3330,N_1937,N_1385);
nor U3331 (N_3331,N_1733,N_2192);
or U3332 (N_3332,N_1864,N_2395);
nor U3333 (N_3333,N_1619,N_1577);
or U3334 (N_3334,N_1314,N_1844);
xnor U3335 (N_3335,N_1930,N_2060);
xor U3336 (N_3336,N_2269,N_1384);
xor U3337 (N_3337,N_1269,N_1234);
nand U3338 (N_3338,N_1619,N_2063);
nand U3339 (N_3339,N_1377,N_2091);
and U3340 (N_3340,N_2012,N_1665);
nor U3341 (N_3341,N_2300,N_2220);
nand U3342 (N_3342,N_1479,N_2127);
nor U3343 (N_3343,N_1231,N_1325);
or U3344 (N_3344,N_1663,N_1972);
xor U3345 (N_3345,N_2263,N_1268);
xor U3346 (N_3346,N_1612,N_1570);
nand U3347 (N_3347,N_1737,N_1622);
xnor U3348 (N_3348,N_1890,N_2057);
nor U3349 (N_3349,N_1890,N_1321);
or U3350 (N_3350,N_1472,N_2232);
nor U3351 (N_3351,N_1304,N_1455);
and U3352 (N_3352,N_1677,N_1733);
nand U3353 (N_3353,N_2371,N_1362);
nand U3354 (N_3354,N_2297,N_2132);
and U3355 (N_3355,N_2141,N_2007);
and U3356 (N_3356,N_1467,N_1651);
and U3357 (N_3357,N_2391,N_1747);
nor U3358 (N_3358,N_2195,N_2211);
nand U3359 (N_3359,N_1303,N_1239);
or U3360 (N_3360,N_1703,N_1588);
xnor U3361 (N_3361,N_2148,N_1735);
xnor U3362 (N_3362,N_1267,N_2211);
nand U3363 (N_3363,N_1882,N_1623);
xor U3364 (N_3364,N_1971,N_1706);
nand U3365 (N_3365,N_2202,N_1544);
and U3366 (N_3366,N_2263,N_2179);
xnor U3367 (N_3367,N_1628,N_1622);
xnor U3368 (N_3368,N_1480,N_1501);
or U3369 (N_3369,N_2144,N_1755);
xor U3370 (N_3370,N_1790,N_1955);
and U3371 (N_3371,N_1681,N_2002);
and U3372 (N_3372,N_2288,N_2018);
nor U3373 (N_3373,N_1301,N_1598);
nor U3374 (N_3374,N_1645,N_1575);
nand U3375 (N_3375,N_2254,N_1685);
or U3376 (N_3376,N_2021,N_1931);
nor U3377 (N_3377,N_2104,N_1374);
nor U3378 (N_3378,N_1205,N_1369);
nand U3379 (N_3379,N_1537,N_1743);
and U3380 (N_3380,N_1429,N_2161);
and U3381 (N_3381,N_1643,N_1820);
nor U3382 (N_3382,N_1628,N_1293);
xor U3383 (N_3383,N_1887,N_2106);
and U3384 (N_3384,N_1492,N_1272);
nor U3385 (N_3385,N_1308,N_1505);
nor U3386 (N_3386,N_1565,N_2280);
xor U3387 (N_3387,N_1858,N_1461);
and U3388 (N_3388,N_1565,N_1719);
xnor U3389 (N_3389,N_1885,N_1975);
and U3390 (N_3390,N_2124,N_2301);
xor U3391 (N_3391,N_1639,N_2225);
nand U3392 (N_3392,N_1643,N_1538);
xor U3393 (N_3393,N_1719,N_2161);
nand U3394 (N_3394,N_1340,N_1927);
nor U3395 (N_3395,N_1711,N_2211);
nor U3396 (N_3396,N_1939,N_1792);
nand U3397 (N_3397,N_1606,N_1303);
nand U3398 (N_3398,N_1804,N_1230);
nor U3399 (N_3399,N_1522,N_1687);
and U3400 (N_3400,N_1586,N_1543);
nand U3401 (N_3401,N_1579,N_2112);
xnor U3402 (N_3402,N_2029,N_1793);
xnor U3403 (N_3403,N_1307,N_2239);
and U3404 (N_3404,N_2075,N_1449);
or U3405 (N_3405,N_2347,N_2344);
and U3406 (N_3406,N_2086,N_1510);
xor U3407 (N_3407,N_1253,N_1522);
and U3408 (N_3408,N_1976,N_1746);
or U3409 (N_3409,N_1779,N_2210);
nor U3410 (N_3410,N_1518,N_1431);
and U3411 (N_3411,N_1793,N_1974);
and U3412 (N_3412,N_1426,N_1444);
xnor U3413 (N_3413,N_1322,N_1638);
and U3414 (N_3414,N_2333,N_1854);
nor U3415 (N_3415,N_2069,N_2003);
nand U3416 (N_3416,N_1453,N_1252);
nor U3417 (N_3417,N_2307,N_1214);
and U3418 (N_3418,N_2099,N_2124);
and U3419 (N_3419,N_1313,N_1734);
nor U3420 (N_3420,N_2160,N_1839);
or U3421 (N_3421,N_1734,N_2310);
nand U3422 (N_3422,N_2250,N_2303);
nand U3423 (N_3423,N_1338,N_1318);
and U3424 (N_3424,N_1791,N_2260);
and U3425 (N_3425,N_1761,N_1457);
xnor U3426 (N_3426,N_2155,N_2071);
and U3427 (N_3427,N_1302,N_1813);
nor U3428 (N_3428,N_2156,N_1751);
and U3429 (N_3429,N_2100,N_2240);
and U3430 (N_3430,N_1671,N_1738);
nor U3431 (N_3431,N_1902,N_1257);
and U3432 (N_3432,N_1379,N_1465);
xor U3433 (N_3433,N_2160,N_1591);
nand U3434 (N_3434,N_2337,N_1421);
and U3435 (N_3435,N_2121,N_1710);
or U3436 (N_3436,N_1228,N_2049);
and U3437 (N_3437,N_2369,N_1617);
nand U3438 (N_3438,N_1793,N_2015);
nor U3439 (N_3439,N_2146,N_1494);
or U3440 (N_3440,N_2319,N_1505);
nor U3441 (N_3441,N_1970,N_1927);
or U3442 (N_3442,N_2256,N_2150);
and U3443 (N_3443,N_2160,N_1475);
nor U3444 (N_3444,N_2221,N_1452);
and U3445 (N_3445,N_2345,N_1922);
xor U3446 (N_3446,N_1691,N_1351);
and U3447 (N_3447,N_1329,N_2088);
nor U3448 (N_3448,N_1328,N_2076);
nor U3449 (N_3449,N_1454,N_1704);
and U3450 (N_3450,N_1968,N_1844);
or U3451 (N_3451,N_1784,N_1850);
xnor U3452 (N_3452,N_1937,N_1323);
and U3453 (N_3453,N_2325,N_2278);
and U3454 (N_3454,N_1478,N_1708);
nand U3455 (N_3455,N_1462,N_1549);
xnor U3456 (N_3456,N_1991,N_2213);
or U3457 (N_3457,N_1208,N_1497);
xnor U3458 (N_3458,N_2136,N_2346);
and U3459 (N_3459,N_1907,N_1649);
nor U3460 (N_3460,N_2320,N_1409);
xnor U3461 (N_3461,N_1473,N_1743);
or U3462 (N_3462,N_2313,N_1335);
nand U3463 (N_3463,N_1751,N_2088);
nor U3464 (N_3464,N_1955,N_1891);
xnor U3465 (N_3465,N_2087,N_1957);
and U3466 (N_3466,N_1373,N_1799);
xor U3467 (N_3467,N_2171,N_1701);
and U3468 (N_3468,N_1816,N_1438);
and U3469 (N_3469,N_2220,N_2376);
xor U3470 (N_3470,N_1460,N_1275);
nand U3471 (N_3471,N_1894,N_1204);
xnor U3472 (N_3472,N_1361,N_1276);
or U3473 (N_3473,N_1334,N_1711);
and U3474 (N_3474,N_2180,N_1360);
xor U3475 (N_3475,N_2199,N_2133);
nand U3476 (N_3476,N_1933,N_1870);
or U3477 (N_3477,N_2096,N_2239);
xnor U3478 (N_3478,N_1288,N_2263);
nor U3479 (N_3479,N_1895,N_1465);
nand U3480 (N_3480,N_1255,N_2368);
and U3481 (N_3481,N_1938,N_2174);
and U3482 (N_3482,N_1765,N_2392);
nand U3483 (N_3483,N_2390,N_1685);
nand U3484 (N_3484,N_1735,N_1708);
xor U3485 (N_3485,N_1649,N_1877);
or U3486 (N_3486,N_1674,N_1560);
and U3487 (N_3487,N_1405,N_1377);
xnor U3488 (N_3488,N_1426,N_2313);
xnor U3489 (N_3489,N_1838,N_1404);
nor U3490 (N_3490,N_1521,N_1216);
nand U3491 (N_3491,N_1938,N_2290);
and U3492 (N_3492,N_1518,N_2155);
xnor U3493 (N_3493,N_1740,N_1761);
xnor U3494 (N_3494,N_1294,N_1818);
xnor U3495 (N_3495,N_2010,N_2086);
xnor U3496 (N_3496,N_2214,N_2069);
nor U3497 (N_3497,N_2364,N_1370);
and U3498 (N_3498,N_1870,N_2085);
xnor U3499 (N_3499,N_1704,N_1234);
or U3500 (N_3500,N_2171,N_1505);
or U3501 (N_3501,N_2073,N_2189);
and U3502 (N_3502,N_1996,N_1816);
nand U3503 (N_3503,N_1904,N_2316);
and U3504 (N_3504,N_1289,N_1538);
or U3505 (N_3505,N_1431,N_1633);
nand U3506 (N_3506,N_1524,N_2317);
or U3507 (N_3507,N_1411,N_2226);
xnor U3508 (N_3508,N_1544,N_1709);
nor U3509 (N_3509,N_2385,N_2177);
nor U3510 (N_3510,N_1297,N_1484);
nand U3511 (N_3511,N_1967,N_1428);
xor U3512 (N_3512,N_2132,N_1949);
xnor U3513 (N_3513,N_1340,N_2322);
and U3514 (N_3514,N_1878,N_1255);
or U3515 (N_3515,N_1274,N_1224);
nor U3516 (N_3516,N_1382,N_1204);
xnor U3517 (N_3517,N_1532,N_2082);
nand U3518 (N_3518,N_2021,N_2103);
and U3519 (N_3519,N_2270,N_1851);
nor U3520 (N_3520,N_1970,N_2208);
nand U3521 (N_3521,N_1255,N_1483);
xnor U3522 (N_3522,N_2261,N_2378);
nand U3523 (N_3523,N_1883,N_1905);
nand U3524 (N_3524,N_2352,N_2239);
nor U3525 (N_3525,N_1718,N_2348);
xor U3526 (N_3526,N_2130,N_1677);
nand U3527 (N_3527,N_1541,N_2390);
and U3528 (N_3528,N_1338,N_1665);
nand U3529 (N_3529,N_1330,N_1982);
nand U3530 (N_3530,N_2365,N_1918);
and U3531 (N_3531,N_1294,N_1637);
nand U3532 (N_3532,N_1836,N_1495);
nand U3533 (N_3533,N_1433,N_1573);
nor U3534 (N_3534,N_2051,N_1461);
xnor U3535 (N_3535,N_1596,N_2186);
nor U3536 (N_3536,N_1593,N_1450);
and U3537 (N_3537,N_1880,N_2293);
xor U3538 (N_3538,N_2342,N_1605);
nand U3539 (N_3539,N_2255,N_1972);
nor U3540 (N_3540,N_2180,N_1660);
nand U3541 (N_3541,N_1679,N_1207);
xor U3542 (N_3542,N_2249,N_1494);
xnor U3543 (N_3543,N_1201,N_1925);
nand U3544 (N_3544,N_1972,N_1960);
and U3545 (N_3545,N_1460,N_1659);
or U3546 (N_3546,N_1606,N_1615);
nand U3547 (N_3547,N_1232,N_2386);
and U3548 (N_3548,N_1615,N_1452);
and U3549 (N_3549,N_1537,N_1583);
nor U3550 (N_3550,N_1556,N_2384);
nor U3551 (N_3551,N_2051,N_2119);
xor U3552 (N_3552,N_1981,N_1219);
or U3553 (N_3553,N_2060,N_2208);
nor U3554 (N_3554,N_1528,N_1266);
xor U3555 (N_3555,N_2283,N_1430);
nand U3556 (N_3556,N_2336,N_2150);
nor U3557 (N_3557,N_1816,N_1264);
nand U3558 (N_3558,N_1473,N_1590);
nor U3559 (N_3559,N_2153,N_1977);
and U3560 (N_3560,N_1300,N_1266);
or U3561 (N_3561,N_1360,N_2100);
or U3562 (N_3562,N_2214,N_2210);
or U3563 (N_3563,N_1466,N_2094);
nor U3564 (N_3564,N_1976,N_2135);
nor U3565 (N_3565,N_1650,N_1956);
and U3566 (N_3566,N_1709,N_1581);
nor U3567 (N_3567,N_2080,N_2259);
and U3568 (N_3568,N_1985,N_2073);
nor U3569 (N_3569,N_1551,N_2179);
xor U3570 (N_3570,N_1616,N_1614);
nand U3571 (N_3571,N_1294,N_1433);
nor U3572 (N_3572,N_1424,N_1557);
nand U3573 (N_3573,N_1615,N_1614);
and U3574 (N_3574,N_1738,N_1247);
or U3575 (N_3575,N_2353,N_1751);
and U3576 (N_3576,N_1489,N_2267);
or U3577 (N_3577,N_1738,N_1910);
xnor U3578 (N_3578,N_1593,N_1788);
or U3579 (N_3579,N_1817,N_1987);
and U3580 (N_3580,N_1323,N_2323);
and U3581 (N_3581,N_1537,N_1227);
and U3582 (N_3582,N_2308,N_1558);
nor U3583 (N_3583,N_2004,N_2332);
or U3584 (N_3584,N_1826,N_2380);
and U3585 (N_3585,N_1971,N_1513);
nand U3586 (N_3586,N_1989,N_2274);
nand U3587 (N_3587,N_2068,N_1762);
and U3588 (N_3588,N_1750,N_1566);
nor U3589 (N_3589,N_2187,N_1920);
nand U3590 (N_3590,N_2341,N_1714);
xnor U3591 (N_3591,N_2357,N_1378);
and U3592 (N_3592,N_1472,N_2350);
or U3593 (N_3593,N_1834,N_1879);
or U3594 (N_3594,N_1431,N_1444);
nand U3595 (N_3595,N_1928,N_1330);
nor U3596 (N_3596,N_1201,N_1663);
nand U3597 (N_3597,N_2219,N_1547);
and U3598 (N_3598,N_1305,N_1729);
or U3599 (N_3599,N_1283,N_2196);
and U3600 (N_3600,N_2741,N_2718);
and U3601 (N_3601,N_3528,N_3390);
nor U3602 (N_3602,N_2753,N_2926);
xnor U3603 (N_3603,N_2964,N_3341);
nand U3604 (N_3604,N_3159,N_3027);
nor U3605 (N_3605,N_3401,N_2966);
nor U3606 (N_3606,N_2884,N_3108);
nor U3607 (N_3607,N_2549,N_3359);
or U3608 (N_3608,N_2871,N_3102);
xnor U3609 (N_3609,N_2878,N_3251);
or U3610 (N_3610,N_2849,N_3060);
nand U3611 (N_3611,N_3020,N_3112);
or U3612 (N_3612,N_3039,N_2591);
and U3613 (N_3613,N_2516,N_2876);
xor U3614 (N_3614,N_3469,N_2571);
xnor U3615 (N_3615,N_2800,N_3491);
nand U3616 (N_3616,N_2761,N_3490);
xor U3617 (N_3617,N_2856,N_3510);
nand U3618 (N_3618,N_3180,N_2424);
nand U3619 (N_3619,N_2507,N_2640);
or U3620 (N_3620,N_2732,N_3275);
or U3621 (N_3621,N_2608,N_3193);
nor U3622 (N_3622,N_3221,N_3555);
nor U3623 (N_3623,N_2406,N_3142);
or U3624 (N_3624,N_3363,N_3071);
or U3625 (N_3625,N_3082,N_3339);
and U3626 (N_3626,N_3048,N_3452);
nor U3627 (N_3627,N_2739,N_2680);
xnor U3628 (N_3628,N_2863,N_3319);
nor U3629 (N_3629,N_2911,N_2728);
or U3630 (N_3630,N_2799,N_3459);
or U3631 (N_3631,N_2559,N_2487);
nor U3632 (N_3632,N_2414,N_3414);
nor U3633 (N_3633,N_3132,N_3432);
or U3634 (N_3634,N_2961,N_3547);
nand U3635 (N_3635,N_2981,N_2552);
nor U3636 (N_3636,N_2913,N_2916);
and U3637 (N_3637,N_2595,N_3161);
nor U3638 (N_3638,N_2442,N_3206);
nand U3639 (N_3639,N_3382,N_3046);
or U3640 (N_3640,N_2982,N_3399);
or U3641 (N_3641,N_2457,N_3535);
or U3642 (N_3642,N_2942,N_2635);
nand U3643 (N_3643,N_2600,N_2580);
nor U3644 (N_3644,N_2658,N_3470);
nor U3645 (N_3645,N_2449,N_3171);
nand U3646 (N_3646,N_2893,N_3538);
xor U3647 (N_3647,N_2874,N_2717);
nand U3648 (N_3648,N_2996,N_3294);
xnor U3649 (N_3649,N_2473,N_3500);
nand U3650 (N_3650,N_3595,N_2777);
or U3651 (N_3651,N_3434,N_2400);
xor U3652 (N_3652,N_2810,N_3322);
or U3653 (N_3653,N_2491,N_3301);
and U3654 (N_3654,N_2788,N_3453);
and U3655 (N_3655,N_2675,N_3278);
nand U3656 (N_3656,N_3077,N_2703);
and U3657 (N_3657,N_2484,N_2809);
and U3658 (N_3658,N_3335,N_2494);
nand U3659 (N_3659,N_3557,N_3466);
and U3660 (N_3660,N_3332,N_3114);
nand U3661 (N_3661,N_3398,N_3389);
nor U3662 (N_3662,N_3391,N_3174);
xnor U3663 (N_3663,N_3521,N_3482);
nand U3664 (N_3664,N_3073,N_2953);
nand U3665 (N_3665,N_2420,N_2505);
or U3666 (N_3666,N_2922,N_2789);
nor U3667 (N_3667,N_3563,N_2662);
or U3668 (N_3668,N_2468,N_2567);
xnor U3669 (N_3669,N_3146,N_2485);
or U3670 (N_3670,N_3006,N_2845);
nor U3671 (N_3671,N_3329,N_2509);
or U3672 (N_3672,N_2985,N_2721);
nor U3673 (N_3673,N_3219,N_2903);
xor U3674 (N_3674,N_3511,N_2607);
and U3675 (N_3675,N_2746,N_3277);
nor U3676 (N_3676,N_2550,N_3014);
or U3677 (N_3677,N_2652,N_3517);
nand U3678 (N_3678,N_3334,N_2632);
xnor U3679 (N_3679,N_2792,N_2476);
nand U3680 (N_3680,N_2489,N_2664);
or U3681 (N_3681,N_3136,N_3549);
or U3682 (N_3682,N_3156,N_2415);
or U3683 (N_3683,N_3472,N_3493);
and U3684 (N_3684,N_2514,N_3587);
nor U3685 (N_3685,N_3581,N_2740);
nand U3686 (N_3686,N_2645,N_3150);
and U3687 (N_3687,N_3366,N_2599);
and U3688 (N_3688,N_3593,N_3525);
nor U3689 (N_3689,N_3323,N_3342);
nor U3690 (N_3690,N_2905,N_2417);
nand U3691 (N_3691,N_2997,N_3138);
nor U3692 (N_3692,N_3530,N_2637);
and U3693 (N_3693,N_3049,N_3099);
nor U3694 (N_3694,N_3464,N_2619);
nor U3695 (N_3695,N_2822,N_3565);
nor U3696 (N_3696,N_3461,N_3418);
xor U3697 (N_3697,N_2682,N_3520);
or U3698 (N_3698,N_3599,N_3368);
nor U3699 (N_3699,N_3243,N_3412);
nand U3700 (N_3700,N_3188,N_3578);
or U3701 (N_3701,N_3078,N_2492);
and U3702 (N_3702,N_3262,N_3479);
xor U3703 (N_3703,N_3239,N_2801);
and U3704 (N_3704,N_3279,N_2586);
or U3705 (N_3705,N_3122,N_2867);
and U3706 (N_3706,N_2584,N_3045);
nor U3707 (N_3707,N_2737,N_3264);
and U3708 (N_3708,N_3238,N_2757);
nand U3709 (N_3709,N_3367,N_2676);
and U3710 (N_3710,N_3253,N_3035);
and U3711 (N_3711,N_2702,N_2413);
or U3712 (N_3712,N_2843,N_3499);
and U3713 (N_3713,N_2882,N_2455);
nand U3714 (N_3714,N_2529,N_3200);
nand U3715 (N_3715,N_3523,N_2855);
nand U3716 (N_3716,N_2610,N_2511);
nand U3717 (N_3717,N_2930,N_3577);
or U3718 (N_3718,N_3559,N_2720);
nor U3719 (N_3719,N_2432,N_3134);
nand U3720 (N_3720,N_2797,N_3568);
nand U3721 (N_3721,N_2766,N_2947);
and U3722 (N_3722,N_3041,N_2502);
or U3723 (N_3723,N_2570,N_3437);
nor U3724 (N_3724,N_3289,N_2431);
and U3725 (N_3725,N_3429,N_2624);
xnor U3726 (N_3726,N_2949,N_2490);
or U3727 (N_3727,N_3233,N_3127);
nand U3728 (N_3728,N_2920,N_2727);
or U3729 (N_3729,N_3369,N_2747);
nor U3730 (N_3730,N_3580,N_3276);
xor U3731 (N_3731,N_2885,N_3282);
or U3732 (N_3732,N_3133,N_3225);
and U3733 (N_3733,N_2959,N_3068);
xor U3734 (N_3734,N_2470,N_3406);
xnor U3735 (N_3735,N_3560,N_2934);
nand U3736 (N_3736,N_2963,N_2850);
or U3737 (N_3737,N_2636,N_3104);
xor U3738 (N_3738,N_3448,N_3495);
nor U3739 (N_3739,N_2939,N_3468);
nor U3740 (N_3740,N_3573,N_3162);
or U3741 (N_3741,N_3269,N_3417);
nor U3742 (N_3742,N_3387,N_2666);
xor U3743 (N_3743,N_3572,N_2488);
nand U3744 (N_3744,N_3316,N_2749);
nor U3745 (N_3745,N_2950,N_3440);
and U3746 (N_3746,N_2465,N_3235);
and U3747 (N_3747,N_2648,N_2450);
or U3748 (N_3748,N_2561,N_3413);
nor U3749 (N_3749,N_3152,N_2554);
or U3750 (N_3750,N_2897,N_2700);
nand U3751 (N_3751,N_3187,N_2630);
or U3752 (N_3752,N_2659,N_3328);
or U3753 (N_3753,N_3280,N_3561);
and U3754 (N_3754,N_3503,N_2919);
nor U3755 (N_3755,N_3485,N_3224);
xor U3756 (N_3756,N_2803,N_3237);
or U3757 (N_3757,N_3218,N_3208);
or U3758 (N_3758,N_2547,N_2602);
xnor U3759 (N_3759,N_3201,N_3331);
xnor U3760 (N_3760,N_3326,N_2612);
nor U3761 (N_3761,N_3596,N_3337);
nor U3762 (N_3762,N_2923,N_2471);
or U3763 (N_3763,N_3119,N_3586);
xor U3764 (N_3764,N_3590,N_3139);
and U3765 (N_3765,N_2458,N_2960);
xor U3766 (N_3766,N_3403,N_2714);
or U3767 (N_3767,N_2725,N_2733);
or U3768 (N_3768,N_3589,N_2412);
or U3769 (N_3769,N_3093,N_2410);
or U3770 (N_3770,N_3259,N_2408);
or U3771 (N_3771,N_2646,N_2790);
nor U3772 (N_3772,N_2945,N_2978);
or U3773 (N_3773,N_3498,N_3098);
xnor U3774 (N_3774,N_2704,N_3421);
nand U3775 (N_3775,N_3011,N_2852);
nand U3776 (N_3776,N_2812,N_3582);
or U3777 (N_3777,N_2781,N_3362);
xnor U3778 (N_3778,N_3542,N_3063);
or U3779 (N_3779,N_2895,N_2528);
nand U3780 (N_3780,N_2708,N_2556);
xor U3781 (N_3781,N_2469,N_3303);
or U3782 (N_3782,N_3009,N_2601);
xnor U3783 (N_3783,N_2642,N_3296);
nor U3784 (N_3784,N_2451,N_3124);
and U3785 (N_3785,N_3502,N_3204);
xor U3786 (N_3786,N_3583,N_2649);
nor U3787 (N_3787,N_2827,N_3058);
nor U3788 (N_3788,N_3443,N_3113);
nor U3789 (N_3789,N_3013,N_2877);
and U3790 (N_3790,N_2841,N_3400);
xor U3791 (N_3791,N_3106,N_2993);
or U3792 (N_3792,N_2446,N_3450);
nor U3793 (N_3793,N_2481,N_2971);
or U3794 (N_3794,N_3105,N_2401);
or U3795 (N_3795,N_2763,N_3494);
and U3796 (N_3796,N_2441,N_2946);
nand U3797 (N_3797,N_3527,N_2938);
nand U3798 (N_3798,N_2907,N_3216);
xor U3799 (N_3799,N_2994,N_2503);
or U3800 (N_3800,N_2752,N_2991);
xor U3801 (N_3801,N_3241,N_3433);
xnor U3802 (N_3802,N_2767,N_3252);
or U3803 (N_3803,N_2536,N_2924);
nand U3804 (N_3804,N_3383,N_2574);
and U3805 (N_3805,N_2979,N_2523);
nand U3806 (N_3806,N_2901,N_3483);
and U3807 (N_3807,N_3148,N_3512);
nor U3808 (N_3808,N_2452,N_2900);
and U3809 (N_3809,N_2872,N_2771);
nor U3810 (N_3810,N_3090,N_3404);
xnor U3811 (N_3811,N_3351,N_2499);
or U3812 (N_3812,N_3436,N_3489);
nand U3813 (N_3813,N_3299,N_3425);
or U3814 (N_3814,N_3524,N_2500);
and U3815 (N_3815,N_2669,N_3381);
nor U3816 (N_3816,N_3385,N_2517);
nor U3817 (N_3817,N_2407,N_3447);
xnor U3818 (N_3818,N_3172,N_3052);
xnor U3819 (N_3819,N_2986,N_2888);
xnor U3820 (N_3820,N_2531,N_3505);
or U3821 (N_3821,N_2501,N_2896);
nor U3822 (N_3822,N_2520,N_2678);
xnor U3823 (N_3823,N_2448,N_2644);
xor U3824 (N_3824,N_3183,N_2764);
nor U3825 (N_3825,N_3576,N_3354);
xnor U3826 (N_3826,N_2638,N_3285);
or U3827 (N_3827,N_2656,N_3091);
nor U3828 (N_3828,N_2833,N_3344);
nor U3829 (N_3829,N_2707,N_2858);
nor U3830 (N_3830,N_3541,N_3408);
or U3831 (N_3831,N_2869,N_3537);
nor U3832 (N_3832,N_3121,N_3182);
or U3833 (N_3833,N_2650,N_2889);
xnor U3834 (N_3834,N_3205,N_3202);
or U3835 (N_3835,N_3175,N_3442);
xor U3836 (N_3836,N_2614,N_3033);
nor U3837 (N_3837,N_2716,N_2689);
xor U3838 (N_3838,N_3357,N_3540);
xor U3839 (N_3839,N_3327,N_3308);
and U3840 (N_3840,N_2824,N_3571);
xnor U3841 (N_3841,N_3379,N_3153);
xor U3842 (N_3842,N_2526,N_2730);
and U3843 (N_3843,N_2527,N_3438);
or U3844 (N_3844,N_3564,N_3173);
and U3845 (N_3845,N_3397,N_2918);
xnor U3846 (N_3846,N_2694,N_3003);
nand U3847 (N_3847,N_2438,N_2904);
nor U3848 (N_3848,N_2954,N_2628);
nor U3849 (N_3849,N_2686,N_3548);
or U3850 (N_3850,N_2854,N_2795);
or U3851 (N_3851,N_3008,N_3240);
and U3852 (N_3852,N_2988,N_2565);
nor U3853 (N_3853,N_2563,N_3446);
and U3854 (N_3854,N_2605,N_3000);
nor U3855 (N_3855,N_2731,N_3476);
and U3856 (N_3856,N_3118,N_3151);
nand U3857 (N_3857,N_3038,N_2404);
and U3858 (N_3858,N_2965,N_2775);
or U3859 (N_3859,N_2620,N_3346);
or U3860 (N_3860,N_3181,N_2639);
or U3861 (N_3861,N_2495,N_2744);
nor U3862 (N_3862,N_3165,N_3290);
nand U3863 (N_3863,N_3002,N_2980);
and U3864 (N_3864,N_3420,N_3488);
or U3865 (N_3865,N_2685,N_2621);
xor U3866 (N_3866,N_2472,N_2932);
xor U3867 (N_3867,N_3598,N_2710);
or U3868 (N_3868,N_3352,N_3522);
xor U3869 (N_3869,N_3467,N_3199);
and U3870 (N_3870,N_3558,N_2890);
nand U3871 (N_3871,N_2736,N_3550);
and U3872 (N_3872,N_2847,N_3195);
nand U3873 (N_3873,N_3287,N_2846);
xnor U3874 (N_3874,N_3076,N_3526);
and U3875 (N_3875,N_2968,N_3242);
nor U3876 (N_3876,N_3422,N_3191);
nor U3877 (N_3877,N_2955,N_2672);
nand U3878 (N_3878,N_3386,N_3380);
nand U3879 (N_3879,N_2560,N_2906);
or U3880 (N_3880,N_2820,N_2544);
xnor U3881 (N_3881,N_2972,N_2784);
xnor U3882 (N_3882,N_2785,N_3178);
xnor U3883 (N_3883,N_2582,N_3591);
and U3884 (N_3884,N_2466,N_2421);
nor U3885 (N_3885,N_3074,N_3217);
nor U3886 (N_3886,N_3141,N_3567);
nand U3887 (N_3887,N_3456,N_3057);
nor U3888 (N_3888,N_3266,N_3075);
or U3889 (N_3889,N_3222,N_3372);
and U3890 (N_3890,N_3257,N_3552);
nand U3891 (N_3891,N_2832,N_3261);
or U3892 (N_3892,N_3394,N_2974);
xnor U3893 (N_3893,N_2750,N_2665);
nor U3894 (N_3894,N_3170,N_2464);
xor U3895 (N_3895,N_2699,N_3026);
xnor U3896 (N_3896,N_2493,N_2461);
or U3897 (N_3897,N_2510,N_2695);
xnor U3898 (N_3898,N_3256,N_3497);
xnor U3899 (N_3899,N_3260,N_3402);
xor U3900 (N_3900,N_3249,N_2403);
or U3901 (N_3901,N_2796,N_3254);
and U3902 (N_3902,N_3270,N_2504);
and U3903 (N_3903,N_2936,N_2791);
nor U3904 (N_3904,N_2453,N_3189);
nor U3905 (N_3905,N_2698,N_2677);
or U3906 (N_3906,N_3444,N_3017);
and U3907 (N_3907,N_2984,N_2976);
xor U3908 (N_3908,N_2925,N_2673);
or U3909 (N_3909,N_3110,N_3309);
or U3910 (N_3910,N_2842,N_2798);
nand U3911 (N_3911,N_2879,N_3131);
and U3912 (N_3912,N_3455,N_2668);
nand U3913 (N_3913,N_3518,N_3306);
nor U3914 (N_3914,N_3248,N_3325);
nand U3915 (N_3915,N_2629,N_2931);
nor U3916 (N_3916,N_2553,N_3016);
xnor U3917 (N_3917,N_3364,N_2829);
or U3918 (N_3918,N_2530,N_3069);
nor U3919 (N_3919,N_3157,N_3330);
and U3920 (N_3920,N_2870,N_3409);
xor U3921 (N_3921,N_2616,N_2723);
and U3922 (N_3922,N_2709,N_3504);
nor U3923 (N_3923,N_2802,N_2426);
nand U3924 (N_3924,N_2447,N_3168);
xor U3925 (N_3925,N_2524,N_3220);
nor U3926 (N_3926,N_2693,N_2683);
nor U3927 (N_3927,N_3245,N_3293);
nand U3928 (N_3928,N_2626,N_3111);
xnor U3929 (N_3929,N_3519,N_2770);
xor U3930 (N_3930,N_3012,N_3236);
nor U3931 (N_3931,N_3286,N_2647);
xor U3932 (N_3932,N_3449,N_3244);
xor U3933 (N_3933,N_3297,N_2825);
xor U3934 (N_3934,N_3506,N_3115);
and U3935 (N_3935,N_3203,N_2713);
nand U3936 (N_3936,N_2804,N_2908);
nor U3937 (N_3937,N_2653,N_2969);
xor U3938 (N_3938,N_2532,N_3336);
xnor U3939 (N_3939,N_2618,N_2782);
and U3940 (N_3940,N_3507,N_3365);
nand U3941 (N_3941,N_3324,N_3036);
nor U3942 (N_3942,N_2593,N_3508);
and U3943 (N_3943,N_3051,N_2837);
and U3944 (N_3944,N_3056,N_2758);
or U3945 (N_3945,N_3307,N_2754);
nor U3946 (N_3946,N_2681,N_2866);
or U3947 (N_3947,N_3004,N_3028);
and U3948 (N_3948,N_2794,N_3288);
nor U3949 (N_3949,N_3460,N_2533);
nand U3950 (N_3950,N_2691,N_3551);
or U3951 (N_3951,N_2899,N_3094);
or U3952 (N_3952,N_3304,N_3154);
nor U3953 (N_3953,N_3478,N_3229);
and U3954 (N_3954,N_3128,N_3545);
nand U3955 (N_3955,N_3474,N_3025);
xor U3956 (N_3956,N_2402,N_3072);
xor U3957 (N_3957,N_2596,N_3393);
xor U3958 (N_3958,N_2823,N_3037);
or U3959 (N_3959,N_3388,N_3378);
and U3960 (N_3960,N_3416,N_2405);
xnor U3961 (N_3961,N_2687,N_3250);
and U3962 (N_3962,N_2557,N_3130);
xor U3963 (N_3963,N_3079,N_3109);
nand U3964 (N_3964,N_3137,N_3441);
xnor U3965 (N_3965,N_2948,N_2615);
nor U3966 (N_3966,N_2859,N_2587);
xor U3967 (N_3967,N_3070,N_3143);
or U3968 (N_3968,N_2512,N_2828);
and U3969 (N_3969,N_2776,N_2418);
xnor U3970 (N_3970,N_3395,N_2562);
and U3971 (N_3971,N_2898,N_3569);
and U3972 (N_3972,N_3155,N_3120);
nor U3973 (N_3973,N_2912,N_3247);
xnor U3974 (N_3974,N_2423,N_3515);
nor U3975 (N_3975,N_2838,N_2496);
nor U3976 (N_3976,N_3465,N_2883);
or U3977 (N_3977,N_2711,N_2805);
nor U3978 (N_3978,N_3043,N_3592);
nor U3979 (N_3979,N_3376,N_2588);
xnor U3980 (N_3980,N_2483,N_2541);
and U3981 (N_3981,N_2937,N_3197);
nor U3982 (N_3982,N_3096,N_2579);
or U3983 (N_3983,N_3430,N_2592);
nand U3984 (N_3984,N_2551,N_2844);
nor U3985 (N_3985,N_2657,N_3164);
nand U3986 (N_3986,N_3274,N_3481);
or U3987 (N_3987,N_2475,N_2674);
xor U3988 (N_3988,N_2439,N_2941);
nor U3989 (N_3989,N_2886,N_2622);
nor U3990 (N_3990,N_2831,N_2857);
and U3991 (N_3991,N_2679,N_2575);
and U3992 (N_3992,N_3546,N_2853);
nand U3993 (N_3993,N_3377,N_2734);
nand U3994 (N_3994,N_3223,N_3356);
xor U3995 (N_3995,N_2428,N_3486);
and U3996 (N_3996,N_2419,N_3370);
nor U3997 (N_3997,N_2909,N_2773);
and U3998 (N_3998,N_2848,N_2430);
nor U3999 (N_3999,N_2958,N_2861);
and U4000 (N_4000,N_3445,N_2548);
or U4001 (N_4001,N_2459,N_3080);
xor U4002 (N_4002,N_2970,N_2778);
or U4003 (N_4003,N_3024,N_2769);
or U4004 (N_4004,N_2623,N_2456);
xor U4005 (N_4005,N_2826,N_2537);
or U4006 (N_4006,N_3575,N_3010);
or U4007 (N_4007,N_2696,N_3475);
xor U4008 (N_4008,N_3281,N_3015);
and U4009 (N_4009,N_2486,N_3353);
or U4010 (N_4010,N_2462,N_2815);
nor U4011 (N_4011,N_2755,N_2440);
or U4012 (N_4012,N_2444,N_3064);
nor U4013 (N_4013,N_2992,N_2522);
and U4014 (N_4014,N_3194,N_3192);
and U4015 (N_4015,N_2604,N_3092);
or U4016 (N_4016,N_3544,N_2542);
nand U4017 (N_4017,N_3427,N_2578);
xor U4018 (N_4018,N_2540,N_3410);
and U4019 (N_4019,N_3361,N_2590);
xor U4020 (N_4020,N_3384,N_3496);
or U4021 (N_4021,N_3129,N_3536);
nand U4022 (N_4022,N_3340,N_2667);
or U4023 (N_4023,N_2808,N_3059);
or U4024 (N_4024,N_2748,N_3230);
xnor U4025 (N_4025,N_3176,N_2597);
or U4026 (N_4026,N_3031,N_2474);
nand U4027 (N_4027,N_2416,N_3424);
xor U4028 (N_4028,N_3019,N_3088);
and U4029 (N_4029,N_3273,N_3283);
or U4030 (N_4030,N_2952,N_2839);
and U4031 (N_4031,N_3333,N_2814);
xnor U4032 (N_4032,N_3298,N_3345);
and U4033 (N_4033,N_3392,N_2821);
and U4034 (N_4034,N_2429,N_2929);
and U4035 (N_4035,N_3407,N_3431);
and U4036 (N_4036,N_2816,N_2606);
nand U4037 (N_4037,N_3310,N_2661);
nor U4038 (N_4038,N_3597,N_3292);
xor U4039 (N_4039,N_2538,N_3584);
nand U4040 (N_4040,N_2573,N_2518);
nand U4041 (N_4041,N_2989,N_3018);
and U4042 (N_4042,N_2564,N_3255);
or U4043 (N_4043,N_3044,N_3167);
nor U4044 (N_4044,N_2774,N_2975);
or U4045 (N_4045,N_2515,N_3179);
nand U4046 (N_4046,N_2962,N_3501);
xor U4047 (N_4047,N_2479,N_3005);
xnor U4048 (N_4048,N_3439,N_3062);
and U4049 (N_4049,N_3190,N_2435);
and U4050 (N_4050,N_2572,N_3458);
nand U4051 (N_4051,N_2706,N_2445);
and U4052 (N_4052,N_3428,N_2436);
or U4053 (N_4053,N_3570,N_2467);
and U4054 (N_4054,N_2873,N_2759);
nor U4055 (N_4055,N_2480,N_3169);
nand U4056 (N_4056,N_3343,N_2598);
xnor U4057 (N_4057,N_3579,N_3258);
and U4058 (N_4058,N_2715,N_2631);
and U4059 (N_4059,N_2881,N_3272);
nand U4060 (N_4060,N_3086,N_2760);
xor U4061 (N_4061,N_2880,N_3100);
nand U4062 (N_4062,N_2660,N_3480);
or U4063 (N_4063,N_2765,N_2806);
nor U4064 (N_4064,N_3147,N_2454);
xor U4065 (N_4065,N_3066,N_3532);
nor U4066 (N_4066,N_2651,N_3032);
nand U4067 (N_4067,N_3040,N_3215);
xor U4068 (N_4068,N_2995,N_3211);
nand U4069 (N_4069,N_3313,N_3097);
or U4070 (N_4070,N_3347,N_2641);
nor U4071 (N_4071,N_3030,N_3207);
nand U4072 (N_4072,N_3135,N_2830);
nor U4073 (N_4073,N_2875,N_2729);
xor U4074 (N_4074,N_2463,N_3084);
nand U4075 (N_4075,N_2745,N_3089);
nand U4076 (N_4076,N_3001,N_3484);
or U4077 (N_4077,N_3457,N_3513);
nand U4078 (N_4078,N_3267,N_3232);
nor U4079 (N_4079,N_3516,N_2724);
nor U4080 (N_4080,N_2868,N_3534);
and U4081 (N_4081,N_2973,N_2910);
and U4082 (N_4082,N_3426,N_3553);
or U4083 (N_4083,N_2772,N_2697);
xnor U4084 (N_4084,N_2990,N_2743);
nor U4085 (N_4085,N_3543,N_2534);
nand U4086 (N_4086,N_2787,N_2634);
xnor U4087 (N_4087,N_2983,N_3349);
and U4088 (N_4088,N_3246,N_3348);
nand U4089 (N_4089,N_3284,N_3023);
nand U4090 (N_4090,N_2999,N_2793);
xnor U4091 (N_4091,N_3473,N_3396);
nor U4092 (N_4092,N_2943,N_2701);
xnor U4093 (N_4093,N_2568,N_3158);
nand U4094 (N_4094,N_3186,N_2688);
nand U4095 (N_4095,N_3423,N_3212);
xnor U4096 (N_4096,N_3107,N_3160);
nor U4097 (N_4097,N_3463,N_2519);
xnor U4098 (N_4098,N_2477,N_3419);
or U4099 (N_4099,N_2535,N_2555);
nand U4100 (N_4100,N_3454,N_2433);
or U4101 (N_4101,N_3462,N_2569);
and U4102 (N_4102,N_2705,N_3085);
and U4103 (N_4103,N_3350,N_2751);
xnor U4104 (N_4104,N_2539,N_2690);
and U4105 (N_4105,N_3050,N_3123);
and U4106 (N_4106,N_2558,N_2409);
xnor U4107 (N_4107,N_3101,N_2902);
nand U4108 (N_4108,N_2521,N_2422);
or U4109 (N_4109,N_3477,N_3061);
nand U4110 (N_4110,N_2840,N_3209);
nand U4111 (N_4111,N_3585,N_2921);
nand U4112 (N_4112,N_3415,N_3268);
nand U4113 (N_4113,N_2655,N_2443);
and U4114 (N_4114,N_3087,N_2762);
and U4115 (N_4115,N_3588,N_3315);
and U4116 (N_4116,N_2633,N_2783);
or U4117 (N_4117,N_2756,N_2807);
nor U4118 (N_4118,N_3291,N_2887);
nand U4119 (N_4119,N_3042,N_3311);
xnor U4120 (N_4120,N_2583,N_3487);
nor U4121 (N_4121,N_3314,N_2603);
xnor U4122 (N_4122,N_3184,N_3451);
nand U4123 (N_4123,N_2411,N_2817);
or U4124 (N_4124,N_3566,N_2594);
or U4125 (N_4125,N_3196,N_3562);
nor U4126 (N_4126,N_3055,N_2434);
nand U4127 (N_4127,N_3103,N_3065);
or U4128 (N_4128,N_2482,N_2786);
or U4129 (N_4129,N_2811,N_3166);
nand U4130 (N_4130,N_2768,N_3539);
and U4131 (N_4131,N_3054,N_2914);
nand U4132 (N_4132,N_2722,N_3317);
or U4133 (N_4133,N_3300,N_3095);
or U4134 (N_4134,N_2585,N_2917);
or U4135 (N_4135,N_3213,N_2726);
xnor U4136 (N_4136,N_2684,N_3529);
nand U4137 (N_4137,N_2506,N_2862);
or U4138 (N_4138,N_2627,N_2956);
nor U4139 (N_4139,N_2497,N_2719);
xnor U4140 (N_4140,N_2735,N_2927);
nand U4141 (N_4141,N_2581,N_3302);
nor U4142 (N_4142,N_2654,N_2663);
or U4143 (N_4143,N_2813,N_3338);
xor U4144 (N_4144,N_2864,N_3234);
or U4145 (N_4145,N_3321,N_3053);
xnor U4146 (N_4146,N_3594,N_3509);
or U4147 (N_4147,N_3492,N_2915);
nand U4148 (N_4148,N_2712,N_3117);
nor U4149 (N_4149,N_2525,N_2957);
or U4150 (N_4150,N_2460,N_2543);
or U4151 (N_4151,N_2589,N_2779);
xnor U4152 (N_4152,N_3140,N_2613);
xnor U4153 (N_4153,N_3471,N_3263);
and U4154 (N_4154,N_3411,N_2427);
xnor U4155 (N_4155,N_2738,N_2425);
and U4156 (N_4156,N_3228,N_3047);
and U4157 (N_4157,N_2834,N_2546);
xnor U4158 (N_4158,N_3081,N_3125);
nand U4159 (N_4159,N_3531,N_2928);
nor U4160 (N_4160,N_3374,N_2577);
nand U4161 (N_4161,N_2894,N_3214);
nor U4162 (N_4162,N_2998,N_3554);
or U4163 (N_4163,N_2933,N_2576);
nor U4164 (N_4164,N_3226,N_3227);
and U4165 (N_4165,N_3149,N_2643);
nor U4166 (N_4166,N_3265,N_2670);
and U4167 (N_4167,N_3231,N_2498);
and U4168 (N_4168,N_3312,N_2437);
nand U4169 (N_4169,N_3029,N_2967);
xor U4170 (N_4170,N_3144,N_2780);
or U4171 (N_4171,N_2508,N_2865);
nor U4172 (N_4172,N_3067,N_2819);
nand U4173 (N_4173,N_3295,N_3358);
xnor U4174 (N_4174,N_2625,N_2891);
or U4175 (N_4175,N_3375,N_3177);
xnor U4176 (N_4176,N_2566,N_3371);
nor U4177 (N_4177,N_3145,N_3198);
nand U4178 (N_4178,N_2935,N_3574);
or U4179 (N_4179,N_2836,N_3556);
and U4180 (N_4180,N_3007,N_3435);
nand U4181 (N_4181,N_2692,N_2478);
or U4182 (N_4182,N_2835,N_3271);
nand U4183 (N_4183,N_3116,N_2671);
or U4184 (N_4184,N_2617,N_2818);
xnor U4185 (N_4185,N_2987,N_3022);
xnor U4186 (N_4186,N_2951,N_2851);
nand U4187 (N_4187,N_3185,N_2977);
nand U4188 (N_4188,N_3034,N_3126);
or U4189 (N_4189,N_2545,N_2940);
nand U4190 (N_4190,N_3021,N_2944);
and U4191 (N_4191,N_3533,N_3163);
xnor U4192 (N_4192,N_2609,N_3514);
nand U4193 (N_4193,N_2892,N_2742);
nand U4194 (N_4194,N_2611,N_3305);
nor U4195 (N_4195,N_3360,N_3373);
nand U4196 (N_4196,N_3210,N_3320);
xor U4197 (N_4197,N_3318,N_3405);
nand U4198 (N_4198,N_2513,N_2860);
or U4199 (N_4199,N_3083,N_3355);
xor U4200 (N_4200,N_2796,N_3513);
and U4201 (N_4201,N_2479,N_3545);
xnor U4202 (N_4202,N_3228,N_3331);
xnor U4203 (N_4203,N_2483,N_3403);
nor U4204 (N_4204,N_2440,N_2835);
xor U4205 (N_4205,N_2871,N_3440);
xor U4206 (N_4206,N_2793,N_3547);
or U4207 (N_4207,N_3103,N_2618);
and U4208 (N_4208,N_2699,N_3470);
or U4209 (N_4209,N_2670,N_2569);
or U4210 (N_4210,N_3159,N_3439);
nor U4211 (N_4211,N_3253,N_3208);
nand U4212 (N_4212,N_3564,N_3140);
nor U4213 (N_4213,N_3404,N_3271);
nor U4214 (N_4214,N_3408,N_3016);
and U4215 (N_4215,N_2772,N_2973);
nand U4216 (N_4216,N_2588,N_3531);
nor U4217 (N_4217,N_3190,N_2493);
and U4218 (N_4218,N_2832,N_2871);
nor U4219 (N_4219,N_2693,N_2435);
or U4220 (N_4220,N_2666,N_2583);
xor U4221 (N_4221,N_2589,N_3590);
nand U4222 (N_4222,N_3117,N_3489);
or U4223 (N_4223,N_3268,N_3278);
nor U4224 (N_4224,N_3567,N_3414);
xor U4225 (N_4225,N_3307,N_3540);
or U4226 (N_4226,N_2680,N_2692);
or U4227 (N_4227,N_2501,N_3202);
nor U4228 (N_4228,N_2609,N_3533);
nor U4229 (N_4229,N_3582,N_3228);
nand U4230 (N_4230,N_2616,N_3260);
xnor U4231 (N_4231,N_3113,N_2449);
nand U4232 (N_4232,N_3042,N_3562);
xnor U4233 (N_4233,N_3393,N_3341);
and U4234 (N_4234,N_3156,N_3506);
xor U4235 (N_4235,N_3176,N_3171);
and U4236 (N_4236,N_3479,N_3214);
xnor U4237 (N_4237,N_2567,N_3583);
xor U4238 (N_4238,N_3221,N_3186);
or U4239 (N_4239,N_2868,N_2540);
xor U4240 (N_4240,N_2523,N_3309);
xor U4241 (N_4241,N_2914,N_3566);
nor U4242 (N_4242,N_2640,N_3493);
nor U4243 (N_4243,N_2948,N_2540);
nor U4244 (N_4244,N_2865,N_3302);
nor U4245 (N_4245,N_3500,N_3066);
and U4246 (N_4246,N_3509,N_2854);
xnor U4247 (N_4247,N_2826,N_2681);
nand U4248 (N_4248,N_2632,N_2611);
nor U4249 (N_4249,N_2494,N_2430);
and U4250 (N_4250,N_2907,N_2725);
xnor U4251 (N_4251,N_3405,N_2725);
or U4252 (N_4252,N_2888,N_2601);
nor U4253 (N_4253,N_2641,N_2775);
or U4254 (N_4254,N_2726,N_2495);
and U4255 (N_4255,N_3592,N_3157);
and U4256 (N_4256,N_2636,N_2888);
and U4257 (N_4257,N_2769,N_3436);
nand U4258 (N_4258,N_3384,N_3320);
and U4259 (N_4259,N_2802,N_3458);
and U4260 (N_4260,N_3218,N_2891);
nor U4261 (N_4261,N_2424,N_3465);
nor U4262 (N_4262,N_2979,N_2531);
nor U4263 (N_4263,N_2791,N_2836);
nand U4264 (N_4264,N_3252,N_2716);
and U4265 (N_4265,N_2808,N_3287);
xnor U4266 (N_4266,N_3316,N_3579);
xor U4267 (N_4267,N_3546,N_3074);
nor U4268 (N_4268,N_2888,N_2646);
and U4269 (N_4269,N_2583,N_2629);
and U4270 (N_4270,N_3159,N_3352);
and U4271 (N_4271,N_3157,N_3443);
nor U4272 (N_4272,N_2600,N_3226);
nor U4273 (N_4273,N_3583,N_2581);
nand U4274 (N_4274,N_3352,N_3240);
and U4275 (N_4275,N_3393,N_2860);
xnor U4276 (N_4276,N_2778,N_2952);
and U4277 (N_4277,N_2889,N_2401);
or U4278 (N_4278,N_3445,N_2476);
and U4279 (N_4279,N_3509,N_2989);
and U4280 (N_4280,N_2966,N_3314);
and U4281 (N_4281,N_2925,N_2446);
nand U4282 (N_4282,N_2832,N_2591);
and U4283 (N_4283,N_3334,N_2578);
nor U4284 (N_4284,N_3303,N_3460);
or U4285 (N_4285,N_2703,N_3266);
or U4286 (N_4286,N_3313,N_2842);
nand U4287 (N_4287,N_2586,N_3380);
nand U4288 (N_4288,N_3553,N_3428);
xor U4289 (N_4289,N_3552,N_3174);
nand U4290 (N_4290,N_3439,N_3120);
and U4291 (N_4291,N_3524,N_3572);
nand U4292 (N_4292,N_2837,N_3520);
and U4293 (N_4293,N_2473,N_3250);
xnor U4294 (N_4294,N_3027,N_2783);
nand U4295 (N_4295,N_3145,N_3207);
and U4296 (N_4296,N_3369,N_3389);
xor U4297 (N_4297,N_2676,N_3587);
and U4298 (N_4298,N_2766,N_3424);
nand U4299 (N_4299,N_2523,N_3574);
or U4300 (N_4300,N_3114,N_3121);
xor U4301 (N_4301,N_2570,N_3344);
xnor U4302 (N_4302,N_2426,N_3550);
nand U4303 (N_4303,N_3367,N_3209);
and U4304 (N_4304,N_3101,N_3124);
xnor U4305 (N_4305,N_3463,N_3340);
nand U4306 (N_4306,N_3240,N_3468);
or U4307 (N_4307,N_2906,N_3102);
xnor U4308 (N_4308,N_3244,N_3518);
nor U4309 (N_4309,N_3049,N_3178);
nor U4310 (N_4310,N_2447,N_2992);
nor U4311 (N_4311,N_2420,N_2427);
xnor U4312 (N_4312,N_3442,N_3284);
xnor U4313 (N_4313,N_2677,N_2475);
xor U4314 (N_4314,N_2578,N_2448);
nor U4315 (N_4315,N_2421,N_3474);
nor U4316 (N_4316,N_2734,N_2430);
nand U4317 (N_4317,N_2402,N_3273);
or U4318 (N_4318,N_3312,N_2849);
xnor U4319 (N_4319,N_2577,N_3549);
and U4320 (N_4320,N_2951,N_3582);
xnor U4321 (N_4321,N_2925,N_2861);
and U4322 (N_4322,N_3132,N_2487);
or U4323 (N_4323,N_3064,N_3027);
nand U4324 (N_4324,N_3458,N_2470);
or U4325 (N_4325,N_2921,N_2583);
nor U4326 (N_4326,N_2709,N_3430);
or U4327 (N_4327,N_3168,N_2471);
or U4328 (N_4328,N_2750,N_2556);
xnor U4329 (N_4329,N_2986,N_3448);
or U4330 (N_4330,N_3433,N_2643);
nand U4331 (N_4331,N_3385,N_3328);
or U4332 (N_4332,N_2508,N_3033);
nand U4333 (N_4333,N_3556,N_3185);
and U4334 (N_4334,N_3365,N_2635);
nor U4335 (N_4335,N_2577,N_3320);
and U4336 (N_4336,N_3236,N_2796);
and U4337 (N_4337,N_2860,N_3109);
or U4338 (N_4338,N_2516,N_3120);
or U4339 (N_4339,N_3557,N_2572);
nor U4340 (N_4340,N_2658,N_3045);
nand U4341 (N_4341,N_2879,N_3239);
xor U4342 (N_4342,N_3087,N_3346);
and U4343 (N_4343,N_2961,N_3045);
xnor U4344 (N_4344,N_2981,N_3262);
nor U4345 (N_4345,N_2616,N_3498);
and U4346 (N_4346,N_3196,N_2751);
xor U4347 (N_4347,N_2593,N_3416);
xnor U4348 (N_4348,N_3206,N_3269);
and U4349 (N_4349,N_2905,N_2671);
nor U4350 (N_4350,N_3477,N_2728);
xnor U4351 (N_4351,N_2908,N_2429);
xnor U4352 (N_4352,N_2754,N_3429);
nand U4353 (N_4353,N_3488,N_3587);
xnor U4354 (N_4354,N_3321,N_3333);
nand U4355 (N_4355,N_3318,N_2659);
or U4356 (N_4356,N_2694,N_3340);
or U4357 (N_4357,N_2527,N_3318);
or U4358 (N_4358,N_3264,N_3020);
nand U4359 (N_4359,N_2450,N_2850);
nand U4360 (N_4360,N_3563,N_3301);
nand U4361 (N_4361,N_3436,N_2974);
nand U4362 (N_4362,N_3222,N_3457);
or U4363 (N_4363,N_2640,N_3540);
and U4364 (N_4364,N_2872,N_3449);
nand U4365 (N_4365,N_3164,N_3133);
or U4366 (N_4366,N_3360,N_3510);
or U4367 (N_4367,N_2978,N_2747);
and U4368 (N_4368,N_3463,N_2649);
and U4369 (N_4369,N_3133,N_2922);
nor U4370 (N_4370,N_3066,N_2847);
nand U4371 (N_4371,N_3289,N_3145);
and U4372 (N_4372,N_2914,N_3009);
nor U4373 (N_4373,N_2599,N_3361);
nor U4374 (N_4374,N_3386,N_2901);
xnor U4375 (N_4375,N_3549,N_3177);
nor U4376 (N_4376,N_2455,N_2507);
xor U4377 (N_4377,N_3527,N_2529);
nand U4378 (N_4378,N_3476,N_2932);
and U4379 (N_4379,N_3428,N_2427);
nand U4380 (N_4380,N_3305,N_2866);
nand U4381 (N_4381,N_2716,N_3247);
nor U4382 (N_4382,N_3004,N_2597);
xnor U4383 (N_4383,N_3177,N_2618);
xnor U4384 (N_4384,N_3497,N_2602);
or U4385 (N_4385,N_3317,N_3489);
xnor U4386 (N_4386,N_3317,N_3355);
xor U4387 (N_4387,N_2419,N_3230);
nor U4388 (N_4388,N_3347,N_3255);
nand U4389 (N_4389,N_2580,N_2936);
xor U4390 (N_4390,N_2515,N_2550);
nand U4391 (N_4391,N_2471,N_2693);
or U4392 (N_4392,N_2712,N_2457);
xor U4393 (N_4393,N_3307,N_2559);
and U4394 (N_4394,N_3472,N_2598);
xor U4395 (N_4395,N_2435,N_3040);
xor U4396 (N_4396,N_2526,N_3153);
nand U4397 (N_4397,N_2675,N_3569);
or U4398 (N_4398,N_3171,N_3518);
nand U4399 (N_4399,N_3275,N_3599);
nand U4400 (N_4400,N_3319,N_3536);
nand U4401 (N_4401,N_2872,N_3441);
xor U4402 (N_4402,N_2437,N_2495);
or U4403 (N_4403,N_3158,N_2440);
or U4404 (N_4404,N_3130,N_2884);
nand U4405 (N_4405,N_3547,N_2675);
nand U4406 (N_4406,N_3229,N_3524);
xor U4407 (N_4407,N_2658,N_3330);
xnor U4408 (N_4408,N_2427,N_2727);
or U4409 (N_4409,N_2777,N_2451);
or U4410 (N_4410,N_3028,N_3085);
nand U4411 (N_4411,N_2517,N_3027);
xnor U4412 (N_4412,N_3587,N_3446);
and U4413 (N_4413,N_2428,N_2983);
nand U4414 (N_4414,N_2925,N_2485);
nand U4415 (N_4415,N_2758,N_3112);
and U4416 (N_4416,N_2471,N_2892);
xnor U4417 (N_4417,N_3098,N_3448);
and U4418 (N_4418,N_2818,N_3354);
nor U4419 (N_4419,N_3550,N_2662);
nor U4420 (N_4420,N_2917,N_2804);
nor U4421 (N_4421,N_2783,N_2408);
nor U4422 (N_4422,N_3438,N_2447);
or U4423 (N_4423,N_2418,N_3053);
nand U4424 (N_4424,N_2553,N_2416);
xnor U4425 (N_4425,N_3076,N_3438);
and U4426 (N_4426,N_3289,N_2847);
or U4427 (N_4427,N_3447,N_2891);
xnor U4428 (N_4428,N_2438,N_3173);
nand U4429 (N_4429,N_2943,N_2885);
nor U4430 (N_4430,N_2966,N_3513);
xnor U4431 (N_4431,N_2750,N_2711);
and U4432 (N_4432,N_3014,N_3366);
nand U4433 (N_4433,N_2878,N_2896);
nor U4434 (N_4434,N_2529,N_3485);
xor U4435 (N_4435,N_3011,N_2525);
and U4436 (N_4436,N_2936,N_3394);
or U4437 (N_4437,N_2759,N_3390);
xor U4438 (N_4438,N_2480,N_2599);
nor U4439 (N_4439,N_3486,N_2458);
nor U4440 (N_4440,N_3418,N_3447);
nand U4441 (N_4441,N_2826,N_2500);
nand U4442 (N_4442,N_3389,N_3270);
or U4443 (N_4443,N_2491,N_2533);
nand U4444 (N_4444,N_2646,N_2819);
nand U4445 (N_4445,N_3173,N_3479);
and U4446 (N_4446,N_2934,N_3469);
and U4447 (N_4447,N_3275,N_2993);
and U4448 (N_4448,N_3524,N_2725);
or U4449 (N_4449,N_2771,N_3407);
and U4450 (N_4450,N_2901,N_2564);
or U4451 (N_4451,N_3003,N_3182);
xor U4452 (N_4452,N_3492,N_2430);
or U4453 (N_4453,N_3475,N_2923);
nand U4454 (N_4454,N_2687,N_2993);
nor U4455 (N_4455,N_3102,N_3498);
or U4456 (N_4456,N_3369,N_2624);
nand U4457 (N_4457,N_2710,N_2533);
nor U4458 (N_4458,N_2419,N_2432);
and U4459 (N_4459,N_3003,N_2617);
and U4460 (N_4460,N_2824,N_3114);
and U4461 (N_4461,N_3203,N_3123);
nor U4462 (N_4462,N_2677,N_2607);
xor U4463 (N_4463,N_2685,N_2566);
nand U4464 (N_4464,N_2472,N_2773);
nor U4465 (N_4465,N_3445,N_2786);
and U4466 (N_4466,N_2857,N_2538);
and U4467 (N_4467,N_2678,N_2500);
or U4468 (N_4468,N_2419,N_3098);
nor U4469 (N_4469,N_3457,N_2880);
xor U4470 (N_4470,N_3465,N_3171);
and U4471 (N_4471,N_3484,N_3494);
nor U4472 (N_4472,N_2614,N_3394);
nor U4473 (N_4473,N_2409,N_3329);
xnor U4474 (N_4474,N_2659,N_3197);
or U4475 (N_4475,N_2709,N_3248);
or U4476 (N_4476,N_3599,N_3294);
or U4477 (N_4477,N_2959,N_2674);
nand U4478 (N_4478,N_3397,N_3136);
or U4479 (N_4479,N_2706,N_3403);
xor U4480 (N_4480,N_3454,N_2883);
xor U4481 (N_4481,N_3081,N_3055);
or U4482 (N_4482,N_2841,N_2558);
nand U4483 (N_4483,N_2402,N_2946);
and U4484 (N_4484,N_2446,N_3227);
or U4485 (N_4485,N_2631,N_2984);
nand U4486 (N_4486,N_2993,N_3254);
xnor U4487 (N_4487,N_2795,N_2887);
nor U4488 (N_4488,N_3165,N_3396);
and U4489 (N_4489,N_3557,N_2542);
or U4490 (N_4490,N_2410,N_2488);
or U4491 (N_4491,N_2632,N_3051);
or U4492 (N_4492,N_2561,N_2732);
nor U4493 (N_4493,N_2886,N_3100);
nand U4494 (N_4494,N_3156,N_2726);
and U4495 (N_4495,N_3010,N_3548);
or U4496 (N_4496,N_3337,N_3548);
nor U4497 (N_4497,N_3178,N_3548);
nand U4498 (N_4498,N_3234,N_2803);
nand U4499 (N_4499,N_2689,N_2662);
or U4500 (N_4500,N_3103,N_3037);
nor U4501 (N_4501,N_2835,N_3073);
xor U4502 (N_4502,N_2962,N_3047);
nand U4503 (N_4503,N_3553,N_3015);
and U4504 (N_4504,N_3023,N_3329);
xnor U4505 (N_4505,N_2670,N_3077);
xor U4506 (N_4506,N_2729,N_2412);
nor U4507 (N_4507,N_2643,N_3091);
or U4508 (N_4508,N_3248,N_2549);
xnor U4509 (N_4509,N_3092,N_3211);
nand U4510 (N_4510,N_2881,N_2556);
and U4511 (N_4511,N_2569,N_2573);
nor U4512 (N_4512,N_3053,N_2764);
nand U4513 (N_4513,N_2745,N_3586);
nand U4514 (N_4514,N_3462,N_2662);
nor U4515 (N_4515,N_2956,N_3090);
and U4516 (N_4516,N_3257,N_2957);
and U4517 (N_4517,N_2893,N_3241);
xor U4518 (N_4518,N_2972,N_3212);
xnor U4519 (N_4519,N_3178,N_2994);
nor U4520 (N_4520,N_3531,N_3594);
xnor U4521 (N_4521,N_3431,N_2691);
nand U4522 (N_4522,N_2678,N_3061);
and U4523 (N_4523,N_2431,N_3447);
or U4524 (N_4524,N_2408,N_3342);
xnor U4525 (N_4525,N_2874,N_2993);
nand U4526 (N_4526,N_2766,N_3078);
nor U4527 (N_4527,N_2772,N_3504);
xor U4528 (N_4528,N_2902,N_3486);
and U4529 (N_4529,N_3395,N_3370);
nor U4530 (N_4530,N_2668,N_2746);
nand U4531 (N_4531,N_3131,N_3212);
nand U4532 (N_4532,N_3151,N_3535);
xnor U4533 (N_4533,N_3436,N_3233);
nand U4534 (N_4534,N_2631,N_3560);
xnor U4535 (N_4535,N_3081,N_2454);
xor U4536 (N_4536,N_3369,N_3234);
xnor U4537 (N_4537,N_2813,N_3423);
nand U4538 (N_4538,N_3116,N_2869);
nand U4539 (N_4539,N_3214,N_3575);
and U4540 (N_4540,N_2978,N_2911);
or U4541 (N_4541,N_2907,N_2867);
nor U4542 (N_4542,N_2790,N_3247);
nand U4543 (N_4543,N_3441,N_3304);
and U4544 (N_4544,N_3532,N_3062);
xor U4545 (N_4545,N_3214,N_3064);
and U4546 (N_4546,N_2537,N_2744);
xor U4547 (N_4547,N_2759,N_3143);
nor U4548 (N_4548,N_3459,N_2802);
nand U4549 (N_4549,N_2725,N_3368);
or U4550 (N_4550,N_2995,N_3510);
or U4551 (N_4551,N_3349,N_2670);
and U4552 (N_4552,N_2456,N_2794);
xor U4553 (N_4553,N_3452,N_3202);
nand U4554 (N_4554,N_3260,N_2494);
nor U4555 (N_4555,N_3269,N_3481);
nor U4556 (N_4556,N_2891,N_3132);
and U4557 (N_4557,N_3480,N_3458);
xnor U4558 (N_4558,N_2614,N_2592);
xnor U4559 (N_4559,N_3286,N_3469);
nor U4560 (N_4560,N_2628,N_2448);
and U4561 (N_4561,N_2826,N_3334);
and U4562 (N_4562,N_2444,N_3269);
or U4563 (N_4563,N_2797,N_2807);
xnor U4564 (N_4564,N_2611,N_3567);
nand U4565 (N_4565,N_3298,N_2823);
nor U4566 (N_4566,N_2658,N_2766);
and U4567 (N_4567,N_3584,N_2909);
or U4568 (N_4568,N_3365,N_2976);
and U4569 (N_4569,N_2419,N_2890);
nor U4570 (N_4570,N_3572,N_3194);
and U4571 (N_4571,N_3563,N_2585);
xor U4572 (N_4572,N_2932,N_2879);
nor U4573 (N_4573,N_3428,N_2472);
or U4574 (N_4574,N_2760,N_2788);
and U4575 (N_4575,N_3257,N_2873);
nor U4576 (N_4576,N_2805,N_2705);
xor U4577 (N_4577,N_2443,N_2881);
nand U4578 (N_4578,N_3556,N_3021);
xor U4579 (N_4579,N_2938,N_3302);
and U4580 (N_4580,N_3045,N_2744);
xor U4581 (N_4581,N_3342,N_3025);
xor U4582 (N_4582,N_3358,N_2655);
nand U4583 (N_4583,N_3563,N_3167);
nand U4584 (N_4584,N_2591,N_3357);
nor U4585 (N_4585,N_2985,N_3282);
and U4586 (N_4586,N_3492,N_3545);
nand U4587 (N_4587,N_3291,N_2594);
and U4588 (N_4588,N_3476,N_3431);
or U4589 (N_4589,N_3065,N_2719);
or U4590 (N_4590,N_3449,N_2420);
nand U4591 (N_4591,N_3487,N_2780);
nand U4592 (N_4592,N_2459,N_3094);
nand U4593 (N_4593,N_2764,N_3085);
or U4594 (N_4594,N_3173,N_2732);
and U4595 (N_4595,N_3087,N_3258);
xor U4596 (N_4596,N_2743,N_3390);
xor U4597 (N_4597,N_2824,N_2864);
and U4598 (N_4598,N_2932,N_3155);
xor U4599 (N_4599,N_3322,N_2584);
nand U4600 (N_4600,N_3587,N_3260);
and U4601 (N_4601,N_2561,N_2592);
or U4602 (N_4602,N_3034,N_3051);
nand U4603 (N_4603,N_2572,N_2995);
or U4604 (N_4604,N_2659,N_2783);
and U4605 (N_4605,N_2459,N_2658);
xnor U4606 (N_4606,N_2737,N_2762);
nor U4607 (N_4607,N_3206,N_3122);
and U4608 (N_4608,N_3536,N_3166);
nor U4609 (N_4609,N_2629,N_3145);
nand U4610 (N_4610,N_3198,N_2913);
nand U4611 (N_4611,N_3340,N_2813);
and U4612 (N_4612,N_3577,N_3405);
nand U4613 (N_4613,N_2527,N_3179);
or U4614 (N_4614,N_3340,N_3185);
or U4615 (N_4615,N_3165,N_3537);
or U4616 (N_4616,N_3198,N_2592);
or U4617 (N_4617,N_2744,N_2560);
xor U4618 (N_4618,N_3099,N_2798);
and U4619 (N_4619,N_2705,N_2751);
nand U4620 (N_4620,N_2814,N_2418);
and U4621 (N_4621,N_3182,N_2924);
or U4622 (N_4622,N_3114,N_2770);
xnor U4623 (N_4623,N_3360,N_2844);
xnor U4624 (N_4624,N_2863,N_2631);
nand U4625 (N_4625,N_3337,N_3159);
xnor U4626 (N_4626,N_3125,N_3378);
nor U4627 (N_4627,N_2647,N_2600);
or U4628 (N_4628,N_3237,N_2776);
or U4629 (N_4629,N_3068,N_2533);
nand U4630 (N_4630,N_2944,N_3226);
and U4631 (N_4631,N_2831,N_3277);
xor U4632 (N_4632,N_2660,N_3173);
or U4633 (N_4633,N_3422,N_3245);
nand U4634 (N_4634,N_2699,N_2670);
xor U4635 (N_4635,N_2614,N_2685);
xnor U4636 (N_4636,N_2771,N_3337);
nand U4637 (N_4637,N_3557,N_2817);
nor U4638 (N_4638,N_2926,N_3372);
and U4639 (N_4639,N_2437,N_2562);
and U4640 (N_4640,N_2926,N_2841);
xnor U4641 (N_4641,N_2731,N_3461);
nand U4642 (N_4642,N_2531,N_2427);
and U4643 (N_4643,N_3152,N_2680);
nor U4644 (N_4644,N_2542,N_2738);
xor U4645 (N_4645,N_2478,N_2463);
nor U4646 (N_4646,N_3203,N_2696);
nor U4647 (N_4647,N_3083,N_3033);
xnor U4648 (N_4648,N_2932,N_3042);
nand U4649 (N_4649,N_2904,N_3400);
xnor U4650 (N_4650,N_3505,N_3049);
or U4651 (N_4651,N_3467,N_3280);
xnor U4652 (N_4652,N_2548,N_2432);
and U4653 (N_4653,N_2517,N_3318);
or U4654 (N_4654,N_2464,N_2709);
xor U4655 (N_4655,N_2729,N_3218);
and U4656 (N_4656,N_2729,N_2869);
nand U4657 (N_4657,N_3409,N_2619);
or U4658 (N_4658,N_3319,N_2835);
and U4659 (N_4659,N_3265,N_2751);
xnor U4660 (N_4660,N_2712,N_3434);
xnor U4661 (N_4661,N_3109,N_3240);
xnor U4662 (N_4662,N_2953,N_2819);
or U4663 (N_4663,N_3468,N_2430);
nor U4664 (N_4664,N_3126,N_2501);
nor U4665 (N_4665,N_2792,N_3046);
or U4666 (N_4666,N_3191,N_3554);
xnor U4667 (N_4667,N_2514,N_3458);
nor U4668 (N_4668,N_3322,N_2829);
xor U4669 (N_4669,N_3146,N_3147);
and U4670 (N_4670,N_3075,N_2609);
xnor U4671 (N_4671,N_2531,N_2866);
xor U4672 (N_4672,N_3544,N_2858);
and U4673 (N_4673,N_2891,N_2627);
or U4674 (N_4674,N_2645,N_2806);
and U4675 (N_4675,N_2675,N_2482);
nand U4676 (N_4676,N_2953,N_3290);
or U4677 (N_4677,N_3346,N_2709);
nor U4678 (N_4678,N_3015,N_2605);
or U4679 (N_4679,N_2995,N_3314);
nor U4680 (N_4680,N_3448,N_3457);
nor U4681 (N_4681,N_3473,N_2897);
xor U4682 (N_4682,N_2994,N_2476);
and U4683 (N_4683,N_2521,N_3410);
and U4684 (N_4684,N_2979,N_2417);
xor U4685 (N_4685,N_3352,N_2407);
and U4686 (N_4686,N_3537,N_3392);
or U4687 (N_4687,N_3116,N_3146);
or U4688 (N_4688,N_3127,N_3463);
nand U4689 (N_4689,N_3541,N_2528);
nor U4690 (N_4690,N_3428,N_2402);
or U4691 (N_4691,N_3195,N_2541);
or U4692 (N_4692,N_3143,N_2673);
nor U4693 (N_4693,N_2486,N_3197);
xnor U4694 (N_4694,N_3389,N_3536);
nand U4695 (N_4695,N_3475,N_3430);
xor U4696 (N_4696,N_3115,N_3106);
xor U4697 (N_4697,N_2654,N_2910);
and U4698 (N_4698,N_2777,N_2942);
nand U4699 (N_4699,N_2868,N_3224);
nand U4700 (N_4700,N_2768,N_2514);
and U4701 (N_4701,N_3546,N_3483);
and U4702 (N_4702,N_3192,N_2511);
nand U4703 (N_4703,N_2904,N_2720);
nor U4704 (N_4704,N_2454,N_2497);
or U4705 (N_4705,N_3023,N_2502);
nand U4706 (N_4706,N_3260,N_2854);
and U4707 (N_4707,N_3416,N_3383);
nand U4708 (N_4708,N_3575,N_2974);
or U4709 (N_4709,N_2610,N_3150);
and U4710 (N_4710,N_2621,N_2675);
xnor U4711 (N_4711,N_2586,N_2854);
or U4712 (N_4712,N_3101,N_2793);
or U4713 (N_4713,N_2463,N_3220);
xor U4714 (N_4714,N_3007,N_3027);
and U4715 (N_4715,N_3170,N_3528);
xor U4716 (N_4716,N_3429,N_2985);
nand U4717 (N_4717,N_2890,N_3307);
or U4718 (N_4718,N_3247,N_3464);
or U4719 (N_4719,N_3222,N_2469);
or U4720 (N_4720,N_2529,N_2639);
nor U4721 (N_4721,N_3217,N_3441);
or U4722 (N_4722,N_3122,N_3445);
nor U4723 (N_4723,N_3213,N_2850);
nor U4724 (N_4724,N_2605,N_2521);
nand U4725 (N_4725,N_2940,N_3299);
xnor U4726 (N_4726,N_2702,N_3099);
nor U4727 (N_4727,N_3391,N_3255);
nor U4728 (N_4728,N_2837,N_3260);
nand U4729 (N_4729,N_2537,N_3345);
and U4730 (N_4730,N_3568,N_2753);
nor U4731 (N_4731,N_2480,N_3137);
nand U4732 (N_4732,N_3172,N_2595);
or U4733 (N_4733,N_3574,N_3301);
or U4734 (N_4734,N_2619,N_3280);
nand U4735 (N_4735,N_3137,N_3081);
and U4736 (N_4736,N_3591,N_3084);
nor U4737 (N_4737,N_2410,N_3500);
nor U4738 (N_4738,N_3436,N_3470);
nor U4739 (N_4739,N_3023,N_2804);
nand U4740 (N_4740,N_2797,N_3589);
or U4741 (N_4741,N_2809,N_3003);
and U4742 (N_4742,N_3576,N_3371);
nor U4743 (N_4743,N_2702,N_3088);
or U4744 (N_4744,N_3448,N_3015);
nor U4745 (N_4745,N_3488,N_3251);
xor U4746 (N_4746,N_3359,N_3075);
or U4747 (N_4747,N_2951,N_3580);
or U4748 (N_4748,N_2947,N_2525);
xnor U4749 (N_4749,N_3440,N_2761);
or U4750 (N_4750,N_3585,N_2485);
xor U4751 (N_4751,N_3255,N_2586);
xor U4752 (N_4752,N_3148,N_2788);
and U4753 (N_4753,N_2758,N_3046);
and U4754 (N_4754,N_2563,N_3408);
nor U4755 (N_4755,N_3269,N_2554);
xor U4756 (N_4756,N_3043,N_2867);
nand U4757 (N_4757,N_3598,N_2432);
or U4758 (N_4758,N_2611,N_3562);
or U4759 (N_4759,N_3232,N_2876);
and U4760 (N_4760,N_3501,N_2400);
nand U4761 (N_4761,N_3177,N_2668);
nand U4762 (N_4762,N_3406,N_3580);
and U4763 (N_4763,N_2531,N_2825);
or U4764 (N_4764,N_3468,N_3135);
or U4765 (N_4765,N_2646,N_3044);
and U4766 (N_4766,N_3301,N_2951);
nor U4767 (N_4767,N_3304,N_2835);
or U4768 (N_4768,N_3421,N_3202);
nor U4769 (N_4769,N_3186,N_3405);
or U4770 (N_4770,N_3098,N_3070);
or U4771 (N_4771,N_2835,N_2796);
nand U4772 (N_4772,N_2839,N_2470);
and U4773 (N_4773,N_3177,N_3252);
and U4774 (N_4774,N_3021,N_3417);
nor U4775 (N_4775,N_3144,N_3266);
xnor U4776 (N_4776,N_3328,N_2835);
and U4777 (N_4777,N_2683,N_2973);
xnor U4778 (N_4778,N_2976,N_2957);
xor U4779 (N_4779,N_3567,N_2414);
or U4780 (N_4780,N_2704,N_3158);
or U4781 (N_4781,N_3258,N_2993);
xnor U4782 (N_4782,N_3049,N_3192);
and U4783 (N_4783,N_2527,N_3402);
nand U4784 (N_4784,N_2724,N_3498);
xnor U4785 (N_4785,N_3034,N_2927);
nor U4786 (N_4786,N_2443,N_2644);
nor U4787 (N_4787,N_2991,N_3113);
or U4788 (N_4788,N_3200,N_3587);
and U4789 (N_4789,N_3237,N_2489);
or U4790 (N_4790,N_2408,N_3451);
and U4791 (N_4791,N_3109,N_3211);
or U4792 (N_4792,N_3373,N_3422);
and U4793 (N_4793,N_3249,N_2633);
nand U4794 (N_4794,N_2845,N_2973);
nor U4795 (N_4795,N_2988,N_3060);
nand U4796 (N_4796,N_2526,N_3446);
or U4797 (N_4797,N_3559,N_3176);
xnor U4798 (N_4798,N_2838,N_3312);
nand U4799 (N_4799,N_2547,N_2958);
or U4800 (N_4800,N_4284,N_3963);
nand U4801 (N_4801,N_4692,N_4635);
nand U4802 (N_4802,N_4526,N_3714);
or U4803 (N_4803,N_4408,N_4787);
nand U4804 (N_4804,N_4769,N_3787);
and U4805 (N_4805,N_4690,N_4420);
nor U4806 (N_4806,N_4114,N_4219);
nor U4807 (N_4807,N_4424,N_4516);
and U4808 (N_4808,N_3668,N_4412);
nor U4809 (N_4809,N_4224,N_4524);
xnor U4810 (N_4810,N_3600,N_4358);
nand U4811 (N_4811,N_3933,N_4538);
xor U4812 (N_4812,N_4044,N_3643);
nor U4813 (N_4813,N_4689,N_4318);
xor U4814 (N_4814,N_4489,N_4392);
nand U4815 (N_4815,N_4419,N_3716);
and U4816 (N_4816,N_3723,N_4167);
and U4817 (N_4817,N_3947,N_4555);
and U4818 (N_4818,N_4055,N_4504);
nand U4819 (N_4819,N_4141,N_3609);
nand U4820 (N_4820,N_3601,N_4462);
and U4821 (N_4821,N_4662,N_4432);
xnor U4822 (N_4822,N_3684,N_3727);
xnor U4823 (N_4823,N_4700,N_4361);
or U4824 (N_4824,N_4716,N_4610);
and U4825 (N_4825,N_4742,N_4630);
xor U4826 (N_4826,N_4456,N_4477);
nor U4827 (N_4827,N_4520,N_4152);
xnor U4828 (N_4828,N_3743,N_3917);
nand U4829 (N_4829,N_4228,N_3769);
nand U4830 (N_4830,N_4046,N_4168);
nand U4831 (N_4831,N_3809,N_4193);
or U4832 (N_4832,N_4666,N_4011);
xor U4833 (N_4833,N_3793,N_3756);
xor U4834 (N_4834,N_3670,N_4080);
nand U4835 (N_4835,N_4104,N_3748);
or U4836 (N_4836,N_4528,N_4235);
nand U4837 (N_4837,N_4664,N_3613);
nand U4838 (N_4838,N_4650,N_4066);
or U4839 (N_4839,N_4745,N_4118);
or U4840 (N_4840,N_3946,N_4058);
and U4841 (N_4841,N_4561,N_3844);
or U4842 (N_4842,N_3970,N_4498);
nand U4843 (N_4843,N_3812,N_4023);
and U4844 (N_4844,N_3894,N_4202);
xnor U4845 (N_4845,N_4337,N_4531);
xor U4846 (N_4846,N_4329,N_3636);
nand U4847 (N_4847,N_4290,N_4435);
xnor U4848 (N_4848,N_4026,N_4161);
xor U4849 (N_4849,N_4427,N_4774);
and U4850 (N_4850,N_4206,N_3721);
xor U4851 (N_4851,N_4410,N_4316);
nor U4852 (N_4852,N_4506,N_4281);
nor U4853 (N_4853,N_4695,N_3945);
nand U4854 (N_4854,N_4325,N_4364);
xnor U4855 (N_4855,N_4301,N_4203);
nor U4856 (N_4856,N_4607,N_4400);
nand U4857 (N_4857,N_3685,N_4214);
or U4858 (N_4858,N_4128,N_3610);
and U4859 (N_4859,N_4215,N_3842);
nand U4860 (N_4860,N_4150,N_3954);
and U4861 (N_4861,N_4580,N_3871);
nor U4862 (N_4862,N_4793,N_3629);
nand U4863 (N_4863,N_4629,N_4048);
or U4864 (N_4864,N_4699,N_4776);
or U4865 (N_4865,N_3914,N_3766);
nor U4866 (N_4866,N_4078,N_4429);
nor U4867 (N_4867,N_3648,N_4166);
nand U4868 (N_4868,N_4094,N_4522);
nand U4869 (N_4869,N_3857,N_4292);
nor U4870 (N_4870,N_4233,N_3885);
or U4871 (N_4871,N_4391,N_3759);
and U4872 (N_4872,N_4602,N_3941);
xnor U4873 (N_4873,N_4025,N_4398);
nor U4874 (N_4874,N_4672,N_4728);
nand U4875 (N_4875,N_3650,N_4190);
and U4876 (N_4876,N_4648,N_4705);
nor U4877 (N_4877,N_3961,N_3700);
or U4878 (N_4878,N_4009,N_4668);
nand U4879 (N_4879,N_4527,N_4688);
and U4880 (N_4880,N_4008,N_3794);
xnor U4881 (N_4881,N_4160,N_3798);
or U4882 (N_4882,N_4075,N_4485);
and U4883 (N_4883,N_3923,N_4343);
xnor U4884 (N_4884,N_3988,N_3697);
xor U4885 (N_4885,N_4523,N_4052);
and U4886 (N_4886,N_4208,N_3654);
xor U4887 (N_4887,N_3972,N_4661);
and U4888 (N_4888,N_3647,N_4680);
and U4889 (N_4889,N_3877,N_4546);
nor U4890 (N_4890,N_3757,N_4632);
xor U4891 (N_4891,N_3915,N_3819);
or U4892 (N_4892,N_4727,N_3804);
nor U4893 (N_4893,N_4714,N_4449);
xnor U4894 (N_4894,N_4162,N_4004);
and U4895 (N_4895,N_4022,N_4441);
xnor U4896 (N_4896,N_3679,N_4642);
or U4897 (N_4897,N_4102,N_3605);
and U4898 (N_4898,N_3918,N_3763);
or U4899 (N_4899,N_4274,N_4671);
nor U4900 (N_4900,N_3925,N_4216);
and U4901 (N_4901,N_4461,N_4431);
or U4902 (N_4902,N_4792,N_3806);
nand U4903 (N_4903,N_3847,N_3637);
and U4904 (N_4904,N_4592,N_4321);
and U4905 (N_4905,N_3775,N_3674);
nand U4906 (N_4906,N_3796,N_3661);
nand U4907 (N_4907,N_4576,N_4288);
or U4908 (N_4908,N_4605,N_4782);
nand U4909 (N_4909,N_4440,N_4260);
or U4910 (N_4910,N_3971,N_3996);
xnor U4911 (N_4911,N_4496,N_4594);
and U4912 (N_4912,N_4480,N_4289);
nor U4913 (N_4913,N_4652,N_4717);
or U4914 (N_4914,N_3864,N_4336);
xor U4915 (N_4915,N_4674,N_4346);
nand U4916 (N_4916,N_3858,N_4283);
nor U4917 (N_4917,N_4384,N_4054);
and U4918 (N_4918,N_3865,N_4194);
or U4919 (N_4919,N_4268,N_4320);
xnor U4920 (N_4920,N_4261,N_4556);
xor U4921 (N_4921,N_4334,N_3626);
nand U4922 (N_4922,N_4693,N_4421);
nand U4923 (N_4923,N_4665,N_4053);
nand U4924 (N_4924,N_3886,N_3976);
or U4925 (N_4925,N_3730,N_4359);
nor U4926 (N_4926,N_3777,N_4124);
and U4927 (N_4927,N_4568,N_4158);
or U4928 (N_4928,N_4579,N_4200);
nor U4929 (N_4929,N_3625,N_4192);
nand U4930 (N_4930,N_4088,N_3978);
nand U4931 (N_4931,N_3876,N_4638);
nand U4932 (N_4932,N_4402,N_4082);
and U4933 (N_4933,N_3772,N_4560);
nor U4934 (N_4934,N_3818,N_3632);
or U4935 (N_4935,N_3628,N_4112);
nor U4936 (N_4936,N_4309,N_4035);
nand U4937 (N_4937,N_3795,N_4731);
xor U4938 (N_4938,N_4375,N_3966);
and U4939 (N_4939,N_3874,N_3994);
or U4940 (N_4940,N_4433,N_3651);
nor U4941 (N_4941,N_4465,N_4582);
and U4942 (N_4942,N_4711,N_4682);
nor U4943 (N_4943,N_4533,N_4795);
nor U4944 (N_4944,N_3943,N_4659);
or U4945 (N_4945,N_4310,N_4209);
and U4946 (N_4946,N_4315,N_4735);
nand U4947 (N_4947,N_3630,N_3872);
xnor U4948 (N_4948,N_4415,N_3753);
nand U4949 (N_4949,N_4511,N_4324);
and U4950 (N_4950,N_4030,N_3764);
nand U4951 (N_4951,N_4157,N_4488);
nand U4952 (N_4952,N_4264,N_3658);
or U4953 (N_4953,N_4417,N_3786);
nor U4954 (N_4954,N_4354,N_3891);
or U4955 (N_4955,N_4684,N_4086);
nor U4956 (N_4956,N_3695,N_4332);
nand U4957 (N_4957,N_4487,N_4558);
or U4958 (N_4958,N_4482,N_3882);
nor U4959 (N_4959,N_4059,N_3694);
or U4960 (N_4960,N_4532,N_4351);
nand U4961 (N_4961,N_4033,N_3986);
nor U4962 (N_4962,N_4207,N_4484);
xor U4963 (N_4963,N_4767,N_4140);
or U4964 (N_4964,N_3672,N_3612);
xor U4965 (N_4965,N_4350,N_4238);
and U4966 (N_4966,N_3949,N_4541);
nor U4967 (N_4967,N_4521,N_3736);
and U4968 (N_4968,N_3724,N_4322);
or U4969 (N_4969,N_3895,N_4418);
xnor U4970 (N_4970,N_3706,N_3659);
xnor U4971 (N_4971,N_4317,N_3646);
and U4972 (N_4972,N_3951,N_4065);
and U4973 (N_4973,N_4414,N_4381);
or U4974 (N_4974,N_3603,N_4399);
or U4975 (N_4975,N_3619,N_4143);
nor U4976 (N_4976,N_4129,N_4411);
nand U4977 (N_4977,N_4464,N_4049);
xor U4978 (N_4978,N_3998,N_4603);
nand U4979 (N_4979,N_4244,N_4236);
nand U4980 (N_4980,N_3981,N_4438);
or U4981 (N_4981,N_4726,N_4308);
nand U4982 (N_4982,N_4515,N_3683);
nand U4983 (N_4983,N_4637,N_3653);
nor U4984 (N_4984,N_3878,N_4172);
nand U4985 (N_4985,N_3762,N_4483);
or U4986 (N_4986,N_3633,N_4117);
nand U4987 (N_4987,N_4734,N_4445);
nor U4988 (N_4988,N_4205,N_4618);
and U4989 (N_4989,N_4108,N_4755);
and U4990 (N_4990,N_4189,N_4019);
and U4991 (N_4991,N_4611,N_4373);
nand U4992 (N_4992,N_3732,N_4481);
xnor U4993 (N_4993,N_4459,N_4762);
or U4994 (N_4994,N_3950,N_3725);
nand U4995 (N_4995,N_3816,N_3948);
xnor U4996 (N_4996,N_4017,N_3749);
xnor U4997 (N_4997,N_4730,N_4146);
and U4998 (N_4998,N_3807,N_4187);
or U4999 (N_4999,N_4447,N_4779);
nor U5000 (N_5000,N_4698,N_4436);
nand U5001 (N_5001,N_4099,N_3935);
or U5002 (N_5002,N_3707,N_3750);
and U5003 (N_5003,N_4071,N_3907);
xor U5004 (N_5004,N_4076,N_4092);
or U5005 (N_5005,N_3718,N_3959);
nor U5006 (N_5006,N_4366,N_3912);
xnor U5007 (N_5007,N_4476,N_3927);
nor U5008 (N_5008,N_4109,N_3870);
nor U5009 (N_5009,N_4712,N_4406);
or U5010 (N_5010,N_4423,N_4644);
nor U5011 (N_5011,N_4703,N_4758);
nand U5012 (N_5012,N_4394,N_4581);
nor U5013 (N_5013,N_4165,N_3731);
or U5014 (N_5014,N_4335,N_3910);
xor U5015 (N_5015,N_4196,N_4565);
and U5016 (N_5016,N_4323,N_4159);
or U5017 (N_5017,N_4016,N_4754);
xnor U5018 (N_5018,N_4372,N_3893);
nor U5019 (N_5019,N_3688,N_4370);
nor U5020 (N_5020,N_4739,N_4249);
nand U5021 (N_5021,N_4069,N_3663);
xnor U5022 (N_5022,N_4353,N_4169);
xor U5023 (N_5023,N_4751,N_3906);
nand U5024 (N_5024,N_3783,N_3792);
xnor U5025 (N_5025,N_4256,N_4466);
nor U5026 (N_5026,N_4401,N_3701);
xnor U5027 (N_5027,N_4171,N_4513);
and U5028 (N_5028,N_4291,N_4210);
and U5029 (N_5029,N_3828,N_3868);
or U5030 (N_5030,N_4497,N_3699);
nand U5031 (N_5031,N_4038,N_3889);
or U5032 (N_5032,N_4537,N_4229);
or U5033 (N_5033,N_3676,N_4027);
nor U5034 (N_5034,N_4454,N_4226);
nand U5035 (N_5035,N_3856,N_4643);
and U5036 (N_5036,N_4340,N_3832);
or U5037 (N_5037,N_4606,N_4654);
or U5038 (N_5038,N_4706,N_4615);
xnor U5039 (N_5039,N_4679,N_4557);
nor U5040 (N_5040,N_4788,N_4585);
and U5041 (N_5041,N_4426,N_4116);
and U5042 (N_5042,N_4562,N_3968);
or U5043 (N_5043,N_4683,N_4694);
nand U5044 (N_5044,N_4744,N_4696);
and U5045 (N_5045,N_3831,N_3929);
nand U5046 (N_5046,N_3703,N_4006);
or U5047 (N_5047,N_4179,N_3892);
xnor U5048 (N_5048,N_4740,N_3788);
nor U5049 (N_5049,N_4790,N_4218);
or U5050 (N_5050,N_3997,N_4542);
or U5051 (N_5051,N_3698,N_4132);
xnor U5052 (N_5052,N_4443,N_3860);
nor U5053 (N_5053,N_3667,N_3754);
xnor U5054 (N_5054,N_3926,N_4012);
or U5055 (N_5055,N_4021,N_3952);
xnor U5056 (N_5056,N_4191,N_4270);
and U5057 (N_5057,N_4089,N_3789);
xor U5058 (N_5058,N_4258,N_4781);
nor U5059 (N_5059,N_4407,N_4110);
nand U5060 (N_5060,N_3621,N_4468);
or U5061 (N_5061,N_4621,N_4448);
or U5062 (N_5062,N_3919,N_4599);
xnor U5063 (N_5063,N_3987,N_4584);
nor U5064 (N_5064,N_3975,N_4741);
and U5065 (N_5065,N_4534,N_4126);
and U5066 (N_5066,N_4718,N_4338);
nor U5067 (N_5067,N_4084,N_4500);
nand U5068 (N_5068,N_4296,N_4772);
and U5069 (N_5069,N_3896,N_3938);
and U5070 (N_5070,N_4339,N_3810);
or U5071 (N_5071,N_4626,N_4434);
nor U5072 (N_5072,N_4732,N_3673);
nor U5073 (N_5073,N_3851,N_3880);
or U5074 (N_5074,N_4062,N_4463);
xor U5075 (N_5075,N_3822,N_4303);
nand U5076 (N_5076,N_4000,N_4595);
nand U5077 (N_5077,N_4614,N_4530);
nand U5078 (N_5078,N_4552,N_4271);
nand U5079 (N_5079,N_4263,N_4357);
and U5080 (N_5080,N_4633,N_3977);
nand U5081 (N_5081,N_4123,N_4266);
and U5082 (N_5082,N_4444,N_4657);
nor U5083 (N_5083,N_3742,N_4707);
nand U5084 (N_5084,N_3645,N_3666);
and U5085 (N_5085,N_4293,N_4355);
xnor U5086 (N_5086,N_3884,N_4243);
nand U5087 (N_5087,N_3755,N_3836);
xnor U5088 (N_5088,N_4242,N_3606);
nand U5089 (N_5089,N_3693,N_4155);
or U5090 (N_5090,N_4573,N_4056);
nor U5091 (N_5091,N_4620,N_3726);
and U5092 (N_5092,N_3834,N_4024);
xor U5093 (N_5093,N_4722,N_3752);
and U5094 (N_5094,N_4697,N_3728);
and U5095 (N_5095,N_4330,N_3909);
nor U5096 (N_5096,N_4486,N_4252);
nor U5097 (N_5097,N_4273,N_4455);
and U5098 (N_5098,N_4136,N_3655);
and U5099 (N_5099,N_4231,N_3973);
nor U5100 (N_5100,N_4656,N_4188);
xnor U5101 (N_5101,N_4622,N_3740);
or U5102 (N_5102,N_4327,N_4760);
nand U5103 (N_5103,N_3622,N_3744);
and U5104 (N_5104,N_4397,N_3823);
nand U5105 (N_5105,N_4195,N_4512);
nand U5106 (N_5106,N_4651,N_3953);
nor U5107 (N_5107,N_3958,N_3932);
xnor U5108 (N_5108,N_3675,N_4536);
xnor U5109 (N_5109,N_3824,N_4153);
nor U5110 (N_5110,N_3678,N_4131);
nor U5111 (N_5111,N_4563,N_4719);
and U5112 (N_5112,N_4380,N_4575);
or U5113 (N_5113,N_4369,N_4331);
and U5114 (N_5114,N_4178,N_4403);
or U5115 (N_5115,N_4276,N_4766);
or U5116 (N_5116,N_4647,N_4472);
or U5117 (N_5117,N_3944,N_3900);
nand U5118 (N_5118,N_3863,N_3602);
and U5119 (N_5119,N_4085,N_3888);
and U5120 (N_5120,N_4428,N_3615);
and U5121 (N_5121,N_4287,N_4569);
nand U5122 (N_5122,N_4458,N_4127);
and U5123 (N_5123,N_4405,N_3746);
nor U5124 (N_5124,N_3989,N_4013);
nor U5125 (N_5125,N_4702,N_4566);
and U5126 (N_5126,N_4031,N_4794);
nor U5127 (N_5127,N_4326,N_4655);
nor U5128 (N_5128,N_3770,N_3939);
nand U5129 (N_5129,N_3830,N_4770);
nand U5130 (N_5130,N_4723,N_4067);
nor U5131 (N_5131,N_3696,N_4043);
and U5132 (N_5132,N_4034,N_4072);
nand U5133 (N_5133,N_4743,N_3631);
nor U5134 (N_5134,N_4250,N_3614);
and U5135 (N_5135,N_4608,N_4265);
or U5136 (N_5136,N_4090,N_4499);
or U5137 (N_5137,N_4388,N_4115);
nand U5138 (N_5138,N_4460,N_4074);
and U5139 (N_5139,N_4600,N_4262);
nor U5140 (N_5140,N_3635,N_3908);
nor U5141 (N_5141,N_3780,N_4245);
or U5142 (N_5142,N_4148,N_4768);
or U5143 (N_5143,N_3761,N_4360);
and U5144 (N_5144,N_4299,N_4184);
nor U5145 (N_5145,N_3771,N_4492);
xnor U5146 (N_5146,N_4625,N_4005);
nor U5147 (N_5147,N_4073,N_4222);
and U5148 (N_5148,N_4544,N_4363);
nand U5149 (N_5149,N_4395,N_4032);
and U5150 (N_5150,N_3644,N_4147);
or U5151 (N_5151,N_4502,N_4393);
nand U5152 (N_5152,N_4098,N_4737);
nand U5153 (N_5153,N_4553,N_3982);
xor U5154 (N_5154,N_3984,N_4183);
or U5155 (N_5155,N_4300,N_3656);
nand U5156 (N_5156,N_4255,N_4785);
nand U5157 (N_5157,N_4685,N_4091);
nand U5158 (N_5158,N_3827,N_4386);
and U5159 (N_5159,N_3937,N_4383);
xor U5160 (N_5160,N_4564,N_4663);
xnor U5161 (N_5161,N_4267,N_4204);
and U5162 (N_5162,N_3642,N_4356);
or U5163 (N_5163,N_4180,N_4640);
or U5164 (N_5164,N_4796,N_4007);
or U5165 (N_5165,N_3985,N_4314);
or U5166 (N_5166,N_3902,N_4387);
and U5167 (N_5167,N_4667,N_4686);
and U5168 (N_5168,N_4548,N_3760);
nor U5169 (N_5169,N_3960,N_4491);
or U5170 (N_5170,N_3850,N_4079);
nand U5171 (N_5171,N_4010,N_4612);
or U5172 (N_5172,N_4624,N_3641);
or U5173 (N_5173,N_3692,N_4660);
xor U5174 (N_5174,N_4678,N_3691);
xor U5175 (N_5175,N_3833,N_3785);
nor U5176 (N_5176,N_3689,N_3680);
xor U5177 (N_5177,N_4634,N_4259);
xor U5178 (N_5178,N_3843,N_3829);
or U5179 (N_5179,N_3911,N_3717);
xnor U5180 (N_5180,N_4154,N_4691);
nand U5181 (N_5181,N_3715,N_3712);
nor U5182 (N_5182,N_4586,N_4442);
or U5183 (N_5183,N_4510,N_4749);
and U5184 (N_5184,N_4232,N_4151);
or U5185 (N_5185,N_3841,N_3660);
or U5186 (N_5186,N_4590,N_3964);
nand U5187 (N_5187,N_3803,N_4041);
nand U5188 (N_5188,N_4060,N_4452);
nand U5189 (N_5189,N_4518,N_3979);
xor U5190 (N_5190,N_3686,N_4628);
and U5191 (N_5191,N_3801,N_3826);
or U5192 (N_5192,N_4295,N_4042);
nand U5193 (N_5193,N_3855,N_4709);
nand U5194 (N_5194,N_4311,N_3916);
nor U5195 (N_5195,N_4623,N_3702);
or U5196 (N_5196,N_3811,N_4014);
or U5197 (N_5197,N_4619,N_4763);
or U5198 (N_5198,N_4404,N_3624);
nand U5199 (N_5199,N_3779,N_4275);
nand U5200 (N_5200,N_3778,N_4508);
nor U5201 (N_5201,N_3733,N_3873);
or U5202 (N_5202,N_4721,N_3846);
nand U5203 (N_5203,N_4780,N_3980);
nand U5204 (N_5204,N_3739,N_3808);
or U5205 (N_5205,N_4239,N_3848);
nand U5206 (N_5206,N_3773,N_4631);
xnor U5207 (N_5207,N_4125,N_4047);
nand U5208 (N_5208,N_4475,N_3634);
xor U5209 (N_5209,N_4764,N_4687);
or U5210 (N_5210,N_3898,N_3617);
nand U5211 (N_5211,N_3657,N_3735);
nor U5212 (N_5212,N_4550,N_4704);
nand U5213 (N_5213,N_3974,N_4713);
and U5214 (N_5214,N_4457,N_4144);
xor U5215 (N_5215,N_4001,N_3709);
or U5216 (N_5216,N_4247,N_4495);
nand U5217 (N_5217,N_4677,N_4029);
xor U5218 (N_5218,N_4439,N_3713);
or U5219 (N_5219,N_3640,N_4589);
nand U5220 (N_5220,N_3758,N_4106);
or U5221 (N_5221,N_4646,N_3616);
and U5222 (N_5222,N_3993,N_4738);
nor U5223 (N_5223,N_4567,N_3607);
nand U5224 (N_5224,N_4096,N_4230);
xor U5225 (N_5225,N_4545,N_4604);
and U5226 (N_5226,N_4601,N_4312);
xor U5227 (N_5227,N_4253,N_3664);
nand U5228 (N_5228,N_3837,N_3784);
nand U5229 (N_5229,N_4759,N_4149);
and U5230 (N_5230,N_3839,N_4122);
nand U5231 (N_5231,N_4450,N_4174);
xor U5232 (N_5232,N_4474,N_4103);
nand U5233 (N_5233,N_4133,N_3825);
nor U5234 (N_5234,N_3669,N_3936);
and U5235 (N_5235,N_4503,N_4617);
nand U5236 (N_5236,N_4598,N_4134);
and U5237 (N_5237,N_4748,N_4120);
and U5238 (N_5238,N_4539,N_3920);
nor U5239 (N_5239,N_4050,N_4577);
and U5240 (N_5240,N_4057,N_4367);
xnor U5241 (N_5241,N_3639,N_4307);
xor U5242 (N_5242,N_4298,N_4348);
nor U5243 (N_5243,N_3738,N_4636);
xor U5244 (N_5244,N_4609,N_4467);
and U5245 (N_5245,N_4297,N_4313);
xnor U5246 (N_5246,N_4639,N_3649);
and U5247 (N_5247,N_4453,N_4105);
nor U5248 (N_5248,N_4077,N_3869);
nor U5249 (N_5249,N_3814,N_4176);
nand U5250 (N_5250,N_4135,N_4396);
or U5251 (N_5251,N_4342,N_4282);
nand U5252 (N_5252,N_3924,N_4753);
nor U5253 (N_5253,N_4587,N_3849);
xor U5254 (N_5254,N_4234,N_3861);
nand U5255 (N_5255,N_3711,N_4280);
or U5256 (N_5256,N_4490,N_4371);
nand U5257 (N_5257,N_3940,N_4305);
nor U5258 (N_5258,N_3838,N_4227);
xor U5259 (N_5259,N_4593,N_3782);
or U5260 (N_5260,N_3729,N_4729);
nand U5261 (N_5261,N_4365,N_3905);
and U5262 (N_5262,N_3710,N_4164);
or U5263 (N_5263,N_3734,N_4509);
or U5264 (N_5264,N_3931,N_4519);
and U5265 (N_5265,N_4430,N_4479);
nand U5266 (N_5266,N_4039,N_4789);
xnor U5267 (N_5267,N_3618,N_3881);
nor U5268 (N_5268,N_4673,N_4591);
nor U5269 (N_5269,N_4220,N_3922);
nand U5270 (N_5270,N_4170,N_4736);
nor U5271 (N_5271,N_4710,N_4045);
nor U5272 (N_5272,N_3835,N_3737);
nor U5273 (N_5273,N_4378,N_4376);
or U5274 (N_5274,N_3747,N_3774);
or U5275 (N_5275,N_4670,N_4653);
or U5276 (N_5276,N_4061,N_3820);
and U5277 (N_5277,N_4302,N_3934);
xnor U5278 (N_5278,N_3765,N_3751);
nor U5279 (N_5279,N_4139,N_3815);
nor U5280 (N_5280,N_4107,N_4554);
nand U5281 (N_5281,N_3928,N_3995);
and U5282 (N_5282,N_3790,N_4570);
or U5283 (N_5283,N_3904,N_4100);
nand U5284 (N_5284,N_4328,N_3682);
or U5285 (N_5285,N_4003,N_4559);
nand U5286 (N_5286,N_4221,N_4756);
and U5287 (N_5287,N_4422,N_4173);
nor U5288 (N_5288,N_3681,N_3930);
xnor U5289 (N_5289,N_4199,N_4720);
and U5290 (N_5290,N_4786,N_4574);
nor U5291 (N_5291,N_4018,N_3805);
and U5292 (N_5292,N_4416,N_3969);
and U5293 (N_5293,N_3767,N_4733);
or U5294 (N_5294,N_3620,N_4237);
and U5295 (N_5295,N_4588,N_4156);
xnor U5296 (N_5296,N_3887,N_3992);
or U5297 (N_5297,N_4362,N_3840);
and U5298 (N_5298,N_3662,N_4036);
xnor U5299 (N_5299,N_4791,N_4181);
nor U5300 (N_5300,N_4725,N_4752);
and U5301 (N_5301,N_3741,N_3627);
or U5302 (N_5302,N_3800,N_4379);
nand U5303 (N_5303,N_4597,N_4130);
and U5304 (N_5304,N_4333,N_4306);
or U5305 (N_5305,N_4413,N_3913);
xnor U5306 (N_5306,N_4175,N_4529);
nor U5307 (N_5307,N_4798,N_4201);
xnor U5308 (N_5308,N_4773,N_4549);
and U5309 (N_5309,N_4547,N_4551);
nand U5310 (N_5310,N_4286,N_3955);
or U5311 (N_5311,N_3853,N_4596);
nand U5312 (N_5312,N_4572,N_4543);
xnor U5313 (N_5313,N_3638,N_4750);
xor U5314 (N_5314,N_3719,N_4070);
and U5315 (N_5315,N_4681,N_4715);
nor U5316 (N_5316,N_4068,N_4269);
nor U5317 (N_5317,N_4319,N_4345);
nand U5318 (N_5318,N_3999,N_4478);
and U5319 (N_5319,N_3671,N_4185);
nand U5320 (N_5320,N_4385,N_4213);
and U5321 (N_5321,N_4211,N_4701);
nand U5322 (N_5322,N_4571,N_3965);
nor U5323 (N_5323,N_3608,N_3768);
or U5324 (N_5324,N_3859,N_4507);
and U5325 (N_5325,N_4501,N_4277);
xnor U5326 (N_5326,N_4248,N_4002);
xnor U5327 (N_5327,N_4145,N_3821);
xnor U5328 (N_5328,N_4797,N_4505);
nand U5329 (N_5329,N_3890,N_4217);
or U5330 (N_5330,N_4279,N_4451);
nor U5331 (N_5331,N_3866,N_4294);
nor U5332 (N_5332,N_3791,N_4613);
nor U5333 (N_5333,N_4389,N_4777);
and U5334 (N_5334,N_4142,N_4627);
or U5335 (N_5335,N_4101,N_3897);
xor U5336 (N_5336,N_4799,N_3956);
or U5337 (N_5337,N_4616,N_4514);
nand U5338 (N_5338,N_4113,N_4037);
or U5339 (N_5339,N_4064,N_4778);
and U5340 (N_5340,N_4177,N_3921);
or U5341 (N_5341,N_3611,N_4437);
xor U5342 (N_5342,N_4341,N_3705);
xnor U5343 (N_5343,N_4368,N_3708);
xor U5344 (N_5344,N_4425,N_4390);
nand U5345 (N_5345,N_4517,N_4223);
nor U5346 (N_5346,N_4254,N_4446);
or U5347 (N_5347,N_4645,N_3687);
nand U5348 (N_5348,N_4111,N_4708);
nand U5349 (N_5349,N_4138,N_4493);
nand U5350 (N_5350,N_3957,N_4285);
nor U5351 (N_5351,N_4409,N_4163);
xor U5352 (N_5352,N_3967,N_4040);
xor U5353 (N_5353,N_4765,N_3690);
or U5354 (N_5354,N_3797,N_4658);
nand U5355 (N_5355,N_4352,N_4761);
or U5356 (N_5356,N_4669,N_3867);
nor U5357 (N_5357,N_3899,N_3845);
nor U5358 (N_5358,N_3652,N_3665);
xor U5359 (N_5359,N_4746,N_3781);
or U5360 (N_5360,N_4063,N_3720);
nor U5361 (N_5361,N_3879,N_4137);
nor U5362 (N_5362,N_3722,N_3604);
nor U5363 (N_5363,N_4225,N_4578);
or U5364 (N_5364,N_3677,N_4212);
nand U5365 (N_5365,N_4304,N_3776);
and U5366 (N_5366,N_4470,N_4198);
and U5367 (N_5367,N_3745,N_3623);
and U5368 (N_5368,N_4015,N_3852);
nor U5369 (N_5369,N_4241,N_3991);
and U5370 (N_5370,N_4251,N_3962);
xnor U5371 (N_5371,N_4747,N_4087);
xnor U5372 (N_5372,N_4757,N_4344);
nor U5373 (N_5373,N_4197,N_4093);
nor U5374 (N_5374,N_3802,N_4771);
nand U5375 (N_5375,N_4272,N_3983);
xnor U5376 (N_5376,N_4097,N_4675);
nor U5377 (N_5377,N_4641,N_4377);
xor U5378 (N_5378,N_4121,N_4525);
or U5379 (N_5379,N_4783,N_4081);
nor U5380 (N_5380,N_4469,N_4240);
nand U5381 (N_5381,N_4382,N_4020);
xnor U5382 (N_5382,N_4051,N_3903);
nor U5383 (N_5383,N_4186,N_4278);
or U5384 (N_5384,N_3875,N_4347);
xor U5385 (N_5385,N_4724,N_3854);
and U5386 (N_5386,N_4473,N_3704);
or U5387 (N_5387,N_4246,N_4649);
and U5388 (N_5388,N_4119,N_4095);
xor U5389 (N_5389,N_3990,N_3799);
or U5390 (N_5390,N_3817,N_3862);
nor U5391 (N_5391,N_4775,N_4257);
nand U5392 (N_5392,N_4535,N_4374);
xor U5393 (N_5393,N_4471,N_4676);
and U5394 (N_5394,N_4583,N_4540);
or U5395 (N_5395,N_3901,N_4028);
nand U5396 (N_5396,N_4349,N_3813);
or U5397 (N_5397,N_4784,N_4494);
nand U5398 (N_5398,N_3883,N_4083);
xor U5399 (N_5399,N_4182,N_3942);
xnor U5400 (N_5400,N_3873,N_4051);
nor U5401 (N_5401,N_3972,N_4728);
nand U5402 (N_5402,N_3921,N_4752);
and U5403 (N_5403,N_4016,N_4546);
xor U5404 (N_5404,N_4178,N_4671);
xor U5405 (N_5405,N_4484,N_4346);
and U5406 (N_5406,N_3699,N_3926);
or U5407 (N_5407,N_4003,N_4157);
and U5408 (N_5408,N_4104,N_4620);
or U5409 (N_5409,N_4706,N_3919);
nor U5410 (N_5410,N_4349,N_4154);
nand U5411 (N_5411,N_4797,N_4711);
nor U5412 (N_5412,N_3723,N_4293);
and U5413 (N_5413,N_4291,N_3721);
nor U5414 (N_5414,N_4297,N_3907);
nand U5415 (N_5415,N_4387,N_4357);
and U5416 (N_5416,N_3934,N_4551);
or U5417 (N_5417,N_4091,N_3838);
xnor U5418 (N_5418,N_4246,N_3818);
or U5419 (N_5419,N_4230,N_4692);
or U5420 (N_5420,N_3815,N_3640);
nor U5421 (N_5421,N_3898,N_3815);
or U5422 (N_5422,N_3688,N_4066);
nand U5423 (N_5423,N_4005,N_4667);
nand U5424 (N_5424,N_4361,N_3635);
and U5425 (N_5425,N_4181,N_4379);
xor U5426 (N_5426,N_4783,N_4744);
xnor U5427 (N_5427,N_3874,N_4616);
nor U5428 (N_5428,N_3829,N_4555);
xnor U5429 (N_5429,N_4674,N_3630);
nor U5430 (N_5430,N_3689,N_3644);
xnor U5431 (N_5431,N_4018,N_3712);
nand U5432 (N_5432,N_3843,N_4238);
nand U5433 (N_5433,N_4415,N_4177);
xnor U5434 (N_5434,N_4724,N_4172);
xnor U5435 (N_5435,N_4571,N_3701);
or U5436 (N_5436,N_4107,N_4655);
nor U5437 (N_5437,N_4397,N_3785);
xnor U5438 (N_5438,N_4555,N_3920);
and U5439 (N_5439,N_4506,N_4186);
nand U5440 (N_5440,N_3837,N_4517);
and U5441 (N_5441,N_3893,N_4715);
xnor U5442 (N_5442,N_4450,N_4682);
and U5443 (N_5443,N_3794,N_3845);
nand U5444 (N_5444,N_4243,N_4722);
nand U5445 (N_5445,N_4487,N_4412);
and U5446 (N_5446,N_4041,N_3955);
and U5447 (N_5447,N_4721,N_4016);
or U5448 (N_5448,N_3889,N_4467);
nor U5449 (N_5449,N_3662,N_3900);
nand U5450 (N_5450,N_3922,N_4573);
xor U5451 (N_5451,N_3947,N_3730);
or U5452 (N_5452,N_4131,N_4446);
xor U5453 (N_5453,N_3871,N_3623);
nor U5454 (N_5454,N_4373,N_4164);
or U5455 (N_5455,N_3824,N_3852);
or U5456 (N_5456,N_4789,N_4322);
or U5457 (N_5457,N_4595,N_3710);
xor U5458 (N_5458,N_4039,N_3772);
nor U5459 (N_5459,N_4348,N_3669);
and U5460 (N_5460,N_4070,N_4336);
and U5461 (N_5461,N_3677,N_3854);
xnor U5462 (N_5462,N_4706,N_4702);
xnor U5463 (N_5463,N_3713,N_4446);
or U5464 (N_5464,N_3621,N_4754);
or U5465 (N_5465,N_3690,N_4705);
or U5466 (N_5466,N_4369,N_4711);
xor U5467 (N_5467,N_4379,N_4638);
xnor U5468 (N_5468,N_3660,N_3721);
nand U5469 (N_5469,N_3802,N_4230);
nand U5470 (N_5470,N_3665,N_4199);
nand U5471 (N_5471,N_4230,N_4455);
or U5472 (N_5472,N_4703,N_4593);
and U5473 (N_5473,N_4168,N_4471);
nor U5474 (N_5474,N_4560,N_4773);
nand U5475 (N_5475,N_4313,N_4503);
nor U5476 (N_5476,N_4704,N_4775);
nand U5477 (N_5477,N_3775,N_4444);
or U5478 (N_5478,N_4133,N_3925);
xnor U5479 (N_5479,N_4193,N_3785);
xnor U5480 (N_5480,N_4273,N_4014);
nand U5481 (N_5481,N_3836,N_4745);
nor U5482 (N_5482,N_3764,N_4195);
nand U5483 (N_5483,N_4636,N_3824);
xnor U5484 (N_5484,N_4250,N_3792);
or U5485 (N_5485,N_4218,N_3669);
xnor U5486 (N_5486,N_4776,N_4676);
xor U5487 (N_5487,N_4654,N_3929);
nor U5488 (N_5488,N_4738,N_3913);
nor U5489 (N_5489,N_3682,N_4598);
or U5490 (N_5490,N_3624,N_3763);
nor U5491 (N_5491,N_3888,N_3707);
xnor U5492 (N_5492,N_4630,N_4372);
nor U5493 (N_5493,N_3651,N_3769);
and U5494 (N_5494,N_3944,N_4438);
nand U5495 (N_5495,N_4008,N_4215);
or U5496 (N_5496,N_4606,N_4518);
or U5497 (N_5497,N_4612,N_3974);
or U5498 (N_5498,N_4248,N_3606);
nand U5499 (N_5499,N_4338,N_4225);
or U5500 (N_5500,N_4087,N_4024);
and U5501 (N_5501,N_3659,N_4236);
xor U5502 (N_5502,N_4183,N_4059);
xor U5503 (N_5503,N_4209,N_4694);
xor U5504 (N_5504,N_4283,N_4109);
xnor U5505 (N_5505,N_3778,N_4641);
or U5506 (N_5506,N_3956,N_3672);
xnor U5507 (N_5507,N_4198,N_3859);
nand U5508 (N_5508,N_4396,N_4051);
nand U5509 (N_5509,N_3924,N_3887);
nand U5510 (N_5510,N_4357,N_4133);
nand U5511 (N_5511,N_4342,N_3663);
and U5512 (N_5512,N_3858,N_3935);
nor U5513 (N_5513,N_3865,N_4261);
xnor U5514 (N_5514,N_3818,N_4471);
or U5515 (N_5515,N_3995,N_4334);
nor U5516 (N_5516,N_4462,N_3676);
nand U5517 (N_5517,N_3603,N_4156);
xor U5518 (N_5518,N_3944,N_4704);
nand U5519 (N_5519,N_3976,N_4408);
nand U5520 (N_5520,N_4302,N_4729);
and U5521 (N_5521,N_3857,N_4053);
or U5522 (N_5522,N_4135,N_4533);
nand U5523 (N_5523,N_4260,N_4363);
or U5524 (N_5524,N_3964,N_4568);
nand U5525 (N_5525,N_4266,N_4524);
xnor U5526 (N_5526,N_4698,N_3754);
nand U5527 (N_5527,N_4398,N_4571);
or U5528 (N_5528,N_3926,N_4034);
nand U5529 (N_5529,N_4766,N_4109);
or U5530 (N_5530,N_3804,N_4746);
nand U5531 (N_5531,N_4719,N_4758);
or U5532 (N_5532,N_4778,N_4722);
nor U5533 (N_5533,N_4377,N_3916);
nand U5534 (N_5534,N_4452,N_4755);
xnor U5535 (N_5535,N_3857,N_4601);
nand U5536 (N_5536,N_4399,N_4076);
and U5537 (N_5537,N_3950,N_4547);
nor U5538 (N_5538,N_4537,N_4251);
xnor U5539 (N_5539,N_3906,N_4482);
nor U5540 (N_5540,N_4364,N_4045);
xor U5541 (N_5541,N_4057,N_4461);
and U5542 (N_5542,N_3630,N_4295);
or U5543 (N_5543,N_4511,N_4393);
or U5544 (N_5544,N_3886,N_4669);
and U5545 (N_5545,N_4343,N_3919);
or U5546 (N_5546,N_4766,N_3739);
and U5547 (N_5547,N_3932,N_3866);
and U5548 (N_5548,N_4739,N_3621);
or U5549 (N_5549,N_3847,N_4790);
xnor U5550 (N_5550,N_3985,N_3691);
and U5551 (N_5551,N_3671,N_3732);
xnor U5552 (N_5552,N_3619,N_4009);
nand U5553 (N_5553,N_4310,N_3920);
or U5554 (N_5554,N_4620,N_4641);
xnor U5555 (N_5555,N_4418,N_4376);
and U5556 (N_5556,N_3999,N_4022);
nor U5557 (N_5557,N_4551,N_3974);
and U5558 (N_5558,N_4543,N_3754);
nand U5559 (N_5559,N_4179,N_4189);
nor U5560 (N_5560,N_3886,N_4070);
and U5561 (N_5561,N_4213,N_4750);
nor U5562 (N_5562,N_4266,N_3973);
or U5563 (N_5563,N_4097,N_4118);
nor U5564 (N_5564,N_4119,N_3913);
nand U5565 (N_5565,N_3780,N_3815);
or U5566 (N_5566,N_4637,N_4491);
nand U5567 (N_5567,N_4755,N_3796);
and U5568 (N_5568,N_4423,N_4290);
and U5569 (N_5569,N_4227,N_4771);
nor U5570 (N_5570,N_4076,N_4400);
nand U5571 (N_5571,N_3718,N_4126);
xnor U5572 (N_5572,N_4116,N_4324);
xnor U5573 (N_5573,N_3880,N_4327);
nand U5574 (N_5574,N_4657,N_4755);
and U5575 (N_5575,N_4733,N_3680);
xnor U5576 (N_5576,N_3602,N_4618);
xor U5577 (N_5577,N_3751,N_4165);
nand U5578 (N_5578,N_4728,N_4659);
or U5579 (N_5579,N_4056,N_4160);
nand U5580 (N_5580,N_4008,N_4520);
or U5581 (N_5581,N_4097,N_4419);
nand U5582 (N_5582,N_4156,N_3755);
xnor U5583 (N_5583,N_3773,N_4621);
or U5584 (N_5584,N_4404,N_3654);
nor U5585 (N_5585,N_4110,N_3867);
or U5586 (N_5586,N_4731,N_4633);
nor U5587 (N_5587,N_4613,N_3786);
xor U5588 (N_5588,N_4477,N_4204);
xor U5589 (N_5589,N_4460,N_3988);
nor U5590 (N_5590,N_4016,N_4455);
and U5591 (N_5591,N_4207,N_3844);
xnor U5592 (N_5592,N_4758,N_3975);
or U5593 (N_5593,N_4418,N_4041);
nand U5594 (N_5594,N_4052,N_4654);
xor U5595 (N_5595,N_3929,N_4102);
nor U5596 (N_5596,N_3650,N_4397);
nand U5597 (N_5597,N_3694,N_4675);
nor U5598 (N_5598,N_4003,N_3870);
and U5599 (N_5599,N_4191,N_3770);
and U5600 (N_5600,N_3836,N_4418);
xor U5601 (N_5601,N_4680,N_4765);
nand U5602 (N_5602,N_4631,N_4063);
and U5603 (N_5603,N_4193,N_4086);
nand U5604 (N_5604,N_4755,N_4367);
nor U5605 (N_5605,N_4474,N_3642);
xor U5606 (N_5606,N_3732,N_4218);
or U5607 (N_5607,N_4610,N_4708);
nand U5608 (N_5608,N_3770,N_3860);
nand U5609 (N_5609,N_3989,N_3800);
and U5610 (N_5610,N_3692,N_3950);
nand U5611 (N_5611,N_3823,N_4136);
and U5612 (N_5612,N_4792,N_4206);
nor U5613 (N_5613,N_3693,N_4568);
and U5614 (N_5614,N_3760,N_3934);
nor U5615 (N_5615,N_4774,N_3924);
xnor U5616 (N_5616,N_4216,N_3608);
nor U5617 (N_5617,N_4757,N_4018);
and U5618 (N_5618,N_3755,N_4335);
and U5619 (N_5619,N_4603,N_4121);
xor U5620 (N_5620,N_3611,N_3722);
and U5621 (N_5621,N_4548,N_3917);
xor U5622 (N_5622,N_4630,N_4509);
xnor U5623 (N_5623,N_4306,N_3741);
xor U5624 (N_5624,N_4141,N_4331);
and U5625 (N_5625,N_4727,N_4491);
nand U5626 (N_5626,N_4231,N_4474);
nand U5627 (N_5627,N_4584,N_3632);
xnor U5628 (N_5628,N_4512,N_3712);
and U5629 (N_5629,N_4567,N_3903);
nand U5630 (N_5630,N_4656,N_4500);
nor U5631 (N_5631,N_3833,N_4544);
nor U5632 (N_5632,N_4602,N_3721);
xor U5633 (N_5633,N_3613,N_4353);
nor U5634 (N_5634,N_3767,N_4341);
or U5635 (N_5635,N_4043,N_4334);
nor U5636 (N_5636,N_3949,N_4054);
or U5637 (N_5637,N_4151,N_3811);
nor U5638 (N_5638,N_4056,N_4734);
xnor U5639 (N_5639,N_4699,N_4496);
nand U5640 (N_5640,N_4551,N_4665);
nor U5641 (N_5641,N_4277,N_3915);
and U5642 (N_5642,N_4731,N_4116);
or U5643 (N_5643,N_4028,N_4783);
and U5644 (N_5644,N_4696,N_4344);
and U5645 (N_5645,N_3995,N_3958);
nand U5646 (N_5646,N_4471,N_3624);
nor U5647 (N_5647,N_4678,N_4293);
and U5648 (N_5648,N_3711,N_4119);
nor U5649 (N_5649,N_4529,N_4237);
xor U5650 (N_5650,N_4281,N_3795);
nand U5651 (N_5651,N_4038,N_4755);
and U5652 (N_5652,N_3986,N_4790);
and U5653 (N_5653,N_4219,N_3958);
nor U5654 (N_5654,N_4456,N_3845);
and U5655 (N_5655,N_4039,N_4643);
nand U5656 (N_5656,N_4483,N_4381);
and U5657 (N_5657,N_4080,N_4129);
xnor U5658 (N_5658,N_4105,N_4605);
or U5659 (N_5659,N_4386,N_4472);
and U5660 (N_5660,N_4158,N_4208);
nand U5661 (N_5661,N_4053,N_3968);
nor U5662 (N_5662,N_4084,N_4630);
nor U5663 (N_5663,N_3885,N_4454);
or U5664 (N_5664,N_3842,N_4022);
or U5665 (N_5665,N_4596,N_4110);
and U5666 (N_5666,N_3861,N_3609);
xor U5667 (N_5667,N_3759,N_3718);
or U5668 (N_5668,N_4423,N_3896);
and U5669 (N_5669,N_3761,N_4214);
xnor U5670 (N_5670,N_4082,N_3824);
xnor U5671 (N_5671,N_4580,N_4525);
xor U5672 (N_5672,N_4177,N_4710);
or U5673 (N_5673,N_3624,N_3650);
nand U5674 (N_5674,N_3931,N_4099);
and U5675 (N_5675,N_4243,N_4359);
nor U5676 (N_5676,N_4403,N_3881);
nand U5677 (N_5677,N_4443,N_3761);
nand U5678 (N_5678,N_4320,N_4375);
nor U5679 (N_5679,N_3627,N_3759);
nor U5680 (N_5680,N_4605,N_4484);
or U5681 (N_5681,N_4548,N_4507);
nor U5682 (N_5682,N_4679,N_3806);
and U5683 (N_5683,N_4635,N_3685);
nor U5684 (N_5684,N_4615,N_4323);
nor U5685 (N_5685,N_4716,N_3895);
xnor U5686 (N_5686,N_4565,N_3660);
or U5687 (N_5687,N_4772,N_4596);
or U5688 (N_5688,N_4224,N_4345);
nand U5689 (N_5689,N_4202,N_4115);
or U5690 (N_5690,N_4494,N_4773);
nor U5691 (N_5691,N_4390,N_4705);
nand U5692 (N_5692,N_4059,N_3997);
and U5693 (N_5693,N_3748,N_4180);
and U5694 (N_5694,N_4371,N_4688);
nand U5695 (N_5695,N_3737,N_3603);
and U5696 (N_5696,N_4771,N_3676);
xnor U5697 (N_5697,N_4082,N_4642);
nor U5698 (N_5698,N_4030,N_4289);
and U5699 (N_5699,N_4380,N_4736);
xor U5700 (N_5700,N_4332,N_4728);
or U5701 (N_5701,N_4157,N_4042);
nor U5702 (N_5702,N_4744,N_4328);
or U5703 (N_5703,N_4180,N_4294);
and U5704 (N_5704,N_4335,N_4694);
xor U5705 (N_5705,N_4343,N_4182);
and U5706 (N_5706,N_4076,N_4340);
or U5707 (N_5707,N_4481,N_4562);
nand U5708 (N_5708,N_3850,N_3989);
nand U5709 (N_5709,N_4109,N_3641);
xnor U5710 (N_5710,N_3942,N_4291);
and U5711 (N_5711,N_3811,N_4067);
xor U5712 (N_5712,N_4650,N_4647);
nand U5713 (N_5713,N_3780,N_4365);
xor U5714 (N_5714,N_3763,N_3818);
nand U5715 (N_5715,N_3859,N_4098);
nor U5716 (N_5716,N_4009,N_4472);
xnor U5717 (N_5717,N_4472,N_3927);
xor U5718 (N_5718,N_3735,N_4283);
nand U5719 (N_5719,N_4290,N_3651);
and U5720 (N_5720,N_4465,N_3688);
xnor U5721 (N_5721,N_4159,N_4098);
and U5722 (N_5722,N_3670,N_3716);
xnor U5723 (N_5723,N_3979,N_4354);
nand U5724 (N_5724,N_4289,N_4200);
xor U5725 (N_5725,N_4575,N_3718);
and U5726 (N_5726,N_4098,N_4538);
and U5727 (N_5727,N_3769,N_3716);
xnor U5728 (N_5728,N_4510,N_4431);
nor U5729 (N_5729,N_4498,N_3663);
and U5730 (N_5730,N_4698,N_4528);
nand U5731 (N_5731,N_3857,N_3626);
nor U5732 (N_5732,N_4521,N_4366);
and U5733 (N_5733,N_3945,N_3901);
nand U5734 (N_5734,N_4052,N_4084);
nor U5735 (N_5735,N_4413,N_4655);
nand U5736 (N_5736,N_3954,N_4308);
nand U5737 (N_5737,N_4109,N_4440);
or U5738 (N_5738,N_4152,N_4340);
nor U5739 (N_5739,N_3800,N_4009);
nor U5740 (N_5740,N_3717,N_3790);
nor U5741 (N_5741,N_4455,N_3697);
xnor U5742 (N_5742,N_3704,N_4423);
xor U5743 (N_5743,N_3939,N_3816);
or U5744 (N_5744,N_3903,N_4421);
xor U5745 (N_5745,N_3757,N_4652);
nand U5746 (N_5746,N_4355,N_4486);
nand U5747 (N_5747,N_4233,N_3741);
and U5748 (N_5748,N_3668,N_3863);
and U5749 (N_5749,N_3833,N_4272);
nand U5750 (N_5750,N_4452,N_3940);
nor U5751 (N_5751,N_3855,N_4355);
nor U5752 (N_5752,N_4376,N_3748);
or U5753 (N_5753,N_4599,N_3891);
xor U5754 (N_5754,N_3653,N_3793);
nor U5755 (N_5755,N_3738,N_3713);
nand U5756 (N_5756,N_4421,N_3946);
nor U5757 (N_5757,N_4279,N_3811);
nand U5758 (N_5758,N_4405,N_4170);
nor U5759 (N_5759,N_4200,N_4479);
or U5760 (N_5760,N_3799,N_3850);
nor U5761 (N_5761,N_4070,N_4073);
xor U5762 (N_5762,N_4164,N_4324);
and U5763 (N_5763,N_3813,N_3858);
xor U5764 (N_5764,N_4543,N_4531);
xor U5765 (N_5765,N_4639,N_4727);
and U5766 (N_5766,N_4041,N_3713);
xnor U5767 (N_5767,N_4781,N_4548);
xnor U5768 (N_5768,N_4139,N_4615);
or U5769 (N_5769,N_4254,N_4406);
xor U5770 (N_5770,N_3984,N_4335);
nor U5771 (N_5771,N_4166,N_4460);
nand U5772 (N_5772,N_3816,N_4004);
nand U5773 (N_5773,N_4745,N_4061);
and U5774 (N_5774,N_4384,N_3782);
and U5775 (N_5775,N_3663,N_4565);
xor U5776 (N_5776,N_3695,N_3859);
or U5777 (N_5777,N_3851,N_3680);
nand U5778 (N_5778,N_4683,N_3658);
nand U5779 (N_5779,N_3774,N_3845);
xor U5780 (N_5780,N_4003,N_4604);
or U5781 (N_5781,N_4182,N_4680);
xnor U5782 (N_5782,N_4235,N_4119);
nand U5783 (N_5783,N_4263,N_4280);
or U5784 (N_5784,N_4177,N_4692);
and U5785 (N_5785,N_3977,N_3633);
or U5786 (N_5786,N_3790,N_4550);
nand U5787 (N_5787,N_4516,N_4164);
and U5788 (N_5788,N_4587,N_4698);
or U5789 (N_5789,N_3714,N_4183);
or U5790 (N_5790,N_4050,N_4047);
and U5791 (N_5791,N_4464,N_4262);
xor U5792 (N_5792,N_3710,N_4046);
nand U5793 (N_5793,N_4544,N_3638);
nand U5794 (N_5794,N_4195,N_3879);
nand U5795 (N_5795,N_4509,N_4104);
xnor U5796 (N_5796,N_4390,N_3973);
or U5797 (N_5797,N_3857,N_4709);
nor U5798 (N_5798,N_3944,N_3796);
nand U5799 (N_5799,N_4638,N_4223);
and U5800 (N_5800,N_4637,N_3611);
and U5801 (N_5801,N_4230,N_4519);
or U5802 (N_5802,N_4593,N_4558);
nand U5803 (N_5803,N_4491,N_4552);
and U5804 (N_5804,N_4688,N_4608);
nand U5805 (N_5805,N_4714,N_4239);
xnor U5806 (N_5806,N_3693,N_4146);
nor U5807 (N_5807,N_4242,N_4354);
and U5808 (N_5808,N_3882,N_4041);
nor U5809 (N_5809,N_3703,N_4685);
or U5810 (N_5810,N_4564,N_4683);
or U5811 (N_5811,N_4356,N_3735);
and U5812 (N_5812,N_4459,N_3773);
nor U5813 (N_5813,N_3847,N_4731);
nor U5814 (N_5814,N_4254,N_4036);
nand U5815 (N_5815,N_3678,N_3794);
nand U5816 (N_5816,N_3924,N_4330);
or U5817 (N_5817,N_4574,N_4022);
xor U5818 (N_5818,N_3917,N_4528);
and U5819 (N_5819,N_3616,N_3996);
xnor U5820 (N_5820,N_4105,N_3800);
or U5821 (N_5821,N_4292,N_3971);
nor U5822 (N_5822,N_3939,N_4333);
xor U5823 (N_5823,N_4239,N_4058);
nor U5824 (N_5824,N_4651,N_3701);
nor U5825 (N_5825,N_3878,N_4522);
nor U5826 (N_5826,N_4033,N_4054);
and U5827 (N_5827,N_4220,N_4140);
xnor U5828 (N_5828,N_3893,N_4663);
and U5829 (N_5829,N_4243,N_3959);
xor U5830 (N_5830,N_4723,N_4554);
or U5831 (N_5831,N_4542,N_4409);
and U5832 (N_5832,N_4321,N_3730);
or U5833 (N_5833,N_3764,N_3868);
and U5834 (N_5834,N_3666,N_4381);
or U5835 (N_5835,N_4179,N_4705);
or U5836 (N_5836,N_3845,N_4445);
or U5837 (N_5837,N_4692,N_4502);
nand U5838 (N_5838,N_4744,N_3762);
nor U5839 (N_5839,N_4641,N_4155);
xnor U5840 (N_5840,N_3895,N_4159);
and U5841 (N_5841,N_4418,N_3732);
xnor U5842 (N_5842,N_3756,N_4749);
xor U5843 (N_5843,N_4620,N_4566);
nor U5844 (N_5844,N_4168,N_4650);
nand U5845 (N_5845,N_3955,N_4015);
nand U5846 (N_5846,N_3945,N_4705);
xnor U5847 (N_5847,N_3866,N_4142);
nand U5848 (N_5848,N_4008,N_4205);
xor U5849 (N_5849,N_4314,N_3840);
or U5850 (N_5850,N_4635,N_3840);
nor U5851 (N_5851,N_3925,N_3807);
or U5852 (N_5852,N_4219,N_3699);
xor U5853 (N_5853,N_4560,N_4112);
and U5854 (N_5854,N_4230,N_3916);
nor U5855 (N_5855,N_4370,N_4794);
nor U5856 (N_5856,N_4336,N_3895);
nor U5857 (N_5857,N_4446,N_3931);
nor U5858 (N_5858,N_3713,N_4702);
nor U5859 (N_5859,N_4703,N_4475);
xor U5860 (N_5860,N_4346,N_4500);
and U5861 (N_5861,N_4234,N_3863);
or U5862 (N_5862,N_3781,N_3858);
xor U5863 (N_5863,N_3652,N_4473);
xnor U5864 (N_5864,N_4692,N_3671);
or U5865 (N_5865,N_4601,N_4294);
xnor U5866 (N_5866,N_3723,N_4077);
nor U5867 (N_5867,N_4651,N_4487);
nor U5868 (N_5868,N_4620,N_4285);
nor U5869 (N_5869,N_4645,N_4724);
nor U5870 (N_5870,N_4155,N_3723);
or U5871 (N_5871,N_3685,N_4333);
nand U5872 (N_5872,N_4444,N_4208);
or U5873 (N_5873,N_4407,N_4243);
and U5874 (N_5874,N_4722,N_4659);
nor U5875 (N_5875,N_4667,N_3623);
nand U5876 (N_5876,N_3665,N_4267);
nand U5877 (N_5877,N_4604,N_4311);
xor U5878 (N_5878,N_4247,N_3984);
or U5879 (N_5879,N_4723,N_3966);
xnor U5880 (N_5880,N_4465,N_4265);
nor U5881 (N_5881,N_4679,N_4486);
nand U5882 (N_5882,N_4011,N_4151);
nor U5883 (N_5883,N_4381,N_4792);
xor U5884 (N_5884,N_4242,N_3832);
and U5885 (N_5885,N_4175,N_4428);
and U5886 (N_5886,N_4437,N_3809);
xnor U5887 (N_5887,N_4340,N_4329);
nand U5888 (N_5888,N_4285,N_3697);
and U5889 (N_5889,N_4641,N_4686);
nor U5890 (N_5890,N_4554,N_4775);
xnor U5891 (N_5891,N_4605,N_4163);
or U5892 (N_5892,N_4727,N_4092);
nor U5893 (N_5893,N_4579,N_4675);
xnor U5894 (N_5894,N_4750,N_4234);
nor U5895 (N_5895,N_4683,N_3969);
nand U5896 (N_5896,N_4504,N_3642);
or U5897 (N_5897,N_4127,N_4199);
nand U5898 (N_5898,N_4402,N_3714);
xor U5899 (N_5899,N_3770,N_3715);
nand U5900 (N_5900,N_4262,N_3616);
and U5901 (N_5901,N_4705,N_4021);
or U5902 (N_5902,N_3842,N_3619);
or U5903 (N_5903,N_4530,N_4406);
and U5904 (N_5904,N_4600,N_4320);
nor U5905 (N_5905,N_4567,N_4536);
and U5906 (N_5906,N_3830,N_3702);
and U5907 (N_5907,N_3832,N_4748);
nand U5908 (N_5908,N_4770,N_4134);
or U5909 (N_5909,N_4136,N_4667);
and U5910 (N_5910,N_3974,N_4390);
nand U5911 (N_5911,N_4286,N_4544);
nand U5912 (N_5912,N_4781,N_4525);
and U5913 (N_5913,N_4386,N_4659);
and U5914 (N_5914,N_3661,N_3812);
nand U5915 (N_5915,N_4628,N_4123);
and U5916 (N_5916,N_4540,N_4044);
nor U5917 (N_5917,N_4517,N_4586);
and U5918 (N_5918,N_3840,N_4000);
nand U5919 (N_5919,N_3695,N_3628);
and U5920 (N_5920,N_3607,N_4014);
nand U5921 (N_5921,N_3618,N_3622);
xnor U5922 (N_5922,N_4243,N_3749);
nand U5923 (N_5923,N_4057,N_4347);
xor U5924 (N_5924,N_4084,N_4197);
and U5925 (N_5925,N_3794,N_4250);
nand U5926 (N_5926,N_4748,N_4506);
xnor U5927 (N_5927,N_4235,N_3616);
nand U5928 (N_5928,N_4701,N_4519);
xor U5929 (N_5929,N_4131,N_3812);
or U5930 (N_5930,N_3736,N_4070);
and U5931 (N_5931,N_3939,N_4658);
nand U5932 (N_5932,N_4567,N_3818);
and U5933 (N_5933,N_3882,N_4032);
xnor U5934 (N_5934,N_4264,N_4083);
xor U5935 (N_5935,N_3967,N_4595);
nand U5936 (N_5936,N_4267,N_4265);
or U5937 (N_5937,N_4368,N_4154);
and U5938 (N_5938,N_4101,N_3943);
or U5939 (N_5939,N_4465,N_4553);
and U5940 (N_5940,N_4419,N_3988);
nor U5941 (N_5941,N_4297,N_4774);
nor U5942 (N_5942,N_3958,N_4703);
xor U5943 (N_5943,N_4779,N_3837);
xnor U5944 (N_5944,N_4029,N_3718);
nor U5945 (N_5945,N_4688,N_4200);
nand U5946 (N_5946,N_4753,N_4140);
xnor U5947 (N_5947,N_4103,N_4241);
nor U5948 (N_5948,N_4533,N_4029);
or U5949 (N_5949,N_3614,N_4477);
and U5950 (N_5950,N_4479,N_3941);
and U5951 (N_5951,N_4724,N_4098);
and U5952 (N_5952,N_3918,N_4696);
and U5953 (N_5953,N_3838,N_4378);
nor U5954 (N_5954,N_3921,N_3913);
nor U5955 (N_5955,N_4598,N_3850);
nor U5956 (N_5956,N_3637,N_4151);
xor U5957 (N_5957,N_4420,N_4606);
nand U5958 (N_5958,N_4527,N_4534);
nand U5959 (N_5959,N_3825,N_4659);
or U5960 (N_5960,N_4309,N_3641);
or U5961 (N_5961,N_4279,N_3764);
nand U5962 (N_5962,N_4024,N_4365);
and U5963 (N_5963,N_3952,N_4797);
xnor U5964 (N_5964,N_3733,N_4253);
and U5965 (N_5965,N_4747,N_4736);
nand U5966 (N_5966,N_4183,N_4266);
nand U5967 (N_5967,N_4400,N_4587);
nor U5968 (N_5968,N_4381,N_4644);
or U5969 (N_5969,N_4066,N_4751);
nor U5970 (N_5970,N_4626,N_4077);
and U5971 (N_5971,N_4198,N_4102);
xnor U5972 (N_5972,N_3936,N_4720);
nand U5973 (N_5973,N_4549,N_4199);
or U5974 (N_5974,N_4536,N_3667);
nand U5975 (N_5975,N_3951,N_4688);
nor U5976 (N_5976,N_4294,N_4546);
and U5977 (N_5977,N_4737,N_4283);
or U5978 (N_5978,N_4786,N_3755);
xnor U5979 (N_5979,N_3943,N_4351);
and U5980 (N_5980,N_3640,N_3990);
or U5981 (N_5981,N_4716,N_4289);
and U5982 (N_5982,N_4143,N_4752);
nor U5983 (N_5983,N_4565,N_3627);
nor U5984 (N_5984,N_3854,N_3814);
nor U5985 (N_5985,N_3664,N_4440);
and U5986 (N_5986,N_4658,N_4647);
nor U5987 (N_5987,N_3674,N_4320);
and U5988 (N_5988,N_4103,N_4440);
nor U5989 (N_5989,N_4392,N_3613);
or U5990 (N_5990,N_3735,N_4739);
xor U5991 (N_5991,N_3841,N_4497);
and U5992 (N_5992,N_4240,N_4668);
nor U5993 (N_5993,N_4040,N_4332);
xnor U5994 (N_5994,N_3834,N_4244);
or U5995 (N_5995,N_4739,N_4157);
and U5996 (N_5996,N_4709,N_4566);
nand U5997 (N_5997,N_4217,N_3738);
nor U5998 (N_5998,N_4730,N_4011);
xnor U5999 (N_5999,N_4689,N_3815);
nand U6000 (N_6000,N_5740,N_5733);
nand U6001 (N_6001,N_5169,N_5593);
xnor U6002 (N_6002,N_5645,N_4845);
and U6003 (N_6003,N_5874,N_5449);
nor U6004 (N_6004,N_5510,N_5338);
nor U6005 (N_6005,N_5866,N_5054);
or U6006 (N_6006,N_5495,N_5195);
and U6007 (N_6007,N_4924,N_5067);
and U6008 (N_6008,N_5774,N_5313);
nor U6009 (N_6009,N_5957,N_5815);
nand U6010 (N_6010,N_5750,N_5948);
xnor U6011 (N_6011,N_4912,N_5395);
or U6012 (N_6012,N_5309,N_5858);
nand U6013 (N_6013,N_5246,N_5226);
or U6014 (N_6014,N_5613,N_5608);
and U6015 (N_6015,N_5812,N_5217);
xor U6016 (N_6016,N_5837,N_5597);
and U6017 (N_6017,N_5787,N_5039);
or U6018 (N_6018,N_5712,N_5411);
nand U6019 (N_6019,N_4903,N_5864);
nor U6020 (N_6020,N_5611,N_5203);
nor U6021 (N_6021,N_5637,N_4989);
nand U6022 (N_6022,N_5382,N_5487);
nand U6023 (N_6023,N_5739,N_4880);
nand U6024 (N_6024,N_5454,N_5022);
nand U6025 (N_6025,N_5137,N_5481);
nand U6026 (N_6026,N_5698,N_5207);
or U6027 (N_6027,N_5244,N_5018);
xnor U6028 (N_6028,N_5933,N_5677);
xnor U6029 (N_6029,N_5624,N_5404);
nor U6030 (N_6030,N_5991,N_5727);
nand U6031 (N_6031,N_5233,N_5861);
nand U6032 (N_6032,N_5354,N_5814);
and U6033 (N_6033,N_5790,N_5311);
or U6034 (N_6034,N_5116,N_5484);
xor U6035 (N_6035,N_5384,N_5072);
or U6036 (N_6036,N_5974,N_5048);
xor U6037 (N_6037,N_5682,N_5989);
xnor U6038 (N_6038,N_5135,N_5346);
nor U6039 (N_6039,N_5823,N_4864);
nor U6040 (N_6040,N_5418,N_5307);
nand U6041 (N_6041,N_5232,N_5860);
xor U6042 (N_6042,N_5589,N_5049);
xnor U6043 (N_6043,N_5051,N_5716);
nand U6044 (N_6044,N_4981,N_5417);
and U6045 (N_6045,N_5743,N_5155);
nor U6046 (N_6046,N_5040,N_5503);
nand U6047 (N_6047,N_5718,N_5450);
xnor U6048 (N_6048,N_5671,N_5000);
and U6049 (N_6049,N_5667,N_5235);
nor U6050 (N_6050,N_4987,N_5271);
or U6051 (N_6051,N_4841,N_5494);
xnor U6052 (N_6052,N_5185,N_5149);
nand U6053 (N_6053,N_5683,N_4809);
nand U6054 (N_6054,N_4829,N_5196);
xor U6055 (N_6055,N_5227,N_5994);
or U6056 (N_6056,N_5315,N_5436);
or U6057 (N_6057,N_5359,N_4871);
xnor U6058 (N_6058,N_5855,N_5024);
or U6059 (N_6059,N_4850,N_5281);
nor U6060 (N_6060,N_5662,N_5761);
xnor U6061 (N_6061,N_5986,N_5835);
or U6062 (N_6062,N_5713,N_5209);
and U6063 (N_6063,N_5635,N_5703);
nor U6064 (N_6064,N_5690,N_5093);
xnor U6065 (N_6065,N_5324,N_5491);
xor U6066 (N_6066,N_5365,N_4805);
or U6067 (N_6067,N_5279,N_5389);
and U6068 (N_6068,N_5117,N_5465);
or U6069 (N_6069,N_4929,N_5610);
xor U6070 (N_6070,N_5900,N_4890);
xor U6071 (N_6071,N_5824,N_5568);
and U6072 (N_6072,N_5385,N_5876);
or U6073 (N_6073,N_5147,N_5922);
or U6074 (N_6074,N_5139,N_4884);
nor U6075 (N_6075,N_5469,N_5646);
xnor U6076 (N_6076,N_5020,N_5950);
or U6077 (N_6077,N_5615,N_5477);
and U6078 (N_6078,N_5799,N_5930);
nor U6079 (N_6079,N_5165,N_5625);
or U6080 (N_6080,N_5546,N_4975);
nand U6081 (N_6081,N_5993,N_5747);
or U6082 (N_6082,N_5172,N_5390);
and U6083 (N_6083,N_5979,N_5161);
nor U6084 (N_6084,N_4916,N_4966);
xnor U6085 (N_6085,N_5729,N_5959);
or U6086 (N_6086,N_5941,N_5705);
and U6087 (N_6087,N_5951,N_4932);
nand U6088 (N_6088,N_4877,N_5518);
or U6089 (N_6089,N_5471,N_5559);
xnor U6090 (N_6090,N_5334,N_5267);
nand U6091 (N_6091,N_5092,N_5350);
and U6092 (N_6092,N_5089,N_5919);
nor U6093 (N_6093,N_5907,N_5914);
nand U6094 (N_6094,N_5845,N_5759);
nand U6095 (N_6095,N_4906,N_5230);
and U6096 (N_6096,N_5191,N_5619);
nor U6097 (N_6097,N_5838,N_4955);
nand U6098 (N_6098,N_5798,N_5283);
nand U6099 (N_6099,N_5153,N_4858);
or U6100 (N_6100,N_5988,N_5983);
xnor U6101 (N_6101,N_5766,N_5152);
nand U6102 (N_6102,N_5833,N_5136);
xor U6103 (N_6103,N_5679,N_5782);
nor U6104 (N_6104,N_4901,N_5173);
xor U6105 (N_6105,N_5100,N_5428);
or U6106 (N_6106,N_5869,N_5581);
nor U6107 (N_6107,N_5325,N_5508);
or U6108 (N_6108,N_4817,N_5490);
and U6109 (N_6109,N_5038,N_5753);
and U6110 (N_6110,N_5547,N_5300);
or U6111 (N_6111,N_5036,N_5781);
nand U6112 (N_6112,N_5783,N_4852);
nand U6113 (N_6113,N_4902,N_5065);
nand U6114 (N_6114,N_5584,N_5273);
or U6115 (N_6115,N_5827,N_5305);
and U6116 (N_6116,N_5694,N_5516);
or U6117 (N_6117,N_5524,N_4872);
nor U6118 (N_6118,N_4960,N_5160);
nor U6119 (N_6119,N_5556,N_5996);
and U6120 (N_6120,N_4873,N_5660);
or U6121 (N_6121,N_4907,N_5200);
nand U6122 (N_6122,N_5170,N_5184);
and U6123 (N_6123,N_5189,N_5243);
nor U6124 (N_6124,N_4946,N_5058);
or U6125 (N_6125,N_5452,N_5035);
nand U6126 (N_6126,N_5374,N_4979);
nand U6127 (N_6127,N_5251,N_5995);
nor U6128 (N_6128,N_5461,N_5587);
nor U6129 (N_6129,N_5641,N_5882);
nand U6130 (N_6130,N_5744,N_4952);
and U6131 (N_6131,N_5956,N_5938);
nor U6132 (N_6132,N_5258,N_5883);
or U6133 (N_6133,N_5586,N_5985);
xor U6134 (N_6134,N_5872,N_5475);
or U6135 (N_6135,N_4888,N_5725);
or U6136 (N_6136,N_5870,N_5242);
and U6137 (N_6137,N_5541,N_5890);
nand U6138 (N_6138,N_4963,N_5924);
nand U6139 (N_6139,N_5061,N_5090);
or U6140 (N_6140,N_5434,N_5999);
nand U6141 (N_6141,N_5737,N_5424);
or U6142 (N_6142,N_5894,N_5561);
nor U6143 (N_6143,N_4949,N_5125);
xnor U6144 (N_6144,N_5777,N_5296);
nor U6145 (N_6145,N_5129,N_4842);
and U6146 (N_6146,N_4943,N_5275);
and U6147 (N_6147,N_4915,N_5383);
xnor U6148 (N_6148,N_5197,N_5651);
nor U6149 (N_6149,N_5778,N_4839);
nand U6150 (N_6150,N_5765,N_5413);
or U6151 (N_6151,N_5911,N_5032);
xor U6152 (N_6152,N_5198,N_5480);
nand U6153 (N_6153,N_5228,N_4832);
nand U6154 (N_6154,N_5528,N_5786);
xor U6155 (N_6155,N_5339,N_5805);
nand U6156 (N_6156,N_4861,N_5844);
and U6157 (N_6157,N_5954,N_5282);
and U6158 (N_6158,N_5987,N_5083);
or U6159 (N_6159,N_4802,N_4860);
nand U6160 (N_6160,N_5763,N_5926);
xnor U6161 (N_6161,N_5272,N_5818);
nor U6162 (N_6162,N_5086,N_5046);
and U6163 (N_6163,N_5081,N_5499);
nand U6164 (N_6164,N_5885,N_4848);
and U6165 (N_6165,N_5199,N_5157);
nor U6166 (N_6166,N_5509,N_5442);
or U6167 (N_6167,N_4885,N_5447);
and U6168 (N_6168,N_5257,N_5665);
or U6169 (N_6169,N_5111,N_5070);
or U6170 (N_6170,N_4847,N_5362);
nand U6171 (N_6171,N_5310,N_5764);
nor U6172 (N_6172,N_5005,N_5483);
nand U6173 (N_6173,N_4942,N_5700);
and U6174 (N_6174,N_5757,N_5695);
and U6175 (N_6175,N_5632,N_4993);
nand U6176 (N_6176,N_5653,N_4957);
and U6177 (N_6177,N_5981,N_4804);
nand U6178 (N_6178,N_5607,N_5298);
nor U6179 (N_6179,N_5293,N_5785);
nand U6180 (N_6180,N_4807,N_5544);
or U6181 (N_6181,N_5467,N_5287);
xor U6182 (N_6182,N_5056,N_5719);
nand U6183 (N_6183,N_5113,N_5735);
xnor U6184 (N_6184,N_5825,N_5274);
or U6185 (N_6185,N_5723,N_5746);
or U6186 (N_6186,N_5564,N_4810);
xor U6187 (N_6187,N_5224,N_5133);
and U6188 (N_6188,N_4995,N_4976);
nor U6189 (N_6189,N_4856,N_5103);
or U6190 (N_6190,N_5306,N_5636);
or U6191 (N_6191,N_5910,N_5333);
nand U6192 (N_6192,N_4908,N_5468);
and U6193 (N_6193,N_5376,N_5952);
xor U6194 (N_6194,N_5539,N_4862);
nand U6195 (N_6195,N_5323,N_5730);
xnor U6196 (N_6196,N_5820,N_5621);
or U6197 (N_6197,N_4821,N_5696);
and U6198 (N_6198,N_5158,N_4937);
nand U6199 (N_6199,N_5268,N_5532);
and U6200 (N_6200,N_5968,N_5453);
nor U6201 (N_6201,N_5895,N_5406);
or U6202 (N_6202,N_5550,N_5433);
and U6203 (N_6203,N_5237,N_5028);
and U6204 (N_6204,N_5967,N_5462);
nand U6205 (N_6205,N_4803,N_5446);
or U6206 (N_6206,N_4881,N_5329);
nand U6207 (N_6207,N_5806,N_5121);
nor U6208 (N_6208,N_5605,N_5030);
and U6209 (N_6209,N_5706,N_5533);
or U6210 (N_6210,N_5720,N_5771);
or U6211 (N_6211,N_4882,N_5557);
nand U6212 (N_6212,N_5931,N_5141);
nand U6213 (N_6213,N_5708,N_4935);
nor U6214 (N_6214,N_5429,N_5511);
nand U6215 (N_6215,N_5409,N_5552);
xnor U6216 (N_6216,N_4851,N_5015);
nor U6217 (N_6217,N_4961,N_5364);
and U6218 (N_6218,N_5650,N_5183);
and U6219 (N_6219,N_5134,N_5962);
xor U6220 (N_6220,N_5127,N_4868);
xnor U6221 (N_6221,N_5913,N_5043);
and U6222 (N_6222,N_5915,N_5692);
or U6223 (N_6223,N_5391,N_5050);
xnor U6224 (N_6224,N_5684,N_5534);
xnor U6225 (N_6225,N_5222,N_5167);
xnor U6226 (N_6226,N_5029,N_4956);
nand U6227 (N_6227,N_4876,N_5617);
nand U6228 (N_6228,N_5724,N_5856);
and U6229 (N_6229,N_5213,N_5571);
nor U6230 (N_6230,N_4824,N_5314);
nor U6231 (N_6231,N_4998,N_5025);
nor U6232 (N_6232,N_5520,N_5810);
and U6233 (N_6233,N_4909,N_4933);
and U6234 (N_6234,N_5977,N_5105);
or U6235 (N_6235,N_4835,N_5891);
nor U6236 (N_6236,N_4997,N_4920);
nor U6237 (N_6237,N_5109,N_5661);
or U6238 (N_6238,N_5801,N_5789);
nand U6239 (N_6239,N_5351,N_5639);
nand U6240 (N_6240,N_5361,N_5201);
and U6241 (N_6241,N_5657,N_5128);
nand U6242 (N_6242,N_5091,N_5179);
xnor U6243 (N_6243,N_5019,N_5375);
nor U6244 (N_6244,N_5772,N_5253);
or U6245 (N_6245,N_5037,N_4918);
or U6246 (N_6246,N_5622,N_5088);
and U6247 (N_6247,N_4926,N_4863);
nand U6248 (N_6248,N_4971,N_5102);
and U6249 (N_6249,N_5905,N_5349);
nor U6250 (N_6250,N_4819,N_5960);
and U6251 (N_6251,N_5563,N_5848);
nand U6252 (N_6252,N_5084,N_5412);
and U6253 (N_6253,N_5939,N_5330);
and U6254 (N_6254,N_5208,N_5360);
or U6255 (N_6255,N_4934,N_5558);
nor U6256 (N_6256,N_5675,N_4944);
or U6257 (N_6257,N_5321,N_5535);
or U6258 (N_6258,N_5863,N_5920);
xnor U6259 (N_6259,N_5145,N_5479);
xnor U6260 (N_6260,N_4816,N_5033);
and U6261 (N_6261,N_5548,N_5800);
nand U6262 (N_6262,N_5337,N_5304);
nor U6263 (N_6263,N_5672,N_5123);
or U6264 (N_6264,N_5669,N_5980);
nand U6265 (N_6265,N_5817,N_5071);
xor U6266 (N_6266,N_5438,N_5752);
nand U6267 (N_6267,N_5488,N_5175);
nor U6268 (N_6268,N_5372,N_5796);
nand U6269 (N_6269,N_5756,N_5717);
xnor U6270 (N_6270,N_5080,N_5041);
or U6271 (N_6271,N_5734,N_5598);
xnor U6272 (N_6272,N_5807,N_5302);
or U6273 (N_6273,N_4859,N_5699);
and U6274 (N_6274,N_5601,N_5249);
or U6275 (N_6275,N_5500,N_5223);
and U6276 (N_6276,N_5654,N_5923);
and U6277 (N_6277,N_5248,N_5400);
nand U6278 (N_6278,N_4990,N_5620);
and U6279 (N_6279,N_5972,N_4867);
nand U6280 (N_6280,N_5573,N_5463);
nand U6281 (N_6281,N_5430,N_5498);
and U6282 (N_6282,N_4844,N_5021);
nor U6283 (N_6283,N_5431,N_5928);
xor U6284 (N_6284,N_4853,N_5347);
and U6285 (N_6285,N_4973,N_5935);
or U6286 (N_6286,N_4875,N_5068);
nand U6287 (N_6287,N_4964,N_5678);
nand U6288 (N_6288,N_4836,N_5537);
nand U6289 (N_6289,N_4895,N_4823);
nand U6290 (N_6290,N_5663,N_4854);
and U6291 (N_6291,N_5936,N_5888);
nand U6292 (N_6292,N_5131,N_5476);
and U6293 (N_6293,N_5403,N_5378);
or U6294 (N_6294,N_5748,N_5371);
or U6295 (N_6295,N_5770,N_5252);
nand U6296 (N_6296,N_5009,N_5523);
xor U6297 (N_6297,N_5240,N_5178);
or U6298 (N_6298,N_5187,N_5691);
and U6299 (N_6299,N_4921,N_5921);
nor U6300 (N_6300,N_5059,N_5368);
nand U6301 (N_6301,N_5414,N_5358);
and U6302 (N_6302,N_5204,N_5205);
nor U6303 (N_6303,N_5388,N_5604);
nand U6304 (N_6304,N_5906,N_5932);
xnor U6305 (N_6305,N_5822,N_5085);
nor U6306 (N_6306,N_5702,N_5647);
nand U6307 (N_6307,N_5640,N_5370);
xor U6308 (N_6308,N_5012,N_5426);
nand U6309 (N_6309,N_4857,N_5241);
xor U6310 (N_6310,N_5808,N_5754);
nor U6311 (N_6311,N_5685,N_5419);
nor U6312 (N_6312,N_5834,N_4917);
and U6313 (N_6313,N_5514,N_5758);
xnor U6314 (N_6314,N_5367,N_5878);
xor U6315 (N_6315,N_5961,N_5773);
xnor U6316 (N_6316,N_5576,N_5964);
or U6317 (N_6317,N_5676,N_5002);
xor U6318 (N_6318,N_5707,N_4919);
xor U6319 (N_6319,N_5410,N_5643);
nand U6320 (N_6320,N_5115,N_5946);
or U6321 (N_6321,N_5852,N_5842);
or U6322 (N_6322,N_5316,N_4965);
nand U6323 (N_6323,N_4813,N_5963);
or U6324 (N_6324,N_5269,N_5373);
nor U6325 (N_6325,N_5633,N_5369);
and U6326 (N_6326,N_5423,N_5689);
and U6327 (N_6327,N_5031,N_4840);
xnor U6328 (N_6328,N_5623,N_5212);
or U6329 (N_6329,N_5513,N_5862);
and U6330 (N_6330,N_5631,N_5343);
nor U6331 (N_6331,N_5775,N_5859);
and U6332 (N_6332,N_5760,N_5506);
nor U6333 (N_6333,N_5577,N_5655);
or U6334 (N_6334,N_5877,N_5401);
xor U6335 (N_6335,N_5344,N_5027);
xnor U6336 (N_6336,N_5585,N_5457);
or U6337 (N_6337,N_5236,N_5104);
xor U6338 (N_6338,N_4977,N_5278);
nand U6339 (N_6339,N_5190,N_5828);
nor U6340 (N_6340,N_5288,N_5762);
nor U6341 (N_6341,N_5319,N_5944);
nor U6342 (N_6342,N_5357,N_5245);
xor U6343 (N_6343,N_5472,N_5231);
or U6344 (N_6344,N_4889,N_5722);
and U6345 (N_6345,N_4914,N_5555);
nand U6346 (N_6346,N_5507,N_5194);
nand U6347 (N_6347,N_5975,N_5816);
and U6348 (N_6348,N_4978,N_5688);
nand U6349 (N_6349,N_5892,N_5515);
and U6350 (N_6350,N_5420,N_5318);
and U6351 (N_6351,N_5206,N_5386);
or U6352 (N_6352,N_5711,N_5943);
xor U6353 (N_6353,N_5148,N_5482);
xor U6354 (N_6354,N_5425,N_4991);
nor U6355 (N_6355,N_4996,N_5399);
nor U6356 (N_6356,N_5501,N_5973);
nand U6357 (N_6357,N_5182,N_4814);
nor U6358 (N_6358,N_5908,N_5057);
xor U6359 (N_6359,N_5074,N_5188);
or U6360 (N_6360,N_5299,N_5784);
and U6361 (N_6361,N_5405,N_5704);
nor U6362 (N_6362,N_5791,N_5693);
or U6363 (N_6363,N_5984,N_5077);
nor U6364 (N_6364,N_5016,N_5794);
nand U6365 (N_6365,N_5902,N_5210);
nand U6366 (N_6366,N_4838,N_5710);
or U6367 (N_6367,N_5875,N_5427);
and U6368 (N_6368,N_4970,N_4897);
nor U6369 (N_6369,N_4808,N_5776);
or U6370 (N_6370,N_5638,N_5893);
nand U6371 (N_6371,N_5879,N_4988);
nand U6372 (N_6372,N_5238,N_5536);
or U6373 (N_6373,N_5470,N_4982);
xnor U6374 (N_6374,N_5966,N_5603);
xor U6375 (N_6375,N_5732,N_5277);
and U6376 (N_6376,N_5211,N_5466);
xor U6377 (N_6377,N_5285,N_5751);
xor U6378 (N_6378,N_4967,N_5830);
nand U6379 (N_6379,N_5998,N_4865);
xnor U6380 (N_6380,N_4843,N_4968);
and U6381 (N_6381,N_5052,N_5478);
and U6382 (N_6382,N_5918,N_4800);
xnor U6383 (N_6383,N_5073,N_5297);
nor U6384 (N_6384,N_5947,N_5076);
nor U6385 (N_6385,N_5408,N_5545);
nor U6386 (N_6386,N_5916,N_4958);
nand U6387 (N_6387,N_5062,N_4939);
and U6388 (N_6388,N_5517,N_5122);
xnor U6389 (N_6389,N_5821,N_5949);
xor U6390 (N_6390,N_5832,N_5697);
nand U6391 (N_6391,N_5075,N_5898);
xnor U6392 (N_6392,N_4849,N_5749);
or U6393 (N_6393,N_5473,N_5353);
nand U6394 (N_6394,N_5927,N_5909);
nor U6395 (N_6395,N_5606,N_5439);
xnor U6396 (N_6396,N_5079,N_5779);
nor U6397 (N_6397,N_4931,N_5502);
xnor U6398 (N_6398,N_4994,N_5320);
nand U6399 (N_6399,N_4833,N_5045);
or U6400 (N_6400,N_5336,N_5925);
xor U6401 (N_6401,N_5579,N_5332);
nand U6402 (N_6402,N_5867,N_5392);
xor U6403 (N_6403,N_5899,N_5095);
xnor U6404 (N_6404,N_5819,N_5276);
nor U6405 (N_6405,N_5110,N_5460);
xnor U6406 (N_6406,N_5687,N_5112);
xnor U6407 (N_6407,N_4874,N_5937);
nor U6408 (N_6408,N_5529,N_5441);
xor U6409 (N_6409,N_5997,N_5574);
and U6410 (N_6410,N_4940,N_4896);
nor U6411 (N_6411,N_5728,N_5250);
nor U6412 (N_6412,N_5387,N_4905);
nor U6413 (N_6413,N_5327,N_5138);
nor U6414 (N_6414,N_5263,N_5456);
nor U6415 (N_6415,N_5124,N_5831);
xnor U6416 (N_6416,N_5459,N_5202);
nor U6417 (N_6417,N_5301,N_5114);
nand U6418 (N_6418,N_5745,N_5560);
and U6419 (N_6419,N_5259,N_4886);
xor U6420 (N_6420,N_5247,N_4891);
nor U6421 (N_6421,N_5982,N_5549);
nor U6422 (N_6422,N_4951,N_5525);
nand U6423 (N_6423,N_5118,N_5168);
or U6424 (N_6424,N_5917,N_5627);
and U6425 (N_6425,N_5255,N_5595);
or U6426 (N_6426,N_5616,N_5393);
nand U6427 (N_6427,N_5596,N_5780);
xnor U6428 (N_6428,N_5013,N_5591);
nand U6429 (N_6429,N_5542,N_5955);
or U6430 (N_6430,N_5873,N_5396);
nand U6431 (N_6431,N_5006,N_5570);
nor U6432 (N_6432,N_5142,N_5652);
nor U6433 (N_6433,N_5670,N_5363);
nor U6434 (N_6434,N_5871,N_5034);
and U6435 (N_6435,N_5140,N_5366);
and U6436 (N_6436,N_5398,N_5254);
nor U6437 (N_6437,N_5341,N_5220);
nor U6438 (N_6438,N_4883,N_5214);
nand U6439 (N_6439,N_5826,N_5099);
nand U6440 (N_6440,N_5126,N_4986);
nand U6441 (N_6441,N_4974,N_5286);
xor U6442 (N_6442,N_5565,N_5648);
nand U6443 (N_6443,N_4938,N_5069);
or U6444 (N_6444,N_5225,N_5380);
and U6445 (N_6445,N_5265,N_4941);
or U6446 (N_6446,N_4969,N_5379);
and U6447 (N_6447,N_4869,N_5990);
nor U6448 (N_6448,N_5171,N_5726);
or U6449 (N_6449,N_5294,N_5458);
nand U6450 (N_6450,N_5853,N_5177);
or U6451 (N_6451,N_4900,N_5176);
nand U6452 (N_6452,N_5489,N_5192);
and U6453 (N_6453,N_5096,N_5234);
nand U6454 (N_6454,N_4899,N_5144);
or U6455 (N_6455,N_5889,N_5680);
and U6456 (N_6456,N_5714,N_5256);
nand U6457 (N_6457,N_4923,N_5101);
and U6458 (N_6458,N_5444,N_5519);
nand U6459 (N_6459,N_5312,N_5464);
nor U6460 (N_6460,N_4992,N_5664);
nand U6461 (N_6461,N_4827,N_5261);
and U6462 (N_6462,N_5011,N_5912);
xnor U6463 (N_6463,N_4928,N_4984);
xnor U6464 (N_6464,N_5897,N_5221);
xnor U6465 (N_6465,N_5886,N_5668);
nand U6466 (N_6466,N_5108,N_5901);
nand U6467 (N_6467,N_5649,N_4815);
xnor U6468 (N_6468,N_5569,N_5394);
xor U6469 (N_6469,N_5813,N_5580);
xor U6470 (N_6470,N_5978,N_4831);
nand U6471 (N_6471,N_5965,N_5792);
nor U6472 (N_6472,N_5609,N_5602);
and U6473 (N_6473,N_5865,N_5451);
and U6474 (N_6474,N_5163,N_4887);
xor U6475 (N_6475,N_4947,N_5673);
and U6476 (N_6476,N_5042,N_5159);
or U6477 (N_6477,N_5934,N_5497);
nand U6478 (N_6478,N_5992,N_5342);
nand U6479 (N_6479,N_4825,N_5162);
and U6480 (N_6480,N_5348,N_5106);
nand U6481 (N_6481,N_5849,N_5001);
nand U6482 (N_6482,N_5284,N_5836);
xnor U6483 (N_6483,N_5493,N_5004);
nor U6484 (N_6484,N_5397,N_4870);
nor U6485 (N_6485,N_4820,N_5970);
and U6486 (N_6486,N_5094,N_4904);
or U6487 (N_6487,N_5066,N_5857);
and U6488 (N_6488,N_4959,N_5448);
xnor U6489 (N_6489,N_5098,N_5229);
xnor U6490 (N_6490,N_5521,N_5219);
nand U6491 (N_6491,N_5328,N_5402);
nand U6492 (N_6492,N_5239,N_4972);
nor U6493 (N_6493,N_4922,N_4950);
xor U6494 (N_6494,N_5715,N_5130);
nand U6495 (N_6495,N_5087,N_5797);
nor U6496 (N_6496,N_5809,N_4945);
or U6497 (N_6497,N_5017,N_4826);
and U6498 (N_6498,N_4980,N_5686);
xor U6499 (N_6499,N_5674,N_5701);
and U6500 (N_6500,N_4893,N_5023);
nor U6501 (N_6501,N_5082,N_4925);
and U6502 (N_6502,N_5644,N_4878);
or U6503 (N_6503,N_5270,N_5280);
or U6504 (N_6504,N_5566,N_5626);
xor U6505 (N_6505,N_5097,N_5156);
xnor U6506 (N_6506,N_5007,N_5958);
or U6507 (N_6507,N_5578,N_5854);
xnor U6508 (N_6508,N_5326,N_5415);
xor U6509 (N_6509,N_5345,N_4846);
xnor U6510 (N_6510,N_5795,N_5811);
or U6511 (N_6511,N_5146,N_5971);
and U6512 (N_6512,N_5562,N_5512);
and U6513 (N_6513,N_5377,N_4936);
and U6514 (N_6514,N_5078,N_5527);
and U6515 (N_6515,N_4948,N_5634);
nor U6516 (N_6516,N_5896,N_5421);
and U6517 (N_6517,N_5215,N_4855);
nand U6518 (N_6518,N_5588,N_4812);
and U6519 (N_6519,N_5903,N_5666);
and U6520 (N_6520,N_5014,N_5166);
nor U6521 (N_6521,N_4962,N_5060);
xnor U6522 (N_6522,N_5572,N_5107);
xnor U6523 (N_6523,N_5969,N_5154);
nor U6524 (N_6524,N_5736,N_5355);
xnor U6525 (N_6525,N_5485,N_5590);
nor U6526 (N_6526,N_5440,N_4818);
and U6527 (N_6527,N_5583,N_5174);
or U6528 (N_6528,N_5193,N_5945);
nand U6529 (N_6529,N_5047,N_5308);
nor U6530 (N_6530,N_4822,N_4898);
or U6531 (N_6531,N_5904,N_5731);
nor U6532 (N_6532,N_5741,N_5445);
nor U6533 (N_6533,N_5614,N_5769);
and U6534 (N_6534,N_5437,N_5681);
or U6535 (N_6535,N_5435,N_5432);
xnor U6536 (N_6536,N_5151,N_5150);
and U6537 (N_6537,N_5292,N_5804);
or U6538 (N_6538,N_5260,N_5767);
nand U6539 (N_6539,N_5884,N_5592);
and U6540 (N_6540,N_5599,N_5492);
and U6541 (N_6541,N_4930,N_5003);
nand U6542 (N_6542,N_5522,N_5340);
or U6543 (N_6543,N_5120,N_5322);
or U6544 (N_6544,N_5504,N_4837);
or U6545 (N_6545,N_5612,N_4983);
xnor U6546 (N_6546,N_5538,N_5422);
or U6547 (N_6547,N_5181,N_4911);
xor U6548 (N_6548,N_5290,N_5486);
or U6549 (N_6549,N_4913,N_4892);
xor U6550 (N_6550,N_5543,N_4830);
nor U6551 (N_6551,N_5505,N_5530);
xor U6552 (N_6552,N_5868,N_5553);
nor U6553 (N_6553,N_5618,N_5053);
nor U6554 (N_6554,N_4894,N_5738);
or U6555 (N_6555,N_5407,N_5180);
xnor U6556 (N_6556,N_5540,N_5356);
nand U6557 (N_6557,N_5317,N_5658);
nand U6558 (N_6558,N_5803,N_5262);
xnor U6559 (N_6559,N_5443,N_5026);
nor U6560 (N_6560,N_5953,N_4999);
and U6561 (N_6561,N_5331,N_5940);
or U6562 (N_6562,N_5594,N_5843);
nand U6563 (N_6563,N_5829,N_5887);
nand U6564 (N_6564,N_5802,N_5629);
and U6565 (N_6565,N_5788,N_5455);
or U6566 (N_6566,N_5416,N_4866);
nor U6567 (N_6567,N_5526,N_5218);
nand U6568 (N_6568,N_5628,N_5929);
nand U6569 (N_6569,N_5008,N_5742);
nor U6570 (N_6570,N_5851,N_5289);
xnor U6571 (N_6571,N_5840,N_4985);
xnor U6572 (N_6572,N_5976,N_5942);
xnor U6573 (N_6573,N_4879,N_5656);
or U6574 (N_6574,N_5847,N_5755);
nor U6575 (N_6575,N_5709,N_5055);
or U6576 (N_6576,N_4910,N_4811);
or U6577 (N_6577,N_5567,N_5531);
xor U6578 (N_6578,N_5295,N_4828);
or U6579 (N_6579,N_4954,N_4927);
and U6580 (N_6580,N_5793,N_5474);
nand U6581 (N_6581,N_5551,N_5768);
nand U6582 (N_6582,N_5381,N_5186);
nand U6583 (N_6583,N_5303,N_5264);
xnor U6584 (N_6584,N_5496,N_5839);
nor U6585 (N_6585,N_4806,N_5850);
and U6586 (N_6586,N_5335,N_5721);
nor U6587 (N_6587,N_5600,N_5216);
or U6588 (N_6588,N_5846,N_5064);
xnor U6589 (N_6589,N_5266,N_4953);
xnor U6590 (N_6590,N_5010,N_5881);
nor U6591 (N_6591,N_5063,N_5582);
or U6592 (N_6592,N_5291,N_5880);
and U6593 (N_6593,N_5642,N_5164);
xor U6594 (N_6594,N_5119,N_5841);
nor U6595 (N_6595,N_5132,N_5630);
xor U6596 (N_6596,N_4834,N_5575);
nor U6597 (N_6597,N_4801,N_5659);
or U6598 (N_6598,N_5352,N_5554);
xnor U6599 (N_6599,N_5044,N_5143);
xnor U6600 (N_6600,N_5229,N_5402);
nor U6601 (N_6601,N_4865,N_5883);
xnor U6602 (N_6602,N_5336,N_5613);
or U6603 (N_6603,N_5848,N_5989);
nor U6604 (N_6604,N_5700,N_5643);
and U6605 (N_6605,N_5555,N_5876);
xnor U6606 (N_6606,N_5823,N_5353);
nor U6607 (N_6607,N_5000,N_4976);
xnor U6608 (N_6608,N_5142,N_5884);
nor U6609 (N_6609,N_4802,N_5072);
nor U6610 (N_6610,N_5322,N_5325);
or U6611 (N_6611,N_5399,N_5082);
xor U6612 (N_6612,N_5928,N_5104);
nor U6613 (N_6613,N_5905,N_4993);
nor U6614 (N_6614,N_5002,N_5746);
xor U6615 (N_6615,N_5516,N_5116);
nand U6616 (N_6616,N_5517,N_5164);
nor U6617 (N_6617,N_4880,N_5145);
nor U6618 (N_6618,N_5052,N_5861);
nor U6619 (N_6619,N_5764,N_5208);
xor U6620 (N_6620,N_4960,N_5513);
or U6621 (N_6621,N_5908,N_5558);
and U6622 (N_6622,N_5639,N_5126);
nand U6623 (N_6623,N_5162,N_5423);
or U6624 (N_6624,N_5968,N_5192);
nor U6625 (N_6625,N_4847,N_4993);
nand U6626 (N_6626,N_5144,N_5932);
nand U6627 (N_6627,N_5619,N_5154);
nand U6628 (N_6628,N_5863,N_5718);
nor U6629 (N_6629,N_4965,N_5903);
or U6630 (N_6630,N_5979,N_4829);
nand U6631 (N_6631,N_5462,N_5915);
nand U6632 (N_6632,N_5958,N_5249);
nand U6633 (N_6633,N_5011,N_5669);
nor U6634 (N_6634,N_4937,N_5512);
or U6635 (N_6635,N_4930,N_5665);
nor U6636 (N_6636,N_5783,N_5481);
xnor U6637 (N_6637,N_4894,N_5241);
nand U6638 (N_6638,N_5621,N_5766);
or U6639 (N_6639,N_5452,N_5175);
and U6640 (N_6640,N_5649,N_5159);
and U6641 (N_6641,N_5819,N_4933);
nand U6642 (N_6642,N_5884,N_5312);
nor U6643 (N_6643,N_5139,N_4895);
nand U6644 (N_6644,N_5693,N_5754);
xor U6645 (N_6645,N_5852,N_5546);
and U6646 (N_6646,N_5473,N_5145);
nor U6647 (N_6647,N_4835,N_5683);
nand U6648 (N_6648,N_5856,N_5741);
and U6649 (N_6649,N_5079,N_5362);
and U6650 (N_6650,N_5148,N_5417);
or U6651 (N_6651,N_5500,N_5871);
and U6652 (N_6652,N_5296,N_5130);
and U6653 (N_6653,N_5442,N_4953);
and U6654 (N_6654,N_5640,N_5932);
and U6655 (N_6655,N_5089,N_5028);
nand U6656 (N_6656,N_5352,N_4963);
or U6657 (N_6657,N_5383,N_5844);
xnor U6658 (N_6658,N_5206,N_5195);
nor U6659 (N_6659,N_4847,N_4920);
nand U6660 (N_6660,N_5754,N_5395);
nand U6661 (N_6661,N_5081,N_5078);
nand U6662 (N_6662,N_5323,N_5155);
or U6663 (N_6663,N_5683,N_5632);
or U6664 (N_6664,N_5011,N_5077);
or U6665 (N_6665,N_5299,N_4899);
or U6666 (N_6666,N_4806,N_5013);
nand U6667 (N_6667,N_5991,N_5857);
or U6668 (N_6668,N_5754,N_5873);
or U6669 (N_6669,N_5405,N_4943);
nand U6670 (N_6670,N_5470,N_5186);
and U6671 (N_6671,N_5197,N_5362);
and U6672 (N_6672,N_5289,N_5649);
nand U6673 (N_6673,N_5374,N_5996);
nor U6674 (N_6674,N_5386,N_5779);
and U6675 (N_6675,N_5796,N_5594);
nor U6676 (N_6676,N_5760,N_5764);
nand U6677 (N_6677,N_5719,N_5126);
nor U6678 (N_6678,N_5136,N_4915);
or U6679 (N_6679,N_5948,N_5154);
and U6680 (N_6680,N_4920,N_4970);
xnor U6681 (N_6681,N_4985,N_5343);
or U6682 (N_6682,N_5548,N_5722);
nor U6683 (N_6683,N_4930,N_5469);
nand U6684 (N_6684,N_5497,N_5642);
and U6685 (N_6685,N_5830,N_5642);
and U6686 (N_6686,N_4923,N_5450);
nand U6687 (N_6687,N_4975,N_5119);
nand U6688 (N_6688,N_5949,N_5025);
xnor U6689 (N_6689,N_5088,N_5964);
nand U6690 (N_6690,N_5088,N_4818);
nor U6691 (N_6691,N_5265,N_5848);
nor U6692 (N_6692,N_4869,N_5805);
nand U6693 (N_6693,N_5478,N_5841);
nand U6694 (N_6694,N_5514,N_5210);
or U6695 (N_6695,N_5770,N_5281);
nor U6696 (N_6696,N_5059,N_5573);
or U6697 (N_6697,N_5468,N_5515);
or U6698 (N_6698,N_5640,N_5505);
or U6699 (N_6699,N_5712,N_5021);
nor U6700 (N_6700,N_5027,N_5087);
and U6701 (N_6701,N_5310,N_4812);
xnor U6702 (N_6702,N_5403,N_5860);
nor U6703 (N_6703,N_5691,N_5790);
xnor U6704 (N_6704,N_5417,N_5894);
nand U6705 (N_6705,N_5061,N_5889);
and U6706 (N_6706,N_5854,N_4983);
nor U6707 (N_6707,N_5172,N_5865);
and U6708 (N_6708,N_5499,N_5861);
nand U6709 (N_6709,N_5770,N_5385);
or U6710 (N_6710,N_4816,N_5530);
and U6711 (N_6711,N_4908,N_5200);
nand U6712 (N_6712,N_5959,N_5989);
nand U6713 (N_6713,N_5954,N_5584);
or U6714 (N_6714,N_5932,N_4983);
or U6715 (N_6715,N_5094,N_5563);
and U6716 (N_6716,N_5244,N_5392);
nand U6717 (N_6717,N_5641,N_5108);
and U6718 (N_6718,N_5275,N_5226);
xnor U6719 (N_6719,N_5762,N_5682);
or U6720 (N_6720,N_4946,N_5812);
xnor U6721 (N_6721,N_5110,N_5500);
xor U6722 (N_6722,N_4896,N_5926);
or U6723 (N_6723,N_5412,N_5745);
xnor U6724 (N_6724,N_5315,N_5839);
nor U6725 (N_6725,N_5140,N_5123);
or U6726 (N_6726,N_5651,N_5770);
or U6727 (N_6727,N_5330,N_5804);
xor U6728 (N_6728,N_4879,N_5354);
nand U6729 (N_6729,N_5396,N_5457);
xnor U6730 (N_6730,N_4892,N_5019);
and U6731 (N_6731,N_5064,N_5235);
nor U6732 (N_6732,N_5517,N_5609);
nor U6733 (N_6733,N_5440,N_5229);
nand U6734 (N_6734,N_5422,N_5241);
or U6735 (N_6735,N_5860,N_4802);
or U6736 (N_6736,N_4901,N_5285);
nand U6737 (N_6737,N_5525,N_5316);
or U6738 (N_6738,N_5885,N_5708);
xor U6739 (N_6739,N_5069,N_5571);
nor U6740 (N_6740,N_5925,N_5659);
xnor U6741 (N_6741,N_5667,N_4832);
and U6742 (N_6742,N_5364,N_5396);
nor U6743 (N_6743,N_5572,N_5897);
and U6744 (N_6744,N_4831,N_5917);
or U6745 (N_6745,N_5864,N_4803);
and U6746 (N_6746,N_5184,N_5968);
and U6747 (N_6747,N_4976,N_5294);
or U6748 (N_6748,N_5141,N_5670);
xnor U6749 (N_6749,N_5384,N_5251);
or U6750 (N_6750,N_4835,N_4864);
nand U6751 (N_6751,N_5144,N_5101);
nand U6752 (N_6752,N_5470,N_5489);
nor U6753 (N_6753,N_5698,N_5019);
nand U6754 (N_6754,N_5414,N_5346);
nor U6755 (N_6755,N_5722,N_4978);
and U6756 (N_6756,N_5934,N_4887);
xnor U6757 (N_6757,N_5076,N_5326);
nor U6758 (N_6758,N_5080,N_5872);
xor U6759 (N_6759,N_5590,N_5781);
or U6760 (N_6760,N_5521,N_5752);
xnor U6761 (N_6761,N_4818,N_5126);
or U6762 (N_6762,N_5249,N_5277);
or U6763 (N_6763,N_5822,N_4930);
xnor U6764 (N_6764,N_5200,N_5360);
nand U6765 (N_6765,N_5690,N_5667);
or U6766 (N_6766,N_5884,N_5750);
or U6767 (N_6767,N_5341,N_5429);
and U6768 (N_6768,N_5201,N_5065);
nand U6769 (N_6769,N_5798,N_5772);
or U6770 (N_6770,N_5758,N_5306);
nand U6771 (N_6771,N_5093,N_5916);
xor U6772 (N_6772,N_4868,N_5159);
xor U6773 (N_6773,N_5749,N_5948);
or U6774 (N_6774,N_5020,N_5828);
and U6775 (N_6775,N_5037,N_5680);
and U6776 (N_6776,N_5341,N_5167);
nand U6777 (N_6777,N_5905,N_5234);
xor U6778 (N_6778,N_5438,N_5539);
xor U6779 (N_6779,N_5890,N_5715);
and U6780 (N_6780,N_5528,N_5688);
or U6781 (N_6781,N_5571,N_5477);
nand U6782 (N_6782,N_5743,N_5705);
xnor U6783 (N_6783,N_5682,N_5926);
xnor U6784 (N_6784,N_4878,N_5400);
nor U6785 (N_6785,N_5433,N_5837);
nor U6786 (N_6786,N_5009,N_5731);
and U6787 (N_6787,N_5684,N_5681);
or U6788 (N_6788,N_5836,N_5883);
nor U6789 (N_6789,N_4953,N_5884);
nor U6790 (N_6790,N_5135,N_5391);
nand U6791 (N_6791,N_5724,N_4937);
or U6792 (N_6792,N_5700,N_4908);
nor U6793 (N_6793,N_5026,N_4814);
nor U6794 (N_6794,N_5453,N_5395);
and U6795 (N_6795,N_5421,N_5014);
nor U6796 (N_6796,N_5521,N_5488);
nor U6797 (N_6797,N_4827,N_5542);
nand U6798 (N_6798,N_5577,N_5788);
nand U6799 (N_6799,N_5066,N_5279);
xnor U6800 (N_6800,N_5916,N_5044);
xnor U6801 (N_6801,N_5228,N_5093);
and U6802 (N_6802,N_5535,N_5877);
xnor U6803 (N_6803,N_5495,N_5966);
nand U6804 (N_6804,N_4844,N_4814);
xor U6805 (N_6805,N_5365,N_5117);
nand U6806 (N_6806,N_5779,N_5320);
nand U6807 (N_6807,N_5698,N_5872);
nor U6808 (N_6808,N_5035,N_5262);
or U6809 (N_6809,N_5389,N_4986);
nor U6810 (N_6810,N_5156,N_5108);
or U6811 (N_6811,N_5657,N_5080);
or U6812 (N_6812,N_5529,N_5302);
nand U6813 (N_6813,N_4829,N_5391);
and U6814 (N_6814,N_5190,N_5155);
nand U6815 (N_6815,N_5155,N_5239);
nand U6816 (N_6816,N_5281,N_4875);
nand U6817 (N_6817,N_5634,N_5681);
nand U6818 (N_6818,N_5537,N_5884);
nand U6819 (N_6819,N_5208,N_5999);
xnor U6820 (N_6820,N_5338,N_5913);
or U6821 (N_6821,N_5652,N_4922);
nor U6822 (N_6822,N_4866,N_5420);
xor U6823 (N_6823,N_5095,N_5043);
or U6824 (N_6824,N_5514,N_5296);
and U6825 (N_6825,N_5065,N_5192);
xor U6826 (N_6826,N_5226,N_5153);
and U6827 (N_6827,N_5158,N_5622);
nor U6828 (N_6828,N_5576,N_5672);
and U6829 (N_6829,N_5178,N_5015);
xor U6830 (N_6830,N_5350,N_5154);
and U6831 (N_6831,N_5782,N_5943);
and U6832 (N_6832,N_5430,N_5746);
nand U6833 (N_6833,N_5391,N_5618);
nand U6834 (N_6834,N_5367,N_5700);
and U6835 (N_6835,N_5963,N_5139);
nand U6836 (N_6836,N_5382,N_5755);
nor U6837 (N_6837,N_5950,N_5686);
or U6838 (N_6838,N_5288,N_5752);
nand U6839 (N_6839,N_4957,N_5469);
nand U6840 (N_6840,N_5220,N_5105);
nand U6841 (N_6841,N_5656,N_5299);
and U6842 (N_6842,N_5273,N_5956);
nand U6843 (N_6843,N_5835,N_5224);
and U6844 (N_6844,N_4899,N_5566);
xnor U6845 (N_6845,N_5665,N_5466);
xor U6846 (N_6846,N_5619,N_5717);
nand U6847 (N_6847,N_5082,N_5521);
xnor U6848 (N_6848,N_5561,N_5171);
and U6849 (N_6849,N_4809,N_5487);
nor U6850 (N_6850,N_5376,N_5217);
or U6851 (N_6851,N_5787,N_5354);
nand U6852 (N_6852,N_5375,N_5568);
and U6853 (N_6853,N_5459,N_5217);
nor U6854 (N_6854,N_5612,N_4832);
nand U6855 (N_6855,N_5858,N_5166);
nor U6856 (N_6856,N_4871,N_5996);
nor U6857 (N_6857,N_5684,N_4818);
nor U6858 (N_6858,N_5199,N_5246);
or U6859 (N_6859,N_5195,N_5373);
nor U6860 (N_6860,N_5971,N_4967);
and U6861 (N_6861,N_5515,N_5859);
xor U6862 (N_6862,N_4910,N_5558);
nand U6863 (N_6863,N_4964,N_5220);
nand U6864 (N_6864,N_4983,N_5320);
or U6865 (N_6865,N_5639,N_5705);
nor U6866 (N_6866,N_5009,N_5500);
and U6867 (N_6867,N_5847,N_4997);
xor U6868 (N_6868,N_5677,N_5499);
nand U6869 (N_6869,N_4832,N_5153);
xnor U6870 (N_6870,N_4994,N_5087);
xor U6871 (N_6871,N_5102,N_5207);
or U6872 (N_6872,N_5347,N_5050);
nor U6873 (N_6873,N_5358,N_5469);
or U6874 (N_6874,N_5851,N_5391);
nor U6875 (N_6875,N_5794,N_5806);
and U6876 (N_6876,N_5027,N_4840);
nor U6877 (N_6877,N_5872,N_5114);
nor U6878 (N_6878,N_5863,N_5680);
nand U6879 (N_6879,N_5872,N_5746);
or U6880 (N_6880,N_5642,N_5777);
nor U6881 (N_6881,N_5581,N_5470);
nand U6882 (N_6882,N_5307,N_5583);
or U6883 (N_6883,N_5457,N_5233);
or U6884 (N_6884,N_5779,N_5069);
xnor U6885 (N_6885,N_5206,N_5685);
nor U6886 (N_6886,N_4902,N_5204);
xor U6887 (N_6887,N_4850,N_5077);
xnor U6888 (N_6888,N_5263,N_5635);
nor U6889 (N_6889,N_5971,N_5507);
and U6890 (N_6890,N_5074,N_5985);
nand U6891 (N_6891,N_5069,N_5450);
and U6892 (N_6892,N_4845,N_4830);
and U6893 (N_6893,N_5993,N_5097);
xnor U6894 (N_6894,N_5043,N_4843);
xor U6895 (N_6895,N_5605,N_4821);
nand U6896 (N_6896,N_5973,N_5843);
or U6897 (N_6897,N_5337,N_5601);
and U6898 (N_6898,N_5750,N_5258);
nand U6899 (N_6899,N_5104,N_5389);
and U6900 (N_6900,N_5328,N_5907);
and U6901 (N_6901,N_5124,N_5409);
xor U6902 (N_6902,N_5684,N_5784);
nand U6903 (N_6903,N_5508,N_5863);
nand U6904 (N_6904,N_4905,N_5362);
xor U6905 (N_6905,N_5450,N_5285);
or U6906 (N_6906,N_5543,N_5189);
or U6907 (N_6907,N_5510,N_5317);
nor U6908 (N_6908,N_5034,N_4985);
nor U6909 (N_6909,N_5759,N_5415);
xnor U6910 (N_6910,N_5428,N_5471);
xnor U6911 (N_6911,N_5345,N_5293);
or U6912 (N_6912,N_5724,N_5148);
or U6913 (N_6913,N_5992,N_5966);
nor U6914 (N_6914,N_5175,N_5533);
nor U6915 (N_6915,N_5995,N_5420);
xnor U6916 (N_6916,N_5229,N_4853);
xor U6917 (N_6917,N_5909,N_5764);
and U6918 (N_6918,N_5508,N_5865);
or U6919 (N_6919,N_5071,N_5207);
and U6920 (N_6920,N_5472,N_5462);
and U6921 (N_6921,N_5494,N_5772);
or U6922 (N_6922,N_5102,N_5039);
nor U6923 (N_6923,N_4865,N_5326);
xor U6924 (N_6924,N_5819,N_5063);
and U6925 (N_6925,N_5882,N_4978);
xnor U6926 (N_6926,N_5906,N_5170);
or U6927 (N_6927,N_4969,N_5387);
and U6928 (N_6928,N_5599,N_4819);
nand U6929 (N_6929,N_5071,N_5068);
nand U6930 (N_6930,N_5829,N_5252);
xor U6931 (N_6931,N_5928,N_5869);
nand U6932 (N_6932,N_5287,N_5508);
xor U6933 (N_6933,N_5832,N_5495);
or U6934 (N_6934,N_5048,N_5321);
nor U6935 (N_6935,N_5428,N_5702);
or U6936 (N_6936,N_4943,N_5538);
nand U6937 (N_6937,N_5875,N_5415);
and U6938 (N_6938,N_5469,N_5801);
xor U6939 (N_6939,N_5573,N_5047);
or U6940 (N_6940,N_4811,N_5466);
and U6941 (N_6941,N_5879,N_4866);
and U6942 (N_6942,N_5133,N_5652);
or U6943 (N_6943,N_5230,N_5950);
or U6944 (N_6944,N_5019,N_5421);
and U6945 (N_6945,N_5290,N_5888);
nor U6946 (N_6946,N_5847,N_5801);
nor U6947 (N_6947,N_5416,N_5046);
and U6948 (N_6948,N_5014,N_5408);
xnor U6949 (N_6949,N_5049,N_5407);
or U6950 (N_6950,N_5278,N_4952);
and U6951 (N_6951,N_5548,N_4810);
and U6952 (N_6952,N_5075,N_5702);
xor U6953 (N_6953,N_5923,N_5608);
nand U6954 (N_6954,N_5322,N_5881);
nor U6955 (N_6955,N_5697,N_5616);
and U6956 (N_6956,N_5007,N_5633);
and U6957 (N_6957,N_4810,N_4906);
nand U6958 (N_6958,N_5406,N_5731);
and U6959 (N_6959,N_5412,N_5457);
nor U6960 (N_6960,N_5327,N_5177);
xnor U6961 (N_6961,N_5886,N_5318);
and U6962 (N_6962,N_5322,N_5934);
nand U6963 (N_6963,N_5283,N_5953);
and U6964 (N_6964,N_4958,N_4915);
nand U6965 (N_6965,N_5981,N_5704);
nand U6966 (N_6966,N_4811,N_5502);
nor U6967 (N_6967,N_5083,N_5552);
nor U6968 (N_6968,N_5207,N_4990);
nor U6969 (N_6969,N_5023,N_5763);
nor U6970 (N_6970,N_5121,N_5690);
or U6971 (N_6971,N_4974,N_5439);
or U6972 (N_6972,N_4816,N_4858);
or U6973 (N_6973,N_5088,N_5326);
xnor U6974 (N_6974,N_4852,N_4903);
and U6975 (N_6975,N_5537,N_5414);
and U6976 (N_6976,N_5331,N_5475);
and U6977 (N_6977,N_5536,N_5116);
xor U6978 (N_6978,N_4821,N_5493);
or U6979 (N_6979,N_5883,N_5037);
nor U6980 (N_6980,N_5519,N_5637);
and U6981 (N_6981,N_5776,N_4887);
or U6982 (N_6982,N_5219,N_5948);
nor U6983 (N_6983,N_5881,N_4955);
xor U6984 (N_6984,N_5856,N_5745);
nor U6985 (N_6985,N_5917,N_5474);
xor U6986 (N_6986,N_4807,N_5108);
and U6987 (N_6987,N_5866,N_5110);
xnor U6988 (N_6988,N_5565,N_5113);
and U6989 (N_6989,N_5024,N_5317);
and U6990 (N_6990,N_5085,N_5776);
or U6991 (N_6991,N_5225,N_5349);
nand U6992 (N_6992,N_5090,N_4994);
or U6993 (N_6993,N_5379,N_5677);
xor U6994 (N_6994,N_5337,N_5314);
nor U6995 (N_6995,N_5494,N_5641);
xnor U6996 (N_6996,N_5541,N_5510);
nor U6997 (N_6997,N_4885,N_5843);
nor U6998 (N_6998,N_4992,N_5859);
nand U6999 (N_6999,N_5284,N_5833);
nor U7000 (N_7000,N_5596,N_4891);
and U7001 (N_7001,N_5256,N_4813);
nor U7002 (N_7002,N_5864,N_4877);
and U7003 (N_7003,N_5761,N_5341);
nor U7004 (N_7004,N_5257,N_5581);
or U7005 (N_7005,N_5018,N_5704);
or U7006 (N_7006,N_5046,N_5272);
and U7007 (N_7007,N_5653,N_5802);
nor U7008 (N_7008,N_5985,N_5493);
nand U7009 (N_7009,N_5729,N_5974);
nand U7010 (N_7010,N_5021,N_5918);
nor U7011 (N_7011,N_5824,N_5834);
nor U7012 (N_7012,N_4863,N_4910);
nand U7013 (N_7013,N_4931,N_4982);
xor U7014 (N_7014,N_5899,N_5096);
nand U7015 (N_7015,N_5519,N_5340);
nor U7016 (N_7016,N_5198,N_4878);
xnor U7017 (N_7017,N_5311,N_5363);
and U7018 (N_7018,N_4841,N_5974);
and U7019 (N_7019,N_5005,N_4983);
nor U7020 (N_7020,N_4999,N_4900);
nor U7021 (N_7021,N_5758,N_5883);
or U7022 (N_7022,N_5871,N_5030);
xor U7023 (N_7023,N_5722,N_5050);
and U7024 (N_7024,N_5751,N_5491);
nor U7025 (N_7025,N_5857,N_5796);
nor U7026 (N_7026,N_5845,N_5704);
nor U7027 (N_7027,N_5865,N_5554);
nand U7028 (N_7028,N_5454,N_5093);
nand U7029 (N_7029,N_5282,N_4800);
xor U7030 (N_7030,N_5976,N_5888);
nand U7031 (N_7031,N_5996,N_4863);
xor U7032 (N_7032,N_5401,N_5058);
nor U7033 (N_7033,N_5009,N_5504);
nor U7034 (N_7034,N_5413,N_5896);
or U7035 (N_7035,N_4919,N_5852);
nor U7036 (N_7036,N_5271,N_5151);
xor U7037 (N_7037,N_5187,N_5353);
nand U7038 (N_7038,N_5130,N_5821);
nor U7039 (N_7039,N_4905,N_5882);
and U7040 (N_7040,N_4906,N_5203);
or U7041 (N_7041,N_5437,N_5967);
and U7042 (N_7042,N_5083,N_5960);
and U7043 (N_7043,N_5285,N_5074);
nand U7044 (N_7044,N_4949,N_5670);
or U7045 (N_7045,N_5068,N_5513);
nand U7046 (N_7046,N_5936,N_5281);
or U7047 (N_7047,N_5441,N_5982);
or U7048 (N_7048,N_5925,N_5568);
nand U7049 (N_7049,N_5645,N_5091);
xnor U7050 (N_7050,N_5610,N_5263);
or U7051 (N_7051,N_5785,N_5749);
nor U7052 (N_7052,N_5984,N_5223);
nor U7053 (N_7053,N_5999,N_5133);
or U7054 (N_7054,N_5200,N_4874);
or U7055 (N_7055,N_5453,N_5573);
and U7056 (N_7056,N_5931,N_5292);
nand U7057 (N_7057,N_5115,N_5352);
and U7058 (N_7058,N_4992,N_5178);
and U7059 (N_7059,N_4999,N_5481);
nor U7060 (N_7060,N_5348,N_5153);
nand U7061 (N_7061,N_5581,N_5830);
and U7062 (N_7062,N_5514,N_4869);
nand U7063 (N_7063,N_5787,N_5105);
and U7064 (N_7064,N_5187,N_5119);
and U7065 (N_7065,N_5664,N_5194);
xor U7066 (N_7066,N_5594,N_5914);
nor U7067 (N_7067,N_5177,N_4897);
nor U7068 (N_7068,N_5022,N_5335);
nand U7069 (N_7069,N_5764,N_5145);
nor U7070 (N_7070,N_5499,N_5988);
or U7071 (N_7071,N_5113,N_5768);
and U7072 (N_7072,N_5738,N_5702);
nand U7073 (N_7073,N_5251,N_5308);
nand U7074 (N_7074,N_5864,N_5018);
nor U7075 (N_7075,N_5523,N_5088);
nor U7076 (N_7076,N_5222,N_5035);
xor U7077 (N_7077,N_5980,N_5600);
xnor U7078 (N_7078,N_5486,N_5836);
xnor U7079 (N_7079,N_5245,N_4974);
nand U7080 (N_7080,N_5002,N_4817);
xnor U7081 (N_7081,N_4964,N_5850);
nand U7082 (N_7082,N_5614,N_5680);
and U7083 (N_7083,N_5055,N_5768);
nor U7084 (N_7084,N_5547,N_5903);
nor U7085 (N_7085,N_4945,N_5469);
nand U7086 (N_7086,N_5535,N_5854);
nor U7087 (N_7087,N_4836,N_5296);
nand U7088 (N_7088,N_4811,N_5435);
xnor U7089 (N_7089,N_5447,N_4969);
nand U7090 (N_7090,N_5108,N_5301);
xnor U7091 (N_7091,N_5678,N_5705);
and U7092 (N_7092,N_5078,N_5135);
and U7093 (N_7093,N_5349,N_5515);
xor U7094 (N_7094,N_5333,N_5511);
and U7095 (N_7095,N_5830,N_4886);
and U7096 (N_7096,N_5032,N_5863);
and U7097 (N_7097,N_5408,N_4885);
nand U7098 (N_7098,N_5964,N_4912);
nor U7099 (N_7099,N_5275,N_5619);
nor U7100 (N_7100,N_5520,N_5959);
or U7101 (N_7101,N_5895,N_5833);
nor U7102 (N_7102,N_5328,N_5903);
xor U7103 (N_7103,N_5337,N_5088);
or U7104 (N_7104,N_5548,N_4844);
xor U7105 (N_7105,N_5493,N_5387);
and U7106 (N_7106,N_5839,N_5506);
nand U7107 (N_7107,N_4984,N_5102);
xnor U7108 (N_7108,N_5771,N_5099);
nand U7109 (N_7109,N_4926,N_4960);
nand U7110 (N_7110,N_5795,N_5911);
nor U7111 (N_7111,N_4869,N_5699);
nor U7112 (N_7112,N_5122,N_5349);
xor U7113 (N_7113,N_4905,N_5063);
or U7114 (N_7114,N_4810,N_5519);
nand U7115 (N_7115,N_5534,N_5060);
nor U7116 (N_7116,N_5739,N_5838);
or U7117 (N_7117,N_5875,N_5042);
nand U7118 (N_7118,N_5262,N_5845);
nor U7119 (N_7119,N_5984,N_4975);
nand U7120 (N_7120,N_5639,N_5050);
xnor U7121 (N_7121,N_5301,N_5891);
xor U7122 (N_7122,N_5864,N_5846);
or U7123 (N_7123,N_5830,N_5533);
xnor U7124 (N_7124,N_4899,N_5199);
and U7125 (N_7125,N_4958,N_4948);
nand U7126 (N_7126,N_5198,N_5290);
nand U7127 (N_7127,N_5693,N_5441);
nor U7128 (N_7128,N_5579,N_5596);
nand U7129 (N_7129,N_5091,N_5868);
and U7130 (N_7130,N_5671,N_5087);
or U7131 (N_7131,N_4939,N_4970);
xnor U7132 (N_7132,N_5222,N_5511);
xnor U7133 (N_7133,N_5195,N_5589);
nand U7134 (N_7134,N_5322,N_5256);
or U7135 (N_7135,N_4815,N_5010);
or U7136 (N_7136,N_5921,N_5561);
xnor U7137 (N_7137,N_5722,N_5670);
and U7138 (N_7138,N_5271,N_5697);
xnor U7139 (N_7139,N_5380,N_5173);
or U7140 (N_7140,N_5985,N_5000);
xnor U7141 (N_7141,N_5774,N_5279);
nor U7142 (N_7142,N_5143,N_5770);
or U7143 (N_7143,N_4949,N_5939);
nor U7144 (N_7144,N_5977,N_5267);
nor U7145 (N_7145,N_5209,N_5583);
and U7146 (N_7146,N_5591,N_5636);
xor U7147 (N_7147,N_5583,N_5087);
xor U7148 (N_7148,N_5968,N_5604);
or U7149 (N_7149,N_5833,N_5801);
or U7150 (N_7150,N_5974,N_5880);
and U7151 (N_7151,N_5462,N_4878);
nand U7152 (N_7152,N_5409,N_5910);
xnor U7153 (N_7153,N_5902,N_5315);
xnor U7154 (N_7154,N_5428,N_5255);
xor U7155 (N_7155,N_5999,N_5515);
nor U7156 (N_7156,N_5655,N_5146);
and U7157 (N_7157,N_5580,N_4805);
and U7158 (N_7158,N_5407,N_4868);
nor U7159 (N_7159,N_5947,N_5351);
nand U7160 (N_7160,N_5134,N_5527);
or U7161 (N_7161,N_4925,N_5966);
nand U7162 (N_7162,N_4982,N_5102);
and U7163 (N_7163,N_5791,N_5808);
or U7164 (N_7164,N_5548,N_5514);
or U7165 (N_7165,N_5876,N_5580);
nor U7166 (N_7166,N_5309,N_5033);
nand U7167 (N_7167,N_5335,N_5906);
nor U7168 (N_7168,N_5068,N_4822);
or U7169 (N_7169,N_4867,N_5983);
nand U7170 (N_7170,N_4848,N_4856);
nor U7171 (N_7171,N_5409,N_5300);
xnor U7172 (N_7172,N_5046,N_5661);
or U7173 (N_7173,N_5347,N_5443);
and U7174 (N_7174,N_5877,N_5556);
and U7175 (N_7175,N_4864,N_5183);
nor U7176 (N_7176,N_5018,N_5464);
and U7177 (N_7177,N_5205,N_5707);
nand U7178 (N_7178,N_5519,N_5493);
xnor U7179 (N_7179,N_5735,N_5088);
xnor U7180 (N_7180,N_5779,N_5746);
or U7181 (N_7181,N_4960,N_5917);
nand U7182 (N_7182,N_5679,N_5870);
nor U7183 (N_7183,N_5650,N_5424);
or U7184 (N_7184,N_5635,N_5393);
nand U7185 (N_7185,N_5935,N_4890);
or U7186 (N_7186,N_5692,N_5523);
nand U7187 (N_7187,N_5247,N_5101);
and U7188 (N_7188,N_5868,N_5293);
nand U7189 (N_7189,N_4858,N_5548);
or U7190 (N_7190,N_4823,N_5446);
nand U7191 (N_7191,N_4894,N_5521);
nor U7192 (N_7192,N_5903,N_5811);
nor U7193 (N_7193,N_5074,N_5714);
nor U7194 (N_7194,N_5046,N_5833);
nand U7195 (N_7195,N_5614,N_4804);
nand U7196 (N_7196,N_5554,N_5479);
nor U7197 (N_7197,N_5800,N_5336);
and U7198 (N_7198,N_4930,N_4836);
nor U7199 (N_7199,N_5313,N_5438);
nor U7200 (N_7200,N_6048,N_6512);
nand U7201 (N_7201,N_6702,N_7174);
nand U7202 (N_7202,N_6737,N_6606);
or U7203 (N_7203,N_6957,N_6570);
nor U7204 (N_7204,N_6477,N_6920);
and U7205 (N_7205,N_6097,N_6880);
and U7206 (N_7206,N_6523,N_6172);
nor U7207 (N_7207,N_6678,N_7047);
nor U7208 (N_7208,N_6826,N_6584);
nand U7209 (N_7209,N_6549,N_6428);
xor U7210 (N_7210,N_6436,N_6771);
or U7211 (N_7211,N_7070,N_6076);
or U7212 (N_7212,N_6065,N_6710);
or U7213 (N_7213,N_6996,N_6390);
or U7214 (N_7214,N_6267,N_6630);
nand U7215 (N_7215,N_6592,N_6786);
and U7216 (N_7216,N_6564,N_6548);
or U7217 (N_7217,N_7161,N_6491);
nor U7218 (N_7218,N_6220,N_6358);
nand U7219 (N_7219,N_6833,N_6940);
nand U7220 (N_7220,N_7065,N_6795);
xor U7221 (N_7221,N_6949,N_6042);
and U7222 (N_7222,N_6945,N_6779);
nand U7223 (N_7223,N_6073,N_6007);
and U7224 (N_7224,N_6655,N_6524);
and U7225 (N_7225,N_6553,N_6603);
nor U7226 (N_7226,N_6251,N_6960);
nand U7227 (N_7227,N_6993,N_6003);
and U7228 (N_7228,N_6250,N_7199);
and U7229 (N_7229,N_6917,N_7057);
nand U7230 (N_7230,N_6219,N_6983);
nor U7231 (N_7231,N_6359,N_6522);
or U7232 (N_7232,N_6284,N_7151);
nand U7233 (N_7233,N_6961,N_7133);
xor U7234 (N_7234,N_6615,N_6486);
nand U7235 (N_7235,N_6914,N_6860);
xnor U7236 (N_7236,N_7190,N_6700);
or U7237 (N_7237,N_6970,N_7004);
or U7238 (N_7238,N_6425,N_6688);
or U7239 (N_7239,N_6823,N_6879);
nor U7240 (N_7240,N_6034,N_6542);
and U7241 (N_7241,N_6560,N_6714);
and U7242 (N_7242,N_6004,N_6598);
xor U7243 (N_7243,N_6239,N_6056);
nor U7244 (N_7244,N_6376,N_6739);
or U7245 (N_7245,N_6127,N_7073);
nor U7246 (N_7246,N_6232,N_6399);
and U7247 (N_7247,N_6723,N_6275);
or U7248 (N_7248,N_6400,N_6478);
or U7249 (N_7249,N_7055,N_7157);
nor U7250 (N_7250,N_6517,N_6035);
nand U7251 (N_7251,N_6104,N_6608);
and U7252 (N_7252,N_6892,N_6883);
and U7253 (N_7253,N_6083,N_6045);
nand U7254 (N_7254,N_6125,N_7132);
nor U7255 (N_7255,N_6255,N_6488);
xnor U7256 (N_7256,N_6939,N_6938);
or U7257 (N_7257,N_6278,N_6263);
nor U7258 (N_7258,N_6314,N_6841);
and U7259 (N_7259,N_6117,N_6270);
xnor U7260 (N_7260,N_7138,N_6618);
xnor U7261 (N_7261,N_6438,N_7056);
nor U7262 (N_7262,N_6385,N_6431);
nand U7263 (N_7263,N_6569,N_6345);
nor U7264 (N_7264,N_7184,N_6504);
nand U7265 (N_7265,N_7107,N_7109);
xnor U7266 (N_7266,N_6855,N_6550);
or U7267 (N_7267,N_6595,N_6266);
and U7268 (N_7268,N_6862,N_6762);
nor U7269 (N_7269,N_6043,N_7134);
xor U7270 (N_7270,N_6333,N_6370);
and U7271 (N_7271,N_7061,N_6760);
or U7272 (N_7272,N_7117,N_6613);
nand U7273 (N_7273,N_7052,N_6306);
nor U7274 (N_7274,N_6360,N_7049);
and U7275 (N_7275,N_7009,N_6759);
nand U7276 (N_7276,N_6093,N_7035);
nand U7277 (N_7277,N_6373,N_6601);
and U7278 (N_7278,N_6330,N_6936);
xor U7279 (N_7279,N_6619,N_6651);
or U7280 (N_7280,N_6672,N_6181);
nor U7281 (N_7281,N_6455,N_6780);
nand U7282 (N_7282,N_6871,N_6470);
and U7283 (N_7283,N_6673,N_6268);
nand U7284 (N_7284,N_6062,N_7054);
or U7285 (N_7285,N_7045,N_6930);
and U7286 (N_7286,N_6616,N_6353);
or U7287 (N_7287,N_6234,N_6120);
or U7288 (N_7288,N_6927,N_6843);
or U7289 (N_7289,N_6393,N_7021);
nand U7290 (N_7290,N_6371,N_7153);
nor U7291 (N_7291,N_6646,N_6767);
xnor U7292 (N_7292,N_6667,N_6769);
nand U7293 (N_7293,N_7016,N_6958);
xor U7294 (N_7294,N_6011,N_6775);
xor U7295 (N_7295,N_6822,N_6893);
and U7296 (N_7296,N_6364,N_6772);
nand U7297 (N_7297,N_6214,N_6622);
nand U7298 (N_7298,N_6139,N_6382);
or U7299 (N_7299,N_6184,N_6933);
xnor U7300 (N_7300,N_6343,N_6866);
and U7301 (N_7301,N_6900,N_6135);
and U7302 (N_7302,N_6674,N_6396);
xor U7303 (N_7303,N_6025,N_6935);
and U7304 (N_7304,N_6080,N_7014);
or U7305 (N_7305,N_6213,N_7002);
or U7306 (N_7306,N_6475,N_6956);
nor U7307 (N_7307,N_6644,N_6877);
nor U7308 (N_7308,N_6221,N_6310);
or U7309 (N_7309,N_6742,N_6583);
xor U7310 (N_7310,N_6963,N_6988);
or U7311 (N_7311,N_6844,N_6785);
xor U7312 (N_7312,N_6567,N_7062);
or U7313 (N_7313,N_6163,N_6694);
or U7314 (N_7314,N_6827,N_6476);
and U7315 (N_7315,N_6487,N_7189);
or U7316 (N_7316,N_6367,N_7029);
nand U7317 (N_7317,N_6401,N_6185);
or U7318 (N_7318,N_6816,N_6562);
and U7319 (N_7319,N_6543,N_6224);
or U7320 (N_7320,N_6577,N_6179);
nor U7321 (N_7321,N_7112,N_6037);
nor U7322 (N_7322,N_6008,N_6212);
nor U7323 (N_7323,N_6864,N_7075);
or U7324 (N_7324,N_6908,N_6555);
nand U7325 (N_7325,N_6623,N_6675);
or U7326 (N_7326,N_6812,N_6439);
and U7327 (N_7327,N_7118,N_6624);
nor U7328 (N_7328,N_6617,N_7091);
or U7329 (N_7329,N_6269,N_6128);
nor U7330 (N_7330,N_6049,N_6433);
nand U7331 (N_7331,N_7180,N_6614);
or U7332 (N_7332,N_6283,N_6208);
nor U7333 (N_7333,N_7089,N_6303);
or U7334 (N_7334,N_6637,N_6151);
xor U7335 (N_7335,N_6334,N_6663);
or U7336 (N_7336,N_6051,N_6755);
or U7337 (N_7337,N_6464,N_6317);
nor U7338 (N_7338,N_6122,N_6799);
nor U7339 (N_7339,N_6471,N_6994);
nor U7340 (N_7340,N_7114,N_6347);
nor U7341 (N_7341,N_6468,N_6490);
nand U7342 (N_7342,N_6660,N_6059);
nor U7343 (N_7343,N_6260,N_6916);
or U7344 (N_7344,N_6017,N_6563);
or U7345 (N_7345,N_6050,N_7003);
or U7346 (N_7346,N_6206,N_6225);
and U7347 (N_7347,N_6964,N_6332);
nor U7348 (N_7348,N_6951,N_6783);
xnor U7349 (N_7349,N_7131,N_6625);
nor U7350 (N_7350,N_6777,N_6261);
nor U7351 (N_7351,N_6946,N_7160);
nand U7352 (N_7352,N_6537,N_6676);
nand U7353 (N_7353,N_6934,N_6680);
or U7354 (N_7354,N_6743,N_7148);
nor U7355 (N_7355,N_6539,N_6254);
and U7356 (N_7356,N_6873,N_6684);
and U7357 (N_7357,N_6797,N_6247);
nor U7358 (N_7358,N_6978,N_6813);
and U7359 (N_7359,N_6718,N_6990);
or U7360 (N_7360,N_6513,N_6108);
nand U7361 (N_7361,N_6324,N_6895);
or U7362 (N_7362,N_6285,N_6015);
nor U7363 (N_7363,N_6599,N_6658);
nor U7364 (N_7364,N_6405,N_6469);
or U7365 (N_7365,N_6001,N_6510);
nor U7366 (N_7366,N_6642,N_6271);
nor U7367 (N_7367,N_6194,N_6540);
and U7368 (N_7368,N_6292,N_6987);
nor U7369 (N_7369,N_6578,N_6369);
xor U7370 (N_7370,N_7159,N_6643);
xnor U7371 (N_7371,N_6046,N_6701);
or U7372 (N_7372,N_6137,N_6919);
nand U7373 (N_7373,N_6495,N_6969);
nand U7374 (N_7374,N_6532,N_6915);
xnor U7375 (N_7375,N_7186,N_6472);
xnor U7376 (N_7376,N_6818,N_6904);
and U7377 (N_7377,N_6559,N_6389);
and U7378 (N_7378,N_7135,N_7121);
and U7379 (N_7379,N_6174,N_6244);
nand U7380 (N_7380,N_6609,N_6350);
or U7381 (N_7381,N_6055,N_6064);
and U7382 (N_7382,N_7092,N_6276);
or U7383 (N_7383,N_6657,N_6384);
nand U7384 (N_7384,N_7042,N_6806);
nand U7385 (N_7385,N_6666,N_6620);
nand U7386 (N_7386,N_6689,N_6547);
and U7387 (N_7387,N_6123,N_7013);
xnor U7388 (N_7388,N_6596,N_6725);
nand U7389 (N_7389,N_6148,N_6849);
nor U7390 (N_7390,N_7071,N_6729);
xnor U7391 (N_7391,N_6773,N_6107);
xnor U7392 (N_7392,N_6754,N_6290);
and U7393 (N_7393,N_6748,N_6852);
xnor U7394 (N_7394,N_7077,N_6200);
nand U7395 (N_7395,N_6294,N_6287);
nor U7396 (N_7396,N_6499,N_6561);
xnor U7397 (N_7397,N_7169,N_6337);
or U7398 (N_7398,N_6650,N_6634);
or U7399 (N_7399,N_6311,N_6661);
nand U7400 (N_7400,N_7156,N_6516);
nand U7401 (N_7401,N_6395,N_7123);
or U7402 (N_7402,N_6552,N_6182);
and U7403 (N_7403,N_6419,N_6236);
nand U7404 (N_7404,N_6098,N_6568);
or U7405 (N_7405,N_6321,N_6440);
nor U7406 (N_7406,N_6834,N_6801);
xor U7407 (N_7407,N_6421,N_6077);
or U7408 (N_7408,N_6581,N_6837);
nand U7409 (N_7409,N_6467,N_6511);
xor U7410 (N_7410,N_6288,N_7129);
nor U7411 (N_7411,N_6538,N_6363);
nor U7412 (N_7412,N_6697,N_6183);
xor U7413 (N_7413,N_6340,N_6848);
nand U7414 (N_7414,N_6096,N_6331);
or U7415 (N_7415,N_6685,N_6227);
and U7416 (N_7416,N_6966,N_6109);
and U7417 (N_7417,N_6918,N_6256);
and U7418 (N_7418,N_6020,N_6106);
and U7419 (N_7419,N_6989,N_6410);
nor U7420 (N_7420,N_6505,N_7187);
or U7421 (N_7421,N_6078,N_6707);
or U7422 (N_7422,N_6901,N_6279);
xnor U7423 (N_7423,N_6836,N_6665);
xor U7424 (N_7424,N_6944,N_6398);
and U7425 (N_7425,N_6351,N_6835);
nor U7426 (N_7426,N_6000,N_6085);
nor U7427 (N_7427,N_6764,N_7194);
and U7428 (N_7428,N_6872,N_7191);
nand U7429 (N_7429,N_6972,N_7149);
nor U7430 (N_7430,N_6721,N_6747);
xor U7431 (N_7431,N_6067,N_6053);
and U7432 (N_7432,N_6089,N_6506);
nand U7433 (N_7433,N_6164,N_6429);
or U7434 (N_7434,N_6361,N_6659);
and U7435 (N_7435,N_6447,N_6272);
xor U7436 (N_7436,N_6088,N_6036);
and U7437 (N_7437,N_6820,N_6210);
nand U7438 (N_7438,N_6289,N_6422);
nor U7439 (N_7439,N_6652,N_6190);
nor U7440 (N_7440,N_6201,N_6962);
and U7441 (N_7441,N_7053,N_7173);
nand U7442 (N_7442,N_6162,N_6329);
nor U7443 (N_7443,N_7110,N_6437);
xor U7444 (N_7444,N_6832,N_7136);
xnor U7445 (N_7445,N_7098,N_6840);
xnor U7446 (N_7446,N_6636,N_6842);
nor U7447 (N_7447,N_6146,N_7176);
or U7448 (N_7448,N_6626,N_6325);
and U7449 (N_7449,N_6002,N_6508);
or U7450 (N_7450,N_6407,N_7111);
or U7451 (N_7451,N_6030,N_6264);
nand U7452 (N_7452,N_6095,N_6061);
nand U7453 (N_7453,N_6341,N_6793);
and U7454 (N_7454,N_7104,N_6662);
and U7455 (N_7455,N_6922,N_6984);
xor U7456 (N_7456,N_6235,N_6168);
nand U7457 (N_7457,N_7080,N_6484);
xnor U7458 (N_7458,N_6991,N_6403);
and U7459 (N_7459,N_6454,N_6355);
nor U7460 (N_7460,N_6905,N_6796);
or U7461 (N_7461,N_6838,N_6903);
xnor U7462 (N_7462,N_6556,N_7005);
or U7463 (N_7463,N_6683,N_6316);
xnor U7464 (N_7464,N_6995,N_7020);
xnor U7465 (N_7465,N_6100,N_6968);
nand U7466 (N_7466,N_7168,N_6992);
nor U7467 (N_7467,N_6830,N_6291);
nand U7468 (N_7468,N_6753,N_6750);
nand U7469 (N_7469,N_6870,N_7001);
xnor U7470 (N_7470,N_6379,N_6604);
and U7471 (N_7471,N_6377,N_7196);
nor U7472 (N_7472,N_6483,N_6829);
or U7473 (N_7473,N_7094,N_6896);
or U7474 (N_7474,N_6889,N_6152);
and U7475 (N_7475,N_7141,N_6752);
nand U7476 (N_7476,N_6633,N_6894);
and U7477 (N_7477,N_6228,N_7158);
nand U7478 (N_7478,N_7048,N_6886);
nor U7479 (N_7479,N_6249,N_7126);
nor U7480 (N_7480,N_7103,N_6302);
nand U7481 (N_7481,N_6485,N_6924);
or U7482 (N_7482,N_6735,N_6142);
xnor U7483 (N_7483,N_6656,N_6515);
nand U7484 (N_7484,N_6189,N_6259);
or U7485 (N_7485,N_7068,N_7183);
or U7486 (N_7486,N_6173,N_6971);
and U7487 (N_7487,N_6166,N_6044);
xnor U7488 (N_7488,N_6815,N_7167);
or U7489 (N_7489,N_6071,N_6891);
nor U7490 (N_7490,N_6932,N_6144);
or U7491 (N_7491,N_6890,N_6640);
xnor U7492 (N_7492,N_6790,N_6509);
nor U7493 (N_7493,N_6241,N_6831);
nor U7494 (N_7494,N_7147,N_6457);
xnor U7495 (N_7495,N_6209,N_6010);
xnor U7496 (N_7496,N_6621,N_6418);
xor U7497 (N_7497,N_7090,N_6867);
nand U7498 (N_7498,N_6408,N_7011);
nor U7499 (N_7499,N_6335,N_6416);
xor U7500 (N_7500,N_6277,N_6372);
nor U7501 (N_7501,N_6388,N_7051);
and U7502 (N_7502,N_6222,N_6998);
xnor U7503 (N_7503,N_6309,N_6315);
xnor U7504 (N_7504,N_6865,N_6923);
nand U7505 (N_7505,N_6397,N_7015);
nor U7506 (N_7506,N_6589,N_6708);
nor U7507 (N_7507,N_6068,N_6653);
and U7508 (N_7508,N_6641,N_6888);
xor U7509 (N_7509,N_6566,N_6082);
or U7510 (N_7510,N_6161,N_6952);
or U7511 (N_7511,N_6380,N_6446);
and U7512 (N_7512,N_6788,N_6420);
nand U7513 (N_7513,N_6459,N_6086);
or U7514 (N_7514,N_7175,N_7027);
and U7515 (N_7515,N_7120,N_6114);
and U7516 (N_7516,N_6012,N_6414);
and U7517 (N_7517,N_6713,N_6943);
and U7518 (N_7518,N_7113,N_6501);
or U7519 (N_7519,N_6591,N_6023);
nor U7520 (N_7520,N_6105,N_6774);
nor U7521 (N_7521,N_6323,N_7119);
and U7522 (N_7522,N_6233,N_6435);
nor U7523 (N_7523,N_6899,N_6925);
and U7524 (N_7524,N_6032,N_7012);
and U7525 (N_7525,N_6745,N_6942);
or U7526 (N_7526,N_6715,N_6463);
xor U7527 (N_7527,N_6734,N_6778);
xnor U7528 (N_7528,N_6448,N_6196);
or U7529 (N_7529,N_6479,N_6937);
xnor U7530 (N_7530,N_6452,N_6804);
nor U7531 (N_7531,N_6973,N_6784);
xnor U7532 (N_7532,N_6632,N_7026);
or U7533 (N_7533,N_6383,N_6521);
and U7534 (N_7534,N_7099,N_6594);
and U7535 (N_7535,N_7178,N_6502);
nor U7536 (N_7536,N_6544,N_6977);
nor U7537 (N_7537,N_6134,N_6014);
nand U7538 (N_7538,N_6557,N_6293);
xnor U7539 (N_7539,N_6198,N_7017);
xor U7540 (N_7540,N_6029,N_6950);
nor U7541 (N_7541,N_6686,N_6462);
nand U7542 (N_7542,N_6911,N_6074);
xnor U7543 (N_7543,N_7019,N_6980);
and U7544 (N_7544,N_6404,N_7101);
and U7545 (N_7545,N_6704,N_7166);
nor U7546 (N_7546,N_6248,N_6282);
nand U7547 (N_7547,N_6580,N_7185);
nor U7548 (N_7548,N_6824,N_6009);
xor U7549 (N_7549,N_6079,N_6298);
xnor U7550 (N_7550,N_7179,N_6781);
or U7551 (N_7551,N_6038,N_6041);
nor U7552 (N_7552,N_6965,N_6197);
and U7553 (N_7553,N_6703,N_7018);
nor U7554 (N_7554,N_6348,N_6295);
nand U7555 (N_7555,N_6926,N_6126);
nor U7556 (N_7556,N_6758,N_6195);
xor U7557 (N_7557,N_6597,N_7164);
or U7558 (N_7558,N_6687,N_6770);
or U7559 (N_7559,N_6300,N_6741);
xnor U7560 (N_7560,N_7124,N_7100);
nor U7561 (N_7561,N_6845,N_7031);
and U7562 (N_7562,N_6541,N_6585);
nand U7563 (N_7563,N_6237,N_6119);
xor U7564 (N_7564,N_6668,N_7188);
or U7565 (N_7565,N_7145,N_6876);
xor U7566 (N_7566,N_6628,N_6024);
or U7567 (N_7567,N_6158,N_6610);
and U7568 (N_7568,N_7155,N_6882);
xnor U7569 (N_7569,N_6075,N_7081);
or U7570 (N_7570,N_6458,N_6546);
or U7571 (N_7571,N_7165,N_6132);
and U7572 (N_7572,N_6216,N_6176);
xor U7573 (N_7573,N_7043,N_6092);
nor U7574 (N_7574,N_6205,N_6474);
and U7575 (N_7575,N_7088,N_6887);
nand U7576 (N_7576,N_6526,N_6814);
and U7577 (N_7577,N_7162,N_6191);
nand U7578 (N_7578,N_7122,N_6514);
xor U7579 (N_7579,N_6536,N_6612);
nand U7580 (N_7580,N_6342,N_6805);
nand U7581 (N_7581,N_7006,N_6465);
xor U7582 (N_7582,N_7039,N_6766);
and U7583 (N_7583,N_6110,N_6297);
xnor U7584 (N_7584,N_7083,N_7038);
nand U7585 (N_7585,N_6013,N_6226);
nor U7586 (N_7586,N_6313,N_6572);
and U7587 (N_7587,N_6576,N_7150);
and U7588 (N_7588,N_6733,N_6186);
and U7589 (N_7589,N_7139,N_6052);
xnor U7590 (N_7590,N_6500,N_6913);
and U7591 (N_7591,N_6118,N_6803);
nor U7592 (N_7592,N_6368,N_6480);
xnor U7593 (N_7593,N_6449,N_6695);
xor U7594 (N_7594,N_6507,N_6141);
nor U7595 (N_7595,N_6286,N_6679);
nand U7596 (N_7596,N_7181,N_6199);
and U7597 (N_7597,N_6473,N_6116);
nand U7598 (N_7598,N_6706,N_6535);
xnor U7599 (N_7599,N_6639,N_6693);
and U7600 (N_7600,N_6482,N_6204);
xor U7601 (N_7601,N_6802,N_6720);
xor U7602 (N_7602,N_6724,N_6554);
nand U7603 (N_7603,N_7096,N_6798);
nor U7604 (N_7604,N_6145,N_6792);
nand U7605 (N_7605,N_7030,N_6344);
nand U7606 (N_7606,N_6853,N_6999);
xor U7607 (N_7607,N_6910,N_6740);
nor U7608 (N_7608,N_6800,N_6021);
xnor U7609 (N_7609,N_6143,N_7087);
nor U7610 (N_7610,N_7146,N_6242);
and U7611 (N_7611,N_6607,N_6717);
xor U7612 (N_7612,N_6527,N_6026);
xnor U7613 (N_7613,N_6902,N_6874);
or U7614 (N_7614,N_6808,N_6647);
nor U7615 (N_7615,N_6129,N_6180);
nand U7616 (N_7616,N_7086,N_6839);
xor U7617 (N_7617,N_7025,N_6534);
and U7618 (N_7618,N_7142,N_6746);
nor U7619 (N_7619,N_6354,N_6202);
nand U7620 (N_7620,N_6153,N_6875);
nor U7621 (N_7621,N_6365,N_7082);
and U7622 (N_7622,N_6811,N_7192);
xor U7623 (N_7623,N_7154,N_7102);
xor U7624 (N_7624,N_6217,N_6336);
and U7625 (N_7625,N_7044,N_6415);
nand U7626 (N_7626,N_6593,N_6600);
or U7627 (N_7627,N_6362,N_7085);
xor U7628 (N_7628,N_6664,N_6060);
nor U7629 (N_7629,N_6413,N_6019);
or U7630 (N_7630,N_6959,N_6305);
xnor U7631 (N_7631,N_6027,N_6375);
xnor U7632 (N_7632,N_6670,N_6582);
or U7633 (N_7633,N_6307,N_6187);
and U7634 (N_7634,N_6520,N_6497);
and U7635 (N_7635,N_6631,N_7198);
or U7636 (N_7636,N_6207,N_6058);
and U7637 (N_7637,N_6709,N_6178);
xnor U7638 (N_7638,N_7144,N_6492);
or U7639 (N_7639,N_6768,N_6136);
or U7640 (N_7640,N_7130,N_6776);
or U7641 (N_7641,N_6409,N_6682);
and U7642 (N_7642,N_6175,N_6346);
nand U7643 (N_7643,N_6821,N_6262);
xor U7644 (N_7644,N_6868,N_6856);
nor U7645 (N_7645,N_6442,N_6671);
and U7646 (N_7646,N_6356,N_7028);
nor U7647 (N_7647,N_7059,N_6846);
nand U7648 (N_7648,N_6434,N_6751);
and U7649 (N_7649,N_6629,N_6327);
nor U7650 (N_7650,N_6955,N_6203);
nand U7651 (N_7651,N_6481,N_6489);
and U7652 (N_7652,N_6063,N_6245);
xor U7653 (N_7653,N_6188,N_6339);
xnor U7654 (N_7654,N_6192,N_6885);
xor U7655 (N_7655,N_7040,N_7058);
and U7656 (N_7656,N_6406,N_6496);
nor U7657 (N_7657,N_6040,N_7069);
and U7658 (N_7658,N_6274,N_6669);
or U7659 (N_7659,N_6722,N_6378);
nor U7660 (N_7660,N_6443,N_6320);
nor U7661 (N_7661,N_6211,N_6881);
nor U7662 (N_7662,N_6518,N_6571);
or U7663 (N_7663,N_6238,N_6986);
nor U7664 (N_7664,N_6975,N_6312);
xnor U7665 (N_7665,N_6016,N_6357);
nor U7666 (N_7666,N_6230,N_6691);
nand U7667 (N_7667,N_7076,N_6696);
nor U7668 (N_7668,N_6727,N_6782);
or U7669 (N_7669,N_7078,N_6402);
or U7670 (N_7670,N_6732,N_6246);
nor U7671 (N_7671,N_6445,N_7193);
xnor U7672 (N_7672,N_6551,N_6140);
nand U7673 (N_7673,N_7008,N_6744);
xnor U7674 (N_7674,N_6265,N_7010);
or U7675 (N_7675,N_7095,N_6133);
xnor U7676 (N_7676,N_6039,N_6681);
nor U7677 (N_7677,N_6280,N_6974);
or U7678 (N_7678,N_7024,N_6177);
nor U7679 (N_7679,N_6645,N_7108);
nand U7680 (N_7680,N_6423,N_6374);
nand U7681 (N_7681,N_6147,N_7140);
or U7682 (N_7682,N_6493,N_6525);
nand U7683 (N_7683,N_6461,N_6113);
or U7684 (N_7684,N_7022,N_6519);
nand U7685 (N_7685,N_7072,N_6635);
or U7686 (N_7686,N_6138,N_6257);
and U7687 (N_7687,N_6528,N_6807);
nor U7688 (N_7688,N_6131,N_6130);
nand U7689 (N_7689,N_6028,N_6498);
xor U7690 (N_7690,N_6545,N_6698);
and U7691 (N_7691,N_6757,N_6941);
nor U7692 (N_7692,N_6586,N_6308);
nand U7693 (N_7693,N_7106,N_6909);
nand U7694 (N_7694,N_6854,N_7033);
or U7695 (N_7695,N_6736,N_6386);
and U7696 (N_7696,N_6654,N_6859);
nor U7697 (N_7697,N_6953,N_6857);
nor U7698 (N_7698,N_6111,N_6115);
nand U7699 (N_7699,N_6193,N_7197);
or U7700 (N_7700,N_6982,N_6756);
and U7701 (N_7701,N_6611,N_6381);
nand U7702 (N_7702,N_6967,N_6090);
xor U7703 (N_7703,N_6087,N_6765);
and U7704 (N_7704,N_7037,N_7128);
or U7705 (N_7705,N_6575,N_6338);
xnor U7706 (N_7706,N_6565,N_6997);
xnor U7707 (N_7707,N_6789,N_6861);
xor U7708 (N_7708,N_6921,N_7046);
xnor U7709 (N_7709,N_6171,N_6124);
xnor U7710 (N_7710,N_6602,N_7050);
nor U7711 (N_7711,N_6427,N_7182);
and U7712 (N_7712,N_6426,N_7152);
nand U7713 (N_7713,N_7105,N_6304);
xor U7714 (N_7714,N_6460,N_6869);
nor U7715 (N_7715,N_6022,N_6573);
xnor U7716 (N_7716,N_6590,N_6858);
xnor U7717 (N_7717,N_6851,N_6155);
or U7718 (N_7718,N_6787,N_6243);
or U7719 (N_7719,N_6690,N_7171);
xor U7720 (N_7720,N_6588,N_6719);
or U7721 (N_7721,N_6453,N_6931);
nor U7722 (N_7722,N_6318,N_6441);
and U7723 (N_7723,N_6031,N_6299);
or U7724 (N_7724,N_7041,N_7007);
nor U7725 (N_7725,N_7177,N_6847);
and U7726 (N_7726,N_6912,N_6387);
and U7727 (N_7727,N_6494,N_7115);
xnor U7728 (N_7728,N_7060,N_6328);
xnor U7729 (N_7729,N_6258,N_6349);
nand U7730 (N_7730,N_6738,N_7023);
nand U7731 (N_7731,N_6531,N_6907);
xnor U7732 (N_7732,N_6828,N_7163);
or U7733 (N_7733,N_6084,N_6094);
or U7734 (N_7734,N_6817,N_6692);
nor U7735 (N_7735,N_6558,N_6579);
and U7736 (N_7736,N_6005,N_7172);
or U7737 (N_7737,N_6529,N_6154);
and U7738 (N_7738,N_6391,N_6072);
or U7739 (N_7739,N_6533,N_7074);
xnor U7740 (N_7740,N_6985,N_6728);
xor U7741 (N_7741,N_6948,N_6165);
nor U7742 (N_7742,N_6102,N_6627);
xnor U7743 (N_7743,N_6047,N_6366);
xor U7744 (N_7744,N_7143,N_7032);
and U7745 (N_7745,N_6450,N_6726);
nor U7746 (N_7746,N_6412,N_7034);
nor U7747 (N_7747,N_6466,N_7125);
or U7748 (N_7748,N_6906,N_6169);
nand U7749 (N_7749,N_6705,N_7170);
xnor U7750 (N_7750,N_7084,N_7116);
xor U7751 (N_7751,N_6159,N_6819);
nor U7752 (N_7752,N_6954,N_6081);
nor U7753 (N_7753,N_6066,N_6884);
nand U7754 (N_7754,N_6392,N_6574);
and U7755 (N_7755,N_6218,N_6167);
and U7756 (N_7756,N_6605,N_6070);
or U7757 (N_7757,N_6587,N_6069);
xor U7758 (N_7758,N_6156,N_6794);
nand U7759 (N_7759,N_6712,N_7093);
xor U7760 (N_7760,N_7127,N_6150);
xor U7761 (N_7761,N_6054,N_6229);
nor U7762 (N_7762,N_7079,N_6223);
or U7763 (N_7763,N_7097,N_7063);
nor U7764 (N_7764,N_6649,N_6976);
or U7765 (N_7765,N_6149,N_6810);
and U7766 (N_7766,N_7067,N_6638);
nor U7767 (N_7767,N_6301,N_6809);
xnor U7768 (N_7768,N_6006,N_6326);
nand U7769 (N_7769,N_7195,N_7137);
nand U7770 (N_7770,N_6091,N_6928);
and U7771 (N_7771,N_6424,N_6296);
nand U7772 (N_7772,N_6979,N_6099);
or U7773 (N_7773,N_6503,N_6411);
nand U7774 (N_7774,N_6319,N_6791);
nand U7775 (N_7775,N_6253,N_6417);
and U7776 (N_7776,N_6281,N_6430);
and U7777 (N_7777,N_6763,N_6057);
nor U7778 (N_7778,N_6677,N_6863);
or U7779 (N_7779,N_6112,N_6215);
nand U7780 (N_7780,N_6170,N_6981);
and U7781 (N_7781,N_6231,N_6240);
xor U7782 (N_7782,N_6716,N_6749);
xor U7783 (N_7783,N_6322,N_6711);
or U7784 (N_7784,N_6456,N_6033);
and U7785 (N_7785,N_6530,N_6157);
or U7786 (N_7786,N_6878,N_6394);
nor U7787 (N_7787,N_6699,N_6897);
nand U7788 (N_7788,N_6648,N_7000);
and U7789 (N_7789,N_6898,N_6947);
or U7790 (N_7790,N_6451,N_7066);
nand U7791 (N_7791,N_6444,N_6018);
nor U7792 (N_7792,N_6273,N_6825);
nor U7793 (N_7793,N_6252,N_6730);
or U7794 (N_7794,N_6731,N_6101);
or U7795 (N_7795,N_6432,N_6850);
nand U7796 (N_7796,N_6121,N_6103);
nor U7797 (N_7797,N_6352,N_7064);
and U7798 (N_7798,N_7036,N_6761);
or U7799 (N_7799,N_6929,N_6160);
xnor U7800 (N_7800,N_6277,N_6318);
xnor U7801 (N_7801,N_6414,N_6071);
nor U7802 (N_7802,N_6076,N_6408);
xor U7803 (N_7803,N_6166,N_6708);
or U7804 (N_7804,N_6187,N_6355);
or U7805 (N_7805,N_6038,N_7025);
nor U7806 (N_7806,N_6324,N_6230);
nor U7807 (N_7807,N_6975,N_6491);
nor U7808 (N_7808,N_7122,N_6866);
or U7809 (N_7809,N_6855,N_6867);
nand U7810 (N_7810,N_6589,N_6923);
nor U7811 (N_7811,N_6334,N_6299);
nand U7812 (N_7812,N_6125,N_7010);
or U7813 (N_7813,N_7092,N_6709);
and U7814 (N_7814,N_6793,N_6256);
xnor U7815 (N_7815,N_6038,N_7175);
and U7816 (N_7816,N_6112,N_6890);
or U7817 (N_7817,N_7096,N_6035);
nor U7818 (N_7818,N_7176,N_7140);
or U7819 (N_7819,N_6401,N_6623);
nand U7820 (N_7820,N_6414,N_6758);
nand U7821 (N_7821,N_6969,N_6392);
or U7822 (N_7822,N_6767,N_6955);
nand U7823 (N_7823,N_6339,N_6539);
and U7824 (N_7824,N_6725,N_7037);
or U7825 (N_7825,N_6267,N_6395);
nand U7826 (N_7826,N_6301,N_6559);
xnor U7827 (N_7827,N_6668,N_6747);
xor U7828 (N_7828,N_6109,N_6878);
nand U7829 (N_7829,N_7199,N_6038);
and U7830 (N_7830,N_6090,N_6845);
nor U7831 (N_7831,N_6330,N_6934);
nand U7832 (N_7832,N_6713,N_6711);
nand U7833 (N_7833,N_6769,N_6860);
nor U7834 (N_7834,N_6851,N_7163);
nand U7835 (N_7835,N_7193,N_6751);
and U7836 (N_7836,N_6488,N_6340);
or U7837 (N_7837,N_6318,N_7009);
xor U7838 (N_7838,N_6276,N_7175);
nand U7839 (N_7839,N_7093,N_6896);
or U7840 (N_7840,N_6259,N_6010);
nor U7841 (N_7841,N_6735,N_6622);
xor U7842 (N_7842,N_7110,N_6679);
nor U7843 (N_7843,N_6665,N_6281);
or U7844 (N_7844,N_6718,N_6443);
nand U7845 (N_7845,N_6818,N_6038);
nor U7846 (N_7846,N_6155,N_6578);
xor U7847 (N_7847,N_7077,N_6114);
and U7848 (N_7848,N_6502,N_6870);
nand U7849 (N_7849,N_6718,N_6665);
or U7850 (N_7850,N_7049,N_6740);
xor U7851 (N_7851,N_6635,N_7044);
xor U7852 (N_7852,N_6633,N_6435);
or U7853 (N_7853,N_6263,N_7119);
nand U7854 (N_7854,N_6219,N_7027);
or U7855 (N_7855,N_6860,N_6369);
and U7856 (N_7856,N_7106,N_6368);
nor U7857 (N_7857,N_7049,N_7069);
and U7858 (N_7858,N_6506,N_7153);
xnor U7859 (N_7859,N_6873,N_6560);
xnor U7860 (N_7860,N_6662,N_6373);
or U7861 (N_7861,N_7191,N_6276);
xnor U7862 (N_7862,N_6200,N_7143);
or U7863 (N_7863,N_6169,N_6192);
and U7864 (N_7864,N_6614,N_6937);
and U7865 (N_7865,N_6902,N_6884);
or U7866 (N_7866,N_6725,N_6498);
nor U7867 (N_7867,N_6472,N_7194);
nand U7868 (N_7868,N_6704,N_6976);
xnor U7869 (N_7869,N_6499,N_7179);
or U7870 (N_7870,N_7143,N_6187);
nor U7871 (N_7871,N_6197,N_6810);
or U7872 (N_7872,N_6426,N_6852);
nor U7873 (N_7873,N_6658,N_6428);
and U7874 (N_7874,N_6489,N_6580);
nor U7875 (N_7875,N_6836,N_6560);
or U7876 (N_7876,N_6039,N_6619);
xor U7877 (N_7877,N_6964,N_7161);
nor U7878 (N_7878,N_7190,N_6454);
and U7879 (N_7879,N_6113,N_6167);
xnor U7880 (N_7880,N_6110,N_6734);
xnor U7881 (N_7881,N_6593,N_6913);
xnor U7882 (N_7882,N_6898,N_6668);
xnor U7883 (N_7883,N_6869,N_6323);
or U7884 (N_7884,N_7039,N_6360);
and U7885 (N_7885,N_7194,N_7185);
or U7886 (N_7886,N_6953,N_6665);
xor U7887 (N_7887,N_6775,N_6273);
and U7888 (N_7888,N_6888,N_6167);
xor U7889 (N_7889,N_7014,N_7006);
or U7890 (N_7890,N_6117,N_6206);
xor U7891 (N_7891,N_6000,N_6824);
xnor U7892 (N_7892,N_6276,N_7093);
xor U7893 (N_7893,N_6318,N_6384);
nor U7894 (N_7894,N_6658,N_6251);
nor U7895 (N_7895,N_6678,N_6604);
and U7896 (N_7896,N_6945,N_6288);
xor U7897 (N_7897,N_6037,N_6017);
xor U7898 (N_7898,N_6472,N_6600);
or U7899 (N_7899,N_6312,N_7088);
and U7900 (N_7900,N_6512,N_6874);
or U7901 (N_7901,N_7036,N_6111);
nand U7902 (N_7902,N_6893,N_7026);
nand U7903 (N_7903,N_6505,N_6879);
or U7904 (N_7904,N_6958,N_6701);
nand U7905 (N_7905,N_6127,N_7146);
xor U7906 (N_7906,N_6224,N_6704);
and U7907 (N_7907,N_6925,N_6153);
and U7908 (N_7908,N_7184,N_6695);
or U7909 (N_7909,N_6547,N_6578);
xnor U7910 (N_7910,N_6530,N_6864);
or U7911 (N_7911,N_6616,N_6901);
nand U7912 (N_7912,N_7053,N_7181);
nand U7913 (N_7913,N_6004,N_6565);
xnor U7914 (N_7914,N_6489,N_7179);
and U7915 (N_7915,N_6848,N_6491);
xnor U7916 (N_7916,N_6507,N_6411);
nor U7917 (N_7917,N_6738,N_6339);
nor U7918 (N_7918,N_6318,N_6868);
or U7919 (N_7919,N_7159,N_6367);
and U7920 (N_7920,N_6950,N_6285);
nand U7921 (N_7921,N_6076,N_7053);
and U7922 (N_7922,N_6996,N_6030);
or U7923 (N_7923,N_6557,N_6825);
nor U7924 (N_7924,N_6726,N_6232);
or U7925 (N_7925,N_6878,N_6378);
xnor U7926 (N_7926,N_6257,N_6339);
nand U7927 (N_7927,N_6414,N_6334);
or U7928 (N_7928,N_6693,N_6963);
xnor U7929 (N_7929,N_6967,N_6390);
nand U7930 (N_7930,N_6328,N_7198);
nand U7931 (N_7931,N_6813,N_6784);
or U7932 (N_7932,N_6743,N_6645);
or U7933 (N_7933,N_6270,N_6909);
xor U7934 (N_7934,N_7195,N_6727);
nand U7935 (N_7935,N_6132,N_7155);
and U7936 (N_7936,N_6767,N_6344);
nand U7937 (N_7937,N_6126,N_7159);
xor U7938 (N_7938,N_6294,N_6752);
xnor U7939 (N_7939,N_6001,N_6417);
and U7940 (N_7940,N_6273,N_6248);
nor U7941 (N_7941,N_6619,N_6516);
xor U7942 (N_7942,N_6486,N_6630);
and U7943 (N_7943,N_6910,N_6259);
and U7944 (N_7944,N_7144,N_6769);
and U7945 (N_7945,N_7133,N_6206);
xor U7946 (N_7946,N_6976,N_6898);
xor U7947 (N_7947,N_6904,N_6401);
nand U7948 (N_7948,N_6925,N_6452);
xor U7949 (N_7949,N_6549,N_6120);
xor U7950 (N_7950,N_6525,N_6572);
nor U7951 (N_7951,N_7070,N_6147);
or U7952 (N_7952,N_6749,N_6405);
xor U7953 (N_7953,N_6163,N_7033);
and U7954 (N_7954,N_6133,N_6077);
or U7955 (N_7955,N_6940,N_6726);
nor U7956 (N_7956,N_7135,N_6260);
xor U7957 (N_7957,N_6019,N_6634);
nor U7958 (N_7958,N_6342,N_6508);
nor U7959 (N_7959,N_6880,N_6784);
nor U7960 (N_7960,N_6372,N_7142);
xnor U7961 (N_7961,N_6011,N_6182);
and U7962 (N_7962,N_6224,N_6391);
nand U7963 (N_7963,N_6083,N_6292);
and U7964 (N_7964,N_6907,N_6814);
or U7965 (N_7965,N_6897,N_6346);
nor U7966 (N_7966,N_6626,N_6540);
nor U7967 (N_7967,N_6618,N_6957);
nand U7968 (N_7968,N_7175,N_7026);
or U7969 (N_7969,N_6504,N_6318);
nand U7970 (N_7970,N_6223,N_6560);
nand U7971 (N_7971,N_6991,N_6528);
nor U7972 (N_7972,N_6977,N_6967);
nor U7973 (N_7973,N_6091,N_6766);
nand U7974 (N_7974,N_7051,N_6196);
xnor U7975 (N_7975,N_7163,N_6978);
xor U7976 (N_7976,N_6513,N_6967);
nand U7977 (N_7977,N_6983,N_6170);
nand U7978 (N_7978,N_6073,N_6648);
or U7979 (N_7979,N_6669,N_7024);
nand U7980 (N_7980,N_6864,N_6480);
nor U7981 (N_7981,N_6804,N_6180);
nor U7982 (N_7982,N_6590,N_6962);
xor U7983 (N_7983,N_6404,N_6050);
xor U7984 (N_7984,N_6956,N_6230);
xnor U7985 (N_7985,N_6875,N_6304);
nand U7986 (N_7986,N_6131,N_6183);
nor U7987 (N_7987,N_7126,N_6231);
nor U7988 (N_7988,N_6164,N_6533);
or U7989 (N_7989,N_6604,N_6921);
nand U7990 (N_7990,N_6354,N_6915);
nand U7991 (N_7991,N_7021,N_6164);
or U7992 (N_7992,N_7147,N_7079);
or U7993 (N_7993,N_6325,N_6990);
xor U7994 (N_7994,N_6880,N_6187);
or U7995 (N_7995,N_6017,N_6382);
and U7996 (N_7996,N_6246,N_7077);
xnor U7997 (N_7997,N_7180,N_7179);
and U7998 (N_7998,N_6930,N_6576);
or U7999 (N_7999,N_6953,N_6341);
nor U8000 (N_8000,N_6317,N_6219);
and U8001 (N_8001,N_6452,N_6879);
nor U8002 (N_8002,N_6965,N_6410);
and U8003 (N_8003,N_6227,N_6266);
nor U8004 (N_8004,N_7178,N_6472);
or U8005 (N_8005,N_6817,N_6787);
or U8006 (N_8006,N_7159,N_7024);
xnor U8007 (N_8007,N_6351,N_6605);
nor U8008 (N_8008,N_6428,N_6072);
xnor U8009 (N_8009,N_6577,N_6190);
and U8010 (N_8010,N_6723,N_6087);
and U8011 (N_8011,N_6784,N_6398);
nor U8012 (N_8012,N_6200,N_6715);
xnor U8013 (N_8013,N_6950,N_6215);
xnor U8014 (N_8014,N_6229,N_6169);
nor U8015 (N_8015,N_6687,N_6023);
and U8016 (N_8016,N_6043,N_6434);
xnor U8017 (N_8017,N_6024,N_7157);
xor U8018 (N_8018,N_7035,N_6360);
nand U8019 (N_8019,N_6150,N_6238);
and U8020 (N_8020,N_7090,N_6898);
nand U8021 (N_8021,N_7098,N_6615);
xor U8022 (N_8022,N_6195,N_7010);
xnor U8023 (N_8023,N_6093,N_6816);
nor U8024 (N_8024,N_6110,N_6495);
nand U8025 (N_8025,N_6746,N_7060);
xnor U8026 (N_8026,N_6355,N_6224);
and U8027 (N_8027,N_6798,N_6290);
and U8028 (N_8028,N_6385,N_6768);
nand U8029 (N_8029,N_6963,N_7152);
and U8030 (N_8030,N_6013,N_6411);
xnor U8031 (N_8031,N_6896,N_6748);
xnor U8032 (N_8032,N_6032,N_6571);
or U8033 (N_8033,N_6997,N_6979);
or U8034 (N_8034,N_6574,N_7087);
or U8035 (N_8035,N_6641,N_6709);
xor U8036 (N_8036,N_7064,N_6685);
and U8037 (N_8037,N_6046,N_6837);
xnor U8038 (N_8038,N_6430,N_6554);
nor U8039 (N_8039,N_6019,N_6116);
nor U8040 (N_8040,N_6710,N_6839);
nand U8041 (N_8041,N_6200,N_6975);
or U8042 (N_8042,N_6697,N_7184);
xor U8043 (N_8043,N_6488,N_7105);
and U8044 (N_8044,N_6717,N_6137);
nor U8045 (N_8045,N_6979,N_6136);
or U8046 (N_8046,N_6417,N_6022);
and U8047 (N_8047,N_6399,N_6756);
and U8048 (N_8048,N_7071,N_6075);
and U8049 (N_8049,N_7119,N_6478);
and U8050 (N_8050,N_6819,N_6742);
nor U8051 (N_8051,N_6145,N_7129);
nand U8052 (N_8052,N_7068,N_7081);
nand U8053 (N_8053,N_6702,N_6872);
nor U8054 (N_8054,N_6810,N_7173);
or U8055 (N_8055,N_7149,N_7062);
nor U8056 (N_8056,N_6119,N_6891);
nor U8057 (N_8057,N_7124,N_7148);
nand U8058 (N_8058,N_6186,N_6299);
or U8059 (N_8059,N_7135,N_6405);
nand U8060 (N_8060,N_7109,N_6704);
xor U8061 (N_8061,N_6950,N_7111);
nand U8062 (N_8062,N_6241,N_6390);
nor U8063 (N_8063,N_7096,N_6940);
nor U8064 (N_8064,N_6530,N_6456);
nand U8065 (N_8065,N_6567,N_6145);
nor U8066 (N_8066,N_6088,N_7069);
and U8067 (N_8067,N_7110,N_6828);
xnor U8068 (N_8068,N_6232,N_6641);
or U8069 (N_8069,N_7199,N_6423);
nor U8070 (N_8070,N_6345,N_6662);
nand U8071 (N_8071,N_6384,N_7098);
or U8072 (N_8072,N_7118,N_6821);
nand U8073 (N_8073,N_6348,N_7165);
and U8074 (N_8074,N_6515,N_7159);
xor U8075 (N_8075,N_6853,N_6991);
xor U8076 (N_8076,N_6775,N_7175);
nor U8077 (N_8077,N_6436,N_6423);
or U8078 (N_8078,N_6993,N_6014);
or U8079 (N_8079,N_7154,N_6157);
nor U8080 (N_8080,N_7159,N_6419);
or U8081 (N_8081,N_6146,N_6992);
and U8082 (N_8082,N_6557,N_6182);
nor U8083 (N_8083,N_7042,N_7047);
and U8084 (N_8084,N_6635,N_6917);
nand U8085 (N_8085,N_6849,N_6421);
or U8086 (N_8086,N_6174,N_6759);
xnor U8087 (N_8087,N_6758,N_6377);
or U8088 (N_8088,N_6113,N_6571);
nor U8089 (N_8089,N_7118,N_6182);
and U8090 (N_8090,N_6995,N_6679);
or U8091 (N_8091,N_6398,N_6820);
and U8092 (N_8092,N_6111,N_6526);
nor U8093 (N_8093,N_6476,N_6473);
or U8094 (N_8094,N_6570,N_6465);
nand U8095 (N_8095,N_6421,N_6859);
and U8096 (N_8096,N_7056,N_6355);
or U8097 (N_8097,N_7058,N_6328);
or U8098 (N_8098,N_6334,N_6395);
nand U8099 (N_8099,N_6582,N_6413);
nand U8100 (N_8100,N_6112,N_7068);
nor U8101 (N_8101,N_7071,N_6703);
nor U8102 (N_8102,N_6204,N_6560);
or U8103 (N_8103,N_6743,N_6335);
or U8104 (N_8104,N_6397,N_6903);
and U8105 (N_8105,N_6132,N_6165);
and U8106 (N_8106,N_6742,N_7035);
xnor U8107 (N_8107,N_6015,N_6388);
nor U8108 (N_8108,N_6464,N_6748);
nand U8109 (N_8109,N_6413,N_6559);
nand U8110 (N_8110,N_6056,N_6686);
or U8111 (N_8111,N_7143,N_7119);
xnor U8112 (N_8112,N_7083,N_6074);
nand U8113 (N_8113,N_6085,N_7196);
nand U8114 (N_8114,N_6283,N_6265);
and U8115 (N_8115,N_6070,N_7142);
nor U8116 (N_8116,N_6304,N_7057);
and U8117 (N_8117,N_6116,N_7191);
nand U8118 (N_8118,N_6313,N_7132);
nand U8119 (N_8119,N_6041,N_6996);
xor U8120 (N_8120,N_7145,N_6063);
or U8121 (N_8121,N_6378,N_6208);
nor U8122 (N_8122,N_6821,N_6370);
and U8123 (N_8123,N_6122,N_6509);
nand U8124 (N_8124,N_6429,N_6423);
xor U8125 (N_8125,N_7108,N_6210);
xor U8126 (N_8126,N_6260,N_6180);
nor U8127 (N_8127,N_6324,N_7071);
nor U8128 (N_8128,N_6635,N_6089);
and U8129 (N_8129,N_6187,N_6632);
nor U8130 (N_8130,N_6657,N_6932);
nand U8131 (N_8131,N_6831,N_6475);
nor U8132 (N_8132,N_6726,N_6140);
or U8133 (N_8133,N_6821,N_7098);
nor U8134 (N_8134,N_6904,N_6315);
xor U8135 (N_8135,N_6486,N_6497);
xnor U8136 (N_8136,N_6351,N_6449);
and U8137 (N_8137,N_6668,N_6871);
nand U8138 (N_8138,N_6141,N_6648);
or U8139 (N_8139,N_6106,N_6744);
xor U8140 (N_8140,N_6234,N_6802);
nand U8141 (N_8141,N_6633,N_7123);
or U8142 (N_8142,N_6318,N_6115);
nor U8143 (N_8143,N_6681,N_6789);
and U8144 (N_8144,N_6110,N_6350);
nand U8145 (N_8145,N_6661,N_6634);
or U8146 (N_8146,N_6523,N_6805);
or U8147 (N_8147,N_6398,N_6894);
nand U8148 (N_8148,N_6774,N_7199);
xor U8149 (N_8149,N_6879,N_6357);
or U8150 (N_8150,N_6506,N_6869);
and U8151 (N_8151,N_6869,N_6495);
and U8152 (N_8152,N_7051,N_6303);
xor U8153 (N_8153,N_6591,N_6429);
nand U8154 (N_8154,N_6118,N_6995);
nor U8155 (N_8155,N_6928,N_6642);
nand U8156 (N_8156,N_6470,N_6452);
or U8157 (N_8157,N_6492,N_6308);
or U8158 (N_8158,N_7007,N_7166);
xnor U8159 (N_8159,N_6595,N_6758);
and U8160 (N_8160,N_7170,N_6682);
and U8161 (N_8161,N_6939,N_6028);
and U8162 (N_8162,N_6334,N_6556);
or U8163 (N_8163,N_6796,N_6242);
nor U8164 (N_8164,N_6689,N_6303);
nand U8165 (N_8165,N_6459,N_6256);
nor U8166 (N_8166,N_7028,N_6165);
nand U8167 (N_8167,N_6725,N_6934);
nand U8168 (N_8168,N_7131,N_6249);
nand U8169 (N_8169,N_6412,N_6913);
nor U8170 (N_8170,N_7100,N_6162);
xor U8171 (N_8171,N_7070,N_6180);
nand U8172 (N_8172,N_6788,N_6936);
xor U8173 (N_8173,N_6349,N_6136);
xor U8174 (N_8174,N_6554,N_6487);
xor U8175 (N_8175,N_6237,N_6620);
xor U8176 (N_8176,N_6839,N_7136);
nor U8177 (N_8177,N_6155,N_6361);
or U8178 (N_8178,N_7035,N_6082);
or U8179 (N_8179,N_6420,N_7185);
or U8180 (N_8180,N_6797,N_6967);
nand U8181 (N_8181,N_6815,N_6652);
nor U8182 (N_8182,N_6591,N_6779);
nor U8183 (N_8183,N_7028,N_6934);
xnor U8184 (N_8184,N_6586,N_6108);
nand U8185 (N_8185,N_6525,N_6097);
or U8186 (N_8186,N_7169,N_6704);
xor U8187 (N_8187,N_6184,N_7146);
or U8188 (N_8188,N_6099,N_6130);
or U8189 (N_8189,N_6222,N_6538);
nor U8190 (N_8190,N_6571,N_6425);
nor U8191 (N_8191,N_6068,N_6471);
and U8192 (N_8192,N_6986,N_6152);
and U8193 (N_8193,N_6016,N_6978);
nand U8194 (N_8194,N_6419,N_6147);
nand U8195 (N_8195,N_6771,N_6157);
nand U8196 (N_8196,N_6697,N_6730);
nor U8197 (N_8197,N_6510,N_6615);
or U8198 (N_8198,N_6329,N_6646);
or U8199 (N_8199,N_6166,N_7117);
or U8200 (N_8200,N_6750,N_6991);
xnor U8201 (N_8201,N_6786,N_6685);
and U8202 (N_8202,N_6829,N_6929);
nor U8203 (N_8203,N_6219,N_6829);
nor U8204 (N_8204,N_6823,N_6442);
xnor U8205 (N_8205,N_6361,N_6804);
and U8206 (N_8206,N_6741,N_6368);
or U8207 (N_8207,N_6971,N_7121);
and U8208 (N_8208,N_6163,N_6859);
nand U8209 (N_8209,N_6641,N_6169);
or U8210 (N_8210,N_6105,N_6002);
nor U8211 (N_8211,N_6323,N_6624);
nand U8212 (N_8212,N_6076,N_6851);
nand U8213 (N_8213,N_6806,N_7147);
nor U8214 (N_8214,N_6634,N_6723);
nor U8215 (N_8215,N_7179,N_6939);
or U8216 (N_8216,N_6305,N_6796);
nand U8217 (N_8217,N_6125,N_6155);
nand U8218 (N_8218,N_6434,N_6389);
and U8219 (N_8219,N_7168,N_7070);
xor U8220 (N_8220,N_6674,N_6498);
nor U8221 (N_8221,N_7109,N_7152);
nor U8222 (N_8222,N_6338,N_7180);
nand U8223 (N_8223,N_6787,N_6881);
nor U8224 (N_8224,N_6763,N_6181);
and U8225 (N_8225,N_6398,N_6445);
and U8226 (N_8226,N_6173,N_7106);
and U8227 (N_8227,N_6674,N_6450);
xnor U8228 (N_8228,N_6151,N_6571);
nand U8229 (N_8229,N_6031,N_6013);
nor U8230 (N_8230,N_7159,N_7014);
and U8231 (N_8231,N_7194,N_6336);
nor U8232 (N_8232,N_6374,N_6734);
and U8233 (N_8233,N_6607,N_6812);
nand U8234 (N_8234,N_6874,N_6029);
or U8235 (N_8235,N_7142,N_6535);
and U8236 (N_8236,N_6502,N_6045);
or U8237 (N_8237,N_6514,N_6470);
nor U8238 (N_8238,N_6109,N_6620);
xor U8239 (N_8239,N_6581,N_7126);
xnor U8240 (N_8240,N_6803,N_6553);
xnor U8241 (N_8241,N_6242,N_7140);
nand U8242 (N_8242,N_6637,N_6634);
nand U8243 (N_8243,N_6824,N_6489);
xor U8244 (N_8244,N_6028,N_6155);
xnor U8245 (N_8245,N_6889,N_6124);
xor U8246 (N_8246,N_6875,N_6518);
xor U8247 (N_8247,N_7029,N_6664);
nor U8248 (N_8248,N_6294,N_6353);
or U8249 (N_8249,N_6568,N_6440);
and U8250 (N_8250,N_6180,N_6675);
xnor U8251 (N_8251,N_6654,N_6014);
xnor U8252 (N_8252,N_6141,N_6912);
xnor U8253 (N_8253,N_6094,N_6238);
xor U8254 (N_8254,N_6133,N_6142);
nand U8255 (N_8255,N_6932,N_6858);
xor U8256 (N_8256,N_6166,N_6838);
xor U8257 (N_8257,N_6769,N_6564);
and U8258 (N_8258,N_7131,N_6633);
or U8259 (N_8259,N_6830,N_6267);
and U8260 (N_8260,N_6513,N_6565);
or U8261 (N_8261,N_6216,N_6004);
or U8262 (N_8262,N_7179,N_6659);
nand U8263 (N_8263,N_6773,N_6211);
nor U8264 (N_8264,N_6613,N_6186);
xnor U8265 (N_8265,N_6191,N_6610);
and U8266 (N_8266,N_6468,N_6997);
nand U8267 (N_8267,N_6621,N_6797);
or U8268 (N_8268,N_6458,N_6196);
nor U8269 (N_8269,N_6021,N_6972);
nand U8270 (N_8270,N_6763,N_6192);
nand U8271 (N_8271,N_6378,N_6116);
and U8272 (N_8272,N_6131,N_6884);
and U8273 (N_8273,N_6567,N_7039);
or U8274 (N_8274,N_6491,N_6035);
and U8275 (N_8275,N_6895,N_7041);
and U8276 (N_8276,N_6471,N_6819);
or U8277 (N_8277,N_7070,N_6869);
nand U8278 (N_8278,N_6916,N_6788);
xnor U8279 (N_8279,N_7150,N_6879);
and U8280 (N_8280,N_6557,N_6639);
nand U8281 (N_8281,N_6928,N_6956);
or U8282 (N_8282,N_6477,N_6463);
nand U8283 (N_8283,N_6816,N_7050);
and U8284 (N_8284,N_6122,N_6663);
or U8285 (N_8285,N_6479,N_6815);
xnor U8286 (N_8286,N_6722,N_6163);
nor U8287 (N_8287,N_6227,N_6055);
nand U8288 (N_8288,N_6588,N_6548);
nand U8289 (N_8289,N_6441,N_6277);
and U8290 (N_8290,N_6827,N_6041);
nor U8291 (N_8291,N_6092,N_6237);
xnor U8292 (N_8292,N_6142,N_7187);
nand U8293 (N_8293,N_6537,N_6587);
or U8294 (N_8294,N_6694,N_6312);
nand U8295 (N_8295,N_6958,N_6193);
or U8296 (N_8296,N_6961,N_6404);
nand U8297 (N_8297,N_7123,N_6599);
or U8298 (N_8298,N_6798,N_6108);
and U8299 (N_8299,N_6698,N_7076);
and U8300 (N_8300,N_6290,N_6585);
nor U8301 (N_8301,N_6242,N_6108);
and U8302 (N_8302,N_6255,N_6040);
xor U8303 (N_8303,N_6350,N_6517);
xor U8304 (N_8304,N_6969,N_6197);
nand U8305 (N_8305,N_6659,N_6038);
nor U8306 (N_8306,N_6265,N_7078);
or U8307 (N_8307,N_6272,N_6135);
or U8308 (N_8308,N_6635,N_6693);
nor U8309 (N_8309,N_6924,N_6154);
nor U8310 (N_8310,N_6811,N_7060);
nor U8311 (N_8311,N_7035,N_6888);
or U8312 (N_8312,N_6175,N_6319);
xor U8313 (N_8313,N_7161,N_6319);
nand U8314 (N_8314,N_6738,N_6914);
xnor U8315 (N_8315,N_6835,N_6179);
and U8316 (N_8316,N_6754,N_6743);
xor U8317 (N_8317,N_6471,N_6687);
or U8318 (N_8318,N_6233,N_6206);
nor U8319 (N_8319,N_6881,N_6525);
and U8320 (N_8320,N_7168,N_6176);
and U8321 (N_8321,N_6083,N_6502);
and U8322 (N_8322,N_7078,N_7119);
or U8323 (N_8323,N_7058,N_6586);
or U8324 (N_8324,N_6242,N_6797);
or U8325 (N_8325,N_6316,N_6928);
or U8326 (N_8326,N_6589,N_6400);
and U8327 (N_8327,N_6364,N_6972);
or U8328 (N_8328,N_6328,N_6340);
or U8329 (N_8329,N_6323,N_6221);
and U8330 (N_8330,N_6048,N_6786);
and U8331 (N_8331,N_6944,N_6729);
and U8332 (N_8332,N_6214,N_6156);
nand U8333 (N_8333,N_7107,N_7025);
or U8334 (N_8334,N_6408,N_6772);
xnor U8335 (N_8335,N_6159,N_6976);
nor U8336 (N_8336,N_6887,N_6285);
xor U8337 (N_8337,N_7002,N_6801);
nor U8338 (N_8338,N_6215,N_6545);
nand U8339 (N_8339,N_6496,N_6724);
nor U8340 (N_8340,N_6261,N_7046);
xnor U8341 (N_8341,N_6939,N_7119);
xnor U8342 (N_8342,N_6256,N_6588);
nand U8343 (N_8343,N_6877,N_6842);
or U8344 (N_8344,N_6209,N_6376);
xor U8345 (N_8345,N_6269,N_6223);
or U8346 (N_8346,N_6335,N_6530);
xnor U8347 (N_8347,N_7101,N_6030);
nor U8348 (N_8348,N_7087,N_7121);
and U8349 (N_8349,N_6324,N_6308);
or U8350 (N_8350,N_6168,N_6580);
and U8351 (N_8351,N_7040,N_6854);
or U8352 (N_8352,N_6584,N_7103);
nand U8353 (N_8353,N_6712,N_6526);
nor U8354 (N_8354,N_6544,N_6359);
nor U8355 (N_8355,N_6964,N_6667);
and U8356 (N_8356,N_6154,N_6018);
or U8357 (N_8357,N_6974,N_6312);
xor U8358 (N_8358,N_6298,N_6820);
nand U8359 (N_8359,N_6047,N_6316);
or U8360 (N_8360,N_6852,N_6881);
nand U8361 (N_8361,N_6539,N_6388);
nand U8362 (N_8362,N_6001,N_6179);
nor U8363 (N_8363,N_6783,N_6119);
nor U8364 (N_8364,N_6838,N_6093);
nand U8365 (N_8365,N_6560,N_6001);
xor U8366 (N_8366,N_6480,N_6023);
and U8367 (N_8367,N_6773,N_6594);
xor U8368 (N_8368,N_6609,N_6530);
and U8369 (N_8369,N_6536,N_6726);
nor U8370 (N_8370,N_6095,N_6628);
nor U8371 (N_8371,N_6818,N_6593);
and U8372 (N_8372,N_6261,N_6495);
xnor U8373 (N_8373,N_7093,N_6734);
nor U8374 (N_8374,N_6602,N_6741);
nand U8375 (N_8375,N_6402,N_6374);
xor U8376 (N_8376,N_7184,N_7109);
or U8377 (N_8377,N_6903,N_6175);
xnor U8378 (N_8378,N_6798,N_6092);
and U8379 (N_8379,N_6237,N_6936);
and U8380 (N_8380,N_6439,N_6899);
nor U8381 (N_8381,N_6424,N_6254);
nand U8382 (N_8382,N_6608,N_7176);
nor U8383 (N_8383,N_6687,N_6966);
and U8384 (N_8384,N_6724,N_6238);
xnor U8385 (N_8385,N_6588,N_6007);
xor U8386 (N_8386,N_6137,N_6038);
or U8387 (N_8387,N_6550,N_6019);
nor U8388 (N_8388,N_6924,N_6059);
or U8389 (N_8389,N_6179,N_6748);
nand U8390 (N_8390,N_6577,N_6665);
nor U8391 (N_8391,N_6882,N_6428);
or U8392 (N_8392,N_6380,N_6758);
or U8393 (N_8393,N_6792,N_6012);
nand U8394 (N_8394,N_6248,N_6637);
nand U8395 (N_8395,N_6091,N_6242);
nand U8396 (N_8396,N_7076,N_7047);
and U8397 (N_8397,N_6918,N_6551);
xor U8398 (N_8398,N_7012,N_7010);
nand U8399 (N_8399,N_7082,N_6414);
and U8400 (N_8400,N_8306,N_7914);
xnor U8401 (N_8401,N_7554,N_7790);
xnor U8402 (N_8402,N_7797,N_7411);
xnor U8403 (N_8403,N_8181,N_7686);
and U8404 (N_8404,N_7526,N_8278);
nor U8405 (N_8405,N_7284,N_7532);
or U8406 (N_8406,N_8310,N_7991);
or U8407 (N_8407,N_7353,N_7871);
nand U8408 (N_8408,N_8084,N_8198);
nor U8409 (N_8409,N_7855,N_8206);
nor U8410 (N_8410,N_7595,N_8060);
xnor U8411 (N_8411,N_7350,N_8133);
nor U8412 (N_8412,N_7715,N_7470);
or U8413 (N_8413,N_8257,N_7947);
and U8414 (N_8414,N_7872,N_7606);
xor U8415 (N_8415,N_8040,N_8345);
nand U8416 (N_8416,N_7419,N_7234);
nand U8417 (N_8417,N_7624,N_8151);
or U8418 (N_8418,N_7553,N_8081);
nand U8419 (N_8419,N_7431,N_7250);
nand U8420 (N_8420,N_7985,N_8317);
and U8421 (N_8421,N_7308,N_7471);
nor U8422 (N_8422,N_7934,N_7734);
and U8423 (N_8423,N_7774,N_7717);
nor U8424 (N_8424,N_7255,N_8245);
xnor U8425 (N_8425,N_7481,N_7748);
and U8426 (N_8426,N_7395,N_7220);
nand U8427 (N_8427,N_7227,N_7927);
nand U8428 (N_8428,N_7360,N_7362);
nor U8429 (N_8429,N_7848,N_7408);
and U8430 (N_8430,N_7887,N_7257);
and U8431 (N_8431,N_8279,N_7815);
nor U8432 (N_8432,N_7915,N_7476);
xor U8433 (N_8433,N_8383,N_8064);
xnor U8434 (N_8434,N_7657,N_7544);
nor U8435 (N_8435,N_7586,N_8185);
xor U8436 (N_8436,N_7499,N_7254);
nand U8437 (N_8437,N_8126,N_8372);
nand U8438 (N_8438,N_7432,N_7484);
nor U8439 (N_8439,N_7824,N_8395);
xnor U8440 (N_8440,N_7922,N_7373);
xor U8441 (N_8441,N_8046,N_8124);
or U8442 (N_8442,N_7518,N_7549);
nand U8443 (N_8443,N_8218,N_7733);
nor U8444 (N_8444,N_7273,N_7483);
xor U8445 (N_8445,N_7442,N_8015);
nor U8446 (N_8446,N_7631,N_7956);
nor U8447 (N_8447,N_7698,N_8009);
nor U8448 (N_8448,N_7520,N_7916);
or U8449 (N_8449,N_7929,N_7955);
and U8450 (N_8450,N_7325,N_7712);
or U8451 (N_8451,N_8076,N_8073);
nand U8452 (N_8452,N_8136,N_7832);
or U8453 (N_8453,N_7923,N_8051);
nand U8454 (N_8454,N_8183,N_7679);
nor U8455 (N_8455,N_7519,N_7806);
and U8456 (N_8456,N_7541,N_7901);
and U8457 (N_8457,N_7959,N_7286);
or U8458 (N_8458,N_7893,N_7641);
nor U8459 (N_8459,N_7556,N_8280);
or U8460 (N_8460,N_7275,N_7473);
nand U8461 (N_8461,N_8252,N_7448);
and U8462 (N_8462,N_8269,N_7665);
and U8463 (N_8463,N_8058,N_7575);
nand U8464 (N_8464,N_7397,N_8347);
and U8465 (N_8465,N_7217,N_7512);
and U8466 (N_8466,N_8026,N_7233);
xor U8467 (N_8467,N_7905,N_8338);
xor U8468 (N_8468,N_8371,N_7767);
xnor U8469 (N_8469,N_8361,N_7844);
or U8470 (N_8470,N_8139,N_7493);
nand U8471 (N_8471,N_8030,N_7917);
nand U8472 (N_8472,N_7266,N_7632);
and U8473 (N_8473,N_8061,N_7913);
or U8474 (N_8474,N_8128,N_7455);
xor U8475 (N_8475,N_7762,N_7332);
nand U8476 (N_8476,N_7351,N_8260);
and U8477 (N_8477,N_8219,N_7691);
and U8478 (N_8478,N_7640,N_7629);
or U8479 (N_8479,N_7772,N_7405);
nand U8480 (N_8480,N_8357,N_7634);
or U8481 (N_8481,N_7576,N_7439);
nand U8482 (N_8482,N_8131,N_7709);
or U8483 (N_8483,N_7625,N_7542);
or U8484 (N_8484,N_7794,N_7999);
and U8485 (N_8485,N_7755,N_8158);
xnor U8486 (N_8486,N_7201,N_7636);
and U8487 (N_8487,N_7357,N_7881);
xor U8488 (N_8488,N_8164,N_7445);
nor U8489 (N_8489,N_7638,N_7642);
nand U8490 (N_8490,N_7465,N_7875);
and U8491 (N_8491,N_7823,N_8167);
xor U8492 (N_8492,N_8069,N_7472);
xnor U8493 (N_8493,N_8171,N_8399);
nor U8494 (N_8494,N_8077,N_7944);
xor U8495 (N_8495,N_8297,N_8014);
nor U8496 (N_8496,N_7530,N_7215);
and U8497 (N_8497,N_7510,N_7525);
nor U8498 (N_8498,N_7851,N_7643);
nand U8499 (N_8499,N_7718,N_8224);
nor U8500 (N_8500,N_7782,N_8266);
or U8501 (N_8501,N_7666,N_8091);
nor U8502 (N_8502,N_8267,N_7813);
nand U8503 (N_8503,N_7730,N_8093);
nor U8504 (N_8504,N_8194,N_7368);
nand U8505 (N_8505,N_7216,N_8346);
and U8506 (N_8506,N_7490,N_7464);
and U8507 (N_8507,N_8148,N_8359);
and U8508 (N_8508,N_7443,N_8217);
xor U8509 (N_8509,N_7995,N_7720);
nor U8510 (N_8510,N_8398,N_7746);
nor U8511 (N_8511,N_8162,N_8094);
nor U8512 (N_8512,N_8106,N_8018);
nor U8513 (N_8513,N_7970,N_8370);
and U8514 (N_8514,N_8320,N_7814);
and U8515 (N_8515,N_7301,N_7950);
or U8516 (N_8516,N_8189,N_8339);
nand U8517 (N_8517,N_7870,N_7336);
nand U8518 (N_8518,N_7516,N_7637);
nand U8519 (N_8519,N_7826,N_8354);
or U8520 (N_8520,N_7507,N_7912);
xnor U8521 (N_8521,N_7452,N_7580);
nand U8522 (N_8522,N_7414,N_7812);
xnor U8523 (N_8523,N_7212,N_7514);
nand U8524 (N_8524,N_8012,N_7551);
nand U8525 (N_8525,N_7825,N_8270);
xnor U8526 (N_8526,N_8022,N_7833);
and U8527 (N_8527,N_7545,N_7547);
nor U8528 (N_8528,N_7874,N_8351);
or U8529 (N_8529,N_8107,N_7393);
nand U8530 (N_8530,N_7335,N_7594);
or U8531 (N_8531,N_7253,N_7271);
nor U8532 (N_8532,N_7365,N_7647);
xor U8533 (N_8533,N_7543,N_7447);
xnor U8534 (N_8534,N_7437,N_7777);
nand U8535 (N_8535,N_7272,N_7805);
nor U8536 (N_8536,N_8385,N_7566);
nor U8537 (N_8537,N_8172,N_7770);
or U8538 (N_8538,N_8344,N_8380);
nand U8539 (N_8539,N_7355,N_7608);
and U8540 (N_8540,N_7567,N_7494);
xnor U8541 (N_8541,N_8104,N_7501);
and U8542 (N_8542,N_8153,N_7311);
nor U8543 (N_8543,N_7769,N_8247);
and U8544 (N_8544,N_8188,N_7675);
nor U8545 (N_8545,N_7428,N_7867);
xnor U8546 (N_8546,N_8039,N_8082);
nor U8547 (N_8547,N_7343,N_7380);
nand U8548 (N_8548,N_7986,N_8373);
or U8549 (N_8549,N_7223,N_7375);
and U8550 (N_8550,N_7693,N_8177);
or U8551 (N_8551,N_8321,N_7939);
or U8552 (N_8552,N_7765,N_8037);
nor U8553 (N_8553,N_8156,N_7620);
and U8554 (N_8554,N_8274,N_7741);
nand U8555 (N_8555,N_7224,N_7558);
nor U8556 (N_8556,N_8105,N_7577);
xnor U8557 (N_8557,N_7583,N_7204);
nand U8558 (N_8558,N_8322,N_7590);
nand U8559 (N_8559,N_7458,N_7672);
nor U8560 (N_8560,N_8368,N_7960);
or U8561 (N_8561,N_8291,N_7988);
and U8562 (N_8562,N_7724,N_7651);
xnor U8563 (N_8563,N_7599,N_8004);
and U8564 (N_8564,N_8284,N_8096);
and U8565 (N_8565,N_7363,N_8062);
xnor U8566 (N_8566,N_7511,N_8089);
nand U8567 (N_8567,N_7427,N_7241);
or U8568 (N_8568,N_7652,N_8259);
nand U8569 (N_8569,N_7868,N_8276);
xor U8570 (N_8570,N_7866,N_8292);
and U8571 (N_8571,N_7971,N_7671);
or U8572 (N_8572,N_8160,N_8350);
nand U8573 (N_8573,N_7391,N_8088);
nand U8574 (N_8574,N_7441,N_7251);
nand U8575 (N_8575,N_8066,N_8027);
or U8576 (N_8576,N_7678,N_8001);
nor U8577 (N_8577,N_8099,N_8200);
nand U8578 (N_8578,N_7635,N_7654);
nor U8579 (N_8579,N_7860,N_8256);
nor U8580 (N_8580,N_8308,N_8289);
nor U8581 (N_8581,N_8235,N_7292);
nand U8582 (N_8582,N_7515,N_7372);
and U8583 (N_8583,N_7274,N_7256);
nor U8584 (N_8584,N_7564,N_7713);
and U8585 (N_8585,N_8142,N_7766);
xnor U8586 (N_8586,N_7649,N_7690);
or U8587 (N_8587,N_7450,N_7843);
nand U8588 (N_8588,N_7940,N_8295);
xor U8589 (N_8589,N_8038,N_8057);
or U8590 (N_8590,N_8019,N_7337);
and U8591 (N_8591,N_7277,N_8296);
and U8592 (N_8592,N_8379,N_7683);
and U8593 (N_8593,N_7412,N_7346);
or U8594 (N_8594,N_7831,N_8166);
or U8595 (N_8595,N_8145,N_8067);
nor U8596 (N_8596,N_7404,N_7398);
and U8597 (N_8597,N_7895,N_7557);
nand U8598 (N_8598,N_7582,N_7981);
nor U8599 (N_8599,N_7705,N_7857);
and U8600 (N_8600,N_7341,N_8343);
or U8601 (N_8601,N_7663,N_8002);
nor U8602 (N_8602,N_8029,N_7816);
and U8603 (N_8603,N_8024,N_7488);
and U8604 (N_8604,N_8285,N_8074);
nor U8605 (N_8605,N_8241,N_7327);
and U8606 (N_8606,N_7861,N_8240);
and U8607 (N_8607,N_7658,N_7919);
nand U8608 (N_8608,N_8244,N_7800);
xnor U8609 (N_8609,N_7742,N_8117);
nand U8610 (N_8610,N_7801,N_7781);
and U8611 (N_8611,N_7723,N_8386);
or U8612 (N_8612,N_8393,N_7559);
nand U8613 (N_8613,N_8178,N_8190);
nand U8614 (N_8614,N_7369,N_7390);
nand U8615 (N_8615,N_8025,N_7664);
and U8616 (N_8616,N_8165,N_7957);
xnor U8617 (N_8617,N_7616,N_7536);
nand U8618 (N_8618,N_7682,N_8250);
and U8619 (N_8619,N_8213,N_7653);
or U8620 (N_8620,N_7349,N_7706);
or U8621 (N_8621,N_7702,N_7381);
and U8622 (N_8622,N_8169,N_8272);
xor U8623 (N_8623,N_8135,N_7764);
nand U8624 (N_8624,N_7975,N_8238);
nor U8625 (N_8625,N_7246,N_7342);
or U8626 (N_8626,N_8195,N_7601);
nor U8627 (N_8627,N_7703,N_7750);
or U8628 (N_8628,N_7768,N_7700);
nand U8629 (N_8629,N_7968,N_7288);
xnor U8630 (N_8630,N_7340,N_8273);
xor U8631 (N_8631,N_7747,N_7280);
xnor U8632 (N_8632,N_8140,N_7538);
nor U8633 (N_8633,N_8288,N_7681);
and U8634 (N_8634,N_7238,N_7495);
xnor U8635 (N_8635,N_7710,N_7298);
nand U8636 (N_8636,N_7935,N_7707);
nand U8637 (N_8637,N_7344,N_8326);
nand U8638 (N_8638,N_7527,N_8087);
nor U8639 (N_8639,N_7306,N_8282);
xnor U8640 (N_8640,N_7791,N_7210);
and U8641 (N_8641,N_7454,N_8356);
and U8642 (N_8642,N_7378,N_7909);
nor U8643 (N_8643,N_7228,N_7854);
xor U8644 (N_8644,N_7680,N_7392);
nor U8645 (N_8645,N_8134,N_7883);
nand U8646 (N_8646,N_7829,N_8391);
or U8647 (N_8647,N_7921,N_7468);
nor U8648 (N_8648,N_7743,N_7760);
and U8649 (N_8649,N_8268,N_7415);
nand U8650 (N_8650,N_7752,N_7820);
and U8651 (N_8651,N_8290,N_8378);
xnor U8652 (N_8652,N_7721,N_7619);
or U8653 (N_8653,N_7291,N_8203);
nor U8654 (N_8654,N_8364,N_8298);
nand U8655 (N_8655,N_7453,N_7330);
or U8656 (N_8656,N_8277,N_8005);
nand U8657 (N_8657,N_8312,N_8182);
nand U8658 (N_8658,N_8032,N_7876);
xnor U8659 (N_8659,N_8020,N_7920);
and U8660 (N_8660,N_7908,N_7303);
xor U8661 (N_8661,N_7585,N_8130);
nand U8662 (N_8662,N_8127,N_8116);
xnor U8663 (N_8663,N_8204,N_7751);
xnor U8664 (N_8664,N_8233,N_8173);
nor U8665 (N_8665,N_8085,N_8249);
xor U8666 (N_8666,N_7839,N_7523);
nor U8667 (N_8667,N_8299,N_7609);
xor U8668 (N_8668,N_7354,N_8042);
nor U8669 (N_8669,N_7788,N_8234);
or U8670 (N_8670,N_8337,N_8147);
nand U8671 (N_8671,N_7877,N_7626);
and U8672 (N_8672,N_7684,N_7822);
nor U8673 (N_8673,N_7745,N_8103);
nand U8674 (N_8674,N_7896,N_7555);
xor U8675 (N_8675,N_7245,N_8003);
nand U8676 (N_8676,N_7729,N_7990);
nand U8677 (N_8677,N_7954,N_7289);
or U8678 (N_8678,N_7930,N_7836);
or U8679 (N_8679,N_7853,N_7374);
nand U8680 (N_8680,N_8086,N_7978);
and U8681 (N_8681,N_7434,N_7497);
or U8682 (N_8682,N_7249,N_8254);
nand U8683 (N_8683,N_7676,N_8318);
and U8684 (N_8684,N_7949,N_7239);
xnor U8685 (N_8685,N_8095,N_7401);
nand U8686 (N_8686,N_8112,N_7206);
nor U8687 (N_8687,N_8281,N_8341);
xnor U8688 (N_8688,N_7463,N_7841);
nand U8689 (N_8689,N_7804,N_7753);
nor U8690 (N_8690,N_7361,N_7244);
and U8691 (N_8691,N_8216,N_8054);
or U8692 (N_8692,N_8307,N_7904);
nor U8693 (N_8693,N_7961,N_8043);
xor U8694 (N_8694,N_8122,N_7907);
nand U8695 (N_8695,N_8382,N_7331);
and U8696 (N_8696,N_7319,N_7297);
xor U8697 (N_8697,N_8114,N_7903);
or U8698 (N_8698,N_8397,N_8141);
xor U8699 (N_8699,N_7982,N_7610);
nor U8700 (N_8700,N_7269,N_8362);
xor U8701 (N_8701,N_7440,N_7205);
nor U8702 (N_8702,N_7202,N_7891);
nor U8703 (N_8703,N_7708,N_8137);
or U8704 (N_8704,N_8193,N_7479);
nand U8705 (N_8705,N_7569,N_7719);
nand U8706 (N_8706,N_8175,N_7486);
nor U8707 (N_8707,N_7648,N_7592);
or U8708 (N_8708,N_8220,N_7505);
or U8709 (N_8709,N_7321,N_7264);
nand U8710 (N_8710,N_7537,N_7602);
and U8711 (N_8711,N_8333,N_8358);
nor U8712 (N_8712,N_7359,N_8226);
nand U8713 (N_8713,N_8340,N_7548);
nand U8714 (N_8714,N_7293,N_7756);
nand U8715 (N_8715,N_7761,N_7247);
xor U8716 (N_8716,N_8186,N_7317);
nor U8717 (N_8717,N_7827,N_7716);
or U8718 (N_8718,N_8275,N_7504);
and U8719 (N_8719,N_7926,N_7902);
or U8720 (N_8720,N_7364,N_7997);
or U8721 (N_8721,N_7316,N_7835);
nand U8722 (N_8722,N_7980,N_7409);
nor U8723 (N_8723,N_7587,N_7203);
xor U8724 (N_8724,N_8143,N_7588);
and U8725 (N_8725,N_7429,N_7945);
nor U8726 (N_8726,N_8271,N_7283);
nand U8727 (N_8727,N_7521,N_8080);
nor U8728 (N_8728,N_8090,N_7461);
xnor U8729 (N_8729,N_7282,N_8229);
and U8730 (N_8730,N_7644,N_7565);
or U8731 (N_8731,N_7617,N_7882);
xor U8732 (N_8732,N_8353,N_7689);
nand U8733 (N_8733,N_8007,N_7531);
and U8734 (N_8734,N_7948,N_7562);
and U8735 (N_8735,N_7252,N_8097);
nand U8736 (N_8736,N_7222,N_7489);
or U8737 (N_8737,N_8392,N_8023);
xor U8738 (N_8738,N_8301,N_7838);
nor U8739 (N_8739,N_7775,N_7615);
and U8740 (N_8740,N_7969,N_8174);
or U8741 (N_8741,N_7951,N_7384);
nor U8742 (N_8742,N_7798,N_7736);
nor U8743 (N_8743,N_8329,N_7697);
or U8744 (N_8744,N_7300,N_8261);
and U8745 (N_8745,N_7714,N_7229);
xnor U8746 (N_8746,N_7323,N_8031);
and U8747 (N_8747,N_7312,N_8286);
or U8748 (N_8748,N_7242,N_8360);
nor U8749 (N_8749,N_7655,N_7992);
and U8750 (N_8750,N_7650,N_8065);
and U8751 (N_8751,N_7552,N_8035);
xnor U8752 (N_8752,N_7400,N_7262);
xnor U8753 (N_8753,N_7840,N_7735);
nor U8754 (N_8754,N_8196,N_8050);
or U8755 (N_8755,N_7972,N_7535);
and U8756 (N_8756,N_7910,N_7834);
or U8757 (N_8757,N_7318,N_7482);
xor U8758 (N_8758,N_7214,N_8201);
xnor U8759 (N_8759,N_7500,N_7506);
and U8760 (N_8760,N_7438,N_7457);
or U8761 (N_8761,N_7696,N_7231);
nor U8762 (N_8762,N_7821,N_7669);
and U8763 (N_8763,N_7633,N_8108);
nor U8764 (N_8764,N_8365,N_7376);
or U8765 (N_8765,N_7613,N_7307);
nor U8766 (N_8766,N_8176,N_8258);
nand U8767 (N_8767,N_8157,N_8192);
or U8768 (N_8768,N_8376,N_7294);
nor U8769 (N_8769,N_7759,N_7732);
or U8770 (N_8770,N_8262,N_8389);
xnor U8771 (N_8771,N_7574,N_7314);
nor U8772 (N_8772,N_7226,N_8113);
xor U8773 (N_8773,N_7315,N_7263);
nand U8774 (N_8774,N_7900,N_7941);
xnor U8775 (N_8775,N_7528,N_7618);
nand U8776 (N_8776,N_7230,N_7417);
xnor U8777 (N_8777,N_7845,N_7925);
xnor U8778 (N_8778,N_7589,N_8366);
or U8779 (N_8779,N_7394,N_7406);
nand U8780 (N_8780,N_7502,N_8070);
and U8781 (N_8781,N_8325,N_8363);
xor U8782 (N_8782,N_7973,N_7383);
and U8783 (N_8783,N_7413,N_7276);
xor U8784 (N_8784,N_7808,N_7783);
xnor U8785 (N_8785,N_7740,N_7347);
nor U8786 (N_8786,N_7849,N_8118);
xnor U8787 (N_8787,N_8111,N_7852);
nand U8788 (N_8788,N_7819,N_7370);
xnor U8789 (N_8789,N_8121,N_8335);
nor U8790 (N_8790,N_8119,N_7737);
nor U8791 (N_8791,N_7600,N_8180);
and U8792 (N_8792,N_7334,N_7568);
nor U8793 (N_8793,N_7546,N_7979);
xnor U8794 (N_8794,N_7603,N_7963);
and U8795 (N_8795,N_7433,N_8208);
or U8796 (N_8796,N_7622,N_7422);
nand U8797 (N_8797,N_8120,N_7402);
and U8798 (N_8798,N_7899,N_7385);
nand U8799 (N_8799,N_7928,N_8149);
nor U8800 (N_8800,N_7572,N_7456);
xor U8801 (N_8801,N_7533,N_7540);
and U8802 (N_8802,N_8068,N_7436);
nor U8803 (N_8803,N_7329,N_8052);
and U8804 (N_8804,N_7859,N_7792);
and U8805 (N_8805,N_8253,N_8036);
xnor U8806 (N_8806,N_7208,N_7911);
xnor U8807 (N_8807,N_7656,N_8053);
nor U8808 (N_8808,N_7830,N_7513);
xnor U8809 (N_8809,N_8101,N_8323);
nor U8810 (N_8810,N_7561,N_7287);
nor U8811 (N_8811,N_7728,N_8079);
nor U8812 (N_8812,N_7209,N_7779);
xnor U8813 (N_8813,N_7889,N_8187);
nand U8814 (N_8814,N_7802,N_7787);
nand U8815 (N_8815,N_8394,N_7550);
xnor U8816 (N_8816,N_8390,N_7906);
xor U8817 (N_8817,N_7758,N_8287);
nor U8818 (N_8818,N_8328,N_7688);
nand U8819 (N_8819,N_7694,N_7776);
xor U8820 (N_8820,N_7987,N_8044);
and U8821 (N_8821,N_7964,N_7221);
and U8822 (N_8822,N_7322,N_8072);
or U8823 (N_8823,N_7270,N_7299);
nor U8824 (N_8824,N_8000,N_8367);
nand U8825 (N_8825,N_7880,N_8109);
nand U8826 (N_8826,N_7711,N_7225);
nand U8827 (N_8827,N_8305,N_7888);
and U8828 (N_8828,N_7699,N_7425);
nand U8829 (N_8829,N_7305,N_7235);
and U8830 (N_8830,N_7524,N_8159);
or U8831 (N_8831,N_7460,N_7674);
xnor U8832 (N_8832,N_8228,N_8314);
xor U8833 (N_8833,N_8348,N_7892);
xor U8834 (N_8834,N_8311,N_8223);
and U8835 (N_8835,N_7864,N_8375);
or U8836 (N_8836,N_7366,N_8125);
or U8837 (N_8837,N_7478,N_7290);
nor U8838 (N_8838,N_7661,N_7846);
nand U8839 (N_8839,N_7503,N_7793);
or U8840 (N_8840,N_7692,N_8327);
nand U8841 (N_8841,N_8209,N_7771);
and U8842 (N_8842,N_8017,N_7958);
nor U8843 (N_8843,N_7444,N_7886);
nor U8844 (N_8844,N_8332,N_8056);
or U8845 (N_8845,N_7508,N_8374);
and U8846 (N_8846,N_8028,N_7924);
or U8847 (N_8847,N_7749,N_7480);
xnor U8848 (N_8848,N_7399,N_8264);
or U8849 (N_8849,N_7623,N_7459);
or U8850 (N_8850,N_7424,N_7560);
or U8851 (N_8851,N_7426,N_7687);
nand U8852 (N_8852,N_7931,N_7496);
xor U8853 (N_8853,N_7862,N_8154);
nor U8854 (N_8854,N_8313,N_7581);
and U8855 (N_8855,N_8138,N_7358);
xor U8856 (N_8856,N_7786,N_7591);
nand U8857 (N_8857,N_7605,N_8239);
xor U8858 (N_8858,N_7573,N_7885);
xnor U8859 (N_8859,N_8300,N_8222);
xnor U8860 (N_8860,N_7738,N_8063);
and U8861 (N_8861,N_7260,N_8263);
xor U8862 (N_8862,N_7850,N_8221);
xnor U8863 (N_8863,N_7933,N_7946);
xnor U8864 (N_8864,N_7996,N_7356);
and U8865 (N_8865,N_7983,N_7869);
nand U8866 (N_8866,N_8211,N_7722);
xnor U8867 (N_8867,N_8184,N_7462);
xor U8868 (N_8868,N_8331,N_8330);
nand U8869 (N_8869,N_7645,N_7407);
and U8870 (N_8870,N_7420,N_7667);
or U8871 (N_8871,N_8242,N_7423);
xnor U8872 (N_8872,N_7673,N_7339);
or U8873 (N_8873,N_7953,N_7809);
or U8874 (N_8874,N_7387,N_7200);
xnor U8875 (N_8875,N_8075,N_7873);
or U8876 (N_8876,N_7937,N_8283);
and U8877 (N_8877,N_8049,N_7898);
nand U8878 (N_8878,N_8006,N_8205);
or U8879 (N_8879,N_7539,N_7304);
or U8880 (N_8880,N_7326,N_8010);
xnor U8881 (N_8881,N_7309,N_8251);
xnor U8882 (N_8882,N_8336,N_7386);
xnor U8883 (N_8883,N_7727,N_8232);
nor U8884 (N_8884,N_8152,N_7281);
nor U8885 (N_8885,N_7236,N_7237);
nand U8886 (N_8886,N_7302,N_7410);
or U8887 (N_8887,N_8210,N_8212);
xor U8888 (N_8888,N_7522,N_7966);
or U8889 (N_8889,N_7279,N_7485);
or U8890 (N_8890,N_8102,N_7630);
and U8891 (N_8891,N_7744,N_8396);
xnor U8892 (N_8892,N_8319,N_7763);
nand U8893 (N_8893,N_7897,N_7828);
nand U8894 (N_8894,N_7596,N_7976);
xor U8895 (N_8895,N_7477,N_7627);
xor U8896 (N_8896,N_8144,N_7492);
xor U8897 (N_8897,N_8303,N_7780);
xnor U8898 (N_8898,N_7847,N_7211);
nor U8899 (N_8899,N_7842,N_8155);
or U8900 (N_8900,N_7371,N_7435);
nand U8901 (N_8901,N_8246,N_8369);
nor U8902 (N_8902,N_7278,N_7345);
nor U8903 (N_8903,N_7571,N_7240);
and U8904 (N_8904,N_7563,N_8083);
and U8905 (N_8905,N_7403,N_7579);
nor U8906 (N_8906,N_7310,N_8078);
nor U8907 (N_8907,N_8013,N_8227);
nand U8908 (N_8908,N_7943,N_8387);
and U8909 (N_8909,N_8132,N_8304);
xnor U8910 (N_8910,N_7817,N_7258);
and U8911 (N_8911,N_7285,N_7977);
nand U8912 (N_8912,N_7942,N_7784);
xnor U8913 (N_8913,N_8033,N_7491);
and U8914 (N_8914,N_8161,N_8179);
nand U8915 (N_8915,N_7612,N_7757);
or U8916 (N_8916,N_8123,N_8352);
nand U8917 (N_8917,N_7377,N_7668);
nor U8918 (N_8918,N_7584,N_8191);
nor U8919 (N_8919,N_7348,N_7418);
nand U8920 (N_8920,N_7795,N_8168);
and U8921 (N_8921,N_8041,N_8384);
and U8922 (N_8922,N_8255,N_7918);
nor U8923 (N_8923,N_7475,N_7207);
or U8924 (N_8924,N_8334,N_7352);
or U8925 (N_8925,N_8047,N_7932);
nor U8926 (N_8926,N_7965,N_7333);
xnor U8927 (N_8927,N_7894,N_7614);
and U8928 (N_8928,N_7731,N_7611);
xor U8929 (N_8929,N_7811,N_8197);
and U8930 (N_8930,N_7517,N_7884);
or U8931 (N_8931,N_8349,N_7267);
or U8932 (N_8932,N_8016,N_7865);
nor U8933 (N_8933,N_7389,N_8237);
or U8934 (N_8934,N_7754,N_8021);
and U8935 (N_8935,N_8110,N_8129);
nand U8936 (N_8936,N_7639,N_7213);
and U8937 (N_8937,N_7218,N_7219);
nand U8938 (N_8938,N_8231,N_7701);
xor U8939 (N_8939,N_7646,N_8265);
and U8940 (N_8940,N_7296,N_8098);
nand U8941 (N_8941,N_8034,N_7570);
and U8942 (N_8942,N_8248,N_8230);
xnor U8943 (N_8943,N_8071,N_7382);
nor U8944 (N_8944,N_7796,N_8059);
nand U8945 (N_8945,N_8146,N_8115);
and U8946 (N_8946,N_7607,N_8150);
and U8947 (N_8947,N_7578,N_7324);
xor U8948 (N_8948,N_7837,N_7498);
or U8949 (N_8949,N_7328,N_8315);
nand U8950 (N_8950,N_8207,N_8302);
xnor U8951 (N_8951,N_7739,N_8324);
or U8952 (N_8952,N_7367,N_7430);
xnor U8953 (N_8953,N_7989,N_7509);
and U8954 (N_8954,N_8377,N_7773);
and U8955 (N_8955,N_8163,N_7320);
or U8956 (N_8956,N_7789,N_7534);
nand U8957 (N_8957,N_7268,N_7593);
nand U8958 (N_8958,N_7416,N_7474);
nand U8959 (N_8959,N_8294,N_7938);
and U8960 (N_8960,N_8342,N_7858);
nor U8961 (N_8961,N_7890,N_7396);
nand U8962 (N_8962,N_7659,N_7295);
xor U8963 (N_8963,N_7878,N_8309);
or U8964 (N_8964,N_7803,N_7261);
nand U8965 (N_8965,N_7662,N_7778);
nand U8966 (N_8966,N_7248,N_8388);
xnor U8967 (N_8967,N_7994,N_8100);
or U8968 (N_8968,N_7879,N_7974);
nand U8969 (N_8969,N_7449,N_7660);
or U8970 (N_8970,N_7451,N_7685);
xnor U8971 (N_8971,N_7421,N_7466);
or U8972 (N_8972,N_7998,N_8055);
and U8973 (N_8973,N_7604,N_7446);
xnor U8974 (N_8974,N_8202,N_7952);
and U8975 (N_8975,N_7529,N_7962);
nand U8976 (N_8976,N_8243,N_7785);
nor U8977 (N_8977,N_8355,N_7232);
and U8978 (N_8978,N_8381,N_7265);
or U8979 (N_8979,N_7243,N_7993);
or U8980 (N_8980,N_7984,N_7677);
xnor U8981 (N_8981,N_7936,N_8316);
nor U8982 (N_8982,N_7338,N_8170);
nor U8983 (N_8983,N_8008,N_7628);
or U8984 (N_8984,N_7695,N_7467);
or U8985 (N_8985,N_7726,N_8045);
nor U8986 (N_8986,N_8215,N_8011);
and U8987 (N_8987,N_7313,N_7704);
and U8988 (N_8988,N_7967,N_7621);
and U8989 (N_8989,N_8236,N_7810);
xor U8990 (N_8990,N_7388,N_7598);
nor U8991 (N_8991,N_7487,N_7799);
or U8992 (N_8992,N_7597,N_8225);
nand U8993 (N_8993,N_7670,N_7818);
nand U8994 (N_8994,N_7469,N_7259);
nor U8995 (N_8995,N_8199,N_7807);
nor U8996 (N_8996,N_8214,N_7379);
nor U8997 (N_8997,N_7863,N_7856);
or U8998 (N_8998,N_8048,N_8092);
or U8999 (N_8999,N_7725,N_8293);
and U9000 (N_9000,N_7572,N_7886);
nor U9001 (N_9001,N_7453,N_7864);
or U9002 (N_9002,N_8156,N_8367);
xor U9003 (N_9003,N_8123,N_8253);
nand U9004 (N_9004,N_8135,N_8255);
nand U9005 (N_9005,N_7374,N_7485);
or U9006 (N_9006,N_8170,N_7548);
xnor U9007 (N_9007,N_8112,N_7810);
nor U9008 (N_9008,N_7461,N_7955);
and U9009 (N_9009,N_8190,N_7213);
xor U9010 (N_9010,N_7377,N_7465);
xnor U9011 (N_9011,N_7237,N_7721);
or U9012 (N_9012,N_8057,N_7882);
nor U9013 (N_9013,N_8161,N_7432);
xnor U9014 (N_9014,N_7832,N_7482);
nand U9015 (N_9015,N_8100,N_8266);
nor U9016 (N_9016,N_7540,N_7283);
and U9017 (N_9017,N_8164,N_7781);
and U9018 (N_9018,N_8151,N_8019);
nand U9019 (N_9019,N_7651,N_7474);
nand U9020 (N_9020,N_8015,N_8166);
or U9021 (N_9021,N_7430,N_7592);
nor U9022 (N_9022,N_8286,N_8304);
xor U9023 (N_9023,N_7796,N_7849);
or U9024 (N_9024,N_8191,N_8207);
or U9025 (N_9025,N_8180,N_8345);
nand U9026 (N_9026,N_7566,N_7866);
or U9027 (N_9027,N_7239,N_7783);
or U9028 (N_9028,N_8307,N_7934);
or U9029 (N_9029,N_7733,N_7912);
xor U9030 (N_9030,N_7571,N_7944);
or U9031 (N_9031,N_7281,N_8102);
xor U9032 (N_9032,N_7614,N_8262);
nand U9033 (N_9033,N_7497,N_8120);
nand U9034 (N_9034,N_8033,N_7244);
or U9035 (N_9035,N_7519,N_7837);
and U9036 (N_9036,N_8214,N_8381);
nand U9037 (N_9037,N_8015,N_7932);
nand U9038 (N_9038,N_7386,N_7441);
xor U9039 (N_9039,N_8345,N_7782);
or U9040 (N_9040,N_8038,N_7999);
or U9041 (N_9041,N_7419,N_7200);
xor U9042 (N_9042,N_8359,N_7962);
or U9043 (N_9043,N_7752,N_8005);
xor U9044 (N_9044,N_7589,N_7974);
or U9045 (N_9045,N_7350,N_7580);
or U9046 (N_9046,N_7471,N_7507);
nand U9047 (N_9047,N_7920,N_7397);
or U9048 (N_9048,N_7361,N_8164);
xnor U9049 (N_9049,N_7912,N_7548);
nor U9050 (N_9050,N_8370,N_7408);
nor U9051 (N_9051,N_7877,N_8151);
or U9052 (N_9052,N_7801,N_7530);
or U9053 (N_9053,N_7495,N_7540);
or U9054 (N_9054,N_7496,N_7651);
nor U9055 (N_9055,N_7216,N_7349);
nand U9056 (N_9056,N_7294,N_7234);
xnor U9057 (N_9057,N_7435,N_7971);
or U9058 (N_9058,N_7971,N_8377);
or U9059 (N_9059,N_7867,N_8094);
and U9060 (N_9060,N_8277,N_8137);
xnor U9061 (N_9061,N_7206,N_7449);
nand U9062 (N_9062,N_7496,N_7639);
nor U9063 (N_9063,N_8262,N_7301);
nand U9064 (N_9064,N_8270,N_7295);
nand U9065 (N_9065,N_7249,N_7386);
or U9066 (N_9066,N_7485,N_7427);
and U9067 (N_9067,N_8380,N_7298);
or U9068 (N_9068,N_8389,N_7472);
and U9069 (N_9069,N_7680,N_8396);
nand U9070 (N_9070,N_8172,N_8027);
nor U9071 (N_9071,N_7377,N_7616);
or U9072 (N_9072,N_7620,N_8327);
or U9073 (N_9073,N_7711,N_7440);
nand U9074 (N_9074,N_8087,N_8105);
or U9075 (N_9075,N_8078,N_7926);
nand U9076 (N_9076,N_8335,N_8354);
or U9077 (N_9077,N_7535,N_7321);
and U9078 (N_9078,N_7501,N_7719);
or U9079 (N_9079,N_7914,N_8363);
nor U9080 (N_9080,N_8116,N_7307);
and U9081 (N_9081,N_7203,N_8197);
xor U9082 (N_9082,N_7417,N_7279);
xor U9083 (N_9083,N_7561,N_7744);
and U9084 (N_9084,N_7779,N_7383);
xnor U9085 (N_9085,N_7359,N_8304);
xnor U9086 (N_9086,N_7941,N_8056);
and U9087 (N_9087,N_7297,N_8364);
xnor U9088 (N_9088,N_7916,N_8179);
xor U9089 (N_9089,N_7471,N_8141);
and U9090 (N_9090,N_7775,N_8329);
nor U9091 (N_9091,N_8203,N_7493);
xor U9092 (N_9092,N_8129,N_7796);
xnor U9093 (N_9093,N_7497,N_8181);
xor U9094 (N_9094,N_7470,N_7647);
nand U9095 (N_9095,N_7382,N_7779);
and U9096 (N_9096,N_7987,N_8065);
nor U9097 (N_9097,N_7595,N_7498);
and U9098 (N_9098,N_8326,N_7258);
nor U9099 (N_9099,N_7691,N_7667);
nand U9100 (N_9100,N_7876,N_8239);
nor U9101 (N_9101,N_7863,N_7544);
nand U9102 (N_9102,N_7708,N_8048);
xnor U9103 (N_9103,N_7739,N_7776);
and U9104 (N_9104,N_8015,N_8054);
nand U9105 (N_9105,N_8314,N_7700);
and U9106 (N_9106,N_8327,N_8186);
xor U9107 (N_9107,N_8026,N_7691);
xor U9108 (N_9108,N_8204,N_8083);
xnor U9109 (N_9109,N_7652,N_7953);
nand U9110 (N_9110,N_8127,N_8066);
nor U9111 (N_9111,N_7425,N_7697);
nor U9112 (N_9112,N_7738,N_7565);
or U9113 (N_9113,N_7953,N_8171);
xnor U9114 (N_9114,N_7565,N_8259);
and U9115 (N_9115,N_7394,N_8358);
and U9116 (N_9116,N_7833,N_7308);
xor U9117 (N_9117,N_8297,N_7932);
nand U9118 (N_9118,N_7263,N_8275);
nor U9119 (N_9119,N_8299,N_7463);
nor U9120 (N_9120,N_7707,N_7496);
xor U9121 (N_9121,N_7392,N_7634);
nor U9122 (N_9122,N_8143,N_7660);
nand U9123 (N_9123,N_7739,N_8059);
and U9124 (N_9124,N_7666,N_7848);
or U9125 (N_9125,N_8368,N_7719);
and U9126 (N_9126,N_8138,N_7516);
or U9127 (N_9127,N_7870,N_7891);
nor U9128 (N_9128,N_8210,N_7870);
nand U9129 (N_9129,N_7482,N_8354);
or U9130 (N_9130,N_7660,N_7895);
xnor U9131 (N_9131,N_7924,N_8140);
xnor U9132 (N_9132,N_7217,N_8100);
xnor U9133 (N_9133,N_8203,N_7761);
xnor U9134 (N_9134,N_7398,N_7830);
nor U9135 (N_9135,N_7477,N_8313);
nor U9136 (N_9136,N_8290,N_7449);
nand U9137 (N_9137,N_7546,N_8273);
nand U9138 (N_9138,N_7226,N_7700);
or U9139 (N_9139,N_7802,N_7682);
xnor U9140 (N_9140,N_7420,N_7540);
or U9141 (N_9141,N_7489,N_8319);
nor U9142 (N_9142,N_8239,N_7885);
or U9143 (N_9143,N_8148,N_7347);
and U9144 (N_9144,N_8356,N_8349);
and U9145 (N_9145,N_8354,N_7738);
nand U9146 (N_9146,N_7727,N_7389);
xor U9147 (N_9147,N_8284,N_7839);
xnor U9148 (N_9148,N_7352,N_7549);
nand U9149 (N_9149,N_7676,N_8188);
or U9150 (N_9150,N_8244,N_7738);
and U9151 (N_9151,N_8172,N_7687);
and U9152 (N_9152,N_7254,N_8062);
nor U9153 (N_9153,N_7247,N_7378);
nand U9154 (N_9154,N_8130,N_7983);
xor U9155 (N_9155,N_7220,N_7680);
or U9156 (N_9156,N_7542,N_7675);
nor U9157 (N_9157,N_7850,N_7557);
xor U9158 (N_9158,N_8009,N_7222);
or U9159 (N_9159,N_7763,N_7605);
and U9160 (N_9160,N_7840,N_8164);
and U9161 (N_9161,N_8101,N_8208);
nor U9162 (N_9162,N_8076,N_7465);
nor U9163 (N_9163,N_7268,N_7380);
nand U9164 (N_9164,N_8344,N_7342);
or U9165 (N_9165,N_8042,N_7824);
nor U9166 (N_9166,N_7219,N_7848);
nand U9167 (N_9167,N_7243,N_7683);
nor U9168 (N_9168,N_8050,N_8143);
and U9169 (N_9169,N_7434,N_7421);
nand U9170 (N_9170,N_8149,N_7557);
xor U9171 (N_9171,N_8036,N_8083);
and U9172 (N_9172,N_7306,N_7607);
nand U9173 (N_9173,N_8099,N_7941);
nand U9174 (N_9174,N_7303,N_8338);
or U9175 (N_9175,N_7979,N_7647);
xor U9176 (N_9176,N_8062,N_7230);
or U9177 (N_9177,N_7735,N_7650);
and U9178 (N_9178,N_8086,N_8142);
nor U9179 (N_9179,N_8057,N_7855);
and U9180 (N_9180,N_7620,N_8113);
nand U9181 (N_9181,N_7310,N_7882);
and U9182 (N_9182,N_8382,N_8002);
or U9183 (N_9183,N_8281,N_8068);
nor U9184 (N_9184,N_7405,N_8067);
or U9185 (N_9185,N_7517,N_7857);
or U9186 (N_9186,N_8159,N_8080);
or U9187 (N_9187,N_8380,N_7964);
nor U9188 (N_9188,N_8172,N_7453);
xor U9189 (N_9189,N_8259,N_7766);
and U9190 (N_9190,N_8059,N_7512);
nand U9191 (N_9191,N_7715,N_7500);
nand U9192 (N_9192,N_7534,N_8352);
or U9193 (N_9193,N_7470,N_7496);
nand U9194 (N_9194,N_7326,N_7982);
or U9195 (N_9195,N_8182,N_7880);
or U9196 (N_9196,N_8112,N_7705);
or U9197 (N_9197,N_7882,N_7281);
nand U9198 (N_9198,N_7758,N_7738);
or U9199 (N_9199,N_7609,N_7912);
xnor U9200 (N_9200,N_8389,N_7408);
xor U9201 (N_9201,N_7968,N_7352);
and U9202 (N_9202,N_8139,N_7503);
nor U9203 (N_9203,N_7431,N_7458);
and U9204 (N_9204,N_8175,N_8161);
xor U9205 (N_9205,N_7675,N_7336);
and U9206 (N_9206,N_7780,N_8353);
nand U9207 (N_9207,N_7790,N_7597);
xnor U9208 (N_9208,N_7740,N_8087);
and U9209 (N_9209,N_7239,N_7465);
nand U9210 (N_9210,N_7790,N_8376);
nand U9211 (N_9211,N_7441,N_8394);
or U9212 (N_9212,N_8003,N_7395);
nor U9213 (N_9213,N_7603,N_8259);
nand U9214 (N_9214,N_7913,N_7605);
and U9215 (N_9215,N_7780,N_8045);
nor U9216 (N_9216,N_7937,N_7750);
xnor U9217 (N_9217,N_7972,N_8146);
xor U9218 (N_9218,N_7811,N_7639);
xor U9219 (N_9219,N_7493,N_7450);
nand U9220 (N_9220,N_7368,N_8082);
nor U9221 (N_9221,N_8320,N_7810);
or U9222 (N_9222,N_7662,N_8135);
nand U9223 (N_9223,N_8368,N_8252);
nor U9224 (N_9224,N_7458,N_8259);
nand U9225 (N_9225,N_7865,N_7860);
xnor U9226 (N_9226,N_7710,N_7969);
nor U9227 (N_9227,N_7520,N_8198);
nand U9228 (N_9228,N_7574,N_8217);
nand U9229 (N_9229,N_7961,N_8185);
xor U9230 (N_9230,N_7572,N_7344);
or U9231 (N_9231,N_7583,N_8223);
or U9232 (N_9232,N_8153,N_7453);
xnor U9233 (N_9233,N_7986,N_7468);
nand U9234 (N_9234,N_8199,N_8103);
and U9235 (N_9235,N_7952,N_7994);
nor U9236 (N_9236,N_7389,N_7422);
xor U9237 (N_9237,N_8068,N_7694);
nor U9238 (N_9238,N_8397,N_7269);
and U9239 (N_9239,N_7643,N_7476);
nor U9240 (N_9240,N_7783,N_7456);
xnor U9241 (N_9241,N_7597,N_7628);
or U9242 (N_9242,N_7755,N_8321);
xnor U9243 (N_9243,N_8223,N_7364);
or U9244 (N_9244,N_7628,N_8215);
xor U9245 (N_9245,N_7255,N_7361);
or U9246 (N_9246,N_7553,N_8359);
and U9247 (N_9247,N_7224,N_8324);
nor U9248 (N_9248,N_8355,N_7974);
nor U9249 (N_9249,N_7390,N_8022);
nor U9250 (N_9250,N_8353,N_7596);
and U9251 (N_9251,N_8270,N_8165);
or U9252 (N_9252,N_7504,N_7702);
or U9253 (N_9253,N_7664,N_7735);
nand U9254 (N_9254,N_8134,N_7251);
xnor U9255 (N_9255,N_7844,N_7564);
nor U9256 (N_9256,N_8090,N_7601);
nand U9257 (N_9257,N_7360,N_7859);
xnor U9258 (N_9258,N_7805,N_7551);
nand U9259 (N_9259,N_7879,N_7507);
nand U9260 (N_9260,N_7228,N_7947);
nor U9261 (N_9261,N_7282,N_7723);
nor U9262 (N_9262,N_8391,N_7438);
xnor U9263 (N_9263,N_7973,N_7472);
xor U9264 (N_9264,N_8000,N_8397);
or U9265 (N_9265,N_7787,N_7908);
and U9266 (N_9266,N_7658,N_8246);
and U9267 (N_9267,N_7583,N_7844);
nand U9268 (N_9268,N_8107,N_8332);
or U9269 (N_9269,N_7261,N_8122);
nand U9270 (N_9270,N_7759,N_7557);
xor U9271 (N_9271,N_8026,N_8109);
or U9272 (N_9272,N_8265,N_7292);
xor U9273 (N_9273,N_7715,N_7571);
or U9274 (N_9274,N_7289,N_7997);
and U9275 (N_9275,N_8384,N_7576);
xor U9276 (N_9276,N_7330,N_7431);
or U9277 (N_9277,N_7947,N_7861);
nand U9278 (N_9278,N_8078,N_7405);
or U9279 (N_9279,N_8213,N_7926);
or U9280 (N_9280,N_7867,N_7866);
and U9281 (N_9281,N_8004,N_8040);
and U9282 (N_9282,N_7485,N_8247);
and U9283 (N_9283,N_7471,N_7222);
nor U9284 (N_9284,N_7436,N_7896);
nor U9285 (N_9285,N_7871,N_8129);
or U9286 (N_9286,N_8378,N_7290);
nor U9287 (N_9287,N_8160,N_7935);
nor U9288 (N_9288,N_7513,N_7297);
nor U9289 (N_9289,N_7347,N_7819);
or U9290 (N_9290,N_8016,N_7266);
or U9291 (N_9291,N_7441,N_7617);
nand U9292 (N_9292,N_8125,N_7794);
and U9293 (N_9293,N_8262,N_7349);
nand U9294 (N_9294,N_7549,N_8174);
or U9295 (N_9295,N_7617,N_8271);
xnor U9296 (N_9296,N_7474,N_8028);
nor U9297 (N_9297,N_7340,N_7987);
nor U9298 (N_9298,N_7911,N_7213);
or U9299 (N_9299,N_7203,N_8258);
and U9300 (N_9300,N_7321,N_7756);
or U9301 (N_9301,N_8368,N_7650);
or U9302 (N_9302,N_7457,N_7990);
nor U9303 (N_9303,N_8086,N_7938);
or U9304 (N_9304,N_8000,N_7816);
and U9305 (N_9305,N_7865,N_7206);
or U9306 (N_9306,N_7317,N_8133);
nor U9307 (N_9307,N_8361,N_7547);
and U9308 (N_9308,N_7866,N_7531);
nand U9309 (N_9309,N_7403,N_7870);
xnor U9310 (N_9310,N_8135,N_7655);
nand U9311 (N_9311,N_8060,N_7454);
nor U9312 (N_9312,N_8372,N_7621);
xor U9313 (N_9313,N_7355,N_7526);
nand U9314 (N_9314,N_7635,N_8208);
xnor U9315 (N_9315,N_7507,N_7561);
xor U9316 (N_9316,N_8235,N_7209);
nand U9317 (N_9317,N_8041,N_7683);
xnor U9318 (N_9318,N_7487,N_7759);
nand U9319 (N_9319,N_7921,N_8167);
nand U9320 (N_9320,N_7742,N_7464);
or U9321 (N_9321,N_7361,N_7518);
and U9322 (N_9322,N_8102,N_7883);
xnor U9323 (N_9323,N_8163,N_8288);
xnor U9324 (N_9324,N_7650,N_8121);
xnor U9325 (N_9325,N_8133,N_8317);
or U9326 (N_9326,N_7524,N_8098);
and U9327 (N_9327,N_7707,N_7915);
nor U9328 (N_9328,N_7640,N_7495);
or U9329 (N_9329,N_8274,N_7307);
nor U9330 (N_9330,N_7489,N_7389);
and U9331 (N_9331,N_7891,N_8024);
nand U9332 (N_9332,N_7417,N_8106);
or U9333 (N_9333,N_7343,N_7316);
nor U9334 (N_9334,N_7585,N_7453);
xnor U9335 (N_9335,N_7809,N_7993);
xor U9336 (N_9336,N_7786,N_8128);
and U9337 (N_9337,N_7495,N_7872);
nor U9338 (N_9338,N_8266,N_8359);
nand U9339 (N_9339,N_7604,N_8362);
nor U9340 (N_9340,N_7972,N_7788);
and U9341 (N_9341,N_7559,N_8239);
nor U9342 (N_9342,N_7819,N_8272);
or U9343 (N_9343,N_7208,N_8152);
nand U9344 (N_9344,N_7584,N_7801);
xnor U9345 (N_9345,N_7352,N_7865);
and U9346 (N_9346,N_8200,N_7715);
or U9347 (N_9347,N_7346,N_7637);
and U9348 (N_9348,N_7693,N_8003);
nor U9349 (N_9349,N_7487,N_7243);
nand U9350 (N_9350,N_8373,N_7586);
nand U9351 (N_9351,N_7360,N_7568);
nor U9352 (N_9352,N_8063,N_7874);
xor U9353 (N_9353,N_7454,N_7709);
or U9354 (N_9354,N_7996,N_7682);
xnor U9355 (N_9355,N_7885,N_7315);
nand U9356 (N_9356,N_7829,N_7224);
and U9357 (N_9357,N_7978,N_8191);
nand U9358 (N_9358,N_7796,N_7327);
and U9359 (N_9359,N_8000,N_7806);
and U9360 (N_9360,N_7447,N_7928);
nor U9361 (N_9361,N_8027,N_7559);
nor U9362 (N_9362,N_7920,N_7808);
nor U9363 (N_9363,N_7732,N_7932);
nand U9364 (N_9364,N_7687,N_7658);
and U9365 (N_9365,N_7374,N_8081);
xnor U9366 (N_9366,N_7846,N_7414);
nor U9367 (N_9367,N_7949,N_8234);
nor U9368 (N_9368,N_8395,N_7442);
xor U9369 (N_9369,N_7252,N_7330);
and U9370 (N_9370,N_8293,N_7814);
nand U9371 (N_9371,N_7355,N_7538);
or U9372 (N_9372,N_7512,N_7763);
nor U9373 (N_9373,N_7925,N_8170);
nand U9374 (N_9374,N_7980,N_7893);
nor U9375 (N_9375,N_7601,N_7340);
nor U9376 (N_9376,N_7607,N_7560);
and U9377 (N_9377,N_7510,N_7309);
and U9378 (N_9378,N_7825,N_8054);
nor U9379 (N_9379,N_7575,N_7470);
xnor U9380 (N_9380,N_8327,N_8336);
or U9381 (N_9381,N_7832,N_7210);
or U9382 (N_9382,N_7525,N_7651);
and U9383 (N_9383,N_7628,N_7431);
or U9384 (N_9384,N_7851,N_7368);
nand U9385 (N_9385,N_8029,N_8296);
nand U9386 (N_9386,N_8383,N_8082);
nor U9387 (N_9387,N_7295,N_7968);
or U9388 (N_9388,N_7707,N_7548);
or U9389 (N_9389,N_7847,N_8397);
nand U9390 (N_9390,N_7823,N_8258);
nand U9391 (N_9391,N_8316,N_7647);
and U9392 (N_9392,N_7834,N_7459);
and U9393 (N_9393,N_8129,N_7984);
or U9394 (N_9394,N_8170,N_7896);
nand U9395 (N_9395,N_7791,N_7835);
nor U9396 (N_9396,N_8350,N_7604);
nand U9397 (N_9397,N_7751,N_7638);
nor U9398 (N_9398,N_7778,N_8321);
nand U9399 (N_9399,N_7240,N_8215);
and U9400 (N_9400,N_7256,N_8242);
nand U9401 (N_9401,N_7367,N_8044);
or U9402 (N_9402,N_7934,N_7523);
or U9403 (N_9403,N_7211,N_7574);
xor U9404 (N_9404,N_7500,N_7611);
xnor U9405 (N_9405,N_7975,N_8335);
xnor U9406 (N_9406,N_7538,N_7919);
or U9407 (N_9407,N_8265,N_7269);
or U9408 (N_9408,N_7241,N_7669);
xnor U9409 (N_9409,N_7780,N_7663);
xnor U9410 (N_9410,N_7913,N_8054);
xor U9411 (N_9411,N_7479,N_7566);
and U9412 (N_9412,N_7379,N_7282);
nand U9413 (N_9413,N_7541,N_7488);
nand U9414 (N_9414,N_7291,N_8294);
nor U9415 (N_9415,N_7735,N_8124);
xor U9416 (N_9416,N_7551,N_7200);
xnor U9417 (N_9417,N_8363,N_7616);
or U9418 (N_9418,N_7675,N_7268);
xor U9419 (N_9419,N_7618,N_7351);
xor U9420 (N_9420,N_8365,N_8050);
xnor U9421 (N_9421,N_7477,N_7505);
xnor U9422 (N_9422,N_8071,N_8184);
and U9423 (N_9423,N_7650,N_8034);
nor U9424 (N_9424,N_7982,N_8070);
xnor U9425 (N_9425,N_7534,N_8250);
and U9426 (N_9426,N_7609,N_8369);
and U9427 (N_9427,N_8091,N_8057);
nand U9428 (N_9428,N_7401,N_8002);
nor U9429 (N_9429,N_7213,N_7215);
and U9430 (N_9430,N_7816,N_7653);
xor U9431 (N_9431,N_8324,N_8255);
or U9432 (N_9432,N_8194,N_7273);
xor U9433 (N_9433,N_7274,N_7655);
nor U9434 (N_9434,N_7738,N_7280);
and U9435 (N_9435,N_7308,N_8041);
and U9436 (N_9436,N_7967,N_8259);
and U9437 (N_9437,N_8082,N_7399);
or U9438 (N_9438,N_7264,N_7720);
nand U9439 (N_9439,N_7294,N_7693);
xor U9440 (N_9440,N_7311,N_8215);
nor U9441 (N_9441,N_7887,N_7856);
or U9442 (N_9442,N_7960,N_7491);
xor U9443 (N_9443,N_7300,N_7410);
nor U9444 (N_9444,N_8174,N_7322);
and U9445 (N_9445,N_7733,N_8303);
and U9446 (N_9446,N_7623,N_7676);
xnor U9447 (N_9447,N_8119,N_7268);
nor U9448 (N_9448,N_7731,N_8271);
xnor U9449 (N_9449,N_7486,N_7938);
xor U9450 (N_9450,N_7989,N_7473);
and U9451 (N_9451,N_7811,N_7499);
or U9452 (N_9452,N_7776,N_8263);
nor U9453 (N_9453,N_7442,N_7596);
nor U9454 (N_9454,N_8310,N_7602);
nand U9455 (N_9455,N_7809,N_8117);
nor U9456 (N_9456,N_8047,N_7842);
and U9457 (N_9457,N_8232,N_8388);
nor U9458 (N_9458,N_7961,N_7903);
nor U9459 (N_9459,N_7673,N_7431);
xor U9460 (N_9460,N_7983,N_7992);
nand U9461 (N_9461,N_7450,N_8243);
and U9462 (N_9462,N_7726,N_7929);
xor U9463 (N_9463,N_8352,N_7999);
xnor U9464 (N_9464,N_8341,N_8206);
nand U9465 (N_9465,N_8221,N_7258);
nor U9466 (N_9466,N_7851,N_8168);
and U9467 (N_9467,N_8329,N_8350);
nor U9468 (N_9468,N_7518,N_8311);
nand U9469 (N_9469,N_7968,N_7851);
nand U9470 (N_9470,N_8061,N_7650);
or U9471 (N_9471,N_7462,N_7204);
xor U9472 (N_9472,N_7279,N_7403);
xor U9473 (N_9473,N_8254,N_7983);
and U9474 (N_9474,N_7862,N_8352);
and U9475 (N_9475,N_7801,N_7997);
nand U9476 (N_9476,N_8186,N_7672);
nand U9477 (N_9477,N_7652,N_7666);
nor U9478 (N_9478,N_8128,N_7842);
nand U9479 (N_9479,N_8186,N_7237);
nand U9480 (N_9480,N_8169,N_8018);
and U9481 (N_9481,N_7483,N_7831);
nand U9482 (N_9482,N_7797,N_7500);
and U9483 (N_9483,N_8051,N_8088);
nand U9484 (N_9484,N_7879,N_7823);
nand U9485 (N_9485,N_8122,N_7580);
xor U9486 (N_9486,N_7944,N_7283);
and U9487 (N_9487,N_7387,N_7586);
and U9488 (N_9488,N_7518,N_7256);
nand U9489 (N_9489,N_7647,N_7542);
nor U9490 (N_9490,N_7645,N_8048);
nor U9491 (N_9491,N_7470,N_7460);
xnor U9492 (N_9492,N_7364,N_8215);
or U9493 (N_9493,N_8222,N_7270);
xor U9494 (N_9494,N_8112,N_7292);
and U9495 (N_9495,N_7318,N_8009);
and U9496 (N_9496,N_7938,N_7435);
nor U9497 (N_9497,N_7691,N_8224);
xnor U9498 (N_9498,N_7680,N_7558);
xor U9499 (N_9499,N_7610,N_7249);
nand U9500 (N_9500,N_7754,N_7364);
and U9501 (N_9501,N_7871,N_7616);
nor U9502 (N_9502,N_7853,N_8296);
xor U9503 (N_9503,N_8094,N_7577);
nand U9504 (N_9504,N_8241,N_7772);
and U9505 (N_9505,N_7446,N_7266);
nor U9506 (N_9506,N_8205,N_8005);
and U9507 (N_9507,N_7402,N_7915);
or U9508 (N_9508,N_7561,N_8327);
or U9509 (N_9509,N_7876,N_7897);
nor U9510 (N_9510,N_7229,N_7657);
nand U9511 (N_9511,N_8196,N_7246);
nand U9512 (N_9512,N_7435,N_7910);
nand U9513 (N_9513,N_7203,N_7407);
xor U9514 (N_9514,N_7669,N_7638);
xor U9515 (N_9515,N_8039,N_7273);
xor U9516 (N_9516,N_8207,N_7956);
xnor U9517 (N_9517,N_7762,N_7661);
xnor U9518 (N_9518,N_7783,N_7211);
xor U9519 (N_9519,N_8394,N_7652);
and U9520 (N_9520,N_7281,N_8164);
nand U9521 (N_9521,N_7420,N_8218);
xor U9522 (N_9522,N_7677,N_7656);
or U9523 (N_9523,N_8208,N_8266);
nand U9524 (N_9524,N_7425,N_8308);
xnor U9525 (N_9525,N_8173,N_7505);
or U9526 (N_9526,N_7285,N_7362);
nor U9527 (N_9527,N_7383,N_8369);
and U9528 (N_9528,N_7642,N_7251);
xor U9529 (N_9529,N_7525,N_7475);
xor U9530 (N_9530,N_7280,N_8113);
or U9531 (N_9531,N_7944,N_7987);
nor U9532 (N_9532,N_8262,N_7499);
nand U9533 (N_9533,N_8129,N_8297);
and U9534 (N_9534,N_7572,N_8065);
xor U9535 (N_9535,N_8373,N_8353);
xnor U9536 (N_9536,N_7272,N_7397);
and U9537 (N_9537,N_8275,N_8245);
xnor U9538 (N_9538,N_7269,N_7389);
and U9539 (N_9539,N_7521,N_7418);
nor U9540 (N_9540,N_8372,N_8290);
and U9541 (N_9541,N_7317,N_8374);
xor U9542 (N_9542,N_7490,N_8182);
or U9543 (N_9543,N_8217,N_7337);
or U9544 (N_9544,N_7655,N_7228);
xor U9545 (N_9545,N_7348,N_7638);
xor U9546 (N_9546,N_7730,N_8265);
and U9547 (N_9547,N_7452,N_7947);
and U9548 (N_9548,N_7867,N_7455);
nand U9549 (N_9549,N_7401,N_8174);
and U9550 (N_9550,N_8062,N_7630);
nand U9551 (N_9551,N_8350,N_8370);
xor U9552 (N_9552,N_8314,N_7301);
xnor U9553 (N_9553,N_7910,N_7724);
or U9554 (N_9554,N_7439,N_7228);
xnor U9555 (N_9555,N_7824,N_8264);
and U9556 (N_9556,N_7707,N_7655);
and U9557 (N_9557,N_8358,N_7666);
nor U9558 (N_9558,N_8046,N_7721);
or U9559 (N_9559,N_7944,N_7289);
nand U9560 (N_9560,N_8124,N_7687);
xnor U9561 (N_9561,N_7332,N_8391);
and U9562 (N_9562,N_7392,N_7804);
nand U9563 (N_9563,N_7934,N_7596);
or U9564 (N_9564,N_7801,N_7284);
nor U9565 (N_9565,N_8233,N_7997);
or U9566 (N_9566,N_8011,N_7646);
xor U9567 (N_9567,N_8065,N_7823);
and U9568 (N_9568,N_7421,N_7727);
nor U9569 (N_9569,N_7851,N_8371);
nand U9570 (N_9570,N_7915,N_8102);
xnor U9571 (N_9571,N_7254,N_7233);
nor U9572 (N_9572,N_8251,N_8258);
xnor U9573 (N_9573,N_7808,N_7738);
and U9574 (N_9574,N_7245,N_7785);
nand U9575 (N_9575,N_7256,N_7657);
xor U9576 (N_9576,N_7706,N_8119);
or U9577 (N_9577,N_7230,N_8220);
nand U9578 (N_9578,N_7364,N_8059);
nand U9579 (N_9579,N_7610,N_7985);
nor U9580 (N_9580,N_8095,N_7293);
or U9581 (N_9581,N_8285,N_7574);
nand U9582 (N_9582,N_7681,N_7442);
xnor U9583 (N_9583,N_7590,N_7233);
xor U9584 (N_9584,N_7958,N_7233);
nand U9585 (N_9585,N_7611,N_8352);
and U9586 (N_9586,N_7822,N_7316);
nand U9587 (N_9587,N_7901,N_7509);
and U9588 (N_9588,N_8091,N_8359);
and U9589 (N_9589,N_8289,N_7977);
nand U9590 (N_9590,N_7377,N_7663);
nand U9591 (N_9591,N_7587,N_7310);
and U9592 (N_9592,N_7588,N_7551);
xor U9593 (N_9593,N_7923,N_7778);
and U9594 (N_9594,N_7972,N_7747);
xor U9595 (N_9595,N_8239,N_7540);
xnor U9596 (N_9596,N_8395,N_7574);
xnor U9597 (N_9597,N_7437,N_7228);
nor U9598 (N_9598,N_7485,N_8333);
xnor U9599 (N_9599,N_7219,N_7281);
nand U9600 (N_9600,N_9550,N_8976);
and U9601 (N_9601,N_8959,N_8771);
nor U9602 (N_9602,N_8729,N_8979);
or U9603 (N_9603,N_8928,N_9314);
or U9604 (N_9604,N_8423,N_8691);
nand U9605 (N_9605,N_8457,N_9052);
nor U9606 (N_9606,N_8692,N_8820);
or U9607 (N_9607,N_9551,N_8527);
nand U9608 (N_9608,N_9020,N_8806);
and U9609 (N_9609,N_8433,N_9050);
or U9610 (N_9610,N_8921,N_9036);
or U9611 (N_9611,N_8802,N_9261);
and U9612 (N_9612,N_9543,N_8980);
or U9613 (N_9613,N_8634,N_9523);
nor U9614 (N_9614,N_9114,N_8572);
nand U9615 (N_9615,N_8695,N_8738);
xor U9616 (N_9616,N_8799,N_9084);
xnor U9617 (N_9617,N_9099,N_9258);
or U9618 (N_9618,N_9026,N_9087);
or U9619 (N_9619,N_9493,N_8599);
or U9620 (N_9620,N_9484,N_8822);
nand U9621 (N_9621,N_9411,N_9363);
xor U9622 (N_9622,N_9143,N_8908);
and U9623 (N_9623,N_9081,N_9358);
nand U9624 (N_9624,N_8580,N_8535);
xnor U9625 (N_9625,N_9098,N_8410);
and U9626 (N_9626,N_9240,N_9175);
or U9627 (N_9627,N_9513,N_8663);
or U9628 (N_9628,N_9279,N_8923);
nor U9629 (N_9629,N_9421,N_9443);
nand U9630 (N_9630,N_8826,N_8918);
xor U9631 (N_9631,N_9217,N_9044);
nor U9632 (N_9632,N_9569,N_9480);
xnor U9633 (N_9633,N_8586,N_8462);
or U9634 (N_9634,N_8636,N_9366);
nor U9635 (N_9635,N_8547,N_8884);
and U9636 (N_9636,N_9268,N_8801);
nand U9637 (N_9637,N_8704,N_9278);
nor U9638 (N_9638,N_9133,N_9365);
xnor U9639 (N_9639,N_9283,N_9341);
and U9640 (N_9640,N_8513,N_9520);
nand U9641 (N_9641,N_9518,N_8606);
nand U9642 (N_9642,N_9066,N_8510);
nand U9643 (N_9643,N_9599,N_9459);
nor U9644 (N_9644,N_9515,N_8879);
and U9645 (N_9645,N_8521,N_9220);
nand U9646 (N_9646,N_9414,N_9121);
nor U9647 (N_9647,N_9410,N_9457);
nor U9648 (N_9648,N_9348,N_9262);
xnor U9649 (N_9649,N_9510,N_9222);
xor U9650 (N_9650,N_8565,N_8772);
and U9651 (N_9651,N_8867,N_8914);
nor U9652 (N_9652,N_9406,N_9325);
xnor U9653 (N_9653,N_9051,N_9159);
xnor U9654 (N_9654,N_8898,N_8966);
nor U9655 (N_9655,N_9548,N_8637);
xor U9656 (N_9656,N_8829,N_9196);
or U9657 (N_9657,N_9106,N_9233);
or U9658 (N_9658,N_8456,N_9445);
nand U9659 (N_9659,N_8983,N_9304);
and U9660 (N_9660,N_9075,N_9473);
nand U9661 (N_9661,N_8870,N_9108);
nor U9662 (N_9662,N_9113,N_8842);
nor U9663 (N_9663,N_8759,N_9500);
or U9664 (N_9664,N_9049,N_9151);
nor U9665 (N_9665,N_8899,N_8640);
and U9666 (N_9666,N_8552,N_9112);
xor U9667 (N_9667,N_8762,N_8485);
and U9668 (N_9668,N_9491,N_9389);
or U9669 (N_9669,N_9057,N_8502);
and U9670 (N_9670,N_8935,N_8698);
and U9671 (N_9671,N_9387,N_8962);
and U9672 (N_9672,N_9572,N_8769);
and U9673 (N_9673,N_8894,N_9489);
or U9674 (N_9674,N_8872,N_9536);
xor U9675 (N_9675,N_9352,N_9012);
and U9676 (N_9676,N_9298,N_9203);
or U9677 (N_9677,N_9176,N_9211);
xnor U9678 (N_9678,N_9091,N_9474);
xnor U9679 (N_9679,N_8434,N_9557);
and U9680 (N_9680,N_8618,N_9360);
nand U9681 (N_9681,N_9527,N_9055);
nor U9682 (N_9682,N_8722,N_8600);
and U9683 (N_9683,N_8517,N_9568);
nor U9684 (N_9684,N_9280,N_9157);
nand U9685 (N_9685,N_8814,N_8533);
nor U9686 (N_9686,N_8505,N_9169);
nand U9687 (N_9687,N_8597,N_9249);
nor U9688 (N_9688,N_8626,N_8913);
nand U9689 (N_9689,N_8825,N_8731);
xnor U9690 (N_9690,N_8590,N_8972);
xor U9691 (N_9691,N_9531,N_8708);
or U9692 (N_9692,N_8654,N_9244);
nor U9693 (N_9693,N_8986,N_9229);
nand U9694 (N_9694,N_8447,N_8699);
xor U9695 (N_9695,N_9228,N_9102);
and U9696 (N_9696,N_9180,N_8649);
nor U9697 (N_9697,N_8668,N_8483);
nor U9698 (N_9698,N_8886,N_9528);
nor U9699 (N_9699,N_9463,N_9533);
xor U9700 (N_9700,N_8922,N_9552);
nor U9701 (N_9701,N_9303,N_9342);
and U9702 (N_9702,N_8897,N_8561);
and U9703 (N_9703,N_8439,N_8556);
nor U9704 (N_9704,N_8581,N_9456);
nand U9705 (N_9705,N_9596,N_9440);
nand U9706 (N_9706,N_8920,N_8763);
nor U9707 (N_9707,N_8819,N_9574);
nand U9708 (N_9708,N_8518,N_8719);
nor U9709 (N_9709,N_9269,N_8460);
and U9710 (N_9710,N_8846,N_9589);
xor U9711 (N_9711,N_8474,N_9183);
or U9712 (N_9712,N_8427,N_8723);
nand U9713 (N_9713,N_9471,N_8416);
nor U9714 (N_9714,N_8896,N_8602);
nand U9715 (N_9715,N_9423,N_8747);
nand U9716 (N_9716,N_9067,N_9093);
nor U9717 (N_9717,N_9582,N_8875);
nand U9718 (N_9718,N_9311,N_8508);
nand U9719 (N_9719,N_9204,N_9148);
and U9720 (N_9720,N_8690,N_8671);
and U9721 (N_9721,N_8868,N_9470);
nor U9722 (N_9722,N_8828,N_8871);
xnor U9723 (N_9723,N_9281,N_9409);
or U9724 (N_9724,N_9320,N_9058);
nand U9725 (N_9725,N_8628,N_8987);
nand U9726 (N_9726,N_8546,N_9018);
xnor U9727 (N_9727,N_9561,N_8481);
xor U9728 (N_9728,N_8638,N_9434);
nor U9729 (N_9729,N_8467,N_9144);
nor U9730 (N_9730,N_9535,N_8707);
and U9731 (N_9731,N_9318,N_9184);
nor U9732 (N_9732,N_8815,N_8993);
nand U9733 (N_9733,N_9152,N_8619);
and U9734 (N_9734,N_9327,N_8499);
xor U9735 (N_9735,N_9210,N_9402);
and U9736 (N_9736,N_8404,N_8865);
and U9737 (N_9737,N_8851,N_8977);
and U9738 (N_9738,N_9002,N_8720);
or U9739 (N_9739,N_8516,N_8412);
and U9740 (N_9740,N_8841,N_8685);
nor U9741 (N_9741,N_9054,N_9138);
nor U9742 (N_9742,N_8680,N_8906);
nand U9743 (N_9743,N_9161,N_8482);
and U9744 (N_9744,N_9401,N_9413);
or U9745 (N_9745,N_9014,N_9154);
xnor U9746 (N_9746,N_9511,N_9442);
or U9747 (N_9747,N_8807,N_9212);
xor U9748 (N_9748,N_8578,N_9068);
or U9749 (N_9749,N_8804,N_8643);
nor U9750 (N_9750,N_8528,N_8893);
nand U9751 (N_9751,N_9499,N_9532);
and U9752 (N_9752,N_9034,N_9408);
xnor U9753 (N_9753,N_8647,N_8553);
xnor U9754 (N_9754,N_8607,N_8971);
xor U9755 (N_9755,N_8682,N_9005);
or U9756 (N_9756,N_8464,N_9386);
nor U9757 (N_9757,N_8453,N_8421);
nand U9758 (N_9758,N_9150,N_8796);
xnor U9759 (N_9759,N_9553,N_9284);
nand U9760 (N_9760,N_8673,N_9469);
nand U9761 (N_9761,N_9255,N_8919);
or U9762 (N_9762,N_8610,N_9243);
nand U9763 (N_9763,N_9416,N_8672);
and U9764 (N_9764,N_8444,N_9396);
and U9765 (N_9765,N_9064,N_9481);
nor U9766 (N_9766,N_9129,N_9179);
or U9767 (N_9767,N_9526,N_9429);
or U9768 (N_9768,N_8902,N_8549);
nor U9769 (N_9769,N_9374,N_9424);
nand U9770 (N_9770,N_8950,N_9251);
nand U9771 (N_9771,N_9156,N_9449);
nor U9772 (N_9772,N_9508,N_9274);
nand U9773 (N_9773,N_9357,N_8495);
and U9774 (N_9774,N_9497,N_9462);
and U9775 (N_9775,N_8443,N_9019);
or U9776 (N_9776,N_8625,N_8570);
nor U9777 (N_9777,N_8728,N_8531);
xor U9778 (N_9778,N_9525,N_9011);
nand U9779 (N_9779,N_9206,N_8784);
nand U9780 (N_9780,N_8895,N_8657);
or U9781 (N_9781,N_8718,N_8938);
nand U9782 (N_9782,N_8587,N_8413);
or U9783 (N_9783,N_8449,N_8835);
nand U9784 (N_9784,N_8681,N_8764);
nor U9785 (N_9785,N_8515,N_9082);
nor U9786 (N_9786,N_9571,N_8730);
and U9787 (N_9787,N_9071,N_8860);
or U9788 (N_9788,N_9017,N_9534);
nand U9789 (N_9789,N_8454,N_9453);
and U9790 (N_9790,N_9090,N_8949);
or U9791 (N_9791,N_8611,N_8645);
or U9792 (N_9792,N_9105,N_9267);
and U9793 (N_9793,N_8770,N_9062);
nand U9794 (N_9794,N_9549,N_9023);
xor U9795 (N_9795,N_8658,N_8970);
xor U9796 (N_9796,N_9297,N_8455);
nand U9797 (N_9797,N_9016,N_9502);
nor U9798 (N_9798,N_9438,N_8544);
nor U9799 (N_9799,N_8800,N_8887);
nor U9800 (N_9800,N_8736,N_8900);
and U9801 (N_9801,N_9422,N_9496);
xnor U9802 (N_9802,N_8543,N_8992);
xnor U9803 (N_9803,N_9448,N_9486);
xor U9804 (N_9804,N_9466,N_8735);
and U9805 (N_9805,N_8727,N_8609);
xor U9806 (N_9806,N_8836,N_8995);
xnor U9807 (N_9807,N_9592,N_9213);
nand U9808 (N_9808,N_9173,N_8538);
nor U9809 (N_9809,N_9001,N_8585);
nand U9810 (N_9810,N_9273,N_8402);
nand U9811 (N_9811,N_9194,N_8952);
or U9812 (N_9812,N_9230,N_8661);
xnor U9813 (N_9813,N_9293,N_9163);
nand U9814 (N_9814,N_9003,N_8700);
nor U9815 (N_9815,N_9364,N_9392);
and U9816 (N_9816,N_9200,N_8984);
nor U9817 (N_9817,N_9123,N_8598);
or U9818 (N_9818,N_9332,N_9588);
xor U9819 (N_9819,N_8582,N_9047);
nand U9820 (N_9820,N_8981,N_9381);
or U9821 (N_9821,N_8562,N_8617);
and U9822 (N_9822,N_8519,N_8997);
and U9823 (N_9823,N_9495,N_8678);
nand U9824 (N_9824,N_8400,N_8750);
nor U9825 (N_9825,N_9485,N_8646);
or U9826 (N_9826,N_8431,N_9346);
or U9827 (N_9827,N_9247,N_9048);
xor U9828 (N_9828,N_9376,N_8666);
nor U9829 (N_9829,N_8808,N_8930);
nor U9830 (N_9830,N_8780,N_8653);
xor U9831 (N_9831,N_9450,N_9333);
nor U9832 (N_9832,N_9007,N_8885);
nand U9833 (N_9833,N_9239,N_9216);
nor U9834 (N_9834,N_8717,N_9288);
nand U9835 (N_9835,N_8667,N_8901);
xnor U9836 (N_9836,N_9107,N_9464);
nor U9837 (N_9837,N_9115,N_9174);
nand U9838 (N_9838,N_8845,N_9033);
and U9839 (N_9839,N_9256,N_9570);
nor U9840 (N_9840,N_8838,N_9029);
and U9841 (N_9841,N_9291,N_9382);
or U9842 (N_9842,N_9286,N_9289);
xor U9843 (N_9843,N_8969,N_8407);
nor U9844 (N_9844,N_8492,N_8737);
and U9845 (N_9845,N_9146,N_8861);
or U9846 (N_9846,N_9336,N_9509);
xor U9847 (N_9847,N_8506,N_9529);
nand U9848 (N_9848,N_9544,N_8855);
nand U9849 (N_9849,N_9403,N_8739);
xnor U9850 (N_9850,N_9324,N_8837);
xnor U9851 (N_9851,N_8624,N_9488);
and U9852 (N_9852,N_8631,N_8493);
or U9853 (N_9853,N_9076,N_8792);
nand U9854 (N_9854,N_9294,N_8560);
xnor U9855 (N_9855,N_9141,N_9328);
xnor U9856 (N_9856,N_9454,N_9516);
nor U9857 (N_9857,N_9323,N_9142);
nand U9858 (N_9858,N_9171,N_9235);
nand U9859 (N_9859,N_8675,N_9172);
or U9860 (N_9860,N_9338,N_8452);
and U9861 (N_9861,N_9501,N_8445);
nand U9862 (N_9862,N_8534,N_8891);
or U9863 (N_9863,N_8583,N_8787);
and U9864 (N_9864,N_9285,N_9162);
and U9865 (N_9865,N_9398,N_8994);
nor U9866 (N_9866,N_8496,N_9306);
xor U9867 (N_9867,N_8881,N_8512);
nor U9868 (N_9868,N_9095,N_9227);
and U9869 (N_9869,N_9420,N_9461);
nor U9870 (N_9870,N_9008,N_9197);
xnor U9871 (N_9871,N_9575,N_9043);
nand U9872 (N_9872,N_8405,N_9242);
xor U9873 (N_9873,N_9475,N_8766);
xnor U9874 (N_9874,N_9132,N_9326);
or U9875 (N_9875,N_8810,N_8864);
or U9876 (N_9876,N_8555,N_9096);
xor U9877 (N_9877,N_9193,N_9140);
or U9878 (N_9878,N_9388,N_9340);
or U9879 (N_9879,N_9158,N_9208);
and U9880 (N_9880,N_9214,N_8797);
xnor U9881 (N_9881,N_9110,N_8978);
or U9882 (N_9882,N_8805,N_8890);
or U9883 (N_9883,N_8406,N_9329);
nor U9884 (N_9884,N_8662,N_8710);
or U9885 (N_9885,N_9103,N_8541);
nand U9886 (N_9886,N_9195,N_9094);
xnor U9887 (N_9887,N_9165,N_9209);
nor U9888 (N_9888,N_9545,N_8594);
or U9889 (N_9889,N_8589,N_8451);
nor U9890 (N_9890,N_8752,N_9584);
and U9891 (N_9891,N_9595,N_8988);
xor U9892 (N_9892,N_8593,N_9554);
xor U9893 (N_9893,N_9476,N_9296);
nor U9894 (N_9894,N_8403,N_8569);
or U9895 (N_9895,N_8478,N_8740);
and U9896 (N_9896,N_9586,N_9125);
xnor U9897 (N_9897,N_8694,N_9519);
nand U9898 (N_9898,N_9149,N_9512);
nor U9899 (N_9899,N_9417,N_8644);
nand U9900 (N_9900,N_9116,N_9562);
and U9901 (N_9901,N_8982,N_9503);
nand U9902 (N_9902,N_9455,N_8847);
or U9903 (N_9903,N_9373,N_8605);
nand U9904 (N_9904,N_8776,N_8854);
nand U9905 (N_9905,N_9577,N_9594);
nand U9906 (N_9906,N_8741,N_9100);
and U9907 (N_9907,N_9547,N_8862);
nand U9908 (N_9908,N_9394,N_8973);
nand U9909 (N_9909,N_8765,N_8470);
nand U9910 (N_9910,N_9038,N_9130);
nor U9911 (N_9911,N_9137,N_9418);
nor U9912 (N_9912,N_8777,N_8999);
nor U9913 (N_9913,N_9271,N_9282);
xor U9914 (N_9914,N_8857,N_9122);
or U9915 (N_9915,N_8912,N_9167);
and U9916 (N_9916,N_8614,N_9343);
xnor U9917 (N_9917,N_8726,N_8967);
or U9918 (N_9918,N_8778,N_8830);
xor U9919 (N_9919,N_9522,N_8848);
or U9920 (N_9920,N_9433,N_9042);
nand U9921 (N_9921,N_8724,N_8612);
xor U9922 (N_9922,N_9590,N_8469);
nor U9923 (N_9923,N_9567,N_8486);
xnor U9924 (N_9924,N_8501,N_9031);
or U9925 (N_9925,N_8448,N_8831);
nor U9926 (N_9926,N_9315,N_8925);
xor U9927 (N_9927,N_8428,N_9539);
and U9928 (N_9928,N_9300,N_9063);
xnor U9929 (N_9929,N_9040,N_8783);
nand U9930 (N_9930,N_9482,N_9128);
xor U9931 (N_9931,N_9065,N_8911);
or U9932 (N_9932,N_8852,N_8441);
nor U9933 (N_9933,N_8859,N_8409);
xor U9934 (N_9934,N_9452,N_8623);
nor U9935 (N_9935,N_8774,N_8715);
xnor U9936 (N_9936,N_8954,N_9467);
or U9937 (N_9937,N_9056,N_9494);
nand U9938 (N_9938,N_9117,N_9419);
and U9939 (N_9939,N_8823,N_8615);
and U9940 (N_9940,N_8839,N_9415);
nand U9941 (N_9941,N_9219,N_9407);
and U9942 (N_9942,N_8748,N_9263);
xor U9943 (N_9943,N_9218,N_9236);
nand U9944 (N_9944,N_9435,N_9560);
or U9945 (N_9945,N_9257,N_8604);
nor U9946 (N_9946,N_8436,N_9565);
nor U9947 (N_9947,N_9556,N_8500);
nor U9948 (N_9948,N_8768,N_9041);
xnor U9949 (N_9949,N_9337,N_9231);
nand U9950 (N_9950,N_8817,N_9277);
nor U9951 (N_9951,N_8514,N_8757);
nor U9952 (N_9952,N_8834,N_9238);
xor U9953 (N_9953,N_8688,N_8917);
or U9954 (N_9954,N_9004,N_8511);
xnor U9955 (N_9955,N_8889,N_8781);
and U9956 (N_9956,N_9182,N_8963);
nor U9957 (N_9957,N_8559,N_9367);
and U9958 (N_9958,N_8964,N_9444);
nor U9959 (N_9959,N_9412,N_9426);
or U9960 (N_9960,N_8670,N_9591);
nand U9961 (N_9961,N_9368,N_8696);
or U9962 (N_9962,N_8761,N_9505);
and U9963 (N_9963,N_8442,N_8713);
nor U9964 (N_9964,N_8705,N_9432);
xnor U9965 (N_9965,N_8480,N_8677);
and U9966 (N_9966,N_8866,N_8721);
or U9967 (N_9967,N_8795,N_8659);
nand U9968 (N_9968,N_8725,N_8960);
nor U9969 (N_9969,N_9436,N_9555);
or U9970 (N_9970,N_9086,N_9395);
nand U9971 (N_9971,N_8803,N_8465);
or U9972 (N_9972,N_9478,N_8429);
or U9973 (N_9973,N_9399,N_9237);
nand U9974 (N_9974,N_8522,N_9524);
and U9975 (N_9975,N_9439,N_8786);
and U9976 (N_9976,N_9380,N_8782);
nor U9977 (N_9977,N_8793,N_8655);
xor U9978 (N_9978,N_9224,N_9379);
and U9979 (N_9979,N_9232,N_8557);
nor U9980 (N_9980,N_9160,N_8509);
or U9981 (N_9981,N_8882,N_9192);
nand U9982 (N_9982,N_9085,N_8932);
xnor U9983 (N_9983,N_8525,N_8990);
and U9984 (N_9984,N_9354,N_8595);
or U9985 (N_9985,N_9223,N_9177);
nor U9986 (N_9986,N_9427,N_9404);
or U9987 (N_9987,N_9088,N_9468);
nor U9988 (N_9988,N_8948,N_9301);
nor U9989 (N_9989,N_8651,N_9207);
xnor U9990 (N_9990,N_8955,N_8697);
or U9991 (N_9991,N_8498,N_8812);
xor U9992 (N_9992,N_9009,N_8743);
xor U9993 (N_9993,N_8459,N_9583);
xnor U9994 (N_9994,N_8532,N_9073);
nor U9995 (N_9995,N_8419,N_8751);
nand U9996 (N_9996,N_9250,N_8648);
and U9997 (N_9997,N_9507,N_9506);
nand U9998 (N_9998,N_9126,N_9101);
xnor U9999 (N_9999,N_9027,N_8975);
or U10000 (N_10000,N_8432,N_9225);
and U10001 (N_10001,N_9135,N_8596);
nand U10002 (N_10002,N_9290,N_9241);
or U10003 (N_10003,N_9292,N_8539);
or U10004 (N_10004,N_8430,N_8484);
xor U10005 (N_10005,N_8703,N_8475);
xor U10006 (N_10006,N_9369,N_9362);
xnor U10007 (N_10007,N_9430,N_8907);
or U10008 (N_10008,N_8622,N_9349);
xnor U10009 (N_10009,N_8758,N_9472);
and U10010 (N_10010,N_8524,N_8903);
xor U10011 (N_10011,N_9356,N_8756);
nand U10012 (N_10012,N_9181,N_9202);
nor U10013 (N_10013,N_9264,N_9564);
nor U10014 (N_10014,N_9542,N_8669);
or U10015 (N_10015,N_8712,N_8507);
nor U10016 (N_10016,N_8746,N_9024);
nand U10017 (N_10017,N_8934,N_8745);
or U10018 (N_10018,N_8620,N_9390);
or U10019 (N_10019,N_9490,N_9437);
and U10020 (N_10020,N_9078,N_9254);
or U10021 (N_10021,N_9347,N_9118);
nand U10022 (N_10022,N_8933,N_8520);
nand U10023 (N_10023,N_9317,N_8754);
nor U10024 (N_10024,N_8536,N_8601);
and U10025 (N_10025,N_9393,N_9322);
nand U10026 (N_10026,N_8813,N_9581);
or U10027 (N_10027,N_8961,N_8686);
or U10028 (N_10028,N_9199,N_8755);
or U10029 (N_10029,N_9309,N_8974);
nor U10030 (N_10030,N_9372,N_9191);
nand U10031 (N_10031,N_8943,N_8956);
nand U10032 (N_10032,N_8650,N_9587);
xnor U10033 (N_10033,N_9385,N_8479);
and U10034 (N_10034,N_9307,N_8711);
and U10035 (N_10035,N_9080,N_9010);
and U10036 (N_10036,N_8489,N_9030);
nor U10037 (N_10037,N_8588,N_9580);
or U10038 (N_10038,N_9053,N_8660);
and U10039 (N_10039,N_8608,N_9546);
and U10040 (N_10040,N_9119,N_9573);
nand U10041 (N_10041,N_9344,N_9425);
or U10042 (N_10042,N_9397,N_9166);
nor U10043 (N_10043,N_9391,N_9313);
nor U10044 (N_10044,N_8575,N_8629);
or U10045 (N_10045,N_8497,N_9245);
nor U10046 (N_10046,N_9310,N_8676);
xnor U10047 (N_10047,N_8942,N_9517);
nor U10048 (N_10048,N_9234,N_8440);
nand U10049 (N_10049,N_8714,N_9089);
xor U10050 (N_10050,N_8450,N_9566);
or U10051 (N_10051,N_9266,N_9120);
and U10052 (N_10052,N_8744,N_8415);
and U10053 (N_10053,N_8577,N_8850);
nor U10054 (N_10054,N_8927,N_9046);
and U10055 (N_10055,N_8947,N_9127);
nor U10056 (N_10056,N_8526,N_8853);
and U10057 (N_10057,N_9465,N_9074);
nand U10058 (N_10058,N_8785,N_8689);
nor U10059 (N_10059,N_9492,N_9097);
nor U10060 (N_10060,N_8566,N_8537);
and U10061 (N_10061,N_8563,N_8833);
nor U10062 (N_10062,N_8953,N_9272);
nand U10063 (N_10063,N_8869,N_9477);
nor U10064 (N_10064,N_9335,N_9032);
xnor U10065 (N_10065,N_8701,N_8422);
xor U10066 (N_10066,N_9308,N_9006);
nor U10067 (N_10067,N_8584,N_8471);
nand U10068 (N_10068,N_9275,N_9483);
or U10069 (N_10069,N_8767,N_9000);
and U10070 (N_10070,N_8488,N_9530);
nor U10071 (N_10071,N_8656,N_9215);
nor U10072 (N_10072,N_9375,N_8627);
xor U10073 (N_10073,N_8466,N_8883);
or U10074 (N_10074,N_9072,N_9060);
nor U10075 (N_10075,N_9331,N_8926);
and U10076 (N_10076,N_8840,N_9538);
and U10077 (N_10077,N_8929,N_8408);
and U10078 (N_10078,N_9384,N_9321);
and U10079 (N_10079,N_9460,N_9541);
nand U10080 (N_10080,N_9164,N_8702);
or U10081 (N_10081,N_9104,N_9059);
or U10082 (N_10082,N_8924,N_8733);
and U10083 (N_10083,N_8591,N_8693);
or U10084 (N_10084,N_9248,N_9521);
nand U10085 (N_10085,N_8679,N_8574);
and U10086 (N_10086,N_8414,N_9037);
nand U10087 (N_10087,N_8821,N_8437);
and U10088 (N_10088,N_9198,N_8642);
nand U10089 (N_10089,N_8827,N_9265);
and U10090 (N_10090,N_8775,N_8844);
xnor U10091 (N_10091,N_9170,N_9371);
and U10092 (N_10092,N_8571,N_9260);
and U10093 (N_10093,N_8939,N_8540);
or U10094 (N_10094,N_8424,N_9186);
nor U10095 (N_10095,N_9147,N_8931);
and U10096 (N_10096,N_9270,N_8426);
nor U10097 (N_10097,N_8568,N_8576);
nand U10098 (N_10098,N_9334,N_8458);
nor U10099 (N_10099,N_8832,N_8550);
nand U10100 (N_10100,N_9124,N_9134);
and U10101 (N_10101,N_8916,N_8791);
and U10102 (N_10102,N_8665,N_8753);
or U10103 (N_10103,N_9319,N_9070);
nor U10104 (N_10104,N_8567,N_9045);
nand U10105 (N_10105,N_8417,N_9537);
or U10106 (N_10106,N_8909,N_8811);
nand U10107 (N_10107,N_9405,N_9446);
xnor U10108 (N_10108,N_9178,N_8749);
xnor U10109 (N_10109,N_8818,N_8683);
xor U10110 (N_10110,N_8888,N_8530);
and U10111 (N_10111,N_8630,N_8674);
or U10112 (N_10112,N_8874,N_8613);
xor U10113 (N_10113,N_8968,N_8989);
nor U10114 (N_10114,N_8732,N_8946);
or U10115 (N_10115,N_8878,N_9109);
nor U10116 (N_10116,N_8788,N_8529);
and U10117 (N_10117,N_8876,N_8504);
xnor U10118 (N_10118,N_9131,N_8463);
xor U10119 (N_10119,N_9441,N_8472);
and U10120 (N_10120,N_9377,N_9593);
and U10121 (N_10121,N_9155,N_8418);
xor U10122 (N_10122,N_9400,N_8773);
nand U10123 (N_10123,N_8554,N_8476);
and U10124 (N_10124,N_9350,N_9190);
and U10125 (N_10125,N_8490,N_8635);
or U10126 (N_10126,N_8632,N_8706);
or U10127 (N_10127,N_8491,N_9359);
or U10128 (N_10128,N_9153,N_8965);
nand U10129 (N_10129,N_9246,N_8816);
or U10130 (N_10130,N_8709,N_9339);
xor U10131 (N_10131,N_9077,N_9585);
and U10132 (N_10132,N_9383,N_8461);
nand U10133 (N_10133,N_9563,N_9498);
or U10134 (N_10134,N_9305,N_8446);
or U10135 (N_10135,N_9145,N_8542);
nand U10136 (N_10136,N_8824,N_9479);
and U10137 (N_10137,N_9035,N_8849);
nand U10138 (N_10138,N_9447,N_8880);
or U10139 (N_10139,N_9345,N_8548);
xnor U10140 (N_10140,N_8798,N_9597);
nor U10141 (N_10141,N_9069,N_8734);
xor U10142 (N_10142,N_9221,N_9428);
xnor U10143 (N_10143,N_8958,N_8633);
xnor U10144 (N_10144,N_9330,N_8425);
or U10145 (N_10145,N_8487,N_9458);
or U10146 (N_10146,N_8401,N_9361);
nor U10147 (N_10147,N_8742,N_8687);
nor U10148 (N_10148,N_9259,N_8941);
nor U10149 (N_10149,N_9504,N_9353);
nor U10150 (N_10150,N_8910,N_9111);
xor U10151 (N_10151,N_9201,N_9559);
and U10152 (N_10152,N_8435,N_9558);
nor U10153 (N_10153,N_8551,N_8621);
and U10154 (N_10154,N_9028,N_9287);
nand U10155 (N_10155,N_8477,N_8998);
and U10156 (N_10156,N_9578,N_8760);
and U10157 (N_10157,N_8473,N_8863);
xnor U10158 (N_10158,N_8592,N_8957);
xor U10159 (N_10159,N_9299,N_9514);
nor U10160 (N_10160,N_9185,N_8411);
nor U10161 (N_10161,N_9039,N_8873);
nor U10162 (N_10162,N_8789,N_9189);
or U10163 (N_10163,N_9540,N_8892);
or U10164 (N_10164,N_8951,N_9136);
and U10165 (N_10165,N_8503,N_8877);
and U10166 (N_10166,N_8468,N_8905);
xor U10167 (N_10167,N_8779,N_9576);
and U10168 (N_10168,N_8936,N_9015);
or U10169 (N_10169,N_8858,N_8985);
xnor U10170 (N_10170,N_8996,N_9451);
xor U10171 (N_10171,N_9487,N_9168);
xnor U10172 (N_10172,N_8991,N_9061);
or U10173 (N_10173,N_9139,N_8438);
nand U10174 (N_10174,N_8545,N_8716);
nand U10175 (N_10175,N_8420,N_9252);
xnor U10176 (N_10176,N_9205,N_8940);
xor U10177 (N_10177,N_9021,N_8904);
or U10178 (N_10178,N_9187,N_9092);
or U10179 (N_10179,N_8856,N_9276);
nand U10180 (N_10180,N_9079,N_9083);
and U10181 (N_10181,N_8794,N_8641);
xor U10182 (N_10182,N_8915,N_9312);
and U10183 (N_10183,N_8843,N_9295);
and U10184 (N_10184,N_9022,N_9226);
and U10185 (N_10185,N_8616,N_9378);
xnor U10186 (N_10186,N_8944,N_8639);
or U10187 (N_10187,N_9579,N_8558);
and U10188 (N_10188,N_9253,N_9302);
and U10189 (N_10189,N_8603,N_9370);
nand U10190 (N_10190,N_8494,N_9598);
xnor U10191 (N_10191,N_9188,N_9025);
nor U10192 (N_10192,N_8652,N_8945);
xnor U10193 (N_10193,N_8937,N_9316);
or U10194 (N_10194,N_8579,N_8664);
nor U10195 (N_10195,N_8523,N_9351);
xnor U10196 (N_10196,N_8684,N_8809);
nor U10197 (N_10197,N_9431,N_8564);
and U10198 (N_10198,N_9355,N_9013);
nand U10199 (N_10199,N_8790,N_8573);
xor U10200 (N_10200,N_8438,N_8904);
and U10201 (N_10201,N_9245,N_9215);
and U10202 (N_10202,N_9309,N_9138);
nand U10203 (N_10203,N_8843,N_8400);
and U10204 (N_10204,N_8990,N_8701);
nor U10205 (N_10205,N_8873,N_8675);
and U10206 (N_10206,N_8764,N_8465);
and U10207 (N_10207,N_8595,N_9098);
and U10208 (N_10208,N_8665,N_8883);
and U10209 (N_10209,N_8578,N_9492);
nand U10210 (N_10210,N_8708,N_8716);
or U10211 (N_10211,N_9311,N_9188);
nand U10212 (N_10212,N_9311,N_8598);
nor U10213 (N_10213,N_8804,N_8911);
and U10214 (N_10214,N_9499,N_9212);
nor U10215 (N_10215,N_9537,N_9088);
xor U10216 (N_10216,N_8771,N_9019);
nand U10217 (N_10217,N_9274,N_8883);
xnor U10218 (N_10218,N_8854,N_8658);
nor U10219 (N_10219,N_8926,N_8819);
nor U10220 (N_10220,N_9026,N_9110);
or U10221 (N_10221,N_9349,N_8743);
xor U10222 (N_10222,N_8543,N_8489);
or U10223 (N_10223,N_8476,N_9190);
and U10224 (N_10224,N_8768,N_8491);
xor U10225 (N_10225,N_9533,N_9478);
or U10226 (N_10226,N_9480,N_9283);
nor U10227 (N_10227,N_8696,N_8822);
xor U10228 (N_10228,N_8982,N_8576);
and U10229 (N_10229,N_9477,N_8978);
or U10230 (N_10230,N_8724,N_8519);
xor U10231 (N_10231,N_8817,N_9037);
xnor U10232 (N_10232,N_8561,N_9095);
or U10233 (N_10233,N_9416,N_9217);
nor U10234 (N_10234,N_8461,N_9158);
nand U10235 (N_10235,N_9192,N_8702);
xor U10236 (N_10236,N_9188,N_9596);
or U10237 (N_10237,N_8835,N_8618);
and U10238 (N_10238,N_8463,N_8780);
nand U10239 (N_10239,N_8516,N_8813);
nor U10240 (N_10240,N_8433,N_9151);
xor U10241 (N_10241,N_8790,N_9215);
xor U10242 (N_10242,N_9341,N_8725);
nor U10243 (N_10243,N_9365,N_9165);
and U10244 (N_10244,N_9377,N_9137);
nand U10245 (N_10245,N_9327,N_9368);
nand U10246 (N_10246,N_8768,N_9292);
xor U10247 (N_10247,N_9164,N_9099);
or U10248 (N_10248,N_9047,N_9465);
nor U10249 (N_10249,N_9464,N_9593);
nor U10250 (N_10250,N_9445,N_9033);
and U10251 (N_10251,N_9329,N_9326);
xor U10252 (N_10252,N_8918,N_9358);
xor U10253 (N_10253,N_9204,N_9267);
nand U10254 (N_10254,N_8846,N_9216);
nor U10255 (N_10255,N_9128,N_8988);
xnor U10256 (N_10256,N_9395,N_9055);
nor U10257 (N_10257,N_9070,N_8959);
nor U10258 (N_10258,N_9103,N_9396);
xor U10259 (N_10259,N_8904,N_9039);
and U10260 (N_10260,N_8689,N_8895);
nand U10261 (N_10261,N_9135,N_9521);
nand U10262 (N_10262,N_9485,N_9305);
nor U10263 (N_10263,N_9577,N_8943);
nor U10264 (N_10264,N_9199,N_8491);
or U10265 (N_10265,N_8656,N_9446);
xor U10266 (N_10266,N_9432,N_9434);
xnor U10267 (N_10267,N_9331,N_8905);
nand U10268 (N_10268,N_9020,N_9528);
or U10269 (N_10269,N_8818,N_8756);
nand U10270 (N_10270,N_8608,N_8781);
nor U10271 (N_10271,N_9065,N_8698);
xor U10272 (N_10272,N_8719,N_9166);
or U10273 (N_10273,N_8595,N_8597);
nand U10274 (N_10274,N_9409,N_9373);
nor U10275 (N_10275,N_8997,N_8748);
or U10276 (N_10276,N_9317,N_9168);
or U10277 (N_10277,N_9465,N_8599);
or U10278 (N_10278,N_8445,N_9114);
xor U10279 (N_10279,N_9589,N_9523);
xnor U10280 (N_10280,N_8670,N_8642);
or U10281 (N_10281,N_9099,N_8428);
xor U10282 (N_10282,N_8491,N_9196);
nor U10283 (N_10283,N_9139,N_8513);
xor U10284 (N_10284,N_8923,N_8629);
nand U10285 (N_10285,N_8697,N_9481);
nand U10286 (N_10286,N_9024,N_9137);
nand U10287 (N_10287,N_9290,N_9556);
nor U10288 (N_10288,N_9192,N_8412);
or U10289 (N_10289,N_9064,N_9334);
or U10290 (N_10290,N_9259,N_9197);
or U10291 (N_10291,N_8495,N_9177);
nand U10292 (N_10292,N_8956,N_8668);
or U10293 (N_10293,N_9540,N_8908);
or U10294 (N_10294,N_8699,N_9061);
nand U10295 (N_10295,N_8450,N_9340);
or U10296 (N_10296,N_9255,N_8497);
and U10297 (N_10297,N_8560,N_9154);
nand U10298 (N_10298,N_8894,N_9379);
or U10299 (N_10299,N_9135,N_8457);
nand U10300 (N_10300,N_8786,N_8708);
xor U10301 (N_10301,N_9292,N_9521);
xor U10302 (N_10302,N_9427,N_8989);
nand U10303 (N_10303,N_9044,N_9568);
nor U10304 (N_10304,N_9120,N_8994);
or U10305 (N_10305,N_8755,N_8907);
or U10306 (N_10306,N_8805,N_9535);
nand U10307 (N_10307,N_8453,N_8739);
or U10308 (N_10308,N_8778,N_8909);
nand U10309 (N_10309,N_9083,N_8828);
and U10310 (N_10310,N_8702,N_9468);
nor U10311 (N_10311,N_9402,N_8612);
and U10312 (N_10312,N_9262,N_8859);
nand U10313 (N_10313,N_9228,N_8747);
xnor U10314 (N_10314,N_9049,N_9311);
and U10315 (N_10315,N_8725,N_8930);
nand U10316 (N_10316,N_9386,N_8623);
xor U10317 (N_10317,N_8763,N_9227);
nor U10318 (N_10318,N_8595,N_8612);
nor U10319 (N_10319,N_8547,N_9403);
and U10320 (N_10320,N_9208,N_8857);
xor U10321 (N_10321,N_9377,N_8663);
and U10322 (N_10322,N_9423,N_9487);
and U10323 (N_10323,N_9581,N_8568);
xor U10324 (N_10324,N_9169,N_8788);
xnor U10325 (N_10325,N_8464,N_8603);
and U10326 (N_10326,N_9253,N_9569);
xor U10327 (N_10327,N_8515,N_9310);
xnor U10328 (N_10328,N_9577,N_8742);
or U10329 (N_10329,N_9084,N_9146);
and U10330 (N_10330,N_9219,N_9270);
nand U10331 (N_10331,N_8564,N_8592);
nor U10332 (N_10332,N_9418,N_9585);
nand U10333 (N_10333,N_8421,N_9083);
and U10334 (N_10334,N_8843,N_8528);
or U10335 (N_10335,N_8500,N_8902);
and U10336 (N_10336,N_9119,N_8578);
nor U10337 (N_10337,N_9389,N_8873);
or U10338 (N_10338,N_9218,N_8707);
and U10339 (N_10339,N_9228,N_8653);
and U10340 (N_10340,N_9330,N_9399);
and U10341 (N_10341,N_9491,N_8701);
and U10342 (N_10342,N_8815,N_8532);
nor U10343 (N_10343,N_8747,N_9457);
or U10344 (N_10344,N_9438,N_8871);
and U10345 (N_10345,N_8722,N_9099);
or U10346 (N_10346,N_8887,N_8897);
or U10347 (N_10347,N_8679,N_9428);
or U10348 (N_10348,N_8556,N_9368);
nor U10349 (N_10349,N_8948,N_9124);
nand U10350 (N_10350,N_8843,N_9143);
xor U10351 (N_10351,N_8951,N_9334);
nand U10352 (N_10352,N_8419,N_9244);
and U10353 (N_10353,N_9011,N_9299);
xnor U10354 (N_10354,N_9317,N_8437);
xnor U10355 (N_10355,N_9495,N_9027);
and U10356 (N_10356,N_9531,N_8760);
nor U10357 (N_10357,N_8492,N_9421);
nor U10358 (N_10358,N_9353,N_8677);
and U10359 (N_10359,N_9382,N_9032);
xnor U10360 (N_10360,N_9169,N_8947);
nand U10361 (N_10361,N_8525,N_9477);
nand U10362 (N_10362,N_8628,N_9234);
xnor U10363 (N_10363,N_9503,N_9211);
nor U10364 (N_10364,N_8681,N_8609);
xor U10365 (N_10365,N_9557,N_8970);
and U10366 (N_10366,N_9119,N_8614);
xnor U10367 (N_10367,N_9490,N_9454);
and U10368 (N_10368,N_8781,N_8830);
and U10369 (N_10369,N_9447,N_8945);
xor U10370 (N_10370,N_9167,N_8721);
xor U10371 (N_10371,N_8586,N_9225);
or U10372 (N_10372,N_9257,N_9156);
nand U10373 (N_10373,N_8704,N_8531);
nor U10374 (N_10374,N_9212,N_9230);
nor U10375 (N_10375,N_8818,N_8880);
nand U10376 (N_10376,N_9075,N_9312);
and U10377 (N_10377,N_8760,N_8547);
nand U10378 (N_10378,N_9107,N_8643);
and U10379 (N_10379,N_8848,N_9502);
xor U10380 (N_10380,N_8941,N_8441);
or U10381 (N_10381,N_9373,N_9584);
xnor U10382 (N_10382,N_9206,N_9176);
nand U10383 (N_10383,N_9500,N_8482);
and U10384 (N_10384,N_9304,N_9568);
or U10385 (N_10385,N_8856,N_9242);
nand U10386 (N_10386,N_8766,N_9470);
and U10387 (N_10387,N_9361,N_9444);
nor U10388 (N_10388,N_8830,N_9269);
and U10389 (N_10389,N_9442,N_8980);
or U10390 (N_10390,N_8839,N_9420);
nor U10391 (N_10391,N_8648,N_9538);
nand U10392 (N_10392,N_9341,N_8845);
xnor U10393 (N_10393,N_8541,N_9571);
xnor U10394 (N_10394,N_9505,N_9104);
or U10395 (N_10395,N_8910,N_9000);
and U10396 (N_10396,N_8616,N_8484);
or U10397 (N_10397,N_8980,N_8589);
nand U10398 (N_10398,N_9342,N_8783);
or U10399 (N_10399,N_8688,N_8711);
nor U10400 (N_10400,N_9510,N_9283);
nor U10401 (N_10401,N_9599,N_9017);
or U10402 (N_10402,N_9361,N_9035);
nor U10403 (N_10403,N_9572,N_9459);
or U10404 (N_10404,N_8653,N_9090);
nor U10405 (N_10405,N_8545,N_9134);
nor U10406 (N_10406,N_8817,N_9004);
or U10407 (N_10407,N_8537,N_9201);
xnor U10408 (N_10408,N_8442,N_9327);
nor U10409 (N_10409,N_8560,N_9064);
xnor U10410 (N_10410,N_8688,N_8864);
or U10411 (N_10411,N_8653,N_9202);
or U10412 (N_10412,N_9249,N_8657);
or U10413 (N_10413,N_9086,N_9152);
nor U10414 (N_10414,N_8565,N_9521);
and U10415 (N_10415,N_8442,N_9316);
nor U10416 (N_10416,N_9437,N_9470);
or U10417 (N_10417,N_9144,N_8609);
or U10418 (N_10418,N_8961,N_8687);
or U10419 (N_10419,N_8472,N_8837);
xor U10420 (N_10420,N_9470,N_9078);
or U10421 (N_10421,N_8749,N_8847);
nor U10422 (N_10422,N_9407,N_8920);
nand U10423 (N_10423,N_9260,N_9018);
nand U10424 (N_10424,N_9070,N_9098);
nor U10425 (N_10425,N_8722,N_9440);
nor U10426 (N_10426,N_8439,N_9191);
nor U10427 (N_10427,N_9199,N_8811);
nand U10428 (N_10428,N_8665,N_8760);
and U10429 (N_10429,N_8430,N_8510);
nor U10430 (N_10430,N_9235,N_8578);
and U10431 (N_10431,N_9295,N_9304);
nor U10432 (N_10432,N_9148,N_9376);
or U10433 (N_10433,N_9176,N_8789);
and U10434 (N_10434,N_9160,N_8557);
nor U10435 (N_10435,N_8929,N_9566);
or U10436 (N_10436,N_9124,N_9495);
or U10437 (N_10437,N_9323,N_8614);
xnor U10438 (N_10438,N_9343,N_9322);
or U10439 (N_10439,N_9366,N_9428);
and U10440 (N_10440,N_9299,N_9269);
nor U10441 (N_10441,N_8923,N_9105);
or U10442 (N_10442,N_9222,N_9175);
nand U10443 (N_10443,N_9242,N_9191);
or U10444 (N_10444,N_8402,N_9186);
or U10445 (N_10445,N_8591,N_9266);
and U10446 (N_10446,N_9499,N_9134);
nand U10447 (N_10447,N_8768,N_8824);
nand U10448 (N_10448,N_9598,N_8740);
and U10449 (N_10449,N_9325,N_9467);
xnor U10450 (N_10450,N_9242,N_8963);
xor U10451 (N_10451,N_9326,N_8621);
or U10452 (N_10452,N_9199,N_8842);
nor U10453 (N_10453,N_8638,N_9272);
nand U10454 (N_10454,N_8677,N_9061);
and U10455 (N_10455,N_9007,N_8877);
xnor U10456 (N_10456,N_9411,N_8587);
and U10457 (N_10457,N_9521,N_8819);
or U10458 (N_10458,N_8858,N_9327);
nand U10459 (N_10459,N_8649,N_9554);
nor U10460 (N_10460,N_8508,N_9035);
xor U10461 (N_10461,N_9300,N_9513);
nand U10462 (N_10462,N_9563,N_8444);
nand U10463 (N_10463,N_8688,N_8763);
nand U10464 (N_10464,N_8543,N_8893);
nor U10465 (N_10465,N_9058,N_9300);
or U10466 (N_10466,N_9218,N_8417);
nor U10467 (N_10467,N_8450,N_8594);
or U10468 (N_10468,N_8969,N_9122);
nor U10469 (N_10469,N_9488,N_9393);
nor U10470 (N_10470,N_8608,N_8938);
and U10471 (N_10471,N_9006,N_9261);
xnor U10472 (N_10472,N_9109,N_9530);
xor U10473 (N_10473,N_9329,N_8593);
and U10474 (N_10474,N_8928,N_8541);
and U10475 (N_10475,N_8652,N_9269);
and U10476 (N_10476,N_9500,N_9543);
nor U10477 (N_10477,N_9412,N_8483);
and U10478 (N_10478,N_9223,N_8835);
nor U10479 (N_10479,N_9508,N_8532);
or U10480 (N_10480,N_8540,N_8400);
nor U10481 (N_10481,N_8618,N_9226);
xnor U10482 (N_10482,N_8438,N_9261);
nor U10483 (N_10483,N_8503,N_8420);
xnor U10484 (N_10484,N_8858,N_9270);
nor U10485 (N_10485,N_9179,N_8766);
nand U10486 (N_10486,N_9571,N_8933);
nand U10487 (N_10487,N_8879,N_8706);
nand U10488 (N_10488,N_9084,N_9467);
nor U10489 (N_10489,N_9196,N_8993);
nand U10490 (N_10490,N_9133,N_8783);
or U10491 (N_10491,N_8733,N_8676);
and U10492 (N_10492,N_9360,N_8540);
or U10493 (N_10493,N_9255,N_9209);
or U10494 (N_10494,N_8664,N_9167);
nor U10495 (N_10495,N_9171,N_9520);
nor U10496 (N_10496,N_9274,N_8657);
xor U10497 (N_10497,N_9349,N_8698);
nor U10498 (N_10498,N_9292,N_9299);
xor U10499 (N_10499,N_9472,N_9530);
xor U10500 (N_10500,N_8799,N_9375);
and U10501 (N_10501,N_8629,N_9100);
and U10502 (N_10502,N_8469,N_8979);
or U10503 (N_10503,N_8775,N_8444);
nand U10504 (N_10504,N_9178,N_8778);
and U10505 (N_10505,N_8803,N_9020);
nor U10506 (N_10506,N_8530,N_9403);
and U10507 (N_10507,N_9358,N_8720);
and U10508 (N_10508,N_9393,N_8768);
xor U10509 (N_10509,N_8781,N_8702);
xnor U10510 (N_10510,N_8591,N_8427);
or U10511 (N_10511,N_8425,N_8990);
nand U10512 (N_10512,N_9212,N_8689);
nor U10513 (N_10513,N_9421,N_9540);
nand U10514 (N_10514,N_8687,N_8904);
xor U10515 (N_10515,N_8993,N_9122);
and U10516 (N_10516,N_9226,N_9409);
and U10517 (N_10517,N_9397,N_9127);
nand U10518 (N_10518,N_8930,N_8416);
and U10519 (N_10519,N_8782,N_8475);
nor U10520 (N_10520,N_8637,N_9200);
nor U10521 (N_10521,N_9198,N_9438);
nor U10522 (N_10522,N_8517,N_9083);
nor U10523 (N_10523,N_9365,N_8686);
nand U10524 (N_10524,N_8962,N_8516);
or U10525 (N_10525,N_9200,N_9444);
nand U10526 (N_10526,N_8734,N_9156);
or U10527 (N_10527,N_8944,N_9511);
or U10528 (N_10528,N_8978,N_8923);
or U10529 (N_10529,N_8583,N_8759);
nand U10530 (N_10530,N_8801,N_9057);
and U10531 (N_10531,N_8594,N_9410);
nand U10532 (N_10532,N_8813,N_9521);
and U10533 (N_10533,N_9175,N_9419);
and U10534 (N_10534,N_9313,N_9589);
and U10535 (N_10535,N_9403,N_8977);
and U10536 (N_10536,N_9371,N_9080);
nor U10537 (N_10537,N_9101,N_9280);
nand U10538 (N_10538,N_9160,N_9210);
and U10539 (N_10539,N_9243,N_9528);
nor U10540 (N_10540,N_9295,N_8584);
nand U10541 (N_10541,N_8789,N_9508);
nor U10542 (N_10542,N_8931,N_9289);
or U10543 (N_10543,N_8555,N_9442);
nor U10544 (N_10544,N_8506,N_8916);
xor U10545 (N_10545,N_9554,N_8502);
xor U10546 (N_10546,N_8733,N_9020);
xor U10547 (N_10547,N_9198,N_9540);
and U10548 (N_10548,N_9312,N_8416);
or U10549 (N_10549,N_9176,N_8989);
xor U10550 (N_10550,N_9291,N_8526);
xnor U10551 (N_10551,N_9303,N_8537);
nor U10552 (N_10552,N_9364,N_9314);
and U10553 (N_10553,N_8631,N_9174);
nor U10554 (N_10554,N_9544,N_9379);
and U10555 (N_10555,N_9565,N_9547);
nand U10556 (N_10556,N_9212,N_8567);
nand U10557 (N_10557,N_9545,N_9230);
xor U10558 (N_10558,N_9551,N_8737);
or U10559 (N_10559,N_8421,N_9558);
nand U10560 (N_10560,N_8548,N_8709);
nand U10561 (N_10561,N_8548,N_8599);
and U10562 (N_10562,N_9384,N_9511);
nand U10563 (N_10563,N_9252,N_8459);
nand U10564 (N_10564,N_8784,N_8880);
xor U10565 (N_10565,N_8492,N_9247);
xor U10566 (N_10566,N_8441,N_8929);
nand U10567 (N_10567,N_9189,N_8689);
or U10568 (N_10568,N_8887,N_9081);
and U10569 (N_10569,N_9285,N_9310);
xor U10570 (N_10570,N_8962,N_9220);
or U10571 (N_10571,N_8758,N_8964);
nor U10572 (N_10572,N_8673,N_8987);
or U10573 (N_10573,N_9030,N_8470);
and U10574 (N_10574,N_9540,N_9283);
or U10575 (N_10575,N_9005,N_8581);
or U10576 (N_10576,N_9106,N_8842);
nand U10577 (N_10577,N_9373,N_8421);
and U10578 (N_10578,N_9255,N_9422);
nand U10579 (N_10579,N_8894,N_9433);
or U10580 (N_10580,N_8403,N_8965);
xnor U10581 (N_10581,N_8642,N_8440);
nor U10582 (N_10582,N_8495,N_8416);
and U10583 (N_10583,N_8912,N_8827);
nand U10584 (N_10584,N_9138,N_8639);
xor U10585 (N_10585,N_9556,N_8475);
xor U10586 (N_10586,N_8553,N_9038);
or U10587 (N_10587,N_9450,N_9063);
nor U10588 (N_10588,N_9557,N_9166);
nor U10589 (N_10589,N_9485,N_8443);
xor U10590 (N_10590,N_9400,N_9554);
and U10591 (N_10591,N_9051,N_8997);
and U10592 (N_10592,N_8448,N_8419);
or U10593 (N_10593,N_9280,N_8824);
nor U10594 (N_10594,N_8951,N_9557);
or U10595 (N_10595,N_8692,N_9012);
or U10596 (N_10596,N_8631,N_8640);
nor U10597 (N_10597,N_8555,N_8981);
xor U10598 (N_10598,N_8751,N_9046);
xnor U10599 (N_10599,N_9361,N_9592);
xor U10600 (N_10600,N_9225,N_9204);
and U10601 (N_10601,N_9470,N_9375);
or U10602 (N_10602,N_8470,N_9094);
and U10603 (N_10603,N_8957,N_8650);
xnor U10604 (N_10604,N_8833,N_9065);
and U10605 (N_10605,N_8981,N_8816);
nor U10606 (N_10606,N_8458,N_8683);
or U10607 (N_10607,N_9262,N_8718);
and U10608 (N_10608,N_9220,N_9583);
and U10609 (N_10609,N_8931,N_8534);
nor U10610 (N_10610,N_8739,N_9147);
or U10611 (N_10611,N_8787,N_9094);
nor U10612 (N_10612,N_8631,N_9277);
nand U10613 (N_10613,N_9102,N_9003);
and U10614 (N_10614,N_9359,N_9444);
xnor U10615 (N_10615,N_8946,N_9365);
xnor U10616 (N_10616,N_9426,N_9005);
or U10617 (N_10617,N_8538,N_9299);
and U10618 (N_10618,N_9154,N_9512);
or U10619 (N_10619,N_9280,N_9193);
nor U10620 (N_10620,N_8805,N_9505);
or U10621 (N_10621,N_9223,N_9553);
or U10622 (N_10622,N_9287,N_9300);
and U10623 (N_10623,N_8705,N_8429);
or U10624 (N_10624,N_9085,N_9290);
nor U10625 (N_10625,N_9585,N_9455);
nor U10626 (N_10626,N_9169,N_8765);
xor U10627 (N_10627,N_8440,N_9206);
and U10628 (N_10628,N_9006,N_9014);
xor U10629 (N_10629,N_8409,N_9001);
xor U10630 (N_10630,N_8542,N_9320);
xnor U10631 (N_10631,N_9001,N_9298);
nand U10632 (N_10632,N_8418,N_9031);
and U10633 (N_10633,N_9458,N_8705);
xor U10634 (N_10634,N_8426,N_9532);
or U10635 (N_10635,N_9169,N_8634);
xor U10636 (N_10636,N_9598,N_8954);
nor U10637 (N_10637,N_8597,N_9223);
and U10638 (N_10638,N_8883,N_8527);
and U10639 (N_10639,N_8602,N_8448);
xor U10640 (N_10640,N_8779,N_9587);
xor U10641 (N_10641,N_9305,N_8968);
nor U10642 (N_10642,N_9499,N_8431);
nand U10643 (N_10643,N_9195,N_9429);
or U10644 (N_10644,N_9101,N_9257);
xnor U10645 (N_10645,N_8931,N_9173);
nand U10646 (N_10646,N_9214,N_9231);
nor U10647 (N_10647,N_8989,N_9454);
or U10648 (N_10648,N_9124,N_9369);
or U10649 (N_10649,N_9441,N_8856);
or U10650 (N_10650,N_9506,N_8475);
nand U10651 (N_10651,N_9544,N_9390);
or U10652 (N_10652,N_9078,N_9145);
nand U10653 (N_10653,N_8506,N_9011);
nor U10654 (N_10654,N_9004,N_8931);
nor U10655 (N_10655,N_9144,N_9007);
or U10656 (N_10656,N_8993,N_9404);
or U10657 (N_10657,N_9351,N_9020);
nand U10658 (N_10658,N_8907,N_9509);
xor U10659 (N_10659,N_8719,N_8710);
xor U10660 (N_10660,N_8590,N_8518);
nor U10661 (N_10661,N_9519,N_8861);
nand U10662 (N_10662,N_9471,N_8678);
or U10663 (N_10663,N_8820,N_8782);
and U10664 (N_10664,N_9062,N_9142);
nand U10665 (N_10665,N_9537,N_9071);
xor U10666 (N_10666,N_9423,N_8752);
nand U10667 (N_10667,N_9000,N_9275);
nand U10668 (N_10668,N_9371,N_9305);
xnor U10669 (N_10669,N_9073,N_8983);
xnor U10670 (N_10670,N_8496,N_9045);
nor U10671 (N_10671,N_9092,N_9369);
or U10672 (N_10672,N_8625,N_8776);
and U10673 (N_10673,N_8553,N_8878);
nor U10674 (N_10674,N_9536,N_8956);
or U10675 (N_10675,N_8660,N_9175);
and U10676 (N_10676,N_8823,N_9015);
nand U10677 (N_10677,N_9489,N_8904);
nor U10678 (N_10678,N_9189,N_8727);
nor U10679 (N_10679,N_9406,N_8518);
xor U10680 (N_10680,N_8889,N_9428);
or U10681 (N_10681,N_8652,N_9404);
nand U10682 (N_10682,N_8802,N_9031);
xor U10683 (N_10683,N_9114,N_9180);
nor U10684 (N_10684,N_8867,N_9301);
xor U10685 (N_10685,N_8737,N_8790);
or U10686 (N_10686,N_8843,N_9111);
and U10687 (N_10687,N_8699,N_8791);
nand U10688 (N_10688,N_9183,N_9048);
nor U10689 (N_10689,N_9306,N_9194);
nor U10690 (N_10690,N_8837,N_9017);
nor U10691 (N_10691,N_9210,N_8407);
or U10692 (N_10692,N_8786,N_8545);
or U10693 (N_10693,N_8734,N_8603);
nand U10694 (N_10694,N_8783,N_8557);
nor U10695 (N_10695,N_8758,N_9027);
and U10696 (N_10696,N_8739,N_9132);
or U10697 (N_10697,N_8867,N_8568);
nor U10698 (N_10698,N_9177,N_9571);
xor U10699 (N_10699,N_8481,N_8543);
nand U10700 (N_10700,N_9532,N_8469);
or U10701 (N_10701,N_8670,N_9567);
and U10702 (N_10702,N_8437,N_8433);
or U10703 (N_10703,N_8970,N_9214);
nor U10704 (N_10704,N_8808,N_9305);
or U10705 (N_10705,N_8962,N_8494);
nand U10706 (N_10706,N_8830,N_8978);
and U10707 (N_10707,N_8740,N_8975);
or U10708 (N_10708,N_8875,N_9009);
xnor U10709 (N_10709,N_9167,N_9564);
nand U10710 (N_10710,N_8764,N_9437);
and U10711 (N_10711,N_8931,N_9141);
and U10712 (N_10712,N_8660,N_8902);
xnor U10713 (N_10713,N_9558,N_9014);
nand U10714 (N_10714,N_9035,N_8646);
and U10715 (N_10715,N_8442,N_8860);
nor U10716 (N_10716,N_8603,N_9228);
nand U10717 (N_10717,N_9169,N_9454);
or U10718 (N_10718,N_8535,N_8767);
xor U10719 (N_10719,N_9549,N_9169);
nand U10720 (N_10720,N_9501,N_8502);
nand U10721 (N_10721,N_9516,N_9411);
nor U10722 (N_10722,N_9400,N_9263);
nand U10723 (N_10723,N_8578,N_9027);
xnor U10724 (N_10724,N_8451,N_9134);
xor U10725 (N_10725,N_9092,N_8530);
xnor U10726 (N_10726,N_9193,N_9576);
and U10727 (N_10727,N_9107,N_8998);
or U10728 (N_10728,N_8598,N_9526);
xnor U10729 (N_10729,N_9071,N_8722);
or U10730 (N_10730,N_8430,N_9592);
xor U10731 (N_10731,N_8674,N_9394);
nor U10732 (N_10732,N_9301,N_8876);
nand U10733 (N_10733,N_9257,N_8418);
nor U10734 (N_10734,N_8607,N_8646);
nand U10735 (N_10735,N_9091,N_9575);
xnor U10736 (N_10736,N_9324,N_8843);
and U10737 (N_10737,N_8808,N_9508);
nand U10738 (N_10738,N_9415,N_8670);
and U10739 (N_10739,N_8438,N_8845);
xnor U10740 (N_10740,N_8841,N_9373);
or U10741 (N_10741,N_8455,N_8652);
nand U10742 (N_10742,N_9149,N_8554);
nor U10743 (N_10743,N_9370,N_9417);
or U10744 (N_10744,N_9109,N_9265);
or U10745 (N_10745,N_8605,N_9340);
or U10746 (N_10746,N_9064,N_8893);
xnor U10747 (N_10747,N_8980,N_9194);
or U10748 (N_10748,N_9586,N_9363);
xor U10749 (N_10749,N_9358,N_9369);
xnor U10750 (N_10750,N_8969,N_9092);
nor U10751 (N_10751,N_9162,N_9172);
nor U10752 (N_10752,N_8740,N_9469);
nand U10753 (N_10753,N_8574,N_8515);
nand U10754 (N_10754,N_9107,N_9440);
nand U10755 (N_10755,N_9246,N_9094);
and U10756 (N_10756,N_9301,N_9520);
xnor U10757 (N_10757,N_8631,N_9057);
xor U10758 (N_10758,N_9200,N_8618);
xor U10759 (N_10759,N_9506,N_9237);
nor U10760 (N_10760,N_9175,N_9093);
and U10761 (N_10761,N_8884,N_8782);
and U10762 (N_10762,N_9522,N_8574);
nand U10763 (N_10763,N_9338,N_9543);
nand U10764 (N_10764,N_9153,N_8721);
and U10765 (N_10765,N_8749,N_9502);
xor U10766 (N_10766,N_8666,N_8814);
and U10767 (N_10767,N_9214,N_8937);
or U10768 (N_10768,N_8624,N_9377);
nand U10769 (N_10769,N_9125,N_9006);
or U10770 (N_10770,N_8737,N_8565);
nor U10771 (N_10771,N_8450,N_9289);
xor U10772 (N_10772,N_9293,N_8482);
nor U10773 (N_10773,N_8782,N_9081);
nor U10774 (N_10774,N_9058,N_8722);
xor U10775 (N_10775,N_9050,N_8799);
nand U10776 (N_10776,N_8476,N_8913);
xor U10777 (N_10777,N_9399,N_8439);
and U10778 (N_10778,N_8506,N_9373);
nor U10779 (N_10779,N_8738,N_8509);
or U10780 (N_10780,N_9449,N_8503);
nand U10781 (N_10781,N_9346,N_8644);
xor U10782 (N_10782,N_8643,N_9064);
or U10783 (N_10783,N_9488,N_8941);
nor U10784 (N_10784,N_9081,N_8794);
nand U10785 (N_10785,N_9339,N_9446);
or U10786 (N_10786,N_8858,N_9271);
and U10787 (N_10787,N_8837,N_9098);
or U10788 (N_10788,N_9163,N_8533);
or U10789 (N_10789,N_9261,N_9579);
and U10790 (N_10790,N_9236,N_8683);
or U10791 (N_10791,N_8442,N_8956);
or U10792 (N_10792,N_9073,N_8538);
nor U10793 (N_10793,N_9525,N_9329);
xor U10794 (N_10794,N_9599,N_9331);
nand U10795 (N_10795,N_9107,N_9480);
and U10796 (N_10796,N_8835,N_8779);
or U10797 (N_10797,N_8490,N_9156);
or U10798 (N_10798,N_9529,N_8443);
nand U10799 (N_10799,N_9004,N_8895);
xnor U10800 (N_10800,N_9718,N_9788);
or U10801 (N_10801,N_9863,N_10498);
or U10802 (N_10802,N_10719,N_9763);
and U10803 (N_10803,N_9710,N_10112);
or U10804 (N_10804,N_9951,N_9671);
nand U10805 (N_10805,N_10680,N_10072);
xor U10806 (N_10806,N_10753,N_10426);
nor U10807 (N_10807,N_9885,N_10672);
or U10808 (N_10808,N_10595,N_9682);
nor U10809 (N_10809,N_9850,N_10623);
xor U10810 (N_10810,N_10665,N_10195);
xor U10811 (N_10811,N_10659,N_9734);
or U10812 (N_10812,N_10250,N_9781);
nor U10813 (N_10813,N_9976,N_10727);
or U10814 (N_10814,N_10502,N_10705);
nand U10815 (N_10815,N_10227,N_10641);
nor U10816 (N_10816,N_10429,N_10054);
or U10817 (N_10817,N_9967,N_10164);
nor U10818 (N_10818,N_10414,N_9805);
and U10819 (N_10819,N_9617,N_10696);
nor U10820 (N_10820,N_9676,N_10673);
and U10821 (N_10821,N_10579,N_9873);
nand U10822 (N_10822,N_10224,N_9772);
or U10823 (N_10823,N_10202,N_10386);
nand U10824 (N_10824,N_10435,N_10326);
or U10825 (N_10825,N_9990,N_9766);
nor U10826 (N_10826,N_9757,N_10678);
xor U10827 (N_10827,N_9620,N_9644);
and U10828 (N_10828,N_10441,N_10522);
or U10829 (N_10829,N_9880,N_10583);
nand U10830 (N_10830,N_10045,N_10071);
xnor U10831 (N_10831,N_10307,N_9623);
or U10832 (N_10832,N_9736,N_10430);
nor U10833 (N_10833,N_9814,N_10764);
xnor U10834 (N_10834,N_10364,N_10629);
nor U10835 (N_10835,N_10682,N_10464);
and U10836 (N_10836,N_10327,N_9981);
nand U10837 (N_10837,N_10702,N_9871);
or U10838 (N_10838,N_10133,N_10110);
and U10839 (N_10839,N_10411,N_9603);
nand U10840 (N_10840,N_10617,N_10466);
and U10841 (N_10841,N_10317,N_10138);
xor U10842 (N_10842,N_10253,N_10225);
nand U10843 (N_10843,N_10457,N_10275);
nand U10844 (N_10844,N_10300,N_10029);
or U10845 (N_10845,N_10402,N_10670);
xor U10846 (N_10846,N_10733,N_10676);
xor U10847 (N_10847,N_10143,N_9777);
and U10848 (N_10848,N_10574,N_10365);
and U10849 (N_10849,N_10248,N_10350);
nor U10850 (N_10850,N_10585,N_10362);
and U10851 (N_10851,N_10545,N_10217);
or U10852 (N_10852,N_10157,N_9765);
nor U10853 (N_10853,N_9614,N_10262);
nand U10854 (N_10854,N_10016,N_9975);
xor U10855 (N_10855,N_10700,N_10575);
or U10856 (N_10856,N_10127,N_10101);
or U10857 (N_10857,N_10632,N_10795);
nor U10858 (N_10858,N_10507,N_10000);
and U10859 (N_10859,N_10452,N_10625);
xor U10860 (N_10860,N_10398,N_10343);
or U10861 (N_10861,N_9669,N_10436);
xor U10862 (N_10862,N_10748,N_10494);
nand U10863 (N_10863,N_10311,N_9997);
or U10864 (N_10864,N_9960,N_10400);
xor U10865 (N_10865,N_9843,N_10111);
and U10866 (N_10866,N_9600,N_10059);
and U10867 (N_10867,N_9618,N_10689);
xor U10868 (N_10868,N_10216,N_10460);
or U10869 (N_10869,N_9635,N_9690);
nor U10870 (N_10870,N_10653,N_9657);
xor U10871 (N_10871,N_9927,N_10105);
or U10872 (N_10872,N_10654,N_10104);
nand U10873 (N_10873,N_9881,N_10396);
nor U10874 (N_10874,N_10776,N_9625);
nor U10875 (N_10875,N_9877,N_9965);
or U10876 (N_10876,N_9692,N_9764);
or U10877 (N_10877,N_10528,N_10085);
and U10878 (N_10878,N_10598,N_10269);
nor U10879 (N_10879,N_10624,N_10099);
and U10880 (N_10880,N_10368,N_10090);
nand U10881 (N_10881,N_9649,N_9861);
or U10882 (N_10882,N_10352,N_9667);
xnor U10883 (N_10883,N_10268,N_10289);
or U10884 (N_10884,N_9898,N_10273);
nor U10885 (N_10885,N_9956,N_9744);
nor U10886 (N_10886,N_10550,N_9979);
xnor U10887 (N_10887,N_10564,N_10660);
or U10888 (N_10888,N_10531,N_10572);
xor U10889 (N_10889,N_9913,N_9659);
nor U10890 (N_10890,N_10231,N_9767);
and U10891 (N_10891,N_10658,N_10760);
or U10892 (N_10892,N_9878,N_9826);
nand U10893 (N_10893,N_10001,N_10146);
xor U10894 (N_10894,N_9911,N_9604);
and U10895 (N_10895,N_9780,N_10605);
xnor U10896 (N_10896,N_10485,N_10197);
nand U10897 (N_10897,N_10006,N_9857);
or U10898 (N_10898,N_9899,N_10515);
nor U10899 (N_10899,N_10043,N_10314);
nand U10900 (N_10900,N_10361,N_10095);
nand U10901 (N_10901,N_9910,N_10416);
nand U10902 (N_10902,N_9816,N_10431);
nor U10903 (N_10903,N_10780,N_10304);
nor U10904 (N_10904,N_9973,N_9828);
and U10905 (N_10905,N_10504,N_10232);
or U10906 (N_10906,N_9714,N_10186);
nor U10907 (N_10907,N_10103,N_10423);
xor U10908 (N_10908,N_9868,N_10633);
or U10909 (N_10909,N_10322,N_10235);
nand U10910 (N_10910,N_9661,N_10473);
nand U10911 (N_10911,N_9648,N_10066);
nand U10912 (N_10912,N_10568,N_9702);
and U10913 (N_10913,N_10712,N_10287);
and U10914 (N_10914,N_10525,N_9611);
and U10915 (N_10915,N_10159,N_10567);
nand U10916 (N_10916,N_10387,N_10695);
nand U10917 (N_10917,N_9647,N_9619);
and U10918 (N_10918,N_10184,N_10474);
nand U10919 (N_10919,N_10087,N_10338);
and U10920 (N_10920,N_10758,N_10272);
and U10921 (N_10921,N_9935,N_9622);
nand U10922 (N_10922,N_9853,N_10663);
and U10923 (N_10923,N_10736,N_10381);
nand U10924 (N_10924,N_10382,N_9691);
and U10925 (N_10925,N_9632,N_9807);
xor U10926 (N_10926,N_10088,N_10173);
xor U10927 (N_10927,N_10497,N_10377);
xor U10928 (N_10928,N_10607,N_9773);
nor U10929 (N_10929,N_10266,N_10487);
nand U10930 (N_10930,N_9808,N_10440);
xnor U10931 (N_10931,N_10076,N_9964);
nor U10932 (N_10932,N_10739,N_9957);
nand U10933 (N_10933,N_9995,N_9797);
xor U10934 (N_10934,N_9723,N_9866);
xnor U10935 (N_10935,N_10005,N_9892);
nand U10936 (N_10936,N_10170,N_10533);
nand U10937 (N_10937,N_10615,N_9947);
nor U10938 (N_10938,N_10578,N_10379);
nand U10939 (N_10939,N_10380,N_10121);
xnor U10940 (N_10940,N_10732,N_9638);
nand U10941 (N_10941,N_10551,N_10245);
xor U10942 (N_10942,N_10030,N_10233);
or U10943 (N_10943,N_10465,N_10628);
and U10944 (N_10944,N_9709,N_10768);
and U10945 (N_10945,N_10378,N_10210);
or U10946 (N_10946,N_10002,N_10067);
and U10947 (N_10947,N_10675,N_10264);
nor U10948 (N_10948,N_9776,N_9607);
and U10949 (N_10949,N_10506,N_9890);
nand U10950 (N_10950,N_10277,N_10614);
or U10951 (N_10951,N_10293,N_9694);
nor U10952 (N_10952,N_9705,N_10310);
xor U10953 (N_10953,N_9738,N_10544);
xor U10954 (N_10954,N_10394,N_9670);
and U10955 (N_10955,N_10309,N_10081);
nor U10956 (N_10956,N_10455,N_9700);
and U10957 (N_10957,N_10655,N_10461);
xor U10958 (N_10958,N_9803,N_10511);
nand U10959 (N_10959,N_10267,N_10150);
nand U10960 (N_10960,N_10622,N_10783);
nand U10961 (N_10961,N_10192,N_10097);
or U10962 (N_10962,N_9674,N_10529);
nor U10963 (N_10963,N_9985,N_10291);
or U10964 (N_10964,N_10599,N_10033);
nor U10965 (N_10965,N_9720,N_10540);
or U10966 (N_10966,N_10745,N_10351);
and U10967 (N_10967,N_9724,N_10573);
nor U10968 (N_10968,N_10722,N_10244);
and U10969 (N_10969,N_10409,N_10031);
or U10970 (N_10970,N_9701,N_9818);
xor U10971 (N_10971,N_9977,N_10306);
or U10972 (N_10972,N_9609,N_10360);
nor U10973 (N_10973,N_10332,N_10189);
or U10974 (N_10974,N_10340,N_10297);
nor U10975 (N_10975,N_10483,N_9988);
nor U10976 (N_10976,N_9769,N_10501);
nand U10977 (N_10977,N_9746,N_9745);
nor U10978 (N_10978,N_10613,N_10039);
xor U10979 (N_10979,N_10369,N_10594);
nand U10980 (N_10980,N_10218,N_10239);
nand U10981 (N_10981,N_10693,N_10299);
nor U10982 (N_10982,N_9945,N_9655);
or U10983 (N_10983,N_10543,N_9693);
and U10984 (N_10984,N_10444,N_10735);
or U10985 (N_10985,N_10301,N_10767);
or U10986 (N_10986,N_10683,N_10620);
nand U10987 (N_10987,N_10731,N_10513);
or U10988 (N_10988,N_10296,N_10056);
nand U10989 (N_10989,N_10089,N_10674);
and U10990 (N_10990,N_10290,N_10754);
and U10991 (N_10991,N_10516,N_10499);
xor U10992 (N_10992,N_10201,N_9834);
xor U10993 (N_10993,N_10661,N_10728);
nor U10994 (N_10994,N_9731,N_10724);
and U10995 (N_10995,N_10182,N_10149);
or U10996 (N_10996,N_10552,N_10404);
nand U10997 (N_10997,N_10451,N_9798);
nand U10998 (N_10998,N_9641,N_10458);
xnor U10999 (N_10999,N_9912,N_10281);
or U11000 (N_11000,N_9616,N_10366);
or U11001 (N_11001,N_10008,N_10491);
nand U11002 (N_11002,N_10757,N_9712);
or U11003 (N_11003,N_9770,N_9882);
or U11004 (N_11004,N_9804,N_9634);
xnor U11005 (N_11005,N_10781,N_10004);
or U11006 (N_11006,N_10706,N_10374);
nand U11007 (N_11007,N_10007,N_10510);
and U11008 (N_11008,N_10563,N_9636);
or U11009 (N_11009,N_10288,N_9858);
nor U11010 (N_11010,N_9897,N_10222);
or U11011 (N_11011,N_9784,N_10590);
xor U11012 (N_11012,N_9932,N_9775);
and U11013 (N_11013,N_10162,N_9683);
xnor U11014 (N_11014,N_9688,N_10075);
xor U11015 (N_11015,N_10256,N_10226);
nor U11016 (N_11016,N_10064,N_9822);
and U11017 (N_11017,N_9789,N_10151);
xor U11018 (N_11018,N_9991,N_10018);
or U11019 (N_11019,N_10597,N_10778);
nor U11020 (N_11020,N_9778,N_9753);
or U11021 (N_11021,N_9922,N_10406);
and U11022 (N_11022,N_9728,N_9840);
or U11023 (N_11023,N_10734,N_10260);
or U11024 (N_11024,N_9656,N_10331);
or U11025 (N_11025,N_10080,N_9963);
or U11026 (N_11026,N_10453,N_10241);
or U11027 (N_11027,N_9729,N_10013);
or U11028 (N_11028,N_10477,N_10315);
nor U11029 (N_11029,N_9953,N_9865);
nand U11030 (N_11030,N_9717,N_9917);
or U11031 (N_11031,N_10098,N_10108);
nor U11032 (N_11032,N_10221,N_10247);
and U11033 (N_11033,N_10492,N_10041);
or U11034 (N_11034,N_10084,N_9968);
and U11035 (N_11035,N_9887,N_10236);
nand U11036 (N_11036,N_9665,N_10353);
xnor U11037 (N_11037,N_9695,N_10621);
and U11038 (N_11038,N_10687,N_10619);
nor U11039 (N_11039,N_10468,N_9790);
xor U11040 (N_11040,N_10725,N_10091);
nor U11041 (N_11041,N_10242,N_10634);
nand U11042 (N_11042,N_9761,N_10166);
xor U11043 (N_11043,N_10630,N_9698);
or U11044 (N_11044,N_10637,N_10626);
and U11045 (N_11045,N_9755,N_10037);
nand U11046 (N_11046,N_10541,N_10219);
xnor U11047 (N_11047,N_9906,N_10488);
nor U11048 (N_11048,N_10782,N_9848);
nand U11049 (N_11049,N_10539,N_10475);
xor U11050 (N_11050,N_10535,N_9859);
nand U11051 (N_11051,N_10167,N_10616);
nand U11052 (N_11052,N_9852,N_9844);
and U11053 (N_11053,N_10180,N_9602);
or U11054 (N_11054,N_10114,N_10526);
and U11055 (N_11055,N_10282,N_10639);
and U11056 (N_11056,N_10022,N_9923);
nor U11057 (N_11057,N_9779,N_10342);
nand U11058 (N_11058,N_10669,N_9664);
and U11059 (N_11059,N_9948,N_9854);
and U11060 (N_11060,N_10171,N_9792);
xor U11061 (N_11061,N_9606,N_10120);
and U11062 (N_11062,N_10668,N_10140);
or U11063 (N_11063,N_10390,N_10463);
nor U11064 (N_11064,N_10715,N_10237);
nor U11065 (N_11065,N_9837,N_10212);
xnor U11066 (N_11066,N_10798,N_10196);
nor U11067 (N_11067,N_10303,N_10527);
nor U11068 (N_11068,N_9942,N_9969);
and U11069 (N_11069,N_10771,N_10716);
xnor U11070 (N_11070,N_10355,N_9743);
or U11071 (N_11071,N_9752,N_10015);
xnor U11072 (N_11072,N_10147,N_9972);
nand U11073 (N_11073,N_9938,N_10420);
nor U11074 (N_11074,N_10769,N_10422);
xnor U11075 (N_11075,N_10337,N_9884);
and U11076 (N_11076,N_9802,N_10557);
xnor U11077 (N_11077,N_9987,N_10376);
xnor U11078 (N_11078,N_10721,N_9943);
or U11079 (N_11079,N_10765,N_10358);
and U11080 (N_11080,N_10762,N_10752);
xnor U11081 (N_11081,N_10666,N_9810);
or U11082 (N_11082,N_10417,N_10163);
or U11083 (N_11083,N_10142,N_9914);
and U11084 (N_11084,N_10009,N_10671);
and U11085 (N_11085,N_10647,N_10657);
nor U11086 (N_11086,N_10229,N_10257);
or U11087 (N_11087,N_10538,N_10508);
or U11088 (N_11088,N_10562,N_9982);
nand U11089 (N_11089,N_10011,N_9799);
nor U11090 (N_11090,N_10593,N_9716);
nand U11091 (N_11091,N_10553,N_9952);
and U11092 (N_11092,N_10383,N_10692);
xnor U11093 (N_11093,N_9894,N_9931);
nor U11094 (N_11094,N_10354,N_10472);
or U11095 (N_11095,N_10230,N_10796);
xnor U11096 (N_11096,N_9707,N_9685);
nand U11097 (N_11097,N_9833,N_10571);
and U11098 (N_11098,N_10471,N_9615);
or U11099 (N_11099,N_10141,N_10608);
xnor U11100 (N_11100,N_10428,N_9787);
nor U11101 (N_11101,N_10481,N_10308);
nor U11102 (N_11102,N_10500,N_10793);
nor U11103 (N_11103,N_10106,N_10737);
or U11104 (N_11104,N_10549,N_10651);
and U11105 (N_11105,N_10012,N_10691);
xnor U11106 (N_11106,N_9986,N_9944);
nand U11107 (N_11107,N_10055,N_10160);
or U11108 (N_11108,N_10349,N_10125);
nor U11109 (N_11109,N_9681,N_10292);
xnor U11110 (N_11110,N_10334,N_10199);
nand U11111 (N_11111,N_10512,N_9992);
or U11112 (N_11112,N_10375,N_10493);
nor U11113 (N_11113,N_9936,N_9642);
xnor U11114 (N_11114,N_10486,N_10434);
or U11115 (N_11115,N_9653,N_10274);
nand U11116 (N_11116,N_9930,N_10456);
or U11117 (N_11117,N_10627,N_10328);
and U11118 (N_11118,N_10174,N_10777);
nor U11119 (N_11119,N_10278,N_10602);
or U11120 (N_11120,N_10690,N_10600);
nor U11121 (N_11121,N_10449,N_10710);
or U11122 (N_11122,N_10794,N_9827);
or U11123 (N_11123,N_9876,N_9962);
nor U11124 (N_11124,N_10580,N_10547);
nand U11125 (N_11125,N_9680,N_10482);
or U11126 (N_11126,N_10205,N_10412);
or U11127 (N_11127,N_9631,N_10118);
and U11128 (N_11128,N_10280,N_10726);
nor U11129 (N_11129,N_10642,N_10178);
and U11130 (N_11130,N_10069,N_10587);
or U11131 (N_11131,N_10356,N_10079);
nor U11132 (N_11132,N_10606,N_10129);
nor U11133 (N_11133,N_10418,N_10645);
xor U11134 (N_11134,N_9796,N_9687);
or U11135 (N_11135,N_10145,N_10206);
nand U11136 (N_11136,N_9901,N_9869);
and U11137 (N_11137,N_10773,N_9786);
or U11138 (N_11138,N_10094,N_10389);
nand U11139 (N_11139,N_9675,N_10130);
xor U11140 (N_11140,N_9737,N_9758);
or U11141 (N_11141,N_9946,N_10419);
nor U11142 (N_11142,N_10704,N_10759);
nor U11143 (N_11143,N_10261,N_10359);
nor U11144 (N_11144,N_9934,N_10523);
nor U11145 (N_11145,N_10329,N_10569);
xnor U11146 (N_11146,N_9862,N_10113);
xnor U11147 (N_11147,N_10312,N_10116);
and U11148 (N_11148,N_9624,N_10612);
nand U11149 (N_11149,N_10667,N_9940);
xnor U11150 (N_11150,N_10115,N_10347);
nand U11151 (N_11151,N_9686,N_10559);
xnor U11152 (N_11152,N_10664,N_10316);
nor U11153 (N_11153,N_9704,N_9905);
nor U11154 (N_11154,N_9909,N_10078);
nor U11155 (N_11155,N_10333,N_10791);
or U11156 (N_11156,N_9708,N_9996);
and U11157 (N_11157,N_9955,N_10799);
and U11158 (N_11158,N_10723,N_9732);
or U11159 (N_11159,N_10747,N_9874);
or U11160 (N_11160,N_10408,N_10074);
nand U11161 (N_11161,N_10638,N_9903);
and U11162 (N_11162,N_10405,N_9628);
xor U11163 (N_11163,N_10447,N_10176);
nor U11164 (N_11164,N_10484,N_9949);
nor U11165 (N_11165,N_10028,N_10478);
or U11166 (N_11166,N_10213,N_10720);
nand U11167 (N_11167,N_9791,N_10470);
and U11168 (N_11168,N_9841,N_10751);
and U11169 (N_11169,N_9612,N_10276);
nand U11170 (N_11170,N_10109,N_10397);
or U11171 (N_11171,N_10586,N_9958);
nor U11172 (N_11172,N_10271,N_9812);
or U11173 (N_11173,N_10254,N_10685);
nand U11174 (N_11174,N_9815,N_10220);
xnor U11175 (N_11175,N_10577,N_9795);
xnor U11176 (N_11176,N_9888,N_9879);
nand U11177 (N_11177,N_10610,N_10467);
or U11178 (N_11178,N_10057,N_9809);
or U11179 (N_11179,N_10524,N_10686);
xnor U11180 (N_11180,N_10652,N_10609);
or U11181 (N_11181,N_10161,N_10644);
xor U11182 (N_11182,N_10454,N_10746);
xor U11183 (N_11183,N_9999,N_9684);
nand U11184 (N_11184,N_9771,N_10177);
xnor U11185 (N_11185,N_10373,N_9856);
or U11186 (N_11186,N_10785,N_10701);
nor U11187 (N_11187,N_10503,N_10787);
or U11188 (N_11188,N_10490,N_9851);
xnor U11189 (N_11189,N_9915,N_10036);
or U11190 (N_11190,N_10792,N_9974);
or U11191 (N_11191,N_9715,N_10656);
or U11192 (N_11192,N_10246,N_10040);
or U11193 (N_11193,N_10677,N_10252);
nor U11194 (N_11194,N_9739,N_10155);
nor U11195 (N_11195,N_10279,N_10789);
and U11196 (N_11196,N_9760,N_9836);
and U11197 (N_11197,N_10203,N_9835);
and U11198 (N_11198,N_10168,N_10576);
or U11199 (N_11199,N_10480,N_9768);
and U11200 (N_11200,N_9697,N_10020);
nand U11201 (N_11201,N_10711,N_10320);
xnor U11202 (N_11202,N_9993,N_10175);
nand U11203 (N_11203,N_9646,N_10603);
nor U11204 (N_11204,N_9933,N_10019);
nand U11205 (N_11205,N_9782,N_10392);
or U11206 (N_11206,N_9762,N_10183);
nor U11207 (N_11207,N_9756,N_10514);
or U11208 (N_11208,N_10432,N_10729);
and U11209 (N_11209,N_9678,N_9846);
nor U11210 (N_11210,N_9630,N_9754);
nor U11211 (N_11211,N_10058,N_10215);
nand U11212 (N_11212,N_10565,N_10649);
and U11213 (N_11213,N_10152,N_10052);
nand U11214 (N_11214,N_9733,N_10640);
nand U11215 (N_11215,N_9983,N_10462);
and U11216 (N_11216,N_9713,N_9939);
xnor U11217 (N_11217,N_10694,N_9699);
nor U11218 (N_11218,N_9929,N_9817);
nand U11219 (N_11219,N_10413,N_10295);
xor U11220 (N_11220,N_10024,N_10259);
nor U11221 (N_11221,N_10169,N_10385);
or U11222 (N_11222,N_10062,N_10198);
xor U11223 (N_11223,N_10443,N_9847);
xnor U11224 (N_11224,N_10536,N_10144);
xor U11225 (N_11225,N_9830,N_10285);
or U11226 (N_11226,N_9902,N_10393);
xor U11227 (N_11227,N_9954,N_10083);
or U11228 (N_11228,N_9845,N_9742);
nor U11229 (N_11229,N_10153,N_10438);
or U11230 (N_11230,N_10318,N_9672);
or U11231 (N_11231,N_10073,N_10284);
nor U11232 (N_11232,N_9959,N_10372);
and U11233 (N_11233,N_10530,N_10707);
and U11234 (N_11234,N_10193,N_10046);
or U11235 (N_11235,N_10243,N_9730);
nor U11236 (N_11236,N_10755,N_10065);
or U11237 (N_11237,N_10698,N_9785);
nor U11238 (N_11238,N_9838,N_10749);
nor U11239 (N_11239,N_9721,N_9740);
and U11240 (N_11240,N_9650,N_10131);
and U11241 (N_11241,N_10249,N_10025);
nand U11242 (N_11242,N_10450,N_10047);
and U11243 (N_11243,N_10399,N_10684);
and U11244 (N_11244,N_10604,N_10697);
and U11245 (N_11245,N_10476,N_10646);
and U11246 (N_11246,N_10068,N_10179);
and U11247 (N_11247,N_10786,N_10790);
or U11248 (N_11248,N_10026,N_9673);
nand U11249 (N_11249,N_9832,N_9811);
and U11250 (N_11250,N_9677,N_9916);
xor U11251 (N_11251,N_10763,N_10100);
nor U11252 (N_11252,N_9689,N_10446);
or U11253 (N_11253,N_9727,N_10348);
and U11254 (N_11254,N_10775,N_10123);
xnor U11255 (N_11255,N_9994,N_10190);
and U11256 (N_11256,N_9819,N_10038);
or U11257 (N_11257,N_9679,N_10035);
or U11258 (N_11258,N_9998,N_10708);
nand U11259 (N_11259,N_10546,N_9748);
xnor U11260 (N_11260,N_10509,N_10137);
nand U11261 (N_11261,N_10044,N_10750);
nand U11262 (N_11262,N_10761,N_10034);
xor U11263 (N_11263,N_10158,N_9924);
nand U11264 (N_11264,N_10223,N_9613);
xnor U11265 (N_11265,N_10558,N_9751);
nor U11266 (N_11266,N_9824,N_10662);
and U11267 (N_11267,N_10718,N_10341);
or U11268 (N_11268,N_9793,N_10325);
nand U11269 (N_11269,N_10107,N_10636);
nand U11270 (N_11270,N_10518,N_10601);
xor U11271 (N_11271,N_10648,N_10425);
or U11272 (N_11272,N_10713,N_10263);
or U11273 (N_11273,N_9907,N_10370);
or U11274 (N_11274,N_10286,N_10495);
and U11275 (N_11275,N_10517,N_10592);
or U11276 (N_11276,N_10742,N_10345);
and U11277 (N_11277,N_9696,N_10554);
xnor U11278 (N_11278,N_10134,N_9741);
nand U11279 (N_11279,N_9823,N_9801);
or U11280 (N_11280,N_10784,N_9668);
nand U11281 (N_11281,N_10496,N_10234);
xnor U11282 (N_11282,N_9639,N_9774);
nand U11283 (N_11283,N_10077,N_10124);
or U11284 (N_11284,N_10181,N_9637);
and U11285 (N_11285,N_9886,N_9864);
nand U11286 (N_11286,N_10395,N_9941);
nand U11287 (N_11287,N_10208,N_9937);
or U11288 (N_11288,N_10391,N_10204);
and U11289 (N_11289,N_10339,N_10415);
nand U11290 (N_11290,N_9626,N_10542);
and U11291 (N_11291,N_10093,N_10102);
xnor U11292 (N_11292,N_10132,N_10427);
nor U11293 (N_11293,N_10194,N_10238);
or U11294 (N_11294,N_10032,N_9813);
nor U11295 (N_11295,N_10319,N_9966);
nor U11296 (N_11296,N_10772,N_10344);
or U11297 (N_11297,N_9970,N_9989);
xnor U11298 (N_11298,N_10321,N_10788);
or U11299 (N_11299,N_10556,N_9870);
nor U11300 (N_11300,N_10532,N_10521);
or U11301 (N_11301,N_10063,N_9783);
nor U11302 (N_11302,N_10743,N_10191);
or U11303 (N_11303,N_10228,N_10187);
or U11304 (N_11304,N_9825,N_10240);
xor U11305 (N_11305,N_10367,N_9722);
and U11306 (N_11306,N_10699,N_10555);
nor U11307 (N_11307,N_10714,N_9725);
xnor U11308 (N_11308,N_9747,N_9961);
xor U11309 (N_11309,N_10582,N_10258);
xnor U11310 (N_11310,N_9919,N_10305);
xor U11311 (N_11311,N_10017,N_9794);
xor U11312 (N_11312,N_10505,N_10681);
xor U11313 (N_11313,N_10119,N_10265);
and U11314 (N_11314,N_9750,N_9629);
nor U11315 (N_11315,N_9800,N_9706);
or U11316 (N_11316,N_9605,N_9711);
xnor U11317 (N_11317,N_9666,N_10363);
xor U11318 (N_11318,N_10596,N_9759);
xnor U11319 (N_11319,N_9735,N_10126);
nand U11320 (N_11320,N_10650,N_10270);
xnor U11321 (N_11321,N_10117,N_9831);
xor U11322 (N_11322,N_10313,N_10357);
nand U11323 (N_11323,N_9896,N_9978);
nor U11324 (N_11324,N_10139,N_10520);
xor U11325 (N_11325,N_9867,N_10053);
nor U11326 (N_11326,N_10445,N_10255);
nor U11327 (N_11327,N_10251,N_9984);
or U11328 (N_11328,N_10756,N_9643);
or U11329 (N_11329,N_10442,N_10324);
nor U11330 (N_11330,N_10709,N_10410);
or U11331 (N_11331,N_10489,N_9621);
nand U11332 (N_11332,N_9855,N_9658);
xor U11333 (N_11333,N_10200,N_9842);
and U11334 (N_11334,N_10581,N_10589);
nor U11335 (N_11335,N_9820,N_9872);
xor U11336 (N_11336,N_9829,N_10122);
or U11337 (N_11337,N_10439,N_10740);
xnor U11338 (N_11338,N_10003,N_10770);
xnor U11339 (N_11339,N_9971,N_10774);
nor U11340 (N_11340,N_10021,N_10744);
nand U11341 (N_11341,N_10741,N_10584);
and U11342 (N_11342,N_9926,N_9645);
xor U11343 (N_11343,N_9719,N_9925);
or U11344 (N_11344,N_10014,N_9610);
or U11345 (N_11345,N_10388,N_9980);
and U11346 (N_11346,N_10631,N_9860);
nor U11347 (N_11347,N_10294,N_10384);
nand U11348 (N_11348,N_10207,N_10407);
and U11349 (N_11349,N_9608,N_9601);
xor U11350 (N_11350,N_10096,N_10703);
or U11351 (N_11351,N_10437,N_10323);
nand U11352 (N_11352,N_9904,N_10042);
and U11353 (N_11353,N_9849,N_10560);
and U11354 (N_11354,N_10156,N_10643);
xor U11355 (N_11355,N_9920,N_10070);
xor U11356 (N_11356,N_10566,N_9895);
xor U11357 (N_11357,N_10611,N_10061);
nand U11358 (N_11358,N_10335,N_9883);
nand U11359 (N_11359,N_10561,N_10459);
and U11360 (N_11360,N_10023,N_10779);
xnor U11361 (N_11361,N_10086,N_10479);
nor U11362 (N_11362,N_10209,N_10302);
nand U11363 (N_11363,N_10679,N_10051);
or U11364 (N_11364,N_9726,N_9900);
or U11365 (N_11365,N_10136,N_10738);
xnor U11366 (N_11366,N_9627,N_9663);
or U11367 (N_11367,N_10519,N_9889);
nand U11368 (N_11368,N_10135,N_10534);
xor U11369 (N_11369,N_10185,N_10448);
nand U11370 (N_11370,N_10371,N_10298);
nand U11371 (N_11371,N_10635,N_10049);
nand U11372 (N_11372,N_9908,N_10618);
nand U11373 (N_11373,N_10688,N_10424);
or U11374 (N_11374,N_10421,N_10717);
and U11375 (N_11375,N_9921,N_10092);
and U11376 (N_11376,N_10050,N_10082);
or U11377 (N_11377,N_10027,N_10060);
or U11378 (N_11378,N_10211,N_9918);
nand U11379 (N_11379,N_10214,N_10172);
or U11380 (N_11380,N_10469,N_10403);
or U11381 (N_11381,N_9652,N_9662);
nand U11382 (N_11382,N_10570,N_9633);
or U11383 (N_11383,N_9660,N_9839);
or U11384 (N_11384,N_10048,N_9640);
or U11385 (N_11385,N_9654,N_10154);
nand U11386 (N_11386,N_10797,N_9891);
and U11387 (N_11387,N_9806,N_9950);
xor U11388 (N_11388,N_10730,N_10165);
nor U11389 (N_11389,N_10548,N_10346);
nor U11390 (N_11390,N_9703,N_10401);
xor U11391 (N_11391,N_10537,N_9893);
nand U11392 (N_11392,N_9651,N_9875);
or U11393 (N_11393,N_10283,N_10588);
nand U11394 (N_11394,N_10766,N_10010);
nand U11395 (N_11395,N_9928,N_10148);
nor U11396 (N_11396,N_10128,N_10336);
nor U11397 (N_11397,N_9749,N_10188);
or U11398 (N_11398,N_9821,N_10433);
and U11399 (N_11399,N_10330,N_10591);
nand U11400 (N_11400,N_10654,N_10312);
nor U11401 (N_11401,N_10647,N_10269);
xnor U11402 (N_11402,N_10373,N_9788);
or U11403 (N_11403,N_10668,N_10362);
and U11404 (N_11404,N_10064,N_9867);
nor U11405 (N_11405,N_10137,N_9852);
nor U11406 (N_11406,N_10758,N_9660);
and U11407 (N_11407,N_10432,N_10202);
nor U11408 (N_11408,N_10784,N_10620);
nand U11409 (N_11409,N_10632,N_10018);
nand U11410 (N_11410,N_10619,N_10312);
and U11411 (N_11411,N_9834,N_9745);
and U11412 (N_11412,N_10429,N_10624);
or U11413 (N_11413,N_10463,N_10651);
or U11414 (N_11414,N_10355,N_10099);
nand U11415 (N_11415,N_10164,N_10335);
and U11416 (N_11416,N_10565,N_9653);
nand U11417 (N_11417,N_10784,N_10552);
nor U11418 (N_11418,N_10059,N_9942);
nor U11419 (N_11419,N_10591,N_10771);
and U11420 (N_11420,N_10359,N_9661);
and U11421 (N_11421,N_10168,N_10198);
and U11422 (N_11422,N_9970,N_10227);
nand U11423 (N_11423,N_10167,N_10113);
nor U11424 (N_11424,N_10532,N_9741);
or U11425 (N_11425,N_9795,N_10462);
nor U11426 (N_11426,N_10386,N_10162);
nand U11427 (N_11427,N_10295,N_9975);
nand U11428 (N_11428,N_10277,N_10011);
nand U11429 (N_11429,N_10737,N_9884);
and U11430 (N_11430,N_10682,N_9985);
or U11431 (N_11431,N_10712,N_9857);
nand U11432 (N_11432,N_10267,N_10122);
nand U11433 (N_11433,N_10659,N_9619);
and U11434 (N_11434,N_10247,N_9670);
nor U11435 (N_11435,N_9803,N_10147);
nand U11436 (N_11436,N_10462,N_10068);
xor U11437 (N_11437,N_10486,N_10366);
and U11438 (N_11438,N_10730,N_9824);
xnor U11439 (N_11439,N_9684,N_10693);
and U11440 (N_11440,N_10638,N_10797);
xnor U11441 (N_11441,N_10620,N_10183);
or U11442 (N_11442,N_10424,N_10765);
or U11443 (N_11443,N_9813,N_10503);
xnor U11444 (N_11444,N_9897,N_9931);
and U11445 (N_11445,N_10474,N_9724);
nand U11446 (N_11446,N_9809,N_10009);
xnor U11447 (N_11447,N_10107,N_10643);
or U11448 (N_11448,N_10232,N_9611);
and U11449 (N_11449,N_10052,N_10786);
nor U11450 (N_11450,N_9716,N_10223);
nor U11451 (N_11451,N_10447,N_10200);
nor U11452 (N_11452,N_10152,N_10231);
and U11453 (N_11453,N_9843,N_10777);
nor U11454 (N_11454,N_10522,N_10540);
and U11455 (N_11455,N_10722,N_10584);
nand U11456 (N_11456,N_10770,N_10099);
and U11457 (N_11457,N_10298,N_10006);
xnor U11458 (N_11458,N_9901,N_10660);
or U11459 (N_11459,N_9668,N_10374);
nand U11460 (N_11460,N_10121,N_10516);
xor U11461 (N_11461,N_9886,N_10502);
and U11462 (N_11462,N_10000,N_10673);
nand U11463 (N_11463,N_9705,N_10725);
nor U11464 (N_11464,N_10086,N_10024);
xnor U11465 (N_11465,N_10150,N_9817);
and U11466 (N_11466,N_9630,N_9913);
and U11467 (N_11467,N_10289,N_9729);
nand U11468 (N_11468,N_10052,N_10779);
nor U11469 (N_11469,N_10778,N_10707);
and U11470 (N_11470,N_10029,N_10076);
or U11471 (N_11471,N_10273,N_10361);
and U11472 (N_11472,N_9856,N_9884);
nand U11473 (N_11473,N_10694,N_10565);
nand U11474 (N_11474,N_10448,N_9661);
nand U11475 (N_11475,N_10401,N_9622);
or U11476 (N_11476,N_10047,N_10586);
and U11477 (N_11477,N_9829,N_10160);
or U11478 (N_11478,N_9899,N_10056);
nand U11479 (N_11479,N_10170,N_10168);
and U11480 (N_11480,N_9912,N_10278);
xnor U11481 (N_11481,N_9722,N_9949);
or U11482 (N_11482,N_10408,N_9611);
nand U11483 (N_11483,N_10182,N_10175);
nand U11484 (N_11484,N_10697,N_9644);
nand U11485 (N_11485,N_9629,N_9735);
or U11486 (N_11486,N_10397,N_10487);
or U11487 (N_11487,N_10247,N_9808);
and U11488 (N_11488,N_10110,N_10356);
xor U11489 (N_11489,N_10732,N_10102);
and U11490 (N_11490,N_10130,N_9909);
nand U11491 (N_11491,N_9788,N_10085);
or U11492 (N_11492,N_10636,N_10456);
nor U11493 (N_11493,N_10705,N_10091);
xor U11494 (N_11494,N_10775,N_10622);
nor U11495 (N_11495,N_10672,N_9738);
nand U11496 (N_11496,N_10585,N_9821);
nand U11497 (N_11497,N_9854,N_10090);
and U11498 (N_11498,N_10631,N_10180);
nor U11499 (N_11499,N_10139,N_10157);
nor U11500 (N_11500,N_9863,N_9682);
nor U11501 (N_11501,N_10765,N_10285);
or U11502 (N_11502,N_10589,N_9728);
nor U11503 (N_11503,N_10122,N_10569);
and U11504 (N_11504,N_10475,N_10305);
or U11505 (N_11505,N_10365,N_10560);
nand U11506 (N_11506,N_9776,N_10095);
xnor U11507 (N_11507,N_9940,N_10302);
and U11508 (N_11508,N_10662,N_10493);
nor U11509 (N_11509,N_9964,N_9912);
nor U11510 (N_11510,N_10433,N_10589);
or U11511 (N_11511,N_9783,N_10451);
nand U11512 (N_11512,N_10344,N_10636);
nand U11513 (N_11513,N_10496,N_10181);
xor U11514 (N_11514,N_9993,N_10298);
and U11515 (N_11515,N_9814,N_10772);
nand U11516 (N_11516,N_9620,N_9641);
nor U11517 (N_11517,N_10401,N_10340);
xnor U11518 (N_11518,N_10041,N_10444);
nand U11519 (N_11519,N_10491,N_10293);
nor U11520 (N_11520,N_10598,N_9698);
nor U11521 (N_11521,N_10731,N_10359);
nand U11522 (N_11522,N_9853,N_10705);
or U11523 (N_11523,N_10488,N_9765);
or U11524 (N_11524,N_10373,N_10309);
xnor U11525 (N_11525,N_10772,N_10725);
or U11526 (N_11526,N_10477,N_10081);
nand U11527 (N_11527,N_10728,N_10009);
nor U11528 (N_11528,N_10120,N_10752);
nor U11529 (N_11529,N_10230,N_10014);
or U11530 (N_11530,N_10619,N_10121);
or U11531 (N_11531,N_9762,N_10387);
nor U11532 (N_11532,N_9912,N_9888);
or U11533 (N_11533,N_9872,N_10531);
and U11534 (N_11534,N_10372,N_10278);
and U11535 (N_11535,N_9627,N_9886);
xor U11536 (N_11536,N_10642,N_9679);
or U11537 (N_11537,N_10441,N_9612);
or U11538 (N_11538,N_10253,N_9645);
xor U11539 (N_11539,N_10691,N_10132);
and U11540 (N_11540,N_10033,N_10032);
and U11541 (N_11541,N_10104,N_10781);
nor U11542 (N_11542,N_10758,N_10515);
and U11543 (N_11543,N_10180,N_10229);
or U11544 (N_11544,N_10460,N_9996);
xor U11545 (N_11545,N_10662,N_10762);
nor U11546 (N_11546,N_9681,N_10445);
and U11547 (N_11547,N_10472,N_10684);
xor U11548 (N_11548,N_10481,N_9921);
or U11549 (N_11549,N_9939,N_10652);
nor U11550 (N_11550,N_10699,N_9992);
and U11551 (N_11551,N_9610,N_10061);
and U11552 (N_11552,N_9705,N_10512);
or U11553 (N_11553,N_10000,N_9959);
nor U11554 (N_11554,N_10379,N_10748);
nor U11555 (N_11555,N_9693,N_9807);
nor U11556 (N_11556,N_10521,N_10163);
xnor U11557 (N_11557,N_10081,N_9666);
xor U11558 (N_11558,N_10154,N_9610);
or U11559 (N_11559,N_10374,N_10401);
xor U11560 (N_11560,N_10700,N_10365);
nand U11561 (N_11561,N_9865,N_10229);
and U11562 (N_11562,N_10421,N_10199);
and U11563 (N_11563,N_9842,N_10349);
or U11564 (N_11564,N_9929,N_10313);
nor U11565 (N_11565,N_10514,N_9824);
xor U11566 (N_11566,N_10527,N_9748);
xnor U11567 (N_11567,N_10443,N_10573);
nand U11568 (N_11568,N_10328,N_9851);
nor U11569 (N_11569,N_9789,N_10557);
xnor U11570 (N_11570,N_9625,N_9889);
nand U11571 (N_11571,N_10735,N_10584);
nand U11572 (N_11572,N_10481,N_10733);
xor U11573 (N_11573,N_10073,N_10141);
and U11574 (N_11574,N_10567,N_10327);
nor U11575 (N_11575,N_10150,N_9670);
nor U11576 (N_11576,N_9930,N_9729);
or U11577 (N_11577,N_10502,N_10128);
xnor U11578 (N_11578,N_10678,N_9937);
or U11579 (N_11579,N_9818,N_9614);
and U11580 (N_11580,N_10557,N_10776);
xor U11581 (N_11581,N_9849,N_10025);
xnor U11582 (N_11582,N_9802,N_9809);
and U11583 (N_11583,N_9611,N_10259);
xor U11584 (N_11584,N_9678,N_9921);
nor U11585 (N_11585,N_9787,N_9801);
xnor U11586 (N_11586,N_9601,N_9826);
or U11587 (N_11587,N_10171,N_9755);
or U11588 (N_11588,N_10247,N_9841);
xnor U11589 (N_11589,N_10042,N_10120);
or U11590 (N_11590,N_10249,N_9617);
and U11591 (N_11591,N_10443,N_9893);
nand U11592 (N_11592,N_10272,N_9673);
nand U11593 (N_11593,N_10524,N_10734);
and U11594 (N_11594,N_10022,N_10300);
and U11595 (N_11595,N_9694,N_9680);
nor U11596 (N_11596,N_10733,N_10008);
xnor U11597 (N_11597,N_10116,N_9890);
and U11598 (N_11598,N_10707,N_9924);
xnor U11599 (N_11599,N_10506,N_10013);
nand U11600 (N_11600,N_10146,N_9633);
nand U11601 (N_11601,N_9837,N_9737);
nor U11602 (N_11602,N_10365,N_9683);
and U11603 (N_11603,N_9900,N_10316);
xor U11604 (N_11604,N_10734,N_10756);
and U11605 (N_11605,N_10212,N_9976);
or U11606 (N_11606,N_10486,N_9734);
or U11607 (N_11607,N_9993,N_10037);
xnor U11608 (N_11608,N_10120,N_9641);
nand U11609 (N_11609,N_10030,N_10079);
nand U11610 (N_11610,N_9670,N_10641);
nand U11611 (N_11611,N_10417,N_9966);
xor U11612 (N_11612,N_10194,N_10437);
xor U11613 (N_11613,N_10312,N_9630);
nor U11614 (N_11614,N_10401,N_10674);
or U11615 (N_11615,N_10075,N_10219);
nor U11616 (N_11616,N_10067,N_9801);
or U11617 (N_11617,N_10605,N_9939);
xnor U11618 (N_11618,N_10233,N_10192);
and U11619 (N_11619,N_10002,N_9614);
nand U11620 (N_11620,N_10451,N_10053);
and U11621 (N_11621,N_10332,N_9794);
or U11622 (N_11622,N_10040,N_10434);
and U11623 (N_11623,N_10231,N_10359);
xnor U11624 (N_11624,N_9712,N_10102);
or U11625 (N_11625,N_9841,N_9755);
nor U11626 (N_11626,N_9662,N_10273);
or U11627 (N_11627,N_10653,N_10023);
nor U11628 (N_11628,N_9719,N_9741);
nor U11629 (N_11629,N_10385,N_10558);
xor U11630 (N_11630,N_9942,N_9796);
xnor U11631 (N_11631,N_9730,N_9818);
or U11632 (N_11632,N_10652,N_10539);
nand U11633 (N_11633,N_10527,N_10287);
and U11634 (N_11634,N_10755,N_10096);
nand U11635 (N_11635,N_9735,N_9760);
or U11636 (N_11636,N_10102,N_10685);
xnor U11637 (N_11637,N_9918,N_10180);
xor U11638 (N_11638,N_9666,N_10149);
nor U11639 (N_11639,N_10086,N_10323);
nor U11640 (N_11640,N_10430,N_10230);
xor U11641 (N_11641,N_10609,N_10561);
nand U11642 (N_11642,N_9939,N_10658);
and U11643 (N_11643,N_9772,N_10703);
nand U11644 (N_11644,N_10327,N_10312);
nand U11645 (N_11645,N_10376,N_10776);
nor U11646 (N_11646,N_10100,N_9887);
nor U11647 (N_11647,N_10545,N_9956);
and U11648 (N_11648,N_9893,N_9909);
and U11649 (N_11649,N_9748,N_9795);
and U11650 (N_11650,N_10037,N_10080);
xnor U11651 (N_11651,N_10139,N_10456);
or U11652 (N_11652,N_9983,N_10650);
nand U11653 (N_11653,N_9745,N_10443);
nor U11654 (N_11654,N_9904,N_10329);
xor U11655 (N_11655,N_10537,N_9635);
nand U11656 (N_11656,N_9836,N_10398);
or U11657 (N_11657,N_10764,N_10408);
and U11658 (N_11658,N_9848,N_10252);
nor U11659 (N_11659,N_10365,N_10053);
or U11660 (N_11660,N_10095,N_10772);
nand U11661 (N_11661,N_10098,N_10595);
and U11662 (N_11662,N_10223,N_10209);
or U11663 (N_11663,N_10722,N_10282);
or U11664 (N_11664,N_10258,N_10041);
and U11665 (N_11665,N_10540,N_9815);
or U11666 (N_11666,N_10299,N_9617);
xnor U11667 (N_11667,N_10372,N_9911);
nand U11668 (N_11668,N_9664,N_9770);
nor U11669 (N_11669,N_10453,N_10732);
xor U11670 (N_11670,N_10029,N_10798);
or U11671 (N_11671,N_10456,N_9906);
nand U11672 (N_11672,N_10667,N_10511);
nand U11673 (N_11673,N_10108,N_10568);
nor U11674 (N_11674,N_10664,N_9985);
xnor U11675 (N_11675,N_9660,N_10465);
xnor U11676 (N_11676,N_9864,N_10396);
xor U11677 (N_11677,N_9960,N_9623);
and U11678 (N_11678,N_10496,N_10350);
nand U11679 (N_11679,N_9643,N_10061);
xnor U11680 (N_11680,N_10706,N_9729);
or U11681 (N_11681,N_9735,N_9655);
and U11682 (N_11682,N_9601,N_10777);
or U11683 (N_11683,N_10277,N_10572);
or U11684 (N_11684,N_10001,N_10086);
xnor U11685 (N_11685,N_10010,N_10176);
nor U11686 (N_11686,N_9965,N_10671);
nand U11687 (N_11687,N_9854,N_10121);
nor U11688 (N_11688,N_10434,N_9878);
nor U11689 (N_11689,N_10188,N_10319);
or U11690 (N_11690,N_9763,N_10524);
xnor U11691 (N_11691,N_9857,N_10324);
and U11692 (N_11692,N_10153,N_10030);
xor U11693 (N_11693,N_10022,N_9862);
nor U11694 (N_11694,N_9644,N_10795);
or U11695 (N_11695,N_10777,N_9759);
nand U11696 (N_11696,N_9864,N_10720);
xnor U11697 (N_11697,N_9609,N_9757);
xor U11698 (N_11698,N_10355,N_9849);
nand U11699 (N_11699,N_9979,N_10367);
or U11700 (N_11700,N_10270,N_9646);
nor U11701 (N_11701,N_9950,N_10140);
or U11702 (N_11702,N_9928,N_9746);
nand U11703 (N_11703,N_9696,N_9872);
and U11704 (N_11704,N_9774,N_10050);
xnor U11705 (N_11705,N_10703,N_10368);
or U11706 (N_11706,N_10780,N_10068);
or U11707 (N_11707,N_9625,N_10168);
and U11708 (N_11708,N_10659,N_10088);
xnor U11709 (N_11709,N_9714,N_10507);
or U11710 (N_11710,N_10020,N_9633);
or U11711 (N_11711,N_9912,N_10194);
xor U11712 (N_11712,N_10533,N_10059);
and U11713 (N_11713,N_10222,N_10314);
xor U11714 (N_11714,N_9907,N_10693);
xor U11715 (N_11715,N_10497,N_9693);
or U11716 (N_11716,N_9902,N_9929);
xor U11717 (N_11717,N_10113,N_9803);
xnor U11718 (N_11718,N_10104,N_9617);
nor U11719 (N_11719,N_10172,N_10548);
or U11720 (N_11720,N_9726,N_9778);
nor U11721 (N_11721,N_10731,N_9646);
nand U11722 (N_11722,N_10753,N_10366);
and U11723 (N_11723,N_10031,N_10778);
nor U11724 (N_11724,N_9913,N_9982);
and U11725 (N_11725,N_10479,N_9998);
and U11726 (N_11726,N_9759,N_10518);
and U11727 (N_11727,N_10014,N_10363);
nor U11728 (N_11728,N_10655,N_9812);
nand U11729 (N_11729,N_10101,N_9979);
nor U11730 (N_11730,N_9988,N_9709);
nor U11731 (N_11731,N_10133,N_10706);
or U11732 (N_11732,N_9843,N_10304);
nor U11733 (N_11733,N_10769,N_10462);
and U11734 (N_11734,N_10030,N_9827);
xnor U11735 (N_11735,N_10214,N_9814);
xnor U11736 (N_11736,N_10598,N_10563);
xor U11737 (N_11737,N_10789,N_9842);
and U11738 (N_11738,N_9685,N_10662);
nor U11739 (N_11739,N_9797,N_9721);
nor U11740 (N_11740,N_10368,N_9805);
or U11741 (N_11741,N_10127,N_10574);
xnor U11742 (N_11742,N_10428,N_10244);
xnor U11743 (N_11743,N_9750,N_10672);
xor U11744 (N_11744,N_10029,N_9821);
nor U11745 (N_11745,N_10715,N_9707);
and U11746 (N_11746,N_10399,N_9720);
xor U11747 (N_11747,N_9891,N_10366);
nor U11748 (N_11748,N_10662,N_9745);
or U11749 (N_11749,N_10414,N_9761);
nand U11750 (N_11750,N_9717,N_9875);
nor U11751 (N_11751,N_9866,N_10272);
nand U11752 (N_11752,N_9604,N_10473);
nor U11753 (N_11753,N_9863,N_10068);
or U11754 (N_11754,N_9749,N_10744);
nor U11755 (N_11755,N_10650,N_10562);
and U11756 (N_11756,N_9763,N_9617);
nand U11757 (N_11757,N_10269,N_9817);
or U11758 (N_11758,N_9601,N_10672);
nor U11759 (N_11759,N_10202,N_10339);
or U11760 (N_11760,N_9724,N_10019);
and U11761 (N_11761,N_10591,N_10751);
or U11762 (N_11762,N_9654,N_10208);
xnor U11763 (N_11763,N_10430,N_10650);
xor U11764 (N_11764,N_9662,N_9661);
or U11765 (N_11765,N_10625,N_9896);
nand U11766 (N_11766,N_10284,N_9675);
nand U11767 (N_11767,N_10490,N_10647);
nor U11768 (N_11768,N_10396,N_10536);
xor U11769 (N_11769,N_9883,N_9745);
xnor U11770 (N_11770,N_9814,N_10162);
and U11771 (N_11771,N_10636,N_10687);
and U11772 (N_11772,N_10286,N_10325);
xor U11773 (N_11773,N_9649,N_10298);
and U11774 (N_11774,N_10678,N_10097);
xnor U11775 (N_11775,N_10231,N_10700);
nor U11776 (N_11776,N_9935,N_10508);
nand U11777 (N_11777,N_10622,N_10022);
nand U11778 (N_11778,N_10626,N_10332);
nor U11779 (N_11779,N_9716,N_10027);
nand U11780 (N_11780,N_10450,N_10790);
and U11781 (N_11781,N_10746,N_9731);
or U11782 (N_11782,N_10797,N_9830);
xnor U11783 (N_11783,N_9606,N_9801);
xnor U11784 (N_11784,N_10708,N_10754);
or U11785 (N_11785,N_9793,N_9659);
nand U11786 (N_11786,N_9802,N_10199);
nor U11787 (N_11787,N_9863,N_9825);
xnor U11788 (N_11788,N_10219,N_10742);
nor U11789 (N_11789,N_10674,N_10067);
or U11790 (N_11790,N_9708,N_10043);
xnor U11791 (N_11791,N_9684,N_10304);
xor U11792 (N_11792,N_10359,N_9805);
or U11793 (N_11793,N_10595,N_10554);
nand U11794 (N_11794,N_10707,N_10047);
or U11795 (N_11795,N_9944,N_10676);
nor U11796 (N_11796,N_9771,N_9702);
nand U11797 (N_11797,N_10393,N_10184);
nor U11798 (N_11798,N_9624,N_10382);
xor U11799 (N_11799,N_10568,N_9892);
xnor U11800 (N_11800,N_9950,N_10172);
xnor U11801 (N_11801,N_9956,N_10790);
xnor U11802 (N_11802,N_9963,N_9674);
nor U11803 (N_11803,N_10089,N_10765);
nor U11804 (N_11804,N_10174,N_10572);
or U11805 (N_11805,N_9874,N_9749);
nand U11806 (N_11806,N_10665,N_10561);
or U11807 (N_11807,N_10050,N_9690);
nand U11808 (N_11808,N_10576,N_10052);
xnor U11809 (N_11809,N_10525,N_9800);
or U11810 (N_11810,N_10103,N_9832);
nand U11811 (N_11811,N_10142,N_9612);
nor U11812 (N_11812,N_9732,N_9602);
xnor U11813 (N_11813,N_10460,N_10582);
and U11814 (N_11814,N_10394,N_10250);
xnor U11815 (N_11815,N_10329,N_10429);
nor U11816 (N_11816,N_10107,N_10124);
and U11817 (N_11817,N_10794,N_9671);
xor U11818 (N_11818,N_10448,N_9996);
xor U11819 (N_11819,N_10133,N_9642);
nand U11820 (N_11820,N_10349,N_10709);
or U11821 (N_11821,N_9654,N_9922);
xor U11822 (N_11822,N_9884,N_10706);
xor U11823 (N_11823,N_10321,N_9745);
nor U11824 (N_11824,N_10295,N_9637);
nand U11825 (N_11825,N_10566,N_9879);
nor U11826 (N_11826,N_10128,N_10540);
and U11827 (N_11827,N_9888,N_9600);
nand U11828 (N_11828,N_9737,N_9750);
or U11829 (N_11829,N_10274,N_10763);
xor U11830 (N_11830,N_10224,N_10431);
or U11831 (N_11831,N_9674,N_10672);
nor U11832 (N_11832,N_10583,N_10460);
xnor U11833 (N_11833,N_10651,N_10150);
and U11834 (N_11834,N_10218,N_10489);
or U11835 (N_11835,N_10177,N_10773);
xnor U11836 (N_11836,N_10210,N_9972);
nor U11837 (N_11837,N_10775,N_9673);
and U11838 (N_11838,N_10520,N_9835);
nor U11839 (N_11839,N_10704,N_10687);
nand U11840 (N_11840,N_10076,N_10117);
xnor U11841 (N_11841,N_9907,N_10467);
and U11842 (N_11842,N_10654,N_10577);
xor U11843 (N_11843,N_10224,N_10550);
nand U11844 (N_11844,N_10583,N_10248);
or U11845 (N_11845,N_9846,N_9703);
or U11846 (N_11846,N_10158,N_9794);
xnor U11847 (N_11847,N_10583,N_10749);
and U11848 (N_11848,N_10098,N_10467);
or U11849 (N_11849,N_10438,N_9836);
xor U11850 (N_11850,N_10239,N_9826);
or U11851 (N_11851,N_9876,N_10374);
nor U11852 (N_11852,N_9660,N_10369);
xor U11853 (N_11853,N_9647,N_9650);
nor U11854 (N_11854,N_10512,N_9636);
and U11855 (N_11855,N_9688,N_10136);
xor U11856 (N_11856,N_10140,N_9863);
or U11857 (N_11857,N_9912,N_9626);
and U11858 (N_11858,N_9760,N_10132);
xnor U11859 (N_11859,N_10594,N_10224);
nand U11860 (N_11860,N_9834,N_9936);
and U11861 (N_11861,N_9646,N_9885);
nor U11862 (N_11862,N_10265,N_9866);
nor U11863 (N_11863,N_10576,N_10077);
and U11864 (N_11864,N_10272,N_9701);
or U11865 (N_11865,N_9786,N_10206);
xnor U11866 (N_11866,N_10045,N_9683);
nand U11867 (N_11867,N_9641,N_9640);
nor U11868 (N_11868,N_10136,N_9675);
xnor U11869 (N_11869,N_10316,N_9910);
or U11870 (N_11870,N_9854,N_10652);
or U11871 (N_11871,N_9637,N_10220);
or U11872 (N_11872,N_9955,N_10768);
or U11873 (N_11873,N_9807,N_10018);
and U11874 (N_11874,N_10601,N_10183);
and U11875 (N_11875,N_10365,N_10760);
nor U11876 (N_11876,N_9966,N_10622);
nand U11877 (N_11877,N_10643,N_9656);
nand U11878 (N_11878,N_9842,N_9937);
nor U11879 (N_11879,N_10168,N_9702);
and U11880 (N_11880,N_9814,N_9908);
or U11881 (N_11881,N_10722,N_9667);
nand U11882 (N_11882,N_10589,N_10252);
or U11883 (N_11883,N_9625,N_10378);
nand U11884 (N_11884,N_9902,N_10576);
xor U11885 (N_11885,N_9636,N_9808);
xor U11886 (N_11886,N_9674,N_10557);
nand U11887 (N_11887,N_10523,N_9774);
xnor U11888 (N_11888,N_10307,N_10661);
nand U11889 (N_11889,N_10408,N_9903);
xor U11890 (N_11890,N_9851,N_10553);
or U11891 (N_11891,N_10118,N_10522);
nor U11892 (N_11892,N_10350,N_9999);
or U11893 (N_11893,N_10703,N_10629);
xor U11894 (N_11894,N_10648,N_10797);
and U11895 (N_11895,N_9812,N_10068);
nand U11896 (N_11896,N_9836,N_10471);
and U11897 (N_11897,N_9766,N_10752);
nand U11898 (N_11898,N_10715,N_10626);
nor U11899 (N_11899,N_10272,N_10218);
and U11900 (N_11900,N_10501,N_10619);
xor U11901 (N_11901,N_9692,N_10148);
or U11902 (N_11902,N_9765,N_10772);
nor U11903 (N_11903,N_9841,N_10677);
or U11904 (N_11904,N_10396,N_9901);
nor U11905 (N_11905,N_10510,N_10167);
xor U11906 (N_11906,N_10023,N_10522);
nor U11907 (N_11907,N_10157,N_9859);
or U11908 (N_11908,N_10252,N_10472);
nand U11909 (N_11909,N_9674,N_10538);
and U11910 (N_11910,N_10313,N_9784);
and U11911 (N_11911,N_10265,N_10002);
nand U11912 (N_11912,N_10010,N_10064);
nand U11913 (N_11913,N_10473,N_10650);
and U11914 (N_11914,N_10797,N_10725);
or U11915 (N_11915,N_9804,N_10325);
and U11916 (N_11916,N_10646,N_10246);
xor U11917 (N_11917,N_9611,N_9770);
and U11918 (N_11918,N_9642,N_10412);
and U11919 (N_11919,N_10397,N_10339);
nand U11920 (N_11920,N_10083,N_10550);
nand U11921 (N_11921,N_10273,N_10394);
xnor U11922 (N_11922,N_9974,N_9762);
xnor U11923 (N_11923,N_10599,N_9923);
or U11924 (N_11924,N_9792,N_10575);
xor U11925 (N_11925,N_9904,N_9765);
or U11926 (N_11926,N_10672,N_10090);
or U11927 (N_11927,N_10229,N_10736);
and U11928 (N_11928,N_9624,N_10571);
nand U11929 (N_11929,N_10108,N_9671);
xor U11930 (N_11930,N_10169,N_10736);
xnor U11931 (N_11931,N_9823,N_9788);
nor U11932 (N_11932,N_9968,N_10640);
or U11933 (N_11933,N_10041,N_9965);
nor U11934 (N_11934,N_9842,N_9985);
nor U11935 (N_11935,N_10382,N_10479);
xnor U11936 (N_11936,N_9921,N_10148);
xnor U11937 (N_11937,N_10454,N_10300);
xnor U11938 (N_11938,N_10528,N_9659);
or U11939 (N_11939,N_10748,N_10217);
nor U11940 (N_11940,N_10382,N_10620);
and U11941 (N_11941,N_10636,N_9820);
nor U11942 (N_11942,N_10735,N_10509);
nand U11943 (N_11943,N_10286,N_9865);
nand U11944 (N_11944,N_10440,N_10723);
xnor U11945 (N_11945,N_10110,N_10433);
nand U11946 (N_11946,N_9615,N_9661);
and U11947 (N_11947,N_9954,N_10705);
xnor U11948 (N_11948,N_10454,N_10563);
nand U11949 (N_11949,N_9939,N_10192);
xor U11950 (N_11950,N_10228,N_10217);
xor U11951 (N_11951,N_10373,N_10407);
xnor U11952 (N_11952,N_9657,N_10127);
xor U11953 (N_11953,N_9743,N_10059);
or U11954 (N_11954,N_10648,N_10311);
nand U11955 (N_11955,N_10648,N_9730);
nor U11956 (N_11956,N_10640,N_10099);
nand U11957 (N_11957,N_10125,N_10472);
xnor U11958 (N_11958,N_10392,N_10246);
nand U11959 (N_11959,N_10212,N_10179);
xor U11960 (N_11960,N_10279,N_10093);
and U11961 (N_11961,N_10051,N_10068);
nor U11962 (N_11962,N_10246,N_9807);
or U11963 (N_11963,N_10442,N_10486);
or U11964 (N_11964,N_9985,N_10300);
nor U11965 (N_11965,N_9958,N_10386);
and U11966 (N_11966,N_10782,N_10548);
nor U11967 (N_11967,N_10312,N_10028);
and U11968 (N_11968,N_9764,N_10654);
xor U11969 (N_11969,N_10223,N_10060);
nand U11970 (N_11970,N_10651,N_9988);
nor U11971 (N_11971,N_10794,N_10430);
xor U11972 (N_11972,N_9896,N_10525);
and U11973 (N_11973,N_10087,N_9721);
nor U11974 (N_11974,N_10518,N_10038);
nand U11975 (N_11975,N_9600,N_9858);
and U11976 (N_11976,N_10443,N_10411);
xor U11977 (N_11977,N_9637,N_9604);
or U11978 (N_11978,N_10379,N_9693);
xor U11979 (N_11979,N_10146,N_10584);
or U11980 (N_11980,N_10298,N_10565);
and U11981 (N_11981,N_9764,N_10622);
nand U11982 (N_11982,N_10146,N_9728);
or U11983 (N_11983,N_9946,N_10388);
nand U11984 (N_11984,N_10704,N_10640);
nor U11985 (N_11985,N_10303,N_9989);
or U11986 (N_11986,N_10134,N_10385);
xor U11987 (N_11987,N_9612,N_10722);
and U11988 (N_11988,N_10346,N_9721);
xor U11989 (N_11989,N_9670,N_10121);
or U11990 (N_11990,N_10428,N_10046);
xnor U11991 (N_11991,N_9894,N_9869);
and U11992 (N_11992,N_10358,N_9976);
nand U11993 (N_11993,N_10123,N_9974);
nand U11994 (N_11994,N_9752,N_10456);
xnor U11995 (N_11995,N_9807,N_10187);
and U11996 (N_11996,N_10428,N_10331);
and U11997 (N_11997,N_10052,N_10745);
and U11998 (N_11998,N_10516,N_9707);
nand U11999 (N_11999,N_9707,N_9906);
nand U12000 (N_12000,N_10894,N_11637);
xor U12001 (N_12001,N_11825,N_11633);
or U12002 (N_12002,N_11618,N_11765);
nand U12003 (N_12003,N_11542,N_11446);
or U12004 (N_12004,N_11305,N_11750);
xnor U12005 (N_12005,N_11128,N_11927);
nand U12006 (N_12006,N_11298,N_10952);
nand U12007 (N_12007,N_11396,N_11784);
nor U12008 (N_12008,N_11878,N_11019);
nor U12009 (N_12009,N_11594,N_11081);
nor U12010 (N_12010,N_11501,N_10804);
nand U12011 (N_12011,N_11476,N_11924);
nand U12012 (N_12012,N_11318,N_10917);
and U12013 (N_12013,N_11808,N_11810);
and U12014 (N_12014,N_11402,N_11068);
nand U12015 (N_12015,N_11003,N_11150);
or U12016 (N_12016,N_11353,N_11778);
nand U12017 (N_12017,N_11741,N_11856);
nor U12018 (N_12018,N_10911,N_11336);
nor U12019 (N_12019,N_11214,N_11945);
xnor U12020 (N_12020,N_11267,N_11204);
and U12021 (N_12021,N_10995,N_11442);
nor U12022 (N_12022,N_11184,N_11883);
nand U12023 (N_12023,N_11950,N_11274);
nor U12024 (N_12024,N_11827,N_11754);
and U12025 (N_12025,N_11839,N_11588);
or U12026 (N_12026,N_11217,N_10964);
or U12027 (N_12027,N_11358,N_10933);
nor U12028 (N_12028,N_10946,N_11270);
xnor U12029 (N_12029,N_10969,N_11246);
and U12030 (N_12030,N_11243,N_11682);
and U12031 (N_12031,N_11419,N_10927);
xnor U12032 (N_12032,N_11958,N_11207);
and U12033 (N_12033,N_11236,N_11212);
nand U12034 (N_12034,N_11561,N_11586);
nor U12035 (N_12035,N_11356,N_11707);
and U12036 (N_12036,N_11711,N_10880);
xnor U12037 (N_12037,N_11040,N_11447);
and U12038 (N_12038,N_11727,N_11604);
and U12039 (N_12039,N_11884,N_11209);
nand U12040 (N_12040,N_11621,N_11263);
nor U12041 (N_12041,N_11905,N_11490);
and U12042 (N_12042,N_11891,N_10943);
or U12043 (N_12043,N_11971,N_11534);
xnor U12044 (N_12044,N_11758,N_11027);
and U12045 (N_12045,N_11287,N_11873);
and U12046 (N_12046,N_11262,N_11355);
nand U12047 (N_12047,N_11533,N_10826);
nand U12048 (N_12048,N_11496,N_10827);
nand U12049 (N_12049,N_11978,N_11089);
nor U12050 (N_12050,N_10997,N_10879);
or U12051 (N_12051,N_11991,N_11530);
and U12052 (N_12052,N_11906,N_11102);
and U12053 (N_12053,N_11590,N_11665);
nor U12054 (N_12054,N_11509,N_11831);
nand U12055 (N_12055,N_11986,N_11807);
xnor U12056 (N_12056,N_11231,N_11504);
and U12057 (N_12057,N_10801,N_10845);
nor U12058 (N_12058,N_10949,N_11956);
or U12059 (N_12059,N_11897,N_11491);
xor U12060 (N_12060,N_11578,N_11805);
or U12061 (N_12061,N_11368,N_10825);
or U12062 (N_12062,N_11281,N_11206);
nand U12063 (N_12063,N_11312,N_10896);
xnor U12064 (N_12064,N_10992,N_11155);
xor U12065 (N_12065,N_11835,N_11297);
nand U12066 (N_12066,N_11187,N_11165);
nor U12067 (N_12067,N_11697,N_11760);
nor U12068 (N_12068,N_11461,N_11421);
nand U12069 (N_12069,N_11988,N_11761);
nand U12070 (N_12070,N_11487,N_11324);
and U12071 (N_12071,N_11826,N_11921);
xnor U12072 (N_12072,N_11319,N_11472);
xnor U12073 (N_12073,N_11712,N_11932);
or U12074 (N_12074,N_10988,N_11218);
nor U12075 (N_12075,N_11609,N_11271);
or U12076 (N_12076,N_11030,N_11359);
or U12077 (N_12077,N_10920,N_11959);
nand U12078 (N_12078,N_11985,N_11821);
and U12079 (N_12079,N_11934,N_11485);
xnor U12080 (N_12080,N_10838,N_11732);
xnor U12081 (N_12081,N_11521,N_11253);
and U12082 (N_12082,N_10921,N_11397);
xnor U12083 (N_12083,N_11532,N_11935);
nor U12084 (N_12084,N_11411,N_11576);
nor U12085 (N_12085,N_10916,N_11215);
nor U12086 (N_12086,N_10830,N_11979);
nand U12087 (N_12087,N_11075,N_11642);
nor U12088 (N_12088,N_11892,N_11361);
xor U12089 (N_12089,N_11000,N_11595);
nand U12090 (N_12090,N_11161,N_11635);
nand U12091 (N_12091,N_11302,N_10841);
nand U12092 (N_12092,N_11235,N_11702);
nor U12093 (N_12093,N_11757,N_11949);
xor U12094 (N_12094,N_11028,N_11669);
nand U12095 (N_12095,N_11050,N_10991);
or U12096 (N_12096,N_11382,N_11678);
xnor U12097 (N_12097,N_11437,N_11681);
xor U12098 (N_12098,N_11481,N_11502);
xor U12099 (N_12099,N_11527,N_11575);
or U12100 (N_12100,N_11422,N_11247);
and U12101 (N_12101,N_11864,N_10955);
xor U12102 (N_12102,N_11254,N_11551);
and U12103 (N_12103,N_11730,N_11202);
and U12104 (N_12104,N_11888,N_11074);
nand U12105 (N_12105,N_11789,N_11234);
or U12106 (N_12106,N_11624,N_11911);
and U12107 (N_12107,N_10970,N_11544);
nor U12108 (N_12108,N_11473,N_10800);
and U12109 (N_12109,N_11648,N_11360);
or U12110 (N_12110,N_11651,N_11479);
nand U12111 (N_12111,N_11109,N_11806);
or U12112 (N_12112,N_11138,N_11049);
xnor U12113 (N_12113,N_11374,N_10929);
or U12114 (N_12114,N_11330,N_11684);
or U12115 (N_12115,N_10863,N_11025);
xnor U12116 (N_12116,N_11763,N_11957);
or U12117 (N_12117,N_11597,N_11980);
nor U12118 (N_12118,N_11334,N_11137);
or U12119 (N_12119,N_11777,N_11002);
and U12120 (N_12120,N_11607,N_11917);
and U12121 (N_12121,N_11749,N_11941);
nand U12122 (N_12122,N_10985,N_11615);
nand U12123 (N_12123,N_10835,N_11098);
or U12124 (N_12124,N_10983,N_11387);
xnor U12125 (N_12125,N_11078,N_11948);
nand U12126 (N_12126,N_11315,N_11193);
and U12127 (N_12127,N_11458,N_10904);
or U12128 (N_12128,N_11415,N_11090);
nand U12129 (N_12129,N_10947,N_11240);
or U12130 (N_12130,N_11123,N_11269);
or U12131 (N_12131,N_11589,N_11518);
nand U12132 (N_12132,N_10822,N_11845);
nand U12133 (N_12133,N_11614,N_11799);
nor U12134 (N_12134,N_11713,N_11284);
nor U12135 (N_12135,N_11014,N_11585);
nor U12136 (N_12136,N_11715,N_10831);
nor U12137 (N_12137,N_10876,N_10887);
nand U12138 (N_12138,N_11967,N_11505);
and U12139 (N_12139,N_11796,N_10857);
xnor U12140 (N_12140,N_11900,N_11179);
or U12141 (N_12141,N_10844,N_11363);
nor U12142 (N_12142,N_11738,N_11288);
and U12143 (N_12143,N_11824,N_11866);
xnor U12144 (N_12144,N_11592,N_11346);
or U12145 (N_12145,N_11838,N_11893);
nor U12146 (N_12146,N_10902,N_11785);
nand U12147 (N_12147,N_10961,N_10971);
nand U12148 (N_12148,N_10813,N_11990);
nand U12149 (N_12149,N_11579,N_11158);
or U12150 (N_12150,N_11091,N_11658);
or U12151 (N_12151,N_10895,N_11685);
and U12152 (N_12152,N_10924,N_11813);
nor U12153 (N_12153,N_11655,N_11167);
nand U12154 (N_12154,N_11339,N_11233);
and U12155 (N_12155,N_11797,N_11006);
or U12156 (N_12156,N_11503,N_11350);
nor U12157 (N_12157,N_11084,N_11022);
nand U12158 (N_12158,N_10834,N_11552);
and U12159 (N_12159,N_11881,N_11337);
nand U12160 (N_12160,N_11018,N_11914);
nor U12161 (N_12161,N_11052,N_11770);
nand U12162 (N_12162,N_11392,N_11673);
nand U12163 (N_12163,N_11423,N_11323);
and U12164 (N_12164,N_11268,N_11105);
or U12165 (N_12165,N_11329,N_11211);
and U12166 (N_12166,N_10873,N_11289);
and U12167 (N_12167,N_11163,N_11365);
xor U12168 (N_12168,N_10854,N_10942);
or U12169 (N_12169,N_11471,N_11060);
and U12170 (N_12170,N_11282,N_11550);
and U12171 (N_12171,N_11567,N_11541);
nand U12172 (N_12172,N_11646,N_11465);
and U12173 (N_12173,N_11039,N_11606);
nand U12174 (N_12174,N_11424,N_11901);
or U12175 (N_12175,N_11118,N_10819);
xor U12176 (N_12176,N_10842,N_11822);
nor U12177 (N_12177,N_11410,N_11823);
or U12178 (N_12178,N_11580,N_11404);
and U12179 (N_12179,N_11279,N_11455);
nand U12180 (N_12180,N_11290,N_11559);
and U12181 (N_12181,N_11656,N_10965);
nor U12182 (N_12182,N_11819,N_11619);
nor U12183 (N_12183,N_11840,N_11097);
nand U12184 (N_12184,N_10816,N_11088);
and U12185 (N_12185,N_11644,N_11889);
xnor U12186 (N_12186,N_11445,N_11721);
and U12187 (N_12187,N_11037,N_10972);
nand U12188 (N_12188,N_11470,N_11774);
or U12189 (N_12189,N_11258,N_11507);
nor U12190 (N_12190,N_11308,N_11020);
and U12191 (N_12191,N_11380,N_11364);
nand U12192 (N_12192,N_11629,N_11065);
nor U12193 (N_12193,N_11641,N_11973);
nand U12194 (N_12194,N_11724,N_11320);
nor U12195 (N_12195,N_10932,N_11033);
nor U12196 (N_12196,N_11186,N_10919);
or U12197 (N_12197,N_10928,N_11260);
nand U12198 (N_12198,N_10889,N_11141);
or U12199 (N_12199,N_11908,N_11428);
nand U12200 (N_12200,N_11616,N_10885);
xnor U12201 (N_12201,N_11425,N_11737);
nand U12202 (N_12202,N_11919,N_11871);
nand U12203 (N_12203,N_11023,N_11766);
or U12204 (N_12204,N_11662,N_11096);
nand U12205 (N_12205,N_11981,N_11228);
xor U12206 (N_12206,N_11879,N_11232);
nand U12207 (N_12207,N_11860,N_11322);
or U12208 (N_12208,N_10855,N_11327);
or U12209 (N_12209,N_11468,N_11788);
or U12210 (N_12210,N_11537,N_11524);
and U12211 (N_12211,N_10976,N_11782);
nor U12212 (N_12212,N_11126,N_11384);
nor U12213 (N_12213,N_11056,N_11861);
or U12214 (N_12214,N_10989,N_10881);
nand U12215 (N_12215,N_11783,N_11944);
nor U12216 (N_12216,N_11326,N_11100);
and U12217 (N_12217,N_11227,N_11649);
and U12218 (N_12218,N_11467,N_11809);
and U12219 (N_12219,N_10923,N_11219);
nand U12220 (N_12220,N_11405,N_11677);
nor U12221 (N_12221,N_11107,N_11786);
and U12222 (N_12222,N_11317,N_11790);
xnor U12223 (N_12223,N_11687,N_11064);
nand U12224 (N_12224,N_10912,N_10907);
nand U12225 (N_12225,N_11577,N_11723);
xor U12226 (N_12226,N_11836,N_11605);
nor U12227 (N_12227,N_10951,N_11178);
or U12228 (N_12228,N_11013,N_11693);
nor U12229 (N_12229,N_11795,N_11440);
nand U12230 (N_12230,N_11373,N_11768);
and U12231 (N_12231,N_10866,N_10824);
and U12232 (N_12232,N_11654,N_11403);
xnor U12233 (N_12233,N_10888,N_11928);
nor U12234 (N_12234,N_11196,N_11855);
xor U12235 (N_12235,N_11703,N_11841);
and U12236 (N_12236,N_11451,N_11194);
xnor U12237 (N_12237,N_11676,N_11047);
or U12238 (N_12238,N_11495,N_10868);
nand U12239 (N_12239,N_11094,N_11497);
nand U12240 (N_12240,N_11131,N_10839);
or U12241 (N_12241,N_11195,N_11010);
xnor U12242 (N_12242,N_11753,N_11237);
or U12243 (N_12243,N_11333,N_11983);
and U12244 (N_12244,N_11812,N_11898);
nor U12245 (N_12245,N_11488,N_11553);
and U12246 (N_12246,N_11872,N_11887);
xnor U12247 (N_12247,N_10935,N_10836);
or U12248 (N_12248,N_11275,N_11452);
nand U12249 (N_12249,N_11059,N_10909);
xnor U12250 (N_12250,N_11513,N_10837);
xor U12251 (N_12251,N_10957,N_11453);
nor U12252 (N_12252,N_11966,N_11943);
or U12253 (N_12253,N_11910,N_11854);
nor U12254 (N_12254,N_11787,N_11516);
nand U12255 (N_12255,N_11216,N_10998);
xor U12256 (N_12256,N_11611,N_11115);
xnor U12257 (N_12257,N_11918,N_11870);
xnor U12258 (N_12258,N_10982,N_11417);
or U12259 (N_12259,N_11394,N_10803);
or U12260 (N_12260,N_10886,N_11032);
or U12261 (N_12261,N_11042,N_11972);
nand U12262 (N_12262,N_11894,N_11515);
nand U12263 (N_12263,N_11444,N_11869);
and U12264 (N_12264,N_11244,N_11147);
nand U12265 (N_12265,N_11241,N_11377);
xnor U12266 (N_12266,N_11370,N_11863);
nand U12267 (N_12267,N_11154,N_11775);
xor U12268 (N_12268,N_11344,N_11295);
and U12269 (N_12269,N_11111,N_11175);
xnor U12270 (N_12270,N_11829,N_10807);
and U12271 (N_12271,N_10918,N_11464);
or U12272 (N_12272,N_11803,N_11208);
xnor U12273 (N_12273,N_11717,N_11016);
nor U12274 (N_12274,N_11546,N_11448);
and U12275 (N_12275,N_11933,N_11923);
and U12276 (N_12276,N_11610,N_11070);
nand U12277 (N_12277,N_11976,N_11291);
or U12278 (N_12278,N_11162,N_11401);
nor U12279 (N_12279,N_11180,N_11744);
xnor U12280 (N_12280,N_11613,N_11095);
nor U12281 (N_12281,N_11061,N_11169);
nor U12282 (N_12282,N_11531,N_11735);
nand U12283 (N_12283,N_11238,N_11354);
xor U12284 (N_12284,N_10940,N_11191);
xnor U12285 (N_12285,N_11469,N_10805);
nand U12286 (N_12286,N_11779,N_11017);
and U12287 (N_12287,N_11007,N_11692);
and U12288 (N_12288,N_11939,N_10906);
xor U12289 (N_12289,N_11628,N_10861);
or U12290 (N_12290,N_11151,N_11572);
nand U12291 (N_12291,N_11248,N_10853);
nand U12292 (N_12292,N_10899,N_11045);
and U12293 (N_12293,N_11817,N_11015);
nand U12294 (N_12294,N_11119,N_11771);
nand U12295 (N_12295,N_11875,N_11596);
xor U12296 (N_12296,N_11647,N_10802);
nand U12297 (N_12297,N_10812,N_11252);
nand U12298 (N_12298,N_11709,N_10892);
nor U12299 (N_12299,N_11843,N_11498);
xnor U12300 (N_12300,N_11961,N_10956);
xnor U12301 (N_12301,N_11256,N_11540);
xnor U12302 (N_12302,N_11156,N_11390);
nand U12303 (N_12303,N_11116,N_11255);
nand U12304 (N_12304,N_11818,N_11913);
nand U12305 (N_12305,N_11865,N_11352);
xnor U12306 (N_12306,N_11837,N_11172);
nand U12307 (N_12307,N_11931,N_11144);
and U12308 (N_12308,N_11535,N_11029);
nand U12309 (N_12309,N_11759,N_10821);
xor U12310 (N_12310,N_11272,N_11832);
and U12311 (N_12311,N_11548,N_10898);
or U12312 (N_12312,N_11413,N_10937);
xor U12313 (N_12313,N_10900,N_11372);
or U12314 (N_12314,N_11283,N_11113);
nor U12315 (N_12315,N_11963,N_11904);
and U12316 (N_12316,N_10828,N_11278);
or U12317 (N_12317,N_11634,N_11408);
nor U12318 (N_12318,N_11953,N_11328);
or U12319 (N_12319,N_10850,N_11519);
nor U12320 (N_12320,N_11631,N_11482);
nor U12321 (N_12321,N_11847,N_10973);
xnor U12322 (N_12322,N_10966,N_11710);
nor U12323 (N_12323,N_11299,N_11514);
or U12324 (N_12324,N_11538,N_11087);
nand U12325 (N_12325,N_11314,N_11828);
nand U12326 (N_12326,N_11937,N_11617);
and U12327 (N_12327,N_11564,N_11054);
or U12328 (N_12328,N_10856,N_11466);
nor U12329 (N_12329,N_11349,N_11951);
nor U12330 (N_12330,N_10963,N_11672);
xor U12331 (N_12331,N_11077,N_11478);
nand U12332 (N_12332,N_11925,N_11205);
and U12333 (N_12333,N_11528,N_11250);
nor U12334 (N_12334,N_10974,N_10858);
and U12335 (N_12335,N_10867,N_11731);
nor U12336 (N_12336,N_11024,N_10922);
nor U12337 (N_12337,N_10962,N_11874);
nand U12338 (N_12338,N_11038,N_10877);
xnor U12339 (N_12339,N_11554,N_10908);
xor U12340 (N_12340,N_10934,N_10833);
or U12341 (N_12341,N_10984,N_10883);
nor U12342 (N_12342,N_11849,N_10897);
xor U12343 (N_12343,N_11791,N_11454);
nor U12344 (N_12344,N_11459,N_11036);
nand U12345 (N_12345,N_11099,N_11970);
xnor U12346 (N_12346,N_11762,N_11500);
and U12347 (N_12347,N_11108,N_11414);
and U12348 (N_12348,N_11200,N_11638);
and U12349 (N_12349,N_11398,N_11746);
nand U12350 (N_12350,N_11430,N_10808);
nand U12351 (N_12351,N_10820,N_11776);
or U12352 (N_12352,N_11044,N_10978);
xnor U12353 (N_12353,N_11170,N_10818);
or U12354 (N_12354,N_11434,N_11376);
or U12355 (N_12355,N_10872,N_11708);
nand U12356 (N_12356,N_11602,N_10869);
and U12357 (N_12357,N_11601,N_11345);
or U12358 (N_12358,N_11342,N_10823);
nand U12359 (N_12359,N_10931,N_11433);
xor U12360 (N_12360,N_11124,N_11720);
nand U12361 (N_12361,N_11026,N_10901);
and U12362 (N_12362,N_10811,N_10981);
xnor U12363 (N_12363,N_11489,N_11800);
and U12364 (N_12364,N_11120,N_10860);
nand U12365 (N_12365,N_10926,N_11183);
xnor U12366 (N_12366,N_11306,N_10893);
nand U12367 (N_12367,N_10905,N_11083);
nand U12368 (N_12368,N_10882,N_11714);
nor U12369 (N_12369,N_11555,N_10810);
xnor U12370 (N_12370,N_11522,N_11474);
xnor U12371 (N_12371,N_11603,N_11483);
or U12372 (N_12372,N_11862,N_11701);
nor U12373 (N_12373,N_11391,N_10849);
and U12374 (N_12374,N_11886,N_11794);
nand U12375 (N_12375,N_11004,N_11176);
xnor U12376 (N_12376,N_10999,N_10871);
nand U12377 (N_12377,N_11351,N_11975);
and U12378 (N_12378,N_11133,N_11303);
nand U12379 (N_12379,N_11031,N_11438);
nand U12380 (N_12380,N_11995,N_11493);
xor U12381 (N_12381,N_11441,N_11834);
xor U12382 (N_12382,N_11675,N_11688);
nor U12383 (N_12383,N_11626,N_11386);
xnor U12384 (N_12384,N_10843,N_11436);
xor U12385 (N_12385,N_11103,N_10986);
nor U12386 (N_12386,N_11276,N_11367);
or U12387 (N_12387,N_11292,N_11130);
nor U12388 (N_12388,N_11159,N_11457);
xor U12389 (N_12389,N_11021,N_11820);
nor U12390 (N_12390,N_11798,N_11666);
nor U12391 (N_12391,N_11427,N_11325);
nand U12392 (N_12392,N_11982,N_10948);
nand U12393 (N_12393,N_10884,N_11999);
or U12394 (N_12394,N_11916,N_11492);
nand U12395 (N_12395,N_11593,N_11942);
or U12396 (N_12396,N_11859,N_11517);
nor U12397 (N_12397,N_11657,N_11185);
nor U12398 (N_12398,N_11851,N_11304);
nand U12399 (N_12399,N_11177,N_11946);
xor U12400 (N_12400,N_11767,N_11393);
nand U12401 (N_12401,N_11198,N_11764);
and U12402 (N_12402,N_11418,N_10914);
xor U12403 (N_12403,N_11239,N_10859);
or U12404 (N_12404,N_11378,N_11815);
xnor U12405 (N_12405,N_11680,N_11456);
nand U12406 (N_12406,N_11608,N_11940);
or U12407 (N_12407,N_11112,N_11716);
xnor U12408 (N_12408,N_11752,N_11293);
nand U12409 (N_12409,N_11145,N_10875);
nand U12410 (N_12410,N_11174,N_11523);
xnor U12411 (N_12411,N_11369,N_11072);
nor U12412 (N_12412,N_11591,N_11426);
nand U12413 (N_12413,N_10925,N_11907);
nor U12414 (N_12414,N_10913,N_11484);
nor U12415 (N_12415,N_11539,N_10862);
nand U12416 (N_12416,N_11149,N_11181);
xor U12417 (N_12417,N_11160,N_11612);
nand U12418 (N_12418,N_11696,N_11968);
and U12419 (N_12419,N_11101,N_11740);
nand U12420 (N_12420,N_11079,N_11080);
nor U12421 (N_12421,N_11375,N_10847);
nand U12422 (N_12422,N_11142,N_11435);
and U12423 (N_12423,N_11858,N_11230);
nand U12424 (N_12424,N_11668,N_11811);
or U12425 (N_12425,N_11506,N_11587);
and U12426 (N_12426,N_11584,N_11989);
nor U12427 (N_12427,N_11011,N_11069);
nand U12428 (N_12428,N_11008,N_11135);
nor U12429 (N_12429,N_10891,N_11416);
nand U12430 (N_12430,N_11188,N_11848);
xor U12431 (N_12431,N_11313,N_11557);
xnor U12432 (N_12432,N_11301,N_11573);
xor U12433 (N_12433,N_11563,N_11719);
nor U12434 (N_12434,N_11140,N_11909);
xnor U12435 (N_12435,N_11792,N_11296);
xor U12436 (N_12436,N_11640,N_11743);
nand U12437 (N_12437,N_11543,N_11477);
xor U12438 (N_12438,N_11736,N_11661);
or U12439 (N_12439,N_11772,N_11622);
and U12440 (N_12440,N_10878,N_11545);
or U12441 (N_12441,N_10864,N_11700);
or U12442 (N_12442,N_11667,N_11954);
nor U12443 (N_12443,N_11340,N_11525);
or U12444 (N_12444,N_10987,N_10967);
nand U12445 (N_12445,N_11071,N_11104);
nand U12446 (N_12446,N_11139,N_11076);
xor U12447 (N_12447,N_10815,N_11264);
and U12448 (N_12448,N_11781,N_11085);
xor U12449 (N_12449,N_11896,N_11300);
nand U12450 (N_12450,N_11547,N_11852);
or U12451 (N_12451,N_11969,N_10953);
xnor U12452 (N_12452,N_10945,N_11146);
nand U12453 (N_12453,N_11733,N_11189);
and U12454 (N_12454,N_11062,N_11494);
and U12455 (N_12455,N_10996,N_11136);
or U12456 (N_12456,N_11066,N_11366);
nor U12457 (N_12457,N_11309,N_11132);
nand U12458 (N_12458,N_11987,N_11257);
xnor U12459 (N_12459,N_10806,N_11420);
xnor U12460 (N_12460,N_11110,N_11265);
or U12461 (N_12461,N_11512,N_11962);
nor U12462 (N_12462,N_11383,N_11462);
nor U12463 (N_12463,N_10975,N_11520);
nand U12464 (N_12464,N_10954,N_11210);
nor U12465 (N_12465,N_11486,N_11053);
nor U12466 (N_12466,N_11242,N_11756);
or U12467 (N_12467,N_10959,N_10994);
nand U12468 (N_12468,N_11245,N_11286);
nor U12469 (N_12469,N_11639,N_10938);
and U12470 (N_12470,N_11912,N_11867);
and U12471 (N_12471,N_11439,N_11992);
and U12472 (N_12472,N_11769,N_11880);
nand U12473 (N_12473,N_10832,N_11357);
nor U12474 (N_12474,N_11341,N_10851);
or U12475 (N_12475,N_11853,N_11362);
nor U12476 (N_12476,N_11742,N_11261);
or U12477 (N_12477,N_11645,N_11220);
and U12478 (N_12478,N_11780,N_11722);
nor U12479 (N_12479,N_11463,N_11034);
or U12480 (N_12480,N_11705,N_11226);
or U12481 (N_12481,N_11073,N_11409);
nor U12482 (N_12482,N_11057,N_11223);
and U12483 (N_12483,N_11385,N_11929);
and U12484 (N_12484,N_11092,N_11734);
or U12485 (N_12485,N_11249,N_11993);
nand U12486 (N_12486,N_10852,N_10930);
xnor U12487 (N_12487,N_11192,N_11748);
and U12488 (N_12488,N_10941,N_11343);
or U12489 (N_12489,N_11674,N_11048);
and U12490 (N_12490,N_11630,N_11850);
xor U12491 (N_12491,N_11046,N_11974);
xnor U12492 (N_12492,N_11558,N_11691);
or U12493 (N_12493,N_11984,N_11093);
xnor U12494 (N_12494,N_11755,N_11035);
xor U12495 (N_12495,N_10950,N_11388);
nand U12496 (N_12496,N_11348,N_11389);
nor U12497 (N_12497,N_11833,N_11664);
or U12498 (N_12498,N_11511,N_11920);
or U12499 (N_12499,N_11429,N_11051);
nand U12500 (N_12500,N_11560,N_11331);
or U12501 (N_12501,N_11751,N_11689);
xnor U12502 (N_12502,N_11679,N_11955);
and U12503 (N_12503,N_11332,N_11846);
and U12504 (N_12504,N_11686,N_10979);
and U12505 (N_12505,N_11449,N_11623);
nand U12506 (N_12506,N_11201,N_11706);
xor U12507 (N_12507,N_11229,N_11114);
nand U12508 (N_12508,N_11307,N_11704);
and U12509 (N_12509,N_11844,N_11570);
nor U12510 (N_12510,N_11729,N_10993);
nor U12511 (N_12511,N_11814,N_11793);
nor U12512 (N_12512,N_11480,N_11510);
nand U12513 (N_12513,N_11379,N_11960);
nor U12514 (N_12514,N_11055,N_11890);
nand U12515 (N_12515,N_11694,N_11994);
or U12516 (N_12516,N_11663,N_11650);
and U12517 (N_12517,N_10870,N_11173);
nor U12518 (N_12518,N_11842,N_10840);
or U12519 (N_12519,N_10968,N_10874);
or U12520 (N_12520,N_11659,N_11121);
or U12521 (N_12521,N_11652,N_11335);
nand U12522 (N_12522,N_11671,N_10977);
nor U12523 (N_12523,N_11728,N_11877);
nand U12524 (N_12524,N_11406,N_11549);
nand U12525 (N_12525,N_10903,N_10848);
or U12526 (N_12526,N_11058,N_10817);
nand U12527 (N_12527,N_11266,N_11964);
nor U12528 (N_12528,N_11475,N_11922);
and U12529 (N_12529,N_11225,N_11224);
and U12530 (N_12530,N_11338,N_11311);
nand U12531 (N_12531,N_11903,N_11660);
and U12532 (N_12532,N_11197,N_11012);
xnor U12533 (N_12533,N_11670,N_11690);
and U12534 (N_12534,N_11569,N_11568);
and U12535 (N_12535,N_11043,N_11347);
and U12536 (N_12536,N_11127,N_11965);
or U12537 (N_12537,N_11117,N_11997);
xnor U12538 (N_12538,N_11182,N_11251);
and U12539 (N_12539,N_11653,N_11371);
nand U12540 (N_12540,N_10890,N_10958);
or U12541 (N_12541,N_11199,N_11745);
or U12542 (N_12542,N_11695,N_11636);
nand U12543 (N_12543,N_11171,N_11166);
nor U12544 (N_12544,N_11571,N_11599);
nor U12545 (N_12545,N_11259,N_11952);
and U12546 (N_12546,N_11804,N_11936);
and U12547 (N_12547,N_11203,N_11157);
xor U12548 (N_12548,N_11683,N_11143);
nor U12549 (N_12549,N_10990,N_11938);
and U12550 (N_12550,N_11816,N_11152);
and U12551 (N_12551,N_11400,N_11998);
nand U12552 (N_12552,N_11063,N_10936);
nand U12553 (N_12553,N_11395,N_11773);
xor U12554 (N_12554,N_11129,N_11830);
xnor U12555 (N_12555,N_10910,N_10939);
nand U12556 (N_12556,N_11412,N_10814);
or U12557 (N_12557,N_11529,N_11460);
xor U12558 (N_12558,N_10829,N_11698);
and U12559 (N_12559,N_11882,N_11566);
and U12560 (N_12560,N_11902,N_11277);
or U12561 (N_12561,N_10915,N_11280);
or U12562 (N_12562,N_11556,N_11508);
xnor U12563 (N_12563,N_11153,N_11285);
and U12564 (N_12564,N_11273,N_11565);
and U12565 (N_12565,N_11526,N_11977);
nor U12566 (N_12566,N_11134,N_10809);
nand U12567 (N_12567,N_11316,N_11868);
and U12568 (N_12568,N_11321,N_11009);
nor U12569 (N_12569,N_11583,N_11168);
nor U12570 (N_12570,N_11718,N_11643);
or U12571 (N_12571,N_10980,N_11190);
or U12572 (N_12572,N_11600,N_11802);
and U12573 (N_12573,N_11310,N_11443);
or U12574 (N_12574,N_11431,N_11148);
nor U12575 (N_12575,N_11947,N_11726);
nor U12576 (N_12576,N_11926,N_11432);
and U12577 (N_12577,N_11499,N_11996);
nor U12578 (N_12578,N_11632,N_11106);
or U12579 (N_12579,N_11930,N_10865);
nor U12580 (N_12580,N_11747,N_10944);
and U12581 (N_12581,N_11801,N_11221);
and U12582 (N_12582,N_11122,N_11895);
nand U12583 (N_12583,N_11562,N_11086);
xnor U12584 (N_12584,N_11857,N_11213);
xor U12585 (N_12585,N_11620,N_11739);
nor U12586 (N_12586,N_11125,N_11625);
nor U12587 (N_12587,N_11399,N_11627);
nand U12588 (N_12588,N_11407,N_11041);
and U12589 (N_12589,N_11536,N_11222);
and U12590 (N_12590,N_11899,N_11876);
and U12591 (N_12591,N_11582,N_10846);
or U12592 (N_12592,N_11381,N_11164);
nor U12593 (N_12593,N_11005,N_11574);
and U12594 (N_12594,N_10960,N_11725);
nand U12595 (N_12595,N_11082,N_11067);
nand U12596 (N_12596,N_11699,N_11450);
nor U12597 (N_12597,N_11581,N_11915);
or U12598 (N_12598,N_11001,N_11294);
nor U12599 (N_12599,N_11885,N_11598);
nor U12600 (N_12600,N_11028,N_11912);
xor U12601 (N_12601,N_11528,N_11125);
and U12602 (N_12602,N_10980,N_11633);
nand U12603 (N_12603,N_11202,N_11315);
or U12604 (N_12604,N_11926,N_11864);
or U12605 (N_12605,N_11143,N_10915);
nor U12606 (N_12606,N_11077,N_11090);
and U12607 (N_12607,N_11484,N_11878);
and U12608 (N_12608,N_10917,N_11666);
or U12609 (N_12609,N_11674,N_10883);
or U12610 (N_12610,N_11529,N_11652);
and U12611 (N_12611,N_11507,N_11862);
or U12612 (N_12612,N_11822,N_11000);
nand U12613 (N_12613,N_11942,N_11505);
or U12614 (N_12614,N_11555,N_11815);
nand U12615 (N_12615,N_11558,N_11481);
xnor U12616 (N_12616,N_11814,N_11324);
and U12617 (N_12617,N_11467,N_10888);
xor U12618 (N_12618,N_11614,N_10909);
nor U12619 (N_12619,N_11195,N_11112);
nand U12620 (N_12620,N_11700,N_10987);
or U12621 (N_12621,N_11082,N_11271);
nor U12622 (N_12622,N_11574,N_11207);
or U12623 (N_12623,N_11726,N_11138);
nor U12624 (N_12624,N_10800,N_11994);
nor U12625 (N_12625,N_11520,N_11491);
nand U12626 (N_12626,N_10989,N_11353);
nor U12627 (N_12627,N_11563,N_11227);
nand U12628 (N_12628,N_11778,N_11238);
or U12629 (N_12629,N_11804,N_11568);
and U12630 (N_12630,N_11081,N_11910);
or U12631 (N_12631,N_11049,N_11359);
and U12632 (N_12632,N_10820,N_11589);
or U12633 (N_12633,N_11490,N_11938);
nand U12634 (N_12634,N_11638,N_10908);
and U12635 (N_12635,N_11952,N_11279);
xnor U12636 (N_12636,N_11280,N_11069);
xnor U12637 (N_12637,N_11000,N_11162);
nand U12638 (N_12638,N_11367,N_11305);
xor U12639 (N_12639,N_11537,N_11655);
nor U12640 (N_12640,N_11893,N_11571);
nand U12641 (N_12641,N_11252,N_10832);
and U12642 (N_12642,N_10898,N_11787);
nand U12643 (N_12643,N_11769,N_10971);
or U12644 (N_12644,N_11137,N_11672);
or U12645 (N_12645,N_11625,N_10928);
nor U12646 (N_12646,N_11828,N_11149);
and U12647 (N_12647,N_10879,N_11173);
and U12648 (N_12648,N_10836,N_11177);
nand U12649 (N_12649,N_11971,N_11232);
nand U12650 (N_12650,N_11183,N_11662);
nor U12651 (N_12651,N_11958,N_11872);
nand U12652 (N_12652,N_11234,N_11954);
and U12653 (N_12653,N_11320,N_11025);
xor U12654 (N_12654,N_11972,N_11986);
nor U12655 (N_12655,N_11452,N_10823);
xnor U12656 (N_12656,N_11898,N_11437);
or U12657 (N_12657,N_11789,N_11884);
xnor U12658 (N_12658,N_11990,N_11108);
nand U12659 (N_12659,N_11252,N_11960);
xnor U12660 (N_12660,N_10933,N_11287);
and U12661 (N_12661,N_11144,N_10937);
nand U12662 (N_12662,N_11016,N_11827);
or U12663 (N_12663,N_11297,N_10843);
or U12664 (N_12664,N_10966,N_11140);
nor U12665 (N_12665,N_11715,N_11933);
and U12666 (N_12666,N_11196,N_11598);
xnor U12667 (N_12667,N_11932,N_11218);
and U12668 (N_12668,N_11228,N_11684);
or U12669 (N_12669,N_11481,N_11255);
or U12670 (N_12670,N_11330,N_11767);
and U12671 (N_12671,N_11942,N_11865);
or U12672 (N_12672,N_10803,N_11359);
nor U12673 (N_12673,N_11050,N_10932);
or U12674 (N_12674,N_10929,N_11167);
and U12675 (N_12675,N_11193,N_11101);
or U12676 (N_12676,N_11560,N_11620);
nand U12677 (N_12677,N_11964,N_11251);
nand U12678 (N_12678,N_11951,N_11145);
and U12679 (N_12679,N_11215,N_11745);
or U12680 (N_12680,N_11740,N_11502);
or U12681 (N_12681,N_11382,N_11352);
nor U12682 (N_12682,N_10820,N_11885);
nand U12683 (N_12683,N_11207,N_11904);
nand U12684 (N_12684,N_11965,N_11284);
nor U12685 (N_12685,N_11068,N_11144);
nand U12686 (N_12686,N_11764,N_10826);
xnor U12687 (N_12687,N_10945,N_11986);
and U12688 (N_12688,N_11946,N_11423);
xor U12689 (N_12689,N_11196,N_11191);
nand U12690 (N_12690,N_11018,N_11838);
xor U12691 (N_12691,N_11022,N_10850);
or U12692 (N_12692,N_11079,N_11192);
nand U12693 (N_12693,N_11616,N_11711);
xnor U12694 (N_12694,N_10814,N_11223);
xor U12695 (N_12695,N_10847,N_11291);
nor U12696 (N_12696,N_10943,N_11094);
and U12697 (N_12697,N_11663,N_11021);
xor U12698 (N_12698,N_11330,N_11876);
xnor U12699 (N_12699,N_11559,N_11169);
and U12700 (N_12700,N_11573,N_11162);
and U12701 (N_12701,N_11357,N_11542);
xnor U12702 (N_12702,N_11200,N_11560);
nor U12703 (N_12703,N_11770,N_10869);
nor U12704 (N_12704,N_11300,N_11914);
or U12705 (N_12705,N_11215,N_10865);
nand U12706 (N_12706,N_11640,N_11930);
nand U12707 (N_12707,N_11536,N_11995);
nor U12708 (N_12708,N_11617,N_11673);
and U12709 (N_12709,N_11876,N_11377);
and U12710 (N_12710,N_11067,N_11506);
nand U12711 (N_12711,N_11687,N_11587);
nor U12712 (N_12712,N_11048,N_11961);
xnor U12713 (N_12713,N_11347,N_11356);
and U12714 (N_12714,N_10942,N_11880);
nand U12715 (N_12715,N_11672,N_11973);
nor U12716 (N_12716,N_11171,N_11227);
nor U12717 (N_12717,N_11795,N_11218);
nand U12718 (N_12718,N_11512,N_11565);
xnor U12719 (N_12719,N_11560,N_11983);
and U12720 (N_12720,N_11940,N_10999);
or U12721 (N_12721,N_11773,N_11522);
nor U12722 (N_12722,N_11514,N_11770);
xnor U12723 (N_12723,N_10808,N_11384);
nor U12724 (N_12724,N_10967,N_11473);
nand U12725 (N_12725,N_11504,N_11821);
and U12726 (N_12726,N_11788,N_11244);
nand U12727 (N_12727,N_11671,N_11025);
xnor U12728 (N_12728,N_11142,N_11248);
or U12729 (N_12729,N_11156,N_11478);
nor U12730 (N_12730,N_11474,N_11797);
xor U12731 (N_12731,N_11905,N_11653);
nand U12732 (N_12732,N_11991,N_11566);
nor U12733 (N_12733,N_10909,N_11283);
xnor U12734 (N_12734,N_11595,N_11011);
xnor U12735 (N_12735,N_11127,N_11171);
xnor U12736 (N_12736,N_10829,N_11369);
and U12737 (N_12737,N_11893,N_11549);
nand U12738 (N_12738,N_11421,N_11674);
and U12739 (N_12739,N_10864,N_10828);
xnor U12740 (N_12740,N_10819,N_11988);
and U12741 (N_12741,N_10837,N_11704);
and U12742 (N_12742,N_11623,N_11176);
nand U12743 (N_12743,N_11441,N_11062);
nand U12744 (N_12744,N_11181,N_11345);
nor U12745 (N_12745,N_10808,N_10896);
and U12746 (N_12746,N_11333,N_11907);
and U12747 (N_12747,N_10873,N_10936);
or U12748 (N_12748,N_11206,N_11991);
nor U12749 (N_12749,N_11819,N_11485);
xor U12750 (N_12750,N_11352,N_11644);
xnor U12751 (N_12751,N_10962,N_11716);
and U12752 (N_12752,N_10906,N_11576);
xnor U12753 (N_12753,N_11058,N_11924);
nand U12754 (N_12754,N_10863,N_11325);
and U12755 (N_12755,N_11351,N_11566);
nor U12756 (N_12756,N_11443,N_11323);
and U12757 (N_12757,N_11361,N_10816);
and U12758 (N_12758,N_11398,N_11428);
nor U12759 (N_12759,N_11998,N_11227);
and U12760 (N_12760,N_11634,N_11729);
and U12761 (N_12761,N_10858,N_11190);
nor U12762 (N_12762,N_10987,N_11734);
or U12763 (N_12763,N_11335,N_11718);
xnor U12764 (N_12764,N_11918,N_11151);
xnor U12765 (N_12765,N_11993,N_11443);
xor U12766 (N_12766,N_11637,N_11937);
nor U12767 (N_12767,N_11148,N_11876);
nand U12768 (N_12768,N_11126,N_11051);
nor U12769 (N_12769,N_11697,N_11190);
nand U12770 (N_12770,N_11796,N_11809);
nor U12771 (N_12771,N_11361,N_11814);
and U12772 (N_12772,N_11780,N_11709);
or U12773 (N_12773,N_10884,N_11112);
or U12774 (N_12774,N_11239,N_11367);
and U12775 (N_12775,N_11286,N_11760);
and U12776 (N_12776,N_11975,N_11823);
and U12777 (N_12777,N_11009,N_11489);
nor U12778 (N_12778,N_11653,N_11537);
nand U12779 (N_12779,N_11542,N_11006);
and U12780 (N_12780,N_11403,N_11718);
nand U12781 (N_12781,N_11910,N_11512);
or U12782 (N_12782,N_11384,N_10863);
nand U12783 (N_12783,N_11430,N_10989);
and U12784 (N_12784,N_11506,N_11683);
and U12785 (N_12785,N_11625,N_10869);
and U12786 (N_12786,N_11460,N_11295);
and U12787 (N_12787,N_10920,N_11355);
nor U12788 (N_12788,N_11388,N_11774);
nor U12789 (N_12789,N_11644,N_11897);
or U12790 (N_12790,N_11123,N_11243);
nor U12791 (N_12791,N_11006,N_11651);
nand U12792 (N_12792,N_11859,N_11610);
nand U12793 (N_12793,N_11180,N_11290);
nor U12794 (N_12794,N_11044,N_11921);
nand U12795 (N_12795,N_11054,N_11272);
or U12796 (N_12796,N_11000,N_11803);
nor U12797 (N_12797,N_11097,N_10864);
nor U12798 (N_12798,N_11146,N_11387);
or U12799 (N_12799,N_11560,N_11377);
and U12800 (N_12800,N_11267,N_11356);
xnor U12801 (N_12801,N_11301,N_10814);
nand U12802 (N_12802,N_11556,N_11247);
and U12803 (N_12803,N_11491,N_10914);
nand U12804 (N_12804,N_11046,N_11078);
nor U12805 (N_12805,N_11313,N_11832);
xor U12806 (N_12806,N_10994,N_10836);
or U12807 (N_12807,N_11009,N_11613);
nand U12808 (N_12808,N_11066,N_11329);
and U12809 (N_12809,N_11649,N_10857);
nand U12810 (N_12810,N_11218,N_11263);
or U12811 (N_12811,N_10969,N_11159);
or U12812 (N_12812,N_11123,N_10880);
nand U12813 (N_12813,N_10809,N_11167);
xor U12814 (N_12814,N_11032,N_11634);
or U12815 (N_12815,N_10911,N_11690);
nor U12816 (N_12816,N_10874,N_10916);
or U12817 (N_12817,N_11474,N_11488);
or U12818 (N_12818,N_11483,N_10996);
nor U12819 (N_12819,N_11712,N_11897);
nor U12820 (N_12820,N_11775,N_11960);
nand U12821 (N_12821,N_11329,N_11585);
xnor U12822 (N_12822,N_11124,N_10970);
and U12823 (N_12823,N_11460,N_10819);
xnor U12824 (N_12824,N_11644,N_11610);
xnor U12825 (N_12825,N_11577,N_11515);
nor U12826 (N_12826,N_11458,N_11861);
nor U12827 (N_12827,N_10946,N_11486);
nor U12828 (N_12828,N_11713,N_11214);
and U12829 (N_12829,N_11946,N_10935);
xnor U12830 (N_12830,N_10888,N_11526);
nor U12831 (N_12831,N_11931,N_11800);
or U12832 (N_12832,N_11392,N_11417);
or U12833 (N_12833,N_11506,N_11999);
xor U12834 (N_12834,N_11504,N_10866);
nand U12835 (N_12835,N_11534,N_11932);
xnor U12836 (N_12836,N_10956,N_11709);
nand U12837 (N_12837,N_11424,N_11761);
xnor U12838 (N_12838,N_11293,N_11561);
xor U12839 (N_12839,N_11609,N_11424);
nor U12840 (N_12840,N_11241,N_11038);
and U12841 (N_12841,N_11657,N_10804);
or U12842 (N_12842,N_11762,N_11824);
nor U12843 (N_12843,N_11314,N_11338);
nand U12844 (N_12844,N_11456,N_11369);
nor U12845 (N_12845,N_11230,N_11297);
xnor U12846 (N_12846,N_11973,N_11305);
nor U12847 (N_12847,N_11025,N_11440);
or U12848 (N_12848,N_11592,N_11584);
nand U12849 (N_12849,N_11274,N_11792);
or U12850 (N_12850,N_11732,N_11930);
or U12851 (N_12851,N_11131,N_11844);
nand U12852 (N_12852,N_11221,N_10849);
xor U12853 (N_12853,N_11677,N_11737);
nand U12854 (N_12854,N_10914,N_11301);
and U12855 (N_12855,N_11183,N_11084);
nor U12856 (N_12856,N_11445,N_11152);
or U12857 (N_12857,N_11476,N_11716);
and U12858 (N_12858,N_11691,N_11111);
nand U12859 (N_12859,N_11343,N_11727);
and U12860 (N_12860,N_11009,N_11322);
and U12861 (N_12861,N_11860,N_11265);
or U12862 (N_12862,N_11746,N_11040);
or U12863 (N_12863,N_11105,N_11606);
or U12864 (N_12864,N_11506,N_11315);
and U12865 (N_12865,N_11938,N_11585);
nor U12866 (N_12866,N_11420,N_11355);
nor U12867 (N_12867,N_10923,N_11242);
or U12868 (N_12868,N_10919,N_11679);
nor U12869 (N_12869,N_11032,N_11474);
nand U12870 (N_12870,N_11504,N_11508);
or U12871 (N_12871,N_10877,N_11545);
nand U12872 (N_12872,N_11722,N_11881);
nand U12873 (N_12873,N_11205,N_11324);
nand U12874 (N_12874,N_10840,N_11979);
nand U12875 (N_12875,N_11711,N_11177);
nor U12876 (N_12876,N_11642,N_10888);
and U12877 (N_12877,N_11711,N_11403);
or U12878 (N_12878,N_11444,N_11300);
nor U12879 (N_12879,N_10829,N_11791);
xor U12880 (N_12880,N_11040,N_11754);
or U12881 (N_12881,N_10803,N_11444);
xor U12882 (N_12882,N_11372,N_11409);
or U12883 (N_12883,N_11791,N_11761);
xnor U12884 (N_12884,N_11962,N_11245);
and U12885 (N_12885,N_11722,N_10935);
and U12886 (N_12886,N_11203,N_11681);
xor U12887 (N_12887,N_11690,N_11857);
nor U12888 (N_12888,N_10890,N_11123);
nand U12889 (N_12889,N_11081,N_10996);
nor U12890 (N_12890,N_10949,N_11872);
nor U12891 (N_12891,N_11094,N_11465);
or U12892 (N_12892,N_11696,N_11014);
and U12893 (N_12893,N_11591,N_10847);
xnor U12894 (N_12894,N_11765,N_11499);
nand U12895 (N_12895,N_11238,N_11219);
and U12896 (N_12896,N_11232,N_11629);
and U12897 (N_12897,N_11084,N_11128);
xor U12898 (N_12898,N_11450,N_11882);
xor U12899 (N_12899,N_11948,N_11848);
and U12900 (N_12900,N_11326,N_11786);
and U12901 (N_12901,N_11909,N_11241);
xnor U12902 (N_12902,N_11035,N_10810);
nor U12903 (N_12903,N_11217,N_11857);
or U12904 (N_12904,N_11974,N_11820);
nor U12905 (N_12905,N_11532,N_11689);
xor U12906 (N_12906,N_11139,N_11065);
xnor U12907 (N_12907,N_11449,N_11741);
xnor U12908 (N_12908,N_11912,N_11677);
nor U12909 (N_12909,N_11512,N_11289);
nor U12910 (N_12910,N_11099,N_10935);
and U12911 (N_12911,N_11952,N_11662);
nor U12912 (N_12912,N_11733,N_11604);
or U12913 (N_12913,N_10908,N_11154);
nor U12914 (N_12914,N_10815,N_10842);
xor U12915 (N_12915,N_11929,N_11149);
nor U12916 (N_12916,N_11401,N_11519);
and U12917 (N_12917,N_11052,N_11428);
or U12918 (N_12918,N_11795,N_11943);
xor U12919 (N_12919,N_11339,N_11870);
xnor U12920 (N_12920,N_11436,N_11713);
nand U12921 (N_12921,N_10912,N_11500);
nor U12922 (N_12922,N_10828,N_11990);
and U12923 (N_12923,N_11682,N_10931);
nor U12924 (N_12924,N_11839,N_11608);
nor U12925 (N_12925,N_11368,N_11192);
xor U12926 (N_12926,N_11551,N_11807);
or U12927 (N_12927,N_11009,N_11222);
or U12928 (N_12928,N_11658,N_11957);
nor U12929 (N_12929,N_11260,N_11971);
nand U12930 (N_12930,N_11640,N_10876);
nor U12931 (N_12931,N_11095,N_11604);
nand U12932 (N_12932,N_11879,N_11270);
xnor U12933 (N_12933,N_11057,N_10996);
xor U12934 (N_12934,N_10863,N_11652);
nand U12935 (N_12935,N_11527,N_11278);
nor U12936 (N_12936,N_11265,N_11435);
nand U12937 (N_12937,N_11843,N_11186);
nand U12938 (N_12938,N_11155,N_11249);
nor U12939 (N_12939,N_11565,N_11562);
or U12940 (N_12940,N_11626,N_10812);
and U12941 (N_12941,N_10929,N_10858);
nand U12942 (N_12942,N_11666,N_10968);
nor U12943 (N_12943,N_11544,N_11253);
nand U12944 (N_12944,N_11186,N_11509);
xnor U12945 (N_12945,N_11190,N_11449);
or U12946 (N_12946,N_11871,N_11791);
nand U12947 (N_12947,N_11791,N_11261);
nor U12948 (N_12948,N_11603,N_11433);
nand U12949 (N_12949,N_11800,N_11863);
nand U12950 (N_12950,N_11538,N_11728);
or U12951 (N_12951,N_11608,N_11099);
nor U12952 (N_12952,N_11609,N_11648);
nor U12953 (N_12953,N_11263,N_11807);
xor U12954 (N_12954,N_10971,N_11668);
or U12955 (N_12955,N_11528,N_10876);
and U12956 (N_12956,N_11631,N_11177);
nand U12957 (N_12957,N_10986,N_10948);
nand U12958 (N_12958,N_11032,N_10943);
xnor U12959 (N_12959,N_11612,N_11079);
and U12960 (N_12960,N_11999,N_11681);
or U12961 (N_12961,N_11636,N_10930);
nor U12962 (N_12962,N_11222,N_11461);
or U12963 (N_12963,N_11430,N_11935);
nor U12964 (N_12964,N_11783,N_11299);
or U12965 (N_12965,N_11202,N_11130);
nand U12966 (N_12966,N_10889,N_11776);
and U12967 (N_12967,N_11942,N_11932);
xor U12968 (N_12968,N_11279,N_11527);
xnor U12969 (N_12969,N_11261,N_10891);
or U12970 (N_12970,N_11630,N_10841);
xor U12971 (N_12971,N_10837,N_11577);
or U12972 (N_12972,N_11807,N_11262);
xnor U12973 (N_12973,N_11977,N_11791);
nor U12974 (N_12974,N_11542,N_11132);
and U12975 (N_12975,N_11266,N_11745);
xnor U12976 (N_12976,N_11885,N_11457);
and U12977 (N_12977,N_11415,N_11279);
xor U12978 (N_12978,N_10947,N_11589);
nor U12979 (N_12979,N_11632,N_11521);
nor U12980 (N_12980,N_11248,N_11000);
xor U12981 (N_12981,N_11413,N_11218);
and U12982 (N_12982,N_11167,N_11120);
and U12983 (N_12983,N_11784,N_11524);
nand U12984 (N_12984,N_11982,N_11876);
nor U12985 (N_12985,N_11271,N_11935);
xor U12986 (N_12986,N_11527,N_11702);
xnor U12987 (N_12987,N_10931,N_11083);
and U12988 (N_12988,N_11887,N_11712);
nor U12989 (N_12989,N_11395,N_11630);
nand U12990 (N_12990,N_11068,N_11861);
or U12991 (N_12991,N_11439,N_11434);
or U12992 (N_12992,N_11060,N_11883);
or U12993 (N_12993,N_10847,N_11459);
or U12994 (N_12994,N_11104,N_11536);
xnor U12995 (N_12995,N_11168,N_11442);
nor U12996 (N_12996,N_11913,N_11868);
xor U12997 (N_12997,N_11285,N_11244);
or U12998 (N_12998,N_10951,N_11776);
or U12999 (N_12999,N_11189,N_11934);
and U13000 (N_13000,N_10902,N_11387);
xor U13001 (N_13001,N_11713,N_11147);
and U13002 (N_13002,N_11606,N_10881);
nor U13003 (N_13003,N_10850,N_11221);
nor U13004 (N_13004,N_11052,N_11930);
xnor U13005 (N_13005,N_11249,N_11906);
or U13006 (N_13006,N_11691,N_11956);
and U13007 (N_13007,N_11868,N_10863);
nor U13008 (N_13008,N_10892,N_11563);
or U13009 (N_13009,N_11055,N_11674);
nor U13010 (N_13010,N_10918,N_10880);
nand U13011 (N_13011,N_11667,N_11131);
nand U13012 (N_13012,N_11671,N_11363);
or U13013 (N_13013,N_11013,N_11427);
and U13014 (N_13014,N_11205,N_11190);
nor U13015 (N_13015,N_11508,N_11689);
or U13016 (N_13016,N_11761,N_11617);
nor U13017 (N_13017,N_10811,N_11004);
xnor U13018 (N_13018,N_11652,N_11285);
nand U13019 (N_13019,N_11827,N_11418);
nand U13020 (N_13020,N_11544,N_11943);
xor U13021 (N_13021,N_11933,N_10802);
nand U13022 (N_13022,N_11436,N_11185);
and U13023 (N_13023,N_11006,N_11074);
nand U13024 (N_13024,N_10895,N_11653);
xor U13025 (N_13025,N_11341,N_11811);
nor U13026 (N_13026,N_10915,N_11296);
nand U13027 (N_13027,N_11019,N_11226);
nand U13028 (N_13028,N_11981,N_11799);
nor U13029 (N_13029,N_11789,N_11579);
nand U13030 (N_13030,N_11483,N_11850);
nand U13031 (N_13031,N_11815,N_11904);
or U13032 (N_13032,N_11117,N_11718);
or U13033 (N_13033,N_10915,N_11066);
or U13034 (N_13034,N_10936,N_11511);
xnor U13035 (N_13035,N_11546,N_11516);
and U13036 (N_13036,N_10854,N_10932);
nand U13037 (N_13037,N_10904,N_11134);
or U13038 (N_13038,N_11108,N_11867);
or U13039 (N_13039,N_11151,N_10997);
nor U13040 (N_13040,N_11754,N_11028);
nor U13041 (N_13041,N_10897,N_11737);
nand U13042 (N_13042,N_11716,N_10833);
nor U13043 (N_13043,N_11573,N_11322);
nor U13044 (N_13044,N_11842,N_11851);
xor U13045 (N_13045,N_11790,N_11307);
nor U13046 (N_13046,N_11821,N_10953);
or U13047 (N_13047,N_10835,N_11114);
or U13048 (N_13048,N_11840,N_11093);
xnor U13049 (N_13049,N_10961,N_11103);
nand U13050 (N_13050,N_10859,N_10877);
xor U13051 (N_13051,N_11240,N_11837);
and U13052 (N_13052,N_11396,N_11726);
xor U13053 (N_13053,N_11435,N_10945);
nor U13054 (N_13054,N_10928,N_11059);
nand U13055 (N_13055,N_11891,N_11371);
and U13056 (N_13056,N_11669,N_11096);
and U13057 (N_13057,N_11369,N_11583);
nand U13058 (N_13058,N_11929,N_11799);
xnor U13059 (N_13059,N_11632,N_10880);
nor U13060 (N_13060,N_10987,N_11673);
or U13061 (N_13061,N_11547,N_11457);
xor U13062 (N_13062,N_11583,N_11121);
nand U13063 (N_13063,N_10895,N_10881);
xnor U13064 (N_13064,N_11142,N_11765);
xor U13065 (N_13065,N_11349,N_11909);
nor U13066 (N_13066,N_11855,N_11641);
nand U13067 (N_13067,N_11314,N_11674);
nor U13068 (N_13068,N_11933,N_11429);
or U13069 (N_13069,N_11757,N_11207);
xor U13070 (N_13070,N_10952,N_11097);
nand U13071 (N_13071,N_11489,N_11107);
xor U13072 (N_13072,N_11588,N_11188);
nor U13073 (N_13073,N_11611,N_11358);
nor U13074 (N_13074,N_11923,N_11708);
or U13075 (N_13075,N_11411,N_11049);
nor U13076 (N_13076,N_11397,N_11850);
xor U13077 (N_13077,N_11711,N_11930);
nor U13078 (N_13078,N_10879,N_11487);
nor U13079 (N_13079,N_11949,N_11638);
nor U13080 (N_13080,N_11514,N_10918);
nor U13081 (N_13081,N_11598,N_11576);
nand U13082 (N_13082,N_11208,N_11742);
and U13083 (N_13083,N_11875,N_11265);
xnor U13084 (N_13084,N_11118,N_11228);
and U13085 (N_13085,N_10886,N_11811);
xor U13086 (N_13086,N_11995,N_10894);
xor U13087 (N_13087,N_11009,N_11583);
nor U13088 (N_13088,N_11200,N_10897);
or U13089 (N_13089,N_10888,N_11146);
or U13090 (N_13090,N_10978,N_11852);
xnor U13091 (N_13091,N_11260,N_11499);
xnor U13092 (N_13092,N_11503,N_11697);
and U13093 (N_13093,N_10871,N_11385);
nor U13094 (N_13094,N_10989,N_11373);
nand U13095 (N_13095,N_11582,N_10990);
xor U13096 (N_13096,N_11503,N_11193);
nor U13097 (N_13097,N_11184,N_10935);
nor U13098 (N_13098,N_11751,N_11336);
nand U13099 (N_13099,N_11885,N_11747);
xnor U13100 (N_13100,N_11425,N_11533);
nor U13101 (N_13101,N_10811,N_11837);
nor U13102 (N_13102,N_11679,N_11128);
or U13103 (N_13103,N_11414,N_10942);
xnor U13104 (N_13104,N_11788,N_11679);
nand U13105 (N_13105,N_10897,N_11274);
nand U13106 (N_13106,N_11824,N_11790);
nand U13107 (N_13107,N_11945,N_11571);
nor U13108 (N_13108,N_11854,N_11016);
and U13109 (N_13109,N_11475,N_11304);
nor U13110 (N_13110,N_11757,N_11656);
xor U13111 (N_13111,N_10886,N_10970);
nand U13112 (N_13112,N_11339,N_11198);
nor U13113 (N_13113,N_11950,N_11266);
or U13114 (N_13114,N_11797,N_11888);
nor U13115 (N_13115,N_11939,N_11710);
or U13116 (N_13116,N_11476,N_11481);
nor U13117 (N_13117,N_11213,N_11267);
and U13118 (N_13118,N_11700,N_11828);
and U13119 (N_13119,N_11390,N_11264);
or U13120 (N_13120,N_11838,N_11449);
xnor U13121 (N_13121,N_10878,N_11456);
nand U13122 (N_13122,N_11340,N_10943);
nand U13123 (N_13123,N_11529,N_10922);
and U13124 (N_13124,N_11823,N_11401);
nor U13125 (N_13125,N_11692,N_11673);
xnor U13126 (N_13126,N_11349,N_11779);
and U13127 (N_13127,N_11222,N_11902);
xnor U13128 (N_13128,N_11390,N_11942);
nand U13129 (N_13129,N_11520,N_11216);
and U13130 (N_13130,N_10996,N_10967);
xnor U13131 (N_13131,N_11901,N_11100);
and U13132 (N_13132,N_11804,N_10810);
nand U13133 (N_13133,N_10915,N_11527);
nor U13134 (N_13134,N_11727,N_11151);
and U13135 (N_13135,N_11833,N_11402);
nor U13136 (N_13136,N_11121,N_11542);
and U13137 (N_13137,N_11570,N_11990);
and U13138 (N_13138,N_10939,N_11607);
and U13139 (N_13139,N_11518,N_11321);
nor U13140 (N_13140,N_11166,N_11100);
nand U13141 (N_13141,N_11721,N_11121);
nand U13142 (N_13142,N_11206,N_11412);
nor U13143 (N_13143,N_11193,N_11558);
or U13144 (N_13144,N_10893,N_11504);
nor U13145 (N_13145,N_11187,N_11498);
nor U13146 (N_13146,N_11802,N_10844);
nor U13147 (N_13147,N_11787,N_11278);
or U13148 (N_13148,N_11489,N_11525);
or U13149 (N_13149,N_11496,N_10853);
nor U13150 (N_13150,N_10987,N_11283);
xor U13151 (N_13151,N_10860,N_11900);
or U13152 (N_13152,N_11979,N_10960);
nand U13153 (N_13153,N_11531,N_10949);
and U13154 (N_13154,N_11771,N_11703);
and U13155 (N_13155,N_11445,N_10908);
nand U13156 (N_13156,N_11741,N_11512);
nand U13157 (N_13157,N_11244,N_11595);
and U13158 (N_13158,N_11212,N_11597);
or U13159 (N_13159,N_11834,N_11006);
and U13160 (N_13160,N_10831,N_11287);
nor U13161 (N_13161,N_11671,N_11111);
nor U13162 (N_13162,N_11036,N_11220);
nand U13163 (N_13163,N_11688,N_11433);
or U13164 (N_13164,N_11906,N_10860);
or U13165 (N_13165,N_11590,N_11802);
and U13166 (N_13166,N_10986,N_11809);
or U13167 (N_13167,N_11279,N_11451);
nor U13168 (N_13168,N_11145,N_10860);
nand U13169 (N_13169,N_11870,N_11353);
or U13170 (N_13170,N_11738,N_11952);
nor U13171 (N_13171,N_10810,N_11388);
nor U13172 (N_13172,N_11615,N_11143);
and U13173 (N_13173,N_10883,N_11633);
nand U13174 (N_13174,N_11838,N_11188);
and U13175 (N_13175,N_11242,N_11088);
nand U13176 (N_13176,N_11746,N_11090);
nand U13177 (N_13177,N_11643,N_10984);
nand U13178 (N_13178,N_11086,N_11331);
and U13179 (N_13179,N_11849,N_11534);
xor U13180 (N_13180,N_10815,N_11822);
nand U13181 (N_13181,N_11414,N_11670);
nand U13182 (N_13182,N_11221,N_11132);
and U13183 (N_13183,N_10911,N_11660);
nor U13184 (N_13184,N_11028,N_11149);
xor U13185 (N_13185,N_11729,N_10904);
xnor U13186 (N_13186,N_11554,N_10952);
nand U13187 (N_13187,N_10981,N_10941);
nor U13188 (N_13188,N_11524,N_11956);
or U13189 (N_13189,N_11878,N_11908);
nor U13190 (N_13190,N_11938,N_11956);
xor U13191 (N_13191,N_11036,N_10968);
nand U13192 (N_13192,N_11356,N_11988);
xnor U13193 (N_13193,N_11323,N_11282);
xnor U13194 (N_13194,N_11715,N_11825);
and U13195 (N_13195,N_10852,N_11291);
nor U13196 (N_13196,N_11462,N_10945);
nor U13197 (N_13197,N_11787,N_11984);
nand U13198 (N_13198,N_11795,N_11078);
and U13199 (N_13199,N_11224,N_11630);
nand U13200 (N_13200,N_12934,N_12534);
nand U13201 (N_13201,N_12923,N_13054);
xnor U13202 (N_13202,N_12769,N_12938);
nand U13203 (N_13203,N_12590,N_13187);
or U13204 (N_13204,N_12883,N_12776);
nand U13205 (N_13205,N_12468,N_12234);
nand U13206 (N_13206,N_13057,N_12749);
xnor U13207 (N_13207,N_12339,N_12895);
and U13208 (N_13208,N_13099,N_12162);
xor U13209 (N_13209,N_12289,N_12086);
nor U13210 (N_13210,N_13112,N_13003);
or U13211 (N_13211,N_12295,N_12135);
nor U13212 (N_13212,N_12038,N_13059);
nand U13213 (N_13213,N_12363,N_12493);
and U13214 (N_13214,N_12958,N_12032);
xnor U13215 (N_13215,N_12773,N_13162);
or U13216 (N_13216,N_12492,N_12526);
nand U13217 (N_13217,N_12543,N_12992);
and U13218 (N_13218,N_12571,N_12637);
or U13219 (N_13219,N_12672,N_13036);
or U13220 (N_13220,N_12561,N_12763);
and U13221 (N_13221,N_12939,N_12301);
nor U13222 (N_13222,N_12267,N_12657);
or U13223 (N_13223,N_12971,N_12781);
xnor U13224 (N_13224,N_12897,N_13015);
or U13225 (N_13225,N_13052,N_12400);
and U13226 (N_13226,N_12891,N_12927);
and U13227 (N_13227,N_12761,N_13080);
nand U13228 (N_13228,N_12683,N_13065);
nor U13229 (N_13229,N_12884,N_12321);
and U13230 (N_13230,N_12556,N_13010);
and U13231 (N_13231,N_12152,N_12096);
or U13232 (N_13232,N_12521,N_12831);
nand U13233 (N_13233,N_12870,N_12060);
nand U13234 (N_13234,N_12899,N_12809);
and U13235 (N_13235,N_12257,N_12642);
or U13236 (N_13236,N_13021,N_12106);
xor U13237 (N_13237,N_12089,N_12671);
nor U13238 (N_13238,N_12632,N_13020);
nand U13239 (N_13239,N_13064,N_12649);
or U13240 (N_13240,N_12501,N_12428);
xnor U13241 (N_13241,N_12906,N_12791);
nor U13242 (N_13242,N_12034,N_12709);
nor U13243 (N_13243,N_13082,N_13132);
nand U13244 (N_13244,N_12111,N_12336);
nand U13245 (N_13245,N_12658,N_12546);
and U13246 (N_13246,N_12879,N_12077);
or U13247 (N_13247,N_12115,N_12221);
nand U13248 (N_13248,N_12767,N_13042);
nor U13249 (N_13249,N_12681,N_12080);
nand U13250 (N_13250,N_12237,N_12648);
and U13251 (N_13251,N_12174,N_12202);
nor U13252 (N_13252,N_12548,N_12586);
nand U13253 (N_13253,N_12194,N_12892);
or U13254 (N_13254,N_12005,N_12297);
xor U13255 (N_13255,N_13086,N_12771);
xor U13256 (N_13256,N_12047,N_12838);
or U13257 (N_13257,N_12965,N_12615);
or U13258 (N_13258,N_12944,N_12667);
xor U13259 (N_13259,N_13053,N_12568);
xnor U13260 (N_13260,N_12102,N_12260);
or U13261 (N_13261,N_12969,N_13079);
nor U13262 (N_13262,N_12631,N_13076);
nor U13263 (N_13263,N_12437,N_12139);
xor U13264 (N_13264,N_12088,N_12835);
nor U13265 (N_13265,N_13175,N_13113);
nor U13266 (N_13266,N_12547,N_12097);
and U13267 (N_13267,N_12833,N_12091);
and U13268 (N_13268,N_13012,N_12012);
or U13269 (N_13269,N_12010,N_12433);
or U13270 (N_13270,N_12553,N_13075);
or U13271 (N_13271,N_12601,N_12007);
nor U13272 (N_13272,N_12154,N_12541);
nor U13273 (N_13273,N_12423,N_13135);
and U13274 (N_13274,N_13172,N_13130);
xor U13275 (N_13275,N_13041,N_13094);
and U13276 (N_13276,N_12853,N_12999);
or U13277 (N_13277,N_12677,N_12031);
and U13278 (N_13278,N_12871,N_12737);
nor U13279 (N_13279,N_12936,N_13145);
nand U13280 (N_13280,N_12026,N_12136);
xnor U13281 (N_13281,N_12226,N_13105);
or U13282 (N_13282,N_13091,N_12470);
or U13283 (N_13283,N_12500,N_12227);
or U13284 (N_13284,N_12126,N_12645);
xnor U13285 (N_13285,N_12448,N_12760);
nor U13286 (N_13286,N_13056,N_12846);
nand U13287 (N_13287,N_13136,N_13163);
nor U13288 (N_13288,N_12818,N_12137);
nor U13289 (N_13289,N_13140,N_12516);
nor U13290 (N_13290,N_12744,N_12788);
xnor U13291 (N_13291,N_12133,N_12371);
or U13292 (N_13292,N_12574,N_12701);
or U13293 (N_13293,N_12765,N_13023);
nand U13294 (N_13294,N_12651,N_12241);
or U13295 (N_13295,N_12262,N_13118);
xnor U13296 (N_13296,N_12462,N_12206);
xor U13297 (N_13297,N_12966,N_12807);
nor U13298 (N_13298,N_12424,N_12018);
nor U13299 (N_13299,N_12399,N_12725);
nand U13300 (N_13300,N_12306,N_13039);
nor U13301 (N_13301,N_12367,N_12741);
or U13302 (N_13302,N_13081,N_12244);
and U13303 (N_13303,N_12125,N_12415);
or U13304 (N_13304,N_12357,N_12254);
nor U13305 (N_13305,N_12555,N_12245);
nor U13306 (N_13306,N_12654,N_12092);
xnor U13307 (N_13307,N_12539,N_12011);
xnor U13308 (N_13308,N_12873,N_12929);
nor U13309 (N_13309,N_12180,N_13134);
and U13310 (N_13310,N_12689,N_12759);
and U13311 (N_13311,N_12618,N_12785);
or U13312 (N_13312,N_12281,N_12940);
xor U13313 (N_13313,N_12140,N_12705);
xor U13314 (N_13314,N_12774,N_12607);
nand U13315 (N_13315,N_12663,N_12549);
nand U13316 (N_13316,N_12266,N_12948);
xor U13317 (N_13317,N_12796,N_12953);
or U13318 (N_13318,N_12410,N_12467);
or U13319 (N_13319,N_12650,N_12003);
nor U13320 (N_13320,N_12141,N_13159);
and U13321 (N_13321,N_13106,N_12915);
nor U13322 (N_13322,N_12350,N_12855);
nor U13323 (N_13323,N_13050,N_12469);
or U13324 (N_13324,N_12232,N_12652);
nor U13325 (N_13325,N_12712,N_12507);
nor U13326 (N_13326,N_12129,N_12730);
or U13327 (N_13327,N_12046,N_12413);
or U13328 (N_13328,N_12042,N_12358);
xnor U13329 (N_13329,N_12921,N_12483);
or U13330 (N_13330,N_12517,N_12806);
nand U13331 (N_13331,N_12075,N_12578);
and U13332 (N_13332,N_12457,N_12177);
nor U13333 (N_13333,N_12624,N_12514);
and U13334 (N_13334,N_12017,N_12256);
nor U13335 (N_13335,N_13033,N_13035);
nor U13336 (N_13336,N_12799,N_12678);
nand U13337 (N_13337,N_12387,N_12317);
nand U13338 (N_13338,N_12304,N_12988);
nor U13339 (N_13339,N_12002,N_13100);
and U13340 (N_13340,N_12973,N_12041);
or U13341 (N_13341,N_13150,N_12181);
or U13342 (N_13342,N_12691,N_12124);
or U13343 (N_13343,N_12907,N_12980);
or U13344 (N_13344,N_12821,N_13046);
nand U13345 (N_13345,N_12219,N_12740);
and U13346 (N_13346,N_12770,N_12207);
or U13347 (N_13347,N_13043,N_12646);
nand U13348 (N_13348,N_12629,N_12798);
xnor U13349 (N_13349,N_13142,N_12713);
and U13350 (N_13350,N_12443,N_12560);
xor U13351 (N_13351,N_12979,N_12307);
or U13352 (N_13352,N_12062,N_12865);
and U13353 (N_13353,N_12272,N_12085);
or U13354 (N_13354,N_12867,N_12957);
and U13355 (N_13355,N_12752,N_12402);
and U13356 (N_13356,N_13058,N_12200);
nand U13357 (N_13357,N_12772,N_12377);
or U13358 (N_13358,N_12425,N_12946);
or U13359 (N_13359,N_12349,N_12998);
or U13360 (N_13360,N_12569,N_12783);
xnor U13361 (N_13361,N_12347,N_12967);
and U13362 (N_13362,N_12679,N_12303);
nor U13363 (N_13363,N_13090,N_13152);
nor U13364 (N_13364,N_12758,N_12393);
nor U13365 (N_13365,N_12169,N_12006);
or U13366 (N_13366,N_12587,N_12461);
nand U13367 (N_13367,N_13108,N_12134);
nor U13368 (N_13368,N_12902,N_13151);
nor U13369 (N_13369,N_12119,N_12736);
xnor U13370 (N_13370,N_12072,N_12104);
xor U13371 (N_13371,N_12641,N_12850);
and U13372 (N_13372,N_12887,N_12621);
xor U13373 (N_13373,N_12360,N_12392);
and U13374 (N_13374,N_13154,N_12680);
and U13375 (N_13375,N_12101,N_12635);
nor U13376 (N_13376,N_12354,N_12156);
or U13377 (N_13377,N_12323,N_12438);
nor U13378 (N_13378,N_12112,N_12690);
xnor U13379 (N_13379,N_12160,N_12734);
nor U13380 (N_13380,N_12431,N_12960);
xnor U13381 (N_13381,N_12058,N_12542);
xnor U13382 (N_13382,N_12337,N_13110);
xnor U13383 (N_13383,N_12447,N_12385);
xnor U13384 (N_13384,N_12171,N_12184);
and U13385 (N_13385,N_12030,N_12386);
xnor U13386 (N_13386,N_12913,N_13019);
nor U13387 (N_13387,N_12813,N_12801);
xnor U13388 (N_13388,N_12361,N_12351);
and U13389 (N_13389,N_12217,N_13137);
and U13390 (N_13390,N_12898,N_12095);
or U13391 (N_13391,N_12660,N_12278);
and U13392 (N_13392,N_12828,N_12411);
xor U13393 (N_13393,N_12849,N_12378);
nand U13394 (N_13394,N_12819,N_13068);
and U13395 (N_13395,N_12283,N_13067);
and U13396 (N_13396,N_12930,N_13128);
and U13397 (N_13397,N_12218,N_12094);
nor U13398 (N_13398,N_12346,N_12343);
nand U13399 (N_13399,N_12951,N_12656);
and U13400 (N_13400,N_12751,N_13025);
and U13401 (N_13401,N_12557,N_12665);
or U13402 (N_13402,N_12997,N_12356);
xnor U13403 (N_13403,N_12285,N_12702);
or U13404 (N_13404,N_12318,N_12529);
or U13405 (N_13405,N_12082,N_12620);
and U13406 (N_13406,N_12764,N_12901);
nor U13407 (N_13407,N_13029,N_12750);
or U13408 (N_13408,N_13088,N_13178);
nor U13409 (N_13409,N_12495,N_12747);
and U13410 (N_13410,N_12239,N_12325);
nor U13411 (N_13411,N_12509,N_13084);
nand U13412 (N_13412,N_12427,N_13066);
xnor U13413 (N_13413,N_12859,N_12877);
nor U13414 (N_13414,N_12477,N_12905);
nor U13415 (N_13415,N_12048,N_12612);
nor U13416 (N_13416,N_12839,N_12908);
or U13417 (N_13417,N_12145,N_12826);
and U13418 (N_13418,N_12976,N_13027);
nand U13419 (N_13419,N_12822,N_12151);
and U13420 (N_13420,N_12231,N_12216);
xnor U13421 (N_13421,N_13155,N_12523);
nor U13422 (N_13422,N_12816,N_13095);
or U13423 (N_13423,N_12837,N_13191);
xnor U13424 (N_13424,N_12943,N_12331);
xor U13425 (N_13425,N_12625,N_12888);
or U13426 (N_13426,N_12931,N_12666);
xor U13427 (N_13427,N_12345,N_12059);
and U13428 (N_13428,N_12937,N_12545);
or U13429 (N_13429,N_12117,N_13028);
and U13430 (N_13430,N_12365,N_12220);
nand U13431 (N_13431,N_12506,N_12474);
nand U13432 (N_13432,N_12330,N_12149);
and U13433 (N_13433,N_12579,N_12173);
nor U13434 (N_13434,N_13119,N_12987);
xor U13435 (N_13435,N_12995,N_12172);
nor U13436 (N_13436,N_12634,N_12904);
nand U13437 (N_13437,N_12869,N_13143);
nor U13438 (N_13438,N_13180,N_12175);
xnor U13439 (N_13439,N_13171,N_12098);
xnor U13440 (N_13440,N_12682,N_12315);
nand U13441 (N_13441,N_12808,N_13192);
xor U13442 (N_13442,N_12868,N_12362);
and U13443 (N_13443,N_12616,N_12049);
and U13444 (N_13444,N_12066,N_13070);
nor U13445 (N_13445,N_12955,N_12567);
and U13446 (N_13446,N_13048,N_12903);
nand U13447 (N_13447,N_13026,N_12728);
xnor U13448 (N_13448,N_13147,N_12355);
or U13449 (N_13449,N_12564,N_13123);
nor U13450 (N_13450,N_12592,N_12199);
and U13451 (N_13451,N_12643,N_13120);
or U13452 (N_13452,N_12381,N_12714);
nor U13453 (N_13453,N_12299,N_12950);
and U13454 (N_13454,N_12147,N_12609);
or U13455 (N_13455,N_12659,N_12480);
nor U13456 (N_13456,N_13101,N_13166);
nand U13457 (N_13457,N_12374,N_12669);
or U13458 (N_13458,N_12986,N_12959);
or U13459 (N_13459,N_12212,N_12426);
xnor U13460 (N_13460,N_12670,N_12617);
xor U13461 (N_13461,N_12834,N_12291);
nor U13462 (N_13462,N_12972,N_12107);
or U13463 (N_13463,N_13098,N_12978);
nor U13464 (N_13464,N_12416,N_12604);
or U13465 (N_13465,N_12384,N_12309);
xnor U13466 (N_13466,N_12033,N_12065);
or U13467 (N_13467,N_12341,N_13073);
nand U13468 (N_13468,N_13157,N_12866);
xor U13469 (N_13469,N_12558,N_12409);
or U13470 (N_13470,N_12213,N_12298);
nand U13471 (N_13471,N_12264,N_13072);
and U13472 (N_13472,N_13190,N_12166);
nand U13473 (N_13473,N_12051,N_13022);
or U13474 (N_13474,N_12606,N_12554);
nor U13475 (N_13475,N_12429,N_12893);
and U13476 (N_13476,N_12186,N_13160);
xnor U13477 (N_13477,N_13158,N_12918);
nor U13478 (N_13478,N_12716,N_12013);
xnor U13479 (N_13479,N_12142,N_12746);
nand U13480 (N_13480,N_12926,N_12840);
nand U13481 (N_13481,N_12081,N_12070);
nor U13482 (N_13482,N_12053,N_12146);
and U13483 (N_13483,N_12738,N_12524);
and U13484 (N_13484,N_12722,N_12814);
nand U13485 (N_13485,N_13184,N_12326);
nand U13486 (N_13486,N_12570,N_12848);
or U13487 (N_13487,N_12430,N_13169);
and U13488 (N_13488,N_12511,N_13133);
xnor U13489 (N_13489,N_12074,N_12756);
or U13490 (N_13490,N_12952,N_12475);
nor U13491 (N_13491,N_12185,N_13185);
nand U13492 (N_13492,N_12757,N_13017);
and U13493 (N_13493,N_12021,N_12842);
or U13494 (N_13494,N_12105,N_13179);
nor U13495 (N_13495,N_12496,N_12249);
xor U13496 (N_13496,N_12168,N_12471);
or U13497 (N_13497,N_12472,N_12721);
or U13498 (N_13498,N_13069,N_12627);
nor U13499 (N_13499,N_12768,N_12600);
nor U13500 (N_13500,N_12197,N_12595);
nand U13501 (N_13501,N_12242,N_12205);
nand U13502 (N_13502,N_12403,N_13182);
nand U13503 (N_13503,N_13131,N_12028);
or U13504 (N_13504,N_12300,N_12164);
or U13505 (N_13505,N_12724,N_12333);
nor U13506 (N_13506,N_12261,N_12512);
nand U13507 (N_13507,N_12407,N_12240);
and U13508 (N_13508,N_13038,N_12847);
or U13509 (N_13509,N_12280,N_12694);
and U13510 (N_13510,N_13096,N_12052);
nor U13511 (N_13511,N_12551,N_12845);
or U13512 (N_13512,N_12014,N_12238);
and U13513 (N_13513,N_12263,N_12023);
nor U13514 (N_13514,N_12956,N_12942);
and U13515 (N_13515,N_12661,N_12800);
and U13516 (N_13516,N_12857,N_13093);
nor U13517 (N_13517,N_13032,N_12584);
nor U13518 (N_13518,N_12103,N_12132);
nor U13519 (N_13519,N_12886,N_12449);
or U13520 (N_13520,N_12179,N_12353);
nand U13521 (N_13521,N_13124,N_12476);
and U13522 (N_13522,N_13060,N_12745);
or U13523 (N_13523,N_12882,N_12708);
or U13524 (N_13524,N_12432,N_12451);
or U13525 (N_13525,N_12390,N_12269);
nand U13526 (N_13526,N_12982,N_12639);
nand U13527 (N_13527,N_12489,N_12338);
nor U13528 (N_13528,N_12490,N_13114);
xnor U13529 (N_13529,N_12247,N_12116);
nand U13530 (N_13530,N_12706,N_12209);
xnor U13531 (N_13531,N_12540,N_12633);
or U13532 (N_13532,N_12864,N_12373);
nor U13533 (N_13533,N_13199,N_12552);
nand U13534 (N_13534,N_12910,N_12076);
nor U13535 (N_13535,N_12487,N_12271);
xor U13536 (N_13536,N_12466,N_12463);
xor U13537 (N_13537,N_12335,N_12382);
xnor U13538 (N_13538,N_13002,N_12110);
and U13539 (N_13539,N_12875,N_12854);
xor U13540 (N_13540,N_12019,N_12874);
or U13541 (N_13541,N_12591,N_12368);
and U13542 (N_13542,N_12093,N_12704);
nor U13543 (N_13543,N_12395,N_13121);
or U13544 (N_13544,N_12919,N_12050);
nand U13545 (N_13545,N_13177,N_12990);
nor U13546 (N_13546,N_12118,N_13097);
and U13547 (N_13547,N_12250,N_13161);
nand U13548 (N_13548,N_12962,N_13138);
or U13549 (N_13549,N_12167,N_12025);
nand U13550 (N_13550,N_12210,N_13127);
nand U13551 (N_13551,N_12676,N_12214);
and U13552 (N_13552,N_12153,N_13197);
or U13553 (N_13553,N_13165,N_12790);
or U13554 (N_13554,N_12924,N_12932);
xor U13555 (N_13555,N_12820,N_13198);
and U13556 (N_13556,N_12063,N_12861);
nor U13557 (N_13557,N_13047,N_12204);
and U13558 (N_13558,N_12812,N_12305);
xor U13559 (N_13559,N_12189,N_12876);
xnor U13560 (N_13560,N_12508,N_12778);
nor U13561 (N_13561,N_12150,N_12889);
nor U13562 (N_13562,N_13186,N_12949);
xnor U13563 (N_13563,N_13011,N_13051);
xor U13564 (N_13564,N_12945,N_12538);
nand U13565 (N_13565,N_12376,N_12054);
nand U13566 (N_13566,N_12596,N_12863);
xor U13567 (N_13567,N_12313,N_12941);
xnor U13568 (N_13568,N_12342,N_13168);
and U13569 (N_13569,N_12302,N_12858);
nor U13570 (N_13570,N_12478,N_12223);
or U13571 (N_13571,N_12379,N_12016);
and U13572 (N_13572,N_12131,N_12314);
nand U13573 (N_13573,N_12832,N_12797);
xor U13574 (N_13574,N_13034,N_12372);
nand U13575 (N_13575,N_13122,N_12527);
nor U13576 (N_13576,N_12138,N_12810);
nand U13577 (N_13577,N_12970,N_12515);
nand U13578 (N_13578,N_12726,N_12610);
nor U13579 (N_13579,N_12572,N_13024);
xnor U13580 (N_13580,N_12440,N_12453);
nand U13581 (N_13581,N_12394,N_12310);
or U13582 (N_13582,N_12748,N_12473);
nand U13583 (N_13583,N_12284,N_12636);
xnor U13584 (N_13584,N_12522,N_12559);
xnor U13585 (N_13585,N_12035,N_13156);
nand U13586 (N_13586,N_12603,N_12099);
xnor U13587 (N_13587,N_12920,N_12001);
nor U13588 (N_13588,N_12401,N_12703);
and U13589 (N_13589,N_12287,N_13144);
nor U13590 (N_13590,N_12605,N_13044);
xor U13591 (N_13591,N_12550,N_12794);
or U13592 (N_13592,N_13196,N_12900);
nand U13593 (N_13593,N_12856,N_12359);
and U13594 (N_13594,N_12000,N_12170);
xor U13595 (N_13595,N_12439,N_12114);
or U13596 (N_13596,N_12593,N_12993);
xor U13597 (N_13597,N_12787,N_12322);
or U13598 (N_13598,N_12348,N_12391);
nand U13599 (N_13599,N_12482,N_12532);
and U13600 (N_13600,N_12989,N_12755);
nand U13601 (N_13601,N_12695,N_13173);
or U13602 (N_13602,N_12159,N_12697);
and U13603 (N_13603,N_12922,N_12732);
and U13604 (N_13604,N_12441,N_13030);
xnor U13605 (N_13605,N_12383,N_12843);
or U13606 (N_13606,N_13194,N_12270);
nor U13607 (N_13607,N_12991,N_12530);
nor U13608 (N_13608,N_12743,N_12040);
xnor U13609 (N_13609,N_12528,N_12630);
or U13610 (N_13610,N_12727,N_12155);
and U13611 (N_13611,N_12215,N_12802);
nor U13612 (N_13612,N_13001,N_12045);
nor U13613 (N_13613,N_12113,N_12366);
nor U13614 (N_13614,N_12519,N_12498);
nand U13615 (N_13615,N_12380,N_12450);
xor U13616 (N_13616,N_13103,N_12626);
and U13617 (N_13617,N_12230,N_12811);
and U13618 (N_13618,N_12255,N_12178);
nor U13619 (N_13619,N_12311,N_12319);
xor U13620 (N_13620,N_12688,N_13189);
or U13621 (N_13621,N_12352,N_12055);
nand U13622 (N_13622,N_12334,N_12421);
xnor U13623 (N_13623,N_12279,N_12504);
nor U13624 (N_13624,N_13037,N_12614);
or U13625 (N_13625,N_12418,N_12435);
nor U13626 (N_13626,N_13116,N_12775);
or U13627 (N_13627,N_12917,N_12653);
nand U13628 (N_13628,N_13176,N_12890);
xnor U13629 (N_13629,N_12144,N_12823);
nor U13630 (N_13630,N_13125,N_12968);
and U13631 (N_13631,N_12158,N_12535);
xnor U13632 (N_13632,N_12036,N_12531);
nand U13633 (N_13633,N_12109,N_12222);
or U13634 (N_13634,N_12259,N_12699);
nor U13635 (N_13635,N_12015,N_12286);
xnor U13636 (N_13636,N_12795,N_12452);
xnor U13637 (N_13637,N_12456,N_13117);
xnor U13638 (N_13638,N_12628,N_12533);
and U13639 (N_13639,N_12084,N_12327);
xnor U13640 (N_13640,N_12163,N_12685);
or U13641 (N_13641,N_12536,N_12497);
nor U13642 (N_13642,N_12720,N_12459);
nand U13643 (N_13643,N_12668,N_13102);
and U13644 (N_13644,N_12161,N_13087);
and U13645 (N_13645,N_12925,N_13109);
xnor U13646 (N_13646,N_12947,N_13008);
or U13647 (N_13647,N_12829,N_12061);
nor U13648 (N_13648,N_12885,N_13141);
xor U13649 (N_13649,N_12404,N_12294);
nand U13650 (N_13650,N_12308,N_12397);
nor U13651 (N_13651,N_12235,N_12275);
xnor U13652 (N_13652,N_12251,N_12408);
and U13653 (N_13653,N_12100,N_12292);
and U13654 (N_13654,N_12422,N_12963);
nand U13655 (N_13655,N_12589,N_12090);
nor U13656 (N_13656,N_13049,N_12731);
xor U13657 (N_13657,N_12779,N_12444);
nor U13658 (N_13658,N_12009,N_12252);
and U13659 (N_13659,N_12460,N_12224);
nor U13660 (N_13660,N_12518,N_12577);
or U13661 (N_13661,N_12537,N_12056);
and U13662 (N_13662,N_12370,N_12852);
nor U13663 (N_13663,N_12598,N_12243);
or U13664 (N_13664,N_12793,N_12841);
nand U13665 (N_13665,N_12611,N_12520);
and U13666 (N_13666,N_12068,N_12201);
xor U13667 (N_13667,N_12193,N_12573);
xnor U13668 (N_13668,N_12825,N_12312);
and U13669 (N_13669,N_12187,N_12583);
nor U13670 (N_13670,N_12465,N_12914);
xor U13671 (N_13671,N_13004,N_12580);
xnor U13672 (N_13672,N_12729,N_12268);
nand U13673 (N_13673,N_12710,N_12954);
or U13674 (N_13674,N_12803,N_12157);
and U13675 (N_13675,N_12503,N_12191);
nor U13676 (N_13676,N_12805,N_12486);
nor U13677 (N_13677,N_12563,N_12419);
or U13678 (N_13678,N_12505,N_12662);
xnor U13679 (N_13679,N_12364,N_12484);
or U13680 (N_13680,N_12405,N_12881);
xor U13681 (N_13681,N_12008,N_12324);
or U13682 (N_13682,N_13031,N_12896);
xnor U13683 (N_13683,N_12981,N_12165);
and U13684 (N_13684,N_12575,N_13063);
or U13685 (N_13685,N_12274,N_12183);
nand U13686 (N_13686,N_12647,N_12935);
nand U13687 (N_13687,N_13061,N_13007);
and U13688 (N_13688,N_12622,N_12644);
nand U13689 (N_13689,N_12491,N_12789);
nor U13690 (N_13690,N_12499,N_12108);
and U13691 (N_13691,N_12073,N_12208);
nor U13692 (N_13692,N_12182,N_12933);
nor U13693 (N_13693,N_12087,N_12544);
nand U13694 (N_13694,N_12619,N_12692);
xnor U13695 (N_13695,N_12719,N_12196);
xor U13696 (N_13696,N_13062,N_12762);
or U13697 (N_13697,N_12711,N_12687);
or U13698 (N_13698,N_12417,N_12229);
nor U13699 (N_13699,N_13107,N_12754);
xor U13700 (N_13700,N_12246,N_12277);
nor U13701 (N_13701,N_13040,N_12502);
and U13702 (N_13702,N_12674,N_12985);
xnor U13703 (N_13703,N_12588,N_12320);
nand U13704 (N_13704,N_12375,N_12454);
nor U13705 (N_13705,N_13089,N_12715);
or U13706 (N_13706,N_12067,N_12961);
xnor U13707 (N_13707,N_12817,N_12700);
and U13708 (N_13708,N_12398,N_13083);
and U13709 (N_13709,N_12827,N_12022);
or U13710 (N_13710,N_13006,N_12777);
nand U13711 (N_13711,N_12442,N_12562);
nand U13712 (N_13712,N_12253,N_12123);
xnor U13713 (N_13713,N_12446,N_12860);
xnor U13714 (N_13714,N_12316,N_12057);
and U13715 (N_13715,N_12894,N_12753);
and U13716 (N_13716,N_12911,N_12078);
and U13717 (N_13717,N_12675,N_12344);
or U13718 (N_13718,N_12328,N_12122);
nand U13719 (N_13719,N_12071,N_13104);
or U13720 (N_13720,N_13153,N_12039);
and U13721 (N_13721,N_12878,N_13014);
and U13722 (N_13722,N_13018,N_12148);
and U13723 (N_13723,N_12696,N_12640);
xor U13724 (N_13724,N_12494,N_12766);
xor U13725 (N_13725,N_13000,N_12083);
and U13726 (N_13726,N_12782,N_12412);
or U13727 (N_13727,N_12290,N_12581);
and U13728 (N_13728,N_12739,N_12613);
nor U13729 (N_13729,N_12485,N_12735);
nand U13730 (N_13730,N_12188,N_12044);
xor U13731 (N_13731,N_13009,N_12195);
or U13732 (N_13732,N_12830,N_12996);
nor U13733 (N_13733,N_12190,N_12655);
or U13734 (N_13734,N_12329,N_12233);
nor U13735 (N_13735,N_12248,N_12027);
nor U13736 (N_13736,N_13055,N_12836);
or U13737 (N_13737,N_12608,N_12176);
and U13738 (N_13738,N_12909,N_12597);
xnor U13739 (N_13739,N_12004,N_13149);
nor U13740 (N_13740,N_12983,N_12396);
nor U13741 (N_13741,N_12037,N_12912);
nor U13742 (N_13742,N_12977,N_12121);
nor U13743 (N_13743,N_12707,N_12020);
xor U13744 (N_13744,N_12388,N_12420);
and U13745 (N_13745,N_12198,N_12069);
nand U13746 (N_13746,N_12684,N_12340);
or U13747 (N_13747,N_12203,N_12192);
or U13748 (N_13748,N_12064,N_13045);
nand U13749 (N_13749,N_12804,N_13183);
nor U13750 (N_13750,N_12844,N_12638);
and U13751 (N_13751,N_12582,N_12576);
xor U13752 (N_13752,N_12974,N_12585);
and U13753 (N_13753,N_12293,N_12664);
nand U13754 (N_13754,N_12964,N_12513);
or U13755 (N_13755,N_13078,N_12862);
nand U13756 (N_13756,N_13126,N_12128);
or U13757 (N_13757,N_12332,N_12488);
and U13758 (N_13758,N_12273,N_12686);
and U13759 (N_13759,N_12872,N_12984);
nand U13760 (N_13760,N_13164,N_13005);
xor U13761 (N_13761,N_13074,N_12225);
nand U13762 (N_13762,N_13077,N_12851);
and U13763 (N_13763,N_12717,N_12236);
nor U13764 (N_13764,N_13129,N_12916);
or U13765 (N_13765,N_12120,N_13181);
or U13766 (N_13766,N_12673,N_12565);
xor U13767 (N_13767,N_12276,N_12127);
or U13768 (N_13768,N_12389,N_12594);
and U13769 (N_13769,N_13148,N_13111);
or U13770 (N_13770,N_12481,N_12258);
or U13771 (N_13771,N_12406,N_12445);
or U13772 (N_13772,N_13139,N_12043);
nor U13773 (N_13773,N_12024,N_12436);
xnor U13774 (N_13774,N_13146,N_12928);
nand U13775 (N_13775,N_12228,N_13092);
xor U13776 (N_13776,N_13013,N_12602);
or U13777 (N_13777,N_13174,N_12566);
xnor U13778 (N_13778,N_12288,N_12369);
nor U13779 (N_13779,N_12815,N_13188);
nand U13780 (N_13780,N_12786,N_12143);
nand U13781 (N_13781,N_12994,N_12479);
nand U13782 (N_13782,N_12434,N_12623);
nand U13783 (N_13783,N_12510,N_13071);
xor U13784 (N_13784,N_12780,N_12525);
nand U13785 (N_13785,N_13115,N_12296);
xnor U13786 (N_13786,N_12130,N_12282);
or U13787 (N_13787,N_13016,N_12975);
and U13788 (N_13788,N_12693,N_12265);
or U13789 (N_13789,N_12029,N_12079);
and U13790 (N_13790,N_13167,N_12599);
or U13791 (N_13791,N_12211,N_13085);
xor U13792 (N_13792,N_12784,N_12455);
xor U13793 (N_13793,N_12733,N_12414);
and U13794 (N_13794,N_13170,N_12464);
nand U13795 (N_13795,N_12880,N_12824);
and U13796 (N_13796,N_12718,N_12742);
or U13797 (N_13797,N_12723,N_12792);
nand U13798 (N_13798,N_13193,N_12458);
xnor U13799 (N_13799,N_12698,N_13195);
nor U13800 (N_13800,N_12016,N_12432);
and U13801 (N_13801,N_12169,N_12252);
and U13802 (N_13802,N_12320,N_12766);
nand U13803 (N_13803,N_13185,N_13077);
and U13804 (N_13804,N_13070,N_13155);
nand U13805 (N_13805,N_12373,N_12015);
nand U13806 (N_13806,N_13031,N_12567);
nor U13807 (N_13807,N_12241,N_12886);
and U13808 (N_13808,N_12810,N_13020);
xnor U13809 (N_13809,N_12585,N_12871);
or U13810 (N_13810,N_12449,N_12486);
or U13811 (N_13811,N_12611,N_13186);
nand U13812 (N_13812,N_13045,N_12039);
nand U13813 (N_13813,N_12555,N_12627);
or U13814 (N_13814,N_12273,N_12382);
xnor U13815 (N_13815,N_13013,N_12211);
and U13816 (N_13816,N_12089,N_12244);
nand U13817 (N_13817,N_13032,N_12336);
or U13818 (N_13818,N_12329,N_12312);
xor U13819 (N_13819,N_12525,N_12720);
nor U13820 (N_13820,N_12999,N_12131);
xor U13821 (N_13821,N_12401,N_13077);
nand U13822 (N_13822,N_12865,N_12435);
xor U13823 (N_13823,N_12625,N_12327);
nor U13824 (N_13824,N_12630,N_12204);
and U13825 (N_13825,N_12489,N_12504);
xnor U13826 (N_13826,N_12143,N_12566);
xor U13827 (N_13827,N_12826,N_12226);
xor U13828 (N_13828,N_12728,N_13138);
nor U13829 (N_13829,N_12374,N_12751);
xnor U13830 (N_13830,N_12365,N_12750);
or U13831 (N_13831,N_12590,N_12192);
nand U13832 (N_13832,N_13098,N_12404);
or U13833 (N_13833,N_12626,N_12848);
and U13834 (N_13834,N_13111,N_13073);
xnor U13835 (N_13835,N_12087,N_12319);
or U13836 (N_13836,N_12875,N_12924);
or U13837 (N_13837,N_12002,N_12683);
or U13838 (N_13838,N_12883,N_12816);
xor U13839 (N_13839,N_12184,N_13071);
and U13840 (N_13840,N_12544,N_12941);
or U13841 (N_13841,N_12259,N_12594);
and U13842 (N_13842,N_12822,N_12955);
and U13843 (N_13843,N_13037,N_12510);
nand U13844 (N_13844,N_13053,N_12223);
or U13845 (N_13845,N_12082,N_12314);
nand U13846 (N_13846,N_12585,N_13194);
nor U13847 (N_13847,N_12660,N_12734);
and U13848 (N_13848,N_12998,N_12936);
or U13849 (N_13849,N_12469,N_12498);
nor U13850 (N_13850,N_12964,N_13091);
nor U13851 (N_13851,N_13122,N_13049);
or U13852 (N_13852,N_12418,N_12105);
nor U13853 (N_13853,N_12970,N_12807);
xnor U13854 (N_13854,N_12833,N_12033);
and U13855 (N_13855,N_12118,N_12873);
xor U13856 (N_13856,N_12126,N_12691);
xnor U13857 (N_13857,N_12503,N_13159);
xor U13858 (N_13858,N_12593,N_12251);
nand U13859 (N_13859,N_12951,N_13147);
or U13860 (N_13860,N_13182,N_12474);
and U13861 (N_13861,N_12560,N_12023);
nor U13862 (N_13862,N_12379,N_12462);
nor U13863 (N_13863,N_13157,N_12607);
xor U13864 (N_13864,N_12625,N_12777);
or U13865 (N_13865,N_12985,N_12299);
xor U13866 (N_13866,N_13174,N_12518);
xor U13867 (N_13867,N_12857,N_12791);
xor U13868 (N_13868,N_12170,N_12832);
or U13869 (N_13869,N_12587,N_12758);
nor U13870 (N_13870,N_12694,N_13166);
nor U13871 (N_13871,N_12496,N_12947);
nor U13872 (N_13872,N_12274,N_12956);
nand U13873 (N_13873,N_12121,N_12492);
nor U13874 (N_13874,N_13021,N_12430);
or U13875 (N_13875,N_12102,N_12993);
nand U13876 (N_13876,N_12205,N_12722);
nor U13877 (N_13877,N_12094,N_13116);
xor U13878 (N_13878,N_12922,N_12688);
xor U13879 (N_13879,N_12318,N_12063);
and U13880 (N_13880,N_12746,N_12493);
xor U13881 (N_13881,N_12972,N_12191);
or U13882 (N_13882,N_13148,N_12612);
xnor U13883 (N_13883,N_12366,N_13092);
or U13884 (N_13884,N_12623,N_12535);
and U13885 (N_13885,N_12562,N_12595);
or U13886 (N_13886,N_13098,N_12788);
and U13887 (N_13887,N_12472,N_12477);
xnor U13888 (N_13888,N_12737,N_13093);
nand U13889 (N_13889,N_12635,N_13017);
and U13890 (N_13890,N_12932,N_13016);
nor U13891 (N_13891,N_12701,N_12332);
and U13892 (N_13892,N_12831,N_12870);
or U13893 (N_13893,N_13071,N_12086);
and U13894 (N_13894,N_12685,N_12752);
nand U13895 (N_13895,N_12150,N_12923);
or U13896 (N_13896,N_12409,N_12617);
xnor U13897 (N_13897,N_12579,N_13077);
and U13898 (N_13898,N_12850,N_12439);
and U13899 (N_13899,N_12222,N_12574);
nor U13900 (N_13900,N_12859,N_12735);
xnor U13901 (N_13901,N_12106,N_12568);
or U13902 (N_13902,N_13068,N_13190);
or U13903 (N_13903,N_12865,N_12972);
nand U13904 (N_13904,N_13154,N_12293);
and U13905 (N_13905,N_12476,N_12070);
xnor U13906 (N_13906,N_13045,N_12813);
or U13907 (N_13907,N_13107,N_12684);
and U13908 (N_13908,N_12527,N_12353);
or U13909 (N_13909,N_12491,N_12326);
or U13910 (N_13910,N_12493,N_12908);
nand U13911 (N_13911,N_13109,N_12095);
xnor U13912 (N_13912,N_12154,N_12919);
or U13913 (N_13913,N_13008,N_12685);
xnor U13914 (N_13914,N_12655,N_13085);
nor U13915 (N_13915,N_12730,N_12057);
and U13916 (N_13916,N_12942,N_13193);
nand U13917 (N_13917,N_12259,N_12067);
or U13918 (N_13918,N_12090,N_13070);
xnor U13919 (N_13919,N_12429,N_13167);
nor U13920 (N_13920,N_12300,N_12355);
nor U13921 (N_13921,N_12586,N_12860);
and U13922 (N_13922,N_12905,N_12773);
and U13923 (N_13923,N_12301,N_13182);
or U13924 (N_13924,N_12529,N_13130);
nor U13925 (N_13925,N_12078,N_12857);
nor U13926 (N_13926,N_12131,N_12825);
nor U13927 (N_13927,N_12392,N_12695);
and U13928 (N_13928,N_13140,N_13024);
nand U13929 (N_13929,N_12231,N_12652);
nor U13930 (N_13930,N_12863,N_12057);
nand U13931 (N_13931,N_12462,N_12909);
and U13932 (N_13932,N_12711,N_12339);
xor U13933 (N_13933,N_12948,N_12513);
and U13934 (N_13934,N_12193,N_12882);
xor U13935 (N_13935,N_13012,N_12900);
nand U13936 (N_13936,N_12245,N_12282);
nand U13937 (N_13937,N_12652,N_12303);
and U13938 (N_13938,N_12099,N_12517);
and U13939 (N_13939,N_12353,N_13028);
and U13940 (N_13940,N_12582,N_12091);
and U13941 (N_13941,N_12782,N_12498);
or U13942 (N_13942,N_12811,N_12455);
and U13943 (N_13943,N_12347,N_12519);
or U13944 (N_13944,N_12555,N_12711);
xor U13945 (N_13945,N_12594,N_12984);
nand U13946 (N_13946,N_12902,N_12651);
or U13947 (N_13947,N_12829,N_12565);
or U13948 (N_13948,N_12172,N_12535);
or U13949 (N_13949,N_12334,N_12311);
or U13950 (N_13950,N_12384,N_12291);
nand U13951 (N_13951,N_12796,N_12921);
xor U13952 (N_13952,N_12629,N_12993);
xnor U13953 (N_13953,N_12028,N_12153);
nor U13954 (N_13954,N_12737,N_12741);
xnor U13955 (N_13955,N_12819,N_12935);
xnor U13956 (N_13956,N_12501,N_12208);
nand U13957 (N_13957,N_12367,N_12360);
xor U13958 (N_13958,N_12770,N_12188);
xor U13959 (N_13959,N_12298,N_12948);
and U13960 (N_13960,N_13179,N_12762);
nor U13961 (N_13961,N_13150,N_12920);
nor U13962 (N_13962,N_12046,N_12911);
or U13963 (N_13963,N_12812,N_13155);
nand U13964 (N_13964,N_12375,N_12151);
xnor U13965 (N_13965,N_12096,N_12190);
xnor U13966 (N_13966,N_12770,N_13139);
nor U13967 (N_13967,N_12569,N_12821);
nand U13968 (N_13968,N_12174,N_12758);
xnor U13969 (N_13969,N_12416,N_12341);
and U13970 (N_13970,N_12008,N_12542);
and U13971 (N_13971,N_12644,N_13168);
xnor U13972 (N_13972,N_12305,N_12161);
nor U13973 (N_13973,N_12460,N_12078);
and U13974 (N_13974,N_12825,N_12958);
and U13975 (N_13975,N_12774,N_12781);
xnor U13976 (N_13976,N_13112,N_13195);
xor U13977 (N_13977,N_12359,N_12128);
nor U13978 (N_13978,N_12653,N_12247);
xnor U13979 (N_13979,N_12899,N_13078);
or U13980 (N_13980,N_12691,N_12817);
and U13981 (N_13981,N_12690,N_12416);
nand U13982 (N_13982,N_13152,N_13146);
nor U13983 (N_13983,N_13091,N_12792);
nand U13984 (N_13984,N_12763,N_12727);
nor U13985 (N_13985,N_12777,N_12989);
and U13986 (N_13986,N_12556,N_12201);
nand U13987 (N_13987,N_12113,N_12052);
nor U13988 (N_13988,N_12324,N_12897);
xnor U13989 (N_13989,N_12787,N_12783);
and U13990 (N_13990,N_12721,N_13176);
xnor U13991 (N_13991,N_12993,N_12847);
and U13992 (N_13992,N_12247,N_12471);
nor U13993 (N_13993,N_12833,N_12214);
nand U13994 (N_13994,N_12637,N_13106);
nand U13995 (N_13995,N_12120,N_12644);
nand U13996 (N_13996,N_13090,N_12282);
or U13997 (N_13997,N_13127,N_12205);
or U13998 (N_13998,N_12689,N_13016);
nor U13999 (N_13999,N_12420,N_12373);
nor U14000 (N_14000,N_12283,N_12772);
or U14001 (N_14001,N_12384,N_13070);
xnor U14002 (N_14002,N_12505,N_12203);
xnor U14003 (N_14003,N_12665,N_12360);
nand U14004 (N_14004,N_13136,N_12161);
nor U14005 (N_14005,N_12323,N_12914);
nand U14006 (N_14006,N_12559,N_12697);
nor U14007 (N_14007,N_12136,N_12018);
nor U14008 (N_14008,N_12081,N_12820);
and U14009 (N_14009,N_12683,N_12251);
nand U14010 (N_14010,N_12812,N_12513);
nand U14011 (N_14011,N_12800,N_12614);
nand U14012 (N_14012,N_12573,N_12029);
xnor U14013 (N_14013,N_12281,N_12152);
and U14014 (N_14014,N_12103,N_12859);
and U14015 (N_14015,N_12104,N_12351);
and U14016 (N_14016,N_12454,N_12416);
xnor U14017 (N_14017,N_12627,N_12547);
and U14018 (N_14018,N_12685,N_12837);
nand U14019 (N_14019,N_13070,N_13052);
nand U14020 (N_14020,N_13183,N_12492);
and U14021 (N_14021,N_13162,N_12541);
xnor U14022 (N_14022,N_13162,N_12128);
xor U14023 (N_14023,N_12084,N_12815);
nand U14024 (N_14024,N_12970,N_12086);
nor U14025 (N_14025,N_12255,N_12186);
nand U14026 (N_14026,N_12417,N_12370);
nand U14027 (N_14027,N_12156,N_12685);
nand U14028 (N_14028,N_12348,N_12124);
nor U14029 (N_14029,N_12923,N_12573);
and U14030 (N_14030,N_12515,N_12016);
nand U14031 (N_14031,N_12880,N_12402);
xnor U14032 (N_14032,N_12951,N_12325);
nor U14033 (N_14033,N_12443,N_12679);
xnor U14034 (N_14034,N_12955,N_12363);
nand U14035 (N_14035,N_12250,N_12766);
and U14036 (N_14036,N_12575,N_12578);
nor U14037 (N_14037,N_12078,N_12966);
or U14038 (N_14038,N_12914,N_12771);
xnor U14039 (N_14039,N_12623,N_12108);
or U14040 (N_14040,N_12330,N_12807);
or U14041 (N_14041,N_12977,N_12561);
and U14042 (N_14042,N_12657,N_12678);
and U14043 (N_14043,N_13076,N_12437);
xnor U14044 (N_14044,N_12909,N_12144);
xor U14045 (N_14045,N_13077,N_12463);
and U14046 (N_14046,N_12202,N_12390);
nand U14047 (N_14047,N_12176,N_12555);
nor U14048 (N_14048,N_13166,N_12123);
or U14049 (N_14049,N_13066,N_12682);
and U14050 (N_14050,N_12431,N_12258);
or U14051 (N_14051,N_12323,N_12394);
nand U14052 (N_14052,N_12893,N_12956);
nor U14053 (N_14053,N_12331,N_12535);
nor U14054 (N_14054,N_12612,N_12387);
or U14055 (N_14055,N_12150,N_13123);
nand U14056 (N_14056,N_12670,N_12482);
and U14057 (N_14057,N_12243,N_12319);
or U14058 (N_14058,N_12908,N_12520);
and U14059 (N_14059,N_12137,N_12492);
nand U14060 (N_14060,N_12507,N_12883);
xor U14061 (N_14061,N_12916,N_12755);
xnor U14062 (N_14062,N_12118,N_13155);
nand U14063 (N_14063,N_13004,N_12973);
and U14064 (N_14064,N_12341,N_12030);
and U14065 (N_14065,N_12165,N_12093);
nor U14066 (N_14066,N_12042,N_12166);
and U14067 (N_14067,N_12499,N_12865);
xnor U14068 (N_14068,N_13155,N_12842);
or U14069 (N_14069,N_12224,N_12907);
nand U14070 (N_14070,N_12272,N_12843);
xnor U14071 (N_14071,N_12271,N_13028);
or U14072 (N_14072,N_12592,N_12006);
xnor U14073 (N_14073,N_12770,N_12499);
nand U14074 (N_14074,N_12929,N_13149);
or U14075 (N_14075,N_12546,N_13159);
nand U14076 (N_14076,N_12931,N_12667);
or U14077 (N_14077,N_12933,N_13199);
and U14078 (N_14078,N_12940,N_12913);
or U14079 (N_14079,N_12241,N_12539);
xor U14080 (N_14080,N_12674,N_12369);
nand U14081 (N_14081,N_12531,N_12268);
nand U14082 (N_14082,N_12255,N_12229);
nor U14083 (N_14083,N_12720,N_12539);
nand U14084 (N_14084,N_12155,N_12462);
nor U14085 (N_14085,N_12200,N_12047);
and U14086 (N_14086,N_12843,N_12134);
and U14087 (N_14087,N_12135,N_12304);
nand U14088 (N_14088,N_12968,N_12095);
or U14089 (N_14089,N_12429,N_12223);
and U14090 (N_14090,N_13132,N_12327);
and U14091 (N_14091,N_13147,N_12691);
or U14092 (N_14092,N_12672,N_12951);
or U14093 (N_14093,N_12114,N_12003);
xor U14094 (N_14094,N_12095,N_12261);
nor U14095 (N_14095,N_13003,N_12942);
or U14096 (N_14096,N_12545,N_12598);
and U14097 (N_14097,N_12841,N_12184);
nand U14098 (N_14098,N_12317,N_12103);
xor U14099 (N_14099,N_12459,N_12173);
or U14100 (N_14100,N_12806,N_12257);
nor U14101 (N_14101,N_12735,N_12374);
nor U14102 (N_14102,N_12126,N_12379);
or U14103 (N_14103,N_12232,N_12488);
xor U14104 (N_14104,N_12257,N_12700);
and U14105 (N_14105,N_12793,N_12565);
nand U14106 (N_14106,N_12433,N_12255);
or U14107 (N_14107,N_12857,N_12919);
nor U14108 (N_14108,N_13116,N_12263);
or U14109 (N_14109,N_12996,N_12931);
and U14110 (N_14110,N_12330,N_12832);
and U14111 (N_14111,N_12310,N_12043);
nand U14112 (N_14112,N_12286,N_12179);
nor U14113 (N_14113,N_12049,N_12795);
nand U14114 (N_14114,N_12501,N_12373);
xor U14115 (N_14115,N_12689,N_12484);
or U14116 (N_14116,N_12638,N_12716);
nand U14117 (N_14117,N_12599,N_12452);
and U14118 (N_14118,N_12832,N_13071);
or U14119 (N_14119,N_12885,N_12882);
and U14120 (N_14120,N_13002,N_12724);
or U14121 (N_14121,N_12773,N_12521);
nand U14122 (N_14122,N_12221,N_12535);
or U14123 (N_14123,N_12514,N_12805);
xor U14124 (N_14124,N_12536,N_12409);
and U14125 (N_14125,N_12171,N_12203);
or U14126 (N_14126,N_12462,N_12866);
nor U14127 (N_14127,N_12218,N_12580);
and U14128 (N_14128,N_12071,N_12856);
or U14129 (N_14129,N_12590,N_12034);
and U14130 (N_14130,N_12674,N_12036);
or U14131 (N_14131,N_12099,N_12409);
or U14132 (N_14132,N_13014,N_12866);
or U14133 (N_14133,N_12358,N_13160);
xor U14134 (N_14134,N_12227,N_12959);
or U14135 (N_14135,N_12855,N_12967);
and U14136 (N_14136,N_12028,N_12092);
or U14137 (N_14137,N_12739,N_12805);
nand U14138 (N_14138,N_12806,N_12950);
or U14139 (N_14139,N_12900,N_13072);
or U14140 (N_14140,N_12753,N_12573);
or U14141 (N_14141,N_12623,N_13088);
or U14142 (N_14142,N_12301,N_12380);
or U14143 (N_14143,N_12496,N_12520);
xor U14144 (N_14144,N_13047,N_12319);
or U14145 (N_14145,N_12546,N_12088);
and U14146 (N_14146,N_12971,N_12958);
or U14147 (N_14147,N_12121,N_12700);
or U14148 (N_14148,N_13071,N_12829);
nand U14149 (N_14149,N_12016,N_12610);
nand U14150 (N_14150,N_12689,N_12723);
or U14151 (N_14151,N_12628,N_12712);
and U14152 (N_14152,N_12223,N_12778);
nor U14153 (N_14153,N_13119,N_12098);
nand U14154 (N_14154,N_12431,N_12654);
nand U14155 (N_14155,N_12167,N_12497);
nand U14156 (N_14156,N_12319,N_12975);
or U14157 (N_14157,N_12539,N_13117);
xor U14158 (N_14158,N_12191,N_12409);
nand U14159 (N_14159,N_12297,N_12461);
xor U14160 (N_14160,N_12281,N_12427);
or U14161 (N_14161,N_13026,N_13022);
nor U14162 (N_14162,N_12011,N_13186);
nor U14163 (N_14163,N_12898,N_12241);
and U14164 (N_14164,N_13003,N_12698);
xnor U14165 (N_14165,N_12819,N_12062);
or U14166 (N_14166,N_12053,N_12389);
or U14167 (N_14167,N_13042,N_12451);
and U14168 (N_14168,N_12217,N_12078);
xnor U14169 (N_14169,N_13176,N_12906);
xnor U14170 (N_14170,N_12799,N_12561);
nor U14171 (N_14171,N_12680,N_12356);
xor U14172 (N_14172,N_12815,N_13116);
or U14173 (N_14173,N_12328,N_12319);
nand U14174 (N_14174,N_13191,N_12782);
and U14175 (N_14175,N_13136,N_12075);
or U14176 (N_14176,N_12255,N_12963);
or U14177 (N_14177,N_12290,N_12421);
nand U14178 (N_14178,N_12646,N_12910);
and U14179 (N_14179,N_12314,N_12277);
and U14180 (N_14180,N_12146,N_12291);
or U14181 (N_14181,N_12465,N_12199);
and U14182 (N_14182,N_12973,N_12608);
nand U14183 (N_14183,N_12055,N_13159);
nand U14184 (N_14184,N_12153,N_12950);
nor U14185 (N_14185,N_12939,N_12100);
and U14186 (N_14186,N_12590,N_12972);
and U14187 (N_14187,N_12604,N_12350);
xnor U14188 (N_14188,N_12472,N_12445);
xor U14189 (N_14189,N_12926,N_12685);
nor U14190 (N_14190,N_12925,N_12757);
and U14191 (N_14191,N_13020,N_13183);
xor U14192 (N_14192,N_12757,N_12544);
xnor U14193 (N_14193,N_12905,N_12439);
nor U14194 (N_14194,N_13104,N_12506);
nand U14195 (N_14195,N_12773,N_12253);
xnor U14196 (N_14196,N_12214,N_13112);
nor U14197 (N_14197,N_13084,N_13134);
xnor U14198 (N_14198,N_12352,N_12732);
and U14199 (N_14199,N_12803,N_12146);
and U14200 (N_14200,N_12008,N_12681);
or U14201 (N_14201,N_12568,N_12793);
xor U14202 (N_14202,N_12949,N_12220);
and U14203 (N_14203,N_12195,N_13184);
xor U14204 (N_14204,N_12120,N_12213);
and U14205 (N_14205,N_12663,N_12675);
or U14206 (N_14206,N_12395,N_13174);
xnor U14207 (N_14207,N_12654,N_12368);
and U14208 (N_14208,N_12509,N_12372);
xnor U14209 (N_14209,N_12405,N_12204);
xor U14210 (N_14210,N_12123,N_12772);
xor U14211 (N_14211,N_12487,N_12136);
nor U14212 (N_14212,N_12940,N_12405);
nor U14213 (N_14213,N_12255,N_13022);
nor U14214 (N_14214,N_12023,N_12551);
nand U14215 (N_14215,N_12536,N_12952);
xor U14216 (N_14216,N_12342,N_12758);
and U14217 (N_14217,N_12470,N_12723);
xnor U14218 (N_14218,N_12035,N_12209);
nand U14219 (N_14219,N_13003,N_12204);
nor U14220 (N_14220,N_12108,N_12030);
nand U14221 (N_14221,N_12058,N_12712);
xnor U14222 (N_14222,N_12507,N_12369);
or U14223 (N_14223,N_12887,N_12893);
or U14224 (N_14224,N_12923,N_13084);
nand U14225 (N_14225,N_12093,N_12804);
nor U14226 (N_14226,N_12370,N_12761);
or U14227 (N_14227,N_13078,N_12972);
nand U14228 (N_14228,N_12096,N_13027);
nor U14229 (N_14229,N_13132,N_12438);
nor U14230 (N_14230,N_12715,N_12389);
xnor U14231 (N_14231,N_12215,N_12243);
or U14232 (N_14232,N_13132,N_12629);
and U14233 (N_14233,N_13172,N_12795);
or U14234 (N_14234,N_12744,N_12444);
xor U14235 (N_14235,N_12374,N_12623);
or U14236 (N_14236,N_12401,N_12492);
and U14237 (N_14237,N_12860,N_12095);
or U14238 (N_14238,N_12423,N_12948);
nor U14239 (N_14239,N_12066,N_12074);
xor U14240 (N_14240,N_12279,N_12305);
or U14241 (N_14241,N_12602,N_13048);
nor U14242 (N_14242,N_12287,N_12809);
and U14243 (N_14243,N_12270,N_12049);
and U14244 (N_14244,N_12107,N_13145);
and U14245 (N_14245,N_12270,N_12335);
and U14246 (N_14246,N_12156,N_12908);
xnor U14247 (N_14247,N_12633,N_12555);
and U14248 (N_14248,N_12776,N_12774);
nor U14249 (N_14249,N_13113,N_12520);
xnor U14250 (N_14250,N_12041,N_12671);
xnor U14251 (N_14251,N_12527,N_12292);
nor U14252 (N_14252,N_12278,N_12196);
or U14253 (N_14253,N_12744,N_13190);
or U14254 (N_14254,N_12420,N_12682);
nand U14255 (N_14255,N_12519,N_12359);
or U14256 (N_14256,N_12970,N_13120);
and U14257 (N_14257,N_12181,N_12274);
nand U14258 (N_14258,N_12210,N_12142);
nor U14259 (N_14259,N_12983,N_12652);
or U14260 (N_14260,N_12028,N_13179);
and U14261 (N_14261,N_13080,N_13136);
or U14262 (N_14262,N_12418,N_13069);
nand U14263 (N_14263,N_12443,N_12928);
and U14264 (N_14264,N_12086,N_12271);
nand U14265 (N_14265,N_13021,N_12939);
nand U14266 (N_14266,N_12517,N_12560);
nand U14267 (N_14267,N_12307,N_12077);
xor U14268 (N_14268,N_12109,N_12252);
xor U14269 (N_14269,N_12144,N_12801);
nand U14270 (N_14270,N_12481,N_13185);
and U14271 (N_14271,N_12656,N_12605);
xor U14272 (N_14272,N_12414,N_12820);
or U14273 (N_14273,N_12963,N_12604);
xor U14274 (N_14274,N_12740,N_12788);
nor U14275 (N_14275,N_12816,N_12220);
and U14276 (N_14276,N_13196,N_12275);
nor U14277 (N_14277,N_12538,N_12896);
xor U14278 (N_14278,N_12728,N_13195);
and U14279 (N_14279,N_12625,N_12279);
xnor U14280 (N_14280,N_12498,N_13187);
or U14281 (N_14281,N_13039,N_12424);
nor U14282 (N_14282,N_12455,N_13198);
nor U14283 (N_14283,N_12321,N_12601);
nand U14284 (N_14284,N_13104,N_12556);
nand U14285 (N_14285,N_12317,N_13044);
xor U14286 (N_14286,N_13008,N_12975);
or U14287 (N_14287,N_13127,N_12170);
nor U14288 (N_14288,N_12164,N_12547);
and U14289 (N_14289,N_12830,N_12575);
nor U14290 (N_14290,N_13121,N_13186);
xnor U14291 (N_14291,N_12037,N_12101);
or U14292 (N_14292,N_12824,N_12431);
or U14293 (N_14293,N_12435,N_12931);
or U14294 (N_14294,N_12031,N_12243);
nand U14295 (N_14295,N_12700,N_12612);
nand U14296 (N_14296,N_12533,N_12564);
nand U14297 (N_14297,N_12859,N_12623);
nor U14298 (N_14298,N_12294,N_12925);
or U14299 (N_14299,N_12237,N_12885);
xor U14300 (N_14300,N_12429,N_12127);
or U14301 (N_14301,N_12508,N_12372);
nor U14302 (N_14302,N_12949,N_13027);
and U14303 (N_14303,N_12623,N_12957);
or U14304 (N_14304,N_12649,N_12993);
nand U14305 (N_14305,N_12390,N_12883);
nor U14306 (N_14306,N_12597,N_12715);
nor U14307 (N_14307,N_12107,N_12569);
nor U14308 (N_14308,N_12562,N_13014);
and U14309 (N_14309,N_12286,N_13020);
or U14310 (N_14310,N_12881,N_13010);
nor U14311 (N_14311,N_12688,N_13151);
or U14312 (N_14312,N_12549,N_13137);
and U14313 (N_14313,N_12752,N_12657);
xnor U14314 (N_14314,N_12298,N_12736);
or U14315 (N_14315,N_13039,N_12376);
xnor U14316 (N_14316,N_12707,N_12838);
or U14317 (N_14317,N_12316,N_12772);
or U14318 (N_14318,N_13179,N_12947);
and U14319 (N_14319,N_12289,N_12808);
nand U14320 (N_14320,N_13115,N_12294);
nor U14321 (N_14321,N_12353,N_12577);
nor U14322 (N_14322,N_12229,N_12696);
or U14323 (N_14323,N_12153,N_12971);
xnor U14324 (N_14324,N_12679,N_12797);
nand U14325 (N_14325,N_12626,N_12240);
nand U14326 (N_14326,N_13157,N_12147);
and U14327 (N_14327,N_13027,N_12383);
nand U14328 (N_14328,N_12201,N_13000);
nor U14329 (N_14329,N_13031,N_12623);
and U14330 (N_14330,N_13144,N_12332);
or U14331 (N_14331,N_12507,N_12013);
xnor U14332 (N_14332,N_12007,N_12864);
nand U14333 (N_14333,N_13094,N_12029);
nand U14334 (N_14334,N_12426,N_12861);
and U14335 (N_14335,N_12463,N_13047);
nor U14336 (N_14336,N_12667,N_12525);
and U14337 (N_14337,N_12856,N_12896);
and U14338 (N_14338,N_12613,N_12516);
nor U14339 (N_14339,N_13188,N_12922);
or U14340 (N_14340,N_12082,N_12727);
nand U14341 (N_14341,N_13084,N_12151);
xnor U14342 (N_14342,N_12417,N_13002);
and U14343 (N_14343,N_12811,N_12797);
or U14344 (N_14344,N_12524,N_13025);
nand U14345 (N_14345,N_13178,N_13132);
nor U14346 (N_14346,N_12025,N_12812);
and U14347 (N_14347,N_12777,N_12749);
and U14348 (N_14348,N_12531,N_12465);
nor U14349 (N_14349,N_12682,N_12569);
nand U14350 (N_14350,N_12600,N_12672);
nor U14351 (N_14351,N_13019,N_12866);
nand U14352 (N_14352,N_12438,N_12094);
xnor U14353 (N_14353,N_12630,N_13178);
xnor U14354 (N_14354,N_12574,N_12135);
or U14355 (N_14355,N_12809,N_12686);
or U14356 (N_14356,N_12040,N_12576);
nand U14357 (N_14357,N_12360,N_12144);
or U14358 (N_14358,N_12561,N_12543);
nor U14359 (N_14359,N_12006,N_12857);
xnor U14360 (N_14360,N_12440,N_12276);
xnor U14361 (N_14361,N_12148,N_12445);
or U14362 (N_14362,N_12065,N_12277);
nor U14363 (N_14363,N_12430,N_12032);
and U14364 (N_14364,N_12398,N_12101);
nor U14365 (N_14365,N_13030,N_12721);
nand U14366 (N_14366,N_13111,N_12548);
nand U14367 (N_14367,N_12159,N_12078);
or U14368 (N_14368,N_13053,N_12714);
nand U14369 (N_14369,N_12928,N_12333);
nor U14370 (N_14370,N_12798,N_13076);
nand U14371 (N_14371,N_13187,N_12745);
nand U14372 (N_14372,N_12037,N_12577);
nand U14373 (N_14373,N_12680,N_12737);
or U14374 (N_14374,N_12982,N_12414);
and U14375 (N_14375,N_13086,N_12860);
xnor U14376 (N_14376,N_13049,N_12249);
nor U14377 (N_14377,N_12462,N_12268);
and U14378 (N_14378,N_12064,N_13115);
nor U14379 (N_14379,N_12578,N_12861);
xnor U14380 (N_14380,N_12487,N_12068);
or U14381 (N_14381,N_12177,N_12168);
or U14382 (N_14382,N_13039,N_12724);
or U14383 (N_14383,N_12346,N_12966);
and U14384 (N_14384,N_12488,N_12403);
and U14385 (N_14385,N_12892,N_13179);
and U14386 (N_14386,N_13065,N_12316);
nor U14387 (N_14387,N_12277,N_12140);
and U14388 (N_14388,N_13149,N_13156);
nor U14389 (N_14389,N_13010,N_12236);
and U14390 (N_14390,N_12197,N_12868);
nand U14391 (N_14391,N_12151,N_12386);
xnor U14392 (N_14392,N_12732,N_12226);
and U14393 (N_14393,N_12917,N_12963);
xnor U14394 (N_14394,N_12734,N_12767);
or U14395 (N_14395,N_12554,N_12591);
and U14396 (N_14396,N_12673,N_12425);
or U14397 (N_14397,N_13006,N_12048);
nor U14398 (N_14398,N_12801,N_13140);
xor U14399 (N_14399,N_12747,N_12324);
and U14400 (N_14400,N_14354,N_14153);
nand U14401 (N_14401,N_13340,N_14246);
or U14402 (N_14402,N_13850,N_14387);
nor U14403 (N_14403,N_13822,N_13350);
nor U14404 (N_14404,N_14189,N_13400);
xnor U14405 (N_14405,N_13616,N_14220);
and U14406 (N_14406,N_13663,N_14398);
or U14407 (N_14407,N_14114,N_13221);
xnor U14408 (N_14408,N_14216,N_13450);
nor U14409 (N_14409,N_14340,N_13301);
and U14410 (N_14410,N_14374,N_14310);
or U14411 (N_14411,N_13511,N_13469);
or U14412 (N_14412,N_14273,N_14098);
or U14413 (N_14413,N_13242,N_14380);
and U14414 (N_14414,N_13364,N_14255);
nor U14415 (N_14415,N_13230,N_13273);
nor U14416 (N_14416,N_13676,N_13836);
nand U14417 (N_14417,N_13247,N_13974);
xnor U14418 (N_14418,N_13713,N_13313);
and U14419 (N_14419,N_13913,N_13250);
nor U14420 (N_14420,N_13943,N_14011);
and U14421 (N_14421,N_13216,N_14119);
nand U14422 (N_14422,N_14036,N_14065);
nor U14423 (N_14423,N_13917,N_13710);
and U14424 (N_14424,N_14203,N_14235);
and U14425 (N_14425,N_13463,N_14370);
and U14426 (N_14426,N_13656,N_13842);
and U14427 (N_14427,N_13362,N_14326);
or U14428 (N_14428,N_13757,N_13420);
or U14429 (N_14429,N_13834,N_14236);
or U14430 (N_14430,N_13925,N_13408);
and U14431 (N_14431,N_13893,N_13764);
xnor U14432 (N_14432,N_13363,N_14288);
nand U14433 (N_14433,N_14146,N_13801);
or U14434 (N_14434,N_13983,N_14061);
and U14435 (N_14435,N_13444,N_13415);
and U14436 (N_14436,N_13767,N_13454);
nand U14437 (N_14437,N_13936,N_13532);
xnor U14438 (N_14438,N_13224,N_14297);
nor U14439 (N_14439,N_13765,N_14004);
nor U14440 (N_14440,N_13335,N_13209);
or U14441 (N_14441,N_13251,N_14126);
and U14442 (N_14442,N_13991,N_13686);
nand U14443 (N_14443,N_13266,N_14184);
nand U14444 (N_14444,N_13583,N_14207);
xor U14445 (N_14445,N_13995,N_13785);
or U14446 (N_14446,N_13491,N_13392);
nand U14447 (N_14447,N_13369,N_14032);
or U14448 (N_14448,N_14303,N_13546);
nand U14449 (N_14449,N_14282,N_13239);
nand U14450 (N_14450,N_14197,N_14269);
xnor U14451 (N_14451,N_13732,N_13257);
or U14452 (N_14452,N_13398,N_14222);
xnor U14453 (N_14453,N_13517,N_13254);
xor U14454 (N_14454,N_13915,N_14328);
xor U14455 (N_14455,N_14162,N_13743);
nor U14456 (N_14456,N_13412,N_13904);
or U14457 (N_14457,N_14103,N_13249);
nand U14458 (N_14458,N_13872,N_13289);
and U14459 (N_14459,N_13946,N_13944);
nand U14460 (N_14460,N_14342,N_13481);
xor U14461 (N_14461,N_14049,N_14059);
or U14462 (N_14462,N_14199,N_14042);
or U14463 (N_14463,N_13712,N_14051);
and U14464 (N_14464,N_14225,N_13968);
nand U14465 (N_14465,N_13645,N_13760);
and U14466 (N_14466,N_13378,N_14137);
xnor U14467 (N_14467,N_14035,N_13496);
xor U14468 (N_14468,N_13865,N_14352);
xnor U14469 (N_14469,N_13278,N_13840);
and U14470 (N_14470,N_13506,N_13593);
and U14471 (N_14471,N_14060,N_13222);
xor U14472 (N_14472,N_13344,N_13678);
xnor U14473 (N_14473,N_14177,N_13963);
xor U14474 (N_14474,N_13595,N_14261);
and U14475 (N_14475,N_13423,N_13553);
xor U14476 (N_14476,N_13898,N_13796);
nand U14477 (N_14477,N_14365,N_13885);
and U14478 (N_14478,N_13629,N_14368);
or U14479 (N_14479,N_13581,N_13942);
xor U14480 (N_14480,N_13555,N_14364);
and U14481 (N_14481,N_13895,N_13550);
xor U14482 (N_14482,N_13219,N_14219);
nand U14483 (N_14483,N_13890,N_14022);
xor U14484 (N_14484,N_13787,N_14240);
and U14485 (N_14485,N_14363,N_14373);
nor U14486 (N_14486,N_14280,N_13750);
nor U14487 (N_14487,N_13702,N_14185);
and U14488 (N_14488,N_13486,N_14268);
and U14489 (N_14489,N_13513,N_14030);
and U14490 (N_14490,N_14205,N_13639);
and U14491 (N_14491,N_13468,N_13906);
or U14492 (N_14492,N_14241,N_14144);
and U14493 (N_14493,N_13780,N_14133);
nor U14494 (N_14494,N_13204,N_13390);
xor U14495 (N_14495,N_13373,N_14272);
or U14496 (N_14496,N_13607,N_13673);
or U14497 (N_14497,N_13888,N_14071);
nor U14498 (N_14498,N_13958,N_13499);
nand U14499 (N_14499,N_13954,N_14139);
nor U14500 (N_14500,N_13279,N_13718);
xnor U14501 (N_14501,N_13923,N_13729);
or U14502 (N_14502,N_13397,N_13891);
nand U14503 (N_14503,N_13835,N_13284);
nor U14504 (N_14504,N_13947,N_13706);
or U14505 (N_14505,N_13296,N_13475);
or U14506 (N_14506,N_14377,N_13280);
nand U14507 (N_14507,N_13728,N_13580);
xnor U14508 (N_14508,N_14068,N_13277);
nand U14509 (N_14509,N_13884,N_13263);
nand U14510 (N_14510,N_14003,N_13874);
xnor U14511 (N_14511,N_13986,N_13805);
and U14512 (N_14512,N_13297,N_13766);
or U14513 (N_14513,N_13514,N_13721);
nor U14514 (N_14514,N_13304,N_14121);
xor U14515 (N_14515,N_13603,N_13281);
nand U14516 (N_14516,N_14001,N_14249);
nor U14517 (N_14517,N_14350,N_13451);
and U14518 (N_14518,N_13815,N_14157);
and U14519 (N_14519,N_13524,N_13324);
or U14520 (N_14520,N_13326,N_14007);
nand U14521 (N_14521,N_13414,N_13554);
and U14522 (N_14522,N_13316,N_13405);
xnor U14523 (N_14523,N_13336,N_13535);
nand U14524 (N_14524,N_14290,N_14025);
xor U14525 (N_14525,N_13588,N_14016);
xnor U14526 (N_14526,N_14090,N_13867);
xor U14527 (N_14527,N_13569,N_13606);
nor U14528 (N_14528,N_14265,N_14078);
and U14529 (N_14529,N_13330,N_13669);
and U14530 (N_14530,N_13537,N_13352);
nor U14531 (N_14531,N_13794,N_14124);
nor U14532 (N_14532,N_13618,N_14172);
xor U14533 (N_14533,N_14117,N_13283);
and U14534 (N_14534,N_13303,N_13410);
nand U14535 (N_14535,N_13223,N_13527);
nor U14536 (N_14536,N_13996,N_13459);
nand U14537 (N_14537,N_13498,N_13520);
and U14538 (N_14538,N_13759,N_13471);
or U14539 (N_14539,N_13816,N_13628);
or U14540 (N_14540,N_14263,N_13594);
and U14541 (N_14541,N_14056,N_14169);
and U14542 (N_14542,N_14191,N_13461);
xor U14543 (N_14543,N_13228,N_14317);
nor U14544 (N_14544,N_13894,N_14385);
xnor U14545 (N_14545,N_14034,N_14170);
xnor U14546 (N_14546,N_14285,N_13417);
nor U14547 (N_14547,N_13876,N_13708);
xor U14548 (N_14548,N_13741,N_13206);
and U14549 (N_14549,N_13311,N_13315);
nand U14550 (N_14550,N_13253,N_13208);
and U14551 (N_14551,N_14047,N_14311);
nand U14552 (N_14552,N_13847,N_13981);
xnor U14553 (N_14553,N_13726,N_13902);
and U14554 (N_14554,N_14353,N_14231);
and U14555 (N_14555,N_13979,N_14064);
or U14556 (N_14556,N_13275,N_14344);
xnor U14557 (N_14557,N_13436,N_14307);
nor U14558 (N_14558,N_13666,N_13771);
and U14559 (N_14559,N_14073,N_13689);
nor U14560 (N_14560,N_14021,N_14101);
nor U14561 (N_14561,N_13552,N_14088);
or U14562 (N_14562,N_14391,N_14204);
xor U14563 (N_14563,N_13659,N_13798);
nand U14564 (N_14564,N_13998,N_13651);
or U14565 (N_14565,N_14319,N_13202);
or U14566 (N_14566,N_14258,N_13619);
or U14567 (N_14567,N_13503,N_13934);
and U14568 (N_14568,N_14077,N_14291);
and U14569 (N_14569,N_13859,N_13755);
or U14570 (N_14570,N_13671,N_14361);
nand U14571 (N_14571,N_14395,N_13259);
and U14572 (N_14572,N_14165,N_13952);
nor U14573 (N_14573,N_13869,N_14388);
nand U14574 (N_14574,N_14367,N_13921);
and U14575 (N_14575,N_13971,N_13899);
xnor U14576 (N_14576,N_13641,N_13292);
nand U14577 (N_14577,N_14322,N_14394);
nor U14578 (N_14578,N_14181,N_13927);
or U14579 (N_14579,N_14239,N_14053);
nand U14580 (N_14580,N_13544,N_13379);
xor U14581 (N_14581,N_13807,N_13654);
and U14582 (N_14582,N_13851,N_14372);
nor U14583 (N_14583,N_14151,N_13573);
xor U14584 (N_14584,N_13497,N_13551);
and U14585 (N_14585,N_14331,N_14332);
and U14586 (N_14586,N_14253,N_13839);
xor U14587 (N_14587,N_13244,N_14194);
or U14588 (N_14588,N_13310,N_14337);
and U14589 (N_14589,N_13227,N_13411);
or U14590 (N_14590,N_13285,N_14338);
xnor U14591 (N_14591,N_13533,N_14366);
nor U14592 (N_14592,N_13539,N_14018);
nand U14593 (N_14593,N_13882,N_13272);
or U14594 (N_14594,N_13799,N_14070);
nor U14595 (N_14595,N_13960,N_13243);
nand U14596 (N_14596,N_13245,N_13852);
nand U14597 (N_14597,N_13416,N_13812);
or U14598 (N_14598,N_13967,N_13664);
nor U14599 (N_14599,N_13866,N_14134);
nand U14600 (N_14600,N_13762,N_13620);
nor U14601 (N_14601,N_14218,N_13791);
nor U14602 (N_14602,N_13797,N_13825);
or U14603 (N_14603,N_13441,N_13282);
nor U14604 (N_14604,N_13783,N_14242);
and U14605 (N_14605,N_13359,N_14214);
and U14606 (N_14606,N_13523,N_13268);
or U14607 (N_14607,N_13776,N_13349);
nor U14608 (N_14608,N_14234,N_13644);
xnor U14609 (N_14609,N_13231,N_13492);
nand U14610 (N_14610,N_13993,N_13515);
nor U14611 (N_14611,N_13670,N_13332);
or U14612 (N_14612,N_14397,N_13413);
xor U14613 (N_14613,N_13932,N_13745);
nor U14614 (N_14614,N_13845,N_13374);
nor U14615 (N_14615,N_13596,N_13687);
xnor U14616 (N_14616,N_13388,N_13333);
and U14617 (N_14617,N_14382,N_13833);
nor U14618 (N_14618,N_13919,N_13218);
xnor U14619 (N_14619,N_14024,N_14150);
and U14620 (N_14620,N_13201,N_13601);
or U14621 (N_14621,N_14336,N_14399);
nor U14622 (N_14622,N_13696,N_14250);
and U14623 (N_14623,N_13602,N_13519);
nand U14624 (N_14624,N_13474,N_14043);
xnor U14625 (N_14625,N_13864,N_14277);
and U14626 (N_14626,N_13810,N_13987);
xor U14627 (N_14627,N_14289,N_13467);
nor U14628 (N_14628,N_13945,N_13627);
and U14629 (N_14629,N_13466,N_13905);
nor U14630 (N_14630,N_13425,N_14276);
nand U14631 (N_14631,N_14356,N_13652);
and U14632 (N_14632,N_13817,N_14045);
and U14633 (N_14633,N_13574,N_13590);
xnor U14634 (N_14634,N_13896,N_14046);
and U14635 (N_14635,N_13742,N_13751);
nand U14636 (N_14636,N_13873,N_13912);
nor U14637 (N_14637,N_13961,N_14301);
nand U14638 (N_14638,N_13556,N_13858);
or U14639 (N_14639,N_14039,N_13341);
nor U14640 (N_14640,N_13453,N_13964);
or U14641 (N_14641,N_13427,N_14318);
nor U14642 (N_14642,N_13226,N_13465);
and U14643 (N_14643,N_13494,N_13440);
nor U14644 (N_14644,N_13938,N_13868);
and U14645 (N_14645,N_13455,N_14211);
xor U14646 (N_14646,N_13542,N_13365);
nand U14647 (N_14647,N_14105,N_13727);
or U14648 (N_14648,N_13831,N_13768);
nand U14649 (N_14649,N_14052,N_14093);
or U14650 (N_14650,N_14306,N_13897);
nor U14651 (N_14651,N_14346,N_13462);
xor U14652 (N_14652,N_14248,N_13337);
nand U14653 (N_14653,N_14089,N_13531);
and U14654 (N_14654,N_14058,N_13225);
nor U14655 (N_14655,N_13608,N_13811);
and U14656 (N_14656,N_14100,N_14257);
nand U14657 (N_14657,N_13770,N_13740);
and U14658 (N_14658,N_13953,N_13737);
xor U14659 (N_14659,N_13857,N_13504);
xnor U14660 (N_14660,N_14274,N_13695);
and U14661 (N_14661,N_13381,N_14014);
or U14662 (N_14662,N_14267,N_14102);
and U14663 (N_14663,N_14108,N_13375);
xnor U14664 (N_14664,N_13447,N_13838);
and U14665 (N_14665,N_13931,N_14213);
nand U14666 (N_14666,N_14069,N_14167);
xor U14667 (N_14667,N_14174,N_13819);
nor U14668 (N_14668,N_13661,N_14123);
or U14669 (N_14669,N_13924,N_14037);
and U14670 (N_14670,N_13256,N_13903);
or U14671 (N_14671,N_13353,N_14321);
nor U14672 (N_14672,N_14115,N_13562);
and U14673 (N_14673,N_14233,N_13738);
nand U14674 (N_14674,N_13725,N_14279);
xnor U14675 (N_14675,N_13386,N_14099);
xnor U14676 (N_14676,N_13308,N_13688);
nand U14677 (N_14677,N_13980,N_14147);
nand U14678 (N_14678,N_13844,N_14357);
nor U14679 (N_14679,N_14057,N_14330);
nand U14680 (N_14680,N_13338,N_13643);
and U14681 (N_14681,N_13662,N_13646);
xnor U14682 (N_14682,N_13978,N_13262);
xnor U14683 (N_14683,N_13401,N_14232);
xnor U14684 (N_14684,N_13269,N_14343);
nand U14685 (N_14685,N_14296,N_13294);
xnor U14686 (N_14686,N_13647,N_13351);
nor U14687 (N_14687,N_13684,N_13545);
xor U14688 (N_14688,N_14080,N_14187);
nand U14689 (N_14689,N_14006,N_13999);
nor U14690 (N_14690,N_13637,N_13667);
and U14691 (N_14691,N_13823,N_14193);
or U14692 (N_14692,N_14384,N_13252);
or U14693 (N_14693,N_14378,N_14148);
nand U14694 (N_14694,N_13992,N_14128);
nand U14695 (N_14695,N_13437,N_13970);
or U14696 (N_14696,N_14221,N_14190);
or U14697 (N_14697,N_13638,N_13265);
or U14698 (N_14698,N_13754,N_14142);
or U14699 (N_14699,N_13212,N_14325);
xor U14700 (N_14700,N_13248,N_13355);
and U14701 (N_14701,N_13325,N_14324);
nor U14702 (N_14702,N_14329,N_13419);
nand U14703 (N_14703,N_14215,N_14302);
or U14704 (N_14704,N_13529,N_13989);
or U14705 (N_14705,N_13880,N_13579);
and U14706 (N_14706,N_14085,N_13238);
and U14707 (N_14707,N_13937,N_13792);
nor U14708 (N_14708,N_14202,N_13356);
nand U14709 (N_14709,N_14125,N_13472);
or U14710 (N_14710,N_13557,N_13298);
or U14711 (N_14711,N_14050,N_14333);
and U14712 (N_14712,N_14314,N_13477);
nor U14713 (N_14713,N_13846,N_13217);
nand U14714 (N_14714,N_14109,N_14351);
xor U14715 (N_14715,N_13559,N_13690);
or U14716 (N_14716,N_14075,N_13331);
and U14717 (N_14717,N_14129,N_13458);
nand U14718 (N_14718,N_13784,N_13853);
nand U14719 (N_14719,N_13343,N_14178);
nand U14720 (N_14720,N_13672,N_13907);
nand U14721 (N_14721,N_13319,N_13399);
and U14722 (N_14722,N_13449,N_13305);
nor U14723 (N_14723,N_13354,N_13929);
nor U14724 (N_14724,N_14295,N_14154);
or U14725 (N_14725,N_14054,N_13808);
and U14726 (N_14726,N_13302,N_13300);
xnor U14727 (N_14727,N_13806,N_13736);
and U14728 (N_14728,N_13470,N_13605);
xnor U14729 (N_14729,N_13572,N_13790);
and U14730 (N_14730,N_13571,N_13200);
nand U14731 (N_14731,N_14104,N_14161);
nand U14732 (N_14732,N_14176,N_13658);
xor U14733 (N_14733,N_14375,N_14284);
xor U14734 (N_14734,N_13404,N_14092);
or U14735 (N_14735,N_14168,N_13977);
nor U14736 (N_14736,N_13630,N_14111);
nand U14737 (N_14737,N_13538,N_13370);
or U14738 (N_14738,N_13649,N_14156);
nand U14739 (N_14739,N_13430,N_14230);
and U14740 (N_14740,N_13788,N_14086);
xor U14741 (N_14741,N_13334,N_13476);
and U14742 (N_14742,N_13774,N_13843);
xnor U14743 (N_14743,N_13509,N_13323);
and U14744 (N_14744,N_14000,N_14029);
xnor U14745 (N_14745,N_14252,N_13582);
nor U14746 (N_14746,N_14381,N_13719);
xor U14747 (N_14747,N_13681,N_13685);
nand U14748 (N_14748,N_13345,N_14251);
nor U14749 (N_14749,N_14048,N_14028);
xnor U14750 (N_14750,N_13426,N_13586);
xor U14751 (N_14751,N_13941,N_13306);
nand U14752 (N_14752,N_13548,N_14188);
nand U14753 (N_14753,N_13976,N_13928);
nand U14754 (N_14754,N_13734,N_13707);
and U14755 (N_14755,N_13814,N_14143);
nand U14756 (N_14756,N_14201,N_14304);
nand U14757 (N_14757,N_13473,N_13448);
xor U14758 (N_14758,N_13479,N_13358);
and U14759 (N_14759,N_14379,N_14359);
nor U14760 (N_14760,N_13403,N_13505);
or U14761 (N_14761,N_13361,N_14062);
nor U14762 (N_14762,N_14118,N_13731);
or U14763 (N_14763,N_13312,N_14116);
nor U14764 (N_14764,N_14309,N_13826);
and U14765 (N_14765,N_13951,N_13910);
and U14766 (N_14766,N_13389,N_13564);
nor U14767 (N_14767,N_13795,N_14223);
and U14768 (N_14768,N_14017,N_14286);
or U14769 (N_14769,N_13597,N_13371);
nor U14770 (N_14770,N_13752,N_13962);
nor U14771 (N_14771,N_14278,N_14009);
and U14772 (N_14772,N_14228,N_14316);
or U14773 (N_14773,N_13959,N_14074);
nand U14774 (N_14774,N_14313,N_13674);
nor U14775 (N_14775,N_13339,N_13510);
xnor U14776 (N_14776,N_13988,N_13507);
nor U14777 (N_14777,N_14095,N_13435);
nand U14778 (N_14778,N_14348,N_13837);
nand U14779 (N_14779,N_14200,N_13985);
or U14780 (N_14780,N_14224,N_14079);
xor U14781 (N_14781,N_14305,N_14087);
nand U14782 (N_14782,N_13862,N_13382);
xor U14783 (N_14783,N_13576,N_13495);
nand U14784 (N_14784,N_13267,N_13488);
nand U14785 (N_14785,N_14358,N_13911);
xnor U14786 (N_14786,N_13322,N_13460);
xor U14787 (N_14787,N_13213,N_13366);
nand U14788 (N_14788,N_13965,N_13600);
nand U14789 (N_14789,N_14081,N_13604);
or U14790 (N_14790,N_14136,N_14149);
or U14791 (N_14791,N_13547,N_14237);
nor U14792 (N_14792,N_14376,N_13883);
xnor U14793 (N_14793,N_14275,N_13804);
nand U14794 (N_14794,N_13528,N_14183);
nor U14795 (N_14795,N_13613,N_14063);
or U14796 (N_14796,N_13778,N_13914);
and U14797 (N_14797,N_13756,N_14164);
or U14798 (N_14798,N_14383,N_14120);
xor U14799 (N_14799,N_13950,N_13802);
and U14800 (N_14800,N_13648,N_13210);
and U14801 (N_14801,N_13623,N_14122);
nand U14802 (N_14802,N_13703,N_13347);
xor U14803 (N_14803,N_13887,N_13614);
and U14804 (N_14804,N_13969,N_13478);
xor U14805 (N_14805,N_13878,N_13761);
or U14806 (N_14806,N_14287,N_13957);
nand U14807 (N_14807,N_13636,N_14362);
or U14808 (N_14808,N_14320,N_13549);
xor U14809 (N_14809,N_13317,N_14012);
and U14810 (N_14810,N_13205,N_13516);
nor U14811 (N_14811,N_14066,N_14033);
or U14812 (N_14812,N_13508,N_13422);
nand U14813 (N_14813,N_13848,N_14173);
xnor U14814 (N_14814,N_13777,N_14091);
nand U14815 (N_14815,N_13653,N_13879);
and U14816 (N_14816,N_13235,N_13935);
nor U14817 (N_14817,N_13642,N_13599);
nand U14818 (N_14818,N_14005,N_13747);
and U14819 (N_14819,N_13735,N_13320);
and U14820 (N_14820,N_14171,N_14355);
nor U14821 (N_14821,N_13585,N_13442);
and U14822 (N_14822,N_13697,N_14270);
xor U14823 (N_14823,N_13329,N_14135);
nor U14824 (N_14824,N_13385,N_14271);
xnor U14825 (N_14825,N_13445,N_13540);
and U14826 (N_14826,N_13715,N_14389);
or U14827 (N_14827,N_13429,N_13722);
xnor U14828 (N_14828,N_14019,N_14010);
nor U14829 (N_14829,N_13485,N_13402);
or U14830 (N_14830,N_14023,N_13693);
and U14831 (N_14831,N_13711,N_13530);
nand U14832 (N_14832,N_13609,N_13626);
xnor U14833 (N_14833,N_14138,N_14140);
nand U14834 (N_14834,N_14152,N_14158);
nor U14835 (N_14835,N_13617,N_13500);
nand U14836 (N_14836,N_14335,N_13293);
nor U14837 (N_14837,N_14020,N_14209);
nand U14838 (N_14838,N_13889,N_13632);
nand U14839 (N_14839,N_13744,N_14227);
nor U14840 (N_14840,N_14141,N_13922);
nor U14841 (N_14841,N_14127,N_14002);
or U14842 (N_14842,N_14256,N_13568);
nand U14843 (N_14843,N_14031,N_13566);
xor U14844 (N_14844,N_14145,N_13861);
and U14845 (N_14845,N_13881,N_13918);
xor U14846 (N_14846,N_13295,N_13525);
xor U14847 (N_14847,N_13575,N_14392);
or U14848 (N_14848,N_14131,N_13789);
and U14849 (N_14849,N_13610,N_14292);
nand U14850 (N_14850,N_13820,N_13698);
nor U14851 (N_14851,N_14013,N_13558);
nand U14852 (N_14852,N_13809,N_14179);
and U14853 (N_14853,N_13452,N_13701);
xor U14854 (N_14854,N_14298,N_13424);
nor U14855 (N_14855,N_13237,N_13824);
nor U14856 (N_14856,N_13901,N_13779);
xnor U14857 (N_14857,N_13930,N_14315);
and U14858 (N_14858,N_13892,N_13521);
and U14859 (N_14859,N_14155,N_13522);
xnor U14860 (N_14860,N_13660,N_14327);
nor U14861 (N_14861,N_13821,N_13327);
nand U14862 (N_14862,N_13829,N_13321);
or U14863 (N_14863,N_14094,N_13360);
and U14864 (N_14864,N_14243,N_13286);
and U14865 (N_14865,N_14247,N_14312);
nor U14866 (N_14866,N_14281,N_13287);
and U14867 (N_14867,N_13484,N_13691);
nand U14868 (N_14868,N_13376,N_13260);
nor U14869 (N_14869,N_13346,N_13368);
nor U14870 (N_14870,N_14371,N_14160);
nand U14871 (N_14871,N_13615,N_13407);
or U14872 (N_14872,N_13357,N_14083);
nor U14873 (N_14873,N_14300,N_13409);
and U14874 (N_14874,N_13699,N_13561);
xnor U14875 (N_14875,N_13348,N_14038);
nand U14876 (N_14876,N_14112,N_14206);
or U14877 (N_14877,N_13717,N_13464);
and U14878 (N_14878,N_13723,N_13939);
xor U14879 (N_14879,N_13748,N_13621);
nor U14880 (N_14880,N_13920,N_14266);
or U14881 (N_14881,N_13434,N_14182);
and U14882 (N_14882,N_13692,N_14245);
nand U14883 (N_14883,N_13439,N_13631);
xor U14884 (N_14884,N_13832,N_13587);
nand U14885 (N_14885,N_14008,N_13203);
and U14886 (N_14886,N_13215,N_14396);
nor U14887 (N_14887,N_13775,N_13860);
nor U14888 (N_14888,N_13446,N_13758);
xor U14889 (N_14889,N_14198,N_13675);
nor U14890 (N_14890,N_13456,N_13665);
and U14891 (N_14891,N_13383,N_13793);
and U14892 (N_14892,N_13694,N_13640);
nor U14893 (N_14893,N_13733,N_13211);
and U14894 (N_14894,N_14208,N_13739);
nor U14895 (N_14895,N_13443,N_13421);
or U14896 (N_14896,N_14159,N_14226);
nor U14897 (N_14897,N_14334,N_13818);
nor U14898 (N_14898,N_14294,N_14180);
nand U14899 (N_14899,N_13480,N_14349);
or U14900 (N_14900,N_14186,N_13457);
xor U14901 (N_14901,N_13830,N_13655);
xnor U14902 (N_14902,N_13849,N_13677);
nand U14903 (N_14903,N_13428,N_13384);
or U14904 (N_14904,N_13394,N_13634);
nand U14905 (N_14905,N_13518,N_13994);
xnor U14906 (N_14906,N_13377,N_13214);
xor U14907 (N_14907,N_14308,N_14386);
nand U14908 (N_14908,N_14238,N_13982);
or U14909 (N_14909,N_13512,N_13577);
nor U14910 (N_14910,N_13589,N_13781);
nand U14911 (N_14911,N_13584,N_14132);
or U14912 (N_14912,N_13916,N_13984);
nand U14913 (N_14913,N_13387,N_13314);
and U14914 (N_14914,N_13433,N_13380);
or U14915 (N_14915,N_13236,N_13622);
nand U14916 (N_14916,N_13909,N_13541);
nand U14917 (N_14917,N_13534,N_13700);
nor U14918 (N_14918,N_13372,N_13578);
or U14919 (N_14919,N_13657,N_13704);
or U14920 (N_14920,N_14339,N_13973);
nor U14921 (N_14921,N_13258,N_13635);
nor U14922 (N_14922,N_14084,N_14212);
and U14923 (N_14923,N_13493,N_13207);
nor U14924 (N_14924,N_13264,N_13241);
and U14925 (N_14925,N_13956,N_14076);
nand U14926 (N_14926,N_13786,N_13487);
or U14927 (N_14927,N_13813,N_13233);
or U14928 (N_14928,N_13720,N_13828);
nand U14929 (N_14929,N_13526,N_14195);
xnor U14930 (N_14930,N_14163,N_13328);
xor U14931 (N_14931,N_14254,N_13724);
and U14932 (N_14932,N_14110,N_14015);
nor U14933 (N_14933,N_13863,N_13875);
xnor U14934 (N_14934,N_13240,N_13997);
nor U14935 (N_14935,N_13854,N_13309);
xnor U14936 (N_14936,N_13955,N_13288);
or U14937 (N_14937,N_13274,N_14260);
and U14938 (N_14938,N_14192,N_14217);
nor U14939 (N_14939,N_13933,N_14096);
xor U14940 (N_14940,N_13841,N_14264);
or U14941 (N_14941,N_13220,N_14175);
nor U14942 (N_14942,N_14097,N_13668);
or U14943 (N_14943,N_14347,N_13307);
nand U14944 (N_14944,N_13680,N_13418);
nor U14945 (N_14945,N_13367,N_13900);
or U14946 (N_14946,N_13714,N_13773);
xor U14947 (N_14947,N_13570,N_14082);
or U14948 (N_14948,N_13299,N_14323);
nor U14949 (N_14949,N_13229,N_13948);
or U14950 (N_14950,N_13391,N_14067);
nand U14951 (N_14951,N_13716,N_13255);
nor U14952 (N_14952,N_13432,N_13563);
and U14953 (N_14953,N_13679,N_13772);
nand U14954 (N_14954,N_14027,N_13611);
or U14955 (N_14955,N_13543,N_14107);
nand U14956 (N_14956,N_13270,N_14345);
and U14957 (N_14957,N_14210,N_13940);
or U14958 (N_14958,N_14262,N_13482);
nand U14959 (N_14959,N_13705,N_13567);
nand U14960 (N_14960,N_13232,N_14244);
nand U14961 (N_14961,N_13490,N_13565);
nand U14962 (N_14962,N_13877,N_14283);
or U14963 (N_14963,N_13406,N_13291);
nand U14964 (N_14964,N_14040,N_14026);
and U14965 (N_14965,N_13870,N_13393);
and U14966 (N_14966,N_13625,N_13483);
or U14967 (N_14967,N_14369,N_13683);
nor U14968 (N_14968,N_14393,N_13246);
and U14969 (N_14969,N_13592,N_13966);
xnor U14970 (N_14970,N_13855,N_14044);
xor U14971 (N_14971,N_13782,N_14113);
nor U14972 (N_14972,N_13431,N_13753);
or U14973 (N_14973,N_13612,N_13633);
nand U14974 (N_14974,N_13990,N_13536);
xor U14975 (N_14975,N_14341,N_13856);
nor U14976 (N_14976,N_13271,N_13489);
or U14977 (N_14977,N_13261,N_13749);
or U14978 (N_14978,N_13871,N_13709);
xnor U14979 (N_14979,N_13318,N_13972);
and U14980 (N_14980,N_13763,N_14259);
or U14981 (N_14981,N_14072,N_13560);
or U14982 (N_14982,N_14229,N_13975);
nand U14983 (N_14983,N_13624,N_13395);
and U14984 (N_14984,N_13800,N_14196);
and U14985 (N_14985,N_13598,N_13591);
nand U14986 (N_14986,N_13276,N_14130);
nor U14987 (N_14987,N_13769,N_14055);
nor U14988 (N_14988,N_13926,N_13886);
and U14989 (N_14989,N_13908,N_13342);
nand U14990 (N_14990,N_14106,N_14293);
xnor U14991 (N_14991,N_13730,N_13682);
xor U14992 (N_14992,N_14360,N_13502);
and U14993 (N_14993,N_13949,N_13650);
nand U14994 (N_14994,N_13396,N_14041);
or U14995 (N_14995,N_13234,N_13438);
nor U14996 (N_14996,N_13746,N_13803);
nor U14997 (N_14997,N_14299,N_14166);
and U14998 (N_14998,N_13827,N_13290);
and U14999 (N_14999,N_13501,N_14390);
nor U15000 (N_15000,N_14153,N_13983);
nand U15001 (N_15001,N_13541,N_14098);
nand U15002 (N_15002,N_14353,N_13390);
nor U15003 (N_15003,N_14290,N_13847);
and U15004 (N_15004,N_13779,N_13433);
nand U15005 (N_15005,N_14302,N_13859);
nor U15006 (N_15006,N_13679,N_13985);
nand U15007 (N_15007,N_13657,N_14129);
xnor U15008 (N_15008,N_14192,N_13645);
or U15009 (N_15009,N_13774,N_14222);
or U15010 (N_15010,N_13818,N_13990);
nor U15011 (N_15011,N_13280,N_14134);
and U15012 (N_15012,N_13704,N_14101);
and U15013 (N_15013,N_13915,N_13240);
nand U15014 (N_15014,N_13851,N_13603);
xor U15015 (N_15015,N_14321,N_14249);
nand U15016 (N_15016,N_14249,N_14099);
and U15017 (N_15017,N_13504,N_13354);
nand U15018 (N_15018,N_13714,N_13271);
xor U15019 (N_15019,N_14169,N_13574);
nand U15020 (N_15020,N_14229,N_13905);
and U15021 (N_15021,N_14326,N_13992);
xor U15022 (N_15022,N_13840,N_14057);
and U15023 (N_15023,N_13787,N_14296);
or U15024 (N_15024,N_13943,N_14171);
xor U15025 (N_15025,N_13988,N_14371);
and U15026 (N_15026,N_14072,N_13811);
or U15027 (N_15027,N_13389,N_14236);
and U15028 (N_15028,N_13735,N_14221);
nor U15029 (N_15029,N_14178,N_14281);
nand U15030 (N_15030,N_13639,N_13551);
xor U15031 (N_15031,N_13403,N_13304);
xnor U15032 (N_15032,N_14197,N_13624);
nand U15033 (N_15033,N_13838,N_13894);
and U15034 (N_15034,N_13542,N_14144);
and U15035 (N_15035,N_13351,N_13799);
xor U15036 (N_15036,N_14235,N_13804);
xor U15037 (N_15037,N_13945,N_14309);
or U15038 (N_15038,N_13587,N_13312);
nand U15039 (N_15039,N_13217,N_13873);
nor U15040 (N_15040,N_13623,N_14173);
nand U15041 (N_15041,N_14326,N_13612);
nor U15042 (N_15042,N_13404,N_13468);
xnor U15043 (N_15043,N_13757,N_14218);
nand U15044 (N_15044,N_13969,N_14036);
xor U15045 (N_15045,N_14020,N_13603);
or U15046 (N_15046,N_14047,N_14283);
nor U15047 (N_15047,N_13707,N_13845);
xor U15048 (N_15048,N_14266,N_13300);
xnor U15049 (N_15049,N_13602,N_13695);
nand U15050 (N_15050,N_14223,N_14047);
nand U15051 (N_15051,N_14165,N_13998);
or U15052 (N_15052,N_13942,N_14376);
nand U15053 (N_15053,N_13228,N_13660);
and U15054 (N_15054,N_14029,N_13838);
xnor U15055 (N_15055,N_13593,N_14361);
nor U15056 (N_15056,N_14259,N_13334);
nand U15057 (N_15057,N_13865,N_13692);
nand U15058 (N_15058,N_14109,N_13415);
or U15059 (N_15059,N_14076,N_14157);
nor U15060 (N_15060,N_13414,N_13933);
xor U15061 (N_15061,N_13448,N_14210);
or U15062 (N_15062,N_13764,N_13750);
nand U15063 (N_15063,N_13544,N_13766);
and U15064 (N_15064,N_13449,N_14147);
nand U15065 (N_15065,N_13931,N_13252);
nand U15066 (N_15066,N_13617,N_14148);
nor U15067 (N_15067,N_13926,N_14341);
and U15068 (N_15068,N_14069,N_13852);
and U15069 (N_15069,N_13617,N_14046);
or U15070 (N_15070,N_13677,N_13464);
xnor U15071 (N_15071,N_13863,N_14152);
nand U15072 (N_15072,N_14124,N_13674);
nor U15073 (N_15073,N_13732,N_13222);
xor U15074 (N_15074,N_13237,N_14212);
xor U15075 (N_15075,N_13869,N_13468);
nand U15076 (N_15076,N_13541,N_13580);
nand U15077 (N_15077,N_13741,N_13892);
nand U15078 (N_15078,N_13572,N_13428);
nand U15079 (N_15079,N_13565,N_13869);
nor U15080 (N_15080,N_13288,N_13988);
nor U15081 (N_15081,N_13630,N_13371);
and U15082 (N_15082,N_14203,N_13520);
or U15083 (N_15083,N_13619,N_13335);
nand U15084 (N_15084,N_14132,N_13968);
nand U15085 (N_15085,N_13845,N_13890);
nor U15086 (N_15086,N_13404,N_13744);
or U15087 (N_15087,N_13588,N_13568);
and U15088 (N_15088,N_13585,N_13634);
nand U15089 (N_15089,N_13930,N_14154);
nand U15090 (N_15090,N_13444,N_13339);
nor U15091 (N_15091,N_14392,N_14226);
xor U15092 (N_15092,N_13861,N_14375);
xnor U15093 (N_15093,N_13284,N_13370);
nor U15094 (N_15094,N_13218,N_14337);
xnor U15095 (N_15095,N_14039,N_13769);
nor U15096 (N_15096,N_13266,N_13223);
nand U15097 (N_15097,N_14255,N_13325);
and U15098 (N_15098,N_13393,N_13879);
or U15099 (N_15099,N_14034,N_13754);
xnor U15100 (N_15100,N_13998,N_13447);
nand U15101 (N_15101,N_14299,N_13759);
nand U15102 (N_15102,N_14366,N_13271);
and U15103 (N_15103,N_14372,N_14095);
xnor U15104 (N_15104,N_14003,N_13516);
and U15105 (N_15105,N_14283,N_13336);
or U15106 (N_15106,N_13888,N_13971);
nor U15107 (N_15107,N_13307,N_14374);
nand U15108 (N_15108,N_13296,N_13393);
nor U15109 (N_15109,N_13214,N_14336);
or U15110 (N_15110,N_13734,N_13522);
or U15111 (N_15111,N_13574,N_14079);
nand U15112 (N_15112,N_13236,N_13458);
and U15113 (N_15113,N_13782,N_13370);
or U15114 (N_15114,N_13560,N_13694);
nand U15115 (N_15115,N_13937,N_13735);
xor U15116 (N_15116,N_14325,N_13291);
xnor U15117 (N_15117,N_14204,N_13955);
and U15118 (N_15118,N_13301,N_13609);
nand U15119 (N_15119,N_13895,N_14274);
nand U15120 (N_15120,N_13480,N_13439);
and U15121 (N_15121,N_14389,N_13399);
or U15122 (N_15122,N_14073,N_13583);
and U15123 (N_15123,N_13470,N_13959);
and U15124 (N_15124,N_13353,N_13396);
xnor U15125 (N_15125,N_13286,N_13984);
nand U15126 (N_15126,N_13211,N_14151);
nor U15127 (N_15127,N_13693,N_13677);
nand U15128 (N_15128,N_13893,N_13233);
xnor U15129 (N_15129,N_14339,N_13472);
nor U15130 (N_15130,N_13380,N_14375);
and U15131 (N_15131,N_14059,N_13280);
xor U15132 (N_15132,N_13505,N_14322);
nor U15133 (N_15133,N_13358,N_13855);
or U15134 (N_15134,N_14330,N_13792);
xnor U15135 (N_15135,N_13545,N_13954);
nor U15136 (N_15136,N_13506,N_13395);
or U15137 (N_15137,N_13670,N_14395);
or U15138 (N_15138,N_13714,N_13403);
or U15139 (N_15139,N_14352,N_13994);
nor U15140 (N_15140,N_13233,N_13375);
xnor U15141 (N_15141,N_13301,N_14388);
and U15142 (N_15142,N_14379,N_14237);
nand U15143 (N_15143,N_13933,N_13318);
nor U15144 (N_15144,N_13302,N_13689);
xnor U15145 (N_15145,N_13539,N_13370);
nor U15146 (N_15146,N_13641,N_14241);
nor U15147 (N_15147,N_13348,N_13852);
and U15148 (N_15148,N_14188,N_13386);
nor U15149 (N_15149,N_13906,N_14262);
nor U15150 (N_15150,N_13849,N_13667);
or U15151 (N_15151,N_13972,N_14083);
nand U15152 (N_15152,N_14054,N_13552);
nand U15153 (N_15153,N_13328,N_13883);
xnor U15154 (N_15154,N_14247,N_14245);
nand U15155 (N_15155,N_13271,N_14080);
nand U15156 (N_15156,N_14075,N_13937);
nor U15157 (N_15157,N_13671,N_13946);
nand U15158 (N_15158,N_13844,N_13872);
nor U15159 (N_15159,N_14377,N_13451);
and U15160 (N_15160,N_13781,N_14208);
or U15161 (N_15161,N_13645,N_13288);
xnor U15162 (N_15162,N_13270,N_14383);
xor U15163 (N_15163,N_13272,N_13968);
nand U15164 (N_15164,N_14148,N_13982);
or U15165 (N_15165,N_14059,N_13360);
or U15166 (N_15166,N_14154,N_13234);
and U15167 (N_15167,N_14398,N_13856);
or U15168 (N_15168,N_14391,N_13989);
or U15169 (N_15169,N_13833,N_13668);
nand U15170 (N_15170,N_13558,N_14061);
nor U15171 (N_15171,N_14216,N_13395);
nor U15172 (N_15172,N_13662,N_14106);
and U15173 (N_15173,N_13482,N_14376);
and U15174 (N_15174,N_13420,N_13948);
and U15175 (N_15175,N_14093,N_14111);
xnor U15176 (N_15176,N_13960,N_13987);
or U15177 (N_15177,N_13603,N_14274);
nand U15178 (N_15178,N_13707,N_13434);
xnor U15179 (N_15179,N_13735,N_13576);
nand U15180 (N_15180,N_13629,N_14088);
xnor U15181 (N_15181,N_13213,N_14157);
nand U15182 (N_15182,N_14038,N_13917);
and U15183 (N_15183,N_14123,N_14114);
nand U15184 (N_15184,N_13967,N_13700);
xor U15185 (N_15185,N_13340,N_14013);
and U15186 (N_15186,N_13743,N_14066);
or U15187 (N_15187,N_14076,N_14107);
nor U15188 (N_15188,N_13212,N_13977);
nor U15189 (N_15189,N_13932,N_14318);
and U15190 (N_15190,N_13747,N_13410);
nor U15191 (N_15191,N_14342,N_13539);
and U15192 (N_15192,N_13965,N_13801);
and U15193 (N_15193,N_13472,N_13727);
xnor U15194 (N_15194,N_13974,N_14025);
nor U15195 (N_15195,N_13846,N_13686);
nor U15196 (N_15196,N_13407,N_14383);
nor U15197 (N_15197,N_13362,N_13865);
nor U15198 (N_15198,N_14377,N_13812);
nor U15199 (N_15199,N_13322,N_13699);
nand U15200 (N_15200,N_13824,N_13675);
nand U15201 (N_15201,N_13837,N_13201);
xnor U15202 (N_15202,N_13643,N_13543);
nand U15203 (N_15203,N_14004,N_14197);
nand U15204 (N_15204,N_14171,N_13736);
xor U15205 (N_15205,N_13398,N_13289);
nor U15206 (N_15206,N_14380,N_14334);
and U15207 (N_15207,N_13797,N_13866);
nand U15208 (N_15208,N_13709,N_13216);
and U15209 (N_15209,N_14036,N_13599);
nand U15210 (N_15210,N_14302,N_13794);
or U15211 (N_15211,N_13862,N_14295);
nor U15212 (N_15212,N_13452,N_14361);
and U15213 (N_15213,N_13292,N_13513);
xnor U15214 (N_15214,N_13430,N_13613);
xnor U15215 (N_15215,N_13955,N_14084);
nand U15216 (N_15216,N_13972,N_13658);
xor U15217 (N_15217,N_13573,N_14090);
or U15218 (N_15218,N_14337,N_13795);
and U15219 (N_15219,N_14195,N_13602);
xor U15220 (N_15220,N_13589,N_13951);
nor U15221 (N_15221,N_14398,N_13538);
or U15222 (N_15222,N_13509,N_14133);
xor U15223 (N_15223,N_13381,N_13603);
or U15224 (N_15224,N_14129,N_13517);
and U15225 (N_15225,N_13824,N_13604);
xor U15226 (N_15226,N_13533,N_14363);
and U15227 (N_15227,N_13237,N_13347);
xnor U15228 (N_15228,N_13677,N_14110);
and U15229 (N_15229,N_13318,N_13437);
or U15230 (N_15230,N_14170,N_13342);
xor U15231 (N_15231,N_13586,N_13662);
nor U15232 (N_15232,N_13505,N_13745);
or U15233 (N_15233,N_13958,N_13680);
or U15234 (N_15234,N_13598,N_14312);
and U15235 (N_15235,N_13513,N_13273);
or U15236 (N_15236,N_14195,N_13693);
nand U15237 (N_15237,N_13353,N_13562);
nor U15238 (N_15238,N_13459,N_13556);
nand U15239 (N_15239,N_14028,N_13925);
or U15240 (N_15240,N_13479,N_13756);
xnor U15241 (N_15241,N_14316,N_13283);
xor U15242 (N_15242,N_13634,N_13641);
nor U15243 (N_15243,N_13899,N_13284);
nor U15244 (N_15244,N_13853,N_13234);
xnor U15245 (N_15245,N_13636,N_13464);
and U15246 (N_15246,N_13206,N_14210);
nor U15247 (N_15247,N_13549,N_14099);
nand U15248 (N_15248,N_13764,N_13251);
nand U15249 (N_15249,N_14392,N_13539);
nor U15250 (N_15250,N_13831,N_14129);
nand U15251 (N_15251,N_13346,N_13505);
nand U15252 (N_15252,N_14362,N_14103);
xor U15253 (N_15253,N_13908,N_13852);
nand U15254 (N_15254,N_13484,N_13695);
xor U15255 (N_15255,N_13492,N_14185);
nand U15256 (N_15256,N_13246,N_14208);
xor U15257 (N_15257,N_13273,N_14215);
or U15258 (N_15258,N_13601,N_13858);
and U15259 (N_15259,N_13565,N_13209);
xor U15260 (N_15260,N_13205,N_14221);
nand U15261 (N_15261,N_13756,N_13995);
nand U15262 (N_15262,N_13763,N_13857);
nor U15263 (N_15263,N_13910,N_13419);
xor U15264 (N_15264,N_13726,N_13346);
or U15265 (N_15265,N_13461,N_14222);
and U15266 (N_15266,N_13992,N_13525);
nand U15267 (N_15267,N_13227,N_14375);
nor U15268 (N_15268,N_14088,N_13472);
nor U15269 (N_15269,N_13438,N_13440);
xor U15270 (N_15270,N_13659,N_13497);
and U15271 (N_15271,N_13403,N_13205);
xor U15272 (N_15272,N_13432,N_14384);
nand U15273 (N_15273,N_14100,N_13895);
or U15274 (N_15274,N_13249,N_14378);
xnor U15275 (N_15275,N_13722,N_13397);
or U15276 (N_15276,N_14064,N_14167);
nand U15277 (N_15277,N_13773,N_13877);
or U15278 (N_15278,N_14064,N_14186);
or U15279 (N_15279,N_14098,N_13351);
or U15280 (N_15280,N_13648,N_13669);
nand U15281 (N_15281,N_14281,N_14266);
nor U15282 (N_15282,N_13564,N_13801);
and U15283 (N_15283,N_14128,N_13719);
xor U15284 (N_15284,N_13968,N_13451);
xnor U15285 (N_15285,N_13850,N_14163);
nand U15286 (N_15286,N_13262,N_13278);
nand U15287 (N_15287,N_13415,N_14312);
and U15288 (N_15288,N_13420,N_13867);
xnor U15289 (N_15289,N_14215,N_14059);
and U15290 (N_15290,N_13593,N_14239);
or U15291 (N_15291,N_13421,N_13567);
nor U15292 (N_15292,N_13483,N_13651);
nor U15293 (N_15293,N_13606,N_13422);
nand U15294 (N_15294,N_13648,N_14159);
nand U15295 (N_15295,N_13256,N_13550);
and U15296 (N_15296,N_14064,N_13935);
nand U15297 (N_15297,N_13344,N_13872);
xnor U15298 (N_15298,N_13340,N_14057);
xor U15299 (N_15299,N_14133,N_13365);
nor U15300 (N_15300,N_13417,N_14110);
nand U15301 (N_15301,N_13922,N_13737);
nor U15302 (N_15302,N_13328,N_13488);
and U15303 (N_15303,N_13215,N_14212);
or U15304 (N_15304,N_13813,N_13744);
or U15305 (N_15305,N_14272,N_13443);
xor U15306 (N_15306,N_13367,N_13778);
and U15307 (N_15307,N_13975,N_13685);
nor U15308 (N_15308,N_13275,N_13646);
and U15309 (N_15309,N_14376,N_13644);
or U15310 (N_15310,N_13316,N_13494);
nand U15311 (N_15311,N_14220,N_14165);
xor U15312 (N_15312,N_13354,N_13204);
nand U15313 (N_15313,N_13432,N_14345);
nand U15314 (N_15314,N_13246,N_14175);
or U15315 (N_15315,N_13673,N_14391);
and U15316 (N_15316,N_14217,N_14313);
and U15317 (N_15317,N_13342,N_14124);
and U15318 (N_15318,N_14254,N_13953);
nor U15319 (N_15319,N_13951,N_13970);
and U15320 (N_15320,N_13783,N_13562);
and U15321 (N_15321,N_14035,N_14313);
nand U15322 (N_15322,N_13674,N_13588);
or U15323 (N_15323,N_14042,N_14028);
nand U15324 (N_15324,N_13439,N_14013);
nand U15325 (N_15325,N_14165,N_13462);
nor U15326 (N_15326,N_13671,N_14234);
or U15327 (N_15327,N_14268,N_14324);
xnor U15328 (N_15328,N_13717,N_13499);
xor U15329 (N_15329,N_13250,N_13232);
nor U15330 (N_15330,N_13257,N_14391);
and U15331 (N_15331,N_13773,N_14107);
xor U15332 (N_15332,N_14270,N_14204);
or U15333 (N_15333,N_13558,N_14031);
or U15334 (N_15334,N_13911,N_13761);
and U15335 (N_15335,N_13788,N_13912);
nand U15336 (N_15336,N_13958,N_14389);
nor U15337 (N_15337,N_13353,N_14086);
and U15338 (N_15338,N_14132,N_13241);
nand U15339 (N_15339,N_13882,N_14328);
or U15340 (N_15340,N_13728,N_14067);
nand U15341 (N_15341,N_13633,N_14268);
xnor U15342 (N_15342,N_13325,N_14259);
nor U15343 (N_15343,N_13929,N_13899);
or U15344 (N_15344,N_13599,N_13727);
or U15345 (N_15345,N_13569,N_14394);
nor U15346 (N_15346,N_13698,N_14320);
nor U15347 (N_15347,N_14325,N_13765);
and U15348 (N_15348,N_13382,N_13626);
or U15349 (N_15349,N_13581,N_13931);
nand U15350 (N_15350,N_13641,N_14068);
or U15351 (N_15351,N_14008,N_13404);
nor U15352 (N_15352,N_13853,N_14161);
and U15353 (N_15353,N_13921,N_13363);
and U15354 (N_15354,N_13679,N_13912);
or U15355 (N_15355,N_13762,N_13313);
and U15356 (N_15356,N_14391,N_13923);
xor U15357 (N_15357,N_14244,N_14398);
or U15358 (N_15358,N_13852,N_14256);
and U15359 (N_15359,N_13354,N_14041);
or U15360 (N_15360,N_13420,N_13938);
or U15361 (N_15361,N_13458,N_13276);
and U15362 (N_15362,N_14188,N_13473);
and U15363 (N_15363,N_13614,N_14101);
xor U15364 (N_15364,N_13747,N_13893);
nor U15365 (N_15365,N_14126,N_13517);
and U15366 (N_15366,N_13853,N_13907);
and U15367 (N_15367,N_13983,N_13782);
and U15368 (N_15368,N_13257,N_14397);
and U15369 (N_15369,N_14135,N_14222);
or U15370 (N_15370,N_14188,N_13928);
or U15371 (N_15371,N_13967,N_14268);
and U15372 (N_15372,N_13524,N_14030);
nor U15373 (N_15373,N_13960,N_13647);
nand U15374 (N_15374,N_13294,N_13471);
or U15375 (N_15375,N_13678,N_14235);
or U15376 (N_15376,N_14020,N_13779);
nor U15377 (N_15377,N_13686,N_13376);
or U15378 (N_15378,N_13913,N_14204);
or U15379 (N_15379,N_14077,N_14046);
nand U15380 (N_15380,N_13946,N_13690);
xor U15381 (N_15381,N_13388,N_13674);
nor U15382 (N_15382,N_13816,N_14008);
nand U15383 (N_15383,N_14254,N_14261);
nor U15384 (N_15384,N_13372,N_13223);
nand U15385 (N_15385,N_13885,N_13479);
or U15386 (N_15386,N_13304,N_13759);
nand U15387 (N_15387,N_13904,N_13428);
xnor U15388 (N_15388,N_14032,N_13853);
and U15389 (N_15389,N_13522,N_13694);
nand U15390 (N_15390,N_14263,N_14177);
or U15391 (N_15391,N_14036,N_13519);
nand U15392 (N_15392,N_13447,N_13264);
and U15393 (N_15393,N_13269,N_13907);
nand U15394 (N_15394,N_14385,N_14327);
nand U15395 (N_15395,N_13989,N_14027);
nand U15396 (N_15396,N_13706,N_13273);
and U15397 (N_15397,N_14326,N_13953);
xor U15398 (N_15398,N_13503,N_13870);
xor U15399 (N_15399,N_13709,N_14300);
or U15400 (N_15400,N_13296,N_14118);
nor U15401 (N_15401,N_14389,N_13786);
or U15402 (N_15402,N_14085,N_13903);
xnor U15403 (N_15403,N_14096,N_13554);
xnor U15404 (N_15404,N_13669,N_13477);
and U15405 (N_15405,N_13417,N_13468);
nor U15406 (N_15406,N_13589,N_14142);
xnor U15407 (N_15407,N_14221,N_13366);
or U15408 (N_15408,N_13769,N_13426);
xnor U15409 (N_15409,N_14166,N_13748);
nor U15410 (N_15410,N_14291,N_13255);
or U15411 (N_15411,N_13344,N_13267);
xnor U15412 (N_15412,N_13608,N_13920);
or U15413 (N_15413,N_13269,N_14348);
and U15414 (N_15414,N_14084,N_13855);
and U15415 (N_15415,N_13881,N_13331);
xnor U15416 (N_15416,N_13884,N_14161);
and U15417 (N_15417,N_13698,N_13365);
and U15418 (N_15418,N_13874,N_13506);
and U15419 (N_15419,N_14350,N_13596);
and U15420 (N_15420,N_13973,N_14337);
xor U15421 (N_15421,N_14011,N_13370);
nand U15422 (N_15422,N_14355,N_13642);
or U15423 (N_15423,N_14008,N_13658);
nor U15424 (N_15424,N_13814,N_14326);
nor U15425 (N_15425,N_13798,N_13326);
or U15426 (N_15426,N_13616,N_13840);
nor U15427 (N_15427,N_14027,N_14232);
nor U15428 (N_15428,N_14151,N_13945);
nor U15429 (N_15429,N_13899,N_13331);
nor U15430 (N_15430,N_14244,N_14000);
nor U15431 (N_15431,N_14027,N_13245);
nor U15432 (N_15432,N_14145,N_13777);
and U15433 (N_15433,N_13924,N_13314);
or U15434 (N_15434,N_14315,N_14181);
and U15435 (N_15435,N_14138,N_14074);
xnor U15436 (N_15436,N_14297,N_13295);
nand U15437 (N_15437,N_13654,N_14256);
nand U15438 (N_15438,N_13227,N_13417);
xor U15439 (N_15439,N_13317,N_13537);
nor U15440 (N_15440,N_13684,N_13809);
or U15441 (N_15441,N_13814,N_14254);
or U15442 (N_15442,N_14099,N_14075);
nor U15443 (N_15443,N_14268,N_13261);
nor U15444 (N_15444,N_14339,N_13612);
nor U15445 (N_15445,N_14080,N_13842);
nor U15446 (N_15446,N_13210,N_13967);
nand U15447 (N_15447,N_13585,N_14267);
or U15448 (N_15448,N_14053,N_13303);
and U15449 (N_15449,N_14204,N_14194);
and U15450 (N_15450,N_13988,N_13687);
nor U15451 (N_15451,N_14335,N_14085);
and U15452 (N_15452,N_14168,N_13709);
or U15453 (N_15453,N_13284,N_13865);
or U15454 (N_15454,N_14378,N_13570);
nor U15455 (N_15455,N_14103,N_13813);
or U15456 (N_15456,N_13873,N_13729);
nand U15457 (N_15457,N_14013,N_13903);
nor U15458 (N_15458,N_13565,N_13690);
xnor U15459 (N_15459,N_13928,N_13745);
and U15460 (N_15460,N_13338,N_13419);
nor U15461 (N_15461,N_13899,N_13271);
nor U15462 (N_15462,N_13654,N_13568);
nand U15463 (N_15463,N_13358,N_13899);
xor U15464 (N_15464,N_14124,N_14388);
nand U15465 (N_15465,N_13363,N_13321);
xor U15466 (N_15466,N_13343,N_13974);
nor U15467 (N_15467,N_13438,N_14049);
nor U15468 (N_15468,N_13753,N_13604);
nor U15469 (N_15469,N_14229,N_13343);
nor U15470 (N_15470,N_14355,N_13879);
xor U15471 (N_15471,N_14110,N_13545);
nor U15472 (N_15472,N_13540,N_13538);
or U15473 (N_15473,N_13532,N_13220);
nor U15474 (N_15474,N_13707,N_14341);
nor U15475 (N_15475,N_14270,N_13597);
nand U15476 (N_15476,N_13726,N_14393);
nor U15477 (N_15477,N_13299,N_13308);
and U15478 (N_15478,N_14105,N_13675);
xnor U15479 (N_15479,N_13871,N_13529);
or U15480 (N_15480,N_14288,N_14247);
nor U15481 (N_15481,N_13913,N_14070);
nor U15482 (N_15482,N_14222,N_14342);
or U15483 (N_15483,N_14179,N_14042);
nor U15484 (N_15484,N_13387,N_13808);
nor U15485 (N_15485,N_13387,N_14181);
or U15486 (N_15486,N_14063,N_13233);
nand U15487 (N_15487,N_14108,N_13714);
nor U15488 (N_15488,N_13673,N_13818);
nand U15489 (N_15489,N_14336,N_13342);
or U15490 (N_15490,N_13764,N_13846);
nor U15491 (N_15491,N_14292,N_14038);
nor U15492 (N_15492,N_13944,N_14145);
and U15493 (N_15493,N_13979,N_13628);
and U15494 (N_15494,N_13335,N_13291);
and U15495 (N_15495,N_13819,N_13780);
nor U15496 (N_15496,N_14352,N_13761);
nor U15497 (N_15497,N_13873,N_13347);
xnor U15498 (N_15498,N_13420,N_14174);
nand U15499 (N_15499,N_13852,N_13258);
and U15500 (N_15500,N_13805,N_14236);
and U15501 (N_15501,N_14323,N_13753);
nor U15502 (N_15502,N_14017,N_14023);
nand U15503 (N_15503,N_13740,N_13852);
and U15504 (N_15504,N_13795,N_13654);
and U15505 (N_15505,N_13201,N_14097);
nand U15506 (N_15506,N_13868,N_14150);
and U15507 (N_15507,N_13218,N_13832);
or U15508 (N_15508,N_13924,N_14164);
and U15509 (N_15509,N_14017,N_13692);
and U15510 (N_15510,N_13325,N_13366);
xnor U15511 (N_15511,N_13703,N_13383);
nor U15512 (N_15512,N_14180,N_14181);
nor U15513 (N_15513,N_14266,N_14029);
and U15514 (N_15514,N_13568,N_14389);
xnor U15515 (N_15515,N_13464,N_13301);
or U15516 (N_15516,N_13261,N_13657);
nand U15517 (N_15517,N_13745,N_13882);
or U15518 (N_15518,N_13977,N_13365);
nand U15519 (N_15519,N_13948,N_14235);
or U15520 (N_15520,N_13530,N_13788);
nor U15521 (N_15521,N_14001,N_13833);
xnor U15522 (N_15522,N_13999,N_14063);
nand U15523 (N_15523,N_14330,N_13379);
or U15524 (N_15524,N_14079,N_14242);
and U15525 (N_15525,N_14359,N_13514);
or U15526 (N_15526,N_13639,N_14313);
nand U15527 (N_15527,N_13306,N_13276);
xnor U15528 (N_15528,N_13381,N_13615);
or U15529 (N_15529,N_13449,N_14123);
nand U15530 (N_15530,N_13513,N_13278);
or U15531 (N_15531,N_14301,N_13916);
nand U15532 (N_15532,N_14296,N_13731);
xor U15533 (N_15533,N_14155,N_13240);
nor U15534 (N_15534,N_14022,N_13867);
nor U15535 (N_15535,N_13624,N_13610);
or U15536 (N_15536,N_13526,N_13647);
nand U15537 (N_15537,N_13816,N_14353);
xor U15538 (N_15538,N_13881,N_13839);
nor U15539 (N_15539,N_14208,N_13269);
or U15540 (N_15540,N_13208,N_14282);
nand U15541 (N_15541,N_14169,N_13754);
nor U15542 (N_15542,N_13826,N_13200);
and U15543 (N_15543,N_13625,N_13332);
and U15544 (N_15544,N_14277,N_14035);
nand U15545 (N_15545,N_13666,N_13500);
xnor U15546 (N_15546,N_13936,N_14393);
nor U15547 (N_15547,N_13947,N_14131);
nor U15548 (N_15548,N_13776,N_13693);
and U15549 (N_15549,N_14043,N_13606);
nor U15550 (N_15550,N_13346,N_14198);
and U15551 (N_15551,N_13505,N_14112);
xor U15552 (N_15552,N_13270,N_14332);
and U15553 (N_15553,N_13941,N_14172);
and U15554 (N_15554,N_13295,N_13841);
nand U15555 (N_15555,N_14003,N_13648);
nand U15556 (N_15556,N_14193,N_14344);
nand U15557 (N_15557,N_13396,N_14222);
nor U15558 (N_15558,N_14246,N_13295);
xnor U15559 (N_15559,N_13359,N_13970);
nand U15560 (N_15560,N_13238,N_13223);
xnor U15561 (N_15561,N_13918,N_13320);
and U15562 (N_15562,N_13639,N_13335);
nand U15563 (N_15563,N_14223,N_14377);
or U15564 (N_15564,N_13744,N_13453);
and U15565 (N_15565,N_14049,N_13693);
and U15566 (N_15566,N_14311,N_13528);
or U15567 (N_15567,N_13583,N_13654);
xor U15568 (N_15568,N_14189,N_13216);
or U15569 (N_15569,N_14180,N_13691);
and U15570 (N_15570,N_14046,N_13239);
xor U15571 (N_15571,N_13217,N_13688);
nor U15572 (N_15572,N_14391,N_13560);
or U15573 (N_15573,N_14127,N_13210);
and U15574 (N_15574,N_13789,N_13936);
or U15575 (N_15575,N_14076,N_13660);
and U15576 (N_15576,N_13974,N_13324);
nor U15577 (N_15577,N_14052,N_14335);
xnor U15578 (N_15578,N_13721,N_13856);
xnor U15579 (N_15579,N_13587,N_13591);
or U15580 (N_15580,N_14066,N_13656);
xor U15581 (N_15581,N_13993,N_13853);
nor U15582 (N_15582,N_13927,N_13403);
and U15583 (N_15583,N_13504,N_14066);
nor U15584 (N_15584,N_14282,N_13855);
xor U15585 (N_15585,N_14344,N_13253);
nor U15586 (N_15586,N_14207,N_14221);
nor U15587 (N_15587,N_14149,N_14142);
or U15588 (N_15588,N_14294,N_14285);
or U15589 (N_15589,N_13370,N_14291);
nand U15590 (N_15590,N_13591,N_13258);
or U15591 (N_15591,N_13958,N_14155);
nand U15592 (N_15592,N_14294,N_13295);
nand U15593 (N_15593,N_14343,N_13707);
xnor U15594 (N_15594,N_14381,N_14350);
and U15595 (N_15595,N_13432,N_13558);
nor U15596 (N_15596,N_13852,N_13285);
nand U15597 (N_15597,N_13678,N_13290);
nand U15598 (N_15598,N_14251,N_13432);
or U15599 (N_15599,N_13673,N_14231);
nand U15600 (N_15600,N_15466,N_14790);
xnor U15601 (N_15601,N_14704,N_14748);
or U15602 (N_15602,N_15535,N_14950);
and U15603 (N_15603,N_15317,N_14799);
or U15604 (N_15604,N_14843,N_14451);
and U15605 (N_15605,N_14459,N_15365);
nand U15606 (N_15606,N_14415,N_15397);
nor U15607 (N_15607,N_14606,N_14924);
and U15608 (N_15608,N_15151,N_15178);
nor U15609 (N_15609,N_15085,N_15084);
xnor U15610 (N_15610,N_15552,N_15050);
and U15611 (N_15611,N_15055,N_15005);
nor U15612 (N_15612,N_15119,N_15006);
or U15613 (N_15613,N_14951,N_15237);
and U15614 (N_15614,N_14677,N_14519);
and U15615 (N_15615,N_14760,N_14825);
nand U15616 (N_15616,N_14873,N_15101);
nand U15617 (N_15617,N_14625,N_14724);
or U15618 (N_15618,N_15033,N_14721);
and U15619 (N_15619,N_14571,N_15459);
and U15620 (N_15620,N_14857,N_15412);
xnor U15621 (N_15621,N_14711,N_15590);
or U15622 (N_15622,N_14646,N_15143);
nor U15623 (N_15623,N_14972,N_15188);
nor U15624 (N_15624,N_15097,N_14653);
nand U15625 (N_15625,N_14822,N_14964);
or U15626 (N_15626,N_14481,N_15514);
xnor U15627 (N_15627,N_15189,N_15304);
xor U15628 (N_15628,N_15423,N_15374);
and U15629 (N_15629,N_14928,N_15471);
nand U15630 (N_15630,N_15594,N_14860);
nand U15631 (N_15631,N_15095,N_14896);
and U15632 (N_15632,N_15254,N_15127);
nor U15633 (N_15633,N_14727,N_14788);
nor U15634 (N_15634,N_14818,N_14626);
or U15635 (N_15635,N_15208,N_15421);
and U15636 (N_15636,N_15405,N_15286);
or U15637 (N_15637,N_14676,N_14439);
nand U15638 (N_15638,N_14448,N_14622);
nand U15639 (N_15639,N_15548,N_15303);
xnor U15640 (N_15640,N_14722,N_14440);
nor U15641 (N_15641,N_15464,N_14856);
or U15642 (N_15642,N_15318,N_14584);
xor U15643 (N_15643,N_14766,N_15001);
xor U15644 (N_15644,N_15149,N_14679);
nor U15645 (N_15645,N_14544,N_15527);
nor U15646 (N_15646,N_14779,N_15462);
nand U15647 (N_15647,N_14661,N_14462);
nor U15648 (N_15648,N_15370,N_14560);
nand U15649 (N_15649,N_15505,N_14968);
nor U15650 (N_15650,N_15394,N_15516);
nor U15651 (N_15651,N_15096,N_15408);
nor U15652 (N_15652,N_15146,N_14594);
xor U15653 (N_15653,N_14884,N_15575);
and U15654 (N_15654,N_15023,N_14740);
xor U15655 (N_15655,N_15571,N_14979);
or U15656 (N_15656,N_14613,N_15078);
xor U15657 (N_15657,N_15118,N_15285);
nor U15658 (N_15658,N_15413,N_14554);
or U15659 (N_15659,N_14791,N_15537);
nor U15660 (N_15660,N_14685,N_15128);
nand U15661 (N_15661,N_14808,N_15198);
and U15662 (N_15662,N_15339,N_14999);
nand U15663 (N_15663,N_14707,N_15551);
nand U15664 (N_15664,N_15214,N_14616);
and U15665 (N_15665,N_15159,N_15418);
and U15666 (N_15666,N_15599,N_15201);
xor U15667 (N_15667,N_15161,N_14890);
xor U15668 (N_15668,N_14658,N_15473);
and U15669 (N_15669,N_14854,N_14620);
and U15670 (N_15670,N_15320,N_15204);
nor U15671 (N_15671,N_14473,N_14934);
and U15672 (N_15672,N_15451,N_14739);
or U15673 (N_15673,N_15569,N_14432);
or U15674 (N_15674,N_15416,N_14744);
xnor U15675 (N_15675,N_15501,N_14590);
xnor U15676 (N_15676,N_14812,N_14819);
xor U15677 (N_15677,N_14773,N_15164);
nand U15678 (N_15678,N_15372,N_15034);
nor U15679 (N_15679,N_14757,N_15430);
or U15680 (N_15680,N_14976,N_14568);
or U15681 (N_15681,N_15327,N_15541);
nand U15682 (N_15682,N_15588,N_15270);
nand U15683 (N_15683,N_15349,N_15566);
xor U15684 (N_15684,N_15137,N_14428);
xor U15685 (N_15685,N_15586,N_14828);
nand U15686 (N_15686,N_15328,N_14863);
nand U15687 (N_15687,N_14602,N_15465);
and U15688 (N_15688,N_14703,N_15426);
nor U15689 (N_15689,N_15260,N_15579);
xor U15690 (N_15690,N_14635,N_14956);
nor U15691 (N_15691,N_14411,N_14689);
nand U15692 (N_15692,N_15207,N_15342);
and U15693 (N_15693,N_15082,N_15313);
nor U15694 (N_15694,N_14629,N_15242);
xnor U15695 (N_15695,N_14702,N_14595);
nor U15696 (N_15696,N_14518,N_15478);
or U15697 (N_15697,N_14971,N_15350);
nor U15698 (N_15698,N_14908,N_14452);
or U15699 (N_15699,N_15296,N_14484);
or U15700 (N_15700,N_15386,N_15446);
xnor U15701 (N_15701,N_15474,N_15246);
nor U15702 (N_15702,N_14930,N_14407);
or U15703 (N_15703,N_15308,N_15062);
xor U15704 (N_15704,N_14787,N_14705);
or U15705 (N_15705,N_14900,N_15597);
nor U15706 (N_15706,N_15112,N_15587);
nand U15707 (N_15707,N_14867,N_14586);
and U15708 (N_15708,N_14615,N_15414);
or U15709 (N_15709,N_14555,N_14585);
or U15710 (N_15710,N_15470,N_14521);
nor U15711 (N_15711,N_15441,N_15472);
xor U15712 (N_15712,N_15449,N_14463);
nand U15713 (N_15713,N_15574,N_14502);
and U15714 (N_15714,N_14531,N_15160);
xor U15715 (N_15715,N_15321,N_14438);
or U15716 (N_15716,N_14796,N_15582);
and U15717 (N_15717,N_14981,N_14641);
and U15718 (N_15718,N_14933,N_15503);
xor U15719 (N_15719,N_14923,N_15513);
or U15720 (N_15720,N_15506,N_14904);
xor U15721 (N_15721,N_14471,N_14751);
and U15722 (N_15722,N_15429,N_14800);
nand U15723 (N_15723,N_14445,N_14441);
xor U15724 (N_15724,N_14888,N_15126);
nand U15725 (N_15725,N_15142,N_14730);
or U15726 (N_15726,N_15382,N_14718);
nor U15727 (N_15727,N_15179,N_14985);
nor U15728 (N_15728,N_15280,N_15015);
nand U15729 (N_15729,N_15522,N_14576);
nand U15730 (N_15730,N_15243,N_15131);
nor U15731 (N_15731,N_15000,N_14894);
and U15732 (N_15732,N_14858,N_15493);
nor U15733 (N_15733,N_14477,N_14430);
or U15734 (N_15734,N_15115,N_15434);
or U15735 (N_15735,N_15197,N_15487);
xor U15736 (N_15736,N_14688,N_14480);
and U15737 (N_15737,N_14522,N_15066);
xnor U15738 (N_15738,N_15031,N_15038);
or U15739 (N_15739,N_14970,N_14823);
and U15740 (N_15740,N_15294,N_14909);
and U15741 (N_15741,N_14807,N_15538);
xor U15742 (N_15742,N_15185,N_15287);
and U15743 (N_15743,N_14424,N_15336);
nand U15744 (N_15744,N_14899,N_15549);
nand U15745 (N_15745,N_15224,N_15592);
nor U15746 (N_15746,N_15064,N_15401);
and U15747 (N_15747,N_14640,N_15199);
xor U15748 (N_15748,N_15297,N_15205);
nand U15749 (N_15749,N_14895,N_14533);
or U15750 (N_15750,N_15377,N_14446);
nand U15751 (N_15751,N_14617,N_14548);
or U15752 (N_15752,N_15043,N_15176);
and U15753 (N_15753,N_14862,N_15099);
nor U15754 (N_15754,N_15113,N_14755);
or U15755 (N_15755,N_14578,N_15329);
and U15756 (N_15756,N_15447,N_15218);
xnor U15757 (N_15757,N_15235,N_14944);
xnor U15758 (N_15758,N_14876,N_14815);
nor U15759 (N_15759,N_15358,N_14527);
xnor U15760 (N_15760,N_14458,N_14906);
xnor U15761 (N_15761,N_15404,N_15054);
or U15762 (N_15762,N_15340,N_15363);
xnor U15763 (N_15763,N_15443,N_14472);
and U15764 (N_15764,N_14804,N_15206);
xor U15765 (N_15765,N_14551,N_15075);
xor U15766 (N_15766,N_14589,N_14805);
or U15767 (N_15767,N_15019,N_15489);
xor U15768 (N_15768,N_14608,N_14660);
and U15769 (N_15769,N_14598,N_14511);
nor U15770 (N_15770,N_14770,N_15067);
and U15771 (N_15771,N_14575,N_14932);
nor U15772 (N_15772,N_14542,N_14793);
nand U15773 (N_15773,N_14992,N_14655);
or U15774 (N_15774,N_14997,N_14887);
xnor U15775 (N_15775,N_15145,N_15315);
nor U15776 (N_15776,N_15483,N_14547);
or U15777 (N_15777,N_14720,N_15162);
xnor U15778 (N_15778,N_15077,N_14729);
xor U15779 (N_15779,N_15212,N_15052);
nand U15780 (N_15780,N_15292,N_14435);
xor U15781 (N_15781,N_14714,N_14662);
xnor U15782 (N_15782,N_14574,N_15591);
xor U15783 (N_15783,N_15102,N_14738);
or U15784 (N_15784,N_15385,N_14678);
nor U15785 (N_15785,N_15236,N_15520);
nand U15786 (N_15786,N_15310,N_14680);
nor U15787 (N_15787,N_15016,N_15251);
nor U15788 (N_15788,N_15562,N_14965);
or U15789 (N_15789,N_15271,N_14572);
xnor U15790 (N_15790,N_14814,N_15532);
or U15791 (N_15791,N_14706,N_15356);
xor U15792 (N_15792,N_14806,N_14422);
nand U15793 (N_15793,N_15152,N_14947);
nand U15794 (N_15794,N_15158,N_14723);
or U15795 (N_15795,N_14499,N_14967);
and U15796 (N_15796,N_14496,N_15435);
nand U15797 (N_15797,N_14449,N_15458);
nand U15798 (N_15798,N_15531,N_15366);
or U15799 (N_15799,N_14565,N_14987);
and U15800 (N_15800,N_15330,N_14874);
or U15801 (N_15801,N_14645,N_15364);
nor U15802 (N_15802,N_14421,N_15529);
and U15803 (N_15803,N_15448,N_14743);
or U15804 (N_15804,N_15316,N_15193);
and U15805 (N_15805,N_15008,N_15182);
or U15806 (N_15806,N_15585,N_15452);
and U15807 (N_15807,N_15593,N_14798);
or U15808 (N_15808,N_15035,N_14975);
xnor U15809 (N_15809,N_15341,N_15378);
and U15810 (N_15810,N_14486,N_15135);
or U15811 (N_15811,N_15040,N_15511);
xor U15812 (N_15812,N_14903,N_14666);
xor U15813 (N_15813,N_15528,N_15504);
nand U15814 (N_15814,N_15192,N_14691);
xnor U15815 (N_15815,N_14937,N_14878);
xnor U15816 (N_15816,N_14945,N_15289);
or U15817 (N_15817,N_14506,N_14623);
xnor U15818 (N_15818,N_15556,N_15295);
xor U15819 (N_15819,N_14621,N_15150);
and U15820 (N_15820,N_15445,N_14986);
and U15821 (N_15821,N_14478,N_14665);
nand U15822 (N_15822,N_14758,N_14582);
nand U15823 (N_15823,N_15577,N_15334);
or U15824 (N_15824,N_15530,N_14960);
or U15825 (N_15825,N_15539,N_14604);
xor U15826 (N_15826,N_15515,N_14902);
nor U15827 (N_15827,N_14514,N_14483);
nand U15828 (N_15828,N_14893,N_15545);
xnor U15829 (N_15829,N_14817,N_15276);
nand U15830 (N_15830,N_15269,N_14919);
nor U15831 (N_15831,N_15589,N_15324);
xnor U15832 (N_15832,N_14786,N_15216);
and U15833 (N_15833,N_14456,N_14918);
nor U15834 (N_15834,N_15578,N_15524);
nor U15835 (N_15835,N_14657,N_15134);
and U15836 (N_15836,N_14603,N_14609);
xor U15837 (N_15837,N_15457,N_14423);
nor U15838 (N_15838,N_14840,N_15036);
xnor U15839 (N_15839,N_15444,N_14474);
nand U15840 (N_15840,N_14713,N_14882);
and U15841 (N_15841,N_14922,N_14675);
nor U15842 (N_15842,N_15110,N_14517);
or U15843 (N_15843,N_14410,N_15573);
nand U15844 (N_15844,N_15438,N_14619);
nor U15845 (N_15845,N_15220,N_15433);
xnor U15846 (N_15846,N_15581,N_15156);
or U15847 (N_15847,N_14417,N_15293);
or U15848 (N_15848,N_14712,N_14509);
xnor U15849 (N_15849,N_15299,N_14450);
and U15850 (N_15850,N_15173,N_14780);
nand U15851 (N_15851,N_14994,N_15094);
nand U15852 (N_15852,N_15463,N_15022);
or U15853 (N_15853,N_15155,N_14583);
nor U15854 (N_15854,N_14405,N_14427);
xor U15855 (N_15855,N_14413,N_15335);
and U15856 (N_15856,N_15076,N_15026);
and U15857 (N_15857,N_14643,N_15311);
nor U15858 (N_15858,N_15298,N_14842);
and U15859 (N_15859,N_14690,N_14859);
xnor U15860 (N_15860,N_14954,N_15042);
xor U15861 (N_15861,N_15027,N_14995);
or U15862 (N_15862,N_15406,N_15253);
nand U15863 (N_15863,N_15017,N_15091);
nand U15864 (N_15864,N_14672,N_15439);
xor U15865 (N_15865,N_14870,N_15277);
xnor U15866 (N_15866,N_14490,N_15547);
nand U15867 (N_15867,N_14813,N_15509);
nor U15868 (N_15868,N_14778,N_14837);
and U15869 (N_15869,N_15490,N_14570);
xnor U15870 (N_15870,N_14694,N_15229);
nor U15871 (N_15871,N_15092,N_14803);
nand U15872 (N_15872,N_14696,N_15512);
xnor U15873 (N_15873,N_14820,N_15526);
and U15874 (N_15874,N_14567,N_14768);
nand U15875 (N_15875,N_14830,N_14824);
nor U15876 (N_15876,N_15380,N_14401);
xor U15877 (N_15877,N_15125,N_15540);
or U15878 (N_15878,N_14540,N_15456);
or U15879 (N_15879,N_15171,N_15010);
nand U15880 (N_15880,N_14756,N_14461);
nor U15881 (N_15881,N_14535,N_15244);
nor U15882 (N_15882,N_15258,N_14493);
xnor U15883 (N_15883,N_14725,N_15352);
xor U15884 (N_15884,N_15454,N_15202);
nor U15885 (N_15885,N_14792,N_15544);
nand U15886 (N_15886,N_14871,N_15124);
nor U15887 (N_15887,N_14901,N_15122);
xnor U15888 (N_15888,N_15248,N_14912);
xor U15889 (N_15889,N_15180,N_14569);
and U15890 (N_15890,N_14507,N_15120);
nor U15891 (N_15891,N_15203,N_14667);
nor U15892 (N_15892,N_14684,N_15012);
and U15893 (N_15893,N_14539,N_15346);
and U15894 (N_15894,N_15411,N_15323);
or U15895 (N_15895,N_14916,N_15268);
nor U15896 (N_15896,N_14605,N_14425);
xnor U15897 (N_15897,N_15059,N_15166);
or U15898 (N_15898,N_15121,N_15139);
or U15899 (N_15899,N_14886,N_15533);
nand U15900 (N_15900,N_15420,N_14630);
nand U15901 (N_15901,N_15147,N_14664);
and U15902 (N_15902,N_15098,N_15056);
nor U15903 (N_15903,N_14774,N_14959);
nand U15904 (N_15904,N_15305,N_15422);
and U15905 (N_15905,N_14767,N_15360);
and U15906 (N_15906,N_15402,N_14416);
nand U15907 (N_15907,N_15554,N_15431);
or U15908 (N_15908,N_14505,N_14949);
and U15909 (N_15909,N_14556,N_15424);
nand U15910 (N_15910,N_14642,N_14716);
nor U15911 (N_15911,N_14731,N_15114);
nand U15912 (N_15912,N_15007,N_15428);
or U15913 (N_15913,N_15045,N_14732);
or U15914 (N_15914,N_14710,N_15028);
or U15915 (N_15915,N_15065,N_14885);
and U15916 (N_15916,N_15497,N_15563);
or U15917 (N_15917,N_15583,N_14797);
xor U15918 (N_15918,N_15263,N_14686);
nand U15919 (N_15919,N_14408,N_14580);
nor U15920 (N_15920,N_15494,N_15157);
and U15921 (N_15921,N_14742,N_14733);
and U15922 (N_15922,N_15089,N_14431);
and U15923 (N_15923,N_15387,N_15407);
xor U15924 (N_15924,N_15234,N_14973);
xor U15925 (N_15925,N_14437,N_14692);
nand U15926 (N_15926,N_14771,N_15278);
nand U15927 (N_15927,N_15020,N_14841);
or U15928 (N_15928,N_15072,N_15359);
and U15929 (N_15929,N_15499,N_15468);
nor U15930 (N_15930,N_14898,N_14697);
xor U15931 (N_15931,N_15502,N_14670);
or U15932 (N_15932,N_14400,N_15274);
nand U15933 (N_15933,N_14802,N_15106);
and U15934 (N_15934,N_14880,N_15314);
nand U15935 (N_15935,N_15174,N_14687);
nor U15936 (N_15936,N_15484,N_15518);
nand U15937 (N_15937,N_15083,N_15267);
nand U15938 (N_15938,N_15331,N_14599);
and U15939 (N_15939,N_15070,N_15553);
nand U15940 (N_15940,N_15261,N_14998);
or U15941 (N_15941,N_14469,N_14736);
nor U15942 (N_15942,N_14487,N_15024);
or U15943 (N_15943,N_14549,N_14782);
nor U15944 (N_15944,N_14877,N_15584);
or U15945 (N_15945,N_14838,N_15259);
nand U15946 (N_15946,N_14591,N_14831);
nand U15947 (N_15947,N_15536,N_14564);
xor U15948 (N_15948,N_15534,N_14980);
and U15949 (N_15949,N_15168,N_15148);
nor U15950 (N_15950,N_14983,N_14861);
or U15951 (N_15951,N_14404,N_14552);
xor U15952 (N_15952,N_14946,N_14753);
xor U15953 (N_15953,N_15351,N_14537);
nor U15954 (N_15954,N_15415,N_15307);
xnor U15955 (N_15955,N_14816,N_14419);
xnor U15956 (N_15956,N_15519,N_14750);
nor U15957 (N_15957,N_14915,N_14869);
nor U15958 (N_15958,N_14845,N_15279);
and U15959 (N_15959,N_15345,N_14488);
nand U15960 (N_15960,N_15500,N_15580);
and U15961 (N_15961,N_14953,N_15598);
nor U15962 (N_15962,N_15181,N_14939);
nor U15963 (N_15963,N_15565,N_14513);
xnor U15964 (N_15964,N_14957,N_15284);
nand U15965 (N_15965,N_15046,N_15461);
or U15966 (N_15966,N_15477,N_15032);
or U15967 (N_15967,N_15371,N_14464);
nand U15968 (N_15968,N_15302,N_14835);
or U15969 (N_15969,N_15343,N_15326);
or U15970 (N_15970,N_15576,N_14512);
or U15971 (N_15971,N_15211,N_15213);
nor U15972 (N_15972,N_15391,N_15495);
or U15973 (N_15973,N_14683,N_14897);
or U15974 (N_15974,N_14777,N_14941);
nor U15975 (N_15975,N_14996,N_14875);
and U15976 (N_15976,N_15368,N_15393);
or U15977 (N_15977,N_14978,N_14628);
or U15978 (N_15978,N_14592,N_14659);
nor U15979 (N_15979,N_15196,N_14961);
xor U15980 (N_15980,N_14699,N_15200);
nand U15981 (N_15981,N_14573,N_14520);
nor U15982 (N_15982,N_15123,N_14601);
or U15983 (N_15983,N_14810,N_15154);
nor U15984 (N_15984,N_14476,N_14546);
xnor U15985 (N_15985,N_14801,N_15090);
xnor U15986 (N_15986,N_15183,N_15309);
nand U15987 (N_15987,N_14865,N_15227);
or U15988 (N_15988,N_15288,N_15596);
and U15989 (N_15989,N_15469,N_14412);
xor U15990 (N_15990,N_14534,N_15088);
and U15991 (N_15991,N_14597,N_15283);
xor U15992 (N_15992,N_14479,N_15481);
nor U15993 (N_15993,N_15132,N_15570);
and U15994 (N_15994,N_14717,N_14631);
nor U15995 (N_15995,N_15319,N_15100);
nand U15996 (N_15996,N_15282,N_15133);
nand U15997 (N_15997,N_14809,N_14434);
and U15998 (N_15998,N_14526,N_14681);
nor U15999 (N_15999,N_15079,N_15567);
nand U16000 (N_16000,N_14455,N_15272);
nor U16001 (N_16001,N_15117,N_15560);
or U16002 (N_16002,N_15256,N_14468);
nand U16003 (N_16003,N_14562,N_15322);
nor U16004 (N_16004,N_14523,N_15029);
nor U16005 (N_16005,N_15510,N_15262);
nand U16006 (N_16006,N_14775,N_14403);
nor U16007 (N_16007,N_14715,N_15442);
or U16008 (N_16008,N_14891,N_15039);
nand U16009 (N_16009,N_14627,N_15144);
or U16010 (N_16010,N_15140,N_14414);
xnor U16011 (N_16011,N_14530,N_15376);
or U16012 (N_16012,N_14700,N_15427);
xnor U16013 (N_16013,N_15080,N_15247);
xor U16014 (N_16014,N_14889,N_14442);
nor U16015 (N_16015,N_14737,N_15488);
nor U16016 (N_16016,N_14913,N_15172);
nand U16017 (N_16017,N_14735,N_15230);
or U16018 (N_16018,N_15111,N_15561);
nand U16019 (N_16019,N_14637,N_15169);
nor U16020 (N_16020,N_15485,N_15003);
and U16021 (N_16021,N_14543,N_14963);
and U16022 (N_16022,N_14647,N_14639);
nand U16023 (N_16023,N_14508,N_14734);
or U16024 (N_16024,N_14776,N_14917);
xor U16025 (N_16025,N_14501,N_15018);
nand U16026 (N_16026,N_14827,N_14881);
and U16027 (N_16027,N_15093,N_15542);
xnor U16028 (N_16028,N_15222,N_15069);
and U16029 (N_16029,N_15013,N_14466);
and U16030 (N_16030,N_14600,N_14849);
and U16031 (N_16031,N_15306,N_14532);
or U16032 (N_16032,N_14610,N_14638);
nor U16033 (N_16033,N_15209,N_14495);
or U16034 (N_16034,N_15241,N_14418);
nand U16035 (N_16035,N_15257,N_14467);
nor U16036 (N_16036,N_15290,N_14529);
nand U16037 (N_16037,N_15396,N_14671);
xor U16038 (N_16038,N_15048,N_15353);
and U16039 (N_16039,N_15250,N_14654);
nor U16040 (N_16040,N_14673,N_15373);
xor U16041 (N_16041,N_14741,N_14650);
nand U16042 (N_16042,N_14545,N_15379);
or U16043 (N_16043,N_15239,N_15049);
or U16044 (N_16044,N_15116,N_14784);
or U16045 (N_16045,N_15060,N_14491);
nand U16046 (N_16046,N_14811,N_14510);
nor U16047 (N_16047,N_14762,N_14632);
nand U16048 (N_16048,N_14851,N_15348);
xor U16049 (N_16049,N_15167,N_14754);
nand U16050 (N_16050,N_14503,N_14772);
or U16051 (N_16051,N_14905,N_15063);
nor U16052 (N_16052,N_14651,N_14765);
xor U16053 (N_16053,N_15068,N_14444);
xnor U16054 (N_16054,N_15498,N_15482);
nor U16055 (N_16055,N_15354,N_15301);
or U16056 (N_16056,N_14420,N_15355);
or U16057 (N_16057,N_15014,N_15264);
or U16058 (N_16058,N_14826,N_14984);
and U16059 (N_16059,N_14541,N_14764);
nand U16060 (N_16060,N_15467,N_14852);
nor U16061 (N_16061,N_14931,N_14515);
nand U16062 (N_16062,N_14794,N_14990);
or U16063 (N_16063,N_14693,N_15086);
nor U16064 (N_16064,N_15187,N_15217);
or U16065 (N_16065,N_14761,N_14485);
and U16066 (N_16066,N_15389,N_15266);
and U16067 (N_16067,N_15333,N_15163);
nand U16068 (N_16068,N_15555,N_14864);
xor U16069 (N_16069,N_15037,N_15194);
xnor U16070 (N_16070,N_15184,N_14524);
xnor U16071 (N_16071,N_14952,N_15523);
or U16072 (N_16072,N_14847,N_14497);
xnor U16073 (N_16073,N_15480,N_15332);
or U16074 (N_16074,N_14566,N_15265);
xnor U16075 (N_16075,N_15232,N_14936);
or U16076 (N_16076,N_15357,N_15177);
xnor U16077 (N_16077,N_15375,N_14848);
and U16078 (N_16078,N_14648,N_14465);
or U16079 (N_16079,N_14429,N_14698);
nor U16080 (N_16080,N_15105,N_14855);
nand U16081 (N_16081,N_15312,N_15507);
nand U16082 (N_16082,N_14433,N_15273);
xor U16083 (N_16083,N_14596,N_14577);
or U16084 (N_16084,N_15170,N_15002);
and U16085 (N_16085,N_14853,N_14669);
and U16086 (N_16086,N_14614,N_15399);
nand U16087 (N_16087,N_15436,N_14844);
nand U16088 (N_16088,N_15362,N_14726);
or U16089 (N_16089,N_15004,N_15476);
or U16090 (N_16090,N_14550,N_15338);
or U16091 (N_16091,N_14977,N_15044);
nand U16092 (N_16092,N_14783,N_15419);
or U16093 (N_16093,N_14879,N_15245);
or U16094 (N_16094,N_15153,N_14553);
or U16095 (N_16095,N_14929,N_15240);
and U16096 (N_16096,N_15425,N_14695);
nand U16097 (N_16097,N_14426,N_14850);
or U16098 (N_16098,N_14839,N_14636);
and U16099 (N_16099,N_14475,N_14557);
nand U16100 (N_16100,N_15103,N_14447);
nand U16101 (N_16101,N_15165,N_15300);
nor U16102 (N_16102,N_15369,N_14579);
nand U16103 (N_16103,N_15337,N_15210);
nand U16104 (N_16104,N_15252,N_15410);
nor U16105 (N_16105,N_15074,N_14538);
or U16106 (N_16106,N_15508,N_14674);
xor U16107 (N_16107,N_15073,N_15453);
xnor U16108 (N_16108,N_14728,N_15395);
xor U16109 (N_16109,N_14454,N_14991);
and U16110 (N_16110,N_14436,N_14498);
or U16111 (N_16111,N_14846,N_14914);
or U16112 (N_16112,N_14892,N_14872);
and U16113 (N_16113,N_15238,N_14866);
and U16114 (N_16114,N_14500,N_14607);
and U16115 (N_16115,N_14832,N_14821);
xor U16116 (N_16116,N_15550,N_14644);
nor U16117 (N_16117,N_15417,N_15543);
nand U16118 (N_16118,N_15190,N_15136);
nor U16119 (N_16119,N_14745,N_14920);
and U16120 (N_16120,N_14561,N_14559);
or U16121 (N_16121,N_14988,N_14868);
or U16122 (N_16122,N_14955,N_15195);
and U16123 (N_16123,N_15525,N_14940);
or U16124 (N_16124,N_15025,N_14935);
xor U16125 (N_16125,N_14482,N_14969);
xnor U16126 (N_16126,N_14781,N_14942);
and U16127 (N_16127,N_14747,N_14962);
and U16128 (N_16128,N_14709,N_15361);
nor U16129 (N_16129,N_14993,N_14834);
xor U16130 (N_16130,N_15521,N_15061);
and U16131 (N_16131,N_14795,N_14656);
xnor U16132 (N_16132,N_14943,N_15440);
xnor U16133 (N_16133,N_15041,N_15233);
xnor U16134 (N_16134,N_15057,N_14883);
nand U16135 (N_16135,N_15546,N_14624);
nor U16136 (N_16136,N_15129,N_15479);
or U16137 (N_16137,N_15030,N_14402);
nor U16138 (N_16138,N_15568,N_14633);
nand U16139 (N_16139,N_15450,N_15011);
nand U16140 (N_16140,N_14581,N_15564);
or U16141 (N_16141,N_15572,N_14558);
nor U16142 (N_16142,N_14833,N_15432);
or U16143 (N_16143,N_15191,N_15231);
xnor U16144 (N_16144,N_15437,N_14789);
or U16145 (N_16145,N_15486,N_15557);
nor U16146 (N_16146,N_14668,N_14528);
and U16147 (N_16147,N_15517,N_14910);
nor U16148 (N_16148,N_15325,N_14409);
nand U16149 (N_16149,N_15475,N_15275);
xor U16150 (N_16150,N_15138,N_14911);
xor U16151 (N_16151,N_15291,N_15175);
nand U16152 (N_16152,N_15384,N_15219);
or U16153 (N_16153,N_15403,N_14406);
and U16154 (N_16154,N_15223,N_15281);
or U16155 (N_16155,N_15221,N_14966);
and U16156 (N_16156,N_15344,N_15058);
xor U16157 (N_16157,N_14982,N_14785);
or U16158 (N_16158,N_14489,N_15109);
nand U16159 (N_16159,N_14634,N_14663);
or U16160 (N_16160,N_14974,N_15367);
nor U16161 (N_16161,N_14769,N_14457);
and U16162 (N_16162,N_15392,N_15249);
or U16163 (N_16163,N_15081,N_14836);
or U16164 (N_16164,N_14504,N_14593);
nor U16165 (N_16165,N_14907,N_15215);
and U16166 (N_16166,N_14829,N_15595);
and U16167 (N_16167,N_14611,N_14470);
nand U16168 (N_16168,N_14649,N_14759);
nor U16169 (N_16169,N_15228,N_14921);
xnor U16170 (N_16170,N_15255,N_15053);
or U16171 (N_16171,N_15226,N_15390);
xor U16172 (N_16172,N_15141,N_14708);
and U16173 (N_16173,N_14563,N_15400);
or U16174 (N_16174,N_15492,N_15108);
nand U16175 (N_16175,N_15087,N_14926);
nor U16176 (N_16176,N_15009,N_14453);
nand U16177 (N_16177,N_15104,N_15383);
and U16178 (N_16178,N_14989,N_15558);
xnor U16179 (N_16179,N_14746,N_15347);
nand U16180 (N_16180,N_14652,N_15130);
or U16181 (N_16181,N_14492,N_15381);
nand U16182 (N_16182,N_15021,N_14682);
nor U16183 (N_16183,N_15398,N_14494);
xnor U16184 (N_16184,N_15047,N_14460);
xor U16185 (N_16185,N_15051,N_14925);
xnor U16186 (N_16186,N_14536,N_15491);
xnor U16187 (N_16187,N_15559,N_15071);
xor U16188 (N_16188,N_15409,N_15107);
or U16189 (N_16189,N_14612,N_14588);
nor U16190 (N_16190,N_14516,N_14701);
or U16191 (N_16191,N_14958,N_14948);
and U16192 (N_16192,N_15496,N_14618);
and U16193 (N_16193,N_14525,N_15225);
and U16194 (N_16194,N_14938,N_15460);
and U16195 (N_16195,N_14927,N_14749);
or U16196 (N_16196,N_14752,N_14763);
nor U16197 (N_16197,N_15186,N_14443);
xor U16198 (N_16198,N_14587,N_15455);
nor U16199 (N_16199,N_15388,N_14719);
xnor U16200 (N_16200,N_14946,N_15395);
or U16201 (N_16201,N_15461,N_14463);
xnor U16202 (N_16202,N_14461,N_15452);
xnor U16203 (N_16203,N_14881,N_14943);
xnor U16204 (N_16204,N_15092,N_15584);
xnor U16205 (N_16205,N_15505,N_15291);
xor U16206 (N_16206,N_15216,N_15562);
nand U16207 (N_16207,N_15451,N_14823);
xnor U16208 (N_16208,N_14565,N_15528);
or U16209 (N_16209,N_15018,N_15046);
or U16210 (N_16210,N_14623,N_15300);
and U16211 (N_16211,N_15117,N_15266);
xor U16212 (N_16212,N_14511,N_14641);
nor U16213 (N_16213,N_14603,N_15344);
xnor U16214 (N_16214,N_14660,N_14499);
and U16215 (N_16215,N_15236,N_14599);
xor U16216 (N_16216,N_14546,N_15265);
xnor U16217 (N_16217,N_15042,N_15301);
nor U16218 (N_16218,N_14588,N_14576);
nor U16219 (N_16219,N_14853,N_15538);
nor U16220 (N_16220,N_15528,N_15301);
or U16221 (N_16221,N_14564,N_15193);
nor U16222 (N_16222,N_14861,N_15270);
nor U16223 (N_16223,N_15373,N_15539);
xor U16224 (N_16224,N_15270,N_15397);
nor U16225 (N_16225,N_15540,N_15516);
and U16226 (N_16226,N_15367,N_15231);
xor U16227 (N_16227,N_14949,N_14849);
xor U16228 (N_16228,N_15585,N_15249);
nor U16229 (N_16229,N_14900,N_15247);
nor U16230 (N_16230,N_15430,N_14988);
or U16231 (N_16231,N_14650,N_15569);
or U16232 (N_16232,N_15560,N_14952);
nand U16233 (N_16233,N_14469,N_14916);
nor U16234 (N_16234,N_14566,N_14545);
xnor U16235 (N_16235,N_15508,N_15445);
nand U16236 (N_16236,N_14472,N_14895);
nand U16237 (N_16237,N_14870,N_15051);
nor U16238 (N_16238,N_15018,N_14497);
xnor U16239 (N_16239,N_15338,N_15308);
xnor U16240 (N_16240,N_15333,N_14852);
xor U16241 (N_16241,N_14479,N_15476);
xor U16242 (N_16242,N_15229,N_14582);
xor U16243 (N_16243,N_14751,N_15289);
xor U16244 (N_16244,N_14466,N_15336);
or U16245 (N_16245,N_14500,N_14515);
nor U16246 (N_16246,N_14516,N_14875);
or U16247 (N_16247,N_15585,N_15235);
or U16248 (N_16248,N_14514,N_15480);
nand U16249 (N_16249,N_15431,N_15344);
and U16250 (N_16250,N_15355,N_15453);
and U16251 (N_16251,N_15279,N_14760);
or U16252 (N_16252,N_15362,N_15209);
and U16253 (N_16253,N_14569,N_15295);
or U16254 (N_16254,N_15264,N_14539);
nand U16255 (N_16255,N_14981,N_14895);
or U16256 (N_16256,N_14539,N_14816);
xnor U16257 (N_16257,N_14843,N_14972);
nor U16258 (N_16258,N_14473,N_14632);
xor U16259 (N_16259,N_14468,N_15009);
xnor U16260 (N_16260,N_15200,N_14931);
xor U16261 (N_16261,N_15477,N_14573);
nand U16262 (N_16262,N_15522,N_14521);
nor U16263 (N_16263,N_14485,N_14665);
or U16264 (N_16264,N_15419,N_15176);
nand U16265 (N_16265,N_14782,N_15558);
and U16266 (N_16266,N_15406,N_15261);
nor U16267 (N_16267,N_15216,N_15214);
nor U16268 (N_16268,N_14616,N_15312);
or U16269 (N_16269,N_14529,N_14716);
nand U16270 (N_16270,N_14484,N_15022);
or U16271 (N_16271,N_15430,N_15152);
and U16272 (N_16272,N_15417,N_15234);
and U16273 (N_16273,N_14432,N_15114);
and U16274 (N_16274,N_15316,N_14401);
nand U16275 (N_16275,N_15502,N_14903);
nand U16276 (N_16276,N_14968,N_15458);
xnor U16277 (N_16277,N_15576,N_15524);
and U16278 (N_16278,N_15100,N_14658);
and U16279 (N_16279,N_14646,N_15121);
and U16280 (N_16280,N_14866,N_15049);
nand U16281 (N_16281,N_14454,N_14939);
and U16282 (N_16282,N_14661,N_14711);
xnor U16283 (N_16283,N_15294,N_15149);
nor U16284 (N_16284,N_15357,N_15471);
nor U16285 (N_16285,N_14527,N_15128);
nand U16286 (N_16286,N_15591,N_14501);
xnor U16287 (N_16287,N_15028,N_15046);
nor U16288 (N_16288,N_15026,N_14960);
xor U16289 (N_16289,N_15386,N_15347);
xor U16290 (N_16290,N_15271,N_15593);
nor U16291 (N_16291,N_14803,N_15124);
xnor U16292 (N_16292,N_15057,N_15202);
nor U16293 (N_16293,N_14683,N_14692);
nor U16294 (N_16294,N_14632,N_15443);
and U16295 (N_16295,N_15343,N_14680);
nor U16296 (N_16296,N_15150,N_15489);
nand U16297 (N_16297,N_14778,N_14581);
nor U16298 (N_16298,N_14956,N_14488);
nand U16299 (N_16299,N_14690,N_15472);
nand U16300 (N_16300,N_14615,N_15072);
and U16301 (N_16301,N_15468,N_15236);
nand U16302 (N_16302,N_14608,N_14909);
nor U16303 (N_16303,N_14449,N_15064);
xor U16304 (N_16304,N_15006,N_15345);
nor U16305 (N_16305,N_15450,N_14797);
xnor U16306 (N_16306,N_15316,N_14884);
nor U16307 (N_16307,N_14759,N_14449);
nand U16308 (N_16308,N_15595,N_15152);
or U16309 (N_16309,N_14451,N_14718);
xnor U16310 (N_16310,N_15429,N_14620);
or U16311 (N_16311,N_14653,N_14406);
xor U16312 (N_16312,N_14670,N_15247);
and U16313 (N_16313,N_15290,N_14773);
nand U16314 (N_16314,N_15374,N_14508);
nor U16315 (N_16315,N_14936,N_15250);
xor U16316 (N_16316,N_14930,N_15227);
nand U16317 (N_16317,N_14683,N_14523);
nand U16318 (N_16318,N_14570,N_15186);
nor U16319 (N_16319,N_15387,N_14907);
and U16320 (N_16320,N_14459,N_15328);
or U16321 (N_16321,N_15256,N_15508);
or U16322 (N_16322,N_15017,N_14847);
or U16323 (N_16323,N_14980,N_15598);
and U16324 (N_16324,N_14920,N_15522);
and U16325 (N_16325,N_14616,N_15463);
nand U16326 (N_16326,N_15189,N_15282);
nand U16327 (N_16327,N_14478,N_14960);
and U16328 (N_16328,N_14687,N_15275);
nand U16329 (N_16329,N_15464,N_14981);
nand U16330 (N_16330,N_14576,N_14955);
and U16331 (N_16331,N_15297,N_14922);
nor U16332 (N_16332,N_15208,N_14830);
nor U16333 (N_16333,N_14661,N_15101);
nor U16334 (N_16334,N_14549,N_14424);
nand U16335 (N_16335,N_15572,N_15221);
xnor U16336 (N_16336,N_15546,N_14719);
and U16337 (N_16337,N_14779,N_15031);
and U16338 (N_16338,N_15382,N_14680);
nand U16339 (N_16339,N_15277,N_15303);
and U16340 (N_16340,N_14810,N_15451);
xor U16341 (N_16341,N_14766,N_14467);
and U16342 (N_16342,N_15479,N_15301);
nor U16343 (N_16343,N_14430,N_14647);
and U16344 (N_16344,N_15420,N_14678);
nor U16345 (N_16345,N_14824,N_14862);
nor U16346 (N_16346,N_15066,N_15378);
xor U16347 (N_16347,N_15123,N_15299);
and U16348 (N_16348,N_15427,N_14609);
xor U16349 (N_16349,N_14508,N_14518);
or U16350 (N_16350,N_15023,N_14949);
nor U16351 (N_16351,N_14406,N_14909);
nand U16352 (N_16352,N_14775,N_14947);
xor U16353 (N_16353,N_14416,N_14914);
nand U16354 (N_16354,N_15490,N_15471);
nand U16355 (N_16355,N_15474,N_15525);
nor U16356 (N_16356,N_14614,N_14609);
and U16357 (N_16357,N_14979,N_15440);
xnor U16358 (N_16358,N_14748,N_15311);
nand U16359 (N_16359,N_14834,N_14639);
nand U16360 (N_16360,N_14433,N_15284);
or U16361 (N_16361,N_14554,N_15512);
nand U16362 (N_16362,N_15135,N_15533);
xor U16363 (N_16363,N_15155,N_15299);
nand U16364 (N_16364,N_14679,N_14574);
nor U16365 (N_16365,N_14675,N_15006);
xor U16366 (N_16366,N_14687,N_15561);
xor U16367 (N_16367,N_15345,N_14484);
nor U16368 (N_16368,N_14916,N_14670);
nand U16369 (N_16369,N_15236,N_15456);
and U16370 (N_16370,N_14893,N_15367);
nand U16371 (N_16371,N_14935,N_14788);
nor U16372 (N_16372,N_14413,N_15373);
nand U16373 (N_16373,N_15046,N_15488);
nor U16374 (N_16374,N_15509,N_15177);
or U16375 (N_16375,N_15406,N_14953);
nand U16376 (N_16376,N_15597,N_15177);
or U16377 (N_16377,N_14911,N_14406);
nand U16378 (N_16378,N_14989,N_14638);
xnor U16379 (N_16379,N_14482,N_14449);
xnor U16380 (N_16380,N_15010,N_14778);
xnor U16381 (N_16381,N_14678,N_15088);
or U16382 (N_16382,N_14865,N_15379);
nand U16383 (N_16383,N_14890,N_15469);
nor U16384 (N_16384,N_14926,N_14738);
nor U16385 (N_16385,N_15325,N_15131);
or U16386 (N_16386,N_15324,N_14488);
or U16387 (N_16387,N_15516,N_15166);
nand U16388 (N_16388,N_14824,N_14507);
and U16389 (N_16389,N_15059,N_14685);
and U16390 (N_16390,N_14707,N_15322);
and U16391 (N_16391,N_15042,N_15188);
or U16392 (N_16392,N_15326,N_15295);
nor U16393 (N_16393,N_14638,N_14841);
or U16394 (N_16394,N_15557,N_15026);
xnor U16395 (N_16395,N_15458,N_15596);
and U16396 (N_16396,N_15075,N_15090);
nor U16397 (N_16397,N_15415,N_14717);
nor U16398 (N_16398,N_14407,N_15430);
and U16399 (N_16399,N_15494,N_14768);
nor U16400 (N_16400,N_14698,N_14640);
nor U16401 (N_16401,N_15181,N_15415);
xnor U16402 (N_16402,N_15378,N_14447);
and U16403 (N_16403,N_15351,N_15444);
xor U16404 (N_16404,N_14574,N_15568);
or U16405 (N_16405,N_15364,N_14928);
xor U16406 (N_16406,N_15309,N_14615);
xor U16407 (N_16407,N_14960,N_14788);
and U16408 (N_16408,N_15312,N_15598);
or U16409 (N_16409,N_15569,N_15235);
xnor U16410 (N_16410,N_15200,N_15553);
nor U16411 (N_16411,N_15276,N_15193);
nand U16412 (N_16412,N_14893,N_15263);
and U16413 (N_16413,N_14670,N_14516);
or U16414 (N_16414,N_15243,N_14412);
xor U16415 (N_16415,N_15318,N_15315);
or U16416 (N_16416,N_15034,N_14638);
nand U16417 (N_16417,N_15137,N_15213);
and U16418 (N_16418,N_14637,N_15165);
nand U16419 (N_16419,N_15089,N_14756);
xor U16420 (N_16420,N_14625,N_14666);
or U16421 (N_16421,N_15143,N_14514);
xnor U16422 (N_16422,N_14470,N_15152);
and U16423 (N_16423,N_15123,N_15095);
and U16424 (N_16424,N_15487,N_14604);
or U16425 (N_16425,N_14933,N_14784);
or U16426 (N_16426,N_14751,N_14629);
xnor U16427 (N_16427,N_15349,N_15101);
nand U16428 (N_16428,N_14550,N_15376);
or U16429 (N_16429,N_14558,N_15575);
or U16430 (N_16430,N_15472,N_15570);
and U16431 (N_16431,N_15481,N_15038);
xnor U16432 (N_16432,N_14706,N_14733);
and U16433 (N_16433,N_14513,N_15528);
and U16434 (N_16434,N_15543,N_14466);
or U16435 (N_16435,N_14909,N_14883);
nor U16436 (N_16436,N_14444,N_14811);
xor U16437 (N_16437,N_15344,N_15567);
nand U16438 (N_16438,N_15187,N_14656);
or U16439 (N_16439,N_14611,N_15146);
or U16440 (N_16440,N_14655,N_14615);
or U16441 (N_16441,N_14897,N_14747);
and U16442 (N_16442,N_14953,N_14728);
nand U16443 (N_16443,N_15500,N_14646);
nand U16444 (N_16444,N_14946,N_15595);
xor U16445 (N_16445,N_14908,N_15395);
and U16446 (N_16446,N_14906,N_14634);
or U16447 (N_16447,N_14482,N_14894);
nand U16448 (N_16448,N_14599,N_14505);
and U16449 (N_16449,N_14993,N_15499);
and U16450 (N_16450,N_15192,N_14539);
nand U16451 (N_16451,N_15084,N_15580);
nor U16452 (N_16452,N_14846,N_14593);
and U16453 (N_16453,N_15565,N_14665);
and U16454 (N_16454,N_14945,N_15021);
nor U16455 (N_16455,N_14811,N_15559);
nor U16456 (N_16456,N_14971,N_15300);
nand U16457 (N_16457,N_14753,N_14634);
nand U16458 (N_16458,N_15123,N_14781);
nand U16459 (N_16459,N_14647,N_14408);
or U16460 (N_16460,N_14934,N_14448);
nor U16461 (N_16461,N_15072,N_14604);
xor U16462 (N_16462,N_14756,N_14757);
and U16463 (N_16463,N_14995,N_15014);
nand U16464 (N_16464,N_15375,N_15597);
and U16465 (N_16465,N_14934,N_14414);
or U16466 (N_16466,N_14616,N_14653);
and U16467 (N_16467,N_14562,N_15349);
nor U16468 (N_16468,N_15337,N_15357);
or U16469 (N_16469,N_15511,N_14669);
and U16470 (N_16470,N_15297,N_14753);
xnor U16471 (N_16471,N_15080,N_15279);
and U16472 (N_16472,N_14875,N_15428);
nand U16473 (N_16473,N_15556,N_14685);
or U16474 (N_16474,N_14977,N_15551);
nor U16475 (N_16475,N_15555,N_14679);
nor U16476 (N_16476,N_15195,N_15027);
and U16477 (N_16477,N_15310,N_14926);
and U16478 (N_16478,N_14762,N_14963);
nor U16479 (N_16479,N_15247,N_15535);
nand U16480 (N_16480,N_14418,N_14545);
or U16481 (N_16481,N_15367,N_14538);
or U16482 (N_16482,N_15087,N_14764);
xnor U16483 (N_16483,N_15144,N_15477);
xnor U16484 (N_16484,N_14631,N_15254);
and U16485 (N_16485,N_15267,N_15376);
xor U16486 (N_16486,N_14411,N_14635);
or U16487 (N_16487,N_15570,N_15467);
or U16488 (N_16488,N_15568,N_15497);
xor U16489 (N_16489,N_14991,N_15497);
xnor U16490 (N_16490,N_15526,N_14734);
or U16491 (N_16491,N_14601,N_15227);
and U16492 (N_16492,N_14448,N_15371);
nand U16493 (N_16493,N_15127,N_14554);
and U16494 (N_16494,N_14522,N_15432);
and U16495 (N_16495,N_14548,N_14802);
nor U16496 (N_16496,N_14821,N_15448);
nand U16497 (N_16497,N_14587,N_14853);
xor U16498 (N_16498,N_15177,N_14871);
or U16499 (N_16499,N_14795,N_14451);
nand U16500 (N_16500,N_15282,N_15086);
and U16501 (N_16501,N_14514,N_15570);
nor U16502 (N_16502,N_14946,N_14732);
nor U16503 (N_16503,N_15410,N_14656);
nand U16504 (N_16504,N_15238,N_14551);
xnor U16505 (N_16505,N_14802,N_15314);
xor U16506 (N_16506,N_14401,N_14964);
and U16507 (N_16507,N_15085,N_14565);
and U16508 (N_16508,N_15588,N_14498);
nand U16509 (N_16509,N_15396,N_15319);
nor U16510 (N_16510,N_15198,N_14652);
xnor U16511 (N_16511,N_14975,N_15257);
and U16512 (N_16512,N_14655,N_15287);
nand U16513 (N_16513,N_15489,N_15202);
or U16514 (N_16514,N_14895,N_15355);
nand U16515 (N_16515,N_15143,N_14998);
xor U16516 (N_16516,N_15278,N_14675);
or U16517 (N_16517,N_14785,N_15217);
or U16518 (N_16518,N_14517,N_14820);
or U16519 (N_16519,N_15109,N_15299);
xor U16520 (N_16520,N_14595,N_14726);
nor U16521 (N_16521,N_14903,N_14583);
xor U16522 (N_16522,N_15475,N_15126);
or U16523 (N_16523,N_14487,N_14848);
nor U16524 (N_16524,N_14915,N_14653);
xnor U16525 (N_16525,N_14509,N_14587);
nand U16526 (N_16526,N_15142,N_15568);
nor U16527 (N_16527,N_14793,N_15028);
and U16528 (N_16528,N_15011,N_15209);
nor U16529 (N_16529,N_14614,N_15363);
nor U16530 (N_16530,N_15022,N_15079);
or U16531 (N_16531,N_15451,N_14417);
and U16532 (N_16532,N_15503,N_14633);
and U16533 (N_16533,N_15413,N_14493);
and U16534 (N_16534,N_14718,N_15175);
xor U16535 (N_16535,N_15186,N_14410);
or U16536 (N_16536,N_15012,N_14936);
or U16537 (N_16537,N_14881,N_14446);
and U16538 (N_16538,N_14908,N_14680);
or U16539 (N_16539,N_15481,N_15011);
nor U16540 (N_16540,N_14824,N_15200);
nand U16541 (N_16541,N_15574,N_14778);
nor U16542 (N_16542,N_15331,N_15462);
xnor U16543 (N_16543,N_14450,N_15304);
or U16544 (N_16544,N_14959,N_15016);
or U16545 (N_16545,N_14829,N_15509);
or U16546 (N_16546,N_15282,N_14777);
or U16547 (N_16547,N_14592,N_15130);
or U16548 (N_16548,N_14894,N_15491);
nand U16549 (N_16549,N_14687,N_14985);
or U16550 (N_16550,N_15022,N_14939);
nand U16551 (N_16551,N_14572,N_15430);
nand U16552 (N_16552,N_15553,N_14741);
or U16553 (N_16553,N_15235,N_14647);
or U16554 (N_16554,N_15188,N_15323);
nand U16555 (N_16555,N_14938,N_15148);
and U16556 (N_16556,N_15095,N_15369);
or U16557 (N_16557,N_15222,N_14668);
or U16558 (N_16558,N_14835,N_15546);
and U16559 (N_16559,N_15527,N_15566);
nand U16560 (N_16560,N_15419,N_14491);
nand U16561 (N_16561,N_15032,N_15462);
or U16562 (N_16562,N_14812,N_14730);
and U16563 (N_16563,N_14401,N_14733);
and U16564 (N_16564,N_14917,N_14890);
and U16565 (N_16565,N_14792,N_15213);
and U16566 (N_16566,N_15173,N_15204);
xor U16567 (N_16567,N_15515,N_14763);
nor U16568 (N_16568,N_15085,N_14858);
and U16569 (N_16569,N_14480,N_15160);
xor U16570 (N_16570,N_15280,N_14807);
and U16571 (N_16571,N_14509,N_14662);
and U16572 (N_16572,N_14900,N_14555);
and U16573 (N_16573,N_15000,N_15322);
xnor U16574 (N_16574,N_15221,N_14483);
or U16575 (N_16575,N_14547,N_14981);
nand U16576 (N_16576,N_14766,N_15189);
xnor U16577 (N_16577,N_15474,N_15308);
nor U16578 (N_16578,N_15459,N_15572);
xor U16579 (N_16579,N_15353,N_15218);
or U16580 (N_16580,N_14669,N_15032);
and U16581 (N_16581,N_15225,N_15249);
nand U16582 (N_16582,N_14666,N_15484);
or U16583 (N_16583,N_15524,N_15241);
nand U16584 (N_16584,N_15155,N_15144);
nand U16585 (N_16585,N_15008,N_14972);
nand U16586 (N_16586,N_14831,N_15092);
xor U16587 (N_16587,N_15257,N_14538);
and U16588 (N_16588,N_14571,N_15020);
or U16589 (N_16589,N_15327,N_15492);
or U16590 (N_16590,N_14698,N_15073);
nor U16591 (N_16591,N_14502,N_14828);
and U16592 (N_16592,N_15492,N_15099);
nand U16593 (N_16593,N_14800,N_14617);
xor U16594 (N_16594,N_14620,N_14644);
xnor U16595 (N_16595,N_15490,N_14426);
xnor U16596 (N_16596,N_14946,N_15535);
nand U16597 (N_16597,N_14797,N_14936);
nand U16598 (N_16598,N_15536,N_14569);
nor U16599 (N_16599,N_15291,N_15255);
and U16600 (N_16600,N_14725,N_14670);
and U16601 (N_16601,N_14537,N_14445);
or U16602 (N_16602,N_15563,N_14644);
xnor U16603 (N_16603,N_15058,N_14554);
nand U16604 (N_16604,N_15297,N_14600);
nor U16605 (N_16605,N_15166,N_15508);
xnor U16606 (N_16606,N_15197,N_15112);
nor U16607 (N_16607,N_15194,N_14732);
xnor U16608 (N_16608,N_14802,N_15107);
nor U16609 (N_16609,N_14899,N_15182);
xor U16610 (N_16610,N_15425,N_14754);
xor U16611 (N_16611,N_15558,N_14435);
and U16612 (N_16612,N_15302,N_14925);
nand U16613 (N_16613,N_14679,N_14469);
and U16614 (N_16614,N_15313,N_14824);
xor U16615 (N_16615,N_15533,N_14958);
nor U16616 (N_16616,N_15308,N_15309);
nand U16617 (N_16617,N_15243,N_14410);
nand U16618 (N_16618,N_14486,N_14724);
nor U16619 (N_16619,N_15267,N_15176);
and U16620 (N_16620,N_15014,N_14423);
and U16621 (N_16621,N_14766,N_14599);
or U16622 (N_16622,N_14602,N_15209);
xnor U16623 (N_16623,N_15364,N_14477);
nor U16624 (N_16624,N_14718,N_15404);
xor U16625 (N_16625,N_14401,N_15194);
and U16626 (N_16626,N_15546,N_15166);
xnor U16627 (N_16627,N_15200,N_14600);
or U16628 (N_16628,N_15022,N_15352);
nand U16629 (N_16629,N_14692,N_14415);
and U16630 (N_16630,N_14432,N_15071);
xnor U16631 (N_16631,N_14563,N_14651);
xor U16632 (N_16632,N_14553,N_15162);
nand U16633 (N_16633,N_14991,N_15112);
nor U16634 (N_16634,N_14752,N_15492);
or U16635 (N_16635,N_15306,N_15357);
nand U16636 (N_16636,N_15030,N_15488);
xnor U16637 (N_16637,N_15472,N_15213);
nor U16638 (N_16638,N_14911,N_15592);
or U16639 (N_16639,N_14801,N_14877);
nand U16640 (N_16640,N_15245,N_14613);
nand U16641 (N_16641,N_14539,N_15422);
xor U16642 (N_16642,N_15391,N_15163);
nand U16643 (N_16643,N_14684,N_14801);
nor U16644 (N_16644,N_15242,N_14450);
nor U16645 (N_16645,N_14589,N_14739);
or U16646 (N_16646,N_15364,N_14968);
or U16647 (N_16647,N_14538,N_14799);
and U16648 (N_16648,N_14710,N_14771);
nand U16649 (N_16649,N_14702,N_14726);
nand U16650 (N_16650,N_14954,N_15342);
nor U16651 (N_16651,N_14867,N_14971);
or U16652 (N_16652,N_14467,N_14542);
nand U16653 (N_16653,N_15423,N_15569);
xor U16654 (N_16654,N_15047,N_15330);
xnor U16655 (N_16655,N_14899,N_15316);
xnor U16656 (N_16656,N_14560,N_15550);
nand U16657 (N_16657,N_15381,N_15042);
xor U16658 (N_16658,N_14727,N_14573);
xor U16659 (N_16659,N_14497,N_14691);
nor U16660 (N_16660,N_14598,N_14474);
nand U16661 (N_16661,N_15058,N_15416);
xor U16662 (N_16662,N_14400,N_14558);
xnor U16663 (N_16663,N_14659,N_14685);
or U16664 (N_16664,N_15478,N_15109);
or U16665 (N_16665,N_14864,N_15273);
xor U16666 (N_16666,N_14457,N_15119);
or U16667 (N_16667,N_15449,N_14429);
xor U16668 (N_16668,N_14531,N_14481);
nor U16669 (N_16669,N_14433,N_15396);
nor U16670 (N_16670,N_15546,N_15343);
or U16671 (N_16671,N_15492,N_15356);
or U16672 (N_16672,N_14978,N_14935);
or U16673 (N_16673,N_15550,N_14902);
and U16674 (N_16674,N_15118,N_14961);
nor U16675 (N_16675,N_14567,N_15105);
or U16676 (N_16676,N_15366,N_14736);
xor U16677 (N_16677,N_14416,N_14712);
nand U16678 (N_16678,N_14903,N_14528);
or U16679 (N_16679,N_15496,N_14960);
xnor U16680 (N_16680,N_14901,N_15283);
or U16681 (N_16681,N_15143,N_15579);
nor U16682 (N_16682,N_14871,N_15578);
or U16683 (N_16683,N_14883,N_14839);
nor U16684 (N_16684,N_14405,N_15062);
and U16685 (N_16685,N_14889,N_15259);
and U16686 (N_16686,N_15081,N_15332);
nand U16687 (N_16687,N_14905,N_15183);
nor U16688 (N_16688,N_15465,N_14420);
or U16689 (N_16689,N_14893,N_14673);
nor U16690 (N_16690,N_14881,N_14687);
xor U16691 (N_16691,N_14968,N_15188);
nand U16692 (N_16692,N_14519,N_15352);
or U16693 (N_16693,N_14524,N_15368);
nand U16694 (N_16694,N_15462,N_15207);
and U16695 (N_16695,N_15330,N_15192);
nand U16696 (N_16696,N_15243,N_15371);
or U16697 (N_16697,N_14651,N_15024);
nor U16698 (N_16698,N_14823,N_15423);
and U16699 (N_16699,N_15525,N_15517);
or U16700 (N_16700,N_15554,N_14598);
xnor U16701 (N_16701,N_14464,N_15476);
and U16702 (N_16702,N_14490,N_14960);
or U16703 (N_16703,N_15197,N_14967);
or U16704 (N_16704,N_14751,N_15511);
xor U16705 (N_16705,N_15110,N_15117);
or U16706 (N_16706,N_15120,N_15589);
and U16707 (N_16707,N_14610,N_15527);
xor U16708 (N_16708,N_15196,N_15359);
xnor U16709 (N_16709,N_14971,N_15262);
or U16710 (N_16710,N_15342,N_14845);
xor U16711 (N_16711,N_15196,N_14692);
nor U16712 (N_16712,N_14646,N_14487);
xnor U16713 (N_16713,N_15289,N_15014);
nand U16714 (N_16714,N_14886,N_14643);
and U16715 (N_16715,N_14830,N_14879);
and U16716 (N_16716,N_15417,N_14772);
nor U16717 (N_16717,N_15305,N_14525);
or U16718 (N_16718,N_14701,N_15521);
and U16719 (N_16719,N_15499,N_15116);
xor U16720 (N_16720,N_14551,N_15064);
nand U16721 (N_16721,N_14997,N_14401);
nor U16722 (N_16722,N_15346,N_14485);
nor U16723 (N_16723,N_15451,N_15236);
nor U16724 (N_16724,N_15275,N_15283);
nor U16725 (N_16725,N_15018,N_14908);
nor U16726 (N_16726,N_14566,N_15515);
or U16727 (N_16727,N_15343,N_15226);
nand U16728 (N_16728,N_14640,N_14869);
nor U16729 (N_16729,N_15458,N_15267);
nor U16730 (N_16730,N_15322,N_15061);
nor U16731 (N_16731,N_14562,N_15565);
nor U16732 (N_16732,N_15365,N_14650);
xnor U16733 (N_16733,N_15445,N_14883);
and U16734 (N_16734,N_15282,N_14522);
nor U16735 (N_16735,N_14537,N_15375);
nor U16736 (N_16736,N_15350,N_15118);
xor U16737 (N_16737,N_14407,N_15217);
nor U16738 (N_16738,N_15580,N_14978);
nor U16739 (N_16739,N_15573,N_14651);
xnor U16740 (N_16740,N_14903,N_14730);
xnor U16741 (N_16741,N_14569,N_15188);
and U16742 (N_16742,N_14860,N_15375);
nor U16743 (N_16743,N_15151,N_14835);
nand U16744 (N_16744,N_15431,N_14960);
or U16745 (N_16745,N_14803,N_15165);
nor U16746 (N_16746,N_14538,N_14741);
nand U16747 (N_16747,N_15422,N_15119);
nand U16748 (N_16748,N_14945,N_14915);
xnor U16749 (N_16749,N_15081,N_15523);
nand U16750 (N_16750,N_14657,N_14816);
nand U16751 (N_16751,N_15507,N_15304);
xnor U16752 (N_16752,N_14998,N_14665);
xnor U16753 (N_16753,N_15463,N_14618);
and U16754 (N_16754,N_14867,N_14991);
nand U16755 (N_16755,N_15052,N_14415);
nand U16756 (N_16756,N_15114,N_15465);
xor U16757 (N_16757,N_14760,N_14890);
or U16758 (N_16758,N_15569,N_15440);
nor U16759 (N_16759,N_15143,N_14808);
nand U16760 (N_16760,N_15152,N_15583);
or U16761 (N_16761,N_15271,N_14512);
xor U16762 (N_16762,N_15264,N_15118);
nor U16763 (N_16763,N_14690,N_14867);
nor U16764 (N_16764,N_15026,N_14972);
nand U16765 (N_16765,N_14671,N_14831);
and U16766 (N_16766,N_14868,N_15382);
nor U16767 (N_16767,N_14909,N_15298);
xor U16768 (N_16768,N_14436,N_14569);
xor U16769 (N_16769,N_15209,N_14974);
nand U16770 (N_16770,N_14911,N_15356);
or U16771 (N_16771,N_14435,N_14617);
nand U16772 (N_16772,N_14885,N_14778);
and U16773 (N_16773,N_15481,N_14945);
xor U16774 (N_16774,N_14869,N_15518);
nand U16775 (N_16775,N_14502,N_15382);
xnor U16776 (N_16776,N_14659,N_14596);
or U16777 (N_16777,N_15233,N_15152);
and U16778 (N_16778,N_15156,N_15554);
or U16779 (N_16779,N_14748,N_15083);
or U16780 (N_16780,N_15044,N_15345);
xnor U16781 (N_16781,N_14455,N_15283);
xnor U16782 (N_16782,N_15525,N_15527);
nand U16783 (N_16783,N_15111,N_15301);
xnor U16784 (N_16784,N_15550,N_15097);
or U16785 (N_16785,N_15190,N_14490);
and U16786 (N_16786,N_15061,N_14586);
nand U16787 (N_16787,N_15261,N_14612);
and U16788 (N_16788,N_14602,N_14572);
and U16789 (N_16789,N_15007,N_14736);
or U16790 (N_16790,N_15349,N_15553);
nand U16791 (N_16791,N_14585,N_15269);
xor U16792 (N_16792,N_14583,N_15546);
nor U16793 (N_16793,N_14861,N_14838);
xnor U16794 (N_16794,N_14964,N_15349);
or U16795 (N_16795,N_14423,N_14686);
nor U16796 (N_16796,N_14512,N_14430);
xor U16797 (N_16797,N_15445,N_15046);
nor U16798 (N_16798,N_15196,N_15307);
or U16799 (N_16799,N_14548,N_15069);
nand U16800 (N_16800,N_16008,N_15632);
nor U16801 (N_16801,N_16139,N_16767);
or U16802 (N_16802,N_16229,N_15819);
nand U16803 (N_16803,N_15823,N_16630);
nand U16804 (N_16804,N_16213,N_15636);
or U16805 (N_16805,N_16769,N_16069);
or U16806 (N_16806,N_16304,N_16063);
and U16807 (N_16807,N_16572,N_16434);
nor U16808 (N_16808,N_15704,N_16297);
nor U16809 (N_16809,N_15779,N_15894);
nand U16810 (N_16810,N_16217,N_15837);
nand U16811 (N_16811,N_15911,N_16556);
nand U16812 (N_16812,N_15771,N_16151);
xnor U16813 (N_16813,N_15964,N_16453);
nor U16814 (N_16814,N_15862,N_16091);
nand U16815 (N_16815,N_16386,N_16746);
or U16816 (N_16816,N_16000,N_15610);
xnor U16817 (N_16817,N_16364,N_15697);
or U16818 (N_16818,N_16457,N_15724);
nor U16819 (N_16819,N_15674,N_16096);
nor U16820 (N_16820,N_15785,N_15878);
or U16821 (N_16821,N_16192,N_16034);
nand U16822 (N_16822,N_15665,N_15608);
nand U16823 (N_16823,N_15846,N_15755);
or U16824 (N_16824,N_16456,N_16638);
nand U16825 (N_16825,N_16058,N_15901);
or U16826 (N_16826,N_16751,N_16658);
nor U16827 (N_16827,N_16724,N_16084);
or U16828 (N_16828,N_16561,N_15938);
and U16829 (N_16829,N_16042,N_16418);
nor U16830 (N_16830,N_15658,N_16774);
nor U16831 (N_16831,N_16283,N_16320);
and U16832 (N_16832,N_16702,N_16708);
xnor U16833 (N_16833,N_16552,N_16621);
and U16834 (N_16834,N_16780,N_16723);
or U16835 (N_16835,N_16009,N_15981);
and U16836 (N_16836,N_16741,N_15640);
nand U16837 (N_16837,N_16228,N_16424);
or U16838 (N_16838,N_15974,N_15836);
nor U16839 (N_16839,N_16133,N_15638);
nand U16840 (N_16840,N_16215,N_16699);
and U16841 (N_16841,N_15692,N_16012);
nand U16842 (N_16842,N_16107,N_16593);
xor U16843 (N_16843,N_15968,N_16585);
xnor U16844 (N_16844,N_16503,N_15866);
or U16845 (N_16845,N_16415,N_15801);
and U16846 (N_16846,N_16794,N_16470);
xnor U16847 (N_16847,N_16580,N_16261);
or U16848 (N_16848,N_16278,N_16485);
nand U16849 (N_16849,N_16006,N_16553);
or U16850 (N_16850,N_16686,N_15813);
nand U16851 (N_16851,N_16035,N_16608);
nor U16852 (N_16852,N_15997,N_15934);
nor U16853 (N_16853,N_15954,N_15988);
and U16854 (N_16854,N_15677,N_16538);
xor U16855 (N_16855,N_15718,N_16212);
nand U16856 (N_16856,N_16607,N_16116);
nor U16857 (N_16857,N_15906,N_16443);
nand U16858 (N_16858,N_16003,N_15935);
xor U16859 (N_16859,N_15826,N_16155);
or U16860 (N_16860,N_15855,N_15942);
and U16861 (N_16861,N_15780,N_15920);
nand U16862 (N_16862,N_16326,N_16557);
or U16863 (N_16863,N_15945,N_16771);
or U16864 (N_16864,N_15991,N_15840);
nand U16865 (N_16865,N_15940,N_16214);
and U16866 (N_16866,N_16233,N_15871);
nand U16867 (N_16867,N_16772,N_15965);
nor U16868 (N_16868,N_16371,N_15772);
and U16869 (N_16869,N_16288,N_16730);
nor U16870 (N_16870,N_16700,N_15802);
xor U16871 (N_16871,N_16584,N_16394);
xnor U16872 (N_16872,N_15881,N_16193);
or U16873 (N_16873,N_16019,N_16799);
nand U16874 (N_16874,N_16509,N_16747);
xnor U16875 (N_16875,N_15725,N_15984);
nor U16876 (N_16876,N_16671,N_16138);
nor U16877 (N_16877,N_16707,N_15687);
or U16878 (N_16878,N_16762,N_16732);
xnor U16879 (N_16879,N_16798,N_16115);
nor U16880 (N_16880,N_15971,N_15660);
xnor U16881 (N_16881,N_15821,N_16211);
nor U16882 (N_16882,N_16651,N_16646);
xnor U16883 (N_16883,N_15627,N_15734);
nor U16884 (N_16884,N_15927,N_15619);
xnor U16885 (N_16885,N_15824,N_15955);
or U16886 (N_16886,N_16525,N_16567);
nor U16887 (N_16887,N_15653,N_16160);
and U16888 (N_16888,N_16491,N_15745);
and U16889 (N_16889,N_15913,N_16347);
nand U16890 (N_16890,N_16372,N_15931);
and U16891 (N_16891,N_16033,N_15889);
xnor U16892 (N_16892,N_16776,N_15728);
xor U16893 (N_16893,N_16273,N_16360);
nand U16894 (N_16894,N_16626,N_16257);
or U16895 (N_16895,N_16264,N_15979);
and U16896 (N_16896,N_15649,N_15962);
xnor U16897 (N_16897,N_16170,N_15973);
nand U16898 (N_16898,N_15750,N_16588);
xnor U16899 (N_16899,N_16382,N_16606);
or U16900 (N_16900,N_16677,N_15630);
nor U16901 (N_16901,N_16186,N_16477);
and U16902 (N_16902,N_15647,N_16059);
or U16903 (N_16903,N_16426,N_15770);
and U16904 (N_16904,N_16691,N_16025);
xor U16905 (N_16905,N_16715,N_15939);
or U16906 (N_16906,N_16539,N_16290);
nor U16907 (N_16907,N_16670,N_15694);
nand U16908 (N_16908,N_16250,N_15903);
nand U16909 (N_16909,N_16359,N_16341);
or U16910 (N_16910,N_16594,N_16452);
nor U16911 (N_16911,N_16647,N_15835);
xor U16912 (N_16912,N_16111,N_16472);
nand U16913 (N_16913,N_15646,N_16163);
and U16914 (N_16914,N_15675,N_15684);
and U16915 (N_16915,N_16450,N_16230);
nor U16916 (N_16916,N_15676,N_15875);
nor U16917 (N_16917,N_16411,N_15621);
and U16918 (N_16918,N_15663,N_16395);
nor U16919 (N_16919,N_15966,N_15877);
nand U16920 (N_16920,N_16239,N_16024);
or U16921 (N_16921,N_15898,N_15696);
and U16922 (N_16922,N_16796,N_15615);
nand U16923 (N_16923,N_15870,N_16196);
nand U16924 (N_16924,N_16660,N_15868);
and U16925 (N_16925,N_16641,N_16259);
nor U16926 (N_16926,N_16602,N_16792);
nand U16927 (N_16927,N_16507,N_16650);
nor U16928 (N_16928,N_15648,N_15672);
or U16929 (N_16929,N_16582,N_16758);
nand U16930 (N_16930,N_16184,N_15683);
or U16931 (N_16931,N_16156,N_15768);
xnor U16932 (N_16932,N_16536,N_15890);
xor U16933 (N_16933,N_16224,N_16225);
xor U16934 (N_16934,N_15944,N_15720);
nor U16935 (N_16935,N_16078,N_16644);
nand U16936 (N_16936,N_16174,N_15776);
and U16937 (N_16937,N_16044,N_16639);
and U16938 (N_16938,N_16094,N_15668);
or U16939 (N_16939,N_15798,N_15831);
xor U16940 (N_16940,N_16194,N_15618);
or U16941 (N_16941,N_16322,N_15716);
nand U16942 (N_16942,N_15787,N_16559);
and U16943 (N_16943,N_16243,N_15743);
and U16944 (N_16944,N_16581,N_16504);
nand U16945 (N_16945,N_16047,N_16248);
xnor U16946 (N_16946,N_16342,N_16759);
and U16947 (N_16947,N_15602,N_16343);
nand U16948 (N_16948,N_16054,N_16770);
xnor U16949 (N_16949,N_15644,N_15709);
nand U16950 (N_16950,N_16124,N_16517);
nand U16951 (N_16951,N_16253,N_16101);
nand U16952 (N_16952,N_16516,N_16281);
and U16953 (N_16953,N_15867,N_15751);
nand U16954 (N_16954,N_16268,N_16181);
nand U16955 (N_16955,N_15839,N_16512);
and U16956 (N_16956,N_16161,N_15695);
and U16957 (N_16957,N_16591,N_16396);
nand U16958 (N_16958,N_16018,N_16483);
xnor U16959 (N_16959,N_16313,N_16595);
xnor U16960 (N_16960,N_16766,N_16449);
nor U16961 (N_16961,N_16179,N_16688);
xor U16962 (N_16962,N_16332,N_15657);
or U16963 (N_16963,N_15722,N_15784);
or U16964 (N_16964,N_16030,N_16502);
xnor U16965 (N_16965,N_15852,N_15742);
xor U16966 (N_16966,N_15698,N_16398);
and U16967 (N_16967,N_16305,N_16383);
or U16968 (N_16968,N_16307,N_15995);
or U16969 (N_16969,N_16755,N_16468);
nand U16970 (N_16970,N_15727,N_16496);
or U16971 (N_16971,N_15858,N_16541);
nor U16972 (N_16972,N_16514,N_15807);
xnor U16973 (N_16973,N_16570,N_16284);
nor U16974 (N_16974,N_16031,N_15705);
and U16975 (N_16975,N_16719,N_15740);
nand U16976 (N_16976,N_15959,N_16569);
and U16977 (N_16977,N_15902,N_16165);
xor U16978 (N_16978,N_16540,N_16123);
and U16979 (N_16979,N_16579,N_16331);
and U16980 (N_16980,N_16462,N_16684);
or U16981 (N_16981,N_16717,N_16108);
nand U16982 (N_16982,N_16350,N_16414);
or U16983 (N_16983,N_16368,N_15983);
or U16984 (N_16984,N_16037,N_16282);
xor U16985 (N_16985,N_16401,N_16038);
and U16986 (N_16986,N_16451,N_16036);
or U16987 (N_16987,N_16546,N_15941);
and U16988 (N_16988,N_15690,N_16324);
and U16989 (N_16989,N_16397,N_16549);
and U16990 (N_16990,N_15633,N_16637);
or U16991 (N_16991,N_16564,N_16623);
nand U16992 (N_16992,N_16010,N_15681);
or U16993 (N_16993,N_16141,N_16045);
nor U16994 (N_16994,N_16506,N_16576);
nand U16995 (N_16995,N_16146,N_16262);
xnor U16996 (N_16996,N_16029,N_16014);
or U16997 (N_16997,N_16187,N_15884);
xor U16998 (N_16998,N_16654,N_15880);
nor U16999 (N_16999,N_16222,N_16448);
xor U17000 (N_17000,N_15822,N_15857);
nand U17001 (N_17001,N_15703,N_16442);
nand U17002 (N_17002,N_15930,N_16176);
nand U17003 (N_17003,N_16587,N_16548);
or U17004 (N_17004,N_15830,N_16466);
nor U17005 (N_17005,N_16032,N_15631);
or U17006 (N_17006,N_16475,N_15818);
or U17007 (N_17007,N_16316,N_16189);
or U17008 (N_17008,N_16596,N_15872);
nand U17009 (N_17009,N_16458,N_16522);
nand U17010 (N_17010,N_16227,N_16765);
xnor U17011 (N_17011,N_16797,N_15629);
nand U17012 (N_17012,N_15928,N_16612);
or U17013 (N_17013,N_16279,N_16002);
nand U17014 (N_17014,N_16731,N_16270);
and U17015 (N_17015,N_16642,N_16735);
nand U17016 (N_17016,N_15869,N_16739);
nand U17017 (N_17017,N_16445,N_15736);
nor U17018 (N_17018,N_15961,N_16526);
nor U17019 (N_17019,N_15730,N_16043);
xor U17020 (N_17020,N_15970,N_16742);
or U17021 (N_17021,N_16256,N_16131);
and U17022 (N_17022,N_16530,N_16791);
and U17023 (N_17023,N_16781,N_16550);
xor U17024 (N_17024,N_15978,N_16387);
xnor U17025 (N_17025,N_16510,N_16221);
xor U17026 (N_17026,N_15827,N_15686);
or U17027 (N_17027,N_16242,N_16345);
nor U17028 (N_17028,N_16464,N_16631);
xnor U17029 (N_17029,N_15958,N_16306);
and U17030 (N_17030,N_15650,N_16653);
xor U17031 (N_17031,N_16761,N_16154);
or U17032 (N_17032,N_16488,N_15760);
nand U17033 (N_17033,N_16754,N_16681);
nor U17034 (N_17034,N_16407,N_16235);
or U17035 (N_17035,N_15765,N_16710);
and U17036 (N_17036,N_15773,N_15833);
xnor U17037 (N_17037,N_16238,N_15605);
nand U17038 (N_17038,N_15609,N_16469);
nor U17039 (N_17039,N_16286,N_16321);
nor U17040 (N_17040,N_16056,N_16244);
and U17041 (N_17041,N_16158,N_16459);
nand U17042 (N_17042,N_15623,N_16075);
xnor U17043 (N_17043,N_16404,N_16447);
and U17044 (N_17044,N_16537,N_16060);
xnor U17045 (N_17045,N_16562,N_16365);
and U17046 (N_17046,N_16611,N_16366);
or U17047 (N_17047,N_15808,N_15712);
nor U17048 (N_17048,N_16634,N_16391);
and U17049 (N_17049,N_16087,N_15996);
nor U17050 (N_17050,N_16640,N_15829);
and U17051 (N_17051,N_16431,N_16790);
xnor U17052 (N_17052,N_16783,N_16666);
xnor U17053 (N_17053,N_15620,N_16388);
and U17054 (N_17054,N_16476,N_16066);
xor U17055 (N_17055,N_15735,N_16337);
nor U17056 (N_17056,N_15899,N_16773);
nand U17057 (N_17057,N_16129,N_16272);
or U17058 (N_17058,N_16501,N_15799);
xnor U17059 (N_17059,N_16628,N_16218);
nor U17060 (N_17060,N_16663,N_16263);
and U17061 (N_17061,N_15754,N_16197);
nand U17062 (N_17062,N_15656,N_16705);
nand U17063 (N_17063,N_15910,N_16097);
nand U17064 (N_17064,N_16455,N_15753);
nor U17065 (N_17065,N_16474,N_15662);
nor U17066 (N_17066,N_16775,N_16441);
xor U17067 (N_17067,N_16020,N_16005);
and U17068 (N_17068,N_15659,N_16277);
or U17069 (N_17069,N_16669,N_16199);
xor U17070 (N_17070,N_16374,N_16667);
nand U17071 (N_17071,N_16620,N_15924);
nand U17072 (N_17072,N_16711,N_16609);
and U17073 (N_17073,N_15601,N_15731);
and U17074 (N_17074,N_16757,N_16309);
or U17075 (N_17075,N_16590,N_16168);
and U17076 (N_17076,N_16276,N_16150);
nand U17077 (N_17077,N_16098,N_16393);
nor U17078 (N_17078,N_16563,N_16727);
xor U17079 (N_17079,N_16499,N_16422);
and U17080 (N_17080,N_16627,N_16004);
nor U17081 (N_17081,N_16247,N_16678);
nor U17082 (N_17082,N_16648,N_16266);
or U17083 (N_17083,N_16258,N_16318);
nand U17084 (N_17084,N_16714,N_16203);
or U17085 (N_17085,N_15849,N_16057);
nand U17086 (N_17086,N_16427,N_16110);
xor U17087 (N_17087,N_16236,N_16375);
nand U17088 (N_17088,N_16643,N_15987);
and U17089 (N_17089,N_16310,N_16055);
or U17090 (N_17090,N_16302,N_16265);
or U17091 (N_17091,N_16473,N_15732);
nor U17092 (N_17092,N_16399,N_16339);
and U17093 (N_17093,N_16148,N_16763);
nor U17094 (N_17094,N_15985,N_16786);
xor U17095 (N_17095,N_16436,N_16430);
nor U17096 (N_17096,N_16298,N_15815);
nand U17097 (N_17097,N_16409,N_16021);
and U17098 (N_17098,N_16208,N_16064);
or U17099 (N_17099,N_16068,N_16049);
and U17100 (N_17100,N_15767,N_16597);
xor U17101 (N_17101,N_15972,N_15963);
and U17102 (N_17102,N_15682,N_16721);
nand U17103 (N_17103,N_15957,N_15882);
nand U17104 (N_17104,N_16729,N_15664);
nand U17105 (N_17105,N_16695,N_16467);
or U17106 (N_17106,N_16789,N_16665);
and U17107 (N_17107,N_16303,N_16768);
and U17108 (N_17108,N_15752,N_16479);
and U17109 (N_17109,N_15741,N_16376);
or U17110 (N_17110,N_16112,N_15786);
and U17111 (N_17111,N_16269,N_16334);
nand U17112 (N_17112,N_16385,N_15655);
or U17113 (N_17113,N_16092,N_15774);
nand U17114 (N_17114,N_16172,N_16795);
or U17115 (N_17115,N_16493,N_16692);
and U17116 (N_17116,N_16128,N_16190);
and U17117 (N_17117,N_16392,N_16209);
nor U17118 (N_17118,N_16175,N_16592);
nand U17119 (N_17119,N_16102,N_16687);
or U17120 (N_17120,N_16389,N_16103);
xor U17121 (N_17121,N_15810,N_15853);
or U17122 (N_17122,N_16171,N_15834);
and U17123 (N_17123,N_15989,N_16565);
nor U17124 (N_17124,N_16413,N_16716);
and U17125 (N_17125,N_15980,N_16142);
and U17126 (N_17126,N_16130,N_16039);
xnor U17127 (N_17127,N_16061,N_16652);
nand U17128 (N_17128,N_16167,N_15952);
nor U17129 (N_17129,N_15782,N_16712);
xnor U17130 (N_17130,N_16555,N_16252);
or U17131 (N_17131,N_15729,N_16500);
nand U17132 (N_17132,N_16577,N_16271);
nor U17133 (N_17133,N_16603,N_15789);
xor U17134 (N_17134,N_15850,N_16071);
or U17135 (N_17135,N_16073,N_16674);
nor U17136 (N_17136,N_15926,N_16050);
nand U17137 (N_17137,N_15763,N_16315);
and U17138 (N_17138,N_16114,N_16545);
nand U17139 (N_17139,N_15886,N_15993);
xnor U17140 (N_17140,N_16680,N_16140);
nand U17141 (N_17141,N_15737,N_16319);
and U17142 (N_17142,N_16173,N_16764);
nand U17143 (N_17143,N_15713,N_15887);
or U17144 (N_17144,N_16157,N_16330);
nand U17145 (N_17145,N_16788,N_16072);
xnor U17146 (N_17146,N_15929,N_16017);
or U17147 (N_17147,N_16351,N_16361);
xor U17148 (N_17148,N_16617,N_16294);
xnor U17149 (N_17149,N_16067,N_15990);
and U17150 (N_17150,N_16080,N_16785);
xor U17151 (N_17151,N_15689,N_15812);
or U17152 (N_17152,N_16198,N_15678);
nor U17153 (N_17153,N_15645,N_16234);
nand U17154 (N_17154,N_15856,N_16346);
xor U17155 (N_17155,N_16159,N_15706);
xnor U17156 (N_17156,N_15794,N_16575);
and U17157 (N_17157,N_16356,N_16125);
nor U17158 (N_17158,N_15748,N_15795);
xor U17159 (N_17159,N_16106,N_16086);
xor U17160 (N_17160,N_16551,N_16529);
and U17161 (N_17161,N_16210,N_16169);
nor U17162 (N_17162,N_16293,N_16335);
and U17163 (N_17163,N_16289,N_16231);
and U17164 (N_17164,N_15876,N_15873);
nor U17165 (N_17165,N_15777,N_16656);
and U17166 (N_17166,N_15986,N_15814);
xnor U17167 (N_17167,N_16241,N_16513);
or U17168 (N_17168,N_15998,N_15845);
and U17169 (N_17169,N_16245,N_16554);
nor U17170 (N_17170,N_15838,N_16301);
and U17171 (N_17171,N_16178,N_16327);
xnor U17172 (N_17172,N_16463,N_16177);
or U17173 (N_17173,N_16357,N_16527);
nor U17174 (N_17174,N_15937,N_16354);
and U17175 (N_17175,N_16377,N_15783);
and U17176 (N_17176,N_16544,N_16438);
or U17177 (N_17177,N_16440,N_16494);
nand U17178 (N_17178,N_16207,N_16323);
xor U17179 (N_17179,N_16149,N_16405);
xnor U17180 (N_17180,N_16752,N_16249);
nor U17181 (N_17181,N_15702,N_16119);
nand U17182 (N_17182,N_16725,N_16524);
and U17183 (N_17183,N_16425,N_15685);
nor U17184 (N_17184,N_16137,N_15628);
xnor U17185 (N_17185,N_15809,N_15922);
xor U17186 (N_17186,N_16625,N_16750);
and U17187 (N_17187,N_15847,N_16077);
and U17188 (N_17188,N_16132,N_16062);
and U17189 (N_17189,N_16523,N_15953);
xor U17190 (N_17190,N_16206,N_16793);
nor U17191 (N_17191,N_16205,N_16299);
nor U17192 (N_17192,N_15949,N_16543);
and U17193 (N_17193,N_15932,N_15891);
or U17194 (N_17194,N_15766,N_16344);
nand U17195 (N_17195,N_16104,N_16201);
nand U17196 (N_17196,N_16349,N_16421);
nand U17197 (N_17197,N_16498,N_16753);
nand U17198 (N_17198,N_15956,N_16661);
nand U17199 (N_17199,N_16685,N_15607);
nor U17200 (N_17200,N_15769,N_15711);
or U17201 (N_17201,N_16088,N_16260);
and U17202 (N_17202,N_16417,N_16492);
and U17203 (N_17203,N_16074,N_16694);
and U17204 (N_17204,N_16013,N_15747);
and U17205 (N_17205,N_15600,N_15762);
or U17206 (N_17206,N_16726,N_16744);
nor U17207 (N_17207,N_15761,N_15710);
nor U17208 (N_17208,N_16100,N_16733);
nor U17209 (N_17209,N_16622,N_16696);
nor U17210 (N_17210,N_15919,N_16676);
xnor U17211 (N_17211,N_16518,N_15933);
xnor U17212 (N_17212,N_16251,N_16329);
and U17213 (N_17213,N_16028,N_16615);
xnor U17214 (N_17214,N_16704,N_16402);
and U17215 (N_17215,N_15885,N_16701);
nor U17216 (N_17216,N_16011,N_15943);
xnor U17217 (N_17217,N_16481,N_15791);
or U17218 (N_17218,N_15757,N_15612);
nand U17219 (N_17219,N_15723,N_16535);
nand U17220 (N_17220,N_16046,N_15708);
nand U17221 (N_17221,N_15851,N_16560);
and U17222 (N_17222,N_16353,N_15946);
nor U17223 (N_17223,N_16079,N_16325);
xnor U17224 (N_17224,N_15921,N_16122);
nand U17225 (N_17225,N_16437,N_16403);
or U17226 (N_17226,N_16740,N_15604);
xnor U17227 (N_17227,N_15925,N_15670);
or U17228 (N_17228,N_16048,N_16380);
nand U17229 (N_17229,N_16683,N_16520);
nor U17230 (N_17230,N_16127,N_16583);
xnor U17231 (N_17231,N_16533,N_16370);
or U17232 (N_17232,N_15666,N_15739);
and U17233 (N_17233,N_16410,N_15775);
or U17234 (N_17234,N_16202,N_16610);
nor U17235 (N_17235,N_16490,N_16182);
or U17236 (N_17236,N_15800,N_16400);
and U17237 (N_17237,N_15843,N_16573);
or U17238 (N_17238,N_16777,N_16624);
or U17239 (N_17239,N_16429,N_16240);
xor U17240 (N_17240,N_15842,N_16428);
or U17241 (N_17241,N_15749,N_15624);
nor U17242 (N_17242,N_16675,N_16317);
or U17243 (N_17243,N_16053,N_16778);
or U17244 (N_17244,N_16531,N_16664);
or U17245 (N_17245,N_15680,N_16355);
nand U17246 (N_17246,N_16668,N_16571);
nor U17247 (N_17247,N_16558,N_16782);
and U17248 (N_17248,N_16287,N_16362);
or U17249 (N_17249,N_16120,N_16027);
and U17250 (N_17250,N_15781,N_15726);
or U17251 (N_17251,N_16649,N_16619);
xnor U17252 (N_17252,N_15643,N_15915);
or U17253 (N_17253,N_15859,N_16614);
nor U17254 (N_17254,N_15744,N_15976);
nand U17255 (N_17255,N_16589,N_15790);
xor U17256 (N_17256,N_16254,N_15948);
nor U17257 (N_17257,N_16166,N_16022);
nand U17258 (N_17258,N_15917,N_16001);
and U17259 (N_17259,N_16336,N_16153);
xor U17260 (N_17260,N_16226,N_16348);
and U17261 (N_17261,N_15667,N_16291);
and U17262 (N_17262,N_16586,N_16358);
nand U17263 (N_17263,N_15806,N_15721);
nor U17264 (N_17264,N_16180,N_16420);
xor U17265 (N_17265,N_16406,N_16734);
and U17266 (N_17266,N_16390,N_16749);
or U17267 (N_17267,N_16135,N_16433);
and U17268 (N_17268,N_16352,N_16508);
or U17269 (N_17269,N_15805,N_16635);
or U17270 (N_17270,N_15918,N_16534);
nand U17271 (N_17271,N_15613,N_16367);
xor U17272 (N_17272,N_16113,N_16662);
xor U17273 (N_17273,N_16378,N_16412);
nor U17274 (N_17274,N_15854,N_16672);
or U17275 (N_17275,N_16041,N_16089);
nor U17276 (N_17276,N_16090,N_15994);
xor U17277 (N_17277,N_16340,N_15778);
nor U17278 (N_17278,N_16237,N_16599);
xor U17279 (N_17279,N_15820,N_15879);
and U17280 (N_17280,N_16743,N_15671);
or U17281 (N_17281,N_16690,N_16216);
xnor U17282 (N_17282,N_16478,N_15892);
nor U17283 (N_17283,N_16134,N_15796);
or U17284 (N_17284,N_16052,N_16748);
nand U17285 (N_17285,N_16162,N_16183);
and U17286 (N_17286,N_16292,N_16188);
nor U17287 (N_17287,N_16446,N_16121);
nand U17288 (N_17288,N_16274,N_15688);
nor U17289 (N_17289,N_15916,N_15947);
nor U17290 (N_17290,N_15622,N_16435);
nor U17291 (N_17291,N_16408,N_15764);
or U17292 (N_17292,N_15654,N_16143);
xnor U17293 (N_17293,N_15639,N_16657);
nor U17294 (N_17294,N_16720,N_16136);
nand U17295 (N_17295,N_16126,N_15975);
or U17296 (N_17296,N_16693,N_15617);
or U17297 (N_17297,N_16416,N_16713);
or U17298 (N_17298,N_16745,N_15616);
nand U17299 (N_17299,N_15900,N_16023);
or U17300 (N_17300,N_15611,N_15714);
or U17301 (N_17301,N_15825,N_15950);
nand U17302 (N_17302,N_15788,N_16363);
or U17303 (N_17303,N_15992,N_16655);
and U17304 (N_17304,N_16480,N_15883);
nand U17305 (N_17305,N_16673,N_15625);
nand U17306 (N_17306,N_16384,N_16519);
nor U17307 (N_17307,N_16679,N_16051);
and U17308 (N_17308,N_16118,N_16026);
or U17309 (N_17309,N_15977,N_16152);
and U17310 (N_17310,N_15603,N_16373);
xor U17311 (N_17311,N_15969,N_15832);
nor U17312 (N_17312,N_16093,N_16454);
and U17313 (N_17313,N_15923,N_16015);
and U17314 (N_17314,N_15909,N_16109);
nor U17315 (N_17315,N_16703,N_15816);
and U17316 (N_17316,N_16486,N_16311);
and U17317 (N_17317,N_16697,N_16728);
nand U17318 (N_17318,N_16369,N_16495);
and U17319 (N_17319,N_16471,N_16085);
nand U17320 (N_17320,N_16636,N_16784);
or U17321 (N_17321,N_16423,N_15715);
or U17322 (N_17322,N_15905,N_15960);
nor U17323 (N_17323,N_15811,N_16105);
nand U17324 (N_17324,N_16285,N_16219);
xor U17325 (N_17325,N_16223,N_15865);
xor U17326 (N_17326,N_16779,N_15651);
nand U17327 (N_17327,N_16419,N_16333);
and U17328 (N_17328,N_16645,N_15828);
nand U17329 (N_17329,N_15691,N_16280);
nand U17330 (N_17330,N_15999,N_16613);
nand U17331 (N_17331,N_15626,N_15642);
xnor U17332 (N_17332,N_15634,N_16381);
nand U17333 (N_17333,N_16547,N_16542);
xnor U17334 (N_17334,N_16296,N_16632);
xnor U17335 (N_17335,N_16787,N_16633);
nand U17336 (N_17336,N_15637,N_16300);
nor U17337 (N_17337,N_16338,N_16016);
or U17338 (N_17338,N_16081,N_16432);
and U17339 (N_17339,N_16497,N_15874);
and U17340 (N_17340,N_16083,N_16144);
and U17341 (N_17341,N_16600,N_16528);
nand U17342 (N_17342,N_15888,N_15817);
nor U17343 (N_17343,N_16145,N_16722);
and U17344 (N_17344,N_15914,N_15841);
or U17345 (N_17345,N_16515,N_15951);
and U17346 (N_17346,N_16065,N_16439);
or U17347 (N_17347,N_15606,N_15717);
nor U17348 (N_17348,N_15700,N_16737);
nand U17349 (N_17349,N_15982,N_16618);
nor U17350 (N_17350,N_16164,N_16040);
nand U17351 (N_17351,N_15635,N_15699);
or U17352 (N_17352,N_16605,N_16220);
xor U17353 (N_17353,N_16007,N_15967);
nor U17354 (N_17354,N_15719,N_15860);
and U17355 (N_17355,N_16706,N_15758);
or U17356 (N_17356,N_15803,N_15912);
xnor U17357 (N_17357,N_16568,N_16195);
or U17358 (N_17358,N_16185,N_16328);
and U17359 (N_17359,N_16246,N_16574);
and U17360 (N_17360,N_16275,N_15804);
and U17361 (N_17361,N_16314,N_15864);
or U17362 (N_17362,N_16295,N_16709);
nor U17363 (N_17363,N_15896,N_16117);
or U17364 (N_17364,N_15746,N_16487);
nor U17365 (N_17365,N_15701,N_16736);
or U17366 (N_17366,N_15797,N_16521);
nor U17367 (N_17367,N_16698,N_16598);
nand U17368 (N_17368,N_16267,N_16312);
nor U17369 (N_17369,N_16760,N_15897);
nor U17370 (N_17370,N_15792,N_16147);
and U17371 (N_17371,N_16738,N_16489);
or U17372 (N_17372,N_16659,N_15848);
and U17373 (N_17373,N_16484,N_15793);
and U17374 (N_17374,N_15893,N_15652);
nor U17375 (N_17375,N_15738,N_15661);
nand U17376 (N_17376,N_16601,N_16511);
nand U17377 (N_17377,N_16082,N_16232);
nor U17378 (N_17378,N_16255,N_16604);
and U17379 (N_17379,N_15641,N_16756);
nor U17380 (N_17380,N_16308,N_16482);
nor U17381 (N_17381,N_16505,N_16689);
or U17382 (N_17382,N_15759,N_16095);
or U17383 (N_17383,N_16070,N_15756);
and U17384 (N_17384,N_16566,N_15861);
xnor U17385 (N_17385,N_15908,N_16682);
or U17386 (N_17386,N_16460,N_16076);
or U17387 (N_17387,N_16578,N_16444);
nor U17388 (N_17388,N_16379,N_16532);
nor U17389 (N_17389,N_16204,N_15679);
nand U17390 (N_17390,N_15707,N_15936);
nand U17391 (N_17391,N_16718,N_16465);
nand U17392 (N_17392,N_15863,N_16461);
nor U17393 (N_17393,N_15907,N_15693);
or U17394 (N_17394,N_16191,N_16616);
and U17395 (N_17395,N_16099,N_16200);
xnor U17396 (N_17396,N_16629,N_15904);
nand U17397 (N_17397,N_15895,N_15614);
and U17398 (N_17398,N_15673,N_15669);
xor U17399 (N_17399,N_15844,N_15733);
xor U17400 (N_17400,N_16367,N_16385);
and U17401 (N_17401,N_16660,N_15850);
xor U17402 (N_17402,N_16424,N_16402);
nand U17403 (N_17403,N_16123,N_16575);
xor U17404 (N_17404,N_15985,N_15772);
nor U17405 (N_17405,N_16401,N_16230);
and U17406 (N_17406,N_15854,N_15752);
xnor U17407 (N_17407,N_15795,N_16609);
and U17408 (N_17408,N_16091,N_16558);
nand U17409 (N_17409,N_15990,N_16527);
nand U17410 (N_17410,N_15979,N_16636);
and U17411 (N_17411,N_16451,N_16546);
or U17412 (N_17412,N_16326,N_16169);
and U17413 (N_17413,N_16387,N_16606);
xnor U17414 (N_17414,N_16479,N_15819);
or U17415 (N_17415,N_16105,N_16084);
xor U17416 (N_17416,N_16661,N_15709);
and U17417 (N_17417,N_16663,N_15885);
or U17418 (N_17418,N_15918,N_16659);
nor U17419 (N_17419,N_15687,N_15643);
and U17420 (N_17420,N_16552,N_16195);
nor U17421 (N_17421,N_15859,N_16188);
and U17422 (N_17422,N_16132,N_16225);
and U17423 (N_17423,N_15683,N_16207);
and U17424 (N_17424,N_16745,N_15816);
and U17425 (N_17425,N_16038,N_15602);
xnor U17426 (N_17426,N_16372,N_16040);
and U17427 (N_17427,N_16499,N_15680);
and U17428 (N_17428,N_16062,N_15681);
xor U17429 (N_17429,N_15787,N_15901);
and U17430 (N_17430,N_15798,N_16282);
or U17431 (N_17431,N_15979,N_15956);
nor U17432 (N_17432,N_15762,N_15643);
nand U17433 (N_17433,N_16355,N_15907);
and U17434 (N_17434,N_16329,N_16153);
and U17435 (N_17435,N_16466,N_16535);
or U17436 (N_17436,N_16334,N_16544);
and U17437 (N_17437,N_16785,N_15819);
nand U17438 (N_17438,N_15620,N_15848);
and U17439 (N_17439,N_15613,N_16293);
and U17440 (N_17440,N_16516,N_16702);
and U17441 (N_17441,N_16282,N_16680);
or U17442 (N_17442,N_16681,N_16387);
and U17443 (N_17443,N_16648,N_16079);
xnor U17444 (N_17444,N_15974,N_16049);
nor U17445 (N_17445,N_16422,N_16557);
nand U17446 (N_17446,N_16570,N_16048);
and U17447 (N_17447,N_15869,N_16401);
and U17448 (N_17448,N_16501,N_16707);
and U17449 (N_17449,N_16047,N_16230);
nand U17450 (N_17450,N_16048,N_16004);
and U17451 (N_17451,N_16181,N_16144);
nand U17452 (N_17452,N_15635,N_15821);
xnor U17453 (N_17453,N_16499,N_16675);
nor U17454 (N_17454,N_16201,N_16406);
nand U17455 (N_17455,N_16409,N_15948);
or U17456 (N_17456,N_16601,N_16666);
and U17457 (N_17457,N_15802,N_16007);
xnor U17458 (N_17458,N_15646,N_16472);
xor U17459 (N_17459,N_16771,N_15898);
and U17460 (N_17460,N_15831,N_16346);
nor U17461 (N_17461,N_16538,N_15992);
xor U17462 (N_17462,N_16670,N_15609);
xnor U17463 (N_17463,N_15719,N_16535);
nand U17464 (N_17464,N_16140,N_16018);
or U17465 (N_17465,N_16690,N_15723);
nand U17466 (N_17466,N_15815,N_15816);
and U17467 (N_17467,N_15651,N_16108);
nand U17468 (N_17468,N_16660,N_16132);
and U17469 (N_17469,N_15944,N_16366);
nor U17470 (N_17470,N_15938,N_16096);
nand U17471 (N_17471,N_16022,N_16787);
xor U17472 (N_17472,N_15870,N_15660);
xnor U17473 (N_17473,N_16756,N_15859);
xor U17474 (N_17474,N_16053,N_16508);
xnor U17475 (N_17475,N_16621,N_16017);
nor U17476 (N_17476,N_15659,N_16320);
xor U17477 (N_17477,N_15618,N_16348);
xor U17478 (N_17478,N_16540,N_16125);
and U17479 (N_17479,N_15664,N_16604);
or U17480 (N_17480,N_16094,N_16256);
or U17481 (N_17481,N_16191,N_16322);
nor U17482 (N_17482,N_16392,N_15831);
nor U17483 (N_17483,N_16586,N_15872);
or U17484 (N_17484,N_16531,N_16075);
nand U17485 (N_17485,N_16643,N_16275);
and U17486 (N_17486,N_16569,N_16767);
nor U17487 (N_17487,N_16794,N_16433);
and U17488 (N_17488,N_15863,N_16097);
and U17489 (N_17489,N_16202,N_16412);
nor U17490 (N_17490,N_16627,N_15792);
nand U17491 (N_17491,N_16128,N_16733);
xor U17492 (N_17492,N_16247,N_15799);
xor U17493 (N_17493,N_16332,N_15866);
nand U17494 (N_17494,N_16438,N_16256);
nand U17495 (N_17495,N_15939,N_16210);
nor U17496 (N_17496,N_15768,N_16706);
or U17497 (N_17497,N_15946,N_16577);
nand U17498 (N_17498,N_16036,N_16057);
xnor U17499 (N_17499,N_16133,N_15647);
or U17500 (N_17500,N_15706,N_16010);
and U17501 (N_17501,N_15687,N_15609);
nor U17502 (N_17502,N_16709,N_16178);
nor U17503 (N_17503,N_16444,N_16308);
or U17504 (N_17504,N_16242,N_16659);
or U17505 (N_17505,N_16111,N_16564);
or U17506 (N_17506,N_16545,N_16244);
and U17507 (N_17507,N_16639,N_16602);
nand U17508 (N_17508,N_16080,N_16473);
nor U17509 (N_17509,N_16501,N_16265);
nor U17510 (N_17510,N_16438,N_15863);
and U17511 (N_17511,N_15949,N_16347);
nor U17512 (N_17512,N_15923,N_16777);
xnor U17513 (N_17513,N_16741,N_15943);
and U17514 (N_17514,N_16771,N_16331);
xnor U17515 (N_17515,N_16405,N_16552);
or U17516 (N_17516,N_16482,N_16137);
xor U17517 (N_17517,N_16033,N_16412);
or U17518 (N_17518,N_16785,N_16099);
nor U17519 (N_17519,N_16537,N_16444);
or U17520 (N_17520,N_15619,N_16468);
nor U17521 (N_17521,N_16795,N_16629);
and U17522 (N_17522,N_16093,N_15995);
and U17523 (N_17523,N_15789,N_16619);
and U17524 (N_17524,N_16723,N_16729);
or U17525 (N_17525,N_16214,N_16162);
nand U17526 (N_17526,N_16641,N_16112);
or U17527 (N_17527,N_16450,N_16550);
or U17528 (N_17528,N_15845,N_15907);
and U17529 (N_17529,N_15702,N_16702);
and U17530 (N_17530,N_16291,N_16253);
nor U17531 (N_17531,N_16749,N_15848);
or U17532 (N_17532,N_16105,N_15686);
or U17533 (N_17533,N_15900,N_16571);
nand U17534 (N_17534,N_16530,N_15833);
or U17535 (N_17535,N_15792,N_16558);
or U17536 (N_17536,N_16664,N_16618);
or U17537 (N_17537,N_16356,N_16127);
nor U17538 (N_17538,N_15862,N_16460);
xor U17539 (N_17539,N_16094,N_16317);
or U17540 (N_17540,N_15908,N_16239);
xnor U17541 (N_17541,N_16397,N_16106);
xnor U17542 (N_17542,N_16237,N_16277);
and U17543 (N_17543,N_16191,N_16000);
xor U17544 (N_17544,N_16124,N_16268);
or U17545 (N_17545,N_16550,N_16009);
nand U17546 (N_17546,N_16146,N_16588);
or U17547 (N_17547,N_16183,N_16475);
or U17548 (N_17548,N_15840,N_16251);
xnor U17549 (N_17549,N_16489,N_16613);
and U17550 (N_17550,N_16034,N_16238);
or U17551 (N_17551,N_15775,N_16218);
xnor U17552 (N_17552,N_15715,N_16746);
or U17553 (N_17553,N_15826,N_16622);
nor U17554 (N_17554,N_15870,N_15603);
xnor U17555 (N_17555,N_16109,N_16693);
and U17556 (N_17556,N_16450,N_15970);
nor U17557 (N_17557,N_16425,N_16739);
nor U17558 (N_17558,N_16560,N_16075);
xnor U17559 (N_17559,N_15962,N_16574);
nor U17560 (N_17560,N_16564,N_15830);
nor U17561 (N_17561,N_15782,N_16194);
and U17562 (N_17562,N_15628,N_15840);
nand U17563 (N_17563,N_16508,N_16198);
or U17564 (N_17564,N_16687,N_16685);
and U17565 (N_17565,N_16575,N_16609);
nand U17566 (N_17566,N_16381,N_16718);
xnor U17567 (N_17567,N_16077,N_16354);
and U17568 (N_17568,N_16697,N_15666);
or U17569 (N_17569,N_15890,N_16730);
or U17570 (N_17570,N_16719,N_16323);
or U17571 (N_17571,N_16205,N_16046);
nor U17572 (N_17572,N_16261,N_15784);
and U17573 (N_17573,N_15998,N_15723);
or U17574 (N_17574,N_16213,N_15648);
nand U17575 (N_17575,N_16429,N_16146);
or U17576 (N_17576,N_16780,N_16195);
or U17577 (N_17577,N_15738,N_15777);
nor U17578 (N_17578,N_15964,N_15751);
nand U17579 (N_17579,N_15969,N_16458);
or U17580 (N_17580,N_15693,N_16379);
nor U17581 (N_17581,N_16325,N_16744);
xor U17582 (N_17582,N_16787,N_16290);
or U17583 (N_17583,N_16065,N_15743);
and U17584 (N_17584,N_16631,N_15827);
xnor U17585 (N_17585,N_16558,N_16259);
or U17586 (N_17586,N_15708,N_16436);
nand U17587 (N_17587,N_16025,N_15648);
nand U17588 (N_17588,N_16407,N_16786);
nand U17589 (N_17589,N_16432,N_15792);
nand U17590 (N_17590,N_16063,N_16228);
nor U17591 (N_17591,N_16412,N_16699);
nor U17592 (N_17592,N_15801,N_15628);
xor U17593 (N_17593,N_15960,N_16089);
and U17594 (N_17594,N_16593,N_15863);
nand U17595 (N_17595,N_15768,N_16551);
and U17596 (N_17596,N_15974,N_16654);
nor U17597 (N_17597,N_15818,N_15928);
or U17598 (N_17598,N_16613,N_16779);
nand U17599 (N_17599,N_16242,N_16326);
nand U17600 (N_17600,N_16009,N_15889);
xnor U17601 (N_17601,N_15872,N_16799);
nand U17602 (N_17602,N_15605,N_16712);
nand U17603 (N_17603,N_15897,N_15861);
or U17604 (N_17604,N_16050,N_16148);
nand U17605 (N_17605,N_16194,N_15831);
xnor U17606 (N_17606,N_16726,N_15643);
and U17607 (N_17607,N_16065,N_16297);
nand U17608 (N_17608,N_16629,N_16623);
nor U17609 (N_17609,N_16282,N_15994);
nand U17610 (N_17610,N_16306,N_16783);
and U17611 (N_17611,N_16119,N_15751);
nor U17612 (N_17612,N_16195,N_15638);
xor U17613 (N_17613,N_16477,N_16068);
or U17614 (N_17614,N_16403,N_16197);
nand U17615 (N_17615,N_16530,N_15886);
xor U17616 (N_17616,N_16674,N_16306);
xnor U17617 (N_17617,N_15762,N_15736);
or U17618 (N_17618,N_15679,N_16210);
or U17619 (N_17619,N_16301,N_15886);
or U17620 (N_17620,N_16529,N_16133);
xnor U17621 (N_17621,N_16369,N_16450);
nand U17622 (N_17622,N_16793,N_15713);
nor U17623 (N_17623,N_16031,N_16022);
and U17624 (N_17624,N_15973,N_16413);
and U17625 (N_17625,N_16191,N_16309);
and U17626 (N_17626,N_16769,N_16192);
nor U17627 (N_17627,N_15663,N_16034);
and U17628 (N_17628,N_16763,N_15726);
nor U17629 (N_17629,N_16201,N_16362);
and U17630 (N_17630,N_16668,N_16629);
nor U17631 (N_17631,N_15930,N_15893);
and U17632 (N_17632,N_15783,N_16651);
nor U17633 (N_17633,N_16666,N_15841);
and U17634 (N_17634,N_16232,N_16615);
nor U17635 (N_17635,N_15992,N_16367);
or U17636 (N_17636,N_16511,N_15767);
xor U17637 (N_17637,N_16353,N_16134);
and U17638 (N_17638,N_16258,N_16783);
nand U17639 (N_17639,N_16752,N_16718);
nor U17640 (N_17640,N_15913,N_16176);
and U17641 (N_17641,N_15662,N_15617);
or U17642 (N_17642,N_16782,N_15633);
xnor U17643 (N_17643,N_15697,N_16660);
and U17644 (N_17644,N_15821,N_16136);
nand U17645 (N_17645,N_15757,N_16180);
or U17646 (N_17646,N_16491,N_16764);
xor U17647 (N_17647,N_16292,N_16555);
xnor U17648 (N_17648,N_16711,N_15789);
nand U17649 (N_17649,N_15884,N_16665);
nor U17650 (N_17650,N_16592,N_16499);
xor U17651 (N_17651,N_16450,N_16374);
xor U17652 (N_17652,N_15815,N_16647);
and U17653 (N_17653,N_15672,N_16115);
or U17654 (N_17654,N_16590,N_16333);
and U17655 (N_17655,N_16207,N_15970);
or U17656 (N_17656,N_16439,N_16384);
xnor U17657 (N_17657,N_16155,N_15644);
nand U17658 (N_17658,N_16073,N_16178);
and U17659 (N_17659,N_15984,N_16249);
and U17660 (N_17660,N_16349,N_15636);
xnor U17661 (N_17661,N_16536,N_16549);
xnor U17662 (N_17662,N_16257,N_16522);
nand U17663 (N_17663,N_16607,N_15769);
or U17664 (N_17664,N_16340,N_16560);
xnor U17665 (N_17665,N_16140,N_16177);
nand U17666 (N_17666,N_16245,N_16724);
nor U17667 (N_17667,N_15786,N_16412);
or U17668 (N_17668,N_15709,N_16715);
nor U17669 (N_17669,N_16220,N_16399);
or U17670 (N_17670,N_16348,N_15743);
nor U17671 (N_17671,N_16001,N_16448);
or U17672 (N_17672,N_15767,N_16451);
xor U17673 (N_17673,N_15975,N_16699);
xnor U17674 (N_17674,N_16188,N_16151);
or U17675 (N_17675,N_16035,N_15891);
xor U17676 (N_17676,N_16417,N_16519);
nand U17677 (N_17677,N_16172,N_15658);
nand U17678 (N_17678,N_15906,N_16756);
nor U17679 (N_17679,N_16657,N_16622);
nand U17680 (N_17680,N_16276,N_15704);
nand U17681 (N_17681,N_16436,N_15602);
nand U17682 (N_17682,N_16783,N_16769);
xor U17683 (N_17683,N_15731,N_16569);
nand U17684 (N_17684,N_16610,N_16117);
or U17685 (N_17685,N_16228,N_16393);
nand U17686 (N_17686,N_16362,N_16346);
and U17687 (N_17687,N_16319,N_15750);
nor U17688 (N_17688,N_16275,N_15611);
nor U17689 (N_17689,N_16266,N_16255);
and U17690 (N_17690,N_16321,N_16240);
nand U17691 (N_17691,N_16009,N_15793);
and U17692 (N_17692,N_15678,N_15630);
and U17693 (N_17693,N_15947,N_15630);
xnor U17694 (N_17694,N_15785,N_16098);
and U17695 (N_17695,N_16773,N_16281);
nand U17696 (N_17696,N_16471,N_16076);
xnor U17697 (N_17697,N_15654,N_15694);
nand U17698 (N_17698,N_16463,N_16794);
nand U17699 (N_17699,N_16610,N_16016);
nor U17700 (N_17700,N_16314,N_16093);
nor U17701 (N_17701,N_16344,N_16736);
nand U17702 (N_17702,N_16671,N_16152);
or U17703 (N_17703,N_16734,N_15706);
or U17704 (N_17704,N_16632,N_16040);
nor U17705 (N_17705,N_16716,N_16048);
xnor U17706 (N_17706,N_15976,N_16722);
or U17707 (N_17707,N_16273,N_16738);
xor U17708 (N_17708,N_16660,N_16502);
nor U17709 (N_17709,N_15744,N_15843);
nor U17710 (N_17710,N_15829,N_16457);
xnor U17711 (N_17711,N_16662,N_16249);
and U17712 (N_17712,N_16731,N_16423);
xnor U17713 (N_17713,N_15973,N_15731);
nor U17714 (N_17714,N_16761,N_16032);
nand U17715 (N_17715,N_16402,N_15722);
nand U17716 (N_17716,N_16125,N_15646);
nor U17717 (N_17717,N_16489,N_16626);
nor U17718 (N_17718,N_16039,N_16376);
xor U17719 (N_17719,N_16028,N_16765);
nor U17720 (N_17720,N_16370,N_16040);
xnor U17721 (N_17721,N_15764,N_15703);
or U17722 (N_17722,N_16475,N_15815);
or U17723 (N_17723,N_16100,N_16076);
and U17724 (N_17724,N_16042,N_16645);
xor U17725 (N_17725,N_16248,N_16229);
nand U17726 (N_17726,N_15937,N_16209);
nor U17727 (N_17727,N_15847,N_16342);
nand U17728 (N_17728,N_16727,N_16420);
or U17729 (N_17729,N_16528,N_16771);
and U17730 (N_17730,N_16507,N_15850);
xor U17731 (N_17731,N_16666,N_16024);
nand U17732 (N_17732,N_15612,N_15931);
nor U17733 (N_17733,N_16728,N_16640);
nand U17734 (N_17734,N_16609,N_16750);
or U17735 (N_17735,N_15618,N_15828);
nand U17736 (N_17736,N_16547,N_16005);
nor U17737 (N_17737,N_16327,N_15917);
xor U17738 (N_17738,N_16098,N_16746);
and U17739 (N_17739,N_15729,N_15786);
nand U17740 (N_17740,N_15937,N_16226);
or U17741 (N_17741,N_16171,N_15981);
nor U17742 (N_17742,N_16576,N_16111);
xor U17743 (N_17743,N_15837,N_15712);
nand U17744 (N_17744,N_16079,N_16394);
or U17745 (N_17745,N_16420,N_16196);
xor U17746 (N_17746,N_16791,N_16430);
or U17747 (N_17747,N_16172,N_16123);
nand U17748 (N_17748,N_16505,N_15697);
xnor U17749 (N_17749,N_16747,N_15646);
nor U17750 (N_17750,N_15986,N_16709);
nor U17751 (N_17751,N_16125,N_15998);
nand U17752 (N_17752,N_16727,N_16159);
or U17753 (N_17753,N_15654,N_16519);
or U17754 (N_17754,N_15654,N_16204);
nor U17755 (N_17755,N_16468,N_16134);
nor U17756 (N_17756,N_16589,N_16523);
xor U17757 (N_17757,N_16261,N_16299);
and U17758 (N_17758,N_16184,N_16167);
xor U17759 (N_17759,N_16063,N_16726);
or U17760 (N_17760,N_16514,N_16249);
xor U17761 (N_17761,N_16438,N_16600);
and U17762 (N_17762,N_16367,N_15995);
xnor U17763 (N_17763,N_16065,N_15884);
nor U17764 (N_17764,N_16789,N_16678);
nor U17765 (N_17765,N_15634,N_15969);
and U17766 (N_17766,N_16013,N_16736);
and U17767 (N_17767,N_16308,N_16404);
or U17768 (N_17768,N_16718,N_15944);
nand U17769 (N_17769,N_15910,N_15729);
xor U17770 (N_17770,N_16020,N_15789);
or U17771 (N_17771,N_15849,N_15607);
nand U17772 (N_17772,N_16774,N_15859);
or U17773 (N_17773,N_16125,N_15911);
or U17774 (N_17774,N_15982,N_16381);
and U17775 (N_17775,N_16048,N_16695);
nor U17776 (N_17776,N_15718,N_15869);
nand U17777 (N_17777,N_16474,N_16092);
and U17778 (N_17778,N_15947,N_15994);
xnor U17779 (N_17779,N_15920,N_16219);
nand U17780 (N_17780,N_16242,N_16561);
nor U17781 (N_17781,N_15638,N_15963);
nor U17782 (N_17782,N_15763,N_15795);
nor U17783 (N_17783,N_16312,N_16340);
or U17784 (N_17784,N_16466,N_16095);
nand U17785 (N_17785,N_16356,N_16088);
xor U17786 (N_17786,N_16741,N_16072);
xor U17787 (N_17787,N_15842,N_16600);
nand U17788 (N_17788,N_16674,N_16184);
and U17789 (N_17789,N_16345,N_16718);
nand U17790 (N_17790,N_16282,N_16074);
nand U17791 (N_17791,N_16595,N_15648);
nor U17792 (N_17792,N_16760,N_16714);
nor U17793 (N_17793,N_15703,N_15758);
nor U17794 (N_17794,N_16474,N_15757);
and U17795 (N_17795,N_16072,N_16530);
and U17796 (N_17796,N_16132,N_15828);
and U17797 (N_17797,N_16276,N_15825);
and U17798 (N_17798,N_16631,N_15623);
or U17799 (N_17799,N_16326,N_16672);
xnor U17800 (N_17800,N_16617,N_15868);
and U17801 (N_17801,N_16465,N_16602);
xnor U17802 (N_17802,N_15783,N_16452);
or U17803 (N_17803,N_16716,N_16304);
or U17804 (N_17804,N_16048,N_15911);
xnor U17805 (N_17805,N_15725,N_15781);
xnor U17806 (N_17806,N_16598,N_15822);
nand U17807 (N_17807,N_15731,N_15953);
or U17808 (N_17808,N_15956,N_16290);
xnor U17809 (N_17809,N_15669,N_15965);
and U17810 (N_17810,N_16027,N_15982);
and U17811 (N_17811,N_16420,N_16612);
nor U17812 (N_17812,N_16230,N_16728);
nand U17813 (N_17813,N_15631,N_16197);
xor U17814 (N_17814,N_16234,N_16240);
nand U17815 (N_17815,N_16382,N_15642);
and U17816 (N_17816,N_15613,N_16023);
xor U17817 (N_17817,N_16444,N_15629);
xor U17818 (N_17818,N_16567,N_15730);
nand U17819 (N_17819,N_15960,N_16246);
nor U17820 (N_17820,N_16399,N_16096);
and U17821 (N_17821,N_16498,N_15867);
xor U17822 (N_17822,N_16331,N_16701);
xnor U17823 (N_17823,N_16426,N_16775);
or U17824 (N_17824,N_15767,N_16483);
xor U17825 (N_17825,N_15618,N_15937);
xor U17826 (N_17826,N_16522,N_15867);
or U17827 (N_17827,N_16532,N_16712);
and U17828 (N_17828,N_16148,N_16295);
xor U17829 (N_17829,N_15997,N_15847);
nand U17830 (N_17830,N_16666,N_16746);
nand U17831 (N_17831,N_15832,N_16256);
and U17832 (N_17832,N_16469,N_15759);
xor U17833 (N_17833,N_16142,N_15760);
nor U17834 (N_17834,N_16448,N_16229);
nor U17835 (N_17835,N_16246,N_16636);
nand U17836 (N_17836,N_15627,N_16540);
or U17837 (N_17837,N_16618,N_15945);
nor U17838 (N_17838,N_16232,N_16010);
xnor U17839 (N_17839,N_16145,N_16012);
or U17840 (N_17840,N_15940,N_15865);
xnor U17841 (N_17841,N_16326,N_15823);
and U17842 (N_17842,N_15750,N_15928);
xnor U17843 (N_17843,N_15838,N_16024);
nor U17844 (N_17844,N_16627,N_16738);
xnor U17845 (N_17845,N_16049,N_16090);
or U17846 (N_17846,N_16745,N_16229);
nor U17847 (N_17847,N_16525,N_16661);
nor U17848 (N_17848,N_16258,N_16650);
and U17849 (N_17849,N_16610,N_16052);
or U17850 (N_17850,N_16451,N_16660);
nand U17851 (N_17851,N_15695,N_16385);
nand U17852 (N_17852,N_16306,N_15918);
nand U17853 (N_17853,N_16045,N_15683);
or U17854 (N_17854,N_16140,N_16217);
or U17855 (N_17855,N_16773,N_16444);
and U17856 (N_17856,N_15825,N_16565);
and U17857 (N_17857,N_16106,N_16666);
xnor U17858 (N_17858,N_16600,N_15626);
nand U17859 (N_17859,N_16287,N_16199);
or U17860 (N_17860,N_16394,N_16189);
xor U17861 (N_17861,N_16592,N_15673);
or U17862 (N_17862,N_16199,N_15853);
xnor U17863 (N_17863,N_16035,N_15871);
or U17864 (N_17864,N_15805,N_16169);
nand U17865 (N_17865,N_16361,N_15992);
nand U17866 (N_17866,N_16246,N_16028);
nand U17867 (N_17867,N_16636,N_16447);
and U17868 (N_17868,N_16431,N_15706);
or U17869 (N_17869,N_16460,N_15863);
nand U17870 (N_17870,N_16189,N_15908);
nand U17871 (N_17871,N_16511,N_15669);
or U17872 (N_17872,N_15997,N_16144);
and U17873 (N_17873,N_15965,N_16291);
or U17874 (N_17874,N_16209,N_16134);
nor U17875 (N_17875,N_16393,N_15905);
and U17876 (N_17876,N_16126,N_16498);
nand U17877 (N_17877,N_16729,N_15724);
nand U17878 (N_17878,N_15885,N_16421);
xor U17879 (N_17879,N_16406,N_16506);
xnor U17880 (N_17880,N_16621,N_16523);
or U17881 (N_17881,N_15746,N_15867);
and U17882 (N_17882,N_16252,N_16610);
nand U17883 (N_17883,N_16439,N_16283);
and U17884 (N_17884,N_15981,N_16495);
or U17885 (N_17885,N_16750,N_16032);
and U17886 (N_17886,N_15886,N_16650);
nand U17887 (N_17887,N_15669,N_16377);
and U17888 (N_17888,N_15619,N_15867);
xnor U17889 (N_17889,N_15665,N_15655);
nand U17890 (N_17890,N_16150,N_16746);
and U17891 (N_17891,N_16132,N_16194);
xor U17892 (N_17892,N_15874,N_16087);
nor U17893 (N_17893,N_15808,N_15986);
xnor U17894 (N_17894,N_15833,N_15716);
xor U17895 (N_17895,N_16078,N_16055);
or U17896 (N_17896,N_16099,N_15622);
nor U17897 (N_17897,N_16098,N_16449);
nor U17898 (N_17898,N_15956,N_16375);
nor U17899 (N_17899,N_15935,N_16616);
nor U17900 (N_17900,N_16637,N_16364);
xor U17901 (N_17901,N_16445,N_16332);
nor U17902 (N_17902,N_15779,N_15649);
nand U17903 (N_17903,N_16423,N_16553);
nor U17904 (N_17904,N_16758,N_15882);
xnor U17905 (N_17905,N_15930,N_16543);
or U17906 (N_17906,N_16406,N_16277);
nand U17907 (N_17907,N_16293,N_15822);
nand U17908 (N_17908,N_16108,N_16147);
and U17909 (N_17909,N_16790,N_15901);
nand U17910 (N_17910,N_15813,N_16412);
or U17911 (N_17911,N_16024,N_16328);
nand U17912 (N_17912,N_16355,N_16097);
nor U17913 (N_17913,N_16505,N_16007);
and U17914 (N_17914,N_16706,N_16142);
nand U17915 (N_17915,N_16359,N_15607);
nor U17916 (N_17916,N_15654,N_15740);
nand U17917 (N_17917,N_16044,N_16296);
xnor U17918 (N_17918,N_16469,N_15931);
or U17919 (N_17919,N_16195,N_16388);
nor U17920 (N_17920,N_16630,N_15699);
or U17921 (N_17921,N_16192,N_15941);
nand U17922 (N_17922,N_16243,N_15716);
xor U17923 (N_17923,N_16675,N_15786);
nand U17924 (N_17924,N_15853,N_16763);
nor U17925 (N_17925,N_16507,N_15950);
xnor U17926 (N_17926,N_16525,N_16166);
nand U17927 (N_17927,N_16756,N_15674);
and U17928 (N_17928,N_16255,N_16288);
or U17929 (N_17929,N_16702,N_15777);
nor U17930 (N_17930,N_15880,N_15799);
nand U17931 (N_17931,N_16038,N_16788);
nand U17932 (N_17932,N_16774,N_16196);
or U17933 (N_17933,N_16262,N_16695);
xor U17934 (N_17934,N_16716,N_16631);
and U17935 (N_17935,N_15752,N_16421);
xor U17936 (N_17936,N_16273,N_15855);
xor U17937 (N_17937,N_16526,N_16128);
xor U17938 (N_17938,N_16633,N_15702);
and U17939 (N_17939,N_16094,N_16589);
nor U17940 (N_17940,N_16016,N_16703);
xnor U17941 (N_17941,N_16360,N_15860);
and U17942 (N_17942,N_16214,N_16541);
or U17943 (N_17943,N_15882,N_16429);
nor U17944 (N_17944,N_15667,N_16185);
and U17945 (N_17945,N_16076,N_15945);
nor U17946 (N_17946,N_16381,N_16185);
xnor U17947 (N_17947,N_16702,N_15787);
nand U17948 (N_17948,N_16138,N_16077);
xor U17949 (N_17949,N_15602,N_16663);
nor U17950 (N_17950,N_16790,N_16540);
or U17951 (N_17951,N_15879,N_15603);
nand U17952 (N_17952,N_15705,N_15752);
xor U17953 (N_17953,N_15798,N_15821);
or U17954 (N_17954,N_16715,N_16393);
and U17955 (N_17955,N_16076,N_16229);
xnor U17956 (N_17956,N_16431,N_16393);
xor U17957 (N_17957,N_15975,N_15718);
xor U17958 (N_17958,N_16577,N_16614);
xor U17959 (N_17959,N_16034,N_16052);
nor U17960 (N_17960,N_15964,N_16666);
nand U17961 (N_17961,N_15746,N_16301);
nor U17962 (N_17962,N_16501,N_15867);
or U17963 (N_17963,N_16132,N_15650);
nand U17964 (N_17964,N_16302,N_16289);
or U17965 (N_17965,N_15603,N_16155);
and U17966 (N_17966,N_16609,N_15928);
or U17967 (N_17967,N_16305,N_16625);
nor U17968 (N_17968,N_16022,N_16394);
nor U17969 (N_17969,N_16634,N_16347);
nor U17970 (N_17970,N_16534,N_15924);
and U17971 (N_17971,N_15719,N_16716);
nand U17972 (N_17972,N_16356,N_16216);
nand U17973 (N_17973,N_15828,N_16623);
nor U17974 (N_17974,N_16159,N_15690);
and U17975 (N_17975,N_16414,N_16579);
or U17976 (N_17976,N_16367,N_16322);
nor U17977 (N_17977,N_16486,N_15604);
and U17978 (N_17978,N_15872,N_15960);
nor U17979 (N_17979,N_16236,N_16510);
nand U17980 (N_17980,N_16463,N_15617);
nor U17981 (N_17981,N_16011,N_16435);
xnor U17982 (N_17982,N_16638,N_15908);
and U17983 (N_17983,N_16382,N_15672);
xor U17984 (N_17984,N_16531,N_15996);
nand U17985 (N_17985,N_16718,N_16515);
and U17986 (N_17986,N_15834,N_15747);
xnor U17987 (N_17987,N_16705,N_16716);
or U17988 (N_17988,N_15613,N_15692);
nor U17989 (N_17989,N_16718,N_16009);
and U17990 (N_17990,N_15854,N_16497);
nand U17991 (N_17991,N_16234,N_16215);
xnor U17992 (N_17992,N_16609,N_16743);
xnor U17993 (N_17993,N_15843,N_16113);
and U17994 (N_17994,N_16185,N_16215);
and U17995 (N_17995,N_16031,N_15972);
nor U17996 (N_17996,N_16268,N_16673);
and U17997 (N_17997,N_15699,N_16459);
nand U17998 (N_17998,N_16424,N_16566);
nor U17999 (N_17999,N_15826,N_16112);
nand U18000 (N_18000,N_17275,N_17369);
xor U18001 (N_18001,N_17302,N_17488);
and U18002 (N_18002,N_17392,N_16803);
xnor U18003 (N_18003,N_17842,N_17944);
nor U18004 (N_18004,N_17777,N_17370);
nor U18005 (N_18005,N_17863,N_17271);
and U18006 (N_18006,N_16857,N_17883);
and U18007 (N_18007,N_17474,N_17606);
and U18008 (N_18008,N_17290,N_17774);
nor U18009 (N_18009,N_16839,N_17267);
nand U18010 (N_18010,N_17330,N_17658);
nor U18011 (N_18011,N_16896,N_17976);
xor U18012 (N_18012,N_17362,N_17455);
or U18013 (N_18013,N_17490,N_17578);
nand U18014 (N_18014,N_17967,N_17304);
nand U18015 (N_18015,N_16954,N_17841);
or U18016 (N_18016,N_17990,N_17270);
xor U18017 (N_18017,N_17377,N_16948);
xor U18018 (N_18018,N_17085,N_17049);
nand U18019 (N_18019,N_17603,N_17688);
and U18020 (N_18020,N_17792,N_17033);
xnor U18021 (N_18021,N_17629,N_17553);
and U18022 (N_18022,N_17957,N_17793);
or U18023 (N_18023,N_17812,N_17943);
nand U18024 (N_18024,N_17926,N_17038);
nor U18025 (N_18025,N_17543,N_17668);
or U18026 (N_18026,N_17700,N_17634);
nor U18027 (N_18027,N_17588,N_17234);
nor U18028 (N_18028,N_17709,N_16846);
nand U18029 (N_18029,N_17401,N_17790);
and U18030 (N_18030,N_17140,N_17419);
xor U18031 (N_18031,N_17139,N_17040);
nor U18032 (N_18032,N_17272,N_16810);
nand U18033 (N_18033,N_16864,N_17174);
xor U18034 (N_18034,N_17004,N_17440);
or U18035 (N_18035,N_16827,N_17879);
and U18036 (N_18036,N_17529,N_17882);
nand U18037 (N_18037,N_17281,N_16808);
xor U18038 (N_18038,N_17924,N_16943);
and U18039 (N_18039,N_16820,N_17978);
and U18040 (N_18040,N_17589,N_17824);
or U18041 (N_18041,N_17326,N_17745);
or U18042 (N_18042,N_16910,N_17482);
or U18043 (N_18043,N_17852,N_17207);
nor U18044 (N_18044,N_16824,N_17911);
xor U18045 (N_18045,N_17050,N_17441);
or U18046 (N_18046,N_17933,N_17783);
nand U18047 (N_18047,N_17143,N_16877);
or U18048 (N_18048,N_16835,N_16904);
and U18049 (N_18049,N_17509,N_17526);
and U18050 (N_18050,N_17374,N_17857);
and U18051 (N_18051,N_17518,N_16855);
and U18052 (N_18052,N_17115,N_17664);
or U18053 (N_18053,N_17400,N_17355);
nand U18054 (N_18054,N_17618,N_17456);
xor U18055 (N_18055,N_17715,N_17604);
or U18056 (N_18056,N_16981,N_17550);
nor U18057 (N_18057,N_17395,N_17895);
xor U18058 (N_18058,N_17546,N_16922);
nand U18059 (N_18059,N_17887,N_17200);
nand U18060 (N_18060,N_16883,N_17402);
or U18061 (N_18061,N_17835,N_17427);
and U18062 (N_18062,N_17849,N_17558);
nor U18063 (N_18063,N_17959,N_17838);
or U18064 (N_18064,N_17818,N_17333);
or U18065 (N_18065,N_17549,N_16964);
nor U18066 (N_18066,N_17391,N_16923);
nor U18067 (N_18067,N_17813,N_17897);
nand U18068 (N_18068,N_17307,N_17547);
and U18069 (N_18069,N_17937,N_16843);
nand U18070 (N_18070,N_17432,N_17577);
or U18071 (N_18071,N_17502,N_17952);
or U18072 (N_18072,N_17878,N_17182);
or U18073 (N_18073,N_16939,N_17136);
nand U18074 (N_18074,N_17834,N_17090);
nand U18075 (N_18075,N_17251,N_16925);
xor U18076 (N_18076,N_17292,N_17196);
nor U18077 (N_18077,N_17872,N_16870);
nand U18078 (N_18078,N_17601,N_17697);
nand U18079 (N_18079,N_17789,N_17364);
and U18080 (N_18080,N_17497,N_17718);
xor U18081 (N_18081,N_17582,N_17757);
xnor U18082 (N_18082,N_17424,N_16933);
and U18083 (N_18083,N_17283,N_17379);
and U18084 (N_18084,N_17367,N_17285);
and U18085 (N_18085,N_17390,N_16814);
nand U18086 (N_18086,N_17172,N_16862);
or U18087 (N_18087,N_17405,N_16965);
nand U18088 (N_18088,N_17189,N_17311);
nor U18089 (N_18089,N_17342,N_16851);
nand U18090 (N_18090,N_17693,N_17956);
and U18091 (N_18091,N_17542,N_17756);
or U18092 (N_18092,N_17845,N_17650);
nor U18093 (N_18093,N_17078,N_17059);
nor U18094 (N_18094,N_17436,N_17516);
nor U18095 (N_18095,N_17562,N_16995);
xor U18096 (N_18096,N_17185,N_17113);
nand U18097 (N_18097,N_17035,N_16853);
and U18098 (N_18098,N_16957,N_17861);
nor U18099 (N_18099,N_16816,N_17315);
or U18100 (N_18100,N_16913,N_17570);
xnor U18101 (N_18101,N_17205,N_16966);
and U18102 (N_18102,N_16998,N_17511);
nor U18103 (N_18103,N_17028,N_17983);
nand U18104 (N_18104,N_17908,N_17929);
or U18105 (N_18105,N_16813,N_17094);
xnor U18106 (N_18106,N_17221,N_16873);
or U18107 (N_18107,N_16976,N_17261);
nor U18108 (N_18108,N_16856,N_17313);
or U18109 (N_18109,N_17387,N_17008);
and U18110 (N_18110,N_17985,N_17396);
nand U18111 (N_18111,N_17788,N_17416);
nand U18112 (N_18112,N_17052,N_17321);
and U18113 (N_18113,N_16825,N_17936);
xor U18114 (N_18114,N_16961,N_17866);
or U18115 (N_18115,N_17042,N_17707);
and U18116 (N_18116,N_17653,N_17660);
xor U18117 (N_18117,N_17760,N_16932);
and U18118 (N_18118,N_17994,N_17471);
nor U18119 (N_18119,N_17692,N_17969);
or U18120 (N_18120,N_17800,N_17736);
or U18121 (N_18121,N_17150,N_17466);
or U18122 (N_18122,N_17593,N_16879);
and U18123 (N_18123,N_17260,N_17157);
and U18124 (N_18124,N_17087,N_17361);
xor U18125 (N_18125,N_17286,N_17968);
nor U18126 (N_18126,N_17032,N_17227);
and U18127 (N_18127,N_17235,N_17651);
xnor U18128 (N_18128,N_17346,N_17590);
xnor U18129 (N_18129,N_17024,N_17327);
xnor U18130 (N_18130,N_17403,N_17850);
nor U18131 (N_18131,N_17460,N_17195);
xor U18132 (N_18132,N_17726,N_17947);
nor U18133 (N_18133,N_16978,N_17619);
nand U18134 (N_18134,N_16905,N_17735);
nand U18135 (N_18135,N_17414,N_16973);
and U18136 (N_18136,N_17884,N_17310);
xor U18137 (N_18137,N_17397,N_17750);
and U18138 (N_18138,N_16980,N_17954);
nand U18139 (N_18139,N_16907,N_17521);
nor U18140 (N_18140,N_17918,N_17254);
and U18141 (N_18141,N_17125,N_17960);
or U18142 (N_18142,N_17406,N_17851);
or U18143 (N_18143,N_17002,N_17472);
nand U18144 (N_18144,N_17439,N_17503);
nand U18145 (N_18145,N_17612,N_17997);
or U18146 (N_18146,N_17206,N_16982);
xnor U18147 (N_18147,N_16867,N_17477);
or U18148 (N_18148,N_17998,N_17739);
xnor U18149 (N_18149,N_17385,N_17015);
xor U18150 (N_18150,N_16991,N_17043);
nor U18151 (N_18151,N_17611,N_17581);
nand U18152 (N_18152,N_17595,N_16833);
nand U18153 (N_18153,N_17422,N_17572);
and U18154 (N_18154,N_16929,N_17678);
and U18155 (N_18155,N_17265,N_17671);
xor U18156 (N_18156,N_17625,N_17345);
and U18157 (N_18157,N_17248,N_17623);
nand U18158 (N_18158,N_17124,N_17661);
nor U18159 (N_18159,N_17076,N_17948);
or U18160 (N_18160,N_17666,N_16916);
or U18161 (N_18161,N_16861,N_17989);
nor U18162 (N_18162,N_16812,N_16847);
nand U18163 (N_18163,N_16866,N_17946);
nor U18164 (N_18164,N_17393,N_17188);
or U18165 (N_18165,N_17628,N_17949);
or U18166 (N_18166,N_17173,N_17092);
and U18167 (N_18167,N_17016,N_17175);
xnor U18168 (N_18168,N_17772,N_17130);
and U18169 (N_18169,N_17714,N_16920);
and U18170 (N_18170,N_17022,N_17411);
and U18171 (N_18171,N_17066,N_16901);
nor U18172 (N_18172,N_16848,N_16823);
xor U18173 (N_18173,N_17586,N_17154);
xnor U18174 (N_18174,N_17031,N_17348);
or U18175 (N_18175,N_17239,N_17498);
nand U18176 (N_18176,N_17571,N_17901);
nor U18177 (N_18177,N_17831,N_17381);
nand U18178 (N_18178,N_17519,N_17843);
nand U18179 (N_18179,N_17241,N_17097);
or U18180 (N_18180,N_17940,N_17149);
nand U18181 (N_18181,N_17111,N_16804);
xor U18182 (N_18182,N_17413,N_17366);
nor U18183 (N_18183,N_16850,N_17686);
xnor U18184 (N_18184,N_17054,N_17334);
or U18185 (N_18185,N_17105,N_17828);
nor U18186 (N_18186,N_17810,N_17089);
xnor U18187 (N_18187,N_17259,N_17303);
nand U18188 (N_18188,N_17447,N_16934);
nand U18189 (N_18189,N_17806,N_17670);
and U18190 (N_18190,N_17430,N_17375);
nand U18191 (N_18191,N_17371,N_17823);
or U18192 (N_18192,N_17600,N_17677);
nor U18193 (N_18193,N_17088,N_17388);
nand U18194 (N_18194,N_17359,N_16881);
xor U18195 (N_18195,N_17891,N_17148);
xnor U18196 (N_18196,N_17126,N_17568);
nand U18197 (N_18197,N_17018,N_17719);
xor U18198 (N_18198,N_17465,N_17565);
nor U18199 (N_18199,N_17525,N_17902);
and U18200 (N_18200,N_17928,N_17190);
and U18201 (N_18201,N_17225,N_17048);
or U18202 (N_18202,N_17457,N_17063);
and U18203 (N_18203,N_17343,N_17825);
and U18204 (N_18204,N_17885,N_16930);
nor U18205 (N_18205,N_17617,N_17860);
nor U18206 (N_18206,N_17844,N_17382);
and U18207 (N_18207,N_16888,N_17627);
nor U18208 (N_18208,N_17080,N_17914);
or U18209 (N_18209,N_17418,N_17036);
nor U18210 (N_18210,N_17277,N_17811);
and U18211 (N_18211,N_17613,N_17494);
and U18212 (N_18212,N_17404,N_17909);
nand U18213 (N_18213,N_17915,N_17514);
nor U18214 (N_18214,N_17047,N_16945);
nor U18215 (N_18215,N_17481,N_17373);
and U18216 (N_18216,N_17833,N_16990);
or U18217 (N_18217,N_17025,N_17041);
or U18218 (N_18218,N_17759,N_17657);
and U18219 (N_18219,N_16918,N_17244);
or U18220 (N_18220,N_16805,N_17412);
and U18221 (N_18221,N_17308,N_17231);
nor U18222 (N_18222,N_16868,N_17006);
xnor U18223 (N_18223,N_17134,N_17615);
nand U18224 (N_18224,N_17433,N_16865);
and U18225 (N_18225,N_17836,N_17508);
nor U18226 (N_18226,N_17058,N_17177);
and U18227 (N_18227,N_17165,N_17945);
nor U18228 (N_18228,N_16906,N_17742);
nor U18229 (N_18229,N_17840,N_16936);
nor U18230 (N_18230,N_16869,N_17871);
nor U18231 (N_18231,N_17691,N_17469);
xnor U18232 (N_18232,N_16967,N_17218);
xor U18233 (N_18233,N_17996,N_16985);
nand U18234 (N_18234,N_16992,N_17821);
nand U18235 (N_18235,N_17110,N_17109);
nor U18236 (N_18236,N_17484,N_17734);
xnor U18237 (N_18237,N_17987,N_16819);
and U18238 (N_18238,N_17725,N_17880);
and U18239 (N_18239,N_17713,N_16997);
xor U18240 (N_18240,N_17923,N_17091);
nor U18241 (N_18241,N_16950,N_17731);
and U18242 (N_18242,N_17753,N_17183);
nand U18243 (N_18243,N_17238,N_17003);
and U18244 (N_18244,N_17922,N_17132);
or U18245 (N_18245,N_16832,N_17564);
and U18246 (N_18246,N_17903,N_17010);
and U18247 (N_18247,N_17011,N_17328);
or U18248 (N_18248,N_17428,N_17684);
nor U18249 (N_18249,N_17696,N_17293);
and U18250 (N_18250,N_17941,N_16893);
and U18251 (N_18251,N_17316,N_17780);
and U18252 (N_18252,N_17191,N_17512);
and U18253 (N_18253,N_17250,N_17782);
or U18254 (N_18254,N_17768,N_17758);
and U18255 (N_18255,N_17893,N_17829);
xnor U18256 (N_18256,N_16884,N_17791);
or U18257 (N_18257,N_16993,N_17730);
nand U18258 (N_18258,N_17483,N_16829);
nand U18259 (N_18259,N_17787,N_16876);
and U18260 (N_18260,N_17991,N_17106);
nor U18261 (N_18261,N_17309,N_17596);
nor U18262 (N_18262,N_17803,N_17973);
nor U18263 (N_18263,N_17434,N_17938);
nand U18264 (N_18264,N_16807,N_16899);
and U18265 (N_18265,N_17253,N_17255);
nand U18266 (N_18266,N_17476,N_17746);
or U18267 (N_18267,N_17338,N_17233);
nor U18268 (N_18268,N_16871,N_17705);
or U18269 (N_18269,N_17877,N_17552);
or U18270 (N_18270,N_17485,N_17269);
xor U18271 (N_18271,N_17649,N_17257);
or U18272 (N_18272,N_17710,N_16898);
or U18273 (N_18273,N_17630,N_17357);
and U18274 (N_18274,N_17569,N_17112);
and U18275 (N_18275,N_17458,N_16872);
nor U18276 (N_18276,N_16858,N_17979);
and U18277 (N_18277,N_17153,N_17012);
nand U18278 (N_18278,N_16818,N_16892);
and U18279 (N_18279,N_17534,N_16996);
xor U18280 (N_18280,N_17305,N_17673);
nor U18281 (N_18281,N_17646,N_17167);
nor U18282 (N_18282,N_17480,N_16989);
and U18283 (N_18283,N_16956,N_17256);
and U18284 (N_18284,N_17662,N_17817);
and U18285 (N_18285,N_17240,N_17168);
or U18286 (N_18286,N_17900,N_17000);
nand U18287 (N_18287,N_17608,N_17682);
nand U18288 (N_18288,N_17284,N_16844);
nor U18289 (N_18289,N_17197,N_17925);
nor U18290 (N_18290,N_17906,N_17119);
and U18291 (N_18291,N_17082,N_17815);
or U18292 (N_18292,N_17489,N_17280);
xnor U18293 (N_18293,N_16972,N_17068);
xnor U18294 (N_18294,N_17556,N_17762);
or U18295 (N_18295,N_17560,N_16987);
nor U18296 (N_18296,N_17717,N_17522);
or U18297 (N_18297,N_17607,N_17169);
xor U18298 (N_18298,N_17778,N_17687);
or U18299 (N_18299,N_17192,N_17096);
or U18300 (N_18300,N_17832,N_17905);
nor U18301 (N_18301,N_17958,N_16822);
nor U18302 (N_18302,N_17770,N_16900);
and U18303 (N_18303,N_17263,N_17030);
or U18304 (N_18304,N_17856,N_17537);
or U18305 (N_18305,N_17984,N_17072);
or U18306 (N_18306,N_17754,N_17219);
or U18307 (N_18307,N_16886,N_17398);
xnor U18308 (N_18308,N_17084,N_17423);
nand U18309 (N_18309,N_17045,N_16838);
or U18310 (N_18310,N_17242,N_17977);
nor U18311 (N_18311,N_17889,N_17868);
nor U18312 (N_18312,N_16951,N_17222);
and U18313 (N_18313,N_17539,N_17317);
and U18314 (N_18314,N_17298,N_16979);
or U18315 (N_18315,N_16841,N_17862);
nor U18316 (N_18316,N_17795,N_16902);
xor U18317 (N_18317,N_17459,N_17276);
nand U18318 (N_18318,N_17609,N_17029);
and U18319 (N_18319,N_17892,N_17340);
nand U18320 (N_18320,N_17118,N_17224);
xor U18321 (N_18321,N_17711,N_17230);
nor U18322 (N_18322,N_17950,N_17626);
nor U18323 (N_18323,N_17386,N_17282);
or U18324 (N_18324,N_17288,N_17749);
nand U18325 (N_18325,N_17733,N_17212);
and U18326 (N_18326,N_17216,N_17732);
or U18327 (N_18327,N_17493,N_17258);
or U18328 (N_18328,N_17801,N_17656);
nand U18329 (N_18329,N_17814,N_17669);
xor U18330 (N_18330,N_17741,N_17487);
xnor U18331 (N_18331,N_17721,N_17594);
xor U18332 (N_18332,N_17435,N_17995);
nor U18333 (N_18333,N_16890,N_17499);
and U18334 (N_18334,N_17468,N_17808);
xor U18335 (N_18335,N_17859,N_17232);
and U18336 (N_18336,N_17591,N_17703);
nor U18337 (N_18337,N_17538,N_17579);
nand U18338 (N_18338,N_17689,N_17152);
nor U18339 (N_18339,N_17443,N_16924);
nand U18340 (N_18340,N_17492,N_17322);
nand U18341 (N_18341,N_17694,N_17384);
or U18342 (N_18342,N_16975,N_17127);
xor U18343 (N_18343,N_16885,N_17086);
nor U18344 (N_18344,N_17580,N_17797);
nand U18345 (N_18345,N_16959,N_17463);
and U18346 (N_18346,N_16960,N_17504);
xor U18347 (N_18347,N_17005,N_16821);
or U18348 (N_18348,N_17784,N_16830);
nor U18349 (N_18349,N_17663,N_16931);
nand U18350 (N_18350,N_17461,N_16811);
nand U18351 (N_18351,N_17799,N_17951);
and U18352 (N_18352,N_17273,N_17654);
xnor U18353 (N_18353,N_17473,N_17816);
nand U18354 (N_18354,N_17548,N_17324);
nand U18355 (N_18355,N_17744,N_17765);
nor U18356 (N_18356,N_17245,N_16955);
xor U18357 (N_18357,N_17417,N_17934);
nor U18358 (N_18358,N_17104,N_17056);
or U18359 (N_18359,N_17160,N_17920);
and U18360 (N_18360,N_17645,N_17121);
nor U18361 (N_18361,N_16926,N_17116);
nand U18362 (N_18362,N_17702,N_16895);
nor U18363 (N_18363,N_17873,N_17513);
nor U18364 (N_18364,N_17993,N_17467);
nor U18365 (N_18365,N_17826,N_17120);
nor U18366 (N_18366,N_17786,N_17114);
nand U18367 (N_18367,N_17510,N_17462);
nor U18368 (N_18368,N_17927,N_17237);
and U18369 (N_18369,N_17583,N_16977);
and U18370 (N_18370,N_17738,N_17243);
xor U18371 (N_18371,N_17720,N_17201);
xnor U18372 (N_18372,N_16999,N_17751);
nor U18373 (N_18373,N_17202,N_17210);
nand U18374 (N_18374,N_17597,N_17318);
and U18375 (N_18375,N_17681,N_17454);
and U18376 (N_18376,N_17869,N_17249);
nand U18377 (N_18377,N_17349,N_17354);
or U18378 (N_18378,N_17426,N_17953);
nand U18379 (N_18379,N_17798,N_17372);
nand U18380 (N_18380,N_17368,N_17541);
xor U18381 (N_18381,N_17637,N_16944);
xor U18382 (N_18382,N_17610,N_17728);
or U18383 (N_18383,N_17021,N_17648);
xor U18384 (N_18384,N_16970,N_17389);
xor U18385 (N_18385,N_17164,N_17181);
xnor U18386 (N_18386,N_17079,N_17351);
nor U18387 (N_18387,N_17986,N_17955);
and U18388 (N_18388,N_16894,N_16878);
xnor U18389 (N_18389,N_16940,N_17363);
nand U18390 (N_18390,N_17699,N_17545);
or U18391 (N_18391,N_17229,N_16953);
nand U18392 (N_18392,N_17331,N_17246);
or U18393 (N_18393,N_17123,N_17640);
nand U18394 (N_18394,N_17639,N_17523);
nor U18395 (N_18395,N_17988,N_17505);
nand U18396 (N_18396,N_17128,N_17533);
nand U18397 (N_18397,N_16958,N_17704);
or U18398 (N_18398,N_17659,N_17159);
nand U18399 (N_18399,N_17767,N_16802);
or U18400 (N_18400,N_17444,N_17574);
or U18401 (N_18401,N_17655,N_17314);
nor U18402 (N_18402,N_17252,N_16891);
xnor U18403 (N_18403,N_17614,N_17198);
nor U18404 (N_18404,N_17535,N_17449);
xor U18405 (N_18405,N_17599,N_17641);
nand U18406 (N_18406,N_17319,N_17060);
xor U18407 (N_18407,N_17561,N_17775);
xnor U18408 (N_18408,N_16882,N_17962);
nand U18409 (N_18409,N_17100,N_17199);
or U18410 (N_18410,N_17446,N_17620);
and U18411 (N_18411,N_17358,N_17500);
xor U18412 (N_18412,N_17966,N_17971);
and U18413 (N_18413,N_17633,N_17685);
xnor U18414 (N_18414,N_17420,N_17724);
or U18415 (N_18415,N_17062,N_17378);
xnor U18416 (N_18416,N_16962,N_17794);
and U18417 (N_18417,N_17407,N_17053);
xor U18418 (N_18418,N_17070,N_17223);
xor U18419 (N_18419,N_17051,N_17044);
nor U18420 (N_18420,N_17020,N_17009);
or U18421 (N_18421,N_17320,N_17819);
nand U18422 (N_18422,N_17870,N_17890);
xor U18423 (N_18423,N_17083,N_17667);
or U18424 (N_18424,N_16903,N_17980);
nor U18425 (N_18425,N_17046,N_16911);
or U18426 (N_18426,N_17769,N_16927);
xor U18427 (N_18427,N_17323,N_17847);
or U18428 (N_18428,N_17266,N_16801);
and U18429 (N_18429,N_17982,N_17796);
xnor U18430 (N_18430,N_17007,N_17208);
xnor U18431 (N_18431,N_17913,N_17972);
nand U18432 (N_18432,N_17352,N_17716);
xor U18433 (N_18433,N_17540,N_17974);
xnor U18434 (N_18434,N_17142,N_17631);
xnor U18435 (N_18435,N_17486,N_16837);
or U18436 (N_18436,N_17771,N_16889);
xnor U18437 (N_18437,N_17300,N_17409);
nand U18438 (N_18438,N_17643,N_16852);
or U18439 (N_18439,N_17448,N_16834);
nor U18440 (N_18440,N_17665,N_17383);
nor U18441 (N_18441,N_17554,N_16942);
or U18442 (N_18442,N_17647,N_17853);
nor U18443 (N_18443,N_17912,N_17932);
nor U18444 (N_18444,N_17065,N_17672);
nor U18445 (N_18445,N_17764,N_17155);
nand U18446 (N_18446,N_17743,N_16988);
xnor U18447 (N_18447,N_17299,N_17635);
nor U18448 (N_18448,N_17855,N_16986);
or U18449 (N_18449,N_16968,N_17585);
xor U18450 (N_18450,N_17779,N_17876);
nand U18451 (N_18451,N_16831,N_17421);
nor U18452 (N_18452,N_17176,N_17761);
nand U18453 (N_18453,N_16809,N_17805);
nand U18454 (N_18454,N_17329,N_16840);
or U18455 (N_18455,N_17394,N_16875);
nor U18456 (N_18456,N_17729,N_17067);
nand U18457 (N_18457,N_17108,N_17527);
xor U18458 (N_18458,N_16983,N_16915);
xor U18459 (N_18459,N_17566,N_17353);
xor U18460 (N_18460,N_17312,N_17587);
xor U18461 (N_18461,N_17921,N_17170);
xor U18462 (N_18462,N_17917,N_17098);
or U18463 (N_18463,N_16880,N_17264);
nor U18464 (N_18464,N_17544,N_17970);
and U18465 (N_18465,N_17675,N_17632);
nand U18466 (N_18466,N_16860,N_17506);
and U18467 (N_18467,N_17350,N_16887);
nand U18468 (N_18468,N_17723,N_16917);
nor U18469 (N_18469,N_17575,N_17592);
nand U18470 (N_18470,N_17129,N_17356);
nor U18471 (N_18471,N_17652,N_17013);
and U18472 (N_18472,N_17144,N_16854);
nand U18473 (N_18473,N_17874,N_16842);
or U18474 (N_18474,N_17999,N_17425);
or U18475 (N_18475,N_17992,N_17807);
and U18476 (N_18476,N_16946,N_17748);
xnor U18477 (N_18477,N_16859,N_17228);
and U18478 (N_18478,N_17848,N_17194);
nand U18479 (N_18479,N_17881,N_17624);
nand U18480 (N_18480,N_17039,N_17274);
nor U18481 (N_18481,N_17528,N_17184);
nor U18482 (N_18482,N_17122,N_16941);
xnor U18483 (N_18483,N_17894,N_16908);
and U18484 (N_18484,N_17961,N_17809);
or U18485 (N_18485,N_17339,N_17706);
nor U18486 (N_18486,N_16984,N_17820);
or U18487 (N_18487,N_17023,N_17584);
nand U18488 (N_18488,N_17151,N_17147);
nor U18489 (N_18489,N_17138,N_17642);
and U18490 (N_18490,N_17804,N_17209);
and U18491 (N_18491,N_17896,N_17268);
nor U18492 (N_18492,N_17220,N_16849);
xnor U18493 (N_18493,N_16909,N_17297);
and U18494 (N_18494,N_17034,N_17964);
xor U18495 (N_18495,N_17559,N_17598);
or U18496 (N_18496,N_17335,N_17163);
nor U18497 (N_18497,N_17524,N_17690);
nor U18498 (N_18498,N_17306,N_17103);
nor U18499 (N_18499,N_17701,N_17875);
and U18500 (N_18500,N_17864,N_17213);
and U18501 (N_18501,N_16845,N_17296);
xor U18502 (N_18502,N_17898,N_17226);
xor U18503 (N_18503,N_16863,N_17453);
nand U18504 (N_18504,N_16971,N_17429);
nand U18505 (N_18505,N_17464,N_16952);
xnor U18506 (N_18506,N_17919,N_17291);
and U18507 (N_18507,N_17939,N_17001);
xnor U18508 (N_18508,N_17061,N_17203);
nor U18509 (N_18509,N_17247,N_16938);
or U18510 (N_18510,N_17837,N_17442);
nor U18511 (N_18511,N_17916,N_17491);
or U18512 (N_18512,N_17014,N_17077);
or U18513 (N_18513,N_17766,N_17278);
or U18514 (N_18514,N_16815,N_16874);
and U18515 (N_18515,N_17496,N_16826);
xnor U18516 (N_18516,N_17095,N_17846);
and U18517 (N_18517,N_17517,N_17075);
or U18518 (N_18518,N_17755,N_16947);
nor U18519 (N_18519,N_17178,N_17156);
xor U18520 (N_18520,N_17365,N_17380);
nor U18521 (N_18521,N_17193,N_17520);
nor U18522 (N_18522,N_17081,N_17567);
or U18523 (N_18523,N_17551,N_17907);
and U18524 (N_18524,N_17336,N_17965);
or U18525 (N_18525,N_17865,N_16897);
xnor U18526 (N_18526,N_17337,N_17935);
xnor U18527 (N_18527,N_16914,N_17341);
xnor U18528 (N_18528,N_17117,N_17325);
nand U18529 (N_18529,N_16937,N_17279);
nand U18530 (N_18530,N_16994,N_17171);
xnor U18531 (N_18531,N_17214,N_17073);
xor U18532 (N_18532,N_16963,N_17162);
nand U18533 (N_18533,N_17531,N_17727);
or U18534 (N_18534,N_17408,N_17942);
nor U18535 (N_18535,N_17822,N_16806);
or U18536 (N_18536,N_17301,N_17479);
or U18537 (N_18537,N_17093,N_17557);
nand U18538 (N_18538,N_16949,N_16935);
xor U18539 (N_18539,N_16919,N_17602);
xor U18540 (N_18540,N_17360,N_17180);
nand U18541 (N_18541,N_17573,N_17507);
xor U18542 (N_18542,N_17347,N_17399);
xor U18543 (N_18543,N_17179,N_17532);
nor U18544 (N_18544,N_17930,N_17431);
or U18545 (N_18545,N_17166,N_17055);
xnor U18546 (N_18546,N_17910,N_17563);
nor U18547 (N_18547,N_17858,N_17638);
nor U18548 (N_18548,N_17470,N_17827);
nand U18549 (N_18549,N_17071,N_17576);
xnor U18550 (N_18550,N_17295,N_17019);
and U18551 (N_18551,N_17722,N_17101);
and U18552 (N_18552,N_16969,N_17644);
nor U18553 (N_18553,N_17839,N_17141);
nor U18554 (N_18554,N_17680,N_17530);
xnor U18555 (N_18555,N_17332,N_17287);
and U18556 (N_18556,N_17204,N_17899);
xor U18557 (N_18557,N_17131,N_17236);
nor U18558 (N_18558,N_16828,N_17785);
nor U18559 (N_18559,N_17344,N_16817);
and U18560 (N_18560,N_17854,N_17037);
or U18561 (N_18561,N_17773,N_17752);
and U18562 (N_18562,N_17747,N_17158);
nor U18563 (N_18563,N_17888,N_17099);
nand U18564 (N_18564,N_17262,N_17605);
nand U18565 (N_18565,N_17161,N_17069);
nand U18566 (N_18566,N_17931,N_17622);
or U18567 (N_18567,N_16921,N_17708);
or U18568 (N_18568,N_17683,N_17886);
nor U18569 (N_18569,N_17975,N_17438);
xor U18570 (N_18570,N_17495,N_17017);
xnor U18571 (N_18571,N_17057,N_17437);
or U18572 (N_18572,N_17451,N_17698);
nor U18573 (N_18573,N_17145,N_17737);
or U18574 (N_18574,N_16836,N_17217);
nor U18575 (N_18575,N_17211,N_17802);
and U18576 (N_18576,N_17981,N_17695);
xor U18577 (N_18577,N_17536,N_17781);
nor U18578 (N_18578,N_17107,N_17410);
or U18579 (N_18579,N_17026,N_17776);
and U18580 (N_18580,N_17450,N_17294);
and U18581 (N_18581,N_17186,N_16974);
nand U18582 (N_18582,N_17289,N_17215);
and U18583 (N_18583,N_17187,N_17616);
nor U18584 (N_18584,N_16912,N_17636);
xnor U18585 (N_18585,N_17763,N_17676);
xnor U18586 (N_18586,N_17376,N_17452);
xnor U18587 (N_18587,N_17621,N_17064);
nand U18588 (N_18588,N_16928,N_17501);
xnor U18589 (N_18589,N_17674,N_17515);
and U18590 (N_18590,N_17102,N_17712);
nor U18591 (N_18591,N_17478,N_17445);
nor U18592 (N_18592,N_17679,N_17867);
nand U18593 (N_18593,N_17074,N_17135);
xnor U18594 (N_18594,N_17475,N_17137);
or U18595 (N_18595,N_17146,N_17904);
nor U18596 (N_18596,N_16800,N_17740);
or U18597 (N_18597,N_17415,N_17963);
nand U18598 (N_18598,N_17027,N_17830);
or U18599 (N_18599,N_17555,N_17133);
and U18600 (N_18600,N_17089,N_17221);
nand U18601 (N_18601,N_17952,N_17884);
xnor U18602 (N_18602,N_16999,N_17898);
nand U18603 (N_18603,N_17651,N_17537);
or U18604 (N_18604,N_17318,N_17319);
nand U18605 (N_18605,N_17718,N_17394);
nor U18606 (N_18606,N_17472,N_17956);
and U18607 (N_18607,N_17294,N_17035);
nand U18608 (N_18608,N_16813,N_17136);
and U18609 (N_18609,N_17740,N_17784);
and U18610 (N_18610,N_17825,N_17592);
and U18611 (N_18611,N_17472,N_17744);
xnor U18612 (N_18612,N_17377,N_17418);
xor U18613 (N_18613,N_17231,N_17133);
nor U18614 (N_18614,N_17769,N_17539);
nand U18615 (N_18615,N_17287,N_16857);
nand U18616 (N_18616,N_16907,N_17129);
and U18617 (N_18617,N_17099,N_16803);
nand U18618 (N_18618,N_16971,N_17736);
or U18619 (N_18619,N_17392,N_17246);
nand U18620 (N_18620,N_17132,N_17680);
nand U18621 (N_18621,N_17509,N_16900);
or U18622 (N_18622,N_17896,N_17330);
nor U18623 (N_18623,N_17719,N_17341);
or U18624 (N_18624,N_17911,N_16800);
nand U18625 (N_18625,N_16886,N_17311);
or U18626 (N_18626,N_17350,N_17287);
nor U18627 (N_18627,N_17477,N_17177);
nand U18628 (N_18628,N_17334,N_17207);
nand U18629 (N_18629,N_17857,N_17552);
nor U18630 (N_18630,N_17312,N_17470);
xor U18631 (N_18631,N_16943,N_17560);
xor U18632 (N_18632,N_17959,N_17453);
xor U18633 (N_18633,N_16909,N_16850);
xor U18634 (N_18634,N_17177,N_17036);
or U18635 (N_18635,N_17517,N_16858);
xor U18636 (N_18636,N_17714,N_17175);
and U18637 (N_18637,N_17354,N_17374);
xnor U18638 (N_18638,N_17928,N_17838);
or U18639 (N_18639,N_17811,N_17292);
and U18640 (N_18640,N_17188,N_17261);
or U18641 (N_18641,N_17081,N_17897);
nor U18642 (N_18642,N_17995,N_17659);
and U18643 (N_18643,N_17708,N_17940);
or U18644 (N_18644,N_17957,N_17541);
xnor U18645 (N_18645,N_17192,N_16913);
nand U18646 (N_18646,N_17419,N_16884);
and U18647 (N_18647,N_16963,N_17786);
nand U18648 (N_18648,N_17345,N_17153);
and U18649 (N_18649,N_17605,N_17835);
nor U18650 (N_18650,N_17887,N_17213);
nand U18651 (N_18651,N_16958,N_16968);
or U18652 (N_18652,N_17884,N_17528);
xnor U18653 (N_18653,N_17303,N_17500);
nand U18654 (N_18654,N_17642,N_17392);
xnor U18655 (N_18655,N_17422,N_17751);
nor U18656 (N_18656,N_17932,N_17616);
nor U18657 (N_18657,N_17761,N_17944);
and U18658 (N_18658,N_17129,N_17327);
xor U18659 (N_18659,N_17861,N_17725);
and U18660 (N_18660,N_17086,N_17522);
or U18661 (N_18661,N_17740,N_17813);
nand U18662 (N_18662,N_17976,N_17676);
or U18663 (N_18663,N_17987,N_17744);
xor U18664 (N_18664,N_17163,N_17055);
nand U18665 (N_18665,N_17804,N_17455);
nand U18666 (N_18666,N_17528,N_17057);
xnor U18667 (N_18667,N_17629,N_16869);
xor U18668 (N_18668,N_17807,N_17392);
xnor U18669 (N_18669,N_17985,N_17223);
and U18670 (N_18670,N_17884,N_17795);
xor U18671 (N_18671,N_17449,N_17818);
xnor U18672 (N_18672,N_16990,N_17958);
or U18673 (N_18673,N_16912,N_17208);
and U18674 (N_18674,N_17735,N_17877);
xnor U18675 (N_18675,N_17151,N_17662);
nor U18676 (N_18676,N_17413,N_17500);
or U18677 (N_18677,N_17573,N_17205);
and U18678 (N_18678,N_16914,N_17467);
nand U18679 (N_18679,N_17379,N_17044);
nor U18680 (N_18680,N_17335,N_17823);
nor U18681 (N_18681,N_16865,N_17025);
xor U18682 (N_18682,N_17046,N_17121);
or U18683 (N_18683,N_17246,N_17835);
nor U18684 (N_18684,N_17552,N_17689);
or U18685 (N_18685,N_17854,N_17478);
or U18686 (N_18686,N_17639,N_17066);
xor U18687 (N_18687,N_17875,N_17957);
nand U18688 (N_18688,N_17318,N_17503);
nand U18689 (N_18689,N_17915,N_17964);
and U18690 (N_18690,N_17761,N_16936);
xor U18691 (N_18691,N_17370,N_17296);
nor U18692 (N_18692,N_17183,N_17292);
or U18693 (N_18693,N_16868,N_17057);
and U18694 (N_18694,N_17087,N_17546);
nand U18695 (N_18695,N_17125,N_17185);
nor U18696 (N_18696,N_17376,N_16921);
nor U18697 (N_18697,N_16924,N_17540);
xnor U18698 (N_18698,N_17786,N_16863);
nand U18699 (N_18699,N_17272,N_17176);
or U18700 (N_18700,N_17094,N_17943);
xor U18701 (N_18701,N_17910,N_17171);
xor U18702 (N_18702,N_17048,N_17143);
nand U18703 (N_18703,N_17660,N_17237);
xor U18704 (N_18704,N_16989,N_17205);
and U18705 (N_18705,N_16800,N_17887);
nand U18706 (N_18706,N_17161,N_17043);
xor U18707 (N_18707,N_17180,N_17061);
xor U18708 (N_18708,N_16979,N_16889);
and U18709 (N_18709,N_17070,N_16818);
xor U18710 (N_18710,N_17925,N_17151);
and U18711 (N_18711,N_17847,N_17818);
or U18712 (N_18712,N_17942,N_17323);
nor U18713 (N_18713,N_17250,N_17756);
or U18714 (N_18714,N_17860,N_17947);
or U18715 (N_18715,N_17170,N_17108);
and U18716 (N_18716,N_16820,N_17328);
nand U18717 (N_18717,N_17157,N_17423);
or U18718 (N_18718,N_17224,N_17367);
xor U18719 (N_18719,N_16857,N_17140);
nor U18720 (N_18720,N_17222,N_17896);
nand U18721 (N_18721,N_17206,N_17351);
xnor U18722 (N_18722,N_17931,N_17718);
nand U18723 (N_18723,N_17620,N_17026);
nor U18724 (N_18724,N_17920,N_16998);
and U18725 (N_18725,N_17529,N_17341);
or U18726 (N_18726,N_17008,N_17480);
xor U18727 (N_18727,N_17795,N_17763);
xnor U18728 (N_18728,N_17105,N_17311);
xor U18729 (N_18729,N_17724,N_17760);
nor U18730 (N_18730,N_17638,N_17920);
nor U18731 (N_18731,N_17953,N_17605);
nand U18732 (N_18732,N_17854,N_16869);
nor U18733 (N_18733,N_17014,N_17675);
or U18734 (N_18734,N_17326,N_17327);
and U18735 (N_18735,N_17123,N_16979);
or U18736 (N_18736,N_17121,N_17722);
nand U18737 (N_18737,N_17577,N_17119);
nor U18738 (N_18738,N_16970,N_17755);
nor U18739 (N_18739,N_17094,N_17716);
and U18740 (N_18740,N_17503,N_17397);
and U18741 (N_18741,N_17392,N_17558);
nor U18742 (N_18742,N_17489,N_17539);
or U18743 (N_18743,N_16816,N_17687);
and U18744 (N_18744,N_17610,N_17186);
or U18745 (N_18745,N_17012,N_16864);
and U18746 (N_18746,N_17599,N_17571);
nor U18747 (N_18747,N_17273,N_17079);
or U18748 (N_18748,N_17714,N_17782);
nor U18749 (N_18749,N_16830,N_17403);
xnor U18750 (N_18750,N_17822,N_17977);
xor U18751 (N_18751,N_17608,N_17370);
or U18752 (N_18752,N_17530,N_17148);
xnor U18753 (N_18753,N_16969,N_17677);
nand U18754 (N_18754,N_16899,N_17914);
nor U18755 (N_18755,N_17266,N_17628);
nand U18756 (N_18756,N_17838,N_17344);
nor U18757 (N_18757,N_17481,N_17121);
xnor U18758 (N_18758,N_17019,N_17979);
nand U18759 (N_18759,N_17929,N_17289);
nand U18760 (N_18760,N_17964,N_17747);
and U18761 (N_18761,N_17724,N_17983);
and U18762 (N_18762,N_17928,N_17286);
nand U18763 (N_18763,N_16862,N_17415);
nand U18764 (N_18764,N_17081,N_17389);
nand U18765 (N_18765,N_17188,N_16912);
and U18766 (N_18766,N_16837,N_16966);
nand U18767 (N_18767,N_16865,N_17222);
xnor U18768 (N_18768,N_17691,N_17157);
or U18769 (N_18769,N_17440,N_17622);
nor U18770 (N_18770,N_17405,N_16852);
and U18771 (N_18771,N_17688,N_17162);
xnor U18772 (N_18772,N_17613,N_17963);
nand U18773 (N_18773,N_17649,N_16992);
xnor U18774 (N_18774,N_17004,N_17536);
xnor U18775 (N_18775,N_16839,N_17577);
nor U18776 (N_18776,N_16903,N_17227);
nand U18777 (N_18777,N_17085,N_16949);
and U18778 (N_18778,N_17206,N_17289);
and U18779 (N_18779,N_17059,N_17957);
nor U18780 (N_18780,N_17097,N_17585);
nand U18781 (N_18781,N_16914,N_17238);
xnor U18782 (N_18782,N_17426,N_17050);
xnor U18783 (N_18783,N_17644,N_17419);
nand U18784 (N_18784,N_17625,N_17124);
xor U18785 (N_18785,N_16831,N_17241);
and U18786 (N_18786,N_17949,N_17692);
nor U18787 (N_18787,N_16913,N_17603);
nand U18788 (N_18788,N_17564,N_17276);
nand U18789 (N_18789,N_17509,N_17630);
and U18790 (N_18790,N_17047,N_16884);
and U18791 (N_18791,N_17417,N_17630);
nor U18792 (N_18792,N_16884,N_16906);
nand U18793 (N_18793,N_17701,N_17523);
or U18794 (N_18794,N_17600,N_17772);
xor U18795 (N_18795,N_17295,N_17064);
xor U18796 (N_18796,N_17391,N_17760);
nor U18797 (N_18797,N_17018,N_17069);
or U18798 (N_18798,N_17849,N_17474);
nand U18799 (N_18799,N_17402,N_17844);
nor U18800 (N_18800,N_17008,N_17887);
and U18801 (N_18801,N_17347,N_17257);
or U18802 (N_18802,N_17648,N_17427);
or U18803 (N_18803,N_17182,N_17151);
or U18804 (N_18804,N_17589,N_17705);
xor U18805 (N_18805,N_17186,N_17409);
and U18806 (N_18806,N_17369,N_16909);
xnor U18807 (N_18807,N_16865,N_17442);
nand U18808 (N_18808,N_16980,N_17806);
and U18809 (N_18809,N_17235,N_17668);
xnor U18810 (N_18810,N_17579,N_17288);
nand U18811 (N_18811,N_17779,N_17636);
nand U18812 (N_18812,N_17596,N_17402);
and U18813 (N_18813,N_17659,N_17805);
and U18814 (N_18814,N_17369,N_17819);
nand U18815 (N_18815,N_17275,N_17256);
nand U18816 (N_18816,N_17352,N_17445);
nand U18817 (N_18817,N_16863,N_17496);
xor U18818 (N_18818,N_16816,N_17355);
nor U18819 (N_18819,N_16893,N_17388);
nand U18820 (N_18820,N_17799,N_17585);
nand U18821 (N_18821,N_16949,N_17077);
and U18822 (N_18822,N_17655,N_17016);
nand U18823 (N_18823,N_17267,N_17215);
or U18824 (N_18824,N_17241,N_16997);
xor U18825 (N_18825,N_17810,N_17474);
xor U18826 (N_18826,N_17735,N_17646);
nor U18827 (N_18827,N_17432,N_16943);
nand U18828 (N_18828,N_17097,N_16884);
xnor U18829 (N_18829,N_17025,N_17927);
nor U18830 (N_18830,N_16803,N_17486);
nor U18831 (N_18831,N_17536,N_16858);
or U18832 (N_18832,N_17401,N_17269);
nand U18833 (N_18833,N_16982,N_17274);
xor U18834 (N_18834,N_16877,N_17009);
or U18835 (N_18835,N_17073,N_17388);
xnor U18836 (N_18836,N_17074,N_16858);
or U18837 (N_18837,N_17654,N_17423);
nand U18838 (N_18838,N_17800,N_17512);
nand U18839 (N_18839,N_17537,N_16869);
nand U18840 (N_18840,N_17087,N_17130);
xor U18841 (N_18841,N_17913,N_17114);
and U18842 (N_18842,N_17220,N_17308);
and U18843 (N_18843,N_17593,N_17484);
nand U18844 (N_18844,N_17425,N_16917);
or U18845 (N_18845,N_17649,N_17518);
nand U18846 (N_18846,N_17848,N_17273);
nand U18847 (N_18847,N_16907,N_16893);
and U18848 (N_18848,N_16924,N_17713);
and U18849 (N_18849,N_17686,N_17993);
or U18850 (N_18850,N_17118,N_17247);
and U18851 (N_18851,N_17788,N_17850);
nor U18852 (N_18852,N_17644,N_17086);
and U18853 (N_18853,N_17469,N_17855);
nand U18854 (N_18854,N_17684,N_16867);
or U18855 (N_18855,N_17429,N_17396);
xor U18856 (N_18856,N_17620,N_17963);
nand U18857 (N_18857,N_17139,N_17960);
nor U18858 (N_18858,N_17371,N_17190);
xnor U18859 (N_18859,N_17263,N_17041);
nand U18860 (N_18860,N_17509,N_17007);
or U18861 (N_18861,N_17700,N_17640);
and U18862 (N_18862,N_17848,N_17168);
xor U18863 (N_18863,N_17879,N_16815);
nor U18864 (N_18864,N_17230,N_17605);
and U18865 (N_18865,N_17242,N_17663);
nand U18866 (N_18866,N_17019,N_17788);
nor U18867 (N_18867,N_17623,N_17987);
xnor U18868 (N_18868,N_17467,N_17942);
nor U18869 (N_18869,N_17564,N_17791);
xnor U18870 (N_18870,N_17635,N_17302);
or U18871 (N_18871,N_16946,N_16976);
nand U18872 (N_18872,N_17501,N_17119);
xnor U18873 (N_18873,N_17920,N_17623);
nor U18874 (N_18874,N_17667,N_17415);
xnor U18875 (N_18875,N_17620,N_17222);
nand U18876 (N_18876,N_17115,N_16922);
nor U18877 (N_18877,N_17741,N_16854);
or U18878 (N_18878,N_17140,N_16838);
nand U18879 (N_18879,N_17624,N_17685);
or U18880 (N_18880,N_17580,N_17854);
and U18881 (N_18881,N_17857,N_16891);
or U18882 (N_18882,N_17922,N_17108);
and U18883 (N_18883,N_17601,N_17508);
and U18884 (N_18884,N_17103,N_16807);
xor U18885 (N_18885,N_17871,N_17013);
nor U18886 (N_18886,N_17334,N_17655);
nor U18887 (N_18887,N_17836,N_17053);
nand U18888 (N_18888,N_17768,N_17508);
nor U18889 (N_18889,N_17521,N_16928);
and U18890 (N_18890,N_17475,N_17331);
or U18891 (N_18891,N_17236,N_17624);
or U18892 (N_18892,N_17587,N_17915);
xnor U18893 (N_18893,N_17099,N_17235);
and U18894 (N_18894,N_17058,N_17523);
or U18895 (N_18895,N_17788,N_17837);
nor U18896 (N_18896,N_17935,N_17157);
nand U18897 (N_18897,N_17201,N_17217);
and U18898 (N_18898,N_17491,N_17881);
or U18899 (N_18899,N_17614,N_17057);
and U18900 (N_18900,N_17550,N_17809);
xnor U18901 (N_18901,N_16964,N_17028);
nor U18902 (N_18902,N_17016,N_17591);
xor U18903 (N_18903,N_17253,N_17094);
xor U18904 (N_18904,N_17047,N_17592);
and U18905 (N_18905,N_17656,N_17326);
and U18906 (N_18906,N_16911,N_17313);
and U18907 (N_18907,N_17189,N_17420);
or U18908 (N_18908,N_17893,N_17348);
or U18909 (N_18909,N_17319,N_17731);
or U18910 (N_18910,N_17532,N_17055);
or U18911 (N_18911,N_17542,N_17263);
xor U18912 (N_18912,N_17193,N_17263);
nand U18913 (N_18913,N_17831,N_17084);
nor U18914 (N_18914,N_17793,N_17797);
and U18915 (N_18915,N_17244,N_16822);
nor U18916 (N_18916,N_17373,N_17524);
or U18917 (N_18917,N_17900,N_17119);
and U18918 (N_18918,N_17752,N_16827);
and U18919 (N_18919,N_17024,N_17301);
nand U18920 (N_18920,N_17590,N_17921);
or U18921 (N_18921,N_16982,N_17719);
nand U18922 (N_18922,N_17137,N_17252);
or U18923 (N_18923,N_16919,N_17591);
and U18924 (N_18924,N_17109,N_17735);
xor U18925 (N_18925,N_16884,N_17058);
nand U18926 (N_18926,N_17390,N_17282);
nor U18927 (N_18927,N_17973,N_17224);
or U18928 (N_18928,N_17762,N_17432);
nor U18929 (N_18929,N_17157,N_17652);
or U18930 (N_18930,N_17123,N_17875);
nand U18931 (N_18931,N_17798,N_17120);
nor U18932 (N_18932,N_17631,N_17904);
nand U18933 (N_18933,N_17258,N_17716);
and U18934 (N_18934,N_17201,N_17931);
nand U18935 (N_18935,N_17818,N_17727);
nor U18936 (N_18936,N_17207,N_17301);
and U18937 (N_18937,N_17950,N_16884);
nor U18938 (N_18938,N_17306,N_17925);
xnor U18939 (N_18939,N_16861,N_17732);
xor U18940 (N_18940,N_17614,N_16817);
nand U18941 (N_18941,N_17574,N_16820);
or U18942 (N_18942,N_17286,N_17846);
or U18943 (N_18943,N_17261,N_17137);
or U18944 (N_18944,N_17630,N_16905);
nand U18945 (N_18945,N_17688,N_17939);
xor U18946 (N_18946,N_17340,N_17525);
and U18947 (N_18947,N_17530,N_17473);
nand U18948 (N_18948,N_17808,N_17234);
and U18949 (N_18949,N_17605,N_16831);
or U18950 (N_18950,N_17339,N_17090);
xnor U18951 (N_18951,N_17775,N_17376);
or U18952 (N_18952,N_16986,N_17570);
or U18953 (N_18953,N_16935,N_17892);
or U18954 (N_18954,N_17430,N_17682);
nand U18955 (N_18955,N_17188,N_17708);
or U18956 (N_18956,N_16800,N_17028);
xnor U18957 (N_18957,N_17361,N_17299);
xor U18958 (N_18958,N_17088,N_17705);
nand U18959 (N_18959,N_17918,N_16876);
nand U18960 (N_18960,N_17967,N_17732);
and U18961 (N_18961,N_17493,N_17588);
xor U18962 (N_18962,N_17624,N_17552);
xnor U18963 (N_18963,N_17199,N_17176);
and U18964 (N_18964,N_17705,N_17306);
nor U18965 (N_18965,N_17892,N_16996);
nor U18966 (N_18966,N_17014,N_17712);
xnor U18967 (N_18967,N_16942,N_16995);
nand U18968 (N_18968,N_17973,N_17502);
or U18969 (N_18969,N_16969,N_17808);
or U18970 (N_18970,N_17741,N_17369);
nand U18971 (N_18971,N_17867,N_17020);
xnor U18972 (N_18972,N_17866,N_17555);
nand U18973 (N_18973,N_17448,N_17095);
and U18974 (N_18974,N_17225,N_17878);
nand U18975 (N_18975,N_17128,N_17426);
or U18976 (N_18976,N_17565,N_17503);
and U18977 (N_18977,N_17250,N_16844);
xnor U18978 (N_18978,N_17422,N_16913);
nand U18979 (N_18979,N_17441,N_16960);
and U18980 (N_18980,N_17713,N_16929);
xnor U18981 (N_18981,N_17155,N_17752);
nand U18982 (N_18982,N_17108,N_17296);
nor U18983 (N_18983,N_17147,N_17815);
and U18984 (N_18984,N_17906,N_17362);
or U18985 (N_18985,N_17871,N_17770);
and U18986 (N_18986,N_17584,N_17902);
or U18987 (N_18987,N_16883,N_17383);
nor U18988 (N_18988,N_17827,N_16889);
and U18989 (N_18989,N_17216,N_16811);
xor U18990 (N_18990,N_17303,N_17160);
and U18991 (N_18991,N_17527,N_16963);
nor U18992 (N_18992,N_17035,N_16843);
and U18993 (N_18993,N_17205,N_17385);
nand U18994 (N_18994,N_17782,N_17486);
xnor U18995 (N_18995,N_17193,N_16992);
nor U18996 (N_18996,N_17181,N_17547);
nand U18997 (N_18997,N_17271,N_17501);
nor U18998 (N_18998,N_17382,N_17326);
nor U18999 (N_18999,N_17294,N_17399);
nand U19000 (N_19000,N_17231,N_16888);
and U19001 (N_19001,N_17892,N_17889);
nor U19002 (N_19002,N_17623,N_17436);
nor U19003 (N_19003,N_17955,N_17295);
xor U19004 (N_19004,N_17557,N_17288);
nand U19005 (N_19005,N_17633,N_17641);
xor U19006 (N_19006,N_16864,N_17053);
and U19007 (N_19007,N_16972,N_17999);
nand U19008 (N_19008,N_17516,N_17207);
xnor U19009 (N_19009,N_17849,N_17916);
and U19010 (N_19010,N_17474,N_17811);
and U19011 (N_19011,N_16957,N_17449);
nor U19012 (N_19012,N_17977,N_16974);
nand U19013 (N_19013,N_17485,N_17043);
or U19014 (N_19014,N_17113,N_17360);
xor U19015 (N_19015,N_17312,N_17670);
nor U19016 (N_19016,N_17502,N_17111);
nand U19017 (N_19017,N_17506,N_17598);
xor U19018 (N_19018,N_17806,N_17218);
nand U19019 (N_19019,N_16851,N_17566);
or U19020 (N_19020,N_17798,N_17008);
or U19021 (N_19021,N_17565,N_17699);
and U19022 (N_19022,N_17667,N_17556);
nand U19023 (N_19023,N_17707,N_17010);
nand U19024 (N_19024,N_17633,N_17743);
and U19025 (N_19025,N_17372,N_17405);
or U19026 (N_19026,N_17415,N_17847);
xnor U19027 (N_19027,N_17248,N_16965);
xnor U19028 (N_19028,N_16845,N_16899);
or U19029 (N_19029,N_17599,N_17354);
nor U19030 (N_19030,N_17662,N_17106);
and U19031 (N_19031,N_17347,N_17494);
or U19032 (N_19032,N_17807,N_17794);
or U19033 (N_19033,N_17997,N_17295);
or U19034 (N_19034,N_16925,N_16892);
or U19035 (N_19035,N_17981,N_17982);
or U19036 (N_19036,N_17154,N_17070);
or U19037 (N_19037,N_17056,N_17346);
or U19038 (N_19038,N_17435,N_17019);
nor U19039 (N_19039,N_17465,N_17484);
nor U19040 (N_19040,N_17910,N_17194);
xnor U19041 (N_19041,N_17735,N_17476);
nor U19042 (N_19042,N_17695,N_17398);
and U19043 (N_19043,N_16877,N_17260);
xnor U19044 (N_19044,N_17814,N_17112);
nand U19045 (N_19045,N_17027,N_17019);
xnor U19046 (N_19046,N_17464,N_17045);
or U19047 (N_19047,N_16929,N_17040);
nor U19048 (N_19048,N_16846,N_17684);
nor U19049 (N_19049,N_16932,N_17749);
nor U19050 (N_19050,N_17969,N_17829);
and U19051 (N_19051,N_17042,N_17053);
or U19052 (N_19052,N_17291,N_17574);
or U19053 (N_19053,N_16843,N_17445);
or U19054 (N_19054,N_17341,N_17392);
or U19055 (N_19055,N_17002,N_17082);
and U19056 (N_19056,N_17633,N_17026);
nand U19057 (N_19057,N_17579,N_17368);
nand U19058 (N_19058,N_17167,N_17928);
nor U19059 (N_19059,N_17586,N_16900);
nor U19060 (N_19060,N_17663,N_17293);
nand U19061 (N_19061,N_16991,N_17028);
nand U19062 (N_19062,N_16966,N_17926);
or U19063 (N_19063,N_17559,N_16876);
nor U19064 (N_19064,N_17148,N_16827);
and U19065 (N_19065,N_17761,N_17214);
and U19066 (N_19066,N_16913,N_17444);
nor U19067 (N_19067,N_17713,N_17246);
or U19068 (N_19068,N_17687,N_17430);
xnor U19069 (N_19069,N_17434,N_16946);
or U19070 (N_19070,N_17842,N_17636);
nand U19071 (N_19071,N_17005,N_17478);
nor U19072 (N_19072,N_16838,N_16979);
nand U19073 (N_19073,N_17370,N_17439);
or U19074 (N_19074,N_17086,N_17811);
xor U19075 (N_19075,N_17935,N_17801);
or U19076 (N_19076,N_17992,N_17352);
and U19077 (N_19077,N_17666,N_17705);
xnor U19078 (N_19078,N_17472,N_17278);
and U19079 (N_19079,N_17335,N_17344);
xnor U19080 (N_19080,N_17276,N_16995);
xor U19081 (N_19081,N_17099,N_17052);
and U19082 (N_19082,N_17394,N_17000);
and U19083 (N_19083,N_17141,N_17959);
nand U19084 (N_19084,N_16917,N_17695);
nor U19085 (N_19085,N_17048,N_17492);
nor U19086 (N_19086,N_17390,N_17770);
and U19087 (N_19087,N_17737,N_17711);
or U19088 (N_19088,N_17326,N_16894);
nand U19089 (N_19089,N_17061,N_16890);
xor U19090 (N_19090,N_17292,N_17971);
and U19091 (N_19091,N_17266,N_17866);
nand U19092 (N_19092,N_17225,N_16802);
nand U19093 (N_19093,N_16967,N_17781);
nor U19094 (N_19094,N_16879,N_17039);
nand U19095 (N_19095,N_17957,N_17480);
nor U19096 (N_19096,N_17675,N_17600);
nand U19097 (N_19097,N_17525,N_17564);
nand U19098 (N_19098,N_17172,N_17977);
or U19099 (N_19099,N_16986,N_17381);
xor U19100 (N_19100,N_17718,N_17470);
and U19101 (N_19101,N_17341,N_17705);
or U19102 (N_19102,N_16962,N_17173);
xnor U19103 (N_19103,N_17855,N_17092);
nand U19104 (N_19104,N_17042,N_17521);
or U19105 (N_19105,N_17909,N_16954);
nor U19106 (N_19106,N_17169,N_17306);
and U19107 (N_19107,N_17494,N_17195);
xnor U19108 (N_19108,N_17205,N_17365);
or U19109 (N_19109,N_17426,N_17665);
nor U19110 (N_19110,N_17532,N_17197);
nand U19111 (N_19111,N_17073,N_17121);
nand U19112 (N_19112,N_16976,N_17501);
nand U19113 (N_19113,N_17455,N_17851);
nand U19114 (N_19114,N_17019,N_17947);
and U19115 (N_19115,N_17583,N_16890);
or U19116 (N_19116,N_17622,N_17618);
xnor U19117 (N_19117,N_17319,N_17702);
nand U19118 (N_19118,N_17241,N_17492);
or U19119 (N_19119,N_17661,N_17366);
nand U19120 (N_19120,N_16807,N_16938);
xnor U19121 (N_19121,N_16905,N_17892);
nand U19122 (N_19122,N_17149,N_17237);
nand U19123 (N_19123,N_17675,N_17146);
xor U19124 (N_19124,N_17732,N_17425);
nor U19125 (N_19125,N_17706,N_17656);
or U19126 (N_19126,N_17404,N_17070);
nand U19127 (N_19127,N_17309,N_17645);
or U19128 (N_19128,N_17107,N_17404);
nor U19129 (N_19129,N_17805,N_17879);
xnor U19130 (N_19130,N_17959,N_17848);
and U19131 (N_19131,N_17695,N_17530);
or U19132 (N_19132,N_17416,N_16914);
and U19133 (N_19133,N_17623,N_17163);
nor U19134 (N_19134,N_17202,N_17250);
xor U19135 (N_19135,N_17831,N_17945);
and U19136 (N_19136,N_17300,N_17606);
and U19137 (N_19137,N_17715,N_17438);
or U19138 (N_19138,N_17495,N_17823);
or U19139 (N_19139,N_17247,N_17687);
nand U19140 (N_19140,N_17971,N_16853);
nand U19141 (N_19141,N_17329,N_17694);
and U19142 (N_19142,N_17233,N_17648);
nand U19143 (N_19143,N_17837,N_17740);
nand U19144 (N_19144,N_17458,N_17349);
or U19145 (N_19145,N_17052,N_17104);
xnor U19146 (N_19146,N_16853,N_17706);
nor U19147 (N_19147,N_17095,N_17379);
and U19148 (N_19148,N_17160,N_17683);
nor U19149 (N_19149,N_17567,N_17339);
and U19150 (N_19150,N_17048,N_17861);
or U19151 (N_19151,N_17993,N_17893);
and U19152 (N_19152,N_17634,N_17916);
and U19153 (N_19153,N_17394,N_16993);
nor U19154 (N_19154,N_17160,N_17542);
xor U19155 (N_19155,N_17662,N_17673);
and U19156 (N_19156,N_17853,N_17058);
nor U19157 (N_19157,N_16824,N_17745);
or U19158 (N_19158,N_16945,N_17083);
nand U19159 (N_19159,N_16982,N_17462);
xor U19160 (N_19160,N_16838,N_16802);
nor U19161 (N_19161,N_16880,N_16896);
or U19162 (N_19162,N_16860,N_17547);
nand U19163 (N_19163,N_17500,N_17774);
nor U19164 (N_19164,N_17857,N_17332);
and U19165 (N_19165,N_17460,N_17386);
nand U19166 (N_19166,N_17689,N_17543);
and U19167 (N_19167,N_17890,N_17968);
nand U19168 (N_19168,N_17376,N_17130);
or U19169 (N_19169,N_17652,N_17696);
nand U19170 (N_19170,N_17213,N_17455);
nor U19171 (N_19171,N_17756,N_17027);
nand U19172 (N_19172,N_17047,N_17505);
nand U19173 (N_19173,N_16996,N_16901);
or U19174 (N_19174,N_17142,N_17837);
nand U19175 (N_19175,N_17274,N_17859);
nand U19176 (N_19176,N_17038,N_17155);
xnor U19177 (N_19177,N_17887,N_17421);
or U19178 (N_19178,N_17843,N_17552);
or U19179 (N_19179,N_17552,N_16955);
and U19180 (N_19180,N_16883,N_17511);
nand U19181 (N_19181,N_17933,N_17910);
xnor U19182 (N_19182,N_17775,N_17320);
nor U19183 (N_19183,N_17356,N_16806);
xnor U19184 (N_19184,N_17636,N_16965);
or U19185 (N_19185,N_16848,N_17281);
nand U19186 (N_19186,N_16907,N_17214);
nand U19187 (N_19187,N_17969,N_17607);
nor U19188 (N_19188,N_17472,N_17290);
nor U19189 (N_19189,N_17703,N_17940);
or U19190 (N_19190,N_17408,N_17155);
and U19191 (N_19191,N_17302,N_17998);
nand U19192 (N_19192,N_17199,N_17156);
nand U19193 (N_19193,N_16895,N_17886);
and U19194 (N_19194,N_17738,N_17218);
or U19195 (N_19195,N_17868,N_17203);
and U19196 (N_19196,N_17452,N_17306);
or U19197 (N_19197,N_17331,N_17551);
nand U19198 (N_19198,N_17699,N_17445);
and U19199 (N_19199,N_17427,N_17041);
or U19200 (N_19200,N_18048,N_18895);
xnor U19201 (N_19201,N_18778,N_19119);
nor U19202 (N_19202,N_18704,N_18663);
or U19203 (N_19203,N_18904,N_18572);
and U19204 (N_19204,N_18364,N_19142);
nand U19205 (N_19205,N_18532,N_18246);
nand U19206 (N_19206,N_18398,N_19088);
or U19207 (N_19207,N_18878,N_18910);
xnor U19208 (N_19208,N_18251,N_18823);
nand U19209 (N_19209,N_18130,N_18254);
and U19210 (N_19210,N_18810,N_18026);
xor U19211 (N_19211,N_19063,N_18589);
nand U19212 (N_19212,N_18454,N_18544);
or U19213 (N_19213,N_18703,N_18536);
nor U19214 (N_19214,N_19086,N_18570);
nand U19215 (N_19215,N_18071,N_18047);
or U19216 (N_19216,N_19067,N_18097);
and U19217 (N_19217,N_19039,N_18072);
xor U19218 (N_19218,N_18371,N_18079);
nor U19219 (N_19219,N_18955,N_18060);
xnor U19220 (N_19220,N_18807,N_18978);
nor U19221 (N_19221,N_19055,N_18187);
nor U19222 (N_19222,N_18287,N_18673);
nand U19223 (N_19223,N_18498,N_19087);
nand U19224 (N_19224,N_18992,N_18147);
nor U19225 (N_19225,N_18576,N_18974);
and U19226 (N_19226,N_18273,N_18864);
xor U19227 (N_19227,N_19115,N_18350);
or U19228 (N_19228,N_18947,N_19076);
nand U19229 (N_19229,N_18317,N_18239);
nor U19230 (N_19230,N_18314,N_19168);
nand U19231 (N_19231,N_19125,N_18737);
nor U19232 (N_19232,N_19051,N_18718);
or U19233 (N_19233,N_19126,N_18804);
and U19234 (N_19234,N_18391,N_18897);
and U19235 (N_19235,N_18915,N_18863);
nor U19236 (N_19236,N_18840,N_18386);
nand U19237 (N_19237,N_18330,N_18943);
and U19238 (N_19238,N_18592,N_18946);
nor U19239 (N_19239,N_18902,N_18162);
nor U19240 (N_19240,N_18841,N_19048);
and U19241 (N_19241,N_18159,N_18742);
or U19242 (N_19242,N_18918,N_18074);
nand U19243 (N_19243,N_19189,N_18000);
xor U19244 (N_19244,N_18020,N_18569);
xnor U19245 (N_19245,N_18883,N_18789);
nand U19246 (N_19246,N_18960,N_18443);
xor U19247 (N_19247,N_18420,N_19114);
and U19248 (N_19248,N_18771,N_18610);
nor U19249 (N_19249,N_18647,N_18214);
nand U19250 (N_19250,N_18265,N_18166);
nor U19251 (N_19251,N_19035,N_18855);
nand U19252 (N_19252,N_18300,N_18361);
nor U19253 (N_19253,N_19010,N_18997);
xor U19254 (N_19254,N_18081,N_18792);
xnor U19255 (N_19255,N_18377,N_18332);
and U19256 (N_19256,N_18652,N_18688);
nand U19257 (N_19257,N_18548,N_18764);
xor U19258 (N_19258,N_18579,N_19038);
nor U19259 (N_19259,N_18933,N_18210);
xor U19260 (N_19260,N_18838,N_18581);
and U19261 (N_19261,N_18866,N_19011);
nor U19262 (N_19262,N_18237,N_19057);
and U19263 (N_19263,N_18721,N_18787);
xnor U19264 (N_19264,N_19150,N_18219);
nor U19265 (N_19265,N_18690,N_18945);
and U19266 (N_19266,N_18451,N_18928);
xor U19267 (N_19267,N_18261,N_18406);
or U19268 (N_19268,N_18759,N_18369);
xor U19269 (N_19269,N_18004,N_19000);
nor U19270 (N_19270,N_18888,N_19054);
xnor U19271 (N_19271,N_18289,N_18188);
and U19272 (N_19272,N_19009,N_18158);
or U19273 (N_19273,N_18775,N_18631);
xor U19274 (N_19274,N_18101,N_18687);
and U19275 (N_19275,N_19097,N_18509);
nor U19276 (N_19276,N_18644,N_18661);
nand U19277 (N_19277,N_18348,N_18405);
nor U19278 (N_19278,N_18926,N_18538);
nor U19279 (N_19279,N_19004,N_18235);
xor U19280 (N_19280,N_18231,N_18606);
and U19281 (N_19281,N_18301,N_18357);
nand U19282 (N_19282,N_18018,N_19194);
and U19283 (N_19283,N_19184,N_18880);
nand U19284 (N_19284,N_18599,N_18714);
and U19285 (N_19285,N_18667,N_18095);
xor U19286 (N_19286,N_18138,N_18354);
and U19287 (N_19287,N_18686,N_18797);
and U19288 (N_19288,N_18689,N_18478);
nor U19289 (N_19289,N_18274,N_18500);
or U19290 (N_19290,N_18655,N_19041);
or U19291 (N_19291,N_18799,N_18365);
and U19292 (N_19292,N_19101,N_18476);
and U19293 (N_19293,N_18298,N_18240);
nand U19294 (N_19294,N_19153,N_18335);
and U19295 (N_19295,N_18806,N_19091);
and U19296 (N_19296,N_18447,N_18875);
xor U19297 (N_19297,N_18399,N_18212);
or U19298 (N_19298,N_18215,N_18931);
nand U19299 (N_19299,N_19135,N_18487);
nand U19300 (N_19300,N_18283,N_18845);
and U19301 (N_19301,N_18173,N_18436);
nor U19302 (N_19302,N_18972,N_18626);
nand U19303 (N_19303,N_18144,N_18731);
nor U19304 (N_19304,N_18013,N_18250);
nand U19305 (N_19305,N_18137,N_18347);
or U19306 (N_19306,N_18956,N_18229);
and U19307 (N_19307,N_18205,N_18139);
nor U19308 (N_19308,N_18781,N_19084);
nor U19309 (N_19309,N_18449,N_18675);
nor U19310 (N_19310,N_19136,N_18477);
nor U19311 (N_19311,N_18226,N_18221);
or U19312 (N_19312,N_19112,N_18203);
and U19313 (N_19313,N_18976,N_18574);
nand U19314 (N_19314,N_18729,N_18893);
xnor U19315 (N_19315,N_18257,N_18939);
or U19316 (N_19316,N_18717,N_18899);
xnor U19317 (N_19317,N_18774,N_18488);
or U19318 (N_19318,N_19036,N_18001);
nand U19319 (N_19319,N_18343,N_19198);
and U19320 (N_19320,N_18328,N_18602);
nor U19321 (N_19321,N_18472,N_18925);
nand U19322 (N_19322,N_19175,N_18453);
nor U19323 (N_19323,N_18043,N_18469);
xnor U19324 (N_19324,N_18959,N_18099);
xnor U19325 (N_19325,N_18094,N_18299);
xnor U19326 (N_19326,N_18847,N_18975);
xor U19327 (N_19327,N_18442,N_18812);
or U19328 (N_19328,N_18501,N_18064);
nand U19329 (N_19329,N_18950,N_18770);
or U19330 (N_19330,N_18515,N_19159);
and U19331 (N_19331,N_19116,N_18558);
xor U19332 (N_19332,N_18954,N_19178);
or U19333 (N_19333,N_18940,N_18934);
xnor U19334 (N_19334,N_19082,N_18403);
xnor U19335 (N_19335,N_19158,N_18112);
nand U19336 (N_19336,N_18474,N_18433);
nor U19337 (N_19337,N_18178,N_18148);
xor U19338 (N_19338,N_18596,N_18635);
xor U19339 (N_19339,N_18773,N_18715);
xor U19340 (N_19340,N_18758,N_18522);
xor U19341 (N_19341,N_18304,N_18525);
xor U19342 (N_19342,N_19019,N_18580);
nor U19343 (N_19343,N_18096,N_18879);
nor U19344 (N_19344,N_18963,N_18705);
nor U19345 (N_19345,N_18681,N_18961);
or U19346 (N_19346,N_18901,N_18410);
nand U19347 (N_19347,N_18165,N_18356);
nand U19348 (N_19348,N_19187,N_18666);
nand U19349 (N_19349,N_18149,N_19106);
xnor U19350 (N_19350,N_19154,N_18584);
xor U19351 (N_19351,N_18186,N_18312);
nand U19352 (N_19352,N_18054,N_18857);
nor U19353 (N_19353,N_18832,N_18850);
or U19354 (N_19354,N_18949,N_18649);
nor U19355 (N_19355,N_18877,N_18318);
and U19356 (N_19356,N_18195,N_18286);
xor U19357 (N_19357,N_18869,N_18540);
nor U19358 (N_19358,N_18645,N_18639);
and U19359 (N_19359,N_18769,N_18916);
nand U19360 (N_19360,N_19167,N_18986);
nor U19361 (N_19361,N_18034,N_19129);
or U19362 (N_19362,N_19148,N_18382);
xnor U19363 (N_19363,N_19029,N_18725);
or U19364 (N_19364,N_18973,N_18217);
nor U19365 (N_19365,N_19092,N_18448);
and U19366 (N_19366,N_18983,N_18700);
nor U19367 (N_19367,N_19023,N_18051);
and U19368 (N_19368,N_18208,N_18562);
xnor U19369 (N_19369,N_18414,N_18865);
or U19370 (N_19370,N_18315,N_18751);
nand U19371 (N_19371,N_18222,N_18648);
and U19372 (N_19372,N_19001,N_18282);
xor U19373 (N_19373,N_18499,N_18121);
or U19374 (N_19374,N_19120,N_19103);
nand U19375 (N_19375,N_19065,N_18046);
nor U19376 (N_19376,N_18952,N_18552);
or U19377 (N_19377,N_18791,N_19030);
and U19378 (N_19378,N_19110,N_19068);
xor U19379 (N_19379,N_18783,N_18323);
and U19380 (N_19380,N_18338,N_18884);
nand U19381 (N_19381,N_18225,N_18795);
xnor U19382 (N_19382,N_18193,N_18255);
nor U19383 (N_19383,N_18003,N_18707);
xor U19384 (N_19384,N_18151,N_18846);
and U19385 (N_19385,N_18133,N_18266);
xor U19386 (N_19386,N_19015,N_18669);
xnor U19387 (N_19387,N_18452,N_19170);
or U19388 (N_19388,N_18892,N_19100);
and U19389 (N_19389,N_18609,N_18803);
nor U19390 (N_19390,N_18075,N_18793);
or U19391 (N_19391,N_18612,N_18944);
and U19392 (N_19392,N_18078,N_18413);
or U19393 (N_19393,N_18938,N_18085);
and U19394 (N_19394,N_18042,N_19006);
or U19395 (N_19395,N_18889,N_18749);
nand U19396 (N_19396,N_18668,N_18024);
or U19397 (N_19397,N_19121,N_19107);
nor U19398 (N_19398,N_18362,N_18224);
or U19399 (N_19399,N_18252,N_18571);
xor U19400 (N_19400,N_18062,N_18073);
or U19401 (N_19401,N_18181,N_18912);
nor U19402 (N_19402,N_18288,N_18128);
and U19403 (N_19403,N_18868,N_18007);
nand U19404 (N_19404,N_18141,N_19032);
nor U19405 (N_19405,N_18041,N_18966);
and U19406 (N_19406,N_18844,N_18534);
nand U19407 (N_19407,N_18109,N_18604);
and U19408 (N_19408,N_18327,N_18941);
xnor U19409 (N_19409,N_18642,N_18613);
nor U19410 (N_19410,N_18110,N_18547);
nand U19411 (N_19411,N_18697,N_19095);
nor U19412 (N_19412,N_18903,N_19113);
or U19413 (N_19413,N_18153,N_18757);
nor U19414 (N_19414,N_18805,N_18489);
nand U19415 (N_19415,N_18713,N_18641);
and U19416 (N_19416,N_19059,N_18468);
nand U19417 (N_19417,N_18417,N_18630);
and U19418 (N_19418,N_18175,N_18305);
and U19419 (N_19419,N_18032,N_18887);
or U19420 (N_19420,N_18794,N_18411);
nor U19421 (N_19421,N_18620,N_18819);
nor U19422 (N_19422,N_18446,N_18066);
xor U19423 (N_19423,N_18524,N_18984);
and U19424 (N_19424,N_19176,N_18076);
nand U19425 (N_19425,N_18461,N_18542);
or U19426 (N_19426,N_18145,N_19173);
xnor U19427 (N_19427,N_18766,N_18293);
or U19428 (N_19428,N_18036,N_18440);
or U19429 (N_19429,N_18513,N_19018);
or U19430 (N_19430,N_18152,N_18553);
xnor U19431 (N_19431,N_18738,N_18502);
xnor U19432 (N_19432,N_18017,N_19077);
or U19433 (N_19433,N_19174,N_18516);
xor U19434 (N_19434,N_18050,N_18852);
xor U19435 (N_19435,N_18375,N_18117);
nand U19436 (N_19436,N_19020,N_18896);
and U19437 (N_19437,N_19008,N_19138);
nand U19438 (N_19438,N_18784,N_18111);
xnor U19439 (N_19439,N_18334,N_18464);
or U19440 (N_19440,N_18651,N_18965);
nand U19441 (N_19441,N_18025,N_18089);
or U19442 (N_19442,N_18129,N_19141);
nor U19443 (N_19443,N_18264,N_18379);
nand U19444 (N_19444,N_19177,N_18504);
and U19445 (N_19445,N_18748,N_19179);
and U19446 (N_19446,N_18837,N_19073);
nand U19447 (N_19447,N_19003,N_18559);
nand U19448 (N_19448,N_19066,N_19190);
nor U19449 (N_19449,N_18745,N_19026);
and U19450 (N_19450,N_18554,N_18023);
and U19451 (N_19451,N_18495,N_18419);
xor U19452 (N_19452,N_18561,N_18990);
and U19453 (N_19453,N_19155,N_18484);
or U19454 (N_19454,N_18458,N_18194);
and U19455 (N_19455,N_18922,N_18565);
nor U19456 (N_19456,N_18481,N_18430);
nor U19457 (N_19457,N_18747,N_19183);
or U19458 (N_19458,N_19162,N_18372);
or U19459 (N_19459,N_18636,N_18971);
nand U19460 (N_19460,N_18015,N_18914);
xor U19461 (N_19461,N_18768,N_19071);
nor U19462 (N_19462,N_18325,N_19104);
xnor U19463 (N_19463,N_18049,N_18765);
xnor U19464 (N_19464,N_18629,N_18640);
nand U19465 (N_19465,N_18633,N_19061);
nand U19466 (N_19466,N_18308,N_18818);
xnor U19467 (N_19467,N_18735,N_18685);
nor U19468 (N_19468,N_18549,N_18012);
and U19469 (N_19469,N_18253,N_18951);
xnor U19470 (N_19470,N_18370,N_18441);
and U19471 (N_19471,N_18063,N_18808);
nand U19472 (N_19472,N_18678,N_18876);
and U19473 (N_19473,N_18233,N_19171);
or U19474 (N_19474,N_19094,N_18900);
xor U19475 (N_19475,N_18677,N_19149);
or U19476 (N_19476,N_18125,N_18662);
or U19477 (N_19477,N_18625,N_18009);
xnor U19478 (N_19478,N_19074,N_18867);
or U19479 (N_19479,N_19070,N_18385);
or U19480 (N_19480,N_19139,N_18753);
or U19481 (N_19481,N_18605,N_18373);
xnor U19482 (N_19482,N_18278,N_19152);
xor U19483 (N_19483,N_18719,N_19047);
nor U19484 (N_19484,N_18744,N_18696);
xnor U19485 (N_19485,N_18466,N_18146);
or U19486 (N_19486,N_18822,N_18276);
or U19487 (N_19487,N_18245,N_18191);
or U19488 (N_19488,N_18909,N_18831);
xor U19489 (N_19489,N_18811,N_18450);
xnor U19490 (N_19490,N_18119,N_18568);
nand U19491 (N_19491,N_19191,N_18752);
nand U19492 (N_19492,N_18722,N_18790);
xor U19493 (N_19493,N_18249,N_18723);
nor U19494 (N_19494,N_18860,N_18762);
xnor U19495 (N_19495,N_19098,N_18211);
and U19496 (N_19496,N_18259,N_18258);
nand U19497 (N_19497,N_19056,N_18324);
xor U19498 (N_19498,N_18336,N_18352);
xor U19499 (N_19499,N_18813,N_18671);
nor U19500 (N_19500,N_18535,N_18767);
nand U19501 (N_19501,N_18829,N_18106);
nand U19502 (N_19502,N_18828,N_18800);
and U19503 (N_19503,N_18825,N_18473);
nor U19504 (N_19504,N_18045,N_18425);
xnor U19505 (N_19505,N_18157,N_18505);
xnor U19506 (N_19506,N_18349,N_18432);
xnor U19507 (N_19507,N_18611,N_18996);
and U19508 (N_19508,N_18209,N_18202);
xor U19509 (N_19509,N_18970,N_18600);
nand U19510 (N_19510,N_18179,N_18002);
xnor U19511 (N_19511,N_18608,N_18670);
nor U19512 (N_19512,N_18394,N_18585);
nor U19513 (N_19513,N_18200,N_19002);
or U19514 (N_19514,N_19081,N_18172);
xor U19515 (N_19515,N_19075,N_18874);
or U19516 (N_19516,N_18463,N_18161);
or U19517 (N_19517,N_18848,N_19064);
nor U19518 (N_19518,N_18363,N_18711);
xnor U19519 (N_19519,N_18389,N_18780);
nor U19520 (N_19520,N_18434,N_18734);
or U19521 (N_19521,N_18329,N_18533);
xnor U19522 (N_19522,N_19166,N_18456);
or U19523 (N_19523,N_18736,N_18701);
xnor U19524 (N_19524,N_19157,N_18695);
or U19525 (N_19525,N_19127,N_18750);
nor U19526 (N_19526,N_18053,N_18123);
nand U19527 (N_19527,N_19180,N_18080);
xor U19528 (N_19528,N_19060,N_18575);
xnor U19529 (N_19529,N_18291,N_19007);
and U19530 (N_19530,N_18615,N_18555);
xnor U19531 (N_19531,N_19128,N_18981);
nor U19532 (N_19532,N_18980,N_18587);
xnor U19533 (N_19533,N_18905,N_18802);
and U19534 (N_19534,N_18199,N_18256);
or U19535 (N_19535,N_18122,N_18948);
nor U19536 (N_19536,N_18407,N_18664);
nor U19537 (N_19537,N_18859,N_18560);
or U19538 (N_19538,N_18184,N_18496);
nor U19539 (N_19539,N_18917,N_18052);
or U19540 (N_19540,N_19111,N_18027);
nor U19541 (N_19541,N_19193,N_18294);
nor U19542 (N_19542,N_18597,N_18871);
nor U19543 (N_19543,N_18862,N_19117);
or U19544 (N_19544,N_18653,N_18416);
nand U19545 (N_19545,N_18491,N_19172);
nand U19546 (N_19546,N_18388,N_18567);
nand U19547 (N_19547,N_18873,N_19037);
xnor U19548 (N_19548,N_18679,N_18506);
nand U19549 (N_19549,N_18307,N_18816);
xor U19550 (N_19550,N_18177,N_18290);
or U19551 (N_19551,N_18228,N_18107);
nor U19552 (N_19552,N_18422,N_18207);
nand U19553 (N_19553,N_18223,N_19196);
nand U19554 (N_19554,N_18160,N_19131);
or U19555 (N_19555,N_18310,N_18262);
nand U19556 (N_19556,N_18964,N_18400);
nand U19557 (N_19557,N_18445,N_18055);
and U19558 (N_19558,N_18680,N_18497);
nand U19559 (N_19559,N_18634,N_18566);
nor U19560 (N_19560,N_18387,N_18786);
and U19561 (N_19561,N_18728,N_18236);
xor U19562 (N_19562,N_18118,N_18989);
and U19563 (N_19563,N_18772,N_18306);
xor U19564 (N_19564,N_18839,N_18779);
and U19565 (N_19565,N_18708,N_18393);
and U19566 (N_19566,N_18284,N_19160);
xor U19567 (N_19567,N_18183,N_18564);
nand U19568 (N_19568,N_18756,N_18782);
and U19569 (N_19569,N_18083,N_18482);
nor U19570 (N_19570,N_18849,N_18331);
nand U19571 (N_19571,N_18556,N_19046);
and U19572 (N_19572,N_18467,N_18514);
nand U19573 (N_19573,N_18418,N_19013);
and U19574 (N_19574,N_18727,N_19080);
xor U19575 (N_19575,N_18995,N_18316);
or U19576 (N_19576,N_19024,N_18134);
nor U19577 (N_19577,N_18872,N_18383);
xnor U19578 (N_19578,N_18637,N_18185);
and U19579 (N_19579,N_18424,N_19096);
nor U19580 (N_19580,N_19043,N_19031);
nand U19581 (N_19581,N_18366,N_18730);
nand U19582 (N_19582,N_18196,N_18135);
and U19583 (N_19583,N_18627,N_18426);
and U19584 (N_19584,N_18824,N_18035);
and U19585 (N_19585,N_18583,N_18699);
nor U19586 (N_19586,N_18190,N_18429);
and U19587 (N_19587,N_18739,N_18404);
xnor U19588 (N_19588,N_18248,N_18455);
or U19589 (N_19589,N_18674,N_18198);
nand U19590 (N_19590,N_18084,N_18924);
xnor U19591 (N_19591,N_18520,N_18531);
or U19592 (N_19592,N_18881,N_18494);
nand U19593 (N_19593,N_18380,N_18741);
nand U19594 (N_19594,N_18962,N_18355);
xor U19595 (N_19595,N_19145,N_18650);
nor U19596 (N_19596,N_18519,N_18539);
or U19597 (N_19597,N_18709,N_18465);
nor U19598 (N_19598,N_19134,N_18777);
nor U19599 (N_19599,N_18345,N_18979);
xor U19600 (N_19600,N_18706,N_18999);
nand U19601 (N_19601,N_19099,N_18057);
nand U19602 (N_19602,N_18268,N_18665);
nand U19603 (N_19603,N_19123,N_18894);
xnor U19604 (N_19604,N_18390,N_18353);
or U19605 (N_19605,N_18131,N_18319);
xnor U19606 (N_19606,N_18619,N_18858);
or U19607 (N_19607,N_19161,N_18140);
or U19608 (N_19608,N_18740,N_18040);
and U19609 (N_19609,N_18092,N_18102);
xnor U19610 (N_19610,N_19078,N_18280);
and U19611 (N_19611,N_18622,N_18788);
or U19612 (N_19612,N_18480,N_19137);
or U19613 (N_19613,N_18167,N_18339);
nand U19614 (N_19614,N_19093,N_18395);
nor U19615 (N_19615,N_18987,N_18241);
nor U19616 (N_19616,N_19181,N_18530);
or U19617 (N_19617,N_18475,N_18618);
xor U19618 (N_19618,N_18333,N_18408);
nand U19619 (N_19619,N_18743,N_19163);
nand U19620 (N_19620,N_18643,N_18037);
xnor U19621 (N_19621,N_18732,N_18590);
and U19622 (N_19622,N_18998,N_19085);
xor U19623 (N_19623,N_18077,N_18923);
nand U19624 (N_19624,N_18132,N_18523);
nand U19625 (N_19625,N_18303,N_18843);
nand U19626 (N_19626,N_18197,N_19079);
nor U19627 (N_19627,N_18724,N_18263);
and U19628 (N_19628,N_18156,N_18270);
nand U19629 (N_19629,N_18898,N_18835);
nand U19630 (N_19630,N_18834,N_18471);
nor U19631 (N_19631,N_18415,N_18326);
nor U19632 (N_19632,N_18016,N_18906);
xor U19633 (N_19633,N_18269,N_18993);
nand U19634 (N_19634,N_18694,N_19044);
and U19635 (N_19635,N_18591,N_18603);
nor U19636 (N_19636,N_18676,N_18033);
or U19637 (N_19637,N_18911,N_18953);
nor U19638 (N_19638,N_18321,N_18503);
nand U19639 (N_19639,N_18216,N_18595);
or U19640 (N_19640,N_18601,N_18103);
nor U19641 (N_19641,N_18116,N_18150);
nand U19642 (N_19642,N_18120,N_18340);
nor U19643 (N_19643,N_18693,N_18763);
nand U19644 (N_19644,N_18100,N_18213);
nand U19645 (N_19645,N_18281,N_18958);
nand U19646 (N_19646,N_18507,N_18392);
nand U19647 (N_19647,N_18105,N_18493);
nand U19648 (N_19648,N_18358,N_18588);
and U19649 (N_19649,N_18067,N_18541);
xnor U19650 (N_19650,N_18518,N_18486);
nand U19651 (N_19651,N_18279,N_18201);
and U19652 (N_19652,N_18796,N_18243);
and U19653 (N_19653,N_18008,N_18313);
nand U19654 (N_19654,N_18098,N_18624);
xor U19655 (N_19655,N_19105,N_19014);
nand U19656 (N_19656,N_18483,N_18309);
xor U19657 (N_19657,N_18378,N_19199);
and U19658 (N_19658,N_18684,N_18919);
nand U19659 (N_19659,N_18232,N_18720);
xnor U19660 (N_19660,N_18292,N_19109);
and U19661 (N_19661,N_18457,N_18529);
nand U19662 (N_19662,N_18657,N_19016);
nand U19663 (N_19663,N_18341,N_18367);
nor U19664 (N_19664,N_18058,N_18271);
and U19665 (N_19665,N_18272,N_18143);
and U19666 (N_19666,N_18761,N_18942);
or U19667 (N_19667,N_18814,N_18545);
or U19668 (N_19668,N_18218,N_18059);
and U19669 (N_19669,N_19124,N_18842);
nor U19670 (N_19670,N_18913,N_19050);
and U19671 (N_19671,N_18104,N_18907);
and U19672 (N_19672,N_18230,N_18563);
or U19673 (N_19673,N_18296,N_18247);
nand U19674 (N_19674,N_18638,N_18320);
nand U19675 (N_19675,N_18346,N_18801);
nor U19676 (N_19676,N_19033,N_18368);
nand U19677 (N_19677,N_18490,N_19186);
and U19678 (N_19678,N_18396,N_18238);
and U19679 (N_19679,N_18492,N_19072);
nand U19680 (N_19680,N_18220,N_19182);
and U19681 (N_19681,N_18322,N_18528);
nand U19682 (N_19682,N_18428,N_18479);
nor U19683 (N_19683,N_18870,N_18168);
nor U19684 (N_19684,N_18038,N_18021);
nand U19685 (N_19685,N_18826,N_18820);
and U19686 (N_19686,N_18242,N_18311);
nand U19687 (N_19687,N_18409,N_19169);
nor U19688 (N_19688,N_19021,N_18660);
nand U19689 (N_19689,N_18169,N_18384);
nor U19690 (N_19690,N_18154,N_18192);
xor U19691 (N_19691,N_18586,N_18068);
xor U19692 (N_19692,N_18598,N_18658);
nor U19693 (N_19693,N_18136,N_18204);
nor U19694 (N_19694,N_19022,N_19012);
or U19695 (N_19695,N_18785,N_18022);
nor U19696 (N_19696,N_18616,N_18755);
nand U19697 (N_19697,N_18011,N_18886);
and U19698 (N_19698,N_18285,N_19192);
nand U19699 (N_19699,N_18628,N_18427);
nor U19700 (N_19700,N_19069,N_18582);
nand U19701 (N_19701,N_18891,N_18360);
or U19702 (N_19702,N_18830,N_18632);
or U19703 (N_19703,N_18189,N_18070);
or U19704 (N_19704,N_18056,N_18882);
xnor U19705 (N_19705,N_18932,N_18851);
nand U19706 (N_19706,N_18672,N_18985);
nor U19707 (N_19707,N_19164,N_18982);
or U19708 (N_19708,N_18234,N_18275);
nand U19709 (N_19709,N_19052,N_18746);
xnor U19710 (N_19710,N_18593,N_19049);
and U19711 (N_19711,N_19025,N_18833);
nor U19712 (N_19712,N_19195,N_19130);
or U19713 (N_19713,N_19146,N_18437);
nand U19714 (N_19714,N_18827,N_18206);
or U19715 (N_19715,N_18019,N_18817);
xor U19716 (N_19716,N_19144,N_18030);
and U19717 (N_19717,N_19188,N_18171);
and U19718 (N_19718,N_18508,N_19165);
nand U19719 (N_19719,N_18435,N_19118);
nor U19720 (N_19720,N_18460,N_18927);
nand U19721 (N_19721,N_18005,N_18614);
nand U19722 (N_19722,N_18698,N_19053);
or U19723 (N_19723,N_18108,N_18344);
nand U19724 (N_19724,N_18127,N_19005);
nand U19725 (N_19725,N_18439,N_19140);
nand U19726 (N_19726,N_18936,N_18930);
nand U19727 (N_19727,N_18082,N_18921);
nand U19728 (N_19728,N_18594,N_18421);
nand U19729 (N_19729,N_18090,N_18733);
nor U19730 (N_19730,N_18853,N_18029);
and U19731 (N_19731,N_18607,N_18935);
and U19732 (N_19732,N_19028,N_18776);
xnor U19733 (N_19733,N_18691,N_18710);
nor U19734 (N_19734,N_18031,N_18908);
and U19735 (N_19735,N_19042,N_19058);
nand U19736 (N_19736,N_18967,N_18142);
xor U19737 (N_19737,N_18088,N_18656);
and U19738 (N_19738,N_18359,N_18155);
nand U19739 (N_19739,N_18537,N_18039);
nand U19740 (N_19740,N_18163,N_18929);
or U19741 (N_19741,N_19027,N_18861);
or U19742 (N_19742,N_18374,N_18124);
xnor U19743 (N_19743,N_18511,N_18623);
nor U19744 (N_19744,N_18069,N_18557);
nor U19745 (N_19745,N_18459,N_18510);
nand U19746 (N_19746,N_18712,N_18423);
nor U19747 (N_19747,N_19062,N_19156);
nor U19748 (N_19748,N_18260,N_19034);
or U19749 (N_19749,N_18617,N_19090);
nand U19750 (N_19750,N_18821,N_18659);
or U19751 (N_19751,N_18028,N_19133);
or U19752 (N_19752,N_18937,N_19017);
or U19753 (N_19753,N_19132,N_18337);
nor U19754 (N_19754,N_18716,N_18646);
or U19755 (N_19755,N_18376,N_18010);
xnor U19756 (N_19756,N_18182,N_18543);
xor U19757 (N_19757,N_18621,N_18044);
or U19758 (N_19758,N_18113,N_18412);
or U19759 (N_19759,N_18115,N_18573);
or U19760 (N_19760,N_19143,N_18815);
and U19761 (N_19761,N_19083,N_19040);
and U19762 (N_19762,N_18342,N_18277);
or U19763 (N_19763,N_18176,N_18297);
nor U19764 (N_19764,N_18126,N_18726);
nor U19765 (N_19765,N_18267,N_18180);
nand U19766 (N_19766,N_18527,N_19045);
and U19767 (N_19767,N_18809,N_18164);
or U19768 (N_19768,N_18065,N_18551);
xnor U19769 (N_19769,N_18760,N_19089);
nor U19770 (N_19770,N_18654,N_18692);
nand U19771 (N_19771,N_18174,N_18550);
nand U19772 (N_19772,N_18431,N_18512);
nor U19773 (N_19773,N_18683,N_18836);
nand U19774 (N_19774,N_19108,N_18086);
and U19775 (N_19775,N_18546,N_18401);
nor U19776 (N_19776,N_18957,N_18087);
and U19777 (N_19777,N_18885,N_18114);
nor U19778 (N_19778,N_18462,N_18977);
nor U19779 (N_19779,N_19197,N_18438);
and U19780 (N_19780,N_18006,N_18402);
or U19781 (N_19781,N_19185,N_18061);
or U19782 (N_19782,N_18397,N_18702);
and U19783 (N_19783,N_19147,N_18578);
or U19784 (N_19784,N_18521,N_18526);
xor U19785 (N_19785,N_18302,N_18994);
nand U19786 (N_19786,N_18093,N_18444);
nor U19787 (N_19787,N_18170,N_18682);
and U19788 (N_19788,N_18091,N_18351);
nand U19789 (N_19789,N_18856,N_18754);
or U19790 (N_19790,N_18969,N_19122);
nand U19791 (N_19791,N_18577,N_18968);
or U19792 (N_19792,N_19151,N_18295);
nand U19793 (N_19793,N_18244,N_18890);
nand U19794 (N_19794,N_18014,N_18227);
nand U19795 (N_19795,N_18485,N_18991);
nand U19796 (N_19796,N_18381,N_18988);
nor U19797 (N_19797,N_18920,N_18517);
nand U19798 (N_19798,N_18798,N_18470);
or U19799 (N_19799,N_18854,N_19102);
nor U19800 (N_19800,N_19149,N_19043);
or U19801 (N_19801,N_18580,N_18163);
and U19802 (N_19802,N_19152,N_18251);
nand U19803 (N_19803,N_18119,N_18790);
nor U19804 (N_19804,N_18833,N_19033);
xor U19805 (N_19805,N_18022,N_18657);
nor U19806 (N_19806,N_19064,N_18475);
nand U19807 (N_19807,N_18709,N_18360);
and U19808 (N_19808,N_19015,N_18626);
xor U19809 (N_19809,N_19199,N_18264);
or U19810 (N_19810,N_18108,N_19028);
nor U19811 (N_19811,N_18807,N_18100);
or U19812 (N_19812,N_18452,N_18661);
xnor U19813 (N_19813,N_18570,N_18993);
xor U19814 (N_19814,N_18896,N_18976);
nand U19815 (N_19815,N_18656,N_18403);
or U19816 (N_19816,N_18117,N_19090);
xnor U19817 (N_19817,N_18810,N_18970);
or U19818 (N_19818,N_19128,N_19006);
nor U19819 (N_19819,N_19156,N_18193);
nor U19820 (N_19820,N_19086,N_18753);
nor U19821 (N_19821,N_18423,N_18594);
xnor U19822 (N_19822,N_18204,N_18051);
or U19823 (N_19823,N_18804,N_19030);
or U19824 (N_19824,N_18385,N_18432);
nor U19825 (N_19825,N_18119,N_18285);
xor U19826 (N_19826,N_18028,N_18574);
xor U19827 (N_19827,N_18328,N_18921);
xnor U19828 (N_19828,N_18985,N_18211);
xor U19829 (N_19829,N_19167,N_19053);
or U19830 (N_19830,N_18215,N_18838);
nor U19831 (N_19831,N_18651,N_18323);
nand U19832 (N_19832,N_18064,N_18174);
and U19833 (N_19833,N_18474,N_19050);
nor U19834 (N_19834,N_18241,N_18202);
xor U19835 (N_19835,N_19188,N_18337);
or U19836 (N_19836,N_18607,N_18732);
xnor U19837 (N_19837,N_18595,N_18787);
nand U19838 (N_19838,N_19183,N_18548);
xor U19839 (N_19839,N_18112,N_19152);
xnor U19840 (N_19840,N_18096,N_18830);
nor U19841 (N_19841,N_18677,N_19063);
and U19842 (N_19842,N_18208,N_18961);
nand U19843 (N_19843,N_18380,N_18381);
or U19844 (N_19844,N_18633,N_18264);
xor U19845 (N_19845,N_19035,N_18456);
and U19846 (N_19846,N_18362,N_19013);
xor U19847 (N_19847,N_18976,N_18137);
xnor U19848 (N_19848,N_18253,N_18168);
nor U19849 (N_19849,N_18283,N_18836);
and U19850 (N_19850,N_18937,N_18581);
or U19851 (N_19851,N_19185,N_18593);
nor U19852 (N_19852,N_19112,N_18236);
and U19853 (N_19853,N_18250,N_18112);
xor U19854 (N_19854,N_18946,N_18599);
or U19855 (N_19855,N_18464,N_18226);
or U19856 (N_19856,N_18248,N_18800);
xnor U19857 (N_19857,N_18450,N_18555);
and U19858 (N_19858,N_18125,N_18362);
nor U19859 (N_19859,N_19191,N_18188);
or U19860 (N_19860,N_18627,N_18301);
and U19861 (N_19861,N_19002,N_18931);
nand U19862 (N_19862,N_18982,N_18652);
xnor U19863 (N_19863,N_18353,N_19173);
or U19864 (N_19864,N_18686,N_18106);
xor U19865 (N_19865,N_18015,N_18176);
nor U19866 (N_19866,N_18048,N_18904);
nand U19867 (N_19867,N_18722,N_18299);
and U19868 (N_19868,N_19128,N_18537);
nor U19869 (N_19869,N_18384,N_18088);
nand U19870 (N_19870,N_18456,N_18541);
nor U19871 (N_19871,N_18736,N_18392);
nand U19872 (N_19872,N_18461,N_18162);
or U19873 (N_19873,N_18856,N_18326);
xnor U19874 (N_19874,N_18815,N_19052);
nand U19875 (N_19875,N_18922,N_18046);
nor U19876 (N_19876,N_18168,N_18163);
nand U19877 (N_19877,N_18138,N_18127);
xor U19878 (N_19878,N_18758,N_18907);
nor U19879 (N_19879,N_19077,N_18490);
nor U19880 (N_19880,N_18405,N_18167);
xnor U19881 (N_19881,N_18667,N_19171);
or U19882 (N_19882,N_18318,N_18468);
or U19883 (N_19883,N_18239,N_18179);
nand U19884 (N_19884,N_18979,N_18970);
and U19885 (N_19885,N_18575,N_18274);
nand U19886 (N_19886,N_18928,N_18289);
or U19887 (N_19887,N_18278,N_18582);
nand U19888 (N_19888,N_18718,N_18501);
xor U19889 (N_19889,N_19001,N_18084);
nand U19890 (N_19890,N_18053,N_18058);
and U19891 (N_19891,N_18535,N_18990);
xnor U19892 (N_19892,N_18051,N_18758);
and U19893 (N_19893,N_18625,N_18879);
nand U19894 (N_19894,N_18776,N_18630);
and U19895 (N_19895,N_18465,N_19058);
nor U19896 (N_19896,N_18891,N_19117);
xnor U19897 (N_19897,N_18290,N_18268);
nor U19898 (N_19898,N_18331,N_18461);
or U19899 (N_19899,N_18797,N_18714);
nor U19900 (N_19900,N_18107,N_18689);
or U19901 (N_19901,N_18044,N_18451);
nor U19902 (N_19902,N_18014,N_18466);
nor U19903 (N_19903,N_19145,N_18561);
or U19904 (N_19904,N_18196,N_18160);
xnor U19905 (N_19905,N_18386,N_18291);
xnor U19906 (N_19906,N_18263,N_18876);
or U19907 (N_19907,N_18237,N_18907);
and U19908 (N_19908,N_18577,N_18439);
nand U19909 (N_19909,N_18287,N_18760);
nor U19910 (N_19910,N_18773,N_18052);
or U19911 (N_19911,N_18889,N_19192);
nor U19912 (N_19912,N_18462,N_18567);
and U19913 (N_19913,N_18815,N_18637);
nand U19914 (N_19914,N_19046,N_18280);
xnor U19915 (N_19915,N_18317,N_19012);
and U19916 (N_19916,N_18304,N_19176);
xor U19917 (N_19917,N_18032,N_19026);
nand U19918 (N_19918,N_18954,N_18567);
nor U19919 (N_19919,N_19171,N_18837);
nor U19920 (N_19920,N_18715,N_18852);
xnor U19921 (N_19921,N_18837,N_18748);
nand U19922 (N_19922,N_19113,N_18115);
xor U19923 (N_19923,N_19123,N_18502);
xnor U19924 (N_19924,N_18972,N_18054);
xor U19925 (N_19925,N_18957,N_18955);
nand U19926 (N_19926,N_18231,N_18253);
and U19927 (N_19927,N_18132,N_18325);
nor U19928 (N_19928,N_18129,N_18864);
nand U19929 (N_19929,N_18351,N_18757);
xnor U19930 (N_19930,N_18106,N_19055);
nor U19931 (N_19931,N_18824,N_18490);
nand U19932 (N_19932,N_18524,N_18593);
xor U19933 (N_19933,N_18949,N_18919);
nand U19934 (N_19934,N_18911,N_18620);
or U19935 (N_19935,N_19184,N_18560);
nor U19936 (N_19936,N_19039,N_18245);
nor U19937 (N_19937,N_18149,N_18645);
xnor U19938 (N_19938,N_18485,N_18844);
nand U19939 (N_19939,N_18536,N_18291);
nor U19940 (N_19940,N_18061,N_18817);
xor U19941 (N_19941,N_18539,N_18058);
nor U19942 (N_19942,N_18629,N_19108);
or U19943 (N_19943,N_18896,N_19026);
or U19944 (N_19944,N_18302,N_19119);
or U19945 (N_19945,N_18499,N_18285);
or U19946 (N_19946,N_18278,N_18206);
nor U19947 (N_19947,N_18327,N_18317);
or U19948 (N_19948,N_18957,N_19005);
nand U19949 (N_19949,N_18673,N_18800);
or U19950 (N_19950,N_18466,N_18255);
and U19951 (N_19951,N_19161,N_18499);
and U19952 (N_19952,N_19027,N_18685);
nand U19953 (N_19953,N_19184,N_18051);
and U19954 (N_19954,N_18316,N_19116);
xnor U19955 (N_19955,N_18751,N_18122);
and U19956 (N_19956,N_18418,N_18150);
and U19957 (N_19957,N_18680,N_18920);
nand U19958 (N_19958,N_18048,N_19042);
and U19959 (N_19959,N_18660,N_18200);
and U19960 (N_19960,N_18202,N_18013);
xor U19961 (N_19961,N_18444,N_18472);
and U19962 (N_19962,N_18463,N_18310);
or U19963 (N_19963,N_19057,N_18645);
nand U19964 (N_19964,N_18428,N_19005);
nand U19965 (N_19965,N_19153,N_18888);
nand U19966 (N_19966,N_18120,N_18164);
or U19967 (N_19967,N_18512,N_18300);
nand U19968 (N_19968,N_18692,N_18182);
nor U19969 (N_19969,N_19161,N_18929);
or U19970 (N_19970,N_19124,N_18373);
nand U19971 (N_19971,N_19185,N_18669);
or U19972 (N_19972,N_18537,N_19012);
nand U19973 (N_19973,N_18855,N_18465);
and U19974 (N_19974,N_19026,N_18031);
nand U19975 (N_19975,N_18156,N_18727);
or U19976 (N_19976,N_18809,N_18952);
or U19977 (N_19977,N_18455,N_18665);
or U19978 (N_19978,N_18667,N_18635);
nor U19979 (N_19979,N_19028,N_18782);
nor U19980 (N_19980,N_18167,N_18745);
xor U19981 (N_19981,N_18400,N_18916);
nand U19982 (N_19982,N_19088,N_18283);
xnor U19983 (N_19983,N_18842,N_18341);
and U19984 (N_19984,N_19087,N_18990);
or U19985 (N_19985,N_18079,N_18810);
xnor U19986 (N_19986,N_18530,N_18441);
and U19987 (N_19987,N_18975,N_18611);
xnor U19988 (N_19988,N_18813,N_18929);
nor U19989 (N_19989,N_18710,N_18495);
or U19990 (N_19990,N_19161,N_18115);
and U19991 (N_19991,N_18671,N_18949);
xnor U19992 (N_19992,N_18926,N_18621);
nand U19993 (N_19993,N_18349,N_19080);
nand U19994 (N_19994,N_19045,N_18070);
nand U19995 (N_19995,N_18122,N_18555);
and U19996 (N_19996,N_18546,N_18025);
or U19997 (N_19997,N_18266,N_18061);
or U19998 (N_19998,N_18360,N_18087);
nor U19999 (N_19999,N_19117,N_18123);
nor U20000 (N_20000,N_19092,N_18507);
nor U20001 (N_20001,N_19169,N_18024);
nor U20002 (N_20002,N_18269,N_19026);
nand U20003 (N_20003,N_18838,N_18719);
xor U20004 (N_20004,N_18394,N_18548);
and U20005 (N_20005,N_18824,N_18641);
and U20006 (N_20006,N_18363,N_18787);
nand U20007 (N_20007,N_19000,N_18303);
nor U20008 (N_20008,N_18836,N_18793);
xor U20009 (N_20009,N_18297,N_19005);
nor U20010 (N_20010,N_19138,N_19074);
nor U20011 (N_20011,N_18261,N_19196);
xor U20012 (N_20012,N_18615,N_18685);
and U20013 (N_20013,N_18350,N_18745);
and U20014 (N_20014,N_18306,N_18535);
and U20015 (N_20015,N_18634,N_18879);
xor U20016 (N_20016,N_18976,N_18827);
nor U20017 (N_20017,N_18874,N_18201);
nor U20018 (N_20018,N_18266,N_18519);
nor U20019 (N_20019,N_18158,N_19145);
and U20020 (N_20020,N_18762,N_18637);
and U20021 (N_20021,N_19027,N_18908);
xnor U20022 (N_20022,N_18832,N_18153);
nor U20023 (N_20023,N_18727,N_18075);
nor U20024 (N_20024,N_18939,N_18840);
nand U20025 (N_20025,N_18749,N_18289);
or U20026 (N_20026,N_18214,N_18838);
nor U20027 (N_20027,N_18695,N_18683);
xor U20028 (N_20028,N_18270,N_19160);
nand U20029 (N_20029,N_18000,N_18488);
xor U20030 (N_20030,N_18520,N_18601);
nor U20031 (N_20031,N_18237,N_19119);
nor U20032 (N_20032,N_18158,N_18137);
nor U20033 (N_20033,N_18866,N_18697);
xnor U20034 (N_20034,N_18066,N_18906);
xnor U20035 (N_20035,N_19072,N_18679);
xor U20036 (N_20036,N_18202,N_18317);
xnor U20037 (N_20037,N_18110,N_19077);
xor U20038 (N_20038,N_18478,N_18920);
nand U20039 (N_20039,N_19021,N_18395);
nand U20040 (N_20040,N_18995,N_19142);
nand U20041 (N_20041,N_18738,N_18466);
nor U20042 (N_20042,N_18715,N_18988);
and U20043 (N_20043,N_18033,N_18517);
and U20044 (N_20044,N_18316,N_18836);
or U20045 (N_20045,N_18177,N_19066);
and U20046 (N_20046,N_18319,N_18649);
nand U20047 (N_20047,N_18054,N_18418);
nand U20048 (N_20048,N_18665,N_18343);
nor U20049 (N_20049,N_18610,N_18780);
xor U20050 (N_20050,N_18291,N_18257);
or U20051 (N_20051,N_18039,N_18091);
xnor U20052 (N_20052,N_18115,N_18430);
xnor U20053 (N_20053,N_18659,N_18478);
and U20054 (N_20054,N_18659,N_18164);
or U20055 (N_20055,N_18749,N_19040);
and U20056 (N_20056,N_18907,N_18620);
and U20057 (N_20057,N_18795,N_18129);
xor U20058 (N_20058,N_19070,N_19111);
xor U20059 (N_20059,N_18163,N_18750);
or U20060 (N_20060,N_18501,N_18936);
or U20061 (N_20061,N_18454,N_18725);
and U20062 (N_20062,N_18796,N_18778);
or U20063 (N_20063,N_18656,N_18438);
nand U20064 (N_20064,N_18961,N_18085);
xnor U20065 (N_20065,N_18251,N_19121);
or U20066 (N_20066,N_18071,N_18945);
xor U20067 (N_20067,N_18455,N_18033);
or U20068 (N_20068,N_19199,N_18891);
nand U20069 (N_20069,N_19006,N_18651);
or U20070 (N_20070,N_18749,N_19191);
nand U20071 (N_20071,N_18239,N_18676);
and U20072 (N_20072,N_19003,N_18977);
or U20073 (N_20073,N_18676,N_18999);
xor U20074 (N_20074,N_18415,N_18967);
xnor U20075 (N_20075,N_18988,N_18548);
nor U20076 (N_20076,N_19012,N_18256);
and U20077 (N_20077,N_18172,N_18612);
and U20078 (N_20078,N_18752,N_18000);
or U20079 (N_20079,N_18728,N_18312);
xor U20080 (N_20080,N_18326,N_18031);
and U20081 (N_20081,N_18043,N_18432);
nand U20082 (N_20082,N_18352,N_18786);
and U20083 (N_20083,N_19107,N_18548);
and U20084 (N_20084,N_18239,N_18746);
nor U20085 (N_20085,N_18947,N_18559);
nor U20086 (N_20086,N_18308,N_18260);
and U20087 (N_20087,N_18824,N_18415);
nand U20088 (N_20088,N_19012,N_19017);
nand U20089 (N_20089,N_18113,N_18629);
nand U20090 (N_20090,N_18376,N_18678);
and U20091 (N_20091,N_18885,N_18328);
and U20092 (N_20092,N_19119,N_18661);
nor U20093 (N_20093,N_18734,N_19148);
nand U20094 (N_20094,N_19062,N_18866);
xor U20095 (N_20095,N_19150,N_18557);
nor U20096 (N_20096,N_18343,N_18957);
nor U20097 (N_20097,N_18830,N_19007);
nor U20098 (N_20098,N_18672,N_18961);
and U20099 (N_20099,N_18632,N_18881);
nor U20100 (N_20100,N_18357,N_19186);
and U20101 (N_20101,N_18360,N_19022);
and U20102 (N_20102,N_18080,N_18138);
or U20103 (N_20103,N_18548,N_18985);
or U20104 (N_20104,N_18073,N_18700);
and U20105 (N_20105,N_18473,N_18084);
and U20106 (N_20106,N_18308,N_18448);
nand U20107 (N_20107,N_18655,N_18712);
and U20108 (N_20108,N_18646,N_19145);
xnor U20109 (N_20109,N_18119,N_18602);
xor U20110 (N_20110,N_18760,N_19194);
or U20111 (N_20111,N_18125,N_19162);
xor U20112 (N_20112,N_19170,N_18796);
nand U20113 (N_20113,N_18689,N_18936);
or U20114 (N_20114,N_18643,N_18551);
or U20115 (N_20115,N_18044,N_18866);
xnor U20116 (N_20116,N_18338,N_18325);
xnor U20117 (N_20117,N_18453,N_18869);
xnor U20118 (N_20118,N_18843,N_18079);
nand U20119 (N_20119,N_18785,N_18163);
xor U20120 (N_20120,N_19118,N_19053);
nand U20121 (N_20121,N_18488,N_18930);
xnor U20122 (N_20122,N_18002,N_18847);
or U20123 (N_20123,N_18895,N_18976);
nor U20124 (N_20124,N_18720,N_18224);
nand U20125 (N_20125,N_19149,N_18003);
nand U20126 (N_20126,N_18971,N_18233);
or U20127 (N_20127,N_18022,N_18165);
nand U20128 (N_20128,N_18053,N_18403);
nor U20129 (N_20129,N_18344,N_18836);
xnor U20130 (N_20130,N_18499,N_18787);
or U20131 (N_20131,N_18579,N_18712);
xor U20132 (N_20132,N_18160,N_19022);
nand U20133 (N_20133,N_18571,N_19093);
nand U20134 (N_20134,N_18761,N_18462);
xor U20135 (N_20135,N_18834,N_18181);
nand U20136 (N_20136,N_18150,N_18903);
or U20137 (N_20137,N_19172,N_18164);
nand U20138 (N_20138,N_18501,N_18001);
xnor U20139 (N_20139,N_18423,N_18593);
nand U20140 (N_20140,N_18230,N_18163);
nor U20141 (N_20141,N_18236,N_18427);
nand U20142 (N_20142,N_18407,N_18539);
or U20143 (N_20143,N_18686,N_19132);
or U20144 (N_20144,N_18913,N_18403);
and U20145 (N_20145,N_18391,N_18310);
or U20146 (N_20146,N_19082,N_18005);
nand U20147 (N_20147,N_19005,N_18615);
xnor U20148 (N_20148,N_18740,N_18923);
nand U20149 (N_20149,N_18629,N_18420);
nand U20150 (N_20150,N_18539,N_18203);
and U20151 (N_20151,N_18453,N_18124);
nor U20152 (N_20152,N_18714,N_18084);
nand U20153 (N_20153,N_18623,N_19095);
nor U20154 (N_20154,N_18007,N_18029);
and U20155 (N_20155,N_19133,N_18673);
xnor U20156 (N_20156,N_19051,N_18998);
or U20157 (N_20157,N_18886,N_18171);
or U20158 (N_20158,N_18398,N_18866);
nor U20159 (N_20159,N_18518,N_18403);
or U20160 (N_20160,N_19063,N_18355);
nand U20161 (N_20161,N_18779,N_18861);
nand U20162 (N_20162,N_18162,N_18602);
and U20163 (N_20163,N_18258,N_18060);
nand U20164 (N_20164,N_19095,N_18478);
nor U20165 (N_20165,N_18911,N_18293);
nor U20166 (N_20166,N_18723,N_19152);
nand U20167 (N_20167,N_19119,N_18499);
nor U20168 (N_20168,N_18272,N_18114);
nand U20169 (N_20169,N_18864,N_18461);
or U20170 (N_20170,N_18212,N_18542);
and U20171 (N_20171,N_18330,N_18236);
and U20172 (N_20172,N_18109,N_18886);
nor U20173 (N_20173,N_18868,N_18569);
nand U20174 (N_20174,N_18462,N_18966);
nand U20175 (N_20175,N_18447,N_18219);
or U20176 (N_20176,N_18364,N_18738);
xnor U20177 (N_20177,N_18620,N_18918);
or U20178 (N_20178,N_18293,N_18916);
nor U20179 (N_20179,N_18253,N_18591);
xor U20180 (N_20180,N_18568,N_18941);
or U20181 (N_20181,N_18797,N_18099);
or U20182 (N_20182,N_18386,N_18409);
nor U20183 (N_20183,N_18829,N_18910);
nand U20184 (N_20184,N_19027,N_18204);
and U20185 (N_20185,N_18838,N_18529);
or U20186 (N_20186,N_19098,N_18753);
xor U20187 (N_20187,N_19189,N_18332);
nand U20188 (N_20188,N_18689,N_19014);
nand U20189 (N_20189,N_18418,N_18682);
nand U20190 (N_20190,N_18801,N_19162);
and U20191 (N_20191,N_19064,N_19065);
nor U20192 (N_20192,N_19056,N_18768);
nor U20193 (N_20193,N_18985,N_19016);
and U20194 (N_20194,N_18252,N_19195);
xnor U20195 (N_20195,N_19136,N_18667);
and U20196 (N_20196,N_18331,N_18942);
nor U20197 (N_20197,N_18674,N_19055);
nand U20198 (N_20198,N_18465,N_18034);
xnor U20199 (N_20199,N_19007,N_18519);
nor U20200 (N_20200,N_18614,N_19167);
nand U20201 (N_20201,N_18807,N_18170);
and U20202 (N_20202,N_18532,N_18643);
and U20203 (N_20203,N_18660,N_19151);
xnor U20204 (N_20204,N_18496,N_18322);
nor U20205 (N_20205,N_18756,N_18814);
xor U20206 (N_20206,N_18561,N_18331);
or U20207 (N_20207,N_18559,N_18785);
nand U20208 (N_20208,N_19011,N_18430);
nand U20209 (N_20209,N_18628,N_18697);
xnor U20210 (N_20210,N_19039,N_18352);
nand U20211 (N_20211,N_19182,N_18645);
and U20212 (N_20212,N_19069,N_18260);
and U20213 (N_20213,N_18014,N_18833);
and U20214 (N_20214,N_18107,N_18170);
or U20215 (N_20215,N_18689,N_18781);
xnor U20216 (N_20216,N_18812,N_19138);
or U20217 (N_20217,N_18519,N_19020);
nand U20218 (N_20218,N_18711,N_18634);
nand U20219 (N_20219,N_18498,N_19040);
nand U20220 (N_20220,N_18293,N_18425);
or U20221 (N_20221,N_18154,N_18207);
xor U20222 (N_20222,N_18356,N_18385);
nor U20223 (N_20223,N_18100,N_18778);
and U20224 (N_20224,N_18448,N_19128);
nor U20225 (N_20225,N_19097,N_18587);
and U20226 (N_20226,N_19004,N_18695);
and U20227 (N_20227,N_18599,N_18745);
or U20228 (N_20228,N_19169,N_18119);
nand U20229 (N_20229,N_18214,N_19120);
nand U20230 (N_20230,N_18663,N_18996);
nand U20231 (N_20231,N_19185,N_18628);
or U20232 (N_20232,N_18273,N_18483);
nor U20233 (N_20233,N_18374,N_18571);
nand U20234 (N_20234,N_18106,N_19093);
or U20235 (N_20235,N_18031,N_18742);
xor U20236 (N_20236,N_19007,N_18951);
and U20237 (N_20237,N_18526,N_18529);
xnor U20238 (N_20238,N_18053,N_18028);
nor U20239 (N_20239,N_18491,N_18485);
or U20240 (N_20240,N_19147,N_18385);
xor U20241 (N_20241,N_18695,N_18693);
and U20242 (N_20242,N_18525,N_18709);
or U20243 (N_20243,N_18191,N_18199);
nor U20244 (N_20244,N_18670,N_18916);
and U20245 (N_20245,N_18810,N_18426);
xnor U20246 (N_20246,N_18400,N_18536);
nand U20247 (N_20247,N_18018,N_18990);
xor U20248 (N_20248,N_18822,N_19040);
xnor U20249 (N_20249,N_18701,N_18499);
or U20250 (N_20250,N_18656,N_19101);
xor U20251 (N_20251,N_18057,N_18585);
nand U20252 (N_20252,N_18900,N_18396);
and U20253 (N_20253,N_18252,N_18606);
and U20254 (N_20254,N_18265,N_18673);
nand U20255 (N_20255,N_18013,N_18848);
or U20256 (N_20256,N_18658,N_18701);
nand U20257 (N_20257,N_18337,N_19145);
and U20258 (N_20258,N_19044,N_19001);
nand U20259 (N_20259,N_18505,N_18277);
or U20260 (N_20260,N_18017,N_18671);
or U20261 (N_20261,N_18967,N_18734);
and U20262 (N_20262,N_18383,N_18678);
and U20263 (N_20263,N_18335,N_18033);
or U20264 (N_20264,N_18946,N_18177);
nand U20265 (N_20265,N_18630,N_18609);
nand U20266 (N_20266,N_18671,N_18335);
nand U20267 (N_20267,N_18339,N_18718);
nor U20268 (N_20268,N_18731,N_18951);
or U20269 (N_20269,N_18891,N_18997);
or U20270 (N_20270,N_18668,N_18835);
or U20271 (N_20271,N_18792,N_18319);
and U20272 (N_20272,N_18562,N_18142);
or U20273 (N_20273,N_18180,N_18235);
xnor U20274 (N_20274,N_18952,N_19113);
and U20275 (N_20275,N_18934,N_18189);
xnor U20276 (N_20276,N_19101,N_18073);
nand U20277 (N_20277,N_18266,N_18130);
or U20278 (N_20278,N_18609,N_18890);
or U20279 (N_20279,N_19185,N_18083);
nor U20280 (N_20280,N_18220,N_18072);
xor U20281 (N_20281,N_18301,N_18312);
and U20282 (N_20282,N_19088,N_18056);
or U20283 (N_20283,N_19048,N_18828);
nor U20284 (N_20284,N_18535,N_18387);
nor U20285 (N_20285,N_18606,N_18499);
nand U20286 (N_20286,N_18482,N_18818);
nand U20287 (N_20287,N_19044,N_18877);
nor U20288 (N_20288,N_19007,N_18430);
or U20289 (N_20289,N_18253,N_18335);
and U20290 (N_20290,N_18607,N_18263);
xor U20291 (N_20291,N_19080,N_18453);
and U20292 (N_20292,N_18902,N_19148);
xnor U20293 (N_20293,N_19048,N_19171);
nand U20294 (N_20294,N_18877,N_18921);
xnor U20295 (N_20295,N_18569,N_18667);
nand U20296 (N_20296,N_19009,N_18876);
nand U20297 (N_20297,N_18884,N_18727);
nand U20298 (N_20298,N_18455,N_19099);
nor U20299 (N_20299,N_18815,N_18423);
xnor U20300 (N_20300,N_19061,N_18825);
nand U20301 (N_20301,N_18702,N_18022);
nor U20302 (N_20302,N_18602,N_18710);
nor U20303 (N_20303,N_18729,N_18607);
or U20304 (N_20304,N_18987,N_18737);
nand U20305 (N_20305,N_19122,N_18054);
xor U20306 (N_20306,N_19116,N_19195);
nor U20307 (N_20307,N_18079,N_18137);
nand U20308 (N_20308,N_19089,N_18774);
or U20309 (N_20309,N_18822,N_18191);
xor U20310 (N_20310,N_18123,N_19004);
xor U20311 (N_20311,N_18921,N_18059);
xor U20312 (N_20312,N_18010,N_18900);
and U20313 (N_20313,N_18650,N_18586);
or U20314 (N_20314,N_18374,N_18625);
xor U20315 (N_20315,N_18433,N_18773);
and U20316 (N_20316,N_18518,N_18856);
nand U20317 (N_20317,N_18577,N_18346);
or U20318 (N_20318,N_18800,N_18290);
nor U20319 (N_20319,N_18659,N_18453);
or U20320 (N_20320,N_18227,N_18015);
nor U20321 (N_20321,N_18984,N_18072);
and U20322 (N_20322,N_18409,N_18947);
xnor U20323 (N_20323,N_18658,N_18217);
nor U20324 (N_20324,N_18203,N_18730);
nor U20325 (N_20325,N_18829,N_18205);
nor U20326 (N_20326,N_18166,N_18760);
and U20327 (N_20327,N_18436,N_19131);
nor U20328 (N_20328,N_18399,N_18494);
nor U20329 (N_20329,N_18491,N_18075);
nor U20330 (N_20330,N_19115,N_18513);
and U20331 (N_20331,N_18230,N_19063);
and U20332 (N_20332,N_19090,N_18261);
nor U20333 (N_20333,N_18793,N_18693);
nand U20334 (N_20334,N_18429,N_18943);
or U20335 (N_20335,N_18673,N_18992);
xnor U20336 (N_20336,N_18719,N_18178);
nand U20337 (N_20337,N_18480,N_19017);
or U20338 (N_20338,N_19127,N_18979);
nand U20339 (N_20339,N_18665,N_18636);
nor U20340 (N_20340,N_18242,N_18502);
nor U20341 (N_20341,N_18031,N_18985);
nor U20342 (N_20342,N_18423,N_18543);
and U20343 (N_20343,N_19091,N_18543);
nor U20344 (N_20344,N_18534,N_18745);
nand U20345 (N_20345,N_18934,N_19162);
or U20346 (N_20346,N_18721,N_18546);
xor U20347 (N_20347,N_19184,N_18065);
xor U20348 (N_20348,N_18622,N_18119);
and U20349 (N_20349,N_18833,N_18907);
nand U20350 (N_20350,N_18039,N_18333);
or U20351 (N_20351,N_18468,N_19004);
nor U20352 (N_20352,N_18511,N_19142);
and U20353 (N_20353,N_18576,N_18463);
nand U20354 (N_20354,N_18477,N_18481);
or U20355 (N_20355,N_18599,N_18467);
nand U20356 (N_20356,N_18713,N_19045);
and U20357 (N_20357,N_18084,N_18531);
nor U20358 (N_20358,N_18320,N_18842);
and U20359 (N_20359,N_18182,N_19179);
or U20360 (N_20360,N_18363,N_18559);
xor U20361 (N_20361,N_18605,N_18266);
nand U20362 (N_20362,N_19157,N_18727);
xor U20363 (N_20363,N_18298,N_18659);
and U20364 (N_20364,N_18067,N_18492);
nand U20365 (N_20365,N_18333,N_19018);
or U20366 (N_20366,N_18113,N_18006);
or U20367 (N_20367,N_18345,N_18466);
xnor U20368 (N_20368,N_18659,N_19077);
or U20369 (N_20369,N_18205,N_18216);
and U20370 (N_20370,N_18366,N_18139);
or U20371 (N_20371,N_18122,N_18444);
or U20372 (N_20372,N_19125,N_18300);
and U20373 (N_20373,N_19007,N_18685);
or U20374 (N_20374,N_18113,N_18333);
nor U20375 (N_20375,N_18064,N_18582);
and U20376 (N_20376,N_18365,N_18793);
nand U20377 (N_20377,N_19139,N_18485);
xor U20378 (N_20378,N_19065,N_18901);
nor U20379 (N_20379,N_19048,N_19169);
and U20380 (N_20380,N_18750,N_18688);
and U20381 (N_20381,N_18512,N_18555);
nor U20382 (N_20382,N_18749,N_18346);
nand U20383 (N_20383,N_18109,N_18860);
xor U20384 (N_20384,N_18403,N_19126);
xnor U20385 (N_20385,N_18725,N_18056);
and U20386 (N_20386,N_18742,N_19114);
xnor U20387 (N_20387,N_18836,N_19088);
nand U20388 (N_20388,N_19000,N_18837);
nor U20389 (N_20389,N_18633,N_18131);
xnor U20390 (N_20390,N_18253,N_18831);
xor U20391 (N_20391,N_18513,N_18715);
nor U20392 (N_20392,N_19096,N_18771);
nor U20393 (N_20393,N_18343,N_18293);
and U20394 (N_20394,N_18779,N_19041);
nand U20395 (N_20395,N_19085,N_18172);
nor U20396 (N_20396,N_18720,N_18213);
nor U20397 (N_20397,N_18443,N_18370);
and U20398 (N_20398,N_18803,N_18101);
nor U20399 (N_20399,N_19106,N_18314);
xnor U20400 (N_20400,N_19518,N_19506);
or U20401 (N_20401,N_19975,N_20289);
or U20402 (N_20402,N_19278,N_19983);
or U20403 (N_20403,N_19366,N_19455);
and U20404 (N_20404,N_19250,N_19402);
and U20405 (N_20405,N_20129,N_19295);
and U20406 (N_20406,N_20100,N_20016);
or U20407 (N_20407,N_19880,N_20150);
or U20408 (N_20408,N_19809,N_19973);
xor U20409 (N_20409,N_19793,N_19474);
and U20410 (N_20410,N_20178,N_19376);
nand U20411 (N_20411,N_19274,N_20003);
or U20412 (N_20412,N_19240,N_19797);
nor U20413 (N_20413,N_19808,N_19993);
xnor U20414 (N_20414,N_19785,N_19755);
nor U20415 (N_20415,N_19919,N_19275);
or U20416 (N_20416,N_20374,N_20064);
nand U20417 (N_20417,N_19368,N_20130);
and U20418 (N_20418,N_19962,N_19675);
and U20419 (N_20419,N_19382,N_20190);
nor U20420 (N_20420,N_19902,N_20062);
nor U20421 (N_20421,N_19338,N_19556);
and U20422 (N_20422,N_19337,N_20164);
xnor U20423 (N_20423,N_19583,N_20339);
xor U20424 (N_20424,N_20136,N_19824);
nand U20425 (N_20425,N_20195,N_19372);
or U20426 (N_20426,N_19231,N_19744);
xnor U20427 (N_20427,N_19497,N_19513);
nand U20428 (N_20428,N_20207,N_19303);
nor U20429 (N_20429,N_20093,N_20181);
and U20430 (N_20430,N_19780,N_19763);
and U20431 (N_20431,N_20364,N_19604);
nand U20432 (N_20432,N_19268,N_19498);
or U20433 (N_20433,N_20302,N_19897);
nor U20434 (N_20434,N_19634,N_19924);
nor U20435 (N_20435,N_20091,N_19784);
or U20436 (N_20436,N_19296,N_19456);
nand U20437 (N_20437,N_20345,N_20312);
xnor U20438 (N_20438,N_19655,N_20066);
nor U20439 (N_20439,N_20162,N_20291);
or U20440 (N_20440,N_19596,N_19531);
xnor U20441 (N_20441,N_19994,N_20223);
nor U20442 (N_20442,N_20191,N_19750);
nand U20443 (N_20443,N_20336,N_20298);
or U20444 (N_20444,N_19798,N_19332);
and U20445 (N_20445,N_19699,N_19917);
nor U20446 (N_20446,N_20173,N_19363);
or U20447 (N_20447,N_19535,N_20358);
or U20448 (N_20448,N_19563,N_20228);
nand U20449 (N_20449,N_19788,N_19595);
and U20450 (N_20450,N_20176,N_19454);
or U20451 (N_20451,N_19626,N_20246);
xnor U20452 (N_20452,N_19986,N_19321);
nor U20453 (N_20453,N_20155,N_19311);
xor U20454 (N_20454,N_19606,N_19555);
nand U20455 (N_20455,N_19777,N_20180);
xor U20456 (N_20456,N_20252,N_19616);
and U20457 (N_20457,N_20069,N_20141);
and U20458 (N_20458,N_19949,N_19249);
or U20459 (N_20459,N_19613,N_20363);
xnor U20460 (N_20460,N_19310,N_19442);
xnor U20461 (N_20461,N_19217,N_19876);
or U20462 (N_20462,N_19682,N_19804);
or U20463 (N_20463,N_19894,N_19377);
and U20464 (N_20464,N_19437,N_19742);
and U20465 (N_20465,N_19668,N_20054);
nor U20466 (N_20466,N_19749,N_19248);
nand U20467 (N_20467,N_19371,N_19812);
or U20468 (N_20468,N_20254,N_20007);
xnor U20469 (N_20469,N_20056,N_20206);
nor U20470 (N_20470,N_19968,N_20037);
or U20471 (N_20471,N_19656,N_19225);
nor U20472 (N_20472,N_20047,N_20184);
xnor U20473 (N_20473,N_19988,N_20186);
nor U20474 (N_20474,N_19731,N_20103);
nand U20475 (N_20475,N_20175,N_19428);
xnor U20476 (N_20476,N_19920,N_20273);
xnor U20477 (N_20477,N_19667,N_19701);
xor U20478 (N_20478,N_20392,N_20219);
nor U20479 (N_20479,N_19642,N_19739);
or U20480 (N_20480,N_19657,N_20380);
and U20481 (N_20481,N_20170,N_19692);
nor U20482 (N_20482,N_20341,N_19598);
nand U20483 (N_20483,N_19503,N_19270);
and U20484 (N_20484,N_20307,N_19233);
and U20485 (N_20485,N_20073,N_19888);
and U20486 (N_20486,N_19805,N_20095);
xnor U20487 (N_20487,N_19290,N_19541);
or U20488 (N_20488,N_20352,N_19416);
or U20489 (N_20489,N_20032,N_19971);
nand U20490 (N_20490,N_19704,N_20147);
nor U20491 (N_20491,N_20010,N_20269);
and U20492 (N_20492,N_20027,N_20031);
nor U20493 (N_20493,N_19773,N_19825);
and U20494 (N_20494,N_19457,N_20247);
xnor U20495 (N_20495,N_19234,N_20264);
xor U20496 (N_20496,N_20058,N_20179);
nor U20497 (N_20497,N_19863,N_19424);
nand U20498 (N_20498,N_19569,N_19680);
and U20499 (N_20499,N_19412,N_20212);
xnor U20500 (N_20500,N_19536,N_20088);
xnor U20501 (N_20501,N_20359,N_19453);
nand U20502 (N_20502,N_20393,N_19935);
xor U20503 (N_20503,N_19410,N_19215);
nor U20504 (N_20504,N_19512,N_20134);
xnor U20505 (N_20505,N_20123,N_20396);
or U20506 (N_20506,N_19212,N_19914);
or U20507 (N_20507,N_20121,N_19426);
xnor U20508 (N_20508,N_19407,N_19911);
and U20509 (N_20509,N_20376,N_19817);
xnor U20510 (N_20510,N_19482,N_20232);
xnor U20511 (N_20511,N_19253,N_19979);
nand U20512 (N_20512,N_20000,N_19671);
and U20513 (N_20513,N_19326,N_19725);
xnor U20514 (N_20514,N_20194,N_19283);
or U20515 (N_20515,N_20024,N_19520);
nand U20516 (N_20516,N_19548,N_19413);
nand U20517 (N_20517,N_20231,N_20131);
and U20518 (N_20518,N_19359,N_19389);
nand U20519 (N_20519,N_19458,N_19411);
nand U20520 (N_20520,N_19459,N_19939);
nand U20521 (N_20521,N_19961,N_20391);
or U20522 (N_20522,N_19833,N_19517);
xnor U20523 (N_20523,N_19877,N_19850);
and U20524 (N_20524,N_20398,N_19965);
nor U20525 (N_20525,N_20048,N_20317);
xor U20526 (N_20526,N_20038,N_19349);
or U20527 (N_20527,N_19844,N_19540);
and U20528 (N_20528,N_20119,N_19907);
xnor U20529 (N_20529,N_20357,N_19216);
nor U20530 (N_20530,N_19473,N_19272);
xnor U20531 (N_20531,N_20140,N_20285);
nand U20532 (N_20532,N_20015,N_19329);
nor U20533 (N_20533,N_20373,N_20059);
xnor U20534 (N_20534,N_19687,N_19855);
or U20535 (N_20535,N_20314,N_20193);
and U20536 (N_20536,N_19207,N_19714);
nor U20537 (N_20537,N_19209,N_20222);
and U20538 (N_20538,N_19460,N_19528);
nand U20539 (N_20539,N_19519,N_19882);
and U20540 (N_20540,N_20294,N_19741);
or U20541 (N_20541,N_19351,N_19846);
or U20542 (N_20542,N_19401,N_20163);
xnor U20543 (N_20543,N_19969,N_20049);
nand U20544 (N_20544,N_19943,N_19251);
nor U20545 (N_20545,N_20267,N_19673);
nand U20546 (N_20546,N_19779,N_19735);
nor U20547 (N_20547,N_19868,N_20125);
nand U20548 (N_20548,N_19334,N_19849);
and U20549 (N_20549,N_19489,N_19345);
or U20550 (N_20550,N_19972,N_19764);
and U20551 (N_20551,N_20282,N_19466);
nor U20552 (N_20552,N_19931,N_20253);
nor U20553 (N_20553,N_19679,N_19417);
nor U20554 (N_20554,N_19461,N_20205);
xnor U20555 (N_20555,N_20310,N_19883);
xor U20556 (N_20556,N_20168,N_19926);
or U20557 (N_20557,N_19355,N_19650);
nand U20558 (N_20558,N_19653,N_19832);
nor U20559 (N_20559,N_19484,N_19645);
or U20560 (N_20560,N_19226,N_19930);
xnor U20561 (N_20561,N_20331,N_20199);
nand U20562 (N_20562,N_19636,N_19342);
and U20563 (N_20563,N_19245,N_20126);
nor U20564 (N_20564,N_19947,N_19383);
xnor U20565 (N_20565,N_20114,N_19759);
nand U20566 (N_20566,N_19840,N_19698);
or U20567 (N_20567,N_19271,N_19490);
or U20568 (N_20568,N_19652,N_19887);
nor U20569 (N_20569,N_20323,N_19745);
and U20570 (N_20570,N_19823,N_19767);
or U20571 (N_20571,N_19669,N_20244);
xor U20572 (N_20572,N_20145,N_20237);
and U20573 (N_20573,N_20337,N_19884);
and U20574 (N_20574,N_19591,N_19238);
nand U20575 (N_20575,N_19862,N_20109);
xnor U20576 (N_20576,N_20258,N_19605);
xor U20577 (N_20577,N_19927,N_20278);
nand U20578 (N_20578,N_19206,N_19452);
and U20579 (N_20579,N_19953,N_19493);
or U20580 (N_20580,N_19553,N_20213);
xnor U20581 (N_20581,N_20096,N_19241);
nand U20582 (N_20582,N_19958,N_20224);
xnor U20583 (N_20583,N_19550,N_19827);
xor U20584 (N_20584,N_20240,N_19500);
and U20585 (N_20585,N_19247,N_19491);
or U20586 (N_20586,N_20152,N_20350);
nor U20587 (N_20587,N_19587,N_19878);
and U20588 (N_20588,N_19752,N_19436);
or U20589 (N_20589,N_20221,N_19478);
or U20590 (N_20590,N_19505,N_19703);
nor U20591 (N_20591,N_19895,N_19463);
and U20592 (N_20592,N_19348,N_19866);
xnor U20593 (N_20593,N_20297,N_19398);
nor U20594 (N_20594,N_19921,N_20166);
nor U20595 (N_20595,N_19721,N_20045);
nand U20596 (N_20596,N_19946,N_19792);
and U20597 (N_20597,N_20292,N_19558);
nand U20598 (N_20598,N_19288,N_20068);
xnor U20599 (N_20599,N_20160,N_19302);
xnor U20600 (N_20600,N_19347,N_19542);
nor U20601 (N_20601,N_20355,N_19663);
nor U20602 (N_20602,N_19783,N_19813);
xnor U20603 (N_20603,N_20375,N_19945);
or U20604 (N_20604,N_19480,N_19942);
nor U20605 (N_20605,N_19632,N_20013);
nand U20606 (N_20606,N_19621,N_20137);
nand U20607 (N_20607,N_19559,N_19423);
or U20608 (N_20608,N_19881,N_19421);
and U20609 (N_20609,N_19904,N_20270);
xnor U20610 (N_20610,N_19638,N_20251);
or U20611 (N_20611,N_20128,N_20177);
nand U20612 (N_20612,N_19434,N_20209);
xor U20613 (N_20613,N_19778,N_20110);
xnor U20614 (N_20614,N_19603,N_20072);
xnor U20615 (N_20615,N_20116,N_19891);
nand U20616 (N_20616,N_19677,N_20395);
xnor U20617 (N_20617,N_19719,N_20120);
nor U20618 (N_20618,N_19370,N_20306);
and U20619 (N_20619,N_19369,N_20020);
or U20620 (N_20620,N_19210,N_19678);
nor U20621 (N_20621,N_19614,N_20148);
or U20622 (N_20622,N_20390,N_19400);
nand U20623 (N_20623,N_19952,N_19765);
and U20624 (N_20624,N_19639,N_19399);
or U20625 (N_20625,N_19537,N_19835);
nor U20626 (N_20626,N_19589,N_20265);
nor U20627 (N_20627,N_19254,N_19425);
nand U20628 (N_20628,N_19590,N_19799);
nor U20629 (N_20629,N_19486,N_19600);
and U20630 (N_20630,N_20012,N_19906);
nand U20631 (N_20631,N_19305,N_19633);
nor U20632 (N_20632,N_19211,N_19847);
nand U20633 (N_20633,N_20284,N_19912);
and U20634 (N_20634,N_19715,N_19859);
nor U20635 (N_20635,N_19774,N_19758);
and U20636 (N_20636,N_20324,N_19405);
nand U20637 (N_20637,N_19918,N_19658);
or U20638 (N_20638,N_20034,N_20085);
nor U20639 (N_20639,N_20234,N_19913);
nor U20640 (N_20640,N_19727,N_20192);
and U20641 (N_20641,N_19432,N_19343);
nor U20642 (N_20642,N_19997,N_19681);
nand U20643 (N_20643,N_19447,N_19397);
or U20644 (N_20644,N_19996,N_19601);
or U20645 (N_20645,N_20262,N_19718);
or U20646 (N_20646,N_19430,N_19893);
or U20647 (N_20647,N_19872,N_19551);
xnor U20648 (N_20648,N_20074,N_19365);
nor U20649 (N_20649,N_20378,N_19854);
and U20650 (N_20650,N_19716,N_20115);
xor U20651 (N_20651,N_19890,N_19230);
or U20652 (N_20652,N_19340,N_20321);
and U20653 (N_20653,N_20379,N_19861);
xor U20654 (N_20654,N_19379,N_20060);
xor U20655 (N_20655,N_20362,N_20102);
and U20656 (N_20656,N_20233,N_19285);
or U20657 (N_20657,N_19282,N_19746);
nor U20658 (N_20658,N_20215,N_19408);
xnor U20659 (N_20659,N_20287,N_19322);
xnor U20660 (N_20660,N_20335,N_20342);
nand U20661 (N_20661,N_20142,N_19409);
nand U20662 (N_20662,N_19403,N_19267);
xnor U20663 (N_20663,N_20005,N_19481);
nand U20664 (N_20664,N_19929,N_20318);
xnor U20665 (N_20665,N_20139,N_19915);
nand U20666 (N_20666,N_19448,N_19415);
or U20667 (N_20667,N_20332,N_19373);
nor U20668 (N_20668,N_19244,N_19469);
xnor U20669 (N_20669,N_20182,N_20260);
nand U20670 (N_20670,N_20344,N_20198);
nand U20671 (N_20671,N_20249,N_19978);
nand U20672 (N_20672,N_19566,N_19853);
and U20673 (N_20673,N_20075,N_19562);
or U20674 (N_20674,N_19393,N_19235);
or U20675 (N_20675,N_19950,N_20320);
or U20676 (N_20676,N_19255,N_20236);
nor U20677 (N_20677,N_19269,N_20356);
or U20678 (N_20678,N_20361,N_20377);
nor U20679 (N_20679,N_19564,N_20227);
nor U20680 (N_20680,N_19350,N_19304);
or U20681 (N_20681,N_19628,N_19602);
or U20682 (N_20682,N_19928,N_19495);
xnor U20683 (N_20683,N_19521,N_20248);
nor U20684 (N_20684,N_19769,N_19567);
and U20685 (N_20685,N_19830,N_20238);
nand U20686 (N_20686,N_19236,N_19710);
and U20687 (N_20687,N_19916,N_20208);
or U20688 (N_20688,N_19574,N_20017);
and U20689 (N_20689,N_19967,N_19510);
nor U20690 (N_20690,N_19896,N_19511);
xor U20691 (N_20691,N_20187,N_19858);
or U20692 (N_20692,N_19843,N_20372);
or U20693 (N_20693,N_19756,N_19957);
or U20694 (N_20694,N_19357,N_20353);
and U20695 (N_20695,N_19790,N_19900);
xor U20696 (N_20696,N_19297,N_19795);
nor U20697 (N_20697,N_20360,N_19406);
xor U20698 (N_20698,N_19289,N_19757);
or U20699 (N_20699,N_20122,N_19509);
nor U20700 (N_20700,N_19529,N_20197);
nand U20701 (N_20701,N_19593,N_19728);
or U20702 (N_20702,N_20280,N_19546);
nand U20703 (N_20703,N_19989,N_20019);
xnor U20704 (N_20704,N_19451,N_19237);
or U20705 (N_20705,N_19787,N_20053);
xor U20706 (N_20706,N_20239,N_20394);
or U20707 (N_20707,N_20347,N_19573);
nor U20708 (N_20708,N_19985,N_20018);
nand U20709 (N_20709,N_19258,N_20283);
or U20710 (N_20710,N_20041,N_19609);
or U20711 (N_20711,N_19584,N_20250);
nor U20712 (N_20712,N_20081,N_19545);
or U20713 (N_20713,N_19525,N_19360);
and U20714 (N_20714,N_19539,N_19284);
nor U20715 (N_20715,N_19472,N_19312);
nand U20716 (N_20716,N_19821,N_19875);
nor U20717 (N_20717,N_19819,N_20300);
and U20718 (N_20718,N_19433,N_19222);
nand U20719 (N_20719,N_20387,N_19966);
xor U20720 (N_20720,N_19361,N_20001);
nor U20721 (N_20721,N_20089,N_19328);
or U20722 (N_20722,N_19910,N_19273);
or U20723 (N_20723,N_20382,N_19676);
or U20724 (N_20724,N_20290,N_19610);
nand U20725 (N_20725,N_19353,N_19324);
nand U20726 (N_20726,N_19292,N_20305);
nand U20727 (N_20727,N_19580,N_20325);
xor U20728 (N_20728,N_19674,N_20006);
or U20729 (N_20729,N_20326,N_20025);
or U20730 (N_20730,N_19316,N_19740);
and U20731 (N_20731,N_19737,N_19445);
xor U20732 (N_20732,N_19816,N_19419);
nor U20733 (N_20733,N_20009,N_20225);
and U20734 (N_20734,N_19625,N_20022);
nor U20735 (N_20735,N_19641,N_19651);
and U20736 (N_20736,N_19483,N_19631);
xor U20737 (N_20737,N_19227,N_19261);
and U20738 (N_20738,N_19314,N_19836);
xor U20739 (N_20739,N_19839,N_19470);
and U20740 (N_20740,N_20214,N_20386);
or U20741 (N_20741,N_20077,N_20189);
and U20742 (N_20742,N_19526,N_19577);
xnor U20743 (N_20743,N_20381,N_19837);
and U20744 (N_20744,N_19747,N_20111);
nand U20745 (N_20745,N_20351,N_20105);
and U20746 (N_20746,N_20098,N_19695);
nor U20747 (N_20747,N_19586,N_19335);
nor U20748 (N_20748,N_19782,N_20296);
or U20749 (N_20749,N_19879,N_19257);
xor U20750 (N_20750,N_19786,N_20055);
nand U20751 (N_20751,N_19909,N_19477);
nand U20752 (N_20752,N_19706,N_19892);
xnor U20753 (N_20753,N_19299,N_20117);
nand U20754 (N_20754,N_19256,N_20080);
nor U20755 (N_20755,N_19803,N_19391);
nand U20756 (N_20756,N_20274,N_19732);
xor U20757 (N_20757,N_19615,N_19970);
and U20758 (N_20758,N_19309,N_19560);
and U20759 (N_20759,N_20349,N_19441);
nand U20760 (N_20760,N_19647,N_20021);
nor U20761 (N_20761,N_20368,N_20002);
xor U20762 (N_20762,N_19834,N_19640);
xor U20763 (N_20763,N_19646,N_20008);
xnor U20764 (N_20764,N_20241,N_19286);
and U20765 (N_20765,N_20385,N_20084);
and U20766 (N_20766,N_19422,N_19374);
xor U20767 (N_20767,N_19940,N_20065);
and U20768 (N_20768,N_19575,N_20295);
or U20769 (N_20769,N_20133,N_20043);
nand U20770 (N_20770,N_19362,N_19934);
nor U20771 (N_20771,N_19205,N_20156);
nor U20772 (N_20772,N_19886,N_19726);
nand U20773 (N_20773,N_19629,N_20050);
xnor U20774 (N_20774,N_19418,N_19870);
and U20775 (N_20775,N_19462,N_20172);
nand U20776 (N_20776,N_20078,N_20046);
and U20777 (N_20777,N_19867,N_19390);
nor U20778 (N_20778,N_20023,N_20067);
and U20779 (N_20779,N_19814,N_19762);
xnor U20780 (N_20780,N_20044,N_19578);
and U20781 (N_20781,N_19694,N_19766);
and U20782 (N_20782,N_19800,N_19828);
xnor U20783 (N_20783,N_19683,N_20322);
nor U20784 (N_20784,N_19775,N_19826);
or U20785 (N_20785,N_20153,N_19307);
or U20786 (N_20786,N_19364,N_19709);
and U20787 (N_20787,N_19533,N_20370);
nand U20788 (N_20788,N_20255,N_20301);
and U20789 (N_20789,N_20201,N_20281);
and U20790 (N_20790,N_19485,N_19807);
or U20791 (N_20791,N_20245,N_19789);
and U20792 (N_20792,N_20303,N_19262);
or U20793 (N_20793,N_19672,N_19937);
xnor U20794 (N_20794,N_19776,N_20333);
or U20795 (N_20795,N_19960,N_19501);
and U20796 (N_20796,N_19330,N_19392);
nand U20797 (N_20797,N_19464,N_19291);
nand U20798 (N_20798,N_19354,N_19246);
or U20799 (N_20799,N_19822,N_19228);
xor U20800 (N_20800,N_20171,N_19339);
or U20801 (N_20801,N_19358,N_19708);
and U20802 (N_20802,N_19543,N_19933);
and U20803 (N_20803,N_20143,N_19630);
and U20804 (N_20804,N_20327,N_19443);
or U20805 (N_20805,N_19523,N_19991);
xor U20806 (N_20806,N_20257,N_20135);
xnor U20807 (N_20807,N_19208,N_20154);
nor U20808 (N_20808,N_20112,N_19869);
or U20809 (N_20809,N_19333,N_19308);
xnor U20810 (N_20810,N_19221,N_20316);
and U20811 (N_20811,N_19252,N_19751);
or U20812 (N_20812,N_19925,N_20200);
xor U20813 (N_20813,N_20242,N_20397);
or U20814 (N_20814,N_20161,N_19874);
xor U20815 (N_20815,N_20159,N_20330);
and U20816 (N_20816,N_19643,N_19707);
xnor U20817 (N_20817,N_19557,N_20061);
or U20818 (N_20818,N_20086,N_19838);
nand U20819 (N_20819,N_20279,N_19885);
nor U20820 (N_20820,N_20203,N_19223);
nand U20821 (N_20821,N_19588,N_19612);
or U20822 (N_20822,N_19565,N_19637);
xor U20823 (N_20823,N_19494,N_20243);
nor U20824 (N_20824,N_19220,N_19956);
and U20825 (N_20825,N_20271,N_20204);
nor U20826 (N_20826,N_19871,N_19815);
nor U20827 (N_20827,N_20315,N_19738);
nand U20828 (N_20828,N_19396,N_20210);
nor U20829 (N_20829,N_20399,N_19218);
xnor U20830 (N_20830,N_19977,N_19748);
and U20831 (N_20831,N_20348,N_19395);
or U20832 (N_20832,N_19923,N_19772);
or U20833 (N_20833,N_20108,N_19903);
nand U20834 (N_20834,N_20169,N_19488);
nor U20835 (N_20835,N_20226,N_19260);
and U20836 (N_20836,N_19955,N_20174);
nand U20837 (N_20837,N_19224,N_19623);
nand U20838 (N_20838,N_20235,N_19857);
nand U20839 (N_20839,N_19507,N_20196);
xnor U20840 (N_20840,N_19277,N_20094);
nand U20841 (N_20841,N_20127,N_19831);
or U20842 (N_20842,N_19331,N_19214);
nor U20843 (N_20843,N_19736,N_19684);
nor U20844 (N_20844,N_19948,N_19554);
and U20845 (N_20845,N_19980,N_19702);
nor U20846 (N_20846,N_19898,N_20149);
and U20847 (N_20847,N_19380,N_19239);
xnor U20848 (N_20848,N_19743,N_19381);
or U20849 (N_20849,N_19514,N_20082);
and U20850 (N_20850,N_19992,N_19524);
or U20851 (N_20851,N_19515,N_19298);
nor U20852 (N_20852,N_19300,N_19502);
nor U20853 (N_20853,N_20124,N_19976);
nor U20854 (N_20854,N_20011,N_19611);
nand U20855 (N_20855,N_19202,N_20158);
nand U20856 (N_20856,N_19508,N_19323);
and U20857 (N_20857,N_19753,N_20083);
or U20858 (N_20858,N_19689,N_19378);
and U20859 (N_20859,N_19999,N_19654);
xor U20860 (N_20860,N_19734,N_20101);
nor U20861 (N_20861,N_19315,N_19781);
or U20862 (N_20862,N_19771,N_20288);
nor U20863 (N_20863,N_19982,N_19908);
and U20864 (N_20864,N_20052,N_20343);
or U20865 (N_20865,N_19346,N_19901);
and U20866 (N_20866,N_19627,N_19889);
nand U20867 (N_20867,N_20218,N_19995);
and U20868 (N_20868,N_19325,N_19344);
xor U20869 (N_20869,N_19665,N_19276);
or U20870 (N_20870,N_19691,N_19530);
nand U20871 (N_20871,N_19487,N_19713);
or U20872 (N_20872,N_19649,N_20113);
and U20873 (N_20873,N_19319,N_19404);
nor U20874 (N_20874,N_19522,N_19499);
nor U20875 (N_20875,N_19845,N_19696);
or U20876 (N_20876,N_19852,N_19243);
xnor U20877 (N_20877,N_19287,N_19317);
and U20878 (N_20878,N_20272,N_19386);
or U20879 (N_20879,N_19794,N_19571);
and U20880 (N_20880,N_19729,N_20346);
xor U20881 (N_20881,N_19444,N_19791);
nor U20882 (N_20882,N_19984,N_20146);
or U20883 (N_20883,N_19301,N_20388);
or U20884 (N_20884,N_19266,N_20220);
and U20885 (N_20885,N_19761,N_19941);
nor U20886 (N_20886,N_19387,N_19905);
nand U20887 (N_20887,N_19547,N_20217);
nor U20888 (N_20888,N_20014,N_19414);
or U20889 (N_20889,N_19607,N_20026);
nand U20890 (N_20890,N_20076,N_19320);
nand U20891 (N_20891,N_19492,N_19219);
or U20892 (N_20892,N_20299,N_19644);
nand U20893 (N_20893,N_19842,N_20216);
xnor U20894 (N_20894,N_19306,N_20151);
or U20895 (N_20895,N_19561,N_19873);
or U20896 (N_20896,N_19468,N_19465);
or U20897 (N_20897,N_19711,N_19951);
nor U20898 (N_20898,N_20167,N_20266);
or U20899 (N_20899,N_19532,N_20329);
nor U20900 (N_20900,N_19229,N_19232);
xor U20901 (N_20901,N_19959,N_20366);
or U20902 (N_20902,N_19720,N_20029);
and U20903 (N_20903,N_19450,N_19659);
and U20904 (N_20904,N_19313,N_19848);
and U20905 (N_20905,N_19899,N_20118);
or U20906 (N_20906,N_19662,N_19856);
xnor U20907 (N_20907,N_20211,N_20107);
nand U20908 (N_20908,N_20371,N_19618);
or U20909 (N_20909,N_19932,N_20230);
nor U20910 (N_20910,N_19730,N_20365);
xor U20911 (N_20911,N_20309,N_19476);
nor U20912 (N_20912,N_19594,N_20097);
and U20913 (N_20913,N_20340,N_19697);
xnor U20914 (N_20914,N_20334,N_19705);
or U20915 (N_20915,N_19435,N_19864);
nand U20916 (N_20916,N_19527,N_19724);
and U20917 (N_20917,N_19624,N_19635);
nor U20918 (N_20918,N_19664,N_19936);
xor U20919 (N_20919,N_20202,N_19981);
and U20920 (N_20920,N_20063,N_19427);
nor U20921 (N_20921,N_19204,N_19811);
and U20922 (N_20922,N_20338,N_19582);
nand U20923 (N_20923,N_19352,N_19356);
nor U20924 (N_20924,N_19475,N_20259);
xnor U20925 (N_20925,N_19964,N_20090);
xor U20926 (N_20926,N_19722,N_20070);
nor U20927 (N_20927,N_19394,N_20071);
nor U20928 (N_20928,N_20293,N_19693);
xnor U20929 (N_20929,N_19585,N_19576);
and U20930 (N_20930,N_19712,N_19440);
nand U20931 (N_20931,N_19568,N_20308);
and U20932 (N_20932,N_19294,N_20087);
and U20933 (N_20933,N_20183,N_19599);
and U20934 (N_20934,N_19686,N_19263);
or U20935 (N_20935,N_19471,N_19384);
nor U20936 (N_20936,N_20099,N_20383);
and U20937 (N_20937,N_20106,N_19754);
nand U20938 (N_20938,N_20004,N_20028);
nand U20939 (N_20939,N_19367,N_20229);
or U20940 (N_20940,N_19341,N_20328);
and U20941 (N_20941,N_19375,N_19572);
xor U20942 (N_20942,N_19818,N_19619);
or U20943 (N_20943,N_19796,N_19922);
or U20944 (N_20944,N_19648,N_19620);
nor U20945 (N_20945,N_19534,N_20036);
or U20946 (N_20946,N_19608,N_19293);
and U20947 (N_20947,N_19259,N_20033);
and U20948 (N_20948,N_19938,N_20286);
nand U20949 (N_20949,N_19579,N_20311);
xnor U20950 (N_20950,N_19770,N_19661);
or U20951 (N_20951,N_19570,N_19336);
xnor U20952 (N_20952,N_19700,N_20319);
and U20953 (N_20953,N_19504,N_20040);
and U20954 (N_20954,N_19449,N_19597);
or U20955 (N_20955,N_19851,N_19829);
and U20956 (N_20956,N_19496,N_19944);
nand U20957 (N_20957,N_19987,N_20138);
nand U20958 (N_20958,N_19860,N_19760);
nor U20959 (N_20959,N_20165,N_19439);
or U20960 (N_20960,N_19420,N_19841);
xor U20961 (N_20961,N_19820,N_20039);
nand U20962 (N_20962,N_20185,N_19690);
nor U20963 (N_20963,N_20263,N_19429);
nand U20964 (N_20964,N_20035,N_19552);
nor U20965 (N_20965,N_19279,N_20369);
nand U20966 (N_20966,N_20104,N_19688);
or U20967 (N_20967,N_19581,N_20157);
nor U20968 (N_20968,N_19516,N_20367);
xor U20969 (N_20969,N_19733,N_19670);
or U20970 (N_20970,N_19213,N_19479);
nor U20971 (N_20971,N_19280,N_20144);
nor U20972 (N_20972,N_19622,N_20042);
and U20973 (N_20973,N_19666,N_19990);
xnor U20974 (N_20974,N_19200,N_19963);
or U20975 (N_20975,N_20313,N_20261);
and U20976 (N_20976,N_19768,N_19592);
nor U20977 (N_20977,N_20030,N_19954);
and U20978 (N_20978,N_20057,N_19974);
nor U20979 (N_20979,N_19281,N_20092);
xnor U20980 (N_20980,N_19544,N_19327);
and U20981 (N_20981,N_19998,N_20276);
and U20982 (N_20982,N_19264,N_19617);
xor U20983 (N_20983,N_20384,N_20132);
or U20984 (N_20984,N_19265,N_20268);
xor U20985 (N_20985,N_19806,N_20051);
and U20986 (N_20986,N_20354,N_19388);
or U20987 (N_20987,N_19467,N_19549);
nor U20988 (N_20988,N_19242,N_19717);
nor U20989 (N_20989,N_19446,N_19660);
nand U20990 (N_20990,N_19203,N_19538);
xnor U20991 (N_20991,N_19723,N_20188);
and U20992 (N_20992,N_20275,N_19201);
or U20993 (N_20993,N_20389,N_20304);
and U20994 (N_20994,N_20256,N_19318);
and U20995 (N_20995,N_19865,N_19431);
and U20996 (N_20996,N_19385,N_20079);
nand U20997 (N_20997,N_19801,N_19685);
nand U20998 (N_20998,N_20277,N_19810);
and U20999 (N_20999,N_19802,N_19438);
nand U21000 (N_21000,N_19532,N_20312);
xnor U21001 (N_21001,N_19685,N_19665);
nand U21002 (N_21002,N_20040,N_19503);
and U21003 (N_21003,N_20121,N_19240);
and U21004 (N_21004,N_20300,N_20164);
xor U21005 (N_21005,N_20212,N_19730);
xor U21006 (N_21006,N_19930,N_19370);
and U21007 (N_21007,N_20037,N_19485);
nor U21008 (N_21008,N_20118,N_20227);
xor U21009 (N_21009,N_19642,N_19385);
nor U21010 (N_21010,N_19500,N_20125);
nor U21011 (N_21011,N_19380,N_19602);
or U21012 (N_21012,N_20339,N_19388);
xnor U21013 (N_21013,N_19260,N_19907);
xor U21014 (N_21014,N_20329,N_20181);
and U21015 (N_21015,N_19938,N_19251);
nor U21016 (N_21016,N_20294,N_19961);
nand U21017 (N_21017,N_20134,N_20079);
xor U21018 (N_21018,N_20322,N_20029);
and U21019 (N_21019,N_20224,N_19659);
or U21020 (N_21020,N_19658,N_19621);
and U21021 (N_21021,N_19950,N_20222);
or U21022 (N_21022,N_19695,N_19204);
or U21023 (N_21023,N_20312,N_19432);
nor U21024 (N_21024,N_19743,N_20392);
and U21025 (N_21025,N_20320,N_19473);
nor U21026 (N_21026,N_19866,N_20227);
nor U21027 (N_21027,N_19416,N_19269);
nor U21028 (N_21028,N_19906,N_19333);
xnor U21029 (N_21029,N_19721,N_19625);
nand U21030 (N_21030,N_19322,N_20310);
nand U21031 (N_21031,N_19822,N_19979);
xnor U21032 (N_21032,N_19476,N_20194);
nand U21033 (N_21033,N_19824,N_19691);
xnor U21034 (N_21034,N_19644,N_19546);
and U21035 (N_21035,N_19407,N_19848);
and U21036 (N_21036,N_19988,N_20208);
and U21037 (N_21037,N_19411,N_19815);
or U21038 (N_21038,N_19733,N_19525);
xnor U21039 (N_21039,N_19916,N_19271);
and U21040 (N_21040,N_19707,N_19724);
xor U21041 (N_21041,N_20199,N_19255);
nand U21042 (N_21042,N_19431,N_19853);
xnor U21043 (N_21043,N_19872,N_19700);
and U21044 (N_21044,N_19478,N_20225);
nor U21045 (N_21045,N_19337,N_19784);
nor U21046 (N_21046,N_19941,N_19472);
and U21047 (N_21047,N_19632,N_19621);
and U21048 (N_21048,N_19215,N_19358);
nand U21049 (N_21049,N_19981,N_20178);
and U21050 (N_21050,N_20211,N_19535);
xnor U21051 (N_21051,N_20275,N_20304);
xor U21052 (N_21052,N_19684,N_19559);
and U21053 (N_21053,N_20046,N_19886);
xor U21054 (N_21054,N_19954,N_19948);
and U21055 (N_21055,N_20388,N_20196);
nand U21056 (N_21056,N_19846,N_19409);
or U21057 (N_21057,N_19368,N_19388);
or U21058 (N_21058,N_20206,N_19651);
xor U21059 (N_21059,N_20291,N_19913);
xor U21060 (N_21060,N_19221,N_19604);
or U21061 (N_21061,N_20322,N_20382);
nor U21062 (N_21062,N_19632,N_19709);
xor U21063 (N_21063,N_19558,N_19209);
nor U21064 (N_21064,N_19861,N_20260);
nor U21065 (N_21065,N_19444,N_19680);
nand U21066 (N_21066,N_19767,N_19424);
nor U21067 (N_21067,N_19407,N_20320);
or U21068 (N_21068,N_19581,N_19905);
or U21069 (N_21069,N_20286,N_19379);
nand U21070 (N_21070,N_19460,N_19993);
or U21071 (N_21071,N_19505,N_19332);
and U21072 (N_21072,N_20259,N_19506);
and U21073 (N_21073,N_19802,N_19852);
and U21074 (N_21074,N_19339,N_19560);
xor U21075 (N_21075,N_19279,N_20126);
xnor U21076 (N_21076,N_19384,N_19832);
xnor U21077 (N_21077,N_19934,N_19823);
or U21078 (N_21078,N_19816,N_19603);
or U21079 (N_21079,N_19795,N_19377);
nor U21080 (N_21080,N_19279,N_19538);
nand U21081 (N_21081,N_19917,N_19638);
nor U21082 (N_21082,N_19695,N_20170);
and U21083 (N_21083,N_20068,N_19972);
or U21084 (N_21084,N_19656,N_20237);
nor U21085 (N_21085,N_19774,N_19286);
or U21086 (N_21086,N_19611,N_19754);
nor U21087 (N_21087,N_19251,N_20166);
xnor U21088 (N_21088,N_20113,N_19679);
and U21089 (N_21089,N_20072,N_19971);
nor U21090 (N_21090,N_19406,N_20314);
or U21091 (N_21091,N_19603,N_19470);
nand U21092 (N_21092,N_20133,N_19670);
nor U21093 (N_21093,N_19273,N_19661);
nand U21094 (N_21094,N_20118,N_20196);
nand U21095 (N_21095,N_20039,N_19818);
or U21096 (N_21096,N_19203,N_20272);
nor U21097 (N_21097,N_20319,N_20384);
xnor U21098 (N_21098,N_20170,N_19265);
nor U21099 (N_21099,N_19538,N_19276);
xnor U21100 (N_21100,N_20009,N_19314);
or U21101 (N_21101,N_20391,N_19783);
nand U21102 (N_21102,N_19311,N_19800);
and U21103 (N_21103,N_19302,N_19702);
nor U21104 (N_21104,N_19298,N_20297);
or U21105 (N_21105,N_19276,N_20177);
and U21106 (N_21106,N_19332,N_20012);
nor U21107 (N_21107,N_20119,N_20058);
or U21108 (N_21108,N_20312,N_19479);
and U21109 (N_21109,N_20007,N_20302);
xor U21110 (N_21110,N_20205,N_19961);
or U21111 (N_21111,N_20120,N_20210);
xnor U21112 (N_21112,N_19923,N_19532);
nand U21113 (N_21113,N_19501,N_19500);
xor U21114 (N_21114,N_19422,N_19603);
nand U21115 (N_21115,N_20087,N_19686);
xor U21116 (N_21116,N_19577,N_20222);
xor U21117 (N_21117,N_19865,N_20094);
nor U21118 (N_21118,N_20187,N_19713);
xnor U21119 (N_21119,N_19815,N_20275);
or U21120 (N_21120,N_19218,N_19324);
and U21121 (N_21121,N_19384,N_19818);
nand U21122 (N_21122,N_19326,N_19635);
and U21123 (N_21123,N_19870,N_19399);
or U21124 (N_21124,N_19244,N_19321);
or U21125 (N_21125,N_20256,N_19528);
and U21126 (N_21126,N_19616,N_20394);
nor U21127 (N_21127,N_19887,N_20056);
xor U21128 (N_21128,N_19424,N_19789);
or U21129 (N_21129,N_19803,N_19588);
xor U21130 (N_21130,N_19730,N_20374);
or U21131 (N_21131,N_19488,N_19865);
xor U21132 (N_21132,N_20140,N_19762);
xnor U21133 (N_21133,N_19533,N_20100);
nor U21134 (N_21134,N_20233,N_19534);
nor U21135 (N_21135,N_19464,N_19463);
and U21136 (N_21136,N_20045,N_19901);
and U21137 (N_21137,N_19830,N_19496);
nor U21138 (N_21138,N_19226,N_19840);
or U21139 (N_21139,N_19282,N_19220);
nand U21140 (N_21140,N_19246,N_19933);
and U21141 (N_21141,N_19791,N_20367);
xor U21142 (N_21142,N_19386,N_19470);
or U21143 (N_21143,N_20158,N_19601);
and U21144 (N_21144,N_19795,N_20059);
xor U21145 (N_21145,N_19738,N_19552);
or U21146 (N_21146,N_19629,N_19860);
and U21147 (N_21147,N_19503,N_19230);
xnor U21148 (N_21148,N_20301,N_20000);
or U21149 (N_21149,N_19403,N_19968);
nor U21150 (N_21150,N_19872,N_19746);
nor U21151 (N_21151,N_20023,N_20089);
nand U21152 (N_21152,N_19977,N_19236);
xnor U21153 (N_21153,N_19942,N_20162);
nand U21154 (N_21154,N_19828,N_19470);
xnor U21155 (N_21155,N_20213,N_19391);
nor U21156 (N_21156,N_19936,N_20360);
nor U21157 (N_21157,N_19722,N_19915);
nand U21158 (N_21158,N_20343,N_19617);
nand U21159 (N_21159,N_19306,N_19312);
and U21160 (N_21160,N_20346,N_19618);
nor U21161 (N_21161,N_19479,N_19311);
nor U21162 (N_21162,N_19244,N_20304);
nand U21163 (N_21163,N_20157,N_20243);
and U21164 (N_21164,N_19234,N_20136);
nor U21165 (N_21165,N_19612,N_20190);
and U21166 (N_21166,N_20387,N_20312);
or U21167 (N_21167,N_19477,N_19828);
nand U21168 (N_21168,N_19658,N_19956);
nand U21169 (N_21169,N_19612,N_20231);
and U21170 (N_21170,N_20389,N_19655);
or U21171 (N_21171,N_20342,N_20249);
xnor U21172 (N_21172,N_20232,N_19478);
and U21173 (N_21173,N_19565,N_19931);
nor U21174 (N_21174,N_19254,N_19699);
nand U21175 (N_21175,N_19969,N_19943);
nand U21176 (N_21176,N_19227,N_20374);
and U21177 (N_21177,N_19462,N_19274);
xor U21178 (N_21178,N_19864,N_20140);
or U21179 (N_21179,N_19834,N_19841);
or U21180 (N_21180,N_19365,N_20076);
nand U21181 (N_21181,N_20319,N_19210);
nor U21182 (N_21182,N_19390,N_19638);
nor U21183 (N_21183,N_20377,N_20157);
nor U21184 (N_21184,N_19982,N_19443);
nor U21185 (N_21185,N_19606,N_19329);
xnor U21186 (N_21186,N_19649,N_19304);
or U21187 (N_21187,N_19460,N_20147);
xnor U21188 (N_21188,N_19605,N_19481);
and U21189 (N_21189,N_20142,N_20272);
xnor U21190 (N_21190,N_19287,N_20126);
nand U21191 (N_21191,N_19902,N_19409);
and U21192 (N_21192,N_19900,N_19943);
or U21193 (N_21193,N_19616,N_20052);
nor U21194 (N_21194,N_19324,N_19279);
or U21195 (N_21195,N_19283,N_19628);
nor U21196 (N_21196,N_20010,N_19590);
and U21197 (N_21197,N_19260,N_20202);
and U21198 (N_21198,N_20100,N_20280);
nor U21199 (N_21199,N_19247,N_20319);
nand U21200 (N_21200,N_19544,N_19733);
xnor U21201 (N_21201,N_19926,N_19304);
xnor U21202 (N_21202,N_20259,N_20209);
nor U21203 (N_21203,N_20123,N_20084);
nand U21204 (N_21204,N_19910,N_19629);
and U21205 (N_21205,N_19205,N_19398);
xor U21206 (N_21206,N_19682,N_19249);
nand U21207 (N_21207,N_19444,N_20134);
nand U21208 (N_21208,N_19974,N_19850);
or U21209 (N_21209,N_19748,N_19761);
nor U21210 (N_21210,N_19754,N_20171);
or U21211 (N_21211,N_19821,N_19441);
and U21212 (N_21212,N_19580,N_19289);
and U21213 (N_21213,N_19480,N_20276);
and U21214 (N_21214,N_20391,N_20389);
xnor U21215 (N_21215,N_19931,N_19965);
and U21216 (N_21216,N_19572,N_20358);
and U21217 (N_21217,N_19888,N_19447);
nor U21218 (N_21218,N_19405,N_19773);
nor U21219 (N_21219,N_20197,N_19263);
and U21220 (N_21220,N_19370,N_19410);
nor U21221 (N_21221,N_20127,N_19216);
and U21222 (N_21222,N_20132,N_19318);
nand U21223 (N_21223,N_19912,N_19605);
nor U21224 (N_21224,N_20149,N_20316);
nand U21225 (N_21225,N_19361,N_19579);
xor U21226 (N_21226,N_20292,N_19528);
or U21227 (N_21227,N_19569,N_20216);
xnor U21228 (N_21228,N_20292,N_19325);
nand U21229 (N_21229,N_19554,N_19985);
nand U21230 (N_21230,N_20342,N_19453);
and U21231 (N_21231,N_19318,N_19568);
nor U21232 (N_21232,N_19593,N_19333);
xor U21233 (N_21233,N_19280,N_20339);
nand U21234 (N_21234,N_20057,N_19913);
nor U21235 (N_21235,N_19916,N_19918);
nor U21236 (N_21236,N_19615,N_19456);
and U21237 (N_21237,N_20133,N_20023);
nor U21238 (N_21238,N_20187,N_19690);
nor U21239 (N_21239,N_19401,N_20245);
or U21240 (N_21240,N_20166,N_20203);
and U21241 (N_21241,N_19309,N_19701);
nor U21242 (N_21242,N_19575,N_20328);
nor U21243 (N_21243,N_20253,N_19660);
or U21244 (N_21244,N_19750,N_20378);
and U21245 (N_21245,N_19703,N_19667);
nand U21246 (N_21246,N_20119,N_19450);
nand U21247 (N_21247,N_19660,N_19764);
and U21248 (N_21248,N_19329,N_19723);
nand U21249 (N_21249,N_20336,N_19899);
nand U21250 (N_21250,N_20332,N_19562);
nor U21251 (N_21251,N_19684,N_20102);
xnor U21252 (N_21252,N_19245,N_19705);
nand U21253 (N_21253,N_19711,N_19428);
nor U21254 (N_21254,N_19831,N_19588);
xnor U21255 (N_21255,N_20259,N_19433);
and U21256 (N_21256,N_19759,N_20393);
nand U21257 (N_21257,N_20071,N_19294);
nand U21258 (N_21258,N_20080,N_20281);
and U21259 (N_21259,N_19681,N_19990);
nor U21260 (N_21260,N_19233,N_19835);
nand U21261 (N_21261,N_20368,N_19911);
nand U21262 (N_21262,N_19752,N_19770);
xor U21263 (N_21263,N_19502,N_19739);
or U21264 (N_21264,N_19535,N_19603);
or U21265 (N_21265,N_19616,N_19766);
or U21266 (N_21266,N_20017,N_19579);
nand U21267 (N_21267,N_20065,N_19643);
and U21268 (N_21268,N_19891,N_20103);
and U21269 (N_21269,N_19561,N_19355);
and U21270 (N_21270,N_19664,N_19522);
nor U21271 (N_21271,N_19226,N_19338);
or U21272 (N_21272,N_20191,N_19896);
or U21273 (N_21273,N_19833,N_19548);
nand U21274 (N_21274,N_19705,N_20233);
xnor U21275 (N_21275,N_19421,N_19271);
or U21276 (N_21276,N_19407,N_19828);
nor U21277 (N_21277,N_19302,N_20043);
xor U21278 (N_21278,N_19376,N_20081);
xor U21279 (N_21279,N_19677,N_20111);
and U21280 (N_21280,N_19844,N_20090);
nand U21281 (N_21281,N_19340,N_19533);
and U21282 (N_21282,N_19947,N_20070);
nand U21283 (N_21283,N_20168,N_19720);
nand U21284 (N_21284,N_20386,N_19335);
or U21285 (N_21285,N_19610,N_20318);
or U21286 (N_21286,N_20280,N_19842);
xor U21287 (N_21287,N_19967,N_20010);
nand U21288 (N_21288,N_19758,N_19448);
nand U21289 (N_21289,N_20074,N_20172);
nor U21290 (N_21290,N_20286,N_20172);
nor U21291 (N_21291,N_19657,N_20014);
or U21292 (N_21292,N_19366,N_19462);
or U21293 (N_21293,N_19575,N_20188);
nand U21294 (N_21294,N_19253,N_19642);
nor U21295 (N_21295,N_19872,N_19848);
nand U21296 (N_21296,N_19882,N_19843);
nor U21297 (N_21297,N_19455,N_19350);
and U21298 (N_21298,N_19970,N_20124);
nor U21299 (N_21299,N_19793,N_19917);
nand U21300 (N_21300,N_19451,N_20379);
or U21301 (N_21301,N_20281,N_19648);
nor U21302 (N_21302,N_19652,N_20178);
xor U21303 (N_21303,N_19516,N_19382);
and U21304 (N_21304,N_19495,N_19891);
and U21305 (N_21305,N_20281,N_19547);
and U21306 (N_21306,N_20367,N_19949);
xnor U21307 (N_21307,N_19276,N_19930);
nor U21308 (N_21308,N_20255,N_19810);
and U21309 (N_21309,N_20032,N_19557);
or U21310 (N_21310,N_19423,N_19513);
nor U21311 (N_21311,N_19228,N_20324);
and U21312 (N_21312,N_19521,N_19323);
nand U21313 (N_21313,N_20329,N_19729);
or U21314 (N_21314,N_19590,N_19238);
or U21315 (N_21315,N_19714,N_20331);
or U21316 (N_21316,N_20088,N_19706);
nand U21317 (N_21317,N_19759,N_19707);
and U21318 (N_21318,N_19376,N_20097);
nor U21319 (N_21319,N_20136,N_19661);
xnor U21320 (N_21320,N_20361,N_19870);
or U21321 (N_21321,N_20229,N_20230);
nand U21322 (N_21322,N_20280,N_20166);
or U21323 (N_21323,N_20004,N_19694);
or U21324 (N_21324,N_20152,N_19297);
and U21325 (N_21325,N_19277,N_20203);
and U21326 (N_21326,N_19773,N_19410);
xnor U21327 (N_21327,N_19445,N_19203);
xnor U21328 (N_21328,N_19980,N_19828);
xnor U21329 (N_21329,N_20024,N_19273);
or U21330 (N_21330,N_19986,N_20354);
or U21331 (N_21331,N_19456,N_20286);
and U21332 (N_21332,N_20019,N_19264);
nor U21333 (N_21333,N_20200,N_19802);
nand U21334 (N_21334,N_20237,N_19997);
and U21335 (N_21335,N_19426,N_19682);
and U21336 (N_21336,N_20252,N_19852);
and U21337 (N_21337,N_19332,N_19788);
nor U21338 (N_21338,N_19518,N_19535);
or U21339 (N_21339,N_19680,N_19273);
or U21340 (N_21340,N_19542,N_20128);
xnor U21341 (N_21341,N_19507,N_19466);
nor U21342 (N_21342,N_19220,N_20255);
xor U21343 (N_21343,N_19988,N_19658);
or U21344 (N_21344,N_19573,N_19358);
nor U21345 (N_21345,N_19424,N_19543);
xnor U21346 (N_21346,N_19523,N_20068);
nand U21347 (N_21347,N_20034,N_19994);
or U21348 (N_21348,N_19293,N_20354);
and U21349 (N_21349,N_19354,N_20339);
or U21350 (N_21350,N_19406,N_19864);
nand U21351 (N_21351,N_19910,N_19592);
or U21352 (N_21352,N_19749,N_19223);
xor U21353 (N_21353,N_19601,N_19523);
or U21354 (N_21354,N_20132,N_19325);
xnor U21355 (N_21355,N_20144,N_19254);
nor U21356 (N_21356,N_20197,N_20364);
or U21357 (N_21357,N_19848,N_19685);
and U21358 (N_21358,N_20289,N_20140);
xnor U21359 (N_21359,N_19549,N_19355);
xor U21360 (N_21360,N_19780,N_19344);
xor U21361 (N_21361,N_19223,N_19872);
and U21362 (N_21362,N_19440,N_20192);
and U21363 (N_21363,N_19579,N_19769);
nand U21364 (N_21364,N_19330,N_19969);
nand U21365 (N_21365,N_19985,N_19293);
and U21366 (N_21366,N_20129,N_20393);
xor U21367 (N_21367,N_19943,N_19248);
xnor U21368 (N_21368,N_19684,N_19727);
nand U21369 (N_21369,N_20334,N_20326);
nand U21370 (N_21370,N_19789,N_19250);
nor U21371 (N_21371,N_19919,N_19421);
nand U21372 (N_21372,N_19975,N_20203);
and U21373 (N_21373,N_19335,N_19344);
and U21374 (N_21374,N_19631,N_19316);
and U21375 (N_21375,N_19625,N_19320);
or U21376 (N_21376,N_19440,N_19901);
nand U21377 (N_21377,N_19323,N_20160);
or U21378 (N_21378,N_20333,N_19334);
or U21379 (N_21379,N_20206,N_19344);
xor U21380 (N_21380,N_19303,N_19896);
and U21381 (N_21381,N_19253,N_19243);
nand U21382 (N_21382,N_20214,N_20019);
nor U21383 (N_21383,N_19570,N_19434);
xor U21384 (N_21384,N_19538,N_20296);
or U21385 (N_21385,N_19735,N_19850);
or U21386 (N_21386,N_19706,N_20287);
xnor U21387 (N_21387,N_20149,N_19289);
and U21388 (N_21388,N_19272,N_19660);
nor U21389 (N_21389,N_19652,N_19773);
nor U21390 (N_21390,N_19637,N_20353);
and U21391 (N_21391,N_20055,N_19959);
nor U21392 (N_21392,N_19476,N_20287);
xnor U21393 (N_21393,N_19764,N_19763);
nand U21394 (N_21394,N_19554,N_20364);
nand U21395 (N_21395,N_19594,N_19501);
and U21396 (N_21396,N_19279,N_20114);
and U21397 (N_21397,N_20214,N_20279);
nand U21398 (N_21398,N_20347,N_20225);
nor U21399 (N_21399,N_19889,N_19982);
and U21400 (N_21400,N_19605,N_20007);
and U21401 (N_21401,N_19802,N_19848);
nor U21402 (N_21402,N_19385,N_20282);
nor U21403 (N_21403,N_19588,N_19300);
nand U21404 (N_21404,N_19556,N_19442);
and U21405 (N_21405,N_19717,N_19936);
nand U21406 (N_21406,N_19675,N_20124);
nand U21407 (N_21407,N_19747,N_20387);
nor U21408 (N_21408,N_20103,N_20192);
nand U21409 (N_21409,N_19608,N_19909);
nor U21410 (N_21410,N_19826,N_20368);
xnor U21411 (N_21411,N_19476,N_20121);
nor U21412 (N_21412,N_20233,N_19465);
or U21413 (N_21413,N_20078,N_19555);
nor U21414 (N_21414,N_19439,N_19691);
nor U21415 (N_21415,N_19861,N_20263);
xor U21416 (N_21416,N_19968,N_20001);
nand U21417 (N_21417,N_19791,N_19845);
and U21418 (N_21418,N_20298,N_19824);
nor U21419 (N_21419,N_19945,N_20320);
or U21420 (N_21420,N_19622,N_19883);
or U21421 (N_21421,N_20143,N_19835);
nor U21422 (N_21422,N_19342,N_19452);
nor U21423 (N_21423,N_19667,N_19384);
and U21424 (N_21424,N_19337,N_20002);
and U21425 (N_21425,N_19836,N_19531);
and U21426 (N_21426,N_19411,N_19992);
xnor U21427 (N_21427,N_19379,N_19223);
nand U21428 (N_21428,N_20204,N_20201);
or U21429 (N_21429,N_20366,N_19356);
and U21430 (N_21430,N_20140,N_19271);
nor U21431 (N_21431,N_20031,N_20152);
or U21432 (N_21432,N_19754,N_20341);
xor U21433 (N_21433,N_19898,N_19603);
nand U21434 (N_21434,N_19367,N_19970);
xor U21435 (N_21435,N_20114,N_19757);
or U21436 (N_21436,N_20369,N_19839);
or U21437 (N_21437,N_20117,N_19761);
and U21438 (N_21438,N_20373,N_19802);
xnor U21439 (N_21439,N_19291,N_20353);
nor U21440 (N_21440,N_19988,N_20310);
nor U21441 (N_21441,N_19980,N_19536);
nand U21442 (N_21442,N_20275,N_20025);
xor U21443 (N_21443,N_19453,N_19446);
or U21444 (N_21444,N_19503,N_20340);
or U21445 (N_21445,N_19458,N_19483);
and U21446 (N_21446,N_19610,N_19777);
and U21447 (N_21447,N_19215,N_19745);
nor U21448 (N_21448,N_19748,N_19723);
and U21449 (N_21449,N_19660,N_19389);
xnor U21450 (N_21450,N_19612,N_19821);
nor U21451 (N_21451,N_19583,N_19446);
nand U21452 (N_21452,N_19887,N_19908);
and U21453 (N_21453,N_20183,N_19618);
and U21454 (N_21454,N_19963,N_19735);
and U21455 (N_21455,N_20208,N_19228);
and U21456 (N_21456,N_19647,N_19314);
xor U21457 (N_21457,N_19237,N_20242);
xnor U21458 (N_21458,N_19836,N_19866);
or U21459 (N_21459,N_19589,N_19638);
nand U21460 (N_21460,N_19934,N_19352);
or U21461 (N_21461,N_19317,N_19235);
or U21462 (N_21462,N_20008,N_19351);
nor U21463 (N_21463,N_19650,N_19843);
and U21464 (N_21464,N_19842,N_19636);
nor U21465 (N_21465,N_19663,N_19965);
xnor U21466 (N_21466,N_19475,N_19855);
xor U21467 (N_21467,N_20184,N_19692);
nand U21468 (N_21468,N_19910,N_20335);
and U21469 (N_21469,N_19700,N_20357);
xnor U21470 (N_21470,N_19424,N_20165);
and U21471 (N_21471,N_20332,N_19263);
nor U21472 (N_21472,N_19296,N_20130);
xnor U21473 (N_21473,N_19791,N_20195);
and U21474 (N_21474,N_19204,N_19543);
or U21475 (N_21475,N_20212,N_19221);
or U21476 (N_21476,N_20112,N_20017);
or U21477 (N_21477,N_20276,N_20287);
or U21478 (N_21478,N_19310,N_19283);
nor U21479 (N_21479,N_19848,N_19956);
and U21480 (N_21480,N_19514,N_19862);
xnor U21481 (N_21481,N_19407,N_19231);
nor U21482 (N_21482,N_19644,N_19446);
nand U21483 (N_21483,N_19262,N_19517);
xnor U21484 (N_21484,N_19398,N_20031);
nor U21485 (N_21485,N_19261,N_20361);
nand U21486 (N_21486,N_20011,N_20253);
and U21487 (N_21487,N_19783,N_19743);
and U21488 (N_21488,N_19631,N_19333);
or U21489 (N_21489,N_19596,N_19303);
and U21490 (N_21490,N_20135,N_20358);
nor U21491 (N_21491,N_20258,N_19623);
xor U21492 (N_21492,N_20156,N_19650);
and U21493 (N_21493,N_19307,N_20119);
xnor U21494 (N_21494,N_19393,N_19398);
and U21495 (N_21495,N_20223,N_20004);
or U21496 (N_21496,N_19371,N_20045);
xnor U21497 (N_21497,N_19977,N_19495);
or U21498 (N_21498,N_19228,N_19855);
nor U21499 (N_21499,N_19366,N_19403);
and U21500 (N_21500,N_19521,N_19329);
xnor U21501 (N_21501,N_19721,N_20314);
xnor U21502 (N_21502,N_20292,N_19732);
and U21503 (N_21503,N_20220,N_19969);
and U21504 (N_21504,N_19476,N_19265);
nor U21505 (N_21505,N_20321,N_19887);
nor U21506 (N_21506,N_19898,N_19605);
or U21507 (N_21507,N_19627,N_19536);
nor U21508 (N_21508,N_19288,N_20191);
nand U21509 (N_21509,N_19547,N_20050);
xnor U21510 (N_21510,N_20210,N_19337);
or U21511 (N_21511,N_20161,N_20268);
and U21512 (N_21512,N_19951,N_20135);
and U21513 (N_21513,N_19382,N_19770);
and U21514 (N_21514,N_19924,N_20200);
nor U21515 (N_21515,N_19798,N_19837);
and U21516 (N_21516,N_20325,N_19200);
and U21517 (N_21517,N_19248,N_19546);
and U21518 (N_21518,N_19864,N_19330);
nand U21519 (N_21519,N_19741,N_19326);
xnor U21520 (N_21520,N_19282,N_19543);
or U21521 (N_21521,N_19578,N_19720);
xnor U21522 (N_21522,N_19583,N_19523);
nor U21523 (N_21523,N_19897,N_19934);
or U21524 (N_21524,N_19332,N_19543);
xor U21525 (N_21525,N_19284,N_20259);
xnor U21526 (N_21526,N_19480,N_20113);
and U21527 (N_21527,N_19645,N_20026);
nor U21528 (N_21528,N_20327,N_19752);
nor U21529 (N_21529,N_19643,N_20218);
xor U21530 (N_21530,N_19801,N_20282);
and U21531 (N_21531,N_20153,N_20251);
nand U21532 (N_21532,N_19518,N_20021);
and U21533 (N_21533,N_20366,N_19747);
nor U21534 (N_21534,N_19973,N_20063);
or U21535 (N_21535,N_19814,N_19616);
and U21536 (N_21536,N_20203,N_19813);
or U21537 (N_21537,N_20363,N_19482);
nand U21538 (N_21538,N_19435,N_20215);
xor U21539 (N_21539,N_20232,N_19345);
or U21540 (N_21540,N_19851,N_20080);
nor U21541 (N_21541,N_20123,N_19660);
nor U21542 (N_21542,N_19647,N_20348);
or U21543 (N_21543,N_19857,N_19611);
or U21544 (N_21544,N_19430,N_19925);
xnor U21545 (N_21545,N_19659,N_20056);
or U21546 (N_21546,N_19630,N_20051);
nand U21547 (N_21547,N_20212,N_20361);
and U21548 (N_21548,N_19224,N_19347);
nor U21549 (N_21549,N_19989,N_19945);
nand U21550 (N_21550,N_20060,N_20285);
nand U21551 (N_21551,N_19358,N_19853);
xor U21552 (N_21552,N_19384,N_19480);
nor U21553 (N_21553,N_19633,N_19333);
or U21554 (N_21554,N_20302,N_19894);
or U21555 (N_21555,N_19598,N_19798);
nor U21556 (N_21556,N_19256,N_20370);
nor U21557 (N_21557,N_20093,N_19870);
or U21558 (N_21558,N_19236,N_19599);
and U21559 (N_21559,N_19455,N_19666);
nor U21560 (N_21560,N_19592,N_19648);
and U21561 (N_21561,N_20164,N_20090);
or U21562 (N_21562,N_20132,N_19705);
xor U21563 (N_21563,N_19658,N_19777);
nand U21564 (N_21564,N_19295,N_20060);
nor U21565 (N_21565,N_20050,N_19232);
and U21566 (N_21566,N_20229,N_19525);
or U21567 (N_21567,N_19547,N_19736);
nand U21568 (N_21568,N_19625,N_20302);
nand U21569 (N_21569,N_19219,N_20301);
or U21570 (N_21570,N_19538,N_19909);
and U21571 (N_21571,N_20095,N_19643);
or U21572 (N_21572,N_20326,N_20188);
xnor U21573 (N_21573,N_19832,N_19535);
or U21574 (N_21574,N_19914,N_19301);
or U21575 (N_21575,N_19804,N_19279);
and U21576 (N_21576,N_20153,N_20112);
or U21577 (N_21577,N_20145,N_19523);
xnor U21578 (N_21578,N_19991,N_19810);
nor U21579 (N_21579,N_19947,N_19703);
nand U21580 (N_21580,N_19929,N_19258);
xnor U21581 (N_21581,N_19777,N_19926);
and U21582 (N_21582,N_19519,N_20153);
and U21583 (N_21583,N_20278,N_19614);
nor U21584 (N_21584,N_19836,N_20163);
nor U21585 (N_21585,N_19972,N_19905);
or U21586 (N_21586,N_19889,N_19200);
and U21587 (N_21587,N_19491,N_19272);
and U21588 (N_21588,N_19616,N_19890);
xor U21589 (N_21589,N_19300,N_19255);
or U21590 (N_21590,N_19395,N_19615);
nor U21591 (N_21591,N_20178,N_20284);
or U21592 (N_21592,N_19791,N_19764);
xor U21593 (N_21593,N_19643,N_20388);
or U21594 (N_21594,N_19755,N_20236);
or U21595 (N_21595,N_19776,N_19720);
or U21596 (N_21596,N_20191,N_19376);
or U21597 (N_21597,N_19660,N_20147);
xor U21598 (N_21598,N_19530,N_19989);
and U21599 (N_21599,N_19582,N_19920);
or U21600 (N_21600,N_21103,N_21115);
xor U21601 (N_21601,N_21205,N_21116);
or U21602 (N_21602,N_21289,N_21000);
nand U21603 (N_21603,N_20704,N_21068);
and U21604 (N_21604,N_20868,N_20424);
nand U21605 (N_21605,N_20827,N_20713);
nor U21606 (N_21606,N_20811,N_21572);
nor U21607 (N_21607,N_21301,N_21251);
nor U21608 (N_21608,N_21361,N_20779);
or U21609 (N_21609,N_20419,N_20563);
or U21610 (N_21610,N_20491,N_20621);
or U21611 (N_21611,N_20833,N_20897);
nor U21612 (N_21612,N_21408,N_20520);
nand U21613 (N_21613,N_20524,N_21333);
and U21614 (N_21614,N_21345,N_20528);
xnor U21615 (N_21615,N_21481,N_20461);
xnor U21616 (N_21616,N_21536,N_20987);
nand U21617 (N_21617,N_21311,N_20402);
nand U21618 (N_21618,N_21001,N_21538);
nor U21619 (N_21619,N_21526,N_20644);
nand U21620 (N_21620,N_21318,N_20872);
nor U21621 (N_21621,N_20942,N_20706);
or U21622 (N_21622,N_21034,N_21183);
and U21623 (N_21623,N_20645,N_21101);
nor U21624 (N_21624,N_20648,N_20663);
xnor U21625 (N_21625,N_21144,N_20913);
nor U21626 (N_21626,N_21139,N_21217);
and U21627 (N_21627,N_21201,N_20581);
and U21628 (N_21628,N_20457,N_21121);
or U21629 (N_21629,N_20616,N_21582);
nand U21630 (N_21630,N_20416,N_20626);
nand U21631 (N_21631,N_20599,N_21310);
and U21632 (N_21632,N_21079,N_21543);
xor U21633 (N_21633,N_20852,N_20583);
xnor U21634 (N_21634,N_21184,N_20697);
nand U21635 (N_21635,N_20537,N_21218);
xnor U21636 (N_21636,N_21281,N_20800);
nor U21637 (N_21637,N_20536,N_21287);
xor U21638 (N_21638,N_20511,N_21192);
nand U21639 (N_21639,N_21241,N_20986);
nand U21640 (N_21640,N_20669,N_20726);
xor U21641 (N_21641,N_20525,N_21261);
nor U21642 (N_21642,N_20611,N_21562);
and U21643 (N_21643,N_21260,N_20518);
xnor U21644 (N_21644,N_21203,N_21323);
nor U21645 (N_21645,N_21568,N_20501);
nor U21646 (N_21646,N_21188,N_20530);
and U21647 (N_21647,N_21457,N_20935);
nor U21648 (N_21648,N_20571,N_20427);
or U21649 (N_21649,N_20719,N_20998);
or U21650 (N_21650,N_21257,N_21247);
nor U21651 (N_21651,N_20956,N_21433);
xor U21652 (N_21652,N_21441,N_21550);
xor U21653 (N_21653,N_21012,N_20995);
and U21654 (N_21654,N_21211,N_21024);
xor U21655 (N_21655,N_20907,N_20957);
nand U21656 (N_21656,N_21169,N_20658);
and U21657 (N_21657,N_21010,N_21038);
nor U21658 (N_21658,N_20912,N_20679);
xor U21659 (N_21659,N_21208,N_21475);
nor U21660 (N_21660,N_21443,N_21422);
nand U21661 (N_21661,N_21372,N_20553);
nand U21662 (N_21662,N_21586,N_20932);
xnor U21663 (N_21663,N_20686,N_20734);
or U21664 (N_21664,N_21109,N_21271);
nor U21665 (N_21665,N_21132,N_21041);
or U21666 (N_21666,N_21339,N_20947);
nand U21667 (N_21667,N_20438,N_21331);
or U21668 (N_21668,N_21053,N_20632);
xor U21669 (N_21669,N_21233,N_21541);
or U21670 (N_21670,N_21084,N_20463);
or U21671 (N_21671,N_20432,N_21356);
nor U21672 (N_21672,N_20573,N_20839);
or U21673 (N_21673,N_21319,N_21357);
nand U21674 (N_21674,N_21086,N_21014);
xnor U21675 (N_21675,N_21039,N_21031);
nand U21676 (N_21676,N_21246,N_20634);
nor U21677 (N_21677,N_21009,N_21344);
nor U21678 (N_21678,N_21314,N_20735);
xnor U21679 (N_21679,N_21081,N_20768);
nor U21680 (N_21680,N_20748,N_21137);
and U21681 (N_21681,N_20561,N_21486);
nor U21682 (N_21682,N_20879,N_21047);
and U21683 (N_21683,N_20804,N_20542);
nor U21684 (N_21684,N_20950,N_20816);
nand U21685 (N_21685,N_20642,N_20417);
xnor U21686 (N_21686,N_21142,N_20989);
xor U21687 (N_21687,N_20934,N_21178);
and U21688 (N_21688,N_21367,N_21552);
nor U21689 (N_21689,N_20628,N_20666);
or U21690 (N_21690,N_21267,N_20836);
xor U21691 (N_21691,N_20850,N_21430);
nor U21692 (N_21692,N_20535,N_21396);
nor U21693 (N_21693,N_21173,N_21273);
or U21694 (N_21694,N_20578,N_20488);
or U21695 (N_21695,N_21565,N_20436);
nand U21696 (N_21696,N_20963,N_20776);
or U21697 (N_21697,N_21368,N_20494);
nor U21698 (N_21698,N_21412,N_21063);
and U21699 (N_21699,N_21378,N_21557);
and U21700 (N_21700,N_20588,N_20778);
and U21701 (N_21701,N_20649,N_20899);
nand U21702 (N_21702,N_21497,N_21005);
xor U21703 (N_21703,N_20925,N_20869);
and U21704 (N_21704,N_21406,N_21397);
nor U21705 (N_21705,N_20717,N_20595);
and U21706 (N_21706,N_21573,N_21500);
nor U21707 (N_21707,N_21228,N_20741);
xor U21708 (N_21708,N_21199,N_21463);
nor U21709 (N_21709,N_20862,N_21119);
or U21710 (N_21710,N_21167,N_20499);
xor U21711 (N_21711,N_21566,N_20490);
nor U21712 (N_21712,N_21265,N_20887);
and U21713 (N_21713,N_21437,N_21304);
xor U21714 (N_21714,N_20538,N_20677);
nor U21715 (N_21715,N_20452,N_21065);
nand U21716 (N_21716,N_20540,N_20609);
and U21717 (N_21717,N_20478,N_20780);
xnor U21718 (N_21718,N_21567,N_21332);
nand U21719 (N_21719,N_20900,N_21384);
and U21720 (N_21720,N_20691,N_21484);
and U21721 (N_21721,N_20858,N_21035);
nand U21722 (N_21722,N_21591,N_20916);
and U21723 (N_21723,N_20714,N_20492);
or U21724 (N_21724,N_20921,N_20973);
or U21725 (N_21725,N_21590,N_20982);
nand U21726 (N_21726,N_21448,N_20637);
xnor U21727 (N_21727,N_21170,N_20939);
and U21728 (N_21728,N_20560,N_21298);
or U21729 (N_21729,N_20830,N_20514);
or U21730 (N_21730,N_21099,N_21232);
and U21731 (N_21731,N_20455,N_20926);
nor U21732 (N_21732,N_21403,N_21229);
nor U21733 (N_21733,N_21411,N_21596);
and U21734 (N_21734,N_20617,N_21542);
or U21735 (N_21735,N_20829,N_21470);
or U21736 (N_21736,N_21425,N_21055);
xor U21737 (N_21737,N_20716,N_21337);
and U21738 (N_21738,N_20664,N_20674);
and U21739 (N_21739,N_20922,N_21512);
nand U21740 (N_21740,N_21460,N_21242);
nand U21741 (N_21741,N_20889,N_21046);
and U21742 (N_21742,N_20624,N_20911);
nand U21743 (N_21743,N_21306,N_20856);
nor U21744 (N_21744,N_21392,N_20974);
or U21745 (N_21745,N_21126,N_21577);
or U21746 (N_21746,N_20978,N_21230);
nand U21747 (N_21747,N_20454,N_21371);
xor U21748 (N_21748,N_21327,N_21299);
and U21749 (N_21749,N_21108,N_21118);
nor U21750 (N_21750,N_20646,N_20808);
nand U21751 (N_21751,N_20786,N_20610);
xnor U21752 (N_21752,N_20760,N_20906);
or U21753 (N_21753,N_20834,N_21186);
or U21754 (N_21754,N_21315,N_20638);
nor U21755 (N_21755,N_20656,N_20742);
nor U21756 (N_21756,N_20782,N_20472);
or U21757 (N_21757,N_20587,N_21467);
nor U21758 (N_21758,N_20791,N_20444);
xor U21759 (N_21759,N_21428,N_21426);
nor U21760 (N_21760,N_20813,N_21025);
nand U21761 (N_21761,N_20841,N_21349);
xor U21762 (N_21762,N_20979,N_21581);
nor U21763 (N_21763,N_20548,N_21405);
nand U21764 (N_21764,N_20812,N_20866);
nor U21765 (N_21765,N_21151,N_21452);
and U21766 (N_21766,N_21593,N_21070);
and U21767 (N_21767,N_21364,N_21131);
nor U21768 (N_21768,N_21098,N_21454);
or U21769 (N_21769,N_20722,N_21283);
and U21770 (N_21770,N_20489,N_20751);
nor U21771 (N_21771,N_21442,N_20411);
xor U21772 (N_21772,N_20967,N_21363);
and U21773 (N_21773,N_20765,N_20640);
nand U21774 (N_21774,N_21177,N_20882);
and U21775 (N_21775,N_20559,N_20789);
nand U21776 (N_21776,N_21381,N_21309);
nor U21777 (N_21777,N_20908,N_21006);
and U21778 (N_21778,N_20737,N_21439);
and U21779 (N_21779,N_21374,N_21166);
nor U21780 (N_21780,N_21588,N_20665);
xnor U21781 (N_21781,N_21506,N_20904);
xnor U21782 (N_21782,N_20802,N_20855);
nor U21783 (N_21783,N_20429,N_20689);
xnor U21784 (N_21784,N_20917,N_21517);
and U21785 (N_21785,N_20988,N_20509);
or U21786 (N_21786,N_20754,N_21539);
xnor U21787 (N_21787,N_20826,N_20614);
xor U21788 (N_21788,N_21200,N_21540);
xnor U21789 (N_21789,N_20678,N_21589);
nand U21790 (N_21790,N_20915,N_21561);
nand U21791 (N_21791,N_21424,N_21061);
nor U21792 (N_21792,N_21158,N_20730);
xor U21793 (N_21793,N_20959,N_20985);
nand U21794 (N_21794,N_21227,N_20774);
or U21795 (N_21795,N_20651,N_20875);
nand U21796 (N_21796,N_21165,N_20512);
or U21797 (N_21797,N_21082,N_20671);
or U21798 (N_21798,N_21110,N_21197);
xor U21799 (N_21799,N_21136,N_20447);
or U21800 (N_21800,N_20857,N_20724);
and U21801 (N_21801,N_21148,N_20712);
xor U21802 (N_21802,N_21163,N_20589);
nor U21803 (N_21803,N_21052,N_21168);
xnor U21804 (N_21804,N_20828,N_21069);
or U21805 (N_21805,N_20552,N_20619);
and U21806 (N_21806,N_21076,N_21495);
nand U21807 (N_21807,N_21248,N_21569);
nor U21808 (N_21808,N_20728,N_21093);
nand U21809 (N_21809,N_20739,N_20568);
nor U21810 (N_21810,N_20814,N_21049);
xor U21811 (N_21811,N_20604,N_20948);
nand U21812 (N_21812,N_20961,N_20924);
nand U21813 (N_21813,N_20688,N_21545);
and U21814 (N_21814,N_21348,N_21546);
or U21815 (N_21815,N_21390,N_21033);
and U21816 (N_21816,N_20675,N_21483);
or U21817 (N_21817,N_20435,N_21421);
and U21818 (N_21818,N_20562,N_20980);
and U21819 (N_21819,N_20662,N_20708);
or U21820 (N_21820,N_20955,N_20733);
or U21821 (N_21821,N_20867,N_21342);
nand U21822 (N_21822,N_20580,N_20937);
xor U21823 (N_21823,N_20820,N_21202);
xnor U21824 (N_21824,N_21402,N_20554);
xor U21825 (N_21825,N_20418,N_21284);
and U21826 (N_21826,N_20977,N_21334);
xor U21827 (N_21827,N_21236,N_21353);
xor U21828 (N_21828,N_21525,N_21105);
xnor U21829 (N_21829,N_21471,N_20483);
or U21830 (N_21830,N_20895,N_20607);
nand U21831 (N_21831,N_20756,N_21491);
nand U21832 (N_21832,N_20414,N_20613);
nor U21833 (N_21833,N_21316,N_20458);
xnor U21834 (N_21834,N_21180,N_20936);
or U21835 (N_21835,N_20749,N_20783);
and U21836 (N_21836,N_20631,N_21007);
xnor U21837 (N_21837,N_21003,N_21329);
nor U21838 (N_21838,N_20612,N_21285);
or U21839 (N_21839,N_21280,N_21535);
nor U21840 (N_21840,N_21191,N_21223);
nor U21841 (N_21841,N_21585,N_20451);
and U21842 (N_21842,N_21258,N_21355);
or U21843 (N_21843,N_21420,N_21027);
or U21844 (N_21844,N_20764,N_21290);
and U21845 (N_21845,N_20927,N_21240);
xor U21846 (N_21846,N_21016,N_21094);
or U21847 (N_21847,N_20844,N_21578);
and U21848 (N_21848,N_21431,N_20598);
nand U21849 (N_21849,N_21048,N_21359);
nor U21850 (N_21850,N_20532,N_20625);
and U21851 (N_21851,N_20539,N_21185);
nor U21852 (N_21852,N_20550,N_20943);
xnor U21853 (N_21853,N_20482,N_21020);
nand U21854 (N_21854,N_21338,N_21485);
nor U21855 (N_21855,N_21449,N_21296);
nor U21856 (N_21856,N_21134,N_21307);
nand U21857 (N_21857,N_21369,N_20840);
and U21858 (N_21858,N_20496,N_20725);
nand U21859 (N_21859,N_20817,N_21564);
nor U21860 (N_21860,N_20443,N_21040);
xor U21861 (N_21861,N_21274,N_21328);
or U21862 (N_21862,N_20672,N_21499);
nor U21863 (N_21863,N_21073,N_20744);
nor U21864 (N_21864,N_21106,N_21436);
xnor U21865 (N_21865,N_21554,N_20430);
or U21866 (N_21866,N_20605,N_21250);
and U21867 (N_21867,N_20676,N_21135);
xnor U21868 (N_21868,N_21571,N_21407);
or U21869 (N_21869,N_20711,N_20775);
xor U21870 (N_21870,N_21075,N_21256);
nor U21871 (N_21871,N_20464,N_21510);
or U21872 (N_21872,N_21152,N_21059);
and U21873 (N_21873,N_21266,N_20412);
xor U21874 (N_21874,N_21330,N_21089);
nand U21875 (N_21875,N_21087,N_21019);
or U21876 (N_21876,N_20896,N_21350);
xnor U21877 (N_21877,N_21130,N_21351);
nand U21878 (N_21878,N_20682,N_21255);
xnor U21879 (N_21879,N_20873,N_21523);
or U21880 (N_21880,N_20515,N_21210);
and U21881 (N_21881,N_20700,N_21204);
xnor U21882 (N_21882,N_21514,N_21558);
xnor U21883 (N_21883,N_21474,N_20401);
nand U21884 (N_21884,N_21107,N_20792);
nor U21885 (N_21885,N_21294,N_20715);
nor U21886 (N_21886,N_21389,N_20738);
or U21887 (N_21887,N_20544,N_20584);
or U21888 (N_21888,N_20832,N_21574);
xnor U21889 (N_21889,N_21291,N_21122);
nor U21890 (N_21890,N_21502,N_20481);
and U21891 (N_21891,N_21221,N_21231);
xor U21892 (N_21892,N_20954,N_21164);
and U21893 (N_21893,N_20745,N_20630);
nor U21894 (N_21894,N_20972,N_20766);
nor U21895 (N_21895,N_20647,N_21219);
and U21896 (N_21896,N_21358,N_20822);
xnor U21897 (N_21897,N_21462,N_21160);
nor U21898 (N_21898,N_21595,N_21279);
or U21899 (N_21899,N_21370,N_21417);
or U21900 (N_21900,N_21579,N_21043);
nand U21901 (N_21901,N_20701,N_20403);
nor U21902 (N_21902,N_21117,N_20968);
and U21903 (N_21903,N_20788,N_20976);
and U21904 (N_21904,N_20400,N_21215);
and U21905 (N_21905,N_21584,N_20831);
xor U21906 (N_21906,N_21277,N_20591);
nand U21907 (N_21907,N_20854,N_20422);
nand U21908 (N_21908,N_21324,N_20890);
nand U21909 (N_21909,N_21592,N_20650);
and U21910 (N_21910,N_20949,N_21551);
and U21911 (N_21911,N_21128,N_21465);
nor U21912 (N_21912,N_20723,N_21057);
xor U21913 (N_21913,N_20838,N_21516);
or U21914 (N_21914,N_20504,N_20752);
and U21915 (N_21915,N_21434,N_21322);
and U21916 (N_21916,N_20860,N_21037);
or U21917 (N_21917,N_21341,N_21147);
nor U21918 (N_21918,N_21295,N_20473);
nor U21919 (N_21919,N_20885,N_20870);
or U21920 (N_21920,N_20582,N_21404);
nand U21921 (N_21921,N_20761,N_20522);
xnor U21922 (N_21922,N_21066,N_21383);
nand U21923 (N_21923,N_20781,N_20657);
xor U21924 (N_21924,N_21129,N_20874);
nor U21925 (N_21925,N_20667,N_21013);
and U21926 (N_21926,N_21455,N_20696);
or U21927 (N_21927,N_20886,N_20958);
and U21928 (N_21928,N_20593,N_20707);
and U21929 (N_21929,N_21138,N_21575);
and U21930 (N_21930,N_21161,N_20865);
nor U21931 (N_21931,N_20953,N_21174);
xor U21932 (N_21932,N_20894,N_20495);
xnor U21933 (N_21933,N_21028,N_21320);
xor U21934 (N_21934,N_20633,N_21021);
nor U21935 (N_21935,N_21493,N_21453);
xnor U21936 (N_21936,N_20805,N_21120);
nand U21937 (N_21937,N_20431,N_21023);
and U21938 (N_21938,N_21401,N_20549);
xnor U21939 (N_21939,N_21212,N_21599);
nor U21940 (N_21940,N_21456,N_21149);
or U21941 (N_21941,N_21088,N_21159);
xnor U21942 (N_21942,N_21410,N_21469);
xor U21943 (N_21943,N_21095,N_21143);
xnor U21944 (N_21944,N_20847,N_21529);
or U21945 (N_21945,N_21518,N_21022);
or U21946 (N_21946,N_21102,N_21409);
or U21947 (N_21947,N_20423,N_21459);
or U21948 (N_21948,N_21501,N_21056);
and U21949 (N_21949,N_21140,N_21388);
xor U21950 (N_21950,N_20966,N_20433);
nand U21951 (N_21951,N_20533,N_20566);
xnor U21952 (N_21952,N_21216,N_20997);
or U21953 (N_21953,N_21297,N_21553);
and U21954 (N_21954,N_20661,N_20919);
nor U21955 (N_21955,N_20462,N_20600);
or U21956 (N_21956,N_20803,N_20846);
or U21957 (N_21957,N_21293,N_20910);
and U21958 (N_21958,N_20821,N_21393);
nor U21959 (N_21959,N_20500,N_20547);
xnor U21960 (N_21960,N_21097,N_21435);
and U21961 (N_21961,N_20601,N_20545);
xnor U21962 (N_21962,N_21524,N_21583);
xnor U21963 (N_21963,N_21507,N_21198);
nand U21964 (N_21964,N_21300,N_21155);
xnor U21965 (N_21965,N_21238,N_20567);
nor U21966 (N_21966,N_20871,N_20851);
and U21967 (N_21967,N_21104,N_21050);
nor U21968 (N_21968,N_20493,N_20590);
xnor U21969 (N_21969,N_20556,N_21530);
xor U21970 (N_21970,N_20815,N_21496);
xor U21971 (N_21971,N_21508,N_21476);
nand U21972 (N_21972,N_21157,N_21498);
nor U21973 (N_21973,N_20727,N_21078);
or U21974 (N_21974,N_21153,N_21513);
nand U21975 (N_21975,N_20798,N_21440);
or U21976 (N_21976,N_20694,N_20476);
xnor U21977 (N_21977,N_20497,N_21288);
xor U21978 (N_21978,N_20806,N_21234);
or U21979 (N_21979,N_20946,N_20747);
and U21980 (N_21980,N_20627,N_20923);
and U21981 (N_21981,N_20695,N_20962);
nand U21982 (N_21982,N_21214,N_20984);
xor U21983 (N_21983,N_21376,N_20602);
or U21984 (N_21984,N_21385,N_20579);
nor U21985 (N_21985,N_20996,N_21598);
or U21986 (N_21986,N_21077,N_21272);
and U21987 (N_21987,N_21032,N_20794);
xnor U21988 (N_21988,N_20606,N_21278);
and U21989 (N_21989,N_21504,N_21519);
and U21990 (N_21990,N_21239,N_20603);
xor U21991 (N_21991,N_20574,N_21045);
nand U21992 (N_21992,N_21187,N_20660);
nor U21993 (N_21993,N_20558,N_20883);
and U21994 (N_21994,N_21195,N_20466);
nand U21995 (N_21995,N_21133,N_20824);
and U21996 (N_21996,N_21312,N_20983);
nor U21997 (N_21997,N_21563,N_20732);
nor U21998 (N_21998,N_20413,N_21362);
nand U21999 (N_21999,N_21394,N_21505);
nor U22000 (N_22000,N_20555,N_20823);
xor U22001 (N_22001,N_21534,N_20785);
and U22002 (N_22002,N_20474,N_20641);
xor U22003 (N_22003,N_21226,N_20456);
xor U22004 (N_22004,N_20639,N_20884);
and U22005 (N_22005,N_21244,N_20835);
or U22006 (N_22006,N_20521,N_21276);
nand U22007 (N_22007,N_21477,N_20410);
nor U22008 (N_22008,N_21427,N_20623);
nand U22009 (N_22009,N_20484,N_21423);
or U22010 (N_22010,N_20763,N_20975);
nand U22011 (N_22011,N_21245,N_21275);
and U22012 (N_22012,N_21473,N_20684);
xnor U22013 (N_22013,N_20807,N_21146);
xnor U22014 (N_22014,N_20546,N_20952);
and U22015 (N_22015,N_20569,N_21321);
xor U22016 (N_22016,N_20944,N_20636);
nor U22017 (N_22017,N_21445,N_20993);
nor U22018 (N_22018,N_20930,N_21123);
xor U22019 (N_22019,N_20507,N_20428);
nand U22020 (N_22020,N_20837,N_21490);
nand U22021 (N_22021,N_20810,N_20964);
nor U22022 (N_22022,N_20769,N_21254);
or U22023 (N_22023,N_20510,N_20516);
or U22024 (N_22024,N_21382,N_20848);
or U22025 (N_22025,N_20409,N_20842);
nand U22026 (N_22026,N_20592,N_20849);
and U22027 (N_22027,N_21354,N_20784);
and U22028 (N_22028,N_20971,N_20843);
or U22029 (N_22029,N_20928,N_20445);
nand U22030 (N_22030,N_21172,N_20878);
nor U22031 (N_22031,N_20450,N_20863);
nor U22032 (N_22032,N_20486,N_20652);
or U22033 (N_22033,N_20608,N_20437);
nand U22034 (N_22034,N_21487,N_20759);
and U22035 (N_22035,N_21377,N_21282);
nor U22036 (N_22036,N_20861,N_21532);
nor U22037 (N_22037,N_21576,N_20479);
and U22038 (N_22038,N_21450,N_21249);
xor U22039 (N_22039,N_20981,N_20692);
xor U22040 (N_22040,N_21305,N_20893);
or U22041 (N_22041,N_21416,N_20508);
or U22042 (N_22042,N_21002,N_21580);
xnor U22043 (N_22043,N_20502,N_21489);
or U22044 (N_22044,N_20877,N_20888);
or U22045 (N_22045,N_20654,N_20909);
and U22046 (N_22046,N_20441,N_21156);
xnor U22047 (N_22047,N_20681,N_20575);
nor U22048 (N_22048,N_20796,N_21559);
or U22049 (N_22049,N_21222,N_20773);
nor U22050 (N_22050,N_20772,N_21375);
or U22051 (N_22051,N_21399,N_21478);
xor U22052 (N_22052,N_21243,N_20557);
or U22053 (N_22053,N_20485,N_20757);
xor U22054 (N_22054,N_21587,N_21391);
or U22055 (N_22055,N_21446,N_20920);
nand U22056 (N_22056,N_21182,N_20470);
nand U22057 (N_22057,N_20938,N_21175);
and U22058 (N_22058,N_21292,N_21386);
and U22059 (N_22059,N_21237,N_20543);
and U22060 (N_22060,N_20683,N_21418);
or U22061 (N_22061,N_21235,N_21286);
and U22062 (N_22062,N_20710,N_20881);
and U22063 (N_22063,N_21270,N_21067);
and U22064 (N_22064,N_20468,N_20498);
nand U22065 (N_22065,N_20755,N_20596);
nand U22066 (N_22066,N_21026,N_21080);
nor U22067 (N_22067,N_21340,N_20693);
nor U22068 (N_22068,N_21415,N_20453);
nor U22069 (N_22069,N_20572,N_20699);
nand U22070 (N_22070,N_20529,N_20594);
and U22071 (N_22071,N_20809,N_20469);
or U22072 (N_22072,N_20777,N_20767);
nand U22073 (N_22073,N_20586,N_20951);
nand U22074 (N_22074,N_21051,N_21225);
and U22075 (N_22075,N_21413,N_21360);
nor U22076 (N_22076,N_20487,N_21262);
or U22077 (N_22077,N_21395,N_20965);
or U22078 (N_22078,N_20999,N_20853);
nor U22079 (N_22079,N_20408,N_21544);
and U22080 (N_22080,N_20787,N_21004);
xnor U22081 (N_22081,N_21213,N_21220);
or U22082 (N_22082,N_21150,N_20635);
nand U22083 (N_22083,N_20407,N_20750);
xnor U22084 (N_22084,N_20891,N_21162);
xor U22085 (N_22085,N_21464,N_20970);
or U22086 (N_22086,N_20513,N_20597);
and U22087 (N_22087,N_20426,N_20503);
and U22088 (N_22088,N_20541,N_21556);
or U22089 (N_22089,N_21029,N_21127);
xor U22090 (N_22090,N_21264,N_21125);
and U22091 (N_22091,N_21548,N_20434);
xor U22092 (N_22092,N_21124,N_20442);
or U22093 (N_22093,N_20685,N_21461);
nand U22094 (N_22094,N_21488,N_20551);
nor U22095 (N_22095,N_20477,N_21326);
and U22096 (N_22096,N_20731,N_20758);
xnor U22097 (N_22097,N_21400,N_21520);
nand U22098 (N_22098,N_21058,N_21018);
and U22099 (N_22099,N_21458,N_21042);
nand U22100 (N_22100,N_21380,N_20762);
or U22101 (N_22101,N_21302,N_20405);
xor U22102 (N_22102,N_20425,N_21398);
and U22103 (N_22103,N_21259,N_20914);
nor U22104 (N_22104,N_20790,N_21224);
xnor U22105 (N_22105,N_20729,N_20960);
xnor U22106 (N_22106,N_21432,N_20519);
nand U22107 (N_22107,N_20629,N_21096);
nor U22108 (N_22108,N_20845,N_21030);
nand U22109 (N_22109,N_21193,N_20439);
nor U22110 (N_22110,N_20898,N_20933);
nand U22111 (N_22111,N_21366,N_21444);
and U22112 (N_22112,N_20404,N_20465);
nor U22113 (N_22113,N_20564,N_21141);
nand U22114 (N_22114,N_21522,N_20467);
and U22115 (N_22115,N_21560,N_20941);
and U22116 (N_22116,N_20690,N_21494);
nand U22117 (N_22117,N_21447,N_21313);
nor U22118 (N_22118,N_21594,N_21365);
and U22119 (N_22119,N_20655,N_21083);
nand U22120 (N_22120,N_20687,N_20653);
and U22121 (N_22121,N_21036,N_20903);
xor U22122 (N_22122,N_21480,N_21479);
xor U22123 (N_22123,N_21194,N_20799);
nor U22124 (N_22124,N_21268,N_20771);
xnor U22125 (N_22125,N_21419,N_20517);
or U22126 (N_22126,N_21528,N_20577);
or U22127 (N_22127,N_21064,N_20523);
nor U22128 (N_22128,N_21206,N_20818);
nor U22129 (N_22129,N_20615,N_21414);
and U22130 (N_22130,N_21466,N_21343);
and U22131 (N_22131,N_20902,N_20622);
or U22132 (N_22132,N_20480,N_20864);
nor U22133 (N_22133,N_21570,N_20534);
xor U22134 (N_22134,N_21060,N_20746);
nor U22135 (N_22135,N_21303,N_21597);
and U22136 (N_22136,N_21515,N_21521);
xnor U22137 (N_22137,N_21325,N_21071);
nor U22138 (N_22138,N_20659,N_20673);
or U22139 (N_22139,N_20448,N_21176);
or U22140 (N_22140,N_20698,N_20705);
nand U22141 (N_22141,N_20670,N_21387);
or U22142 (N_22142,N_21263,N_21335);
or U22143 (N_22143,N_21533,N_20585);
nor U22144 (N_22144,N_20859,N_21527);
xor U22145 (N_22145,N_21112,N_20475);
nor U22146 (N_22146,N_21062,N_20797);
nor U22147 (N_22147,N_20471,N_21472);
or U22148 (N_22148,N_21482,N_21181);
nand U22149 (N_22149,N_20703,N_21179);
xnor U22150 (N_22150,N_21190,N_21492);
and U22151 (N_22151,N_21011,N_21531);
xor U22152 (N_22152,N_20892,N_20460);
xnor U22153 (N_22153,N_20991,N_20990);
nor U22154 (N_22154,N_20918,N_21308);
or U22155 (N_22155,N_20415,N_21189);
nor U22156 (N_22156,N_21113,N_20876);
nor U22157 (N_22157,N_20420,N_21207);
or U22158 (N_22158,N_20740,N_20825);
nand U22159 (N_22159,N_20931,N_21196);
and U22160 (N_22160,N_20795,N_20421);
or U22161 (N_22161,N_21509,N_20618);
nor U22162 (N_22162,N_21091,N_21252);
and U22163 (N_22163,N_20819,N_20994);
nor U22164 (N_22164,N_21054,N_20643);
nand U22165 (N_22165,N_20901,N_21008);
and U22166 (N_22166,N_21154,N_21100);
or U22167 (N_22167,N_20945,N_21145);
nor U22168 (N_22168,N_21015,N_20793);
and U22169 (N_22169,N_21074,N_20905);
or U22170 (N_22170,N_20940,N_21549);
xor U22171 (N_22171,N_21072,N_20526);
and U22172 (N_22172,N_21209,N_21429);
nand U22173 (N_22173,N_20992,N_20440);
nand U22174 (N_22174,N_21537,N_20446);
or U22175 (N_22175,N_20449,N_21352);
and U22176 (N_22176,N_21347,N_21547);
nand U22177 (N_22177,N_20801,N_20721);
or U22178 (N_22178,N_20668,N_21017);
xor U22179 (N_22179,N_21111,N_21092);
nor U22180 (N_22180,N_21253,N_20718);
or U22181 (N_22181,N_20506,N_20680);
nand U22182 (N_22182,N_20770,N_20929);
nor U22183 (N_22183,N_20880,N_20565);
or U22184 (N_22184,N_20459,N_20753);
and U22185 (N_22185,N_21044,N_20505);
nor U22186 (N_22186,N_20576,N_20743);
nor U22187 (N_22187,N_21503,N_21317);
or U22188 (N_22188,N_21468,N_20620);
or U22189 (N_22189,N_21171,N_20736);
and U22190 (N_22190,N_20527,N_21555);
nor U22191 (N_22191,N_21451,N_21085);
nor U22192 (N_22192,N_21114,N_20570);
and U22193 (N_22193,N_21438,N_20702);
xnor U22194 (N_22194,N_21269,N_20709);
nor U22195 (N_22195,N_20531,N_20406);
or U22196 (N_22196,N_21346,N_21511);
nor U22197 (N_22197,N_21090,N_21379);
and U22198 (N_22198,N_21373,N_20969);
xor U22199 (N_22199,N_20720,N_21336);
or U22200 (N_22200,N_20414,N_21001);
nor U22201 (N_22201,N_20552,N_21131);
and U22202 (N_22202,N_20962,N_20825);
xor U22203 (N_22203,N_20901,N_21084);
or U22204 (N_22204,N_20531,N_21311);
or U22205 (N_22205,N_21535,N_20538);
xnor U22206 (N_22206,N_20518,N_20487);
or U22207 (N_22207,N_21257,N_21118);
nand U22208 (N_22208,N_20776,N_21249);
xnor U22209 (N_22209,N_21077,N_20505);
xnor U22210 (N_22210,N_21109,N_20670);
and U22211 (N_22211,N_21523,N_21232);
and U22212 (N_22212,N_20705,N_20446);
xor U22213 (N_22213,N_20970,N_21376);
nor U22214 (N_22214,N_21488,N_20799);
xor U22215 (N_22215,N_21197,N_20948);
and U22216 (N_22216,N_20635,N_20693);
nand U22217 (N_22217,N_21251,N_20980);
xor U22218 (N_22218,N_21386,N_20979);
nor U22219 (N_22219,N_21332,N_21169);
or U22220 (N_22220,N_21285,N_21520);
xor U22221 (N_22221,N_20530,N_21155);
or U22222 (N_22222,N_21544,N_20652);
nor U22223 (N_22223,N_20654,N_20406);
or U22224 (N_22224,N_20427,N_20846);
xor U22225 (N_22225,N_20899,N_20533);
and U22226 (N_22226,N_21047,N_20758);
xnor U22227 (N_22227,N_20821,N_21227);
xor U22228 (N_22228,N_21018,N_20523);
and U22229 (N_22229,N_20457,N_21463);
and U22230 (N_22230,N_21132,N_21296);
nor U22231 (N_22231,N_21465,N_21200);
nand U22232 (N_22232,N_20650,N_20974);
nand U22233 (N_22233,N_20449,N_21121);
or U22234 (N_22234,N_21265,N_21354);
nor U22235 (N_22235,N_20438,N_20951);
or U22236 (N_22236,N_20415,N_21056);
nor U22237 (N_22237,N_21161,N_20567);
xor U22238 (N_22238,N_21272,N_20747);
or U22239 (N_22239,N_21318,N_21165);
nand U22240 (N_22240,N_20403,N_20783);
xor U22241 (N_22241,N_20931,N_21275);
and U22242 (N_22242,N_20786,N_21311);
nand U22243 (N_22243,N_20409,N_21340);
nand U22244 (N_22244,N_20431,N_21165);
or U22245 (N_22245,N_20956,N_21358);
nor U22246 (N_22246,N_20955,N_20832);
nand U22247 (N_22247,N_21209,N_21521);
or U22248 (N_22248,N_20833,N_20420);
nor U22249 (N_22249,N_20968,N_20657);
xor U22250 (N_22250,N_20939,N_20504);
nor U22251 (N_22251,N_21290,N_20811);
or U22252 (N_22252,N_21443,N_20541);
xnor U22253 (N_22253,N_20836,N_21308);
and U22254 (N_22254,N_20622,N_20881);
xor U22255 (N_22255,N_20654,N_20659);
xnor U22256 (N_22256,N_21349,N_20987);
xor U22257 (N_22257,N_20756,N_21588);
nand U22258 (N_22258,N_21155,N_20804);
or U22259 (N_22259,N_20728,N_21478);
nor U22260 (N_22260,N_21284,N_21163);
or U22261 (N_22261,N_21390,N_21503);
xnor U22262 (N_22262,N_21155,N_21162);
nand U22263 (N_22263,N_20643,N_21305);
or U22264 (N_22264,N_21276,N_21155);
and U22265 (N_22265,N_20908,N_20719);
and U22266 (N_22266,N_21213,N_20678);
and U22267 (N_22267,N_20562,N_21340);
or U22268 (N_22268,N_21522,N_21064);
nand U22269 (N_22269,N_20494,N_21489);
xor U22270 (N_22270,N_21418,N_20968);
xnor U22271 (N_22271,N_20679,N_21088);
and U22272 (N_22272,N_21225,N_20412);
nor U22273 (N_22273,N_20455,N_21458);
nor U22274 (N_22274,N_20653,N_21144);
or U22275 (N_22275,N_21308,N_21570);
nor U22276 (N_22276,N_21593,N_21511);
or U22277 (N_22277,N_20849,N_20496);
nand U22278 (N_22278,N_21065,N_21370);
nor U22279 (N_22279,N_21549,N_21339);
xor U22280 (N_22280,N_21067,N_20470);
or U22281 (N_22281,N_21090,N_20409);
nor U22282 (N_22282,N_20578,N_20538);
and U22283 (N_22283,N_21405,N_21209);
xor U22284 (N_22284,N_20485,N_20461);
and U22285 (N_22285,N_20594,N_21476);
nor U22286 (N_22286,N_20843,N_20732);
and U22287 (N_22287,N_20659,N_21470);
or U22288 (N_22288,N_20764,N_20700);
nor U22289 (N_22289,N_20851,N_21121);
nor U22290 (N_22290,N_21308,N_20951);
nand U22291 (N_22291,N_21577,N_20646);
or U22292 (N_22292,N_21489,N_21096);
xor U22293 (N_22293,N_21563,N_21158);
or U22294 (N_22294,N_20529,N_21077);
and U22295 (N_22295,N_21225,N_20603);
nand U22296 (N_22296,N_20455,N_21334);
nand U22297 (N_22297,N_20605,N_21053);
or U22298 (N_22298,N_20535,N_21332);
nor U22299 (N_22299,N_20541,N_20661);
nand U22300 (N_22300,N_20857,N_21410);
nand U22301 (N_22301,N_20657,N_20432);
and U22302 (N_22302,N_21376,N_20475);
or U22303 (N_22303,N_20914,N_21352);
nand U22304 (N_22304,N_21045,N_20520);
and U22305 (N_22305,N_20631,N_21511);
and U22306 (N_22306,N_20598,N_20949);
or U22307 (N_22307,N_21253,N_21573);
xor U22308 (N_22308,N_21476,N_21392);
nor U22309 (N_22309,N_21447,N_21121);
nand U22310 (N_22310,N_20504,N_21032);
nand U22311 (N_22311,N_21010,N_21401);
nand U22312 (N_22312,N_20969,N_20437);
or U22313 (N_22313,N_21016,N_21571);
nand U22314 (N_22314,N_20874,N_21444);
nand U22315 (N_22315,N_21595,N_20423);
or U22316 (N_22316,N_21146,N_21342);
or U22317 (N_22317,N_21158,N_20852);
or U22318 (N_22318,N_20607,N_20896);
nor U22319 (N_22319,N_21208,N_21265);
nor U22320 (N_22320,N_20811,N_21553);
or U22321 (N_22321,N_20807,N_21247);
xor U22322 (N_22322,N_21025,N_20504);
nor U22323 (N_22323,N_20534,N_21205);
nand U22324 (N_22324,N_20976,N_20460);
nor U22325 (N_22325,N_21552,N_21211);
nand U22326 (N_22326,N_20719,N_21135);
and U22327 (N_22327,N_21109,N_20822);
xnor U22328 (N_22328,N_20622,N_20718);
or U22329 (N_22329,N_20893,N_20863);
nand U22330 (N_22330,N_21414,N_20989);
and U22331 (N_22331,N_20800,N_20976);
xnor U22332 (N_22332,N_21139,N_20571);
nor U22333 (N_22333,N_21553,N_21331);
xnor U22334 (N_22334,N_20907,N_21138);
xnor U22335 (N_22335,N_21066,N_20784);
xor U22336 (N_22336,N_20739,N_20911);
or U22337 (N_22337,N_20521,N_21097);
or U22338 (N_22338,N_21292,N_21478);
nand U22339 (N_22339,N_21134,N_21376);
xnor U22340 (N_22340,N_21394,N_21509);
xor U22341 (N_22341,N_21435,N_20920);
nor U22342 (N_22342,N_21380,N_21409);
or U22343 (N_22343,N_21177,N_21508);
nand U22344 (N_22344,N_20560,N_21591);
nand U22345 (N_22345,N_20990,N_21355);
xor U22346 (N_22346,N_20835,N_21179);
and U22347 (N_22347,N_20401,N_21489);
nand U22348 (N_22348,N_21238,N_21091);
or U22349 (N_22349,N_21382,N_21243);
or U22350 (N_22350,N_21550,N_20887);
nor U22351 (N_22351,N_21490,N_20644);
and U22352 (N_22352,N_21228,N_21135);
or U22353 (N_22353,N_20920,N_20449);
nand U22354 (N_22354,N_21007,N_20686);
and U22355 (N_22355,N_21581,N_21361);
nand U22356 (N_22356,N_20819,N_21426);
and U22357 (N_22357,N_21301,N_20408);
nand U22358 (N_22358,N_21325,N_20897);
and U22359 (N_22359,N_21518,N_20463);
and U22360 (N_22360,N_21486,N_21513);
nor U22361 (N_22361,N_21525,N_20494);
nand U22362 (N_22362,N_20453,N_20913);
or U22363 (N_22363,N_20777,N_20819);
nor U22364 (N_22364,N_21323,N_21230);
xor U22365 (N_22365,N_20831,N_21560);
and U22366 (N_22366,N_20469,N_21519);
and U22367 (N_22367,N_21306,N_20472);
nand U22368 (N_22368,N_20741,N_20939);
xor U22369 (N_22369,N_20721,N_21561);
nor U22370 (N_22370,N_21500,N_20494);
or U22371 (N_22371,N_21526,N_20821);
nand U22372 (N_22372,N_20474,N_21261);
nor U22373 (N_22373,N_20437,N_20907);
or U22374 (N_22374,N_20795,N_21092);
and U22375 (N_22375,N_21166,N_20639);
nor U22376 (N_22376,N_20768,N_21292);
and U22377 (N_22377,N_21457,N_21166);
nand U22378 (N_22378,N_20675,N_21159);
nor U22379 (N_22379,N_20554,N_21414);
or U22380 (N_22380,N_20939,N_21596);
and U22381 (N_22381,N_20844,N_21472);
nand U22382 (N_22382,N_20966,N_21402);
and U22383 (N_22383,N_21134,N_20862);
nand U22384 (N_22384,N_21538,N_21487);
nand U22385 (N_22385,N_21378,N_20824);
nor U22386 (N_22386,N_21599,N_21353);
nand U22387 (N_22387,N_21374,N_21424);
and U22388 (N_22388,N_20908,N_21499);
nor U22389 (N_22389,N_21427,N_20516);
or U22390 (N_22390,N_21533,N_20406);
nand U22391 (N_22391,N_20511,N_20931);
and U22392 (N_22392,N_21219,N_21051);
xor U22393 (N_22393,N_20841,N_21357);
nor U22394 (N_22394,N_21059,N_21144);
nor U22395 (N_22395,N_20476,N_20596);
and U22396 (N_22396,N_21523,N_21176);
and U22397 (N_22397,N_20522,N_20631);
nor U22398 (N_22398,N_21119,N_21446);
nor U22399 (N_22399,N_21112,N_20809);
and U22400 (N_22400,N_21553,N_20783);
nand U22401 (N_22401,N_20928,N_20857);
nor U22402 (N_22402,N_20420,N_21513);
nor U22403 (N_22403,N_21461,N_20920);
and U22404 (N_22404,N_20582,N_20769);
nor U22405 (N_22405,N_20430,N_21190);
nand U22406 (N_22406,N_21215,N_20626);
xor U22407 (N_22407,N_21401,N_21419);
and U22408 (N_22408,N_21261,N_21307);
and U22409 (N_22409,N_21171,N_20481);
and U22410 (N_22410,N_20932,N_20580);
and U22411 (N_22411,N_21592,N_20749);
and U22412 (N_22412,N_21073,N_20748);
or U22413 (N_22413,N_21142,N_21016);
xor U22414 (N_22414,N_20591,N_21046);
nor U22415 (N_22415,N_21237,N_20426);
or U22416 (N_22416,N_20811,N_21335);
xnor U22417 (N_22417,N_21118,N_20747);
nand U22418 (N_22418,N_21133,N_21066);
or U22419 (N_22419,N_21425,N_21589);
and U22420 (N_22420,N_20772,N_21203);
or U22421 (N_22421,N_21578,N_21214);
or U22422 (N_22422,N_21121,N_21248);
nand U22423 (N_22423,N_20825,N_20729);
xor U22424 (N_22424,N_21363,N_20604);
and U22425 (N_22425,N_21168,N_20686);
nor U22426 (N_22426,N_21343,N_21536);
nand U22427 (N_22427,N_20470,N_20590);
and U22428 (N_22428,N_21353,N_20589);
nand U22429 (N_22429,N_21050,N_21062);
and U22430 (N_22430,N_21195,N_21447);
and U22431 (N_22431,N_20985,N_21413);
and U22432 (N_22432,N_21443,N_21020);
nor U22433 (N_22433,N_20522,N_21476);
xor U22434 (N_22434,N_20816,N_21545);
xnor U22435 (N_22435,N_21285,N_21592);
nor U22436 (N_22436,N_20761,N_20908);
or U22437 (N_22437,N_20728,N_20597);
nor U22438 (N_22438,N_21471,N_20645);
and U22439 (N_22439,N_20889,N_20913);
xor U22440 (N_22440,N_21389,N_21289);
or U22441 (N_22441,N_20723,N_20917);
nand U22442 (N_22442,N_20807,N_20939);
xnor U22443 (N_22443,N_21562,N_20872);
and U22444 (N_22444,N_20720,N_20546);
or U22445 (N_22445,N_21050,N_20995);
nor U22446 (N_22446,N_20737,N_20728);
nand U22447 (N_22447,N_20627,N_21541);
nor U22448 (N_22448,N_21398,N_21088);
xnor U22449 (N_22449,N_21330,N_20478);
and U22450 (N_22450,N_21035,N_21123);
xnor U22451 (N_22451,N_20868,N_21299);
and U22452 (N_22452,N_20678,N_20838);
nor U22453 (N_22453,N_20902,N_20437);
and U22454 (N_22454,N_21230,N_20686);
or U22455 (N_22455,N_21445,N_21261);
nor U22456 (N_22456,N_21121,N_20836);
and U22457 (N_22457,N_20762,N_20455);
nor U22458 (N_22458,N_20461,N_20971);
xnor U22459 (N_22459,N_21548,N_20417);
nand U22460 (N_22460,N_20678,N_21460);
nor U22461 (N_22461,N_20783,N_21090);
and U22462 (N_22462,N_21419,N_20786);
or U22463 (N_22463,N_21442,N_20790);
xor U22464 (N_22464,N_20825,N_21142);
and U22465 (N_22465,N_21005,N_20570);
nand U22466 (N_22466,N_21102,N_20462);
or U22467 (N_22467,N_21099,N_21395);
and U22468 (N_22468,N_20937,N_20455);
xor U22469 (N_22469,N_20524,N_20995);
nor U22470 (N_22470,N_20772,N_20452);
or U22471 (N_22471,N_21360,N_21480);
xor U22472 (N_22472,N_20857,N_21596);
xnor U22473 (N_22473,N_20850,N_21461);
or U22474 (N_22474,N_20616,N_21284);
nand U22475 (N_22475,N_21179,N_20592);
or U22476 (N_22476,N_21450,N_21248);
nand U22477 (N_22477,N_21144,N_21593);
xnor U22478 (N_22478,N_21500,N_21052);
nor U22479 (N_22479,N_21594,N_20817);
nor U22480 (N_22480,N_21195,N_21508);
nor U22481 (N_22481,N_20949,N_20635);
xor U22482 (N_22482,N_21472,N_20424);
nor U22483 (N_22483,N_20855,N_21144);
or U22484 (N_22484,N_20577,N_21513);
and U22485 (N_22485,N_21325,N_20484);
nor U22486 (N_22486,N_20931,N_21307);
or U22487 (N_22487,N_20757,N_21134);
or U22488 (N_22488,N_20679,N_21562);
nand U22489 (N_22489,N_20445,N_20553);
nor U22490 (N_22490,N_21038,N_20770);
nand U22491 (N_22491,N_21014,N_21130);
nor U22492 (N_22492,N_20455,N_20862);
xnor U22493 (N_22493,N_21193,N_21239);
nand U22494 (N_22494,N_20425,N_20749);
xor U22495 (N_22495,N_20809,N_21185);
nand U22496 (N_22496,N_20736,N_20400);
nand U22497 (N_22497,N_20769,N_21520);
nand U22498 (N_22498,N_21309,N_21380);
or U22499 (N_22499,N_21023,N_20704);
xnor U22500 (N_22500,N_21489,N_21514);
and U22501 (N_22501,N_20976,N_20539);
nand U22502 (N_22502,N_20834,N_21480);
or U22503 (N_22503,N_21582,N_21089);
and U22504 (N_22504,N_21039,N_20442);
and U22505 (N_22505,N_21061,N_20657);
or U22506 (N_22506,N_21429,N_21343);
and U22507 (N_22507,N_21482,N_21247);
nand U22508 (N_22508,N_21457,N_20843);
nand U22509 (N_22509,N_20833,N_21299);
xnor U22510 (N_22510,N_21597,N_21012);
nor U22511 (N_22511,N_21432,N_21008);
and U22512 (N_22512,N_21202,N_20655);
nand U22513 (N_22513,N_20593,N_20926);
or U22514 (N_22514,N_21367,N_20940);
xnor U22515 (N_22515,N_20701,N_20962);
or U22516 (N_22516,N_21239,N_20896);
nand U22517 (N_22517,N_21279,N_21592);
nor U22518 (N_22518,N_20710,N_21471);
nand U22519 (N_22519,N_21556,N_21427);
and U22520 (N_22520,N_21489,N_20472);
nor U22521 (N_22521,N_20824,N_20450);
nand U22522 (N_22522,N_20817,N_21365);
and U22523 (N_22523,N_21491,N_21192);
xor U22524 (N_22524,N_20711,N_21323);
or U22525 (N_22525,N_21541,N_21424);
and U22526 (N_22526,N_20722,N_21001);
nor U22527 (N_22527,N_20798,N_20603);
and U22528 (N_22528,N_20638,N_20963);
and U22529 (N_22529,N_20946,N_21186);
or U22530 (N_22530,N_21079,N_21385);
nand U22531 (N_22531,N_20458,N_20835);
or U22532 (N_22532,N_21171,N_20513);
nor U22533 (N_22533,N_20683,N_20625);
and U22534 (N_22534,N_21422,N_20786);
xor U22535 (N_22535,N_21485,N_20613);
nand U22536 (N_22536,N_21434,N_21512);
xnor U22537 (N_22537,N_21213,N_21022);
nand U22538 (N_22538,N_20864,N_21508);
or U22539 (N_22539,N_20544,N_20422);
and U22540 (N_22540,N_20952,N_21228);
xnor U22541 (N_22541,N_20723,N_21581);
nand U22542 (N_22542,N_20586,N_20592);
or U22543 (N_22543,N_20677,N_21148);
or U22544 (N_22544,N_20757,N_20687);
nand U22545 (N_22545,N_20679,N_20852);
and U22546 (N_22546,N_21508,N_20643);
nand U22547 (N_22547,N_20950,N_21166);
nor U22548 (N_22548,N_21342,N_20959);
and U22549 (N_22549,N_20444,N_20547);
nor U22550 (N_22550,N_20785,N_20741);
xnor U22551 (N_22551,N_21247,N_20434);
nand U22552 (N_22552,N_20641,N_21027);
nand U22553 (N_22553,N_20871,N_21359);
nor U22554 (N_22554,N_21140,N_20588);
or U22555 (N_22555,N_21505,N_21466);
or U22556 (N_22556,N_20421,N_21070);
or U22557 (N_22557,N_20419,N_21135);
and U22558 (N_22558,N_21084,N_21431);
nor U22559 (N_22559,N_20899,N_21228);
and U22560 (N_22560,N_20464,N_20789);
or U22561 (N_22561,N_20430,N_21566);
nor U22562 (N_22562,N_20819,N_20596);
nand U22563 (N_22563,N_21045,N_20412);
nand U22564 (N_22564,N_20962,N_20992);
and U22565 (N_22565,N_20453,N_20537);
nor U22566 (N_22566,N_20872,N_20880);
nor U22567 (N_22567,N_20735,N_20617);
or U22568 (N_22568,N_20407,N_20861);
nand U22569 (N_22569,N_21041,N_20538);
or U22570 (N_22570,N_21180,N_20846);
and U22571 (N_22571,N_20735,N_20463);
nand U22572 (N_22572,N_20769,N_21352);
nor U22573 (N_22573,N_21587,N_20831);
nor U22574 (N_22574,N_20587,N_21235);
nor U22575 (N_22575,N_21276,N_20538);
nor U22576 (N_22576,N_21459,N_21413);
nand U22577 (N_22577,N_20898,N_20718);
nand U22578 (N_22578,N_21597,N_21217);
xnor U22579 (N_22579,N_21495,N_21386);
nor U22580 (N_22580,N_21404,N_21415);
and U22581 (N_22581,N_20922,N_21330);
or U22582 (N_22582,N_20978,N_20664);
xnor U22583 (N_22583,N_21141,N_21428);
nor U22584 (N_22584,N_21570,N_21494);
nand U22585 (N_22585,N_21091,N_20433);
or U22586 (N_22586,N_21200,N_20480);
nand U22587 (N_22587,N_20464,N_20576);
xor U22588 (N_22588,N_21019,N_20639);
xnor U22589 (N_22589,N_20552,N_21426);
xnor U22590 (N_22590,N_20715,N_21144);
or U22591 (N_22591,N_20782,N_21414);
xor U22592 (N_22592,N_20759,N_21269);
or U22593 (N_22593,N_21344,N_20944);
nand U22594 (N_22594,N_20725,N_21307);
nor U22595 (N_22595,N_20442,N_21298);
or U22596 (N_22596,N_21131,N_20403);
and U22597 (N_22597,N_21553,N_21531);
xor U22598 (N_22598,N_20823,N_20634);
or U22599 (N_22599,N_20415,N_21447);
or U22600 (N_22600,N_21553,N_21567);
nor U22601 (N_22601,N_20582,N_20439);
nor U22602 (N_22602,N_21066,N_21289);
nand U22603 (N_22603,N_20690,N_20907);
and U22604 (N_22604,N_20854,N_20483);
nor U22605 (N_22605,N_21592,N_20442);
nor U22606 (N_22606,N_21126,N_20820);
nand U22607 (N_22607,N_21510,N_21487);
xor U22608 (N_22608,N_20860,N_20720);
xor U22609 (N_22609,N_21485,N_20642);
or U22610 (N_22610,N_20676,N_21438);
xnor U22611 (N_22611,N_20564,N_21568);
or U22612 (N_22612,N_21340,N_20958);
and U22613 (N_22613,N_20983,N_20600);
nand U22614 (N_22614,N_21278,N_20797);
xor U22615 (N_22615,N_20732,N_20450);
xnor U22616 (N_22616,N_20920,N_21521);
or U22617 (N_22617,N_21549,N_20480);
or U22618 (N_22618,N_20987,N_21181);
and U22619 (N_22619,N_20716,N_20803);
and U22620 (N_22620,N_21235,N_21293);
nor U22621 (N_22621,N_21495,N_21182);
nand U22622 (N_22622,N_20439,N_21336);
and U22623 (N_22623,N_21444,N_21598);
xnor U22624 (N_22624,N_21123,N_20540);
or U22625 (N_22625,N_21109,N_20961);
and U22626 (N_22626,N_20621,N_21122);
and U22627 (N_22627,N_20566,N_21195);
xor U22628 (N_22628,N_21014,N_21008);
nand U22629 (N_22629,N_20755,N_20532);
and U22630 (N_22630,N_20424,N_21597);
nand U22631 (N_22631,N_20856,N_20895);
xor U22632 (N_22632,N_20795,N_20721);
and U22633 (N_22633,N_21161,N_21058);
and U22634 (N_22634,N_21433,N_21541);
or U22635 (N_22635,N_20560,N_20415);
or U22636 (N_22636,N_21436,N_21475);
nor U22637 (N_22637,N_20630,N_20871);
nand U22638 (N_22638,N_20711,N_20886);
nand U22639 (N_22639,N_20786,N_21000);
nand U22640 (N_22640,N_20538,N_21530);
nand U22641 (N_22641,N_20405,N_20557);
or U22642 (N_22642,N_21410,N_20576);
and U22643 (N_22643,N_20487,N_21160);
nand U22644 (N_22644,N_20828,N_21079);
or U22645 (N_22645,N_21066,N_20729);
nor U22646 (N_22646,N_21356,N_20857);
or U22647 (N_22647,N_21249,N_21140);
and U22648 (N_22648,N_20884,N_20936);
nand U22649 (N_22649,N_21095,N_21569);
or U22650 (N_22650,N_21210,N_21245);
and U22651 (N_22651,N_20887,N_21293);
xor U22652 (N_22652,N_20704,N_21142);
and U22653 (N_22653,N_20932,N_21304);
and U22654 (N_22654,N_20961,N_21392);
or U22655 (N_22655,N_21307,N_20565);
nor U22656 (N_22656,N_21370,N_20519);
nand U22657 (N_22657,N_20762,N_21393);
nand U22658 (N_22658,N_20501,N_20409);
xnor U22659 (N_22659,N_20744,N_20834);
xor U22660 (N_22660,N_20501,N_20447);
or U22661 (N_22661,N_20877,N_21204);
and U22662 (N_22662,N_20712,N_20670);
xor U22663 (N_22663,N_20873,N_21517);
and U22664 (N_22664,N_21363,N_20813);
xnor U22665 (N_22665,N_21539,N_21040);
nand U22666 (N_22666,N_20418,N_21084);
or U22667 (N_22667,N_21310,N_20405);
xnor U22668 (N_22668,N_21226,N_21266);
xnor U22669 (N_22669,N_20952,N_20805);
nor U22670 (N_22670,N_21564,N_20820);
nor U22671 (N_22671,N_20869,N_21011);
and U22672 (N_22672,N_21033,N_21202);
xor U22673 (N_22673,N_20587,N_20499);
nor U22674 (N_22674,N_20472,N_21139);
nor U22675 (N_22675,N_21104,N_20884);
nand U22676 (N_22676,N_21511,N_21544);
or U22677 (N_22677,N_20547,N_20443);
or U22678 (N_22678,N_20672,N_20786);
nor U22679 (N_22679,N_21469,N_21280);
xor U22680 (N_22680,N_21274,N_20470);
or U22681 (N_22681,N_21440,N_21595);
xnor U22682 (N_22682,N_21582,N_21130);
xnor U22683 (N_22683,N_20510,N_21142);
nand U22684 (N_22684,N_21191,N_21547);
or U22685 (N_22685,N_21475,N_21339);
or U22686 (N_22686,N_20537,N_21349);
or U22687 (N_22687,N_20951,N_20605);
nor U22688 (N_22688,N_21598,N_20799);
xor U22689 (N_22689,N_21123,N_20562);
nor U22690 (N_22690,N_20842,N_20963);
and U22691 (N_22691,N_21420,N_20803);
nand U22692 (N_22692,N_20805,N_21496);
and U22693 (N_22693,N_21332,N_21150);
xor U22694 (N_22694,N_21585,N_20780);
and U22695 (N_22695,N_20827,N_20531);
nand U22696 (N_22696,N_21355,N_20646);
nand U22697 (N_22697,N_21313,N_21390);
or U22698 (N_22698,N_20867,N_21523);
and U22699 (N_22699,N_20727,N_20413);
and U22700 (N_22700,N_20767,N_21400);
nand U22701 (N_22701,N_21154,N_21315);
or U22702 (N_22702,N_21588,N_20997);
or U22703 (N_22703,N_21318,N_20498);
nand U22704 (N_22704,N_20906,N_20759);
xnor U22705 (N_22705,N_20625,N_20400);
xnor U22706 (N_22706,N_20966,N_20605);
or U22707 (N_22707,N_20949,N_21461);
nor U22708 (N_22708,N_20501,N_21338);
and U22709 (N_22709,N_20657,N_21130);
nand U22710 (N_22710,N_21591,N_21223);
or U22711 (N_22711,N_20512,N_20528);
nand U22712 (N_22712,N_21043,N_20423);
nand U22713 (N_22713,N_21342,N_20503);
or U22714 (N_22714,N_20567,N_21183);
or U22715 (N_22715,N_21241,N_20755);
nor U22716 (N_22716,N_20676,N_20779);
or U22717 (N_22717,N_21311,N_20703);
and U22718 (N_22718,N_21294,N_20978);
or U22719 (N_22719,N_20755,N_21538);
xnor U22720 (N_22720,N_21142,N_21208);
nor U22721 (N_22721,N_21151,N_20830);
or U22722 (N_22722,N_20743,N_21586);
and U22723 (N_22723,N_20952,N_20424);
or U22724 (N_22724,N_21155,N_21016);
nor U22725 (N_22725,N_21394,N_20537);
or U22726 (N_22726,N_20564,N_20711);
and U22727 (N_22727,N_20542,N_21164);
xor U22728 (N_22728,N_20508,N_20860);
nor U22729 (N_22729,N_20817,N_21133);
xnor U22730 (N_22730,N_20996,N_21154);
nor U22731 (N_22731,N_20745,N_21397);
nor U22732 (N_22732,N_21122,N_20414);
and U22733 (N_22733,N_20488,N_21160);
or U22734 (N_22734,N_21429,N_21150);
or U22735 (N_22735,N_21037,N_20836);
nand U22736 (N_22736,N_20406,N_21321);
nand U22737 (N_22737,N_21222,N_20859);
or U22738 (N_22738,N_21191,N_21006);
and U22739 (N_22739,N_21313,N_20704);
nand U22740 (N_22740,N_21066,N_21496);
nand U22741 (N_22741,N_20499,N_21424);
or U22742 (N_22742,N_20471,N_20686);
and U22743 (N_22743,N_20924,N_20666);
and U22744 (N_22744,N_20669,N_20454);
xor U22745 (N_22745,N_20720,N_20653);
or U22746 (N_22746,N_20785,N_20620);
nor U22747 (N_22747,N_21238,N_20563);
or U22748 (N_22748,N_21165,N_20923);
xnor U22749 (N_22749,N_20837,N_20574);
and U22750 (N_22750,N_21450,N_20669);
and U22751 (N_22751,N_21497,N_20832);
xor U22752 (N_22752,N_21452,N_21564);
or U22753 (N_22753,N_20723,N_21224);
or U22754 (N_22754,N_20712,N_21253);
and U22755 (N_22755,N_21168,N_21314);
nor U22756 (N_22756,N_20890,N_21121);
nand U22757 (N_22757,N_21158,N_21539);
or U22758 (N_22758,N_20872,N_21552);
and U22759 (N_22759,N_20770,N_20545);
nand U22760 (N_22760,N_20971,N_21285);
and U22761 (N_22761,N_21512,N_21595);
xor U22762 (N_22762,N_21511,N_21061);
nand U22763 (N_22763,N_21578,N_20749);
xor U22764 (N_22764,N_21078,N_20880);
xor U22765 (N_22765,N_21461,N_20743);
nor U22766 (N_22766,N_20782,N_20710);
and U22767 (N_22767,N_21447,N_20765);
and U22768 (N_22768,N_20947,N_21120);
and U22769 (N_22769,N_20815,N_21231);
and U22770 (N_22770,N_20463,N_20962);
xor U22771 (N_22771,N_21017,N_21006);
nor U22772 (N_22772,N_21573,N_20616);
or U22773 (N_22773,N_21338,N_20871);
and U22774 (N_22774,N_20898,N_21048);
nor U22775 (N_22775,N_21027,N_20424);
and U22776 (N_22776,N_21129,N_21303);
and U22777 (N_22777,N_20477,N_21269);
xor U22778 (N_22778,N_21303,N_20407);
nor U22779 (N_22779,N_20765,N_21136);
and U22780 (N_22780,N_21596,N_20740);
or U22781 (N_22781,N_21275,N_20436);
nand U22782 (N_22782,N_21024,N_21069);
and U22783 (N_22783,N_20863,N_20825);
and U22784 (N_22784,N_20813,N_20401);
xor U22785 (N_22785,N_21541,N_20694);
or U22786 (N_22786,N_20594,N_21353);
nand U22787 (N_22787,N_20793,N_21027);
and U22788 (N_22788,N_21191,N_20509);
nor U22789 (N_22789,N_20907,N_20477);
xnor U22790 (N_22790,N_21101,N_20787);
nor U22791 (N_22791,N_21592,N_20739);
nand U22792 (N_22792,N_21502,N_20600);
nor U22793 (N_22793,N_21307,N_20973);
or U22794 (N_22794,N_21397,N_20940);
or U22795 (N_22795,N_20566,N_21580);
or U22796 (N_22796,N_20602,N_21188);
or U22797 (N_22797,N_21060,N_20806);
nand U22798 (N_22798,N_20537,N_20845);
nor U22799 (N_22799,N_21177,N_21358);
and U22800 (N_22800,N_21694,N_21946);
nand U22801 (N_22801,N_22117,N_22779);
and U22802 (N_22802,N_22138,N_21721);
nor U22803 (N_22803,N_22163,N_22394);
or U22804 (N_22804,N_21658,N_22061);
xnor U22805 (N_22805,N_22609,N_22716);
and U22806 (N_22806,N_22194,N_22282);
and U22807 (N_22807,N_21808,N_21827);
nor U22808 (N_22808,N_22104,N_22726);
xnor U22809 (N_22809,N_21720,N_22788);
nand U22810 (N_22810,N_21732,N_21977);
nand U22811 (N_22811,N_21943,N_21743);
nor U22812 (N_22812,N_22276,N_22401);
nand U22813 (N_22813,N_22233,N_21918);
nor U22814 (N_22814,N_22483,N_21930);
nor U22815 (N_22815,N_21723,N_22680);
and U22816 (N_22816,N_22247,N_21844);
nor U22817 (N_22817,N_22546,N_22457);
nand U22818 (N_22818,N_22717,N_22371);
or U22819 (N_22819,N_22008,N_22407);
or U22820 (N_22820,N_22441,N_22711);
xnor U22821 (N_22821,N_21874,N_21708);
and U22822 (N_22822,N_22571,N_22622);
or U22823 (N_22823,N_22387,N_22792);
and U22824 (N_22824,N_21843,N_22206);
xor U22825 (N_22825,N_21901,N_22604);
and U22826 (N_22826,N_22314,N_22340);
and U22827 (N_22827,N_22473,N_21745);
xor U22828 (N_22828,N_22587,N_22029);
xnor U22829 (N_22829,N_21957,N_22542);
or U22830 (N_22830,N_22730,N_21979);
nand U22831 (N_22831,N_22383,N_22057);
xnor U22832 (N_22832,N_22005,N_22279);
or U22833 (N_22833,N_22082,N_22491);
nand U22834 (N_22834,N_21631,N_21606);
xnor U22835 (N_22835,N_22060,N_22582);
or U22836 (N_22836,N_22151,N_21832);
nor U22837 (N_22837,N_22762,N_22778);
nand U22838 (N_22838,N_22493,N_22770);
and U22839 (N_22839,N_21639,N_21651);
or U22840 (N_22840,N_21705,N_21965);
nand U22841 (N_22841,N_22180,N_22280);
nor U22842 (N_22842,N_22443,N_22537);
xnor U22843 (N_22843,N_22187,N_22369);
or U22844 (N_22844,N_22162,N_21649);
nor U22845 (N_22845,N_22055,N_22793);
and U22846 (N_22846,N_22456,N_21933);
nand U22847 (N_22847,N_22649,N_21913);
xnor U22848 (N_22848,N_22112,N_22025);
xor U22849 (N_22849,N_22244,N_22004);
nand U22850 (N_22850,N_22523,N_21703);
or U22851 (N_22851,N_22093,N_21896);
nor U22852 (N_22852,N_21948,N_22050);
and U22853 (N_22853,N_22591,N_21941);
nand U22854 (N_22854,N_22467,N_21994);
nor U22855 (N_22855,N_21895,N_21771);
nand U22856 (N_22856,N_21886,N_22500);
and U22857 (N_22857,N_22507,N_22704);
xor U22858 (N_22858,N_22439,N_22254);
nor U22859 (N_22859,N_21750,N_21877);
or U22860 (N_22860,N_21812,N_22414);
xor U22861 (N_22861,N_22627,N_21902);
nand U22862 (N_22862,N_22035,N_22389);
or U22863 (N_22863,N_22201,N_22746);
nor U22864 (N_22864,N_22406,N_21780);
or U22865 (N_22865,N_22777,N_22193);
nor U22866 (N_22866,N_22196,N_22429);
xnor U22867 (N_22867,N_22402,N_22326);
xnor U22868 (N_22868,N_21984,N_22696);
nand U22869 (N_22869,N_22040,N_22111);
nor U22870 (N_22870,N_21791,N_22653);
xnor U22871 (N_22871,N_21897,N_21833);
xor U22872 (N_22872,N_22219,N_22337);
or U22873 (N_22873,N_21730,N_22228);
nand U22874 (N_22874,N_21648,N_22742);
and U22875 (N_22875,N_22304,N_22287);
and U22876 (N_22876,N_21635,N_22095);
xor U22877 (N_22877,N_22092,N_22434);
or U22878 (N_22878,N_22141,N_22397);
or U22879 (N_22879,N_22221,N_22678);
or U22880 (N_22880,N_22787,N_22548);
and U22881 (N_22881,N_22422,N_22318);
and U22882 (N_22882,N_22416,N_21688);
or U22883 (N_22883,N_21914,N_22642);
nand U22884 (N_22884,N_22789,N_21835);
nor U22885 (N_22885,N_22713,N_21711);
and U22886 (N_22886,N_21959,N_22675);
or U22887 (N_22887,N_22066,N_22010);
nand U22888 (N_22888,N_22661,N_22094);
nor U22889 (N_22889,N_22300,N_22056);
and U22890 (N_22890,N_22695,N_22765);
or U22891 (N_22891,N_22698,N_21935);
nor U22892 (N_22892,N_22692,N_21638);
and U22893 (N_22893,N_22574,N_22553);
or U22894 (N_22894,N_21970,N_21675);
or U22895 (N_22895,N_22305,N_21868);
nand U22896 (N_22896,N_22226,N_22712);
or U22897 (N_22897,N_22544,N_22269);
nand U22898 (N_22898,N_22223,N_22699);
or U22899 (N_22899,N_22207,N_21857);
xnor U22900 (N_22900,N_21867,N_21706);
nand U22901 (N_22901,N_22393,N_22688);
nor U22902 (N_22902,N_22465,N_22189);
nand U22903 (N_22903,N_22464,N_22623);
and U22904 (N_22904,N_21873,N_21625);
or U22905 (N_22905,N_22026,N_22767);
or U22906 (N_22906,N_22488,N_21630);
and U22907 (N_22907,N_21802,N_21936);
nand U22908 (N_22908,N_22472,N_22188);
nor U22909 (N_22909,N_21790,N_21747);
nand U22910 (N_22910,N_22323,N_21769);
xnor U22911 (N_22911,N_22174,N_22199);
and U22912 (N_22912,N_22633,N_22107);
xor U22913 (N_22913,N_22265,N_22255);
nor U22914 (N_22914,N_21626,N_22073);
or U22915 (N_22915,N_21679,N_21982);
nand U22916 (N_22916,N_21871,N_21963);
and U22917 (N_22917,N_21923,N_22612);
or U22918 (N_22918,N_21861,N_22186);
nor U22919 (N_22919,N_22164,N_22132);
xor U22920 (N_22920,N_22277,N_22703);
and U22921 (N_22921,N_22631,N_22710);
and U22922 (N_22922,N_21829,N_21967);
or U22923 (N_22923,N_21824,N_22736);
nand U22924 (N_22924,N_22030,N_21917);
nor U22925 (N_22925,N_22118,N_21981);
nor U22926 (N_22926,N_21777,N_22192);
nand U22927 (N_22927,N_22123,N_21697);
nor U22928 (N_22928,N_22175,N_21954);
nor U22929 (N_22929,N_21773,N_22156);
xnor U22930 (N_22930,N_21787,N_22610);
nor U22931 (N_22931,N_21905,N_22745);
nor U22932 (N_22932,N_21945,N_22496);
nor U22933 (N_22933,N_21667,N_21803);
xnor U22934 (N_22934,N_21840,N_21972);
xor U22935 (N_22935,N_22485,N_21784);
nor U22936 (N_22936,N_21920,N_22691);
or U22937 (N_22937,N_22366,N_22385);
nand U22938 (N_22938,N_22062,N_22741);
xnor U22939 (N_22939,N_21695,N_22235);
nand U22940 (N_22940,N_22774,N_22743);
xnor U22941 (N_22941,N_21922,N_22053);
nand U22942 (N_22942,N_21793,N_21789);
nand U22943 (N_22943,N_22074,N_22545);
nand U22944 (N_22944,N_21885,N_22288);
and U22945 (N_22945,N_22510,N_22084);
nand U22946 (N_22946,N_22278,N_22139);
nand U22947 (N_22947,N_22486,N_21774);
nand U22948 (N_22948,N_21612,N_21894);
nand U22949 (N_22949,N_21644,N_22463);
nand U22950 (N_22950,N_21615,N_22602);
or U22951 (N_22951,N_21713,N_22142);
xor U22952 (N_22952,N_21704,N_22701);
xnor U22953 (N_22953,N_21849,N_21942);
and U22954 (N_22954,N_22733,N_22136);
or U22955 (N_22955,N_22780,N_22363);
nand U22956 (N_22956,N_22532,N_22274);
and U22957 (N_22957,N_22033,N_21969);
and U22958 (N_22958,N_22652,N_22259);
nor U22959 (N_22959,N_22558,N_22447);
xnor U22960 (N_22960,N_22783,N_22513);
and U22961 (N_22961,N_21903,N_22459);
nand U22962 (N_22962,N_22738,N_22249);
nand U22963 (N_22963,N_21692,N_21729);
nand U22964 (N_22964,N_21681,N_22417);
and U22965 (N_22965,N_21865,N_22209);
nand U22966 (N_22966,N_22285,N_21724);
and U22967 (N_22967,N_21908,N_21759);
nand U22968 (N_22968,N_22215,N_21937);
or U22969 (N_22969,N_21701,N_22297);
xor U22970 (N_22970,N_22351,N_21788);
nand U22971 (N_22971,N_22538,N_22605);
nand U22972 (N_22972,N_21689,N_22324);
xor U22973 (N_22973,N_22109,N_22098);
nor U22974 (N_22974,N_22617,N_22122);
xor U22975 (N_22975,N_22144,N_22531);
nand U22976 (N_22976,N_22755,N_22706);
nor U22977 (N_22977,N_21627,N_22428);
nand U22978 (N_22978,N_22495,N_21846);
nand U22979 (N_22979,N_22114,N_22355);
and U22980 (N_22980,N_21607,N_22615);
or U22981 (N_22981,N_21673,N_21636);
xor U22982 (N_22982,N_21960,N_21900);
xnor U22983 (N_22983,N_22568,N_21820);
xor U22984 (N_22984,N_22409,N_22566);
nor U22985 (N_22985,N_22275,N_22487);
and U22986 (N_22986,N_22625,N_21655);
xor U22987 (N_22987,N_22438,N_22036);
and U22988 (N_22988,N_21768,N_21749);
nor U22989 (N_22989,N_22674,N_22231);
nand U22990 (N_22990,N_22178,N_21799);
xor U22991 (N_22991,N_22758,N_22448);
or U22992 (N_22992,N_21702,N_22127);
nor U22993 (N_22993,N_21637,N_22567);
nor U22994 (N_22994,N_21949,N_21640);
and U22995 (N_22995,N_22502,N_21940);
nor U22996 (N_22996,N_21955,N_22197);
or U22997 (N_22997,N_21653,N_22088);
xnor U22998 (N_22998,N_22013,N_22796);
and U22999 (N_22999,N_22613,N_21601);
and U23000 (N_23000,N_22167,N_22191);
and U23001 (N_23001,N_22398,N_22311);
nor U23002 (N_23002,N_22070,N_21966);
nor U23003 (N_23003,N_22651,N_22508);
and U23004 (N_23004,N_22518,N_21893);
nand U23005 (N_23005,N_21854,N_22411);
and U23006 (N_23006,N_22593,N_22667);
nor U23007 (N_23007,N_22342,N_21751);
nand U23008 (N_23008,N_22395,N_21842);
nor U23009 (N_23009,N_22450,N_22046);
nand U23010 (N_23010,N_22024,N_22694);
nor U23011 (N_23011,N_22552,N_22404);
nor U23012 (N_23012,N_21719,N_21792);
and U23013 (N_23013,N_22639,N_22316);
and U23014 (N_23014,N_21932,N_22064);
nand U23015 (N_23015,N_22433,N_22019);
or U23016 (N_23016,N_22754,N_22782);
nor U23017 (N_23017,N_21677,N_21752);
or U23018 (N_23018,N_22541,N_22252);
and U23019 (N_23019,N_22799,N_22427);
and U23020 (N_23020,N_22350,N_21864);
and U23021 (N_23021,N_22536,N_21608);
and U23022 (N_23022,N_21735,N_22596);
nor U23023 (N_23023,N_22760,N_21797);
nor U23024 (N_23024,N_21696,N_21712);
nand U23025 (N_23025,N_22099,N_22470);
xor U23026 (N_23026,N_22262,N_21869);
nor U23027 (N_23027,N_21736,N_22150);
nand U23028 (N_23028,N_22266,N_21807);
xor U23029 (N_23029,N_21847,N_21939);
and U23030 (N_23030,N_22002,N_22636);
nand U23031 (N_23031,N_22528,N_22216);
or U23032 (N_23032,N_22068,N_22159);
nand U23033 (N_23033,N_21938,N_22468);
and U23034 (N_23034,N_22784,N_22618);
or U23035 (N_23035,N_22682,N_22374);
nand U23036 (N_23036,N_21678,N_21983);
or U23037 (N_23037,N_22790,N_21974);
and U23038 (N_23038,N_22590,N_22251);
nor U23039 (N_23039,N_22607,N_22290);
xor U23040 (N_23040,N_21986,N_22145);
nor U23041 (N_23041,N_21964,N_22453);
nor U23042 (N_23042,N_21815,N_21614);
or U23043 (N_23043,N_22700,N_21670);
and U23044 (N_23044,N_22579,N_22125);
nor U23045 (N_23045,N_22437,N_22090);
nor U23046 (N_23046,N_22110,N_22535);
nand U23047 (N_23047,N_22133,N_22480);
nor U23048 (N_23048,N_22478,N_22534);
and U23049 (N_23049,N_22603,N_22103);
or U23050 (N_23050,N_22065,N_22202);
nand U23051 (N_23051,N_21962,N_22009);
nor U23052 (N_23052,N_22578,N_22031);
nor U23053 (N_23053,N_22509,N_21665);
nand U23054 (N_23054,N_21746,N_21993);
or U23055 (N_23055,N_21693,N_22348);
nor U23056 (N_23056,N_21811,N_22183);
or U23057 (N_23057,N_22237,N_21810);
nor U23058 (N_23058,N_22388,N_21848);
and U23059 (N_23059,N_22135,N_22184);
or U23060 (N_23060,N_22616,N_22365);
nor U23061 (N_23061,N_22671,N_21652);
nor U23062 (N_23062,N_21909,N_21958);
and U23063 (N_23063,N_21907,N_22224);
nor U23064 (N_23064,N_22446,N_22078);
xor U23065 (N_23065,N_22134,N_21911);
or U23066 (N_23066,N_22006,N_22551);
nand U23067 (N_23067,N_21934,N_21783);
nand U23068 (N_23068,N_22379,N_22321);
and U23069 (N_23069,N_22238,N_22662);
and U23070 (N_23070,N_22797,N_21875);
and U23071 (N_23071,N_22045,N_22349);
nor U23072 (N_23072,N_22330,N_22550);
nor U23073 (N_23073,N_21728,N_22339);
xnor U23074 (N_23074,N_22506,N_22239);
or U23075 (N_23075,N_22021,N_21887);
nand U23076 (N_23076,N_21707,N_21646);
nor U23077 (N_23077,N_22268,N_21760);
xnor U23078 (N_23078,N_21668,N_22236);
nor U23079 (N_23079,N_22273,N_22298);
or U23080 (N_23080,N_22512,N_22672);
nor U23081 (N_23081,N_22559,N_21828);
nand U23082 (N_23082,N_21919,N_21879);
and U23083 (N_23083,N_21690,N_21726);
and U23084 (N_23084,N_22377,N_22214);
nand U23085 (N_23085,N_22734,N_22729);
and U23086 (N_23086,N_22461,N_22709);
nand U23087 (N_23087,N_21613,N_22442);
xnor U23088 (N_23088,N_21813,N_22449);
xor U23089 (N_23089,N_21669,N_21992);
and U23090 (N_23090,N_22751,N_21632);
nor U23091 (N_23091,N_22158,N_22015);
and U23092 (N_23092,N_22648,N_22659);
xor U23093 (N_23093,N_22412,N_22430);
xor U23094 (N_23094,N_22663,N_21800);
nand U23095 (N_23095,N_22032,N_22530);
nor U23096 (N_23096,N_22647,N_21804);
nand U23097 (N_23097,N_22786,N_22329);
and U23098 (N_23098,N_22757,N_22511);
or U23099 (N_23099,N_21860,N_22182);
or U23100 (N_23100,N_22283,N_21927);
and U23101 (N_23101,N_21662,N_21647);
nand U23102 (N_23102,N_22517,N_21779);
or U23103 (N_23103,N_22034,N_22205);
nand U23104 (N_23104,N_22381,N_22681);
and U23105 (N_23105,N_21691,N_21826);
and U23106 (N_23106,N_22308,N_22059);
or U23107 (N_23107,N_22091,N_22725);
nor U23108 (N_23108,N_22769,N_21889);
xor U23109 (N_23109,N_21785,N_21611);
nor U23110 (N_23110,N_22773,N_22505);
xnor U23111 (N_23111,N_22764,N_22153);
and U23112 (N_23112,N_22650,N_22529);
xor U23113 (N_23113,N_22435,N_21798);
or U23114 (N_23114,N_22299,N_21766);
or U23115 (N_23115,N_21859,N_22358);
nor U23116 (N_23116,N_22737,N_22018);
or U23117 (N_23117,N_21845,N_22229);
or U23118 (N_23118,N_21622,N_21880);
or U23119 (N_23119,N_22225,N_22657);
or U23120 (N_23120,N_22160,N_22335);
nor U23121 (N_23121,N_22514,N_22772);
nand U23122 (N_23122,N_22527,N_22471);
and U23123 (N_23123,N_22169,N_22577);
nand U23124 (N_23124,N_22727,N_22312);
nand U23125 (N_23125,N_22732,N_22242);
nand U23126 (N_23126,N_22785,N_22455);
or U23127 (N_23127,N_21947,N_22309);
nor U23128 (N_23128,N_22027,N_21755);
or U23129 (N_23129,N_22763,N_22359);
xor U23130 (N_23130,N_21621,N_22272);
or U23131 (N_23131,N_21910,N_22481);
or U23132 (N_23132,N_22479,N_22119);
or U23133 (N_23133,N_22436,N_22166);
xnor U23134 (N_23134,N_21674,N_22423);
xnor U23135 (N_23135,N_22597,N_22346);
nand U23136 (N_23136,N_22687,N_21657);
or U23137 (N_23137,N_22565,N_21744);
and U23138 (N_23138,N_21600,N_21956);
nor U23139 (N_23139,N_22645,N_21618);
or U23140 (N_23140,N_22198,N_22102);
nand U23141 (N_23141,N_22044,N_22391);
nor U23142 (N_23142,N_22686,N_21838);
or U23143 (N_23143,N_21998,N_21682);
xnor U23144 (N_23144,N_22105,N_21818);
xor U23145 (N_23145,N_22260,N_21822);
or U23146 (N_23146,N_22515,N_22322);
nor U23147 (N_23147,N_22354,N_22220);
and U23148 (N_23148,N_22356,N_21650);
and U23149 (N_23149,N_22594,N_22775);
or U23150 (N_23150,N_22599,N_21892);
xor U23151 (N_23151,N_21772,N_22204);
and U23152 (N_23152,N_22608,N_21764);
nor U23153 (N_23153,N_22685,N_22452);
and U23154 (N_23154,N_22116,N_21931);
xnor U23155 (N_23155,N_22173,N_22143);
nor U23156 (N_23156,N_21757,N_21676);
nand U23157 (N_23157,N_21995,N_22331);
xor U23158 (N_23158,N_22575,N_22085);
nand U23159 (N_23159,N_22576,N_22294);
and U23160 (N_23160,N_22646,N_21700);
or U23161 (N_23161,N_22328,N_21906);
nor U23162 (N_23162,N_22161,N_22628);
and U23163 (N_23163,N_21740,N_22759);
and U23164 (N_23164,N_22384,N_22336);
or U23165 (N_23165,N_22580,N_22043);
or U23166 (N_23166,N_22217,N_21671);
nand U23167 (N_23167,N_21753,N_21872);
or U23168 (N_23168,N_22664,N_22157);
nand U23169 (N_23169,N_22362,N_22611);
nand U23170 (N_23170,N_21727,N_22600);
or U23171 (N_23171,N_21725,N_22677);
nand U23172 (N_23172,N_22492,N_22146);
and U23173 (N_23173,N_21610,N_21870);
xnor U23174 (N_23174,N_21722,N_22286);
and U23175 (N_23175,N_22332,N_22563);
and U23176 (N_23176,N_22724,N_21786);
or U23177 (N_23177,N_22000,N_21738);
nor U23178 (N_23178,N_22668,N_22619);
xor U23179 (N_23179,N_22128,N_21988);
and U23180 (N_23180,N_22306,N_22595);
nor U23181 (N_23181,N_22632,N_21620);
or U23182 (N_23182,N_21912,N_21685);
and U23183 (N_23183,N_21989,N_22720);
nand U23184 (N_23184,N_22140,N_21796);
nor U23185 (N_23185,N_21990,N_21619);
nor U23186 (N_23186,N_22564,N_21841);
nor U23187 (N_23187,N_22670,N_22357);
nand U23188 (N_23188,N_21767,N_22474);
and U23189 (N_23189,N_22179,N_21778);
or U23190 (N_23190,N_22292,N_22170);
xnor U23191 (N_23191,N_22240,N_21883);
nor U23192 (N_23192,N_22719,N_22028);
xnor U23193 (N_23193,N_22347,N_22753);
nor U23194 (N_23194,N_22747,N_22271);
nor U23195 (N_23195,N_22705,N_21605);
nor U23196 (N_23196,N_22243,N_22106);
nor U23197 (N_23197,N_22315,N_22016);
nand U23198 (N_23198,N_22644,N_22200);
nor U23199 (N_23199,N_22234,N_22011);
xnor U23200 (N_23200,N_22660,N_22629);
nand U23201 (N_23201,N_22327,N_22372);
xor U23202 (N_23202,N_22115,N_22638);
xnor U23203 (N_23203,N_22425,N_22748);
nand U23204 (N_23204,N_22022,N_22794);
xor U23205 (N_23205,N_22477,N_22598);
or U23206 (N_23206,N_22410,N_22444);
nor U23207 (N_23207,N_22586,N_22606);
nor U23208 (N_23208,N_22232,N_21634);
xor U23209 (N_23209,N_22707,N_21775);
nand U23210 (N_23210,N_22525,N_22498);
nor U23211 (N_23211,N_21899,N_21801);
or U23212 (N_23212,N_22475,N_22466);
xnor U23213 (N_23213,N_22124,N_21991);
nand U23214 (N_23214,N_22076,N_21973);
or U23215 (N_23215,N_22640,N_21742);
xnor U23216 (N_23216,N_22702,N_21961);
xnor U23217 (N_23217,N_21951,N_22370);
nand U23218 (N_23218,N_22284,N_22071);
xnor U23219 (N_23219,N_21795,N_22561);
or U23220 (N_23220,N_22573,N_22258);
nor U23221 (N_23221,N_22360,N_22054);
and U23222 (N_23222,N_22364,N_22250);
nor U23223 (N_23223,N_22003,N_22310);
or U23224 (N_23224,N_22499,N_22126);
and U23225 (N_23225,N_22176,N_22655);
nand U23226 (N_23226,N_22690,N_22462);
nor U23227 (N_23227,N_22524,N_22405);
nor U23228 (N_23228,N_22519,N_22386);
xor U23229 (N_23229,N_22165,N_21609);
nor U23230 (N_23230,N_22476,N_21816);
xnor U23231 (N_23231,N_22554,N_22041);
nor U23232 (N_23232,N_22267,N_22752);
xor U23233 (N_23233,N_22121,N_21733);
xor U23234 (N_23234,N_21762,N_22291);
nor U23235 (N_23235,N_21731,N_21718);
xnor U23236 (N_23236,N_21806,N_22113);
xor U23237 (N_23237,N_22079,N_22654);
and U23238 (N_23238,N_22503,N_21975);
xnor U23239 (N_23239,N_21855,N_21717);
xnor U23240 (N_23240,N_22408,N_22658);
nor U23241 (N_23241,N_22708,N_21836);
nand U23242 (N_23242,N_21944,N_21862);
or U23243 (N_23243,N_21834,N_22281);
or U23244 (N_23244,N_22684,N_21863);
or U23245 (N_23245,N_22211,N_21904);
nand U23246 (N_23246,N_21698,N_22781);
nand U23247 (N_23247,N_22744,N_21926);
nor U23248 (N_23248,N_21971,N_22722);
and U23249 (N_23249,N_21754,N_21781);
nand U23250 (N_23250,N_21888,N_22087);
or U23251 (N_23251,N_21925,N_22047);
or U23252 (N_23252,N_22083,N_22320);
nand U23253 (N_23253,N_22418,N_22080);
xor U23254 (N_23254,N_22403,N_22637);
xnor U23255 (N_23255,N_22338,N_21661);
and U23256 (N_23256,N_22494,N_22673);
or U23257 (N_23257,N_21823,N_22361);
nand U23258 (N_23258,N_22042,N_22172);
xor U23259 (N_23259,N_22570,N_22641);
and U23260 (N_23260,N_22375,N_22185);
and U23261 (N_23261,N_22614,N_21666);
nand U23262 (N_23262,N_21890,N_22795);
or U23263 (N_23263,N_22353,N_22583);
and U23264 (N_23264,N_22037,N_22679);
nor U23265 (N_23265,N_22007,N_21782);
nor U23266 (N_23266,N_22431,N_21898);
nand U23267 (N_23267,N_22307,N_21680);
or U23268 (N_23268,N_22440,N_22313);
or U23269 (N_23269,N_22390,N_22222);
xor U23270 (N_23270,N_22293,N_22380);
xor U23271 (N_23271,N_22584,N_21687);
or U23272 (N_23272,N_21602,N_22750);
or U23273 (N_23273,N_22522,N_22556);
nor U23274 (N_23274,N_22768,N_22131);
or U23275 (N_23275,N_22761,N_22063);
nand U23276 (N_23276,N_21737,N_22432);
nor U23277 (N_23277,N_22592,N_21628);
and U23278 (N_23278,N_21876,N_22334);
nor U23279 (N_23279,N_22129,N_21663);
and U23280 (N_23280,N_22296,N_21851);
xor U23281 (N_23281,N_22001,N_21976);
xnor U23282 (N_23282,N_21878,N_22560);
nand U23283 (N_23283,N_22521,N_22458);
nand U23284 (N_23284,N_22072,N_22218);
nor U23285 (N_23285,N_21624,N_22352);
and U23286 (N_23286,N_22038,N_22497);
nand U23287 (N_23287,N_21831,N_22152);
nand U23288 (N_23288,N_22693,N_21852);
xor U23289 (N_23289,N_22624,N_22689);
and U23290 (N_23290,N_22739,N_21716);
xor U23291 (N_23291,N_22270,N_22020);
and U23292 (N_23292,N_22343,N_21987);
and U23293 (N_23293,N_21629,N_21809);
or U23294 (N_23294,N_22798,N_21603);
and U23295 (N_23295,N_22396,N_22039);
and U23296 (N_23296,N_21756,N_22721);
nor U23297 (N_23297,N_21604,N_22376);
nand U23298 (N_23298,N_22227,N_21921);
and U23299 (N_23299,N_22301,N_21714);
or U23300 (N_23300,N_22154,N_21660);
xor U23301 (N_23301,N_22714,N_21950);
nand U23302 (N_23302,N_22213,N_22208);
nor U23303 (N_23303,N_22626,N_22230);
nand U23304 (N_23304,N_22451,N_21709);
and U23305 (N_23305,N_21978,N_21924);
nor U23306 (N_23306,N_22081,N_21617);
and U23307 (N_23307,N_22177,N_21664);
and U23308 (N_23308,N_22557,N_22665);
or U23309 (N_23309,N_22771,N_22533);
xnor U23310 (N_23310,N_22014,N_22656);
xor U23311 (N_23311,N_22373,N_21891);
and U23312 (N_23312,N_21968,N_22245);
nor U23313 (N_23313,N_22634,N_22181);
and U23314 (N_23314,N_22572,N_22052);
and U23315 (N_23315,N_21881,N_21805);
and U23316 (N_23316,N_21683,N_22399);
xnor U23317 (N_23317,N_21641,N_22100);
and U23318 (N_23318,N_22378,N_22501);
xnor U23319 (N_23319,N_22017,N_22581);
or U23320 (N_23320,N_22715,N_21659);
and U23321 (N_23321,N_22295,N_22420);
and U23322 (N_23322,N_22520,N_22289);
nand U23323 (N_23323,N_22248,N_22482);
or U23324 (N_23324,N_22058,N_22212);
nor U23325 (N_23325,N_22749,N_22246);
or U23326 (N_23326,N_21821,N_22445);
nor U23327 (N_23327,N_22489,N_21866);
nor U23328 (N_23328,N_22740,N_21996);
xor U23329 (N_23329,N_22147,N_21853);
nand U23330 (N_23330,N_21763,N_22210);
or U23331 (N_23331,N_22089,N_22547);
nor U23332 (N_23332,N_22130,N_22149);
nand U23333 (N_23333,N_22539,N_22562);
nor U23334 (N_23334,N_21884,N_22137);
xor U23335 (N_23335,N_21739,N_21928);
nor U23336 (N_23336,N_22621,N_22490);
nor U23337 (N_23337,N_21761,N_22148);
xor U23338 (N_23338,N_21686,N_22723);
xor U23339 (N_23339,N_22735,N_21980);
xor U23340 (N_23340,N_22012,N_22120);
nand U23341 (N_23341,N_21758,N_22756);
nand U23342 (N_23342,N_21997,N_21741);
nor U23343 (N_23343,N_22516,N_22049);
or U23344 (N_23344,N_22195,N_22555);
nor U23345 (N_23345,N_22097,N_22264);
and U23346 (N_23346,N_21710,N_22048);
or U23347 (N_23347,N_21858,N_21819);
nor U23348 (N_23348,N_21916,N_22791);
nor U23349 (N_23349,N_21814,N_21765);
xnor U23350 (N_23350,N_22155,N_21929);
and U23351 (N_23351,N_22469,N_22261);
or U23352 (N_23352,N_21748,N_21850);
xnor U23353 (N_23353,N_21642,N_22669);
and U23354 (N_23354,N_22069,N_21672);
or U23355 (N_23355,N_22101,N_22424);
or U23356 (N_23356,N_22051,N_22718);
and U23357 (N_23357,N_22543,N_22067);
nand U23358 (N_23358,N_21915,N_22086);
nand U23359 (N_23359,N_21794,N_22601);
or U23360 (N_23360,N_21770,N_22630);
nor U23361 (N_23361,N_22776,N_22303);
and U23362 (N_23362,N_22325,N_22190);
xnor U23363 (N_23363,N_22683,N_22666);
nor U23364 (N_23364,N_22697,N_22540);
nand U23365 (N_23365,N_21699,N_22302);
nor U23366 (N_23366,N_22203,N_22319);
or U23367 (N_23367,N_22023,N_22077);
and U23368 (N_23368,N_21882,N_22263);
or U23369 (N_23369,N_22484,N_22589);
nand U23370 (N_23370,N_22415,N_22635);
nand U23371 (N_23371,N_22620,N_21985);
and U23372 (N_23372,N_21837,N_22168);
xor U23373 (N_23373,N_21830,N_22400);
nor U23374 (N_23374,N_21645,N_21616);
and U23375 (N_23375,N_22526,N_21776);
nor U23376 (N_23376,N_22096,N_22317);
nor U23377 (N_23377,N_22588,N_22344);
or U23378 (N_23378,N_22345,N_22504);
or U23379 (N_23379,N_21654,N_21953);
and U23380 (N_23380,N_22766,N_22426);
or U23381 (N_23381,N_21825,N_22585);
nand U23382 (N_23382,N_21952,N_21643);
nor U23383 (N_23383,N_22108,N_22454);
nor U23384 (N_23384,N_21633,N_22367);
and U23385 (N_23385,N_22460,N_22333);
nand U23386 (N_23386,N_22341,N_22075);
or U23387 (N_23387,N_22419,N_22421);
or U23388 (N_23388,N_21839,N_22676);
xor U23389 (N_23389,N_21999,N_21684);
nand U23390 (N_23390,N_22368,N_21856);
nor U23391 (N_23391,N_22392,N_22256);
nand U23392 (N_23392,N_21734,N_22728);
nand U23393 (N_23393,N_22731,N_22241);
and U23394 (N_23394,N_22643,N_22549);
xor U23395 (N_23395,N_21817,N_21623);
nand U23396 (N_23396,N_22569,N_22413);
nand U23397 (N_23397,N_22382,N_21715);
or U23398 (N_23398,N_22171,N_21656);
and U23399 (N_23399,N_22253,N_22257);
and U23400 (N_23400,N_21796,N_22382);
xor U23401 (N_23401,N_21966,N_22303);
xor U23402 (N_23402,N_22316,N_21843);
xnor U23403 (N_23403,N_22050,N_22480);
and U23404 (N_23404,N_21718,N_22062);
xnor U23405 (N_23405,N_22112,N_22263);
and U23406 (N_23406,N_22562,N_21795);
xor U23407 (N_23407,N_21672,N_21782);
or U23408 (N_23408,N_22640,N_21982);
nor U23409 (N_23409,N_22175,N_22579);
or U23410 (N_23410,N_22632,N_21928);
nor U23411 (N_23411,N_21982,N_22449);
nand U23412 (N_23412,N_22496,N_22342);
xor U23413 (N_23413,N_22436,N_21956);
and U23414 (N_23414,N_22174,N_22693);
xor U23415 (N_23415,N_22687,N_22348);
and U23416 (N_23416,N_22652,N_21826);
nor U23417 (N_23417,N_22299,N_22600);
or U23418 (N_23418,N_22573,N_22426);
or U23419 (N_23419,N_22360,N_22775);
nand U23420 (N_23420,N_22341,N_22032);
and U23421 (N_23421,N_22471,N_21758);
or U23422 (N_23422,N_22773,N_22716);
nand U23423 (N_23423,N_22783,N_21613);
or U23424 (N_23424,N_22703,N_22751);
xor U23425 (N_23425,N_22233,N_22132);
or U23426 (N_23426,N_22165,N_21861);
nor U23427 (N_23427,N_21718,N_22009);
nor U23428 (N_23428,N_21902,N_21605);
and U23429 (N_23429,N_22166,N_22341);
nor U23430 (N_23430,N_21819,N_22625);
xnor U23431 (N_23431,N_22274,N_22594);
or U23432 (N_23432,N_22661,N_22102);
or U23433 (N_23433,N_22260,N_21707);
xnor U23434 (N_23434,N_22497,N_22711);
nor U23435 (N_23435,N_21706,N_21603);
or U23436 (N_23436,N_21970,N_21745);
xor U23437 (N_23437,N_21601,N_22747);
nand U23438 (N_23438,N_22208,N_22270);
nor U23439 (N_23439,N_21828,N_22576);
xnor U23440 (N_23440,N_22649,N_22281);
nand U23441 (N_23441,N_22520,N_21979);
nand U23442 (N_23442,N_21982,N_22335);
and U23443 (N_23443,N_22118,N_22412);
nand U23444 (N_23444,N_21856,N_22285);
and U23445 (N_23445,N_21623,N_22206);
xor U23446 (N_23446,N_22523,N_22353);
or U23447 (N_23447,N_21612,N_22583);
and U23448 (N_23448,N_22231,N_21605);
xnor U23449 (N_23449,N_22179,N_22791);
nor U23450 (N_23450,N_21702,N_21724);
and U23451 (N_23451,N_22310,N_22767);
xnor U23452 (N_23452,N_22318,N_22005);
and U23453 (N_23453,N_22595,N_21849);
and U23454 (N_23454,N_21794,N_21915);
and U23455 (N_23455,N_22577,N_22504);
xor U23456 (N_23456,N_22300,N_22317);
or U23457 (N_23457,N_22266,N_21766);
or U23458 (N_23458,N_21886,N_21678);
or U23459 (N_23459,N_21820,N_22261);
or U23460 (N_23460,N_21735,N_22204);
xor U23461 (N_23461,N_22111,N_21753);
and U23462 (N_23462,N_21996,N_21614);
xor U23463 (N_23463,N_22005,N_22239);
xor U23464 (N_23464,N_21654,N_22509);
and U23465 (N_23465,N_22251,N_22677);
nand U23466 (N_23466,N_22410,N_21885);
nand U23467 (N_23467,N_22240,N_22363);
nand U23468 (N_23468,N_22154,N_22331);
nand U23469 (N_23469,N_22080,N_22558);
or U23470 (N_23470,N_22344,N_22024);
nand U23471 (N_23471,N_22354,N_22143);
xor U23472 (N_23472,N_22617,N_21664);
xor U23473 (N_23473,N_22730,N_22548);
xnor U23474 (N_23474,N_21736,N_21660);
and U23475 (N_23475,N_21784,N_22465);
nor U23476 (N_23476,N_22590,N_21681);
and U23477 (N_23477,N_21639,N_22653);
xor U23478 (N_23478,N_22495,N_22476);
xnor U23479 (N_23479,N_22373,N_22695);
nand U23480 (N_23480,N_22098,N_22397);
xor U23481 (N_23481,N_21724,N_21689);
and U23482 (N_23482,N_21694,N_22263);
nor U23483 (N_23483,N_22515,N_22721);
or U23484 (N_23484,N_22528,N_22047);
and U23485 (N_23485,N_21763,N_22492);
and U23486 (N_23486,N_21604,N_21914);
or U23487 (N_23487,N_21841,N_21620);
nor U23488 (N_23488,N_22602,N_22343);
nor U23489 (N_23489,N_22651,N_22370);
or U23490 (N_23490,N_22763,N_21620);
xnor U23491 (N_23491,N_22548,N_21842);
or U23492 (N_23492,N_22656,N_22109);
and U23493 (N_23493,N_21761,N_21917);
nand U23494 (N_23494,N_21850,N_21818);
and U23495 (N_23495,N_21944,N_21670);
nand U23496 (N_23496,N_21940,N_22486);
nor U23497 (N_23497,N_22594,N_22722);
and U23498 (N_23498,N_21691,N_22234);
and U23499 (N_23499,N_22773,N_22268);
or U23500 (N_23500,N_22178,N_22369);
or U23501 (N_23501,N_22498,N_22324);
or U23502 (N_23502,N_21616,N_22192);
nor U23503 (N_23503,N_22581,N_22775);
or U23504 (N_23504,N_22277,N_22513);
or U23505 (N_23505,N_22048,N_22230);
xor U23506 (N_23506,N_22302,N_22555);
or U23507 (N_23507,N_22677,N_22132);
nand U23508 (N_23508,N_21953,N_21797);
xor U23509 (N_23509,N_22716,N_22097);
xor U23510 (N_23510,N_22150,N_22568);
nand U23511 (N_23511,N_22454,N_21855);
xnor U23512 (N_23512,N_22134,N_22692);
or U23513 (N_23513,N_21894,N_22138);
nor U23514 (N_23514,N_21978,N_22390);
or U23515 (N_23515,N_21952,N_22424);
xnor U23516 (N_23516,N_22773,N_22060);
or U23517 (N_23517,N_22609,N_22592);
nand U23518 (N_23518,N_22731,N_22612);
nor U23519 (N_23519,N_22616,N_22332);
and U23520 (N_23520,N_22523,N_22416);
nand U23521 (N_23521,N_22138,N_22454);
nor U23522 (N_23522,N_22291,N_22707);
nor U23523 (N_23523,N_22355,N_22730);
nor U23524 (N_23524,N_21671,N_21622);
nand U23525 (N_23525,N_22083,N_22679);
and U23526 (N_23526,N_22640,N_22028);
nor U23527 (N_23527,N_21883,N_22161);
or U23528 (N_23528,N_22002,N_22232);
nor U23529 (N_23529,N_22098,N_22033);
xor U23530 (N_23530,N_22187,N_22328);
and U23531 (N_23531,N_22571,N_22443);
or U23532 (N_23532,N_22789,N_22658);
and U23533 (N_23533,N_21612,N_22412);
or U23534 (N_23534,N_22142,N_22284);
or U23535 (N_23535,N_21754,N_22228);
or U23536 (N_23536,N_21948,N_22315);
nand U23537 (N_23537,N_22162,N_22490);
xnor U23538 (N_23538,N_21796,N_22456);
nor U23539 (N_23539,N_22659,N_22516);
and U23540 (N_23540,N_22593,N_22008);
nand U23541 (N_23541,N_21701,N_22493);
or U23542 (N_23542,N_22137,N_22450);
or U23543 (N_23543,N_22086,N_21719);
and U23544 (N_23544,N_21824,N_22136);
nor U23545 (N_23545,N_22538,N_21937);
nand U23546 (N_23546,N_22280,N_22202);
nor U23547 (N_23547,N_21884,N_21811);
and U23548 (N_23548,N_21663,N_21616);
xor U23549 (N_23549,N_22024,N_22580);
nor U23550 (N_23550,N_22657,N_22694);
nand U23551 (N_23551,N_22752,N_22637);
or U23552 (N_23552,N_21883,N_22597);
or U23553 (N_23553,N_22514,N_22017);
nand U23554 (N_23554,N_22383,N_22594);
nand U23555 (N_23555,N_22369,N_22706);
nor U23556 (N_23556,N_22041,N_22160);
or U23557 (N_23557,N_22111,N_22739);
nand U23558 (N_23558,N_22044,N_22092);
and U23559 (N_23559,N_22559,N_22581);
nand U23560 (N_23560,N_22554,N_22115);
xnor U23561 (N_23561,N_22158,N_22164);
xor U23562 (N_23562,N_22305,N_22326);
xor U23563 (N_23563,N_22008,N_22537);
nor U23564 (N_23564,N_21601,N_21846);
nand U23565 (N_23565,N_22012,N_22034);
nor U23566 (N_23566,N_22236,N_21870);
and U23567 (N_23567,N_21632,N_22536);
and U23568 (N_23568,N_21780,N_21657);
xor U23569 (N_23569,N_21714,N_21829);
nand U23570 (N_23570,N_21872,N_21900);
or U23571 (N_23571,N_22556,N_22425);
nand U23572 (N_23572,N_22708,N_22140);
nand U23573 (N_23573,N_21749,N_21890);
or U23574 (N_23574,N_22197,N_21918);
or U23575 (N_23575,N_22076,N_21928);
or U23576 (N_23576,N_21899,N_21662);
nor U23577 (N_23577,N_22699,N_22272);
nor U23578 (N_23578,N_22191,N_22648);
nand U23579 (N_23579,N_22274,N_22635);
and U23580 (N_23580,N_21888,N_21870);
nand U23581 (N_23581,N_22520,N_22274);
nand U23582 (N_23582,N_22611,N_22190);
and U23583 (N_23583,N_22452,N_22316);
nand U23584 (N_23584,N_22369,N_22605);
and U23585 (N_23585,N_21900,N_21916);
and U23586 (N_23586,N_21609,N_21678);
and U23587 (N_23587,N_21775,N_22229);
and U23588 (N_23588,N_21735,N_22628);
nand U23589 (N_23589,N_22131,N_22312);
nor U23590 (N_23590,N_22419,N_22080);
xor U23591 (N_23591,N_22019,N_22661);
nand U23592 (N_23592,N_22668,N_22239);
nor U23593 (N_23593,N_22634,N_22579);
and U23594 (N_23594,N_22030,N_22341);
nand U23595 (N_23595,N_22626,N_22656);
and U23596 (N_23596,N_21950,N_22022);
nand U23597 (N_23597,N_22413,N_22253);
and U23598 (N_23598,N_21890,N_22762);
and U23599 (N_23599,N_22355,N_22053);
or U23600 (N_23600,N_22448,N_22449);
or U23601 (N_23601,N_22133,N_22019);
xor U23602 (N_23602,N_21675,N_22304);
nor U23603 (N_23603,N_22660,N_22118);
nand U23604 (N_23604,N_22115,N_21918);
nor U23605 (N_23605,N_21809,N_22280);
nand U23606 (N_23606,N_22181,N_21650);
and U23607 (N_23607,N_21701,N_22002);
or U23608 (N_23608,N_22683,N_22687);
nor U23609 (N_23609,N_22503,N_21885);
nand U23610 (N_23610,N_22624,N_22241);
or U23611 (N_23611,N_22556,N_22755);
xor U23612 (N_23612,N_22260,N_22541);
nand U23613 (N_23613,N_22544,N_22449);
or U23614 (N_23614,N_22666,N_22423);
nor U23615 (N_23615,N_21668,N_21755);
and U23616 (N_23616,N_22690,N_21621);
nor U23617 (N_23617,N_22494,N_22704);
or U23618 (N_23618,N_21709,N_22114);
nor U23619 (N_23619,N_21829,N_22710);
nand U23620 (N_23620,N_22720,N_22169);
or U23621 (N_23621,N_21772,N_22656);
nor U23622 (N_23622,N_22463,N_22655);
nor U23623 (N_23623,N_21970,N_22450);
nand U23624 (N_23624,N_21708,N_21782);
nor U23625 (N_23625,N_22025,N_22384);
nand U23626 (N_23626,N_22555,N_21619);
nor U23627 (N_23627,N_21949,N_22449);
xnor U23628 (N_23628,N_22209,N_22676);
nor U23629 (N_23629,N_21973,N_21835);
nand U23630 (N_23630,N_22761,N_22642);
and U23631 (N_23631,N_22191,N_22719);
or U23632 (N_23632,N_22132,N_22759);
and U23633 (N_23633,N_22639,N_21870);
nor U23634 (N_23634,N_22069,N_22080);
xor U23635 (N_23635,N_21707,N_22497);
and U23636 (N_23636,N_21718,N_21847);
and U23637 (N_23637,N_22624,N_21915);
nor U23638 (N_23638,N_21681,N_22540);
nor U23639 (N_23639,N_22342,N_22794);
or U23640 (N_23640,N_22355,N_21992);
nand U23641 (N_23641,N_21911,N_22642);
xnor U23642 (N_23642,N_21681,N_22308);
nand U23643 (N_23643,N_22198,N_21880);
nand U23644 (N_23644,N_21809,N_21616);
nor U23645 (N_23645,N_21675,N_22411);
xor U23646 (N_23646,N_21756,N_22792);
or U23647 (N_23647,N_22688,N_21853);
nand U23648 (N_23648,N_22284,N_22627);
xnor U23649 (N_23649,N_22707,N_21956);
xor U23650 (N_23650,N_21794,N_21709);
nor U23651 (N_23651,N_21724,N_22562);
xor U23652 (N_23652,N_21915,N_22488);
and U23653 (N_23653,N_22066,N_21966);
or U23654 (N_23654,N_22377,N_21604);
or U23655 (N_23655,N_22111,N_21827);
xnor U23656 (N_23656,N_22457,N_21853);
xnor U23657 (N_23657,N_22493,N_21653);
nor U23658 (N_23658,N_22540,N_22488);
nand U23659 (N_23659,N_22355,N_21688);
or U23660 (N_23660,N_21955,N_21622);
and U23661 (N_23661,N_21661,N_22748);
nor U23662 (N_23662,N_22510,N_22040);
nand U23663 (N_23663,N_22637,N_22042);
and U23664 (N_23664,N_22184,N_22566);
xor U23665 (N_23665,N_22165,N_22632);
nand U23666 (N_23666,N_22778,N_22132);
xor U23667 (N_23667,N_22242,N_22486);
nor U23668 (N_23668,N_22753,N_22401);
or U23669 (N_23669,N_22117,N_22096);
nand U23670 (N_23670,N_22301,N_22327);
or U23671 (N_23671,N_22484,N_21652);
xor U23672 (N_23672,N_21733,N_22263);
nand U23673 (N_23673,N_21753,N_22778);
and U23674 (N_23674,N_21983,N_21961);
nand U23675 (N_23675,N_22011,N_21987);
xor U23676 (N_23676,N_22417,N_22784);
and U23677 (N_23677,N_22135,N_22541);
nand U23678 (N_23678,N_22509,N_22603);
nand U23679 (N_23679,N_21848,N_22315);
and U23680 (N_23680,N_22589,N_21925);
nand U23681 (N_23681,N_22308,N_22547);
and U23682 (N_23682,N_21620,N_22770);
or U23683 (N_23683,N_22216,N_22086);
xor U23684 (N_23684,N_22086,N_21795);
and U23685 (N_23685,N_21907,N_22007);
nand U23686 (N_23686,N_22510,N_21772);
or U23687 (N_23687,N_21829,N_22585);
nand U23688 (N_23688,N_22664,N_22105);
nor U23689 (N_23689,N_22514,N_22679);
nand U23690 (N_23690,N_22344,N_22612);
xnor U23691 (N_23691,N_22070,N_21650);
nand U23692 (N_23692,N_22211,N_22143);
or U23693 (N_23693,N_21612,N_22560);
and U23694 (N_23694,N_22670,N_22345);
or U23695 (N_23695,N_22610,N_22167);
nor U23696 (N_23696,N_22603,N_22318);
nor U23697 (N_23697,N_22146,N_22304);
xnor U23698 (N_23698,N_22329,N_21725);
and U23699 (N_23699,N_21672,N_22453);
nor U23700 (N_23700,N_22152,N_21625);
nor U23701 (N_23701,N_22087,N_22781);
nor U23702 (N_23702,N_22129,N_22640);
nor U23703 (N_23703,N_22011,N_21621);
nand U23704 (N_23704,N_22718,N_21756);
and U23705 (N_23705,N_22091,N_22175);
xnor U23706 (N_23706,N_21941,N_22150);
nand U23707 (N_23707,N_22217,N_22618);
and U23708 (N_23708,N_22406,N_22431);
and U23709 (N_23709,N_22796,N_22735);
nand U23710 (N_23710,N_21929,N_22574);
and U23711 (N_23711,N_22067,N_22775);
and U23712 (N_23712,N_22691,N_22348);
xnor U23713 (N_23713,N_21777,N_22289);
nor U23714 (N_23714,N_22059,N_22378);
xnor U23715 (N_23715,N_21782,N_22365);
nor U23716 (N_23716,N_21884,N_22150);
and U23717 (N_23717,N_22589,N_22721);
nor U23718 (N_23718,N_22627,N_22444);
or U23719 (N_23719,N_22061,N_22534);
and U23720 (N_23720,N_22623,N_22132);
xnor U23721 (N_23721,N_22706,N_22689);
and U23722 (N_23722,N_22779,N_21859);
nor U23723 (N_23723,N_22054,N_21697);
nor U23724 (N_23724,N_22690,N_22382);
xnor U23725 (N_23725,N_22723,N_22407);
nand U23726 (N_23726,N_22348,N_22209);
xor U23727 (N_23727,N_21939,N_22641);
nor U23728 (N_23728,N_22475,N_21830);
or U23729 (N_23729,N_21952,N_22746);
and U23730 (N_23730,N_22589,N_21991);
or U23731 (N_23731,N_22494,N_22404);
nand U23732 (N_23732,N_22367,N_21700);
nor U23733 (N_23733,N_22730,N_22153);
or U23734 (N_23734,N_22297,N_22526);
nand U23735 (N_23735,N_21657,N_21671);
nor U23736 (N_23736,N_22519,N_22568);
nor U23737 (N_23737,N_22522,N_22775);
or U23738 (N_23738,N_22575,N_21766);
or U23739 (N_23739,N_22043,N_21629);
or U23740 (N_23740,N_22420,N_21879);
and U23741 (N_23741,N_21941,N_22582);
nand U23742 (N_23742,N_22253,N_22132);
nand U23743 (N_23743,N_22114,N_21767);
nor U23744 (N_23744,N_21624,N_21762);
xnor U23745 (N_23745,N_22030,N_22502);
nand U23746 (N_23746,N_21788,N_22552);
nand U23747 (N_23747,N_22718,N_22742);
nor U23748 (N_23748,N_22405,N_22076);
nand U23749 (N_23749,N_21905,N_21953);
nor U23750 (N_23750,N_22091,N_21759);
nand U23751 (N_23751,N_22750,N_21674);
xnor U23752 (N_23752,N_22264,N_21973);
nor U23753 (N_23753,N_21826,N_22078);
and U23754 (N_23754,N_21915,N_21902);
nor U23755 (N_23755,N_22697,N_22713);
or U23756 (N_23756,N_22445,N_22464);
nand U23757 (N_23757,N_22674,N_22141);
xnor U23758 (N_23758,N_22527,N_21956);
nand U23759 (N_23759,N_22329,N_22495);
or U23760 (N_23760,N_21755,N_22520);
nor U23761 (N_23761,N_21787,N_21650);
nor U23762 (N_23762,N_22294,N_21760);
or U23763 (N_23763,N_21920,N_21820);
or U23764 (N_23764,N_22101,N_22587);
nand U23765 (N_23765,N_22222,N_21705);
nand U23766 (N_23766,N_22593,N_22505);
or U23767 (N_23767,N_22260,N_22654);
and U23768 (N_23768,N_22089,N_21682);
nor U23769 (N_23769,N_22119,N_21839);
and U23770 (N_23770,N_22034,N_22243);
nand U23771 (N_23771,N_22316,N_22003);
and U23772 (N_23772,N_21617,N_21973);
nor U23773 (N_23773,N_22561,N_22440);
xnor U23774 (N_23774,N_22056,N_22505);
nor U23775 (N_23775,N_22394,N_22201);
and U23776 (N_23776,N_22564,N_22592);
and U23777 (N_23777,N_22519,N_22208);
nand U23778 (N_23778,N_22062,N_21864);
nor U23779 (N_23779,N_21885,N_22192);
or U23780 (N_23780,N_21941,N_21614);
nor U23781 (N_23781,N_22127,N_22084);
nand U23782 (N_23782,N_21848,N_21710);
nand U23783 (N_23783,N_22205,N_21838);
and U23784 (N_23784,N_21988,N_21896);
nor U23785 (N_23785,N_22118,N_22447);
nand U23786 (N_23786,N_21887,N_21650);
and U23787 (N_23787,N_22310,N_21812);
and U23788 (N_23788,N_21795,N_22507);
nand U23789 (N_23789,N_21749,N_22484);
xor U23790 (N_23790,N_22689,N_21924);
or U23791 (N_23791,N_22379,N_21934);
or U23792 (N_23792,N_22651,N_21647);
nor U23793 (N_23793,N_22168,N_22259);
or U23794 (N_23794,N_22706,N_21956);
and U23795 (N_23795,N_21631,N_22568);
xnor U23796 (N_23796,N_21731,N_22560);
nor U23797 (N_23797,N_21648,N_22464);
or U23798 (N_23798,N_22504,N_22366);
or U23799 (N_23799,N_22346,N_22770);
and U23800 (N_23800,N_21689,N_21902);
xnor U23801 (N_23801,N_22521,N_22734);
nor U23802 (N_23802,N_22467,N_22518);
nor U23803 (N_23803,N_22142,N_21888);
and U23804 (N_23804,N_22491,N_22640);
nor U23805 (N_23805,N_22435,N_22003);
nand U23806 (N_23806,N_22173,N_21652);
nand U23807 (N_23807,N_21708,N_21813);
nand U23808 (N_23808,N_22796,N_21961);
and U23809 (N_23809,N_21837,N_22398);
and U23810 (N_23810,N_21696,N_22025);
xor U23811 (N_23811,N_21806,N_22388);
or U23812 (N_23812,N_22618,N_22281);
xnor U23813 (N_23813,N_22417,N_21717);
nor U23814 (N_23814,N_22035,N_22234);
and U23815 (N_23815,N_21761,N_22567);
or U23816 (N_23816,N_21962,N_22627);
nor U23817 (N_23817,N_21626,N_22619);
xnor U23818 (N_23818,N_21776,N_22697);
or U23819 (N_23819,N_21815,N_22163);
xor U23820 (N_23820,N_21948,N_22613);
or U23821 (N_23821,N_21709,N_21990);
nand U23822 (N_23822,N_22047,N_22341);
nor U23823 (N_23823,N_21750,N_22046);
or U23824 (N_23824,N_22786,N_22268);
or U23825 (N_23825,N_21975,N_22555);
xor U23826 (N_23826,N_22300,N_22548);
nor U23827 (N_23827,N_22030,N_22276);
nand U23828 (N_23828,N_22476,N_22381);
and U23829 (N_23829,N_22790,N_22671);
and U23830 (N_23830,N_22576,N_22535);
and U23831 (N_23831,N_22173,N_21806);
xnor U23832 (N_23832,N_21839,N_22176);
or U23833 (N_23833,N_22342,N_22205);
or U23834 (N_23834,N_22669,N_21940);
and U23835 (N_23835,N_21651,N_21706);
or U23836 (N_23836,N_22174,N_22146);
or U23837 (N_23837,N_22368,N_22585);
nor U23838 (N_23838,N_21963,N_21988);
nor U23839 (N_23839,N_22184,N_22266);
nor U23840 (N_23840,N_22760,N_21646);
nor U23841 (N_23841,N_22067,N_22281);
xor U23842 (N_23842,N_22138,N_21660);
nor U23843 (N_23843,N_22791,N_22199);
nand U23844 (N_23844,N_22336,N_21803);
and U23845 (N_23845,N_21701,N_21611);
nor U23846 (N_23846,N_22252,N_22442);
or U23847 (N_23847,N_22781,N_21612);
xnor U23848 (N_23848,N_22417,N_22579);
and U23849 (N_23849,N_21655,N_22282);
nand U23850 (N_23850,N_22167,N_22091);
nor U23851 (N_23851,N_22315,N_22050);
and U23852 (N_23852,N_21850,N_21685);
or U23853 (N_23853,N_22423,N_22569);
or U23854 (N_23854,N_22519,N_21950);
nor U23855 (N_23855,N_22217,N_21833);
nand U23856 (N_23856,N_21866,N_22033);
nor U23857 (N_23857,N_22722,N_22570);
or U23858 (N_23858,N_22001,N_21856);
and U23859 (N_23859,N_22712,N_21715);
nor U23860 (N_23860,N_22147,N_22594);
xor U23861 (N_23861,N_22719,N_22397);
xnor U23862 (N_23862,N_21690,N_22489);
nor U23863 (N_23863,N_21662,N_22260);
nand U23864 (N_23864,N_22164,N_22181);
nand U23865 (N_23865,N_22664,N_21614);
nand U23866 (N_23866,N_22638,N_21784);
and U23867 (N_23867,N_22779,N_22110);
or U23868 (N_23868,N_21749,N_21829);
xor U23869 (N_23869,N_21990,N_22067);
xnor U23870 (N_23870,N_22760,N_22391);
xor U23871 (N_23871,N_22470,N_22148);
nand U23872 (N_23872,N_22383,N_22543);
nand U23873 (N_23873,N_22798,N_22465);
and U23874 (N_23874,N_22073,N_22530);
nor U23875 (N_23875,N_22469,N_22772);
nand U23876 (N_23876,N_22756,N_22230);
xor U23877 (N_23877,N_22160,N_22726);
and U23878 (N_23878,N_22765,N_21798);
xor U23879 (N_23879,N_21671,N_21885);
nor U23880 (N_23880,N_22299,N_21644);
nor U23881 (N_23881,N_22279,N_22436);
and U23882 (N_23882,N_22563,N_22361);
xor U23883 (N_23883,N_21621,N_21958);
nand U23884 (N_23884,N_22436,N_22381);
or U23885 (N_23885,N_21948,N_22366);
nor U23886 (N_23886,N_21601,N_22327);
or U23887 (N_23887,N_22253,N_22321);
xnor U23888 (N_23888,N_22321,N_22648);
and U23889 (N_23889,N_22128,N_22737);
and U23890 (N_23890,N_22067,N_22041);
nor U23891 (N_23891,N_22435,N_22012);
nand U23892 (N_23892,N_22458,N_22577);
xor U23893 (N_23893,N_22188,N_22260);
and U23894 (N_23894,N_22342,N_21829);
nor U23895 (N_23895,N_21912,N_22147);
xor U23896 (N_23896,N_22522,N_22516);
or U23897 (N_23897,N_21997,N_22437);
or U23898 (N_23898,N_22280,N_22763);
xor U23899 (N_23899,N_22450,N_22688);
nor U23900 (N_23900,N_22530,N_21717);
nand U23901 (N_23901,N_21947,N_22441);
nor U23902 (N_23902,N_21964,N_22554);
or U23903 (N_23903,N_21871,N_21833);
nor U23904 (N_23904,N_22304,N_22161);
and U23905 (N_23905,N_21795,N_22217);
nand U23906 (N_23906,N_22575,N_22669);
or U23907 (N_23907,N_22595,N_21946);
and U23908 (N_23908,N_22759,N_22055);
nand U23909 (N_23909,N_22576,N_21908);
nand U23910 (N_23910,N_21920,N_22551);
nor U23911 (N_23911,N_22270,N_22788);
xnor U23912 (N_23912,N_22542,N_22168);
xnor U23913 (N_23913,N_22653,N_22763);
nand U23914 (N_23914,N_21778,N_21879);
nor U23915 (N_23915,N_22257,N_22582);
nand U23916 (N_23916,N_22723,N_21963);
nand U23917 (N_23917,N_21869,N_21706);
or U23918 (N_23918,N_22532,N_22716);
or U23919 (N_23919,N_21614,N_21868);
nor U23920 (N_23920,N_21804,N_22458);
nor U23921 (N_23921,N_21882,N_22455);
and U23922 (N_23922,N_22624,N_21727);
or U23923 (N_23923,N_22704,N_22398);
and U23924 (N_23924,N_22190,N_22639);
or U23925 (N_23925,N_21624,N_21946);
and U23926 (N_23926,N_21877,N_22527);
and U23927 (N_23927,N_22726,N_22531);
and U23928 (N_23928,N_21697,N_22230);
and U23929 (N_23929,N_22076,N_22592);
or U23930 (N_23930,N_22572,N_21870);
nand U23931 (N_23931,N_22309,N_21786);
nor U23932 (N_23932,N_22414,N_21965);
nand U23933 (N_23933,N_22115,N_22160);
xnor U23934 (N_23934,N_22108,N_21939);
and U23935 (N_23935,N_21787,N_22709);
nand U23936 (N_23936,N_21783,N_22305);
nor U23937 (N_23937,N_22204,N_22744);
or U23938 (N_23938,N_22723,N_22215);
or U23939 (N_23939,N_22162,N_22057);
or U23940 (N_23940,N_22669,N_22011);
or U23941 (N_23941,N_22410,N_22087);
nor U23942 (N_23942,N_21794,N_22151);
or U23943 (N_23943,N_21880,N_22666);
nor U23944 (N_23944,N_21787,N_22385);
and U23945 (N_23945,N_21816,N_22206);
xor U23946 (N_23946,N_22382,N_22353);
nor U23947 (N_23947,N_21696,N_21744);
xnor U23948 (N_23948,N_21946,N_22154);
nand U23949 (N_23949,N_22532,N_22188);
nand U23950 (N_23950,N_21621,N_22253);
nand U23951 (N_23951,N_22254,N_21627);
xor U23952 (N_23952,N_22155,N_22426);
and U23953 (N_23953,N_21640,N_22330);
and U23954 (N_23954,N_21877,N_21934);
and U23955 (N_23955,N_22051,N_22076);
nand U23956 (N_23956,N_21951,N_22602);
nand U23957 (N_23957,N_21946,N_22688);
xor U23958 (N_23958,N_22190,N_21790);
or U23959 (N_23959,N_22574,N_22743);
xor U23960 (N_23960,N_21623,N_22165);
nand U23961 (N_23961,N_21902,N_22293);
nor U23962 (N_23962,N_21855,N_22427);
or U23963 (N_23963,N_21680,N_22360);
and U23964 (N_23964,N_21817,N_21744);
nor U23965 (N_23965,N_22298,N_21925);
or U23966 (N_23966,N_22260,N_22336);
xnor U23967 (N_23967,N_22113,N_22191);
and U23968 (N_23968,N_22094,N_22386);
nor U23969 (N_23969,N_22587,N_21696);
nor U23970 (N_23970,N_22609,N_21750);
xnor U23971 (N_23971,N_22326,N_22449);
xor U23972 (N_23972,N_22019,N_22467);
or U23973 (N_23973,N_22451,N_22180);
and U23974 (N_23974,N_21642,N_21717);
nor U23975 (N_23975,N_22173,N_21955);
nand U23976 (N_23976,N_21965,N_22660);
nor U23977 (N_23977,N_22099,N_22241);
xor U23978 (N_23978,N_22366,N_22117);
nand U23979 (N_23979,N_22048,N_22294);
nand U23980 (N_23980,N_22302,N_22165);
nand U23981 (N_23981,N_22043,N_21865);
nor U23982 (N_23982,N_22035,N_21867);
or U23983 (N_23983,N_22125,N_22671);
nand U23984 (N_23984,N_22254,N_22617);
nand U23985 (N_23985,N_22749,N_22000);
nand U23986 (N_23986,N_21761,N_22406);
xor U23987 (N_23987,N_22554,N_22253);
xor U23988 (N_23988,N_21883,N_22697);
and U23989 (N_23989,N_22266,N_22251);
nand U23990 (N_23990,N_22699,N_21876);
and U23991 (N_23991,N_22350,N_22106);
and U23992 (N_23992,N_21638,N_21958);
xnor U23993 (N_23993,N_22005,N_22389);
xor U23994 (N_23994,N_22682,N_22737);
nor U23995 (N_23995,N_22137,N_22354);
and U23996 (N_23996,N_22776,N_21823);
xnor U23997 (N_23997,N_22107,N_22691);
or U23998 (N_23998,N_22701,N_21790);
or U23999 (N_23999,N_22224,N_22324);
nor U24000 (N_24000,N_23705,N_23204);
nor U24001 (N_24001,N_23458,N_23602);
xnor U24002 (N_24002,N_23987,N_23018);
nor U24003 (N_24003,N_23314,N_23603);
xnor U24004 (N_24004,N_23468,N_23744);
xnor U24005 (N_24005,N_23818,N_23733);
nand U24006 (N_24006,N_23456,N_23230);
nand U24007 (N_24007,N_23627,N_23763);
nor U24008 (N_24008,N_22983,N_22821);
nor U24009 (N_24009,N_22952,N_23779);
nand U24010 (N_24010,N_23301,N_23296);
nand U24011 (N_24011,N_23369,N_23422);
and U24012 (N_24012,N_23546,N_22845);
nand U24013 (N_24013,N_23170,N_23439);
or U24014 (N_24014,N_23393,N_22830);
and U24015 (N_24015,N_22837,N_23073);
or U24016 (N_24016,N_22930,N_23759);
or U24017 (N_24017,N_23995,N_23955);
nand U24018 (N_24018,N_23832,N_23021);
nand U24019 (N_24019,N_23711,N_23923);
nor U24020 (N_24020,N_23402,N_23063);
nor U24021 (N_24021,N_23707,N_23640);
or U24022 (N_24022,N_22899,N_23616);
nor U24023 (N_24023,N_23996,N_23452);
xor U24024 (N_24024,N_23827,N_23467);
and U24025 (N_24025,N_23713,N_23377);
nor U24026 (N_24026,N_23310,N_22907);
or U24027 (N_24027,N_23993,N_22824);
nand U24028 (N_24028,N_23044,N_23428);
xor U24029 (N_24029,N_22802,N_23852);
or U24030 (N_24030,N_23281,N_23365);
nor U24031 (N_24031,N_22999,N_23188);
or U24032 (N_24032,N_23504,N_22886);
xnor U24033 (N_24033,N_22946,N_23644);
and U24034 (N_24034,N_23838,N_22924);
nand U24035 (N_24035,N_23801,N_23734);
nor U24036 (N_24036,N_22892,N_23283);
nor U24037 (N_24037,N_22973,N_23808);
nor U24038 (N_24038,N_23828,N_23473);
nor U24039 (N_24039,N_23237,N_22902);
and U24040 (N_24040,N_23258,N_23342);
or U24041 (N_24041,N_23182,N_23517);
xor U24042 (N_24042,N_23229,N_23806);
xnor U24043 (N_24043,N_23581,N_22887);
nor U24044 (N_24044,N_23459,N_23540);
nand U24045 (N_24045,N_23986,N_23522);
or U24046 (N_24046,N_23972,N_22928);
and U24047 (N_24047,N_23742,N_23814);
and U24048 (N_24048,N_23450,N_23278);
xnor U24049 (N_24049,N_22863,N_23408);
and U24050 (N_24050,N_23169,N_22848);
and U24051 (N_24051,N_23297,N_23211);
xnor U24052 (N_24052,N_22874,N_23110);
and U24053 (N_24053,N_23645,N_22955);
or U24054 (N_24054,N_22914,N_23495);
nor U24055 (N_24055,N_23017,N_23129);
xor U24056 (N_24056,N_23846,N_22953);
xor U24057 (N_24057,N_23153,N_23174);
or U24058 (N_24058,N_22811,N_23290);
and U24059 (N_24059,N_23072,N_23222);
or U24060 (N_24060,N_23698,N_23884);
nor U24061 (N_24061,N_22982,N_23775);
nand U24062 (N_24062,N_23090,N_23712);
nor U24063 (N_24063,N_22843,N_23925);
and U24064 (N_24064,N_23117,N_23354);
nor U24065 (N_24065,N_23317,N_23082);
and U24066 (N_24066,N_23471,N_23465);
nand U24067 (N_24067,N_23735,N_23445);
nor U24068 (N_24068,N_23954,N_23399);
nand U24069 (N_24069,N_23662,N_22950);
nor U24070 (N_24070,N_23489,N_23798);
nor U24071 (N_24071,N_23554,N_23032);
nor U24072 (N_24072,N_23877,N_23717);
xor U24073 (N_24073,N_22947,N_23280);
and U24074 (N_24074,N_23898,N_23218);
nor U24075 (N_24075,N_23526,N_23124);
xnor U24076 (N_24076,N_23694,N_23145);
or U24077 (N_24077,N_23958,N_23931);
nand U24078 (N_24078,N_23669,N_23558);
nand U24079 (N_24079,N_23765,N_23638);
xor U24080 (N_24080,N_23804,N_22877);
nand U24081 (N_24081,N_23689,N_23532);
nand U24082 (N_24082,N_22851,N_23223);
xnor U24083 (N_24083,N_22968,N_23825);
and U24084 (N_24084,N_23515,N_23924);
nor U24085 (N_24085,N_23490,N_23295);
xnor U24086 (N_24086,N_23180,N_23887);
xor U24087 (N_24087,N_23362,N_23658);
nor U24088 (N_24088,N_23686,N_23027);
or U24089 (N_24089,N_23696,N_22980);
nand U24090 (N_24090,N_23646,N_22822);
nand U24091 (N_24091,N_23156,N_23811);
and U24092 (N_24092,N_23071,N_23816);
or U24093 (N_24093,N_23136,N_23692);
xnor U24094 (N_24094,N_23064,N_23305);
xor U24095 (N_24095,N_23580,N_23331);
xnor U24096 (N_24096,N_23328,N_23879);
nor U24097 (N_24097,N_23922,N_23477);
or U24098 (N_24098,N_23433,N_23654);
and U24099 (N_24099,N_23831,N_23535);
nor U24100 (N_24100,N_23441,N_23181);
nand U24101 (N_24101,N_23960,N_23701);
nand U24102 (N_24102,N_23578,N_23030);
or U24103 (N_24103,N_22849,N_23584);
nor U24104 (N_24104,N_22948,N_23327);
nor U24105 (N_24105,N_23661,N_23994);
or U24106 (N_24106,N_23731,N_22862);
nand U24107 (N_24107,N_23394,N_23529);
nor U24108 (N_24108,N_23805,N_23943);
and U24109 (N_24109,N_23053,N_23411);
nor U24110 (N_24110,N_22970,N_23361);
or U24111 (N_24111,N_22963,N_22926);
xor U24112 (N_24112,N_23697,N_23962);
nand U24113 (N_24113,N_23881,N_23829);
nand U24114 (N_24114,N_23464,N_22856);
nand U24115 (N_24115,N_23285,N_23065);
nor U24116 (N_24116,N_23483,N_23074);
and U24117 (N_24117,N_23083,N_23423);
nand U24118 (N_24118,N_22945,N_23363);
and U24119 (N_24119,N_23446,N_23764);
and U24120 (N_24120,N_23872,N_22997);
nand U24121 (N_24121,N_23319,N_23453);
and U24122 (N_24122,N_23956,N_23245);
xnor U24123 (N_24123,N_23338,N_23513);
or U24124 (N_24124,N_23166,N_23118);
nand U24125 (N_24125,N_23966,N_23984);
or U24126 (N_24126,N_23325,N_23760);
and U24127 (N_24127,N_23860,N_23928);
xnor U24128 (N_24128,N_23810,N_23196);
nand U24129 (N_24129,N_23306,N_22844);
or U24130 (N_24130,N_22814,N_23238);
nor U24131 (N_24131,N_23777,N_22978);
and U24132 (N_24132,N_23867,N_22831);
xor U24133 (N_24133,N_23279,N_23219);
and U24134 (N_24134,N_23186,N_23300);
nand U24135 (N_24135,N_23934,N_23563);
xor U24136 (N_24136,N_23198,N_23102);
nand U24137 (N_24137,N_23845,N_23287);
xnor U24138 (N_24138,N_23719,N_23275);
nor U24139 (N_24139,N_23424,N_22855);
and U24140 (N_24140,N_22905,N_23795);
nor U24141 (N_24141,N_23461,N_23699);
nand U24142 (N_24142,N_23594,N_23988);
nor U24143 (N_24143,N_23747,N_22827);
and U24144 (N_24144,N_23493,N_23103);
nor U24145 (N_24145,N_23585,N_23405);
xnor U24146 (N_24146,N_23990,N_22893);
xor U24147 (N_24147,N_23676,N_22909);
or U24148 (N_24148,N_23026,N_23350);
nor U24149 (N_24149,N_22916,N_23187);
nor U24150 (N_24150,N_23056,N_23417);
and U24151 (N_24151,N_23635,N_23142);
and U24152 (N_24152,N_23757,N_22943);
nor U24153 (N_24153,N_23729,N_23911);
or U24154 (N_24154,N_23335,N_23982);
or U24155 (N_24155,N_23214,N_23551);
xnor U24156 (N_24156,N_23787,N_23380);
nor U24157 (N_24157,N_23938,N_23946);
or U24158 (N_24158,N_23854,N_23703);
xor U24159 (N_24159,N_23973,N_22932);
nand U24160 (N_24160,N_23793,N_23632);
nor U24161 (N_24161,N_23171,N_23309);
nand U24162 (N_24162,N_23313,N_23481);
nor U24163 (N_24163,N_23388,N_23998);
and U24164 (N_24164,N_23137,N_23351);
nor U24165 (N_24165,N_23462,N_23057);
nand U24166 (N_24166,N_23284,N_23571);
nand U24167 (N_24167,N_23674,N_23857);
or U24168 (N_24168,N_23918,N_22941);
or U24169 (N_24169,N_22860,N_23190);
and U24170 (N_24170,N_23203,N_23660);
xor U24171 (N_24171,N_23488,N_23500);
xnor U24172 (N_24172,N_23631,N_23050);
nor U24173 (N_24173,N_23786,N_23649);
xor U24174 (N_24174,N_23950,N_23527);
nor U24175 (N_24175,N_22993,N_23677);
nand U24176 (N_24176,N_23837,N_23963);
or U24177 (N_24177,N_23055,N_23045);
nand U24178 (N_24178,N_23671,N_22803);
or U24179 (N_24179,N_23629,N_23407);
nor U24180 (N_24180,N_23965,N_22897);
xor U24181 (N_24181,N_23304,N_23160);
xnor U24182 (N_24182,N_23609,N_23114);
and U24183 (N_24183,N_22890,N_23792);
and U24184 (N_24184,N_22959,N_23431);
nand U24185 (N_24185,N_23151,N_23067);
nand U24186 (N_24186,N_22921,N_23672);
nand U24187 (N_24187,N_23207,N_23200);
xor U24188 (N_24188,N_23656,N_23652);
nand U24189 (N_24189,N_22871,N_23937);
nor U24190 (N_24190,N_23908,N_22813);
and U24191 (N_24191,N_23648,N_23384);
xnor U24192 (N_24192,N_22835,N_23443);
nand U24193 (N_24193,N_23655,N_23101);
xor U24194 (N_24194,N_23058,N_23345);
xnor U24195 (N_24195,N_23667,N_23511);
nand U24196 (N_24196,N_22918,N_22991);
xnor U24197 (N_24197,N_23555,N_23244);
nand U24198 (N_24198,N_23574,N_22884);
nand U24199 (N_24199,N_22939,N_23567);
nor U24200 (N_24200,N_23463,N_23311);
nor U24201 (N_24201,N_23125,N_23600);
nand U24202 (N_24202,N_23113,N_23066);
xor U24203 (N_24203,N_23028,N_23324);
or U24204 (N_24204,N_23016,N_23980);
xor U24205 (N_24205,N_23721,N_22917);
nor U24206 (N_24206,N_23914,N_23842);
nand U24207 (N_24207,N_23812,N_23364);
nor U24208 (N_24208,N_23005,N_22880);
or U24209 (N_24209,N_23193,N_22998);
nand U24210 (N_24210,N_23498,N_23221);
and U24211 (N_24211,N_23208,N_23289);
xnor U24212 (N_24212,N_22958,N_22865);
and U24213 (N_24213,N_23940,N_22976);
xnor U24214 (N_24214,N_23587,N_22913);
nand U24215 (N_24215,N_23605,N_23374);
and U24216 (N_24216,N_22937,N_23025);
or U24217 (N_24217,N_23748,N_23553);
and U24218 (N_24218,N_23243,N_23081);
xnor U24219 (N_24219,N_22858,N_23143);
nor U24220 (N_24220,N_22833,N_23144);
or U24221 (N_24221,N_23782,N_23562);
and U24222 (N_24222,N_23732,N_23861);
nor U24223 (N_24223,N_23564,N_23897);
xor U24224 (N_24224,N_23547,N_23496);
nand U24225 (N_24225,N_23094,N_23167);
nand U24226 (N_24226,N_23132,N_23583);
and U24227 (N_24227,N_22817,N_23409);
or U24228 (N_24228,N_22872,N_23619);
or U24229 (N_24229,N_22942,N_23385);
nor U24230 (N_24230,N_23647,N_23395);
or U24231 (N_24231,N_23178,N_23308);
nor U24232 (N_24232,N_23680,N_23261);
nand U24233 (N_24233,N_23932,N_23163);
nand U24234 (N_24234,N_23282,N_23704);
nand U24235 (N_24235,N_23119,N_23541);
and U24236 (N_24236,N_23612,N_23606);
or U24237 (N_24237,N_23944,N_23097);
nor U24238 (N_24238,N_23069,N_23514);
xor U24239 (N_24239,N_22915,N_22935);
nor U24240 (N_24240,N_23109,N_22852);
nand U24241 (N_24241,N_23576,N_23383);
and U24242 (N_24242,N_23010,N_23949);
nand U24243 (N_24243,N_22891,N_22806);
or U24244 (N_24244,N_23639,N_22800);
or U24245 (N_24245,N_23874,N_23217);
nand U24246 (N_24246,N_23176,N_23199);
xor U24247 (N_24247,N_22894,N_23358);
or U24248 (N_24248,N_23368,N_23068);
nor U24249 (N_24249,N_23903,N_22846);
xnor U24250 (N_24250,N_23893,N_22966);
or U24251 (N_24251,N_23840,N_23778);
nand U24252 (N_24252,N_23856,N_23220);
xor U24253 (N_24253,N_23249,N_23826);
and U24254 (N_24254,N_23184,N_23608);
xnor U24255 (N_24255,N_23620,N_23771);
nor U24256 (N_24256,N_23915,N_23194);
nand U24257 (N_24257,N_22819,N_23716);
and U24258 (N_24258,N_22961,N_23386);
nor U24259 (N_24259,N_23336,N_23008);
or U24260 (N_24260,N_22826,N_23939);
and U24261 (N_24261,N_22944,N_22988);
and U24262 (N_24262,N_23839,N_23271);
and U24263 (N_24263,N_23549,N_23185);
or U24264 (N_24264,N_23286,N_23141);
xor U24265 (N_24265,N_23892,N_23589);
and U24266 (N_24266,N_23543,N_23077);
nand U24267 (N_24267,N_23265,N_23273);
and U24268 (N_24268,N_23231,N_23034);
nand U24269 (N_24269,N_23098,N_23862);
xnor U24270 (N_24270,N_23228,N_23321);
and U24271 (N_24271,N_22840,N_23851);
xor U24272 (N_24272,N_22870,N_23693);
and U24273 (N_24273,N_22828,N_23343);
nor U24274 (N_24274,N_23569,N_23930);
nor U24275 (N_24275,N_23623,N_23312);
or U24276 (N_24276,N_23435,N_23436);
nand U24277 (N_24277,N_23430,N_23189);
nand U24278 (N_24278,N_23382,N_23079);
and U24279 (N_24279,N_23334,N_23687);
and U24280 (N_24280,N_23138,N_22873);
xor U24281 (N_24281,N_23389,N_23085);
or U24282 (N_24282,N_23613,N_23991);
or U24283 (N_24283,N_23533,N_23323);
nor U24284 (N_24284,N_23344,N_22805);
nand U24285 (N_24285,N_23148,N_23545);
and U24286 (N_24286,N_22964,N_23896);
nand U24287 (N_24287,N_23033,N_23899);
nand U24288 (N_24288,N_23418,N_22834);
nand U24289 (N_24289,N_23889,N_23019);
and U24290 (N_24290,N_23873,N_23849);
or U24291 (N_24291,N_23126,N_23227);
or U24292 (N_24292,N_23476,N_22904);
nand U24293 (N_24293,N_23177,N_23294);
and U24294 (N_24294,N_23597,N_23084);
and U24295 (N_24295,N_23339,N_23905);
xnor U24296 (N_24296,N_23349,N_23078);
xor U24297 (N_24297,N_23414,N_23506);
and U24298 (N_24298,N_22812,N_23260);
and U24299 (N_24299,N_23761,N_23725);
and U24300 (N_24300,N_23738,N_23981);
and U24301 (N_24301,N_22934,N_23685);
nor U24302 (N_24302,N_22923,N_23060);
and U24303 (N_24303,N_23355,N_23791);
nor U24304 (N_24304,N_23983,N_22816);
xor U24305 (N_24305,N_23678,N_22954);
nor U24306 (N_24306,N_23853,N_22967);
nand U24307 (N_24307,N_22857,N_23502);
and U24308 (N_24308,N_23337,N_22908);
or U24309 (N_24309,N_23728,N_23212);
and U24310 (N_24310,N_23121,N_23768);
xnor U24311 (N_24311,N_23438,N_23357);
xnor U24312 (N_24312,N_23878,N_23610);
or U24313 (N_24313,N_23108,N_23075);
nor U24314 (N_24314,N_23233,N_23528);
nor U24315 (N_24315,N_23819,N_22854);
xnor U24316 (N_24316,N_23061,N_23259);
and U24317 (N_24317,N_23750,N_23318);
or U24318 (N_24318,N_23226,N_23150);
and U24319 (N_24319,N_23538,N_23758);
xor U24320 (N_24320,N_23642,N_22879);
xor U24321 (N_24321,N_23668,N_23501);
nand U24322 (N_24322,N_23216,N_23088);
nand U24323 (N_24323,N_23876,N_23641);
or U24324 (N_24324,N_23967,N_23413);
and U24325 (N_24325,N_23745,N_23131);
nor U24326 (N_24326,N_23935,N_22920);
and U24327 (N_24327,N_23420,N_23333);
and U24328 (N_24328,N_23266,N_23246);
or U24329 (N_24329,N_23087,N_23859);
or U24330 (N_24330,N_23048,N_23929);
or U24331 (N_24331,N_23598,N_22969);
xor U24332 (N_24332,N_23906,N_23379);
nand U24333 (N_24333,N_23499,N_23800);
and U24334 (N_24334,N_22867,N_23781);
nand U24335 (N_24335,N_22804,N_23622);
xor U24336 (N_24336,N_22979,N_22927);
or U24337 (N_24337,N_23128,N_23002);
nand U24338 (N_24338,N_23096,N_23519);
and U24339 (N_24339,N_23051,N_23679);
nand U24340 (N_24340,N_23272,N_23040);
nor U24341 (N_24341,N_23969,N_22842);
nand U24342 (N_24342,N_23004,N_23945);
or U24343 (N_24343,N_23920,N_22975);
nand U24344 (N_24344,N_23902,N_23895);
nand U24345 (N_24345,N_23469,N_23375);
and U24346 (N_24346,N_22885,N_23059);
nand U24347 (N_24347,N_23270,N_23695);
and U24348 (N_24348,N_23794,N_23883);
xor U24349 (N_24349,N_23039,N_23139);
nor U24350 (N_24350,N_23173,N_23210);
xor U24351 (N_24351,N_23159,N_23807);
nand U24352 (N_24352,N_23157,N_23123);
nor U24353 (N_24353,N_23036,N_23790);
nand U24354 (N_24354,N_23291,N_23521);
nand U24355 (N_24355,N_23263,N_23885);
nand U24356 (N_24356,N_23834,N_22807);
or U24357 (N_24357,N_23657,N_23257);
and U24358 (N_24358,N_23046,N_23251);
nand U24359 (N_24359,N_23421,N_23947);
nor U24360 (N_24360,N_23403,N_23340);
xnor U24361 (N_24361,N_23298,N_23835);
or U24362 (N_24362,N_23534,N_23715);
xnor U24363 (N_24363,N_23844,N_23823);
nor U24364 (N_24364,N_23348,N_23548);
xor U24365 (N_24365,N_23014,N_23556);
or U24366 (N_24366,N_23637,N_23977);
nand U24367 (N_24367,N_23618,N_23236);
nand U24368 (N_24368,N_23232,N_23953);
or U24369 (N_24369,N_23788,N_22815);
nor U24370 (N_24370,N_22996,N_23936);
xor U24371 (N_24371,N_23891,N_23041);
nor U24372 (N_24372,N_23454,N_23643);
nor U24373 (N_24373,N_23213,N_23442);
nor U24374 (N_24374,N_22818,N_22977);
and U24375 (N_24375,N_23723,N_22985);
xor U24376 (N_24376,N_23706,N_22931);
nor U24377 (N_24377,N_23215,N_23447);
and U24378 (N_24378,N_23557,N_22888);
or U24379 (N_24379,N_23663,N_23913);
nand U24380 (N_24380,N_23460,N_23970);
nor U24381 (N_24381,N_23809,N_22995);
nand U24382 (N_24382,N_23080,N_23948);
xnor U24383 (N_24383,N_22981,N_23444);
or U24384 (N_24384,N_23172,N_23783);
xor U24385 (N_24385,N_22882,N_23855);
nor U24386 (N_24386,N_23485,N_23042);
xnor U24387 (N_24387,N_23882,N_23326);
xor U24388 (N_24388,N_23372,N_23880);
nand U24389 (N_24389,N_23951,N_23330);
xnor U24390 (N_24390,N_23665,N_23673);
and U24391 (N_24391,N_23821,N_22951);
xor U24392 (N_24392,N_23523,N_23225);
and U24393 (N_24393,N_23921,N_23907);
nor U24394 (N_24394,N_22919,N_23037);
xor U24395 (N_24395,N_23843,N_23487);
and U24396 (N_24396,N_23242,N_23047);
or U24397 (N_24397,N_23796,N_23653);
nor U24398 (N_24398,N_23542,N_23617);
xor U24399 (N_24399,N_23933,N_22895);
nor U24400 (N_24400,N_23552,N_23659);
nand U24401 (N_24401,N_23866,N_23941);
xnor U24402 (N_24402,N_23961,N_23205);
xnor U24403 (N_24403,N_22901,N_23293);
xnor U24404 (N_24404,N_23890,N_23105);
xnor U24405 (N_24405,N_23234,N_23772);
nand U24406 (N_24406,N_23352,N_23700);
xor U24407 (N_24407,N_23347,N_22925);
xor U24408 (N_24408,N_23155,N_23978);
nand U24409 (N_24409,N_23730,N_23909);
or U24410 (N_24410,N_23106,N_23122);
nand U24411 (N_24411,N_23727,N_23510);
nand U24412 (N_24412,N_23024,N_23315);
or U24413 (N_24413,N_23833,N_23165);
or U24414 (N_24414,N_23590,N_23474);
and U24415 (N_24415,N_22864,N_23651);
and U24416 (N_24416,N_23015,N_23575);
nand U24417 (N_24417,N_23964,N_23754);
nor U24418 (N_24418,N_23415,N_23095);
nor U24419 (N_24419,N_23815,N_23292);
or U24420 (N_24420,N_23746,N_23100);
or U24421 (N_24421,N_23753,N_22829);
or U24422 (N_24422,N_23307,N_23989);
nor U24423 (N_24423,N_23724,N_23817);
xor U24424 (N_24424,N_23478,N_22898);
xor U24425 (N_24425,N_23371,N_23332);
nor U24426 (N_24426,N_23470,N_23070);
nor U24427 (N_24427,N_23250,N_23007);
xnor U24428 (N_24428,N_23472,N_23111);
or U24429 (N_24429,N_23592,N_23869);
xnor U24430 (N_24430,N_23572,N_23550);
or U24431 (N_24431,N_23202,N_23029);
nand U24432 (N_24432,N_22990,N_23086);
xor U24433 (N_24433,N_22820,N_23870);
nor U24434 (N_24434,N_23848,N_23091);
xnor U24435 (N_24435,N_23482,N_23797);
and U24436 (N_24436,N_23404,N_23518);
nor U24437 (N_24437,N_23952,N_23049);
xor U24438 (N_24438,N_22861,N_23038);
and U24439 (N_24439,N_23267,N_23524);
nor U24440 (N_24440,N_23288,N_23168);
xnor U24441 (N_24441,N_23426,N_23916);
nand U24442 (N_24442,N_23636,N_23112);
nor U24443 (N_24443,N_23256,N_22957);
xnor U24444 (N_24444,N_23979,N_23591);
and U24445 (N_24445,N_23255,N_23670);
nor U24446 (N_24446,N_22896,N_22878);
nor U24447 (N_24447,N_23582,N_23247);
nor U24448 (N_24448,N_23802,N_23912);
nand U24449 (N_24449,N_23752,N_22847);
xnor U24450 (N_24450,N_23366,N_22838);
xor U24451 (N_24451,N_23427,N_23161);
xnor U24452 (N_24452,N_23868,N_23135);
xor U24453 (N_24453,N_23376,N_23691);
nand U24454 (N_24454,N_23628,N_23209);
or U24455 (N_24455,N_23799,N_23455);
nor U24456 (N_24456,N_23820,N_23756);
and U24457 (N_24457,N_23926,N_23957);
or U24458 (N_24458,N_23006,N_23560);
xnor U24459 (N_24459,N_23179,N_23822);
and U24460 (N_24460,N_23864,N_23917);
or U24461 (N_24461,N_23531,N_22832);
nor U24462 (N_24462,N_23191,N_22989);
and U24463 (N_24463,N_23904,N_23381);
nor U24464 (N_24464,N_23149,N_23491);
or U24465 (N_24465,N_23052,N_22810);
nand U24466 (N_24466,N_23992,N_23865);
nand U24467 (N_24467,N_22836,N_23942);
xnor U24468 (N_24468,N_23373,N_23419);
nor U24469 (N_24469,N_23633,N_23277);
nor U24470 (N_24470,N_23601,N_23577);
xor U24471 (N_24471,N_23240,N_23755);
or U24472 (N_24472,N_22906,N_23116);
nor U24473 (N_24473,N_23378,N_23975);
nor U24474 (N_24474,N_23900,N_22933);
or U24475 (N_24475,N_23276,N_23824);
nand U24476 (N_24476,N_22987,N_23830);
nand U24477 (N_24477,N_23099,N_23736);
xnor U24478 (N_24478,N_23115,N_23076);
nand U24479 (N_24479,N_23684,N_23726);
xnor U24480 (N_24480,N_23614,N_23570);
and U24481 (N_24481,N_23396,N_22903);
nand U24482 (N_24482,N_23440,N_23505);
nor U24483 (N_24483,N_23743,N_23432);
nand U24484 (N_24484,N_23525,N_23625);
nand U24485 (N_24485,N_22809,N_23023);
nand U24486 (N_24486,N_23847,N_23011);
nor U24487 (N_24487,N_23359,N_22910);
nor U24488 (N_24488,N_23062,N_23536);
nor U24489 (N_24489,N_23492,N_23302);
or U24490 (N_24490,N_23607,N_23107);
xnor U24491 (N_24491,N_23985,N_23720);
and U24492 (N_24492,N_22965,N_23497);
and U24493 (N_24493,N_23565,N_23484);
nor U24494 (N_24494,N_22929,N_23886);
or U24495 (N_24495,N_23356,N_23813);
nor U24496 (N_24496,N_23367,N_22883);
or U24497 (N_24497,N_23681,N_23391);
and U24498 (N_24498,N_23741,N_22922);
or U24499 (N_24499,N_23675,N_23773);
nor U24500 (N_24500,N_23416,N_23089);
xnor U24501 (N_24501,N_23959,N_22825);
nor U24502 (N_24502,N_23709,N_23624);
and U24503 (N_24503,N_23568,N_23769);
and U24504 (N_24504,N_23593,N_23449);
nand U24505 (N_24505,N_23054,N_23009);
and U24506 (N_24506,N_23714,N_22912);
or U24507 (N_24507,N_23316,N_23586);
xor U24508 (N_24508,N_23248,N_22839);
and U24509 (N_24509,N_23013,N_23360);
and U24510 (N_24510,N_23274,N_23000);
nand U24511 (N_24511,N_22992,N_23392);
or U24512 (N_24512,N_23434,N_23762);
nor U24513 (N_24513,N_23252,N_22962);
or U24514 (N_24514,N_23195,N_23774);
or U24515 (N_24515,N_22801,N_22960);
nand U24516 (N_24516,N_23634,N_23020);
xnor U24517 (N_24517,N_22972,N_23400);
and U24518 (N_24518,N_23708,N_23262);
xor U24519 (N_24519,N_23516,N_23269);
xnor U24520 (N_24520,N_22911,N_23927);
nor U24521 (N_24521,N_23154,N_23561);
xor U24522 (N_24522,N_23001,N_23626);
or U24523 (N_24523,N_23164,N_23406);
nor U24524 (N_24524,N_23588,N_23457);
and U24525 (N_24525,N_23664,N_23650);
and U24526 (N_24526,N_23871,N_23971);
nor U24527 (N_24527,N_23599,N_22868);
nor U24528 (N_24528,N_23206,N_23264);
or U24529 (N_24529,N_22940,N_23322);
and U24530 (N_24530,N_23451,N_23875);
and U24531 (N_24531,N_23503,N_23999);
xnor U24532 (N_24532,N_23539,N_23390);
and U24533 (N_24533,N_23401,N_23201);
and U24534 (N_24534,N_23688,N_23162);
xnor U24535 (N_24535,N_22938,N_23370);
nor U24536 (N_24536,N_23475,N_23239);
nand U24537 (N_24537,N_23850,N_23303);
and U24538 (N_24538,N_23043,N_23780);
or U24539 (N_24539,N_23329,N_22859);
nor U24540 (N_24540,N_23702,N_23509);
nand U24541 (N_24541,N_23718,N_23093);
nor U24542 (N_24542,N_23486,N_23412);
nand U24543 (N_24543,N_23919,N_23740);
nand U24544 (N_24544,N_23480,N_22876);
or U24545 (N_24545,N_23133,N_23183);
or U24546 (N_24546,N_23320,N_23770);
or U24547 (N_24547,N_23092,N_23863);
nand U24548 (N_24548,N_23630,N_23530);
or U24549 (N_24549,N_23566,N_23968);
nor U24550 (N_24550,N_23573,N_23690);
xnor U24551 (N_24551,N_23710,N_23254);
xor U24552 (N_24552,N_23784,N_23134);
nand U24553 (N_24553,N_23479,N_23437);
nand U24554 (N_24554,N_23299,N_22984);
nor U24555 (N_24555,N_23507,N_23682);
nand U24556 (N_24556,N_23596,N_22974);
nor U24557 (N_24557,N_23398,N_23429);
xnor U24558 (N_24558,N_22869,N_23512);
nand U24559 (N_24559,N_23766,N_23241);
and U24560 (N_24560,N_23767,N_23888);
xnor U24561 (N_24561,N_23666,N_23341);
nand U24562 (N_24562,N_22994,N_23425);
or U24563 (N_24563,N_22875,N_23776);
nand U24564 (N_24564,N_23268,N_23253);
nand U24565 (N_24565,N_23120,N_23031);
nand U24566 (N_24566,N_23158,N_23894);
nor U24567 (N_24567,N_22949,N_23022);
nand U24568 (N_24568,N_23611,N_22936);
or U24569 (N_24569,N_23127,N_23858);
nor U24570 (N_24570,N_23224,N_23494);
xor U24571 (N_24571,N_23130,N_23997);
xnor U24572 (N_24572,N_22850,N_22881);
nand U24573 (N_24573,N_23520,N_23146);
nand U24574 (N_24574,N_23749,N_23235);
nand U24575 (N_24575,N_22889,N_23152);
nand U24576 (N_24576,N_23974,N_23910);
and U24577 (N_24577,N_23621,N_22823);
xnor U24578 (N_24578,N_23785,N_23615);
and U24579 (N_24579,N_23448,N_23537);
nand U24580 (N_24580,N_23737,N_23197);
nand U24581 (N_24581,N_23346,N_22900);
nor U24582 (N_24582,N_23035,N_23466);
xnor U24583 (N_24583,N_23192,N_22866);
or U24584 (N_24584,N_23544,N_22841);
or U24585 (N_24585,N_23579,N_23722);
or U24586 (N_24586,N_23803,N_23387);
nand U24587 (N_24587,N_22956,N_23901);
xnor U24588 (N_24588,N_22808,N_23739);
and U24589 (N_24589,N_22853,N_23595);
xor U24590 (N_24590,N_23353,N_23104);
nor U24591 (N_24591,N_23175,N_23559);
xnor U24592 (N_24592,N_23841,N_23147);
or U24593 (N_24593,N_23397,N_23003);
xnor U24594 (N_24594,N_23976,N_22986);
nand U24595 (N_24595,N_23683,N_23508);
or U24596 (N_24596,N_23836,N_22971);
nor U24597 (N_24597,N_23140,N_23410);
nor U24598 (N_24598,N_23012,N_23789);
or U24599 (N_24599,N_23751,N_23604);
nor U24600 (N_24600,N_22985,N_23667);
nand U24601 (N_24601,N_23687,N_23910);
and U24602 (N_24602,N_23971,N_22943);
xnor U24603 (N_24603,N_23135,N_23904);
nor U24604 (N_24604,N_23670,N_23341);
or U24605 (N_24605,N_23491,N_22837);
nor U24606 (N_24606,N_22883,N_23765);
or U24607 (N_24607,N_23844,N_23334);
xnor U24608 (N_24608,N_22959,N_23156);
xnor U24609 (N_24609,N_22956,N_23641);
or U24610 (N_24610,N_23281,N_23090);
nor U24611 (N_24611,N_22830,N_23184);
and U24612 (N_24612,N_23906,N_23628);
xor U24613 (N_24613,N_23190,N_23687);
nand U24614 (N_24614,N_23073,N_23665);
nand U24615 (N_24615,N_23480,N_23853);
or U24616 (N_24616,N_23978,N_22850);
and U24617 (N_24617,N_23071,N_23534);
nor U24618 (N_24618,N_23739,N_23133);
nor U24619 (N_24619,N_22902,N_23084);
nand U24620 (N_24620,N_23623,N_22810);
and U24621 (N_24621,N_22876,N_23051);
nand U24622 (N_24622,N_23371,N_23991);
nor U24623 (N_24623,N_23084,N_23836);
nand U24624 (N_24624,N_23588,N_22825);
xnor U24625 (N_24625,N_23359,N_23903);
and U24626 (N_24626,N_23882,N_23230);
and U24627 (N_24627,N_23205,N_23868);
xnor U24628 (N_24628,N_23789,N_23693);
nand U24629 (N_24629,N_23380,N_23539);
nand U24630 (N_24630,N_23964,N_23231);
nor U24631 (N_24631,N_23524,N_23739);
and U24632 (N_24632,N_23845,N_23166);
nand U24633 (N_24633,N_23197,N_23909);
and U24634 (N_24634,N_23347,N_23046);
nor U24635 (N_24635,N_23204,N_23429);
and U24636 (N_24636,N_23422,N_23907);
nor U24637 (N_24637,N_23761,N_23570);
or U24638 (N_24638,N_22994,N_22822);
xor U24639 (N_24639,N_22975,N_22957);
nor U24640 (N_24640,N_23188,N_23889);
nand U24641 (N_24641,N_23656,N_23048);
or U24642 (N_24642,N_23808,N_22908);
xor U24643 (N_24643,N_23213,N_22811);
nand U24644 (N_24644,N_23002,N_23497);
nor U24645 (N_24645,N_23848,N_23250);
xnor U24646 (N_24646,N_23917,N_23158);
nor U24647 (N_24647,N_23446,N_23674);
xnor U24648 (N_24648,N_22856,N_23898);
and U24649 (N_24649,N_23242,N_23157);
xnor U24650 (N_24650,N_23882,N_23851);
xnor U24651 (N_24651,N_23148,N_23410);
nor U24652 (N_24652,N_23499,N_22836);
nand U24653 (N_24653,N_23594,N_22857);
nor U24654 (N_24654,N_23589,N_23600);
nor U24655 (N_24655,N_23176,N_23238);
or U24656 (N_24656,N_23602,N_23118);
nand U24657 (N_24657,N_23383,N_23134);
nor U24658 (N_24658,N_22883,N_22904);
xnor U24659 (N_24659,N_22993,N_23508);
nand U24660 (N_24660,N_23463,N_22865);
xnor U24661 (N_24661,N_23846,N_23273);
nand U24662 (N_24662,N_22985,N_23021);
xor U24663 (N_24663,N_22861,N_22852);
xor U24664 (N_24664,N_23745,N_23438);
and U24665 (N_24665,N_22833,N_23874);
xor U24666 (N_24666,N_23962,N_23432);
nor U24667 (N_24667,N_23153,N_22838);
or U24668 (N_24668,N_23222,N_23644);
or U24669 (N_24669,N_23872,N_23887);
nand U24670 (N_24670,N_23382,N_23135);
or U24671 (N_24671,N_23271,N_23927);
and U24672 (N_24672,N_23561,N_23317);
or U24673 (N_24673,N_23458,N_23791);
and U24674 (N_24674,N_23078,N_23021);
and U24675 (N_24675,N_23051,N_23345);
xor U24676 (N_24676,N_22839,N_23357);
and U24677 (N_24677,N_23017,N_23466);
nand U24678 (N_24678,N_22930,N_23636);
nor U24679 (N_24679,N_23368,N_22893);
xor U24680 (N_24680,N_23660,N_23609);
xnor U24681 (N_24681,N_23653,N_23264);
and U24682 (N_24682,N_23636,N_23863);
xnor U24683 (N_24683,N_22812,N_23277);
nor U24684 (N_24684,N_22888,N_23235);
nand U24685 (N_24685,N_22889,N_22967);
and U24686 (N_24686,N_22878,N_22836);
xnor U24687 (N_24687,N_23052,N_23449);
or U24688 (N_24688,N_23826,N_23378);
nand U24689 (N_24689,N_22894,N_23404);
or U24690 (N_24690,N_23883,N_23389);
and U24691 (N_24691,N_22971,N_23792);
nand U24692 (N_24692,N_23366,N_23469);
nand U24693 (N_24693,N_23948,N_23713);
nor U24694 (N_24694,N_23612,N_23927);
or U24695 (N_24695,N_23354,N_22810);
and U24696 (N_24696,N_22802,N_23101);
nor U24697 (N_24697,N_23926,N_23053);
xnor U24698 (N_24698,N_23764,N_22804);
or U24699 (N_24699,N_22822,N_22853);
nor U24700 (N_24700,N_22855,N_22911);
xor U24701 (N_24701,N_23629,N_23641);
nor U24702 (N_24702,N_23861,N_22969);
nand U24703 (N_24703,N_23937,N_23746);
nand U24704 (N_24704,N_23771,N_23243);
xor U24705 (N_24705,N_23245,N_22855);
xnor U24706 (N_24706,N_22837,N_22937);
xor U24707 (N_24707,N_22899,N_23993);
nor U24708 (N_24708,N_22868,N_23193);
nor U24709 (N_24709,N_22948,N_23654);
xnor U24710 (N_24710,N_23829,N_22862);
nand U24711 (N_24711,N_23642,N_23145);
xnor U24712 (N_24712,N_23121,N_23673);
or U24713 (N_24713,N_23663,N_23334);
nor U24714 (N_24714,N_23786,N_22910);
or U24715 (N_24715,N_23472,N_23029);
nand U24716 (N_24716,N_23512,N_23164);
xnor U24717 (N_24717,N_23221,N_23270);
or U24718 (N_24718,N_23035,N_23515);
nand U24719 (N_24719,N_23025,N_23280);
nor U24720 (N_24720,N_23455,N_23276);
nand U24721 (N_24721,N_23499,N_23793);
xnor U24722 (N_24722,N_23127,N_23808);
and U24723 (N_24723,N_23389,N_23277);
and U24724 (N_24724,N_23518,N_23409);
and U24725 (N_24725,N_23845,N_23699);
and U24726 (N_24726,N_23119,N_22852);
nor U24727 (N_24727,N_23209,N_23013);
and U24728 (N_24728,N_23808,N_22852);
nor U24729 (N_24729,N_23896,N_23243);
or U24730 (N_24730,N_23897,N_23607);
xor U24731 (N_24731,N_23001,N_23419);
or U24732 (N_24732,N_23944,N_23926);
xnor U24733 (N_24733,N_23505,N_23986);
and U24734 (N_24734,N_23315,N_23668);
nand U24735 (N_24735,N_23696,N_23413);
and U24736 (N_24736,N_23617,N_23183);
or U24737 (N_24737,N_23016,N_23541);
and U24738 (N_24738,N_23344,N_23776);
xor U24739 (N_24739,N_23086,N_23781);
xor U24740 (N_24740,N_23405,N_23100);
or U24741 (N_24741,N_23382,N_23387);
nand U24742 (N_24742,N_22812,N_23679);
nand U24743 (N_24743,N_23512,N_23051);
and U24744 (N_24744,N_23017,N_23528);
nor U24745 (N_24745,N_23183,N_23240);
or U24746 (N_24746,N_23163,N_23002);
nor U24747 (N_24747,N_22864,N_23599);
xor U24748 (N_24748,N_23522,N_23240);
and U24749 (N_24749,N_23271,N_22927);
nand U24750 (N_24750,N_23842,N_23396);
and U24751 (N_24751,N_23295,N_22837);
nor U24752 (N_24752,N_23948,N_23975);
xnor U24753 (N_24753,N_23626,N_23983);
and U24754 (N_24754,N_23933,N_23770);
nor U24755 (N_24755,N_23654,N_23283);
and U24756 (N_24756,N_23643,N_23146);
or U24757 (N_24757,N_22990,N_23267);
xnor U24758 (N_24758,N_23221,N_23358);
xor U24759 (N_24759,N_23823,N_23165);
nand U24760 (N_24760,N_23724,N_22884);
xor U24761 (N_24761,N_23619,N_22839);
and U24762 (N_24762,N_23848,N_23601);
xnor U24763 (N_24763,N_23828,N_23939);
nor U24764 (N_24764,N_23227,N_22875);
xnor U24765 (N_24765,N_23512,N_23845);
and U24766 (N_24766,N_22889,N_23512);
xnor U24767 (N_24767,N_23065,N_23195);
xnor U24768 (N_24768,N_23150,N_22925);
xor U24769 (N_24769,N_23923,N_23798);
and U24770 (N_24770,N_22840,N_23082);
xnor U24771 (N_24771,N_23430,N_23617);
nor U24772 (N_24772,N_23936,N_23723);
xor U24773 (N_24773,N_23137,N_23533);
nand U24774 (N_24774,N_22868,N_23508);
or U24775 (N_24775,N_22945,N_23959);
nor U24776 (N_24776,N_23775,N_23748);
nor U24777 (N_24777,N_23276,N_23352);
nor U24778 (N_24778,N_23974,N_23525);
or U24779 (N_24779,N_23341,N_23224);
nand U24780 (N_24780,N_23364,N_23176);
or U24781 (N_24781,N_23075,N_23450);
xnor U24782 (N_24782,N_22907,N_23114);
nor U24783 (N_24783,N_23931,N_22965);
or U24784 (N_24784,N_23239,N_23015);
nand U24785 (N_24785,N_23728,N_23895);
and U24786 (N_24786,N_23208,N_23918);
and U24787 (N_24787,N_23235,N_23841);
nor U24788 (N_24788,N_23300,N_23704);
or U24789 (N_24789,N_23992,N_23496);
nand U24790 (N_24790,N_22971,N_23076);
or U24791 (N_24791,N_23715,N_23834);
or U24792 (N_24792,N_23029,N_23215);
nor U24793 (N_24793,N_23555,N_22859);
nand U24794 (N_24794,N_23468,N_23387);
nor U24795 (N_24795,N_23302,N_23670);
nand U24796 (N_24796,N_23037,N_23248);
nand U24797 (N_24797,N_23172,N_23036);
nor U24798 (N_24798,N_23806,N_23191);
nor U24799 (N_24799,N_23578,N_23637);
xor U24800 (N_24800,N_23198,N_22986);
nand U24801 (N_24801,N_23487,N_22955);
and U24802 (N_24802,N_23682,N_23900);
xor U24803 (N_24803,N_23425,N_23147);
or U24804 (N_24804,N_23835,N_23852);
or U24805 (N_24805,N_23135,N_23016);
xnor U24806 (N_24806,N_23995,N_23871);
or U24807 (N_24807,N_23127,N_23162);
nand U24808 (N_24808,N_23723,N_23842);
or U24809 (N_24809,N_23386,N_23034);
and U24810 (N_24810,N_23515,N_23966);
nor U24811 (N_24811,N_23178,N_23486);
or U24812 (N_24812,N_23378,N_23208);
xor U24813 (N_24813,N_23933,N_23052);
xor U24814 (N_24814,N_23146,N_23839);
and U24815 (N_24815,N_23324,N_23531);
and U24816 (N_24816,N_23698,N_23245);
or U24817 (N_24817,N_23892,N_23926);
or U24818 (N_24818,N_23803,N_23094);
nand U24819 (N_24819,N_23710,N_23120);
or U24820 (N_24820,N_23138,N_23636);
nand U24821 (N_24821,N_23502,N_23373);
xnor U24822 (N_24822,N_23787,N_23383);
nor U24823 (N_24823,N_22873,N_23943);
xor U24824 (N_24824,N_23080,N_22964);
and U24825 (N_24825,N_23089,N_23093);
and U24826 (N_24826,N_23920,N_23510);
or U24827 (N_24827,N_23392,N_23618);
xor U24828 (N_24828,N_22860,N_22930);
xor U24829 (N_24829,N_22945,N_23705);
nor U24830 (N_24830,N_23964,N_22917);
nand U24831 (N_24831,N_22907,N_23368);
and U24832 (N_24832,N_23196,N_23670);
nor U24833 (N_24833,N_22886,N_23652);
xor U24834 (N_24834,N_23225,N_22908);
xor U24835 (N_24835,N_22877,N_22934);
and U24836 (N_24836,N_23219,N_23173);
or U24837 (N_24837,N_22834,N_23293);
nand U24838 (N_24838,N_23074,N_23574);
nor U24839 (N_24839,N_23706,N_22954);
xor U24840 (N_24840,N_23866,N_23830);
nor U24841 (N_24841,N_23457,N_23442);
nand U24842 (N_24842,N_22918,N_23315);
or U24843 (N_24843,N_23826,N_23347);
xor U24844 (N_24844,N_22856,N_23404);
nor U24845 (N_24845,N_23425,N_23019);
and U24846 (N_24846,N_23701,N_23005);
xor U24847 (N_24847,N_23509,N_23517);
and U24848 (N_24848,N_23313,N_23370);
or U24849 (N_24849,N_23995,N_23374);
or U24850 (N_24850,N_23674,N_23440);
nor U24851 (N_24851,N_23668,N_23016);
xnor U24852 (N_24852,N_23224,N_23725);
nor U24853 (N_24853,N_22891,N_23311);
or U24854 (N_24854,N_23074,N_23885);
or U24855 (N_24855,N_23077,N_22989);
xor U24856 (N_24856,N_23473,N_23834);
or U24857 (N_24857,N_23318,N_23877);
or U24858 (N_24858,N_23295,N_23127);
or U24859 (N_24859,N_23028,N_23944);
nor U24860 (N_24860,N_23908,N_23034);
xnor U24861 (N_24861,N_23927,N_23677);
and U24862 (N_24862,N_22931,N_23318);
nor U24863 (N_24863,N_22818,N_23234);
and U24864 (N_24864,N_23778,N_23400);
nand U24865 (N_24865,N_22950,N_23578);
xnor U24866 (N_24866,N_23263,N_22936);
or U24867 (N_24867,N_23830,N_23325);
and U24868 (N_24868,N_23507,N_23367);
or U24869 (N_24869,N_23390,N_23407);
nor U24870 (N_24870,N_23064,N_23115);
xnor U24871 (N_24871,N_23162,N_23220);
nor U24872 (N_24872,N_23262,N_23651);
or U24873 (N_24873,N_23914,N_23861);
nor U24874 (N_24874,N_23759,N_23041);
xor U24875 (N_24875,N_23995,N_23496);
or U24876 (N_24876,N_23575,N_23941);
nor U24877 (N_24877,N_23120,N_23334);
xnor U24878 (N_24878,N_23120,N_23141);
and U24879 (N_24879,N_23533,N_23582);
and U24880 (N_24880,N_23291,N_23985);
nand U24881 (N_24881,N_23620,N_23875);
nor U24882 (N_24882,N_23614,N_22869);
nand U24883 (N_24883,N_23365,N_22832);
nor U24884 (N_24884,N_23876,N_22991);
and U24885 (N_24885,N_22852,N_23982);
or U24886 (N_24886,N_23046,N_23560);
or U24887 (N_24887,N_23924,N_22837);
or U24888 (N_24888,N_22860,N_23596);
nand U24889 (N_24889,N_22931,N_23877);
and U24890 (N_24890,N_23776,N_23606);
and U24891 (N_24891,N_23416,N_23302);
xnor U24892 (N_24892,N_23280,N_23474);
and U24893 (N_24893,N_23408,N_23484);
xnor U24894 (N_24894,N_23403,N_23928);
or U24895 (N_24895,N_23403,N_23475);
nor U24896 (N_24896,N_23457,N_23610);
xor U24897 (N_24897,N_22952,N_23683);
nor U24898 (N_24898,N_22844,N_23913);
xor U24899 (N_24899,N_23987,N_23677);
nor U24900 (N_24900,N_23729,N_23779);
or U24901 (N_24901,N_23539,N_22927);
nand U24902 (N_24902,N_23424,N_23059);
xor U24903 (N_24903,N_23625,N_23450);
nand U24904 (N_24904,N_23235,N_23048);
and U24905 (N_24905,N_23929,N_23616);
or U24906 (N_24906,N_23682,N_23266);
nand U24907 (N_24907,N_23095,N_23597);
nor U24908 (N_24908,N_22926,N_23855);
or U24909 (N_24909,N_22937,N_23100);
or U24910 (N_24910,N_23119,N_23219);
xor U24911 (N_24911,N_23239,N_23303);
and U24912 (N_24912,N_22814,N_23201);
nand U24913 (N_24913,N_23252,N_23020);
or U24914 (N_24914,N_23732,N_23089);
nand U24915 (N_24915,N_23677,N_23680);
xnor U24916 (N_24916,N_23286,N_23630);
nor U24917 (N_24917,N_22853,N_23777);
and U24918 (N_24918,N_23402,N_23962);
and U24919 (N_24919,N_22998,N_23168);
or U24920 (N_24920,N_22968,N_23077);
nor U24921 (N_24921,N_23714,N_23175);
and U24922 (N_24922,N_23142,N_23763);
or U24923 (N_24923,N_23072,N_23681);
nor U24924 (N_24924,N_23433,N_23234);
and U24925 (N_24925,N_23030,N_23366);
nor U24926 (N_24926,N_23350,N_23270);
or U24927 (N_24927,N_23952,N_23419);
nand U24928 (N_24928,N_23007,N_23417);
or U24929 (N_24929,N_23207,N_23597);
or U24930 (N_24930,N_23091,N_23748);
and U24931 (N_24931,N_23805,N_23657);
nor U24932 (N_24932,N_23313,N_22903);
nand U24933 (N_24933,N_23669,N_22985);
nand U24934 (N_24934,N_23737,N_23678);
nand U24935 (N_24935,N_23209,N_23306);
and U24936 (N_24936,N_23074,N_22994);
xnor U24937 (N_24937,N_23510,N_23852);
xnor U24938 (N_24938,N_23849,N_22817);
nor U24939 (N_24939,N_23117,N_23280);
nor U24940 (N_24940,N_23114,N_23010);
nor U24941 (N_24941,N_23386,N_23689);
nor U24942 (N_24942,N_23881,N_23105);
xor U24943 (N_24943,N_23235,N_23408);
and U24944 (N_24944,N_23625,N_23172);
and U24945 (N_24945,N_22882,N_23267);
or U24946 (N_24946,N_23843,N_23184);
nand U24947 (N_24947,N_23915,N_23981);
nand U24948 (N_24948,N_22915,N_23349);
or U24949 (N_24949,N_22849,N_23855);
xor U24950 (N_24950,N_23545,N_23368);
nor U24951 (N_24951,N_23932,N_23997);
or U24952 (N_24952,N_23932,N_23120);
nor U24953 (N_24953,N_22859,N_23982);
and U24954 (N_24954,N_23605,N_23273);
and U24955 (N_24955,N_23565,N_22869);
or U24956 (N_24956,N_23684,N_23629);
xnor U24957 (N_24957,N_23763,N_23519);
nor U24958 (N_24958,N_22947,N_22834);
or U24959 (N_24959,N_23519,N_23281);
and U24960 (N_24960,N_23126,N_23050);
nor U24961 (N_24961,N_22893,N_23605);
nor U24962 (N_24962,N_23137,N_23968);
or U24963 (N_24963,N_23432,N_23745);
and U24964 (N_24964,N_23369,N_23941);
or U24965 (N_24965,N_23567,N_23566);
nor U24966 (N_24966,N_23953,N_23794);
and U24967 (N_24967,N_23400,N_23100);
or U24968 (N_24968,N_23552,N_23112);
and U24969 (N_24969,N_23886,N_23631);
nor U24970 (N_24970,N_23676,N_23680);
xor U24971 (N_24971,N_23416,N_23534);
and U24972 (N_24972,N_23856,N_23625);
or U24973 (N_24973,N_23070,N_23293);
or U24974 (N_24974,N_22823,N_23346);
and U24975 (N_24975,N_23326,N_23075);
nand U24976 (N_24976,N_23544,N_23384);
xor U24977 (N_24977,N_23481,N_23161);
nor U24978 (N_24978,N_23224,N_23353);
and U24979 (N_24979,N_23066,N_23552);
nand U24980 (N_24980,N_23353,N_23864);
and U24981 (N_24981,N_23961,N_23041);
nand U24982 (N_24982,N_22903,N_23770);
nand U24983 (N_24983,N_23455,N_23701);
and U24984 (N_24984,N_23784,N_23377);
nor U24985 (N_24985,N_23964,N_23753);
nor U24986 (N_24986,N_23666,N_23304);
and U24987 (N_24987,N_23804,N_23654);
and U24988 (N_24988,N_23014,N_22954);
xor U24989 (N_24989,N_23923,N_23797);
nand U24990 (N_24990,N_23819,N_23524);
and U24991 (N_24991,N_23563,N_22815);
and U24992 (N_24992,N_23446,N_23573);
xor U24993 (N_24993,N_23373,N_23687);
nand U24994 (N_24994,N_23183,N_22861);
nand U24995 (N_24995,N_23705,N_23263);
nand U24996 (N_24996,N_23915,N_23623);
and U24997 (N_24997,N_22860,N_23931);
nor U24998 (N_24998,N_23793,N_23238);
and U24999 (N_24999,N_23823,N_23499);
xnor U25000 (N_25000,N_22893,N_23183);
and U25001 (N_25001,N_23189,N_23617);
nand U25002 (N_25002,N_23613,N_22854);
and U25003 (N_25003,N_23885,N_23862);
nand U25004 (N_25004,N_23019,N_23913);
nand U25005 (N_25005,N_23021,N_22806);
xnor U25006 (N_25006,N_23348,N_22843);
and U25007 (N_25007,N_23372,N_22904);
nand U25008 (N_25008,N_23122,N_23920);
xor U25009 (N_25009,N_22801,N_23558);
nor U25010 (N_25010,N_23783,N_22829);
or U25011 (N_25011,N_22950,N_23722);
and U25012 (N_25012,N_22990,N_23300);
nor U25013 (N_25013,N_23588,N_23544);
xor U25014 (N_25014,N_23391,N_23400);
xor U25015 (N_25015,N_23447,N_23078);
or U25016 (N_25016,N_23040,N_23981);
nand U25017 (N_25017,N_23270,N_23680);
or U25018 (N_25018,N_23244,N_23791);
or U25019 (N_25019,N_22952,N_23119);
or U25020 (N_25020,N_23535,N_23077);
nor U25021 (N_25021,N_22923,N_23640);
nor U25022 (N_25022,N_23149,N_23076);
nor U25023 (N_25023,N_23959,N_23660);
nor U25024 (N_25024,N_22831,N_23937);
or U25025 (N_25025,N_23112,N_23747);
nor U25026 (N_25026,N_23206,N_23984);
xor U25027 (N_25027,N_23753,N_23764);
and U25028 (N_25028,N_23537,N_23426);
or U25029 (N_25029,N_23332,N_23349);
and U25030 (N_25030,N_23854,N_23908);
nor U25031 (N_25031,N_23506,N_23792);
nand U25032 (N_25032,N_23198,N_22976);
or U25033 (N_25033,N_23872,N_23792);
nor U25034 (N_25034,N_23723,N_23319);
nor U25035 (N_25035,N_23403,N_23985);
nand U25036 (N_25036,N_23933,N_23070);
xor U25037 (N_25037,N_23570,N_23616);
xor U25038 (N_25038,N_23091,N_23423);
nand U25039 (N_25039,N_22893,N_23188);
nand U25040 (N_25040,N_23373,N_23657);
nor U25041 (N_25041,N_23967,N_23281);
xnor U25042 (N_25042,N_22846,N_23151);
xor U25043 (N_25043,N_23277,N_23861);
xor U25044 (N_25044,N_23049,N_23443);
xnor U25045 (N_25045,N_22865,N_23165);
or U25046 (N_25046,N_23574,N_23747);
and U25047 (N_25047,N_22872,N_23502);
nor U25048 (N_25048,N_23246,N_23598);
nand U25049 (N_25049,N_23918,N_22954);
xnor U25050 (N_25050,N_23900,N_23016);
and U25051 (N_25051,N_23866,N_23849);
nand U25052 (N_25052,N_23960,N_23504);
nand U25053 (N_25053,N_23222,N_23865);
or U25054 (N_25054,N_23467,N_23866);
nand U25055 (N_25055,N_23655,N_22925);
nor U25056 (N_25056,N_23134,N_23790);
nand U25057 (N_25057,N_23401,N_23480);
or U25058 (N_25058,N_23980,N_22975);
and U25059 (N_25059,N_23056,N_23164);
and U25060 (N_25060,N_23209,N_23820);
nand U25061 (N_25061,N_23312,N_23267);
nand U25062 (N_25062,N_23774,N_23521);
or U25063 (N_25063,N_22837,N_23481);
and U25064 (N_25064,N_22983,N_22931);
nand U25065 (N_25065,N_23197,N_23421);
and U25066 (N_25066,N_23755,N_23979);
xor U25067 (N_25067,N_23121,N_23853);
nand U25068 (N_25068,N_23648,N_23612);
and U25069 (N_25069,N_22965,N_23512);
or U25070 (N_25070,N_23257,N_23388);
nor U25071 (N_25071,N_23529,N_22937);
or U25072 (N_25072,N_23479,N_23007);
xnor U25073 (N_25073,N_23243,N_23235);
nand U25074 (N_25074,N_23672,N_23512);
or U25075 (N_25075,N_23728,N_23361);
or U25076 (N_25076,N_22931,N_22927);
nand U25077 (N_25077,N_22991,N_23974);
nor U25078 (N_25078,N_23180,N_22808);
or U25079 (N_25079,N_23590,N_23381);
xor U25080 (N_25080,N_23710,N_22869);
or U25081 (N_25081,N_23930,N_23651);
or U25082 (N_25082,N_23095,N_23491);
or U25083 (N_25083,N_23438,N_23530);
and U25084 (N_25084,N_23644,N_23097);
xor U25085 (N_25085,N_23911,N_23566);
or U25086 (N_25086,N_22932,N_23682);
nand U25087 (N_25087,N_23859,N_22895);
nand U25088 (N_25088,N_23909,N_23198);
or U25089 (N_25089,N_23896,N_23692);
xnor U25090 (N_25090,N_23479,N_23898);
and U25091 (N_25091,N_23992,N_23021);
and U25092 (N_25092,N_23598,N_23444);
xor U25093 (N_25093,N_23669,N_23933);
or U25094 (N_25094,N_23691,N_23285);
or U25095 (N_25095,N_23204,N_23979);
or U25096 (N_25096,N_23720,N_23307);
nand U25097 (N_25097,N_23780,N_23560);
xor U25098 (N_25098,N_22819,N_23127);
or U25099 (N_25099,N_23083,N_23955);
or U25100 (N_25100,N_23483,N_23060);
xor U25101 (N_25101,N_23173,N_23398);
nor U25102 (N_25102,N_23254,N_23160);
nor U25103 (N_25103,N_23440,N_23135);
xnor U25104 (N_25104,N_23048,N_23017);
and U25105 (N_25105,N_23798,N_23240);
nor U25106 (N_25106,N_23159,N_23053);
and U25107 (N_25107,N_23221,N_23843);
nor U25108 (N_25108,N_23180,N_23838);
xor U25109 (N_25109,N_23319,N_23974);
nand U25110 (N_25110,N_23714,N_23979);
or U25111 (N_25111,N_23783,N_23470);
or U25112 (N_25112,N_23214,N_22948);
nor U25113 (N_25113,N_23930,N_23881);
nor U25114 (N_25114,N_23933,N_22992);
nand U25115 (N_25115,N_23775,N_23025);
or U25116 (N_25116,N_23777,N_22911);
nand U25117 (N_25117,N_23488,N_23807);
and U25118 (N_25118,N_22901,N_23861);
nand U25119 (N_25119,N_23167,N_23528);
nand U25120 (N_25120,N_23021,N_23172);
nand U25121 (N_25121,N_23261,N_23216);
nand U25122 (N_25122,N_23746,N_22955);
nor U25123 (N_25123,N_23908,N_23281);
nor U25124 (N_25124,N_23095,N_23055);
xnor U25125 (N_25125,N_23675,N_23653);
nand U25126 (N_25126,N_23627,N_23545);
and U25127 (N_25127,N_23109,N_23548);
or U25128 (N_25128,N_23194,N_23044);
nor U25129 (N_25129,N_23910,N_23830);
xnor U25130 (N_25130,N_23100,N_22826);
nor U25131 (N_25131,N_23828,N_23845);
nor U25132 (N_25132,N_23917,N_23626);
nand U25133 (N_25133,N_23638,N_23850);
and U25134 (N_25134,N_23341,N_23507);
nand U25135 (N_25135,N_23415,N_23574);
or U25136 (N_25136,N_23246,N_23971);
xor U25137 (N_25137,N_22998,N_23355);
and U25138 (N_25138,N_23723,N_23771);
xnor U25139 (N_25139,N_23015,N_23801);
nand U25140 (N_25140,N_22918,N_23529);
xnor U25141 (N_25141,N_23015,N_23951);
nand U25142 (N_25142,N_22890,N_23529);
nand U25143 (N_25143,N_22861,N_23586);
and U25144 (N_25144,N_23814,N_23165);
xnor U25145 (N_25145,N_22804,N_23525);
nor U25146 (N_25146,N_22813,N_23872);
or U25147 (N_25147,N_23415,N_22852);
and U25148 (N_25148,N_23684,N_23111);
and U25149 (N_25149,N_22867,N_23175);
or U25150 (N_25150,N_23449,N_23543);
xnor U25151 (N_25151,N_23495,N_23297);
nand U25152 (N_25152,N_23075,N_23444);
xnor U25153 (N_25153,N_22861,N_23257);
nand U25154 (N_25154,N_23618,N_23051);
nor U25155 (N_25155,N_23367,N_23554);
nor U25156 (N_25156,N_22991,N_23523);
xor U25157 (N_25157,N_23115,N_23380);
nand U25158 (N_25158,N_23201,N_23446);
nand U25159 (N_25159,N_23823,N_23478);
and U25160 (N_25160,N_23043,N_23978);
and U25161 (N_25161,N_23157,N_23830);
nor U25162 (N_25162,N_23488,N_23367);
and U25163 (N_25163,N_23050,N_23271);
nand U25164 (N_25164,N_23144,N_23090);
and U25165 (N_25165,N_23320,N_23544);
nand U25166 (N_25166,N_22905,N_23308);
nor U25167 (N_25167,N_23719,N_23118);
nand U25168 (N_25168,N_23765,N_23585);
or U25169 (N_25169,N_23943,N_23728);
nor U25170 (N_25170,N_23520,N_23357);
nor U25171 (N_25171,N_23983,N_23203);
or U25172 (N_25172,N_23828,N_23918);
xnor U25173 (N_25173,N_22987,N_23870);
and U25174 (N_25174,N_23070,N_22994);
nor U25175 (N_25175,N_23354,N_22994);
and U25176 (N_25176,N_23833,N_23123);
nand U25177 (N_25177,N_23229,N_23328);
nor U25178 (N_25178,N_23730,N_23803);
xor U25179 (N_25179,N_23717,N_23134);
nor U25180 (N_25180,N_23044,N_22960);
xor U25181 (N_25181,N_23782,N_23770);
nor U25182 (N_25182,N_22921,N_23779);
nor U25183 (N_25183,N_23052,N_23022);
xnor U25184 (N_25184,N_23091,N_23256);
nor U25185 (N_25185,N_23798,N_23351);
nand U25186 (N_25186,N_23971,N_23227);
and U25187 (N_25187,N_23592,N_23507);
nand U25188 (N_25188,N_23099,N_23053);
nand U25189 (N_25189,N_23028,N_23568);
and U25190 (N_25190,N_23159,N_22963);
nor U25191 (N_25191,N_23017,N_23014);
or U25192 (N_25192,N_23251,N_23869);
or U25193 (N_25193,N_23069,N_23599);
nor U25194 (N_25194,N_23011,N_23971);
xnor U25195 (N_25195,N_23161,N_23556);
nor U25196 (N_25196,N_23916,N_23391);
or U25197 (N_25197,N_23769,N_23360);
xor U25198 (N_25198,N_23677,N_23688);
nor U25199 (N_25199,N_23909,N_23972);
or U25200 (N_25200,N_24960,N_24115);
nor U25201 (N_25201,N_24045,N_24971);
xnor U25202 (N_25202,N_25043,N_24356);
nor U25203 (N_25203,N_24242,N_25019);
and U25204 (N_25204,N_24615,N_24667);
nor U25205 (N_25205,N_24110,N_24152);
and U25206 (N_25206,N_24124,N_24583);
or U25207 (N_25207,N_24228,N_25012);
nand U25208 (N_25208,N_24871,N_24284);
and U25209 (N_25209,N_25114,N_25130);
nor U25210 (N_25210,N_24037,N_24103);
and U25211 (N_25211,N_25091,N_24217);
and U25212 (N_25212,N_24928,N_24294);
or U25213 (N_25213,N_24264,N_24560);
and U25214 (N_25214,N_24655,N_24180);
and U25215 (N_25215,N_24307,N_24186);
and U25216 (N_25216,N_25067,N_24590);
xnor U25217 (N_25217,N_24755,N_24748);
or U25218 (N_25218,N_24163,N_24922);
and U25219 (N_25219,N_24129,N_24378);
or U25220 (N_25220,N_24641,N_24023);
nand U25221 (N_25221,N_24681,N_24568);
nor U25222 (N_25222,N_24089,N_24704);
nand U25223 (N_25223,N_24792,N_24466);
or U25224 (N_25224,N_24310,N_24467);
or U25225 (N_25225,N_24628,N_24739);
and U25226 (N_25226,N_24104,N_24738);
and U25227 (N_25227,N_24967,N_25156);
or U25228 (N_25228,N_24819,N_24489);
or U25229 (N_25229,N_24741,N_24365);
nor U25230 (N_25230,N_24977,N_24181);
and U25231 (N_25231,N_24844,N_24592);
nor U25232 (N_25232,N_25190,N_24571);
nor U25233 (N_25233,N_24085,N_24627);
or U25234 (N_25234,N_24100,N_24697);
nand U25235 (N_25235,N_24731,N_24052);
xor U25236 (N_25236,N_24506,N_24788);
and U25237 (N_25237,N_24914,N_24551);
or U25238 (N_25238,N_24652,N_24858);
nor U25239 (N_25239,N_25003,N_25016);
and U25240 (N_25240,N_25137,N_25182);
xor U25241 (N_25241,N_25142,N_24584);
nor U25242 (N_25242,N_24501,N_24268);
xor U25243 (N_25243,N_25001,N_25113);
or U25244 (N_25244,N_24328,N_25093);
nand U25245 (N_25245,N_24708,N_25079);
nor U25246 (N_25246,N_24249,N_25052);
nor U25247 (N_25247,N_24398,N_25184);
or U25248 (N_25248,N_24850,N_24505);
nor U25249 (N_25249,N_24799,N_24985);
nand U25250 (N_25250,N_25053,N_24822);
or U25251 (N_25251,N_24281,N_24892);
xnor U25252 (N_25252,N_25089,N_24435);
and U25253 (N_25253,N_24326,N_24849);
xnor U25254 (N_25254,N_24155,N_24827);
nand U25255 (N_25255,N_24083,N_24750);
or U25256 (N_25256,N_25076,N_25074);
or U25257 (N_25257,N_24255,N_24274);
xnor U25258 (N_25258,N_24904,N_24202);
and U25259 (N_25259,N_24261,N_24982);
or U25260 (N_25260,N_24962,N_24385);
or U25261 (N_25261,N_24717,N_24433);
and U25262 (N_25262,N_24753,N_24642);
nor U25263 (N_25263,N_25119,N_24425);
and U25264 (N_25264,N_24875,N_24477);
nand U25265 (N_25265,N_24724,N_24696);
nand U25266 (N_25266,N_25042,N_24051);
xor U25267 (N_25267,N_24920,N_24886);
xor U25268 (N_25268,N_25134,N_24107);
nor U25269 (N_25269,N_25180,N_24387);
nor U25270 (N_25270,N_24332,N_24431);
or U25271 (N_25271,N_25013,N_24245);
and U25272 (N_25272,N_24867,N_24057);
nand U25273 (N_25273,N_24823,N_24338);
and U25274 (N_25274,N_24493,N_24040);
and U25275 (N_25275,N_24794,N_24919);
or U25276 (N_25276,N_25021,N_24744);
and U25277 (N_25277,N_24830,N_24607);
xor U25278 (N_25278,N_24324,N_24544);
nor U25279 (N_25279,N_24013,N_25133);
nor U25280 (N_25280,N_24804,N_24291);
nor U25281 (N_25281,N_25041,N_24557);
nor U25282 (N_25282,N_24301,N_24150);
and U25283 (N_25283,N_25092,N_24727);
and U25284 (N_25284,N_24025,N_24890);
and U25285 (N_25285,N_24570,N_24815);
or U25286 (N_25286,N_24781,N_24128);
nor U25287 (N_25287,N_24063,N_25115);
xor U25288 (N_25288,N_24495,N_24721);
nand U25289 (N_25289,N_24841,N_24447);
nand U25290 (N_25290,N_24676,N_24980);
xnor U25291 (N_25291,N_24192,N_24476);
or U25292 (N_25292,N_24975,N_24730);
or U25293 (N_25293,N_25186,N_24900);
and U25294 (N_25294,N_25065,N_24578);
xor U25295 (N_25295,N_24567,N_24077);
nand U25296 (N_25296,N_24604,N_24649);
or U25297 (N_25297,N_24981,N_24771);
or U25298 (N_25298,N_24270,N_24359);
nor U25299 (N_25299,N_24066,N_24934);
and U25300 (N_25300,N_24253,N_25191);
nor U25301 (N_25301,N_24213,N_24747);
nor U25302 (N_25302,N_24295,N_24381);
xnor U25303 (N_25303,N_24836,N_24761);
xor U25304 (N_25304,N_25005,N_25108);
xor U25305 (N_25305,N_24483,N_24439);
and U25306 (N_25306,N_24327,N_24151);
or U25307 (N_25307,N_24906,N_24885);
or U25308 (N_25308,N_24701,N_24860);
xnor U25309 (N_25309,N_24436,N_24068);
xor U25310 (N_25310,N_24674,N_24248);
nand U25311 (N_25311,N_24366,N_25070);
or U25312 (N_25312,N_24108,N_25124);
or U25313 (N_25313,N_24773,N_25196);
or U25314 (N_25314,N_24139,N_24035);
nand U25315 (N_25315,N_24569,N_24322);
nor U25316 (N_25316,N_24308,N_25015);
xnor U25317 (N_25317,N_24498,N_25006);
nor U25318 (N_25318,N_24130,N_24158);
nor U25319 (N_25319,N_24137,N_24879);
nor U25320 (N_25320,N_24342,N_24972);
or U25321 (N_25321,N_24015,N_25032);
or U25322 (N_25322,N_24712,N_25116);
nand U25323 (N_25323,N_24575,N_24525);
and U25324 (N_25324,N_24599,N_24671);
xnor U25325 (N_25325,N_24621,N_24558);
and U25326 (N_25326,N_24889,N_24177);
nand U25327 (N_25327,N_24603,N_24033);
xnor U25328 (N_25328,N_24516,N_24807);
nor U25329 (N_25329,N_25028,N_24167);
or U25330 (N_25330,N_24367,N_24993);
xnor U25331 (N_25331,N_25171,N_24340);
xor U25332 (N_25332,N_24899,N_24491);
nand U25333 (N_25333,N_24208,N_24863);
nor U25334 (N_25334,N_24749,N_24648);
xnor U25335 (N_25335,N_24350,N_24053);
nor U25336 (N_25336,N_24382,N_24097);
xnor U25337 (N_25337,N_25158,N_24147);
or U25338 (N_25338,N_25029,N_25058);
nand U25339 (N_25339,N_24273,N_24050);
and U25340 (N_25340,N_24723,N_24984);
nand U25341 (N_25341,N_24663,N_24594);
and U25342 (N_25342,N_24534,N_24028);
or U25343 (N_25343,N_24757,N_25047);
or U25344 (N_25344,N_24026,N_25055);
and U25345 (N_25345,N_24669,N_24957);
nor U25346 (N_25346,N_24252,N_24496);
or U25347 (N_25347,N_24418,N_24176);
and U25348 (N_25348,N_24421,N_24715);
xnor U25349 (N_25349,N_24397,N_24591);
nor U25350 (N_25350,N_25025,N_24331);
nor U25351 (N_25351,N_25037,N_24582);
nor U25352 (N_25352,N_25034,N_24256);
or U25353 (N_25353,N_24559,N_24518);
nand U25354 (N_25354,N_24441,N_24776);
and U25355 (N_25355,N_24574,N_24358);
and U25356 (N_25356,N_25095,N_24304);
or U25357 (N_25357,N_24178,N_24758);
nand U25358 (N_25358,N_24318,N_24801);
and U25359 (N_25359,N_25144,N_24405);
or U25360 (N_25360,N_25036,N_24247);
nor U25361 (N_25361,N_24938,N_24031);
xor U25362 (N_25362,N_24692,N_24657);
or U25363 (N_25363,N_24043,N_25164);
nor U25364 (N_25364,N_24046,N_24874);
and U25365 (N_25365,N_24027,N_24532);
xnor U25366 (N_25366,N_24834,N_24924);
or U25367 (N_25367,N_24996,N_24352);
and U25368 (N_25368,N_24145,N_24321);
or U25369 (N_25369,N_25123,N_25062);
nand U25370 (N_25370,N_24945,N_24995);
nor U25371 (N_25371,N_24926,N_24872);
and U25372 (N_25372,N_24913,N_24458);
xor U25373 (N_25373,N_24054,N_25049);
or U25374 (N_25374,N_25138,N_24067);
xor U25375 (N_25375,N_24787,N_24580);
nor U25376 (N_25376,N_24062,N_24259);
nor U25377 (N_25377,N_24099,N_24653);
nand U25378 (N_25378,N_25148,N_24445);
or U25379 (N_25379,N_25050,N_25072);
nor U25380 (N_25380,N_25031,N_24207);
and U25381 (N_25381,N_24154,N_24565);
xnor U25382 (N_25382,N_25198,N_25088);
or U25383 (N_25383,N_24539,N_24878);
nor U25384 (N_25384,N_24393,N_24095);
nand U25385 (N_25385,N_24826,N_24726);
xnor U25386 (N_25386,N_25010,N_24897);
or U25387 (N_25387,N_24226,N_24702);
nor U25388 (N_25388,N_24930,N_24214);
and U25389 (N_25389,N_24537,N_24456);
or U25390 (N_25390,N_24293,N_24643);
nand U25391 (N_25391,N_24277,N_24530);
and U25392 (N_25392,N_24231,N_24891);
nand U25393 (N_25393,N_25185,N_24236);
and U25394 (N_25394,N_24825,N_24832);
nand U25395 (N_25395,N_24953,N_25097);
xor U25396 (N_25396,N_24464,N_25096);
or U25397 (N_25397,N_24585,N_24374);
xor U25398 (N_25398,N_24392,N_24379);
nor U25399 (N_25399,N_24883,N_25199);
and U25400 (N_25400,N_24636,N_24553);
nand U25401 (N_25401,N_24997,N_24243);
and U25402 (N_25402,N_24958,N_24685);
or U25403 (N_25403,N_24101,N_24184);
or U25404 (N_25404,N_25035,N_24131);
nand U25405 (N_25405,N_24665,N_24695);
and U25406 (N_25406,N_24169,N_24229);
or U25407 (N_25407,N_24556,N_24973);
or U25408 (N_25408,N_24080,N_25039);
and U25409 (N_25409,N_24682,N_24593);
and U25410 (N_25410,N_24283,N_25181);
nor U25411 (N_25411,N_24543,N_25008);
nand U25412 (N_25412,N_25018,N_24637);
nand U25413 (N_25413,N_24743,N_24372);
nor U25414 (N_25414,N_24857,N_24700);
and U25415 (N_25415,N_24437,N_24148);
xnor U25416 (N_25416,N_24514,N_24640);
nor U25417 (N_25417,N_24220,N_25112);
or U25418 (N_25418,N_24589,N_24196);
xnor U25419 (N_25419,N_24078,N_24651);
xor U25420 (N_25420,N_24762,N_24915);
xor U25421 (N_25421,N_24357,N_24198);
and U25422 (N_25422,N_24317,N_24865);
nand U25423 (N_25423,N_24851,N_24502);
and U25424 (N_25424,N_24939,N_24634);
nor U25425 (N_25425,N_24286,N_24122);
nor U25426 (N_25426,N_24468,N_24380);
and U25427 (N_25427,N_24140,N_25046);
nand U25428 (N_25428,N_24588,N_24517);
and U25429 (N_25429,N_24774,N_24542);
nor U25430 (N_25430,N_24917,N_24183);
nand U25431 (N_25431,N_24106,N_24449);
or U25432 (N_25432,N_24444,N_24497);
nand U25433 (N_25433,N_24710,N_24146);
nand U25434 (N_25434,N_24339,N_24390);
and U25435 (N_25435,N_24446,N_24361);
and U25436 (N_25436,N_24978,N_24474);
nor U25437 (N_25437,N_25038,N_25111);
or U25438 (N_25438,N_24969,N_24824);
nand U25439 (N_25439,N_24333,N_24923);
and U25440 (N_25440,N_25064,N_25085);
or U25441 (N_25441,N_24786,N_24729);
nand U25442 (N_25442,N_25135,N_25176);
and U25443 (N_25443,N_24839,N_24404);
nor U25444 (N_25444,N_24290,N_24413);
xor U25445 (N_25445,N_24803,N_24135);
xnor U25446 (N_25446,N_24086,N_25120);
nand U25447 (N_25447,N_25128,N_24098);
and U25448 (N_25448,N_24271,N_25030);
and U25449 (N_25449,N_24618,N_24805);
or U25450 (N_25450,N_24384,N_24937);
nand U25451 (N_25451,N_24706,N_25083);
nor U25452 (N_25452,N_24596,N_24126);
nor U25453 (N_25453,N_24668,N_24679);
nand U25454 (N_25454,N_25139,N_25100);
and U25455 (N_25455,N_24048,N_24531);
or U25456 (N_25456,N_24768,N_24733);
nand U25457 (N_25457,N_25140,N_24204);
or U25458 (N_25458,N_25069,N_24816);
nand U25459 (N_25459,N_24305,N_24002);
nor U25460 (N_25460,N_24864,N_24096);
nor U25461 (N_25461,N_25166,N_25109);
nand U25462 (N_25462,N_24507,N_24143);
xnor U25463 (N_25463,N_24838,N_24011);
nand U25464 (N_25464,N_24344,N_25122);
and U25465 (N_25465,N_25054,N_24699);
xnor U25466 (N_25466,N_24039,N_24470);
nor U25467 (N_25467,N_24383,N_24541);
and U25468 (N_25468,N_24267,N_24887);
nand U25469 (N_25469,N_24123,N_24888);
xnor U25470 (N_25470,N_24767,N_24395);
nor U25471 (N_25471,N_24854,N_24144);
or U25472 (N_25472,N_24116,N_24644);
nor U25473 (N_25473,N_24275,N_24313);
and U25474 (N_25474,N_24044,N_24386);
nor U25475 (N_25475,N_24989,N_24988);
and U25476 (N_25476,N_24457,N_24638);
nor U25477 (N_25477,N_24494,N_24341);
and U25478 (N_25478,N_24510,N_24772);
or U25479 (N_25479,N_24798,N_24650);
nand U25480 (N_25480,N_25170,N_24426);
xnor U25481 (N_25481,N_24209,N_24414);
nand U25482 (N_25482,N_24300,N_24992);
or U25483 (N_25483,N_24079,N_24598);
nor U25484 (N_25484,N_24478,N_24951);
and U25485 (N_25485,N_24334,N_24818);
nand U25486 (N_25486,N_24289,N_24861);
nand U25487 (N_25487,N_24954,N_24377);
nand U25488 (N_25488,N_24263,N_24241);
xor U25489 (N_25489,N_24950,N_24112);
xor U25490 (N_25490,N_24927,N_24720);
or U25491 (N_25491,N_24354,N_25084);
nand U25492 (N_25492,N_24955,N_24443);
xnor U25493 (N_25493,N_24412,N_24791);
and U25494 (N_25494,N_24533,N_24287);
or U25495 (N_25495,N_24656,N_24084);
nor U25496 (N_25496,N_24369,N_24548);
and U25497 (N_25497,N_24428,N_24072);
nand U25498 (N_25498,N_25073,N_24554);
or U25499 (N_25499,N_25009,N_24373);
xor U25500 (N_25500,N_24629,N_24908);
xor U25501 (N_25501,N_24552,N_25159);
xnor U25502 (N_25502,N_25066,N_24793);
nor U25503 (N_25503,N_24965,N_24329);
xor U25504 (N_25504,N_24216,N_24024);
xnor U25505 (N_25505,N_25132,N_24881);
and U25506 (N_25506,N_24408,N_24343);
nor U25507 (N_25507,N_24894,N_24141);
or U25508 (N_25508,N_24219,N_24610);
and U25509 (N_25509,N_25007,N_24232);
or U25510 (N_25510,N_24898,N_24309);
nor U25511 (N_25511,N_24120,N_24424);
xnor U25512 (N_25512,N_24952,N_24173);
and U25513 (N_25513,N_24417,N_24092);
nand U25514 (N_25514,N_24986,N_24512);
nand U25515 (N_25515,N_24355,N_24463);
nor U25516 (N_25516,N_24164,N_24315);
xor U25517 (N_25517,N_24740,N_24368);
or U25518 (N_25518,N_24855,N_24711);
xor U25519 (N_25519,N_24964,N_24746);
xor U25520 (N_25520,N_24728,N_25026);
xnor U25521 (N_25521,N_24735,N_24006);
xnor U25522 (N_25522,N_24940,N_24963);
or U25523 (N_25523,N_24966,N_24808);
or U25524 (N_25524,N_24111,N_25187);
nor U25525 (N_25525,N_24519,N_24500);
nor U25526 (N_25526,N_24041,N_25126);
xnor U25527 (N_25527,N_24983,N_24840);
or U25528 (N_25528,N_24484,N_25195);
xnor U25529 (N_25529,N_24422,N_24306);
or U25530 (N_25530,N_24189,N_25172);
or U25531 (N_25531,N_24873,N_25061);
and U25532 (N_25532,N_24672,N_24946);
xor U25533 (N_25533,N_24348,N_24659);
xor U25534 (N_25534,N_24225,N_24019);
or U25535 (N_25535,N_24234,N_24561);
and U25536 (N_25536,N_24427,N_24631);
or U25537 (N_25537,N_24278,N_24415);
and U25538 (N_25538,N_24763,N_24809);
xor U25539 (N_25539,N_24215,N_24550);
and U25540 (N_25540,N_24959,N_24018);
nor U25541 (N_25541,N_24754,N_24736);
and U25542 (N_25542,N_24288,N_24479);
nand U25543 (N_25543,N_24707,N_25033);
xor U25544 (N_25544,N_24187,N_25082);
and U25545 (N_25545,N_24555,N_24311);
or U25546 (N_25546,N_24943,N_24075);
and U25547 (N_25547,N_24769,N_24626);
or U25548 (N_25548,N_25002,N_24316);
or U25549 (N_25549,N_24410,N_24527);
or U25550 (N_25550,N_24499,N_25121);
nand U25551 (N_25551,N_24438,N_24759);
and U25552 (N_25552,N_24779,N_24684);
or U25553 (N_25553,N_24901,N_25004);
nor U25554 (N_25554,N_24459,N_24683);
or U25555 (N_25555,N_24933,N_24713);
and U25556 (N_25556,N_24709,N_24814);
nand U25557 (N_25557,N_24511,N_25068);
and U25558 (N_25558,N_24703,N_24602);
and U25559 (N_25559,N_25169,N_25051);
nand U25560 (N_25560,N_24279,N_24581);
xnor U25561 (N_25561,N_24576,N_24921);
xor U25562 (N_25562,N_25014,N_25071);
nand U25563 (N_25563,N_24292,N_25057);
or U25564 (N_25564,N_25127,N_24999);
and U25565 (N_25565,N_24869,N_24998);
xnor U25566 (N_25566,N_24087,N_24893);
or U25567 (N_25567,N_24925,N_24817);
nand U25568 (N_25568,N_25101,N_24388);
nand U25569 (N_25569,N_24070,N_24742);
or U25570 (N_25570,N_24162,N_24007);
nor U25571 (N_25571,N_25175,N_24091);
and U25572 (N_25572,N_24828,N_25023);
nand U25573 (N_25573,N_24948,N_24910);
or U25574 (N_25574,N_24302,N_24325);
and U25575 (N_25575,N_24811,N_24775);
xnor U25576 (N_25576,N_24931,N_24175);
xnor U25577 (N_25577,N_24401,N_25174);
and U25578 (N_25578,N_24481,N_24406);
and U25579 (N_25579,N_24462,N_24471);
nand U25580 (N_25580,N_24991,N_24632);
nand U25581 (N_25581,N_24005,N_24718);
xnor U25582 (N_25582,N_24852,N_24034);
xnor U25583 (N_25583,N_24090,N_24064);
and U25584 (N_25584,N_25078,N_24635);
and U25585 (N_25585,N_24764,N_25147);
and U25586 (N_25586,N_24990,N_24944);
xor U25587 (N_25587,N_24237,N_24142);
nor U25588 (N_25588,N_24136,N_24929);
and U25589 (N_25589,N_25188,N_24949);
and U25590 (N_25590,N_24513,N_24161);
xor U25591 (N_25591,N_24210,N_24319);
nor U25592 (N_25592,N_24895,N_24349);
and U25593 (N_25593,N_24250,N_24276);
and U25594 (N_25594,N_24687,N_24535);
or U25595 (N_25595,N_24876,N_24257);
nand U25596 (N_25596,N_24778,N_24974);
nor U25597 (N_25597,N_24630,N_24272);
nand U25598 (N_25598,N_24639,N_24492);
nor U25599 (N_25599,N_24932,N_24536);
or U25600 (N_25600,N_24093,N_24049);
nor U25601 (N_25601,N_25020,N_25048);
xnor U25602 (N_25602,N_24239,N_24391);
xor U25603 (N_25603,N_24529,N_25192);
or U25604 (N_25604,N_24074,N_24847);
nand U25605 (N_25605,N_24058,N_24299);
or U25606 (N_25606,N_24722,N_24453);
xor U25607 (N_25607,N_24469,N_24012);
nand U25608 (N_25608,N_25024,N_25077);
xnor U25609 (N_25609,N_24664,N_25125);
or U25610 (N_25610,N_24407,N_24625);
xor U25611 (N_25611,N_24573,N_24780);
or U25612 (N_25612,N_24454,N_24546);
nand U25613 (N_25613,N_24191,N_24364);
nand U25614 (N_25614,N_24347,N_25117);
or U25615 (N_25615,N_24800,N_24363);
and U25616 (N_25616,N_24486,N_25178);
nand U25617 (N_25617,N_24320,N_24118);
nor U25618 (N_25618,N_25143,N_24235);
and U25619 (N_25619,N_24201,N_25163);
xnor U25620 (N_25620,N_24677,N_24218);
and U25621 (N_25621,N_24662,N_24430);
nor U25622 (N_25622,N_24605,N_24022);
and U25623 (N_25623,N_24166,N_24416);
or U25624 (N_25624,N_24109,N_25161);
or U25625 (N_25625,N_25017,N_24689);
or U25626 (N_25626,N_24688,N_25000);
and U25627 (N_25627,N_24149,N_24523);
xnor U25628 (N_25628,N_24094,N_24419);
nor U25629 (N_25629,N_24224,N_25150);
xnor U25630 (N_25630,N_24482,N_24601);
nand U25631 (N_25631,N_24509,N_24911);
nor U25632 (N_25632,N_25165,N_25173);
and U25633 (N_25633,N_25154,N_24624);
nand U25634 (N_25634,N_24056,N_24646);
or U25635 (N_25635,N_24829,N_24200);
or U25636 (N_25636,N_24918,N_24055);
and U25637 (N_25637,N_24678,N_24528);
nor U25638 (N_25638,N_25027,N_25087);
nand U25639 (N_25639,N_24038,N_24784);
xnor U25640 (N_25640,N_24812,N_24994);
xnor U25641 (N_25641,N_24572,N_24030);
and U25642 (N_25642,N_24612,N_24008);
or U25643 (N_25643,N_24705,N_24698);
and U25644 (N_25644,N_24193,N_25099);
xor U25645 (N_25645,N_25167,N_24777);
nor U25646 (N_25646,N_24936,N_24783);
xor U25647 (N_25647,N_24345,N_25063);
and U25648 (N_25648,N_25136,N_24199);
xor U25649 (N_25649,N_24153,N_24907);
nand U25650 (N_25650,N_25081,N_24620);
and U25651 (N_25651,N_24460,N_25153);
nor U25652 (N_25652,N_24206,N_24691);
or U25653 (N_25653,N_24138,N_24595);
and U25654 (N_25654,N_24884,N_24538);
xor U25655 (N_25655,N_24790,N_24654);
xnor U25656 (N_25656,N_24195,N_24473);
and U25657 (N_25657,N_24323,N_24508);
and U25658 (N_25658,N_24670,N_24760);
nand U25659 (N_25659,N_24194,N_24061);
nor U25660 (N_25660,N_24611,N_24905);
nor U25661 (N_25661,N_24848,N_25160);
nand U25662 (N_25662,N_24719,N_24227);
or U25663 (N_25663,N_25131,N_24756);
xnor U25664 (N_25664,N_24912,N_24597);
nor U25665 (N_25665,N_24125,N_25040);
and U25666 (N_25666,N_24240,N_24335);
or U25667 (N_25667,N_25162,N_24622);
nand U25668 (N_25668,N_24806,N_24360);
nor U25669 (N_25669,N_24238,N_24614);
or U25670 (N_25670,N_24411,N_25145);
and U25671 (N_25671,N_24396,N_24586);
or U25672 (N_25672,N_24452,N_24262);
nor U25673 (N_25673,N_25179,N_24114);
and U25674 (N_25674,N_24880,N_24842);
or U25675 (N_25675,N_24203,N_24172);
and U25676 (N_25676,N_24694,N_24402);
nor U25677 (N_25677,N_24020,N_24480);
and U25678 (N_25678,N_24269,N_24001);
and U25679 (N_25679,N_24549,N_24947);
xnor U25680 (N_25680,N_24420,N_24609);
nor U25681 (N_25681,N_24613,N_24297);
xor U25682 (N_25682,N_25103,N_24060);
or U25683 (N_25683,N_24156,N_24956);
nand U25684 (N_25684,N_24003,N_24862);
nor U25685 (N_25685,N_24076,N_24902);
nand U25686 (N_25686,N_24521,N_24190);
and U25687 (N_25687,N_25060,N_25168);
nor U25688 (N_25688,N_24976,N_24680);
xnor U25689 (N_25689,N_25044,N_24211);
or U25690 (N_25690,N_25194,N_24725);
nor U25691 (N_25691,N_24440,N_24221);
nand U25692 (N_25692,N_24059,N_24014);
or U25693 (N_25693,N_24942,N_24265);
xnor U25694 (N_25694,N_24314,N_24617);
or U25695 (N_25695,N_24409,N_24222);
and U25696 (N_25696,N_24258,N_24119);
and U25697 (N_25697,N_25011,N_24647);
and U25698 (N_25698,N_24429,N_24547);
nor U25699 (N_25699,N_24021,N_24843);
nor U25700 (N_25700,N_24520,N_24540);
nand U25701 (N_25701,N_24587,N_24423);
nand U25702 (N_25702,N_24485,N_24065);
nand U25703 (N_25703,N_24337,N_24102);
and U25704 (N_25704,N_25110,N_24660);
nor U25705 (N_25705,N_24661,N_24434);
nor U25706 (N_25706,N_24903,N_24159);
xnor U25707 (N_25707,N_25090,N_24400);
or U25708 (N_25708,N_24403,N_24675);
nor U25709 (N_25709,N_24600,N_24009);
nor U25710 (N_25710,N_24353,N_24782);
xor U25711 (N_25711,N_24577,N_24205);
xnor U25712 (N_25712,N_24877,N_24503);
and U25713 (N_25713,N_24036,N_24916);
nand U25714 (N_25714,N_24690,N_24029);
nand U25715 (N_25715,N_24526,N_24047);
or U25716 (N_25716,N_25107,N_25106);
nand U25717 (N_25717,N_24370,N_24770);
and U25718 (N_25718,N_24821,N_24088);
nand U25719 (N_25719,N_25141,N_24608);
or U25720 (N_25720,N_24351,N_24017);
xnor U25721 (N_25721,N_24371,N_25045);
and U25722 (N_25722,N_24032,N_24069);
nor U25723 (N_25723,N_24802,N_25149);
nand U25724 (N_25724,N_24968,N_24185);
or U25725 (N_25725,N_24515,N_24686);
xnor U25726 (N_25726,N_25146,N_24935);
nand U25727 (N_25727,N_24168,N_25118);
and U25728 (N_25728,N_24266,N_24455);
or U25729 (N_25729,N_24716,N_24254);
and U25730 (N_25730,N_24859,N_24961);
nor U25731 (N_25731,N_24896,N_24837);
nor U25732 (N_25732,N_24171,N_24941);
xor U25733 (N_25733,N_24465,N_24566);
and U25734 (N_25734,N_25102,N_24562);
and U25735 (N_25735,N_24165,N_24450);
nand U25736 (N_25736,N_24170,N_25080);
nand U25737 (N_25737,N_24796,N_25197);
xor U25738 (N_25738,N_24745,N_24000);
nor U25739 (N_25739,N_24174,N_24432);
and U25740 (N_25740,N_24752,N_25129);
or U25741 (N_25741,N_25105,N_25151);
and U25742 (N_25742,N_24789,N_24448);
nand U25743 (N_25743,N_24765,N_25189);
and U25744 (N_25744,N_24833,N_24673);
or U25745 (N_25745,N_24524,N_24797);
and U25746 (N_25746,N_24490,N_24734);
xnor U25747 (N_25747,N_24737,N_24522);
or U25748 (N_25748,N_24545,N_25155);
and U25749 (N_25749,N_24223,N_25183);
nand U25750 (N_25750,N_24298,N_24285);
nor U25751 (N_25751,N_24389,N_25152);
nand U25752 (N_25752,N_24251,N_24134);
nand U25753 (N_25753,N_24472,N_24987);
xnor U25754 (N_25754,N_24071,N_24579);
nand U25755 (N_25755,N_24362,N_24645);
and U25756 (N_25756,N_25056,N_24212);
nand U25757 (N_25757,N_24113,N_24246);
xnor U25758 (N_25758,N_24845,N_24751);
nand U25759 (N_25759,N_24813,N_24606);
or U25760 (N_25760,N_24188,N_25098);
nand U25761 (N_25761,N_24244,N_24127);
nand U25762 (N_25762,N_24346,N_24133);
xnor U25763 (N_25763,N_24399,N_24616);
xor U25764 (N_25764,N_24121,N_24658);
nand U25765 (N_25765,N_24820,N_24004);
and U25766 (N_25766,N_24846,N_24280);
nand U25767 (N_25767,N_24623,N_24233);
nand U25768 (N_25768,N_24666,N_24081);
nor U25769 (N_25769,N_24870,N_24714);
nor U25770 (N_25770,N_24016,N_24132);
nand U25771 (N_25771,N_25104,N_24442);
nand U25772 (N_25772,N_25094,N_24461);
or U25773 (N_25773,N_24451,N_24866);
or U25774 (N_25774,N_24810,N_25177);
or U25775 (N_25775,N_24766,N_24282);
or U25776 (N_25776,N_24785,N_24979);
or U25777 (N_25777,N_25059,N_24197);
nand U25778 (N_25778,N_24260,N_24182);
and U25779 (N_25779,N_24312,N_24868);
nor U25780 (N_25780,N_24853,N_24619);
nand U25781 (N_25781,N_24487,N_25022);
nor U25782 (N_25782,N_25075,N_25086);
nor U25783 (N_25783,N_24330,N_24160);
or U25784 (N_25784,N_24831,N_24179);
nor U25785 (N_25785,N_24693,N_24882);
xor U25786 (N_25786,N_24504,N_24376);
and U25787 (N_25787,N_24835,N_24564);
or U25788 (N_25788,N_24296,N_24394);
and U25789 (N_25789,N_24970,N_24488);
nand U25790 (N_25790,N_24856,N_24375);
nor U25791 (N_25791,N_24336,N_25193);
nand U25792 (N_25792,N_24073,N_24475);
xor U25793 (N_25793,N_24230,N_24563);
nor U25794 (N_25794,N_24117,N_24732);
or U25795 (N_25795,N_24042,N_24909);
or U25796 (N_25796,N_24010,N_24105);
nand U25797 (N_25797,N_24795,N_24082);
nor U25798 (N_25798,N_25157,N_24303);
and U25799 (N_25799,N_24157,N_24633);
xor U25800 (N_25800,N_24942,N_24218);
and U25801 (N_25801,N_25008,N_24629);
and U25802 (N_25802,N_24025,N_25049);
and U25803 (N_25803,N_24869,N_24760);
nand U25804 (N_25804,N_24671,N_24451);
nand U25805 (N_25805,N_24645,N_25155);
xnor U25806 (N_25806,N_25099,N_25106);
nor U25807 (N_25807,N_24915,N_25145);
xnor U25808 (N_25808,N_24409,N_24141);
nor U25809 (N_25809,N_24289,N_24833);
nand U25810 (N_25810,N_24659,N_24531);
and U25811 (N_25811,N_24746,N_24523);
or U25812 (N_25812,N_24507,N_24236);
xnor U25813 (N_25813,N_24011,N_24405);
or U25814 (N_25814,N_24173,N_24248);
or U25815 (N_25815,N_24180,N_24623);
or U25816 (N_25816,N_24021,N_25004);
and U25817 (N_25817,N_24644,N_24357);
xor U25818 (N_25818,N_24913,N_24251);
nor U25819 (N_25819,N_24354,N_25121);
xnor U25820 (N_25820,N_24733,N_25030);
nor U25821 (N_25821,N_24086,N_24150);
or U25822 (N_25822,N_24162,N_24327);
and U25823 (N_25823,N_25175,N_24169);
nor U25824 (N_25824,N_24007,N_24866);
xnor U25825 (N_25825,N_24117,N_24158);
nor U25826 (N_25826,N_25196,N_24605);
nand U25827 (N_25827,N_24222,N_24044);
nand U25828 (N_25828,N_24291,N_24847);
nand U25829 (N_25829,N_24694,N_24979);
or U25830 (N_25830,N_24588,N_24140);
and U25831 (N_25831,N_24080,N_24598);
and U25832 (N_25832,N_24093,N_24727);
nand U25833 (N_25833,N_24836,N_24719);
xor U25834 (N_25834,N_24025,N_24368);
and U25835 (N_25835,N_24821,N_24916);
nand U25836 (N_25836,N_24620,N_24860);
xor U25837 (N_25837,N_24568,N_24415);
nor U25838 (N_25838,N_24252,N_24247);
nand U25839 (N_25839,N_24592,N_24901);
nor U25840 (N_25840,N_24264,N_24900);
and U25841 (N_25841,N_24435,N_24995);
xnor U25842 (N_25842,N_24701,N_24313);
nor U25843 (N_25843,N_24560,N_24937);
nor U25844 (N_25844,N_24847,N_25042);
and U25845 (N_25845,N_24263,N_24522);
or U25846 (N_25846,N_24166,N_24462);
nand U25847 (N_25847,N_24492,N_24329);
and U25848 (N_25848,N_24168,N_24778);
nand U25849 (N_25849,N_24578,N_24091);
or U25850 (N_25850,N_24561,N_24069);
nand U25851 (N_25851,N_24800,N_24386);
nor U25852 (N_25852,N_24297,N_24850);
nor U25853 (N_25853,N_24497,N_24936);
or U25854 (N_25854,N_24687,N_24581);
nand U25855 (N_25855,N_24490,N_24447);
nand U25856 (N_25856,N_24798,N_24749);
nand U25857 (N_25857,N_24721,N_24705);
nand U25858 (N_25858,N_25182,N_24015);
or U25859 (N_25859,N_24655,N_24087);
or U25860 (N_25860,N_24093,N_24625);
and U25861 (N_25861,N_24594,N_25198);
or U25862 (N_25862,N_24323,N_24756);
nor U25863 (N_25863,N_24893,N_24113);
nand U25864 (N_25864,N_24486,N_24876);
and U25865 (N_25865,N_25088,N_24358);
and U25866 (N_25866,N_24203,N_24819);
or U25867 (N_25867,N_24118,N_24651);
nand U25868 (N_25868,N_24383,N_24596);
xor U25869 (N_25869,N_24916,N_24458);
xnor U25870 (N_25870,N_24164,N_25188);
and U25871 (N_25871,N_24641,N_24260);
and U25872 (N_25872,N_25042,N_24268);
and U25873 (N_25873,N_24373,N_24840);
xnor U25874 (N_25874,N_24071,N_24330);
nor U25875 (N_25875,N_24114,N_24305);
and U25876 (N_25876,N_24262,N_25093);
nor U25877 (N_25877,N_24837,N_25077);
xnor U25878 (N_25878,N_24177,N_25061);
or U25879 (N_25879,N_24385,N_24051);
nor U25880 (N_25880,N_24692,N_24342);
or U25881 (N_25881,N_24726,N_24927);
or U25882 (N_25882,N_24978,N_25061);
xnor U25883 (N_25883,N_24642,N_24183);
or U25884 (N_25884,N_24359,N_24861);
nand U25885 (N_25885,N_24258,N_24394);
and U25886 (N_25886,N_24891,N_24397);
or U25887 (N_25887,N_25127,N_24161);
and U25888 (N_25888,N_25167,N_24552);
xor U25889 (N_25889,N_24427,N_24240);
xor U25890 (N_25890,N_25072,N_24544);
nor U25891 (N_25891,N_24673,N_24239);
xor U25892 (N_25892,N_24095,N_24700);
xnor U25893 (N_25893,N_24490,N_24899);
and U25894 (N_25894,N_24313,N_24398);
or U25895 (N_25895,N_24489,N_24793);
and U25896 (N_25896,N_24693,N_24507);
xor U25897 (N_25897,N_25047,N_25074);
nor U25898 (N_25898,N_24752,N_24467);
or U25899 (N_25899,N_24937,N_24439);
nand U25900 (N_25900,N_25046,N_24337);
nand U25901 (N_25901,N_25036,N_24744);
or U25902 (N_25902,N_24145,N_24425);
nand U25903 (N_25903,N_25171,N_24806);
nand U25904 (N_25904,N_24628,N_24176);
or U25905 (N_25905,N_25139,N_24830);
and U25906 (N_25906,N_25067,N_24876);
xnor U25907 (N_25907,N_24892,N_24696);
nand U25908 (N_25908,N_24039,N_25149);
nor U25909 (N_25909,N_25110,N_24643);
and U25910 (N_25910,N_24057,N_24199);
or U25911 (N_25911,N_24213,N_24707);
nor U25912 (N_25912,N_25191,N_24659);
xor U25913 (N_25913,N_24556,N_24170);
xor U25914 (N_25914,N_24465,N_24070);
nor U25915 (N_25915,N_24968,N_24860);
xor U25916 (N_25916,N_24337,N_24064);
and U25917 (N_25917,N_25014,N_25174);
nor U25918 (N_25918,N_25172,N_25073);
and U25919 (N_25919,N_25133,N_24815);
nand U25920 (N_25920,N_24790,N_25022);
or U25921 (N_25921,N_25130,N_24424);
nor U25922 (N_25922,N_25162,N_24965);
and U25923 (N_25923,N_24425,N_24371);
nor U25924 (N_25924,N_24366,N_24298);
nor U25925 (N_25925,N_24719,N_24705);
nor U25926 (N_25926,N_24458,N_24379);
and U25927 (N_25927,N_24188,N_24139);
and U25928 (N_25928,N_25076,N_24564);
and U25929 (N_25929,N_24547,N_24952);
xor U25930 (N_25930,N_24999,N_24834);
and U25931 (N_25931,N_24460,N_24569);
xnor U25932 (N_25932,N_24700,N_24198);
nand U25933 (N_25933,N_25175,N_24165);
or U25934 (N_25934,N_24477,N_24741);
or U25935 (N_25935,N_24149,N_24178);
and U25936 (N_25936,N_24637,N_24122);
and U25937 (N_25937,N_24937,N_24538);
xor U25938 (N_25938,N_24503,N_24615);
and U25939 (N_25939,N_24261,N_24907);
nor U25940 (N_25940,N_25172,N_24610);
xor U25941 (N_25941,N_25165,N_24920);
or U25942 (N_25942,N_24286,N_24721);
nor U25943 (N_25943,N_24311,N_24238);
nor U25944 (N_25944,N_24954,N_24093);
nor U25945 (N_25945,N_24599,N_24263);
or U25946 (N_25946,N_24722,N_24000);
and U25947 (N_25947,N_24357,N_25160);
nor U25948 (N_25948,N_25066,N_25179);
nand U25949 (N_25949,N_24462,N_25081);
and U25950 (N_25950,N_24981,N_24366);
or U25951 (N_25951,N_24348,N_24029);
xnor U25952 (N_25952,N_24076,N_24921);
xnor U25953 (N_25953,N_24986,N_24935);
nand U25954 (N_25954,N_24984,N_25112);
or U25955 (N_25955,N_24038,N_24230);
nor U25956 (N_25956,N_24401,N_24772);
nand U25957 (N_25957,N_24990,N_24709);
or U25958 (N_25958,N_24873,N_24900);
or U25959 (N_25959,N_24224,N_24469);
nand U25960 (N_25960,N_25128,N_24868);
or U25961 (N_25961,N_24745,N_24773);
or U25962 (N_25962,N_25067,N_24145);
xnor U25963 (N_25963,N_24214,N_24305);
nor U25964 (N_25964,N_24384,N_24079);
or U25965 (N_25965,N_24794,N_24462);
xnor U25966 (N_25966,N_25004,N_25156);
xor U25967 (N_25967,N_24636,N_24570);
nor U25968 (N_25968,N_25081,N_24966);
and U25969 (N_25969,N_25067,N_24991);
xor U25970 (N_25970,N_24419,N_25086);
nand U25971 (N_25971,N_24796,N_24597);
xor U25972 (N_25972,N_24705,N_24838);
nand U25973 (N_25973,N_24815,N_24392);
nand U25974 (N_25974,N_24351,N_24230);
nand U25975 (N_25975,N_24207,N_24564);
nor U25976 (N_25976,N_24443,N_24084);
or U25977 (N_25977,N_24943,N_24142);
nor U25978 (N_25978,N_24326,N_24089);
nand U25979 (N_25979,N_24145,N_24434);
xnor U25980 (N_25980,N_24781,N_24362);
nand U25981 (N_25981,N_25187,N_24836);
or U25982 (N_25982,N_24801,N_24374);
nand U25983 (N_25983,N_25016,N_24677);
xnor U25984 (N_25984,N_24975,N_24726);
nor U25985 (N_25985,N_24583,N_24201);
and U25986 (N_25986,N_24679,N_24706);
nor U25987 (N_25987,N_24932,N_25005);
or U25988 (N_25988,N_24941,N_24766);
or U25989 (N_25989,N_25005,N_24236);
or U25990 (N_25990,N_25192,N_24989);
nand U25991 (N_25991,N_25170,N_24635);
and U25992 (N_25992,N_24680,N_24276);
and U25993 (N_25993,N_24577,N_24772);
xor U25994 (N_25994,N_25131,N_24322);
or U25995 (N_25995,N_24939,N_24086);
xor U25996 (N_25996,N_24268,N_24094);
nand U25997 (N_25997,N_24045,N_24682);
nand U25998 (N_25998,N_24675,N_24871);
nor U25999 (N_25999,N_24855,N_24832);
or U26000 (N_26000,N_25102,N_24144);
or U26001 (N_26001,N_25104,N_24208);
or U26002 (N_26002,N_24562,N_24978);
nand U26003 (N_26003,N_24209,N_24440);
xor U26004 (N_26004,N_24223,N_24315);
or U26005 (N_26005,N_24214,N_25076);
or U26006 (N_26006,N_25019,N_24109);
or U26007 (N_26007,N_24665,N_25104);
xnor U26008 (N_26008,N_24501,N_24412);
or U26009 (N_26009,N_24723,N_24806);
nor U26010 (N_26010,N_24101,N_24059);
or U26011 (N_26011,N_24239,N_25102);
nand U26012 (N_26012,N_24394,N_25043);
or U26013 (N_26013,N_24006,N_25044);
nor U26014 (N_26014,N_24870,N_24602);
xnor U26015 (N_26015,N_24228,N_25109);
xor U26016 (N_26016,N_24612,N_24614);
xnor U26017 (N_26017,N_25128,N_24862);
and U26018 (N_26018,N_24970,N_24281);
nand U26019 (N_26019,N_24354,N_24291);
or U26020 (N_26020,N_25187,N_24186);
nand U26021 (N_26021,N_24160,N_24205);
nor U26022 (N_26022,N_24004,N_24504);
or U26023 (N_26023,N_24990,N_24590);
and U26024 (N_26024,N_24278,N_24442);
nand U26025 (N_26025,N_24158,N_24697);
or U26026 (N_26026,N_24059,N_25127);
xnor U26027 (N_26027,N_24893,N_24326);
nor U26028 (N_26028,N_25108,N_24834);
nor U26029 (N_26029,N_24162,N_24225);
or U26030 (N_26030,N_24700,N_24694);
nand U26031 (N_26031,N_24708,N_24082);
and U26032 (N_26032,N_24626,N_24349);
xor U26033 (N_26033,N_25163,N_24125);
xnor U26034 (N_26034,N_24344,N_24802);
and U26035 (N_26035,N_24990,N_24229);
nand U26036 (N_26036,N_24521,N_24055);
and U26037 (N_26037,N_24202,N_24934);
xnor U26038 (N_26038,N_24732,N_24120);
or U26039 (N_26039,N_25052,N_24571);
nand U26040 (N_26040,N_24084,N_24796);
nor U26041 (N_26041,N_24014,N_24515);
xnor U26042 (N_26042,N_24066,N_24075);
and U26043 (N_26043,N_24510,N_24970);
or U26044 (N_26044,N_24814,N_24669);
and U26045 (N_26045,N_24498,N_24821);
nand U26046 (N_26046,N_24493,N_24940);
and U26047 (N_26047,N_24257,N_24326);
nand U26048 (N_26048,N_24667,N_24506);
nor U26049 (N_26049,N_24574,N_24281);
xnor U26050 (N_26050,N_25165,N_25124);
nand U26051 (N_26051,N_24462,N_24103);
or U26052 (N_26052,N_24903,N_24466);
nand U26053 (N_26053,N_24497,N_24302);
xor U26054 (N_26054,N_25010,N_24419);
xnor U26055 (N_26055,N_24616,N_24621);
nand U26056 (N_26056,N_24033,N_25195);
and U26057 (N_26057,N_25196,N_24238);
nand U26058 (N_26058,N_24167,N_25106);
xnor U26059 (N_26059,N_24320,N_24414);
nor U26060 (N_26060,N_25169,N_24556);
xor U26061 (N_26061,N_24460,N_24391);
nor U26062 (N_26062,N_24246,N_24854);
or U26063 (N_26063,N_24709,N_24049);
and U26064 (N_26064,N_24816,N_24338);
nor U26065 (N_26065,N_24211,N_25075);
nand U26066 (N_26066,N_24509,N_24512);
nand U26067 (N_26067,N_25031,N_25079);
nand U26068 (N_26068,N_24121,N_24874);
or U26069 (N_26069,N_24555,N_24904);
or U26070 (N_26070,N_24810,N_24520);
and U26071 (N_26071,N_25090,N_25166);
nand U26072 (N_26072,N_24465,N_24148);
and U26073 (N_26073,N_24263,N_24588);
and U26074 (N_26074,N_24403,N_24412);
and U26075 (N_26075,N_24827,N_25186);
nor U26076 (N_26076,N_24009,N_24261);
or U26077 (N_26077,N_25137,N_24065);
and U26078 (N_26078,N_24038,N_24159);
xor U26079 (N_26079,N_24367,N_24681);
nand U26080 (N_26080,N_24688,N_25016);
xor U26081 (N_26081,N_24941,N_25018);
or U26082 (N_26082,N_24515,N_24022);
nand U26083 (N_26083,N_24388,N_24571);
xor U26084 (N_26084,N_24523,N_24167);
nor U26085 (N_26085,N_24869,N_24639);
or U26086 (N_26086,N_24979,N_25135);
xor U26087 (N_26087,N_24677,N_24679);
and U26088 (N_26088,N_24681,N_24197);
nand U26089 (N_26089,N_24997,N_24667);
nand U26090 (N_26090,N_24562,N_24314);
xor U26091 (N_26091,N_24455,N_24711);
and U26092 (N_26092,N_24587,N_24303);
xor U26093 (N_26093,N_24977,N_24170);
or U26094 (N_26094,N_25144,N_24261);
or U26095 (N_26095,N_25026,N_24687);
and U26096 (N_26096,N_24643,N_24103);
or U26097 (N_26097,N_24122,N_24173);
nand U26098 (N_26098,N_24544,N_25151);
or U26099 (N_26099,N_24373,N_24910);
and U26100 (N_26100,N_24211,N_24058);
xor U26101 (N_26101,N_25084,N_24688);
nor U26102 (N_26102,N_24156,N_24305);
xnor U26103 (N_26103,N_24957,N_24624);
nand U26104 (N_26104,N_24989,N_24358);
and U26105 (N_26105,N_24478,N_24346);
nand U26106 (N_26106,N_24297,N_24512);
xnor U26107 (N_26107,N_24248,N_24761);
nor U26108 (N_26108,N_24733,N_24565);
nand U26109 (N_26109,N_24341,N_24908);
or U26110 (N_26110,N_24683,N_24493);
nand U26111 (N_26111,N_24496,N_24044);
nand U26112 (N_26112,N_24269,N_24745);
and U26113 (N_26113,N_24905,N_24247);
nand U26114 (N_26114,N_24544,N_24971);
and U26115 (N_26115,N_24722,N_24276);
or U26116 (N_26116,N_24406,N_25178);
or U26117 (N_26117,N_25125,N_24330);
nand U26118 (N_26118,N_24590,N_25135);
nand U26119 (N_26119,N_25080,N_24671);
xor U26120 (N_26120,N_24681,N_24513);
or U26121 (N_26121,N_24318,N_24955);
xor U26122 (N_26122,N_24180,N_24731);
xnor U26123 (N_26123,N_24247,N_24258);
nand U26124 (N_26124,N_25104,N_25123);
nor U26125 (N_26125,N_24504,N_24567);
and U26126 (N_26126,N_25005,N_24282);
nand U26127 (N_26127,N_25196,N_24695);
nand U26128 (N_26128,N_24718,N_24919);
xor U26129 (N_26129,N_24403,N_24829);
xnor U26130 (N_26130,N_24510,N_24741);
or U26131 (N_26131,N_24245,N_24309);
nor U26132 (N_26132,N_24794,N_24854);
or U26133 (N_26133,N_24958,N_24394);
xnor U26134 (N_26134,N_24762,N_24619);
or U26135 (N_26135,N_24851,N_24685);
xor U26136 (N_26136,N_24464,N_24202);
nor U26137 (N_26137,N_24923,N_24610);
nand U26138 (N_26138,N_24258,N_24561);
nand U26139 (N_26139,N_24841,N_24863);
and U26140 (N_26140,N_24194,N_24598);
xor U26141 (N_26141,N_24154,N_24708);
nand U26142 (N_26142,N_24560,N_25076);
xnor U26143 (N_26143,N_24592,N_24257);
or U26144 (N_26144,N_24798,N_24866);
nor U26145 (N_26145,N_24889,N_24319);
xnor U26146 (N_26146,N_24323,N_24235);
and U26147 (N_26147,N_25115,N_24931);
or U26148 (N_26148,N_24550,N_24777);
nor U26149 (N_26149,N_25011,N_24121);
and U26150 (N_26150,N_25000,N_25093);
nand U26151 (N_26151,N_24972,N_24176);
and U26152 (N_26152,N_24666,N_24510);
nor U26153 (N_26153,N_24527,N_24665);
xnor U26154 (N_26154,N_24056,N_24721);
nand U26155 (N_26155,N_24604,N_25031);
or U26156 (N_26156,N_24581,N_24407);
or U26157 (N_26157,N_24346,N_24744);
nor U26158 (N_26158,N_24868,N_25124);
xor U26159 (N_26159,N_24031,N_24334);
xnor U26160 (N_26160,N_25095,N_25176);
nor U26161 (N_26161,N_25146,N_25043);
nor U26162 (N_26162,N_24087,N_24964);
or U26163 (N_26163,N_25150,N_24960);
nor U26164 (N_26164,N_24770,N_24389);
or U26165 (N_26165,N_25125,N_24049);
nor U26166 (N_26166,N_24034,N_24050);
xnor U26167 (N_26167,N_24358,N_24602);
and U26168 (N_26168,N_24039,N_24090);
nor U26169 (N_26169,N_24014,N_25037);
xor U26170 (N_26170,N_24284,N_25054);
nor U26171 (N_26171,N_24436,N_24264);
nand U26172 (N_26172,N_24066,N_24197);
xnor U26173 (N_26173,N_24107,N_25064);
or U26174 (N_26174,N_24051,N_25182);
and U26175 (N_26175,N_24094,N_24479);
nand U26176 (N_26176,N_24623,N_24226);
xor U26177 (N_26177,N_25179,N_24426);
nor U26178 (N_26178,N_24651,N_24329);
nor U26179 (N_26179,N_24418,N_24069);
nor U26180 (N_26180,N_24814,N_24033);
nor U26181 (N_26181,N_24530,N_24179);
and U26182 (N_26182,N_25151,N_24512);
and U26183 (N_26183,N_25150,N_24474);
nand U26184 (N_26184,N_24060,N_24541);
or U26185 (N_26185,N_24383,N_24117);
or U26186 (N_26186,N_25023,N_24365);
or U26187 (N_26187,N_24780,N_25061);
nor U26188 (N_26188,N_25087,N_24750);
nand U26189 (N_26189,N_24080,N_24078);
nand U26190 (N_26190,N_24936,N_24399);
and U26191 (N_26191,N_24019,N_24904);
or U26192 (N_26192,N_25151,N_24160);
xnor U26193 (N_26193,N_24583,N_24270);
and U26194 (N_26194,N_25101,N_24068);
nor U26195 (N_26195,N_24243,N_25168);
xnor U26196 (N_26196,N_24130,N_24208);
nand U26197 (N_26197,N_24108,N_24528);
and U26198 (N_26198,N_24833,N_24019);
or U26199 (N_26199,N_24594,N_24029);
or U26200 (N_26200,N_24617,N_24555);
and U26201 (N_26201,N_24896,N_25067);
and U26202 (N_26202,N_24201,N_24614);
xor U26203 (N_26203,N_25128,N_25115);
xor U26204 (N_26204,N_24215,N_24177);
or U26205 (N_26205,N_24748,N_24542);
nor U26206 (N_26206,N_24732,N_24461);
nor U26207 (N_26207,N_24079,N_24186);
nand U26208 (N_26208,N_24097,N_24549);
nand U26209 (N_26209,N_24614,N_24126);
or U26210 (N_26210,N_24473,N_24119);
nand U26211 (N_26211,N_25130,N_24199);
xor U26212 (N_26212,N_25018,N_24252);
nor U26213 (N_26213,N_24208,N_24708);
and U26214 (N_26214,N_24185,N_24460);
or U26215 (N_26215,N_24650,N_24314);
xor U26216 (N_26216,N_24347,N_24353);
or U26217 (N_26217,N_24753,N_24357);
xor U26218 (N_26218,N_24515,N_24534);
nand U26219 (N_26219,N_24287,N_24385);
nor U26220 (N_26220,N_25027,N_24386);
xnor U26221 (N_26221,N_24814,N_24454);
or U26222 (N_26222,N_24060,N_24832);
or U26223 (N_26223,N_24085,N_24422);
nand U26224 (N_26224,N_25166,N_24270);
or U26225 (N_26225,N_24237,N_24737);
nor U26226 (N_26226,N_25071,N_24356);
nand U26227 (N_26227,N_24730,N_24931);
nor U26228 (N_26228,N_24038,N_24150);
nand U26229 (N_26229,N_24571,N_24824);
nand U26230 (N_26230,N_24370,N_24419);
or U26231 (N_26231,N_24838,N_24731);
nand U26232 (N_26232,N_24798,N_24710);
nand U26233 (N_26233,N_24634,N_24902);
nor U26234 (N_26234,N_24025,N_25029);
nor U26235 (N_26235,N_24818,N_24839);
nand U26236 (N_26236,N_24846,N_24319);
nor U26237 (N_26237,N_24475,N_24994);
and U26238 (N_26238,N_24705,N_24127);
nand U26239 (N_26239,N_24525,N_24265);
nor U26240 (N_26240,N_24132,N_24386);
nand U26241 (N_26241,N_24499,N_24906);
or U26242 (N_26242,N_25144,N_24527);
nor U26243 (N_26243,N_24137,N_24890);
nor U26244 (N_26244,N_24452,N_24689);
nand U26245 (N_26245,N_24520,N_25077);
nand U26246 (N_26246,N_24886,N_24414);
nor U26247 (N_26247,N_24673,N_24934);
nand U26248 (N_26248,N_24840,N_24863);
nor U26249 (N_26249,N_24761,N_24264);
nand U26250 (N_26250,N_24374,N_24368);
or U26251 (N_26251,N_24954,N_24845);
and U26252 (N_26252,N_24822,N_24975);
and U26253 (N_26253,N_24504,N_24645);
xor U26254 (N_26254,N_24395,N_24790);
and U26255 (N_26255,N_24848,N_24814);
and U26256 (N_26256,N_25179,N_25018);
and U26257 (N_26257,N_24896,N_25041);
or U26258 (N_26258,N_24846,N_24960);
and U26259 (N_26259,N_24201,N_24668);
xnor U26260 (N_26260,N_24760,N_24435);
and U26261 (N_26261,N_24798,N_24139);
nand U26262 (N_26262,N_24363,N_25159);
nor U26263 (N_26263,N_24816,N_24479);
xor U26264 (N_26264,N_24584,N_24332);
nor U26265 (N_26265,N_24774,N_24441);
nor U26266 (N_26266,N_24825,N_24925);
nor U26267 (N_26267,N_24957,N_24832);
or U26268 (N_26268,N_25119,N_24529);
nor U26269 (N_26269,N_24907,N_24706);
and U26270 (N_26270,N_25026,N_24602);
nor U26271 (N_26271,N_24519,N_24483);
or U26272 (N_26272,N_24311,N_24610);
and U26273 (N_26273,N_24026,N_24115);
nand U26274 (N_26274,N_24245,N_24373);
and U26275 (N_26275,N_24151,N_24806);
nor U26276 (N_26276,N_24930,N_25084);
xor U26277 (N_26277,N_24932,N_24712);
xor U26278 (N_26278,N_25041,N_24246);
or U26279 (N_26279,N_24489,N_24329);
nor U26280 (N_26280,N_24203,N_24419);
or U26281 (N_26281,N_24787,N_24074);
and U26282 (N_26282,N_24576,N_24405);
or U26283 (N_26283,N_24061,N_25042);
nand U26284 (N_26284,N_24550,N_24363);
nor U26285 (N_26285,N_25044,N_25122);
and U26286 (N_26286,N_24245,N_24998);
and U26287 (N_26287,N_24948,N_24224);
nand U26288 (N_26288,N_24573,N_24945);
and U26289 (N_26289,N_24027,N_24557);
nor U26290 (N_26290,N_24916,N_24202);
nand U26291 (N_26291,N_24974,N_24274);
nor U26292 (N_26292,N_24232,N_24280);
or U26293 (N_26293,N_24073,N_24968);
xor U26294 (N_26294,N_24129,N_24731);
and U26295 (N_26295,N_24796,N_25021);
nand U26296 (N_26296,N_25178,N_24734);
or U26297 (N_26297,N_24791,N_24676);
and U26298 (N_26298,N_24063,N_25134);
xor U26299 (N_26299,N_24164,N_24736);
nand U26300 (N_26300,N_24945,N_24769);
and U26301 (N_26301,N_24504,N_24413);
xnor U26302 (N_26302,N_24768,N_24651);
xnor U26303 (N_26303,N_24977,N_24695);
or U26304 (N_26304,N_24970,N_24536);
nand U26305 (N_26305,N_24241,N_24649);
nand U26306 (N_26306,N_24939,N_25035);
nor U26307 (N_26307,N_24526,N_24736);
or U26308 (N_26308,N_24353,N_24151);
nor U26309 (N_26309,N_24289,N_24764);
nand U26310 (N_26310,N_24835,N_24926);
and U26311 (N_26311,N_24396,N_24725);
xor U26312 (N_26312,N_25031,N_24981);
nor U26313 (N_26313,N_24287,N_25129);
nand U26314 (N_26314,N_25076,N_24613);
and U26315 (N_26315,N_24425,N_24239);
nand U26316 (N_26316,N_24354,N_24127);
or U26317 (N_26317,N_24674,N_25013);
and U26318 (N_26318,N_24416,N_24944);
nand U26319 (N_26319,N_24046,N_24360);
xnor U26320 (N_26320,N_24903,N_25036);
xor U26321 (N_26321,N_25026,N_24897);
or U26322 (N_26322,N_24165,N_25180);
or U26323 (N_26323,N_24219,N_24892);
xor U26324 (N_26324,N_24642,N_24873);
nor U26325 (N_26325,N_25126,N_25133);
xor U26326 (N_26326,N_24581,N_24162);
xor U26327 (N_26327,N_24892,N_24227);
or U26328 (N_26328,N_24207,N_24483);
and U26329 (N_26329,N_24642,N_24586);
nor U26330 (N_26330,N_24713,N_24392);
nand U26331 (N_26331,N_25036,N_24118);
nor U26332 (N_26332,N_24334,N_24203);
xnor U26333 (N_26333,N_24327,N_24903);
nor U26334 (N_26334,N_24823,N_25188);
nand U26335 (N_26335,N_24487,N_25131);
nor U26336 (N_26336,N_25130,N_24721);
nand U26337 (N_26337,N_25079,N_25192);
xnor U26338 (N_26338,N_24629,N_25144);
or U26339 (N_26339,N_24764,N_25132);
xnor U26340 (N_26340,N_24505,N_24625);
or U26341 (N_26341,N_24652,N_24474);
or U26342 (N_26342,N_24660,N_24028);
or U26343 (N_26343,N_24259,N_24368);
or U26344 (N_26344,N_24529,N_24437);
xor U26345 (N_26345,N_24810,N_24378);
or U26346 (N_26346,N_24678,N_24758);
xnor U26347 (N_26347,N_24365,N_24728);
and U26348 (N_26348,N_24413,N_24963);
xnor U26349 (N_26349,N_25192,N_24638);
nor U26350 (N_26350,N_24719,N_24438);
and U26351 (N_26351,N_24829,N_24078);
nor U26352 (N_26352,N_24078,N_25113);
nand U26353 (N_26353,N_24501,N_24648);
or U26354 (N_26354,N_24264,N_24512);
and U26355 (N_26355,N_24057,N_24539);
nor U26356 (N_26356,N_25184,N_24671);
xnor U26357 (N_26357,N_25150,N_24318);
nand U26358 (N_26358,N_24498,N_25181);
or U26359 (N_26359,N_24431,N_24929);
nand U26360 (N_26360,N_24675,N_24639);
nand U26361 (N_26361,N_24964,N_24077);
and U26362 (N_26362,N_24710,N_24931);
nor U26363 (N_26363,N_24139,N_24314);
xor U26364 (N_26364,N_24197,N_24383);
nor U26365 (N_26365,N_24691,N_25100);
nor U26366 (N_26366,N_25170,N_24297);
and U26367 (N_26367,N_24494,N_24691);
xnor U26368 (N_26368,N_24847,N_24528);
or U26369 (N_26369,N_25066,N_24568);
or U26370 (N_26370,N_25160,N_24336);
nor U26371 (N_26371,N_24258,N_24752);
xnor U26372 (N_26372,N_24529,N_24884);
nor U26373 (N_26373,N_24266,N_24618);
or U26374 (N_26374,N_25138,N_25039);
nor U26375 (N_26375,N_24099,N_24938);
nand U26376 (N_26376,N_24828,N_25167);
or U26377 (N_26377,N_24689,N_24496);
and U26378 (N_26378,N_24825,N_24387);
xnor U26379 (N_26379,N_24438,N_24270);
and U26380 (N_26380,N_24468,N_24825);
nand U26381 (N_26381,N_24325,N_24461);
xnor U26382 (N_26382,N_24804,N_24567);
nand U26383 (N_26383,N_24009,N_24023);
and U26384 (N_26384,N_24223,N_24380);
nand U26385 (N_26385,N_24852,N_24436);
nor U26386 (N_26386,N_24536,N_24567);
nand U26387 (N_26387,N_24489,N_25030);
nand U26388 (N_26388,N_24528,N_24434);
nor U26389 (N_26389,N_24977,N_24990);
nor U26390 (N_26390,N_24257,N_24854);
or U26391 (N_26391,N_24221,N_24075);
xor U26392 (N_26392,N_24269,N_25039);
nor U26393 (N_26393,N_25177,N_25144);
or U26394 (N_26394,N_24106,N_24302);
nand U26395 (N_26395,N_24161,N_25190);
nor U26396 (N_26396,N_24400,N_24022);
nor U26397 (N_26397,N_24320,N_24819);
or U26398 (N_26398,N_24461,N_24261);
and U26399 (N_26399,N_24051,N_24686);
nand U26400 (N_26400,N_26389,N_25790);
nand U26401 (N_26401,N_25233,N_26095);
and U26402 (N_26402,N_25384,N_25682);
xnor U26403 (N_26403,N_25912,N_26265);
and U26404 (N_26404,N_26032,N_25488);
nand U26405 (N_26405,N_25509,N_26307);
nand U26406 (N_26406,N_25497,N_25681);
nand U26407 (N_26407,N_25683,N_25436);
or U26408 (N_26408,N_26266,N_25717);
nor U26409 (N_26409,N_25966,N_26010);
and U26410 (N_26410,N_25555,N_25578);
and U26411 (N_26411,N_25301,N_25923);
xor U26412 (N_26412,N_25930,N_25324);
nor U26413 (N_26413,N_26379,N_25244);
xor U26414 (N_26414,N_25518,N_25872);
nand U26415 (N_26415,N_25772,N_26334);
and U26416 (N_26416,N_25726,N_26114);
and U26417 (N_26417,N_25937,N_25973);
nor U26418 (N_26418,N_26272,N_25900);
and U26419 (N_26419,N_25315,N_25481);
nor U26420 (N_26420,N_26018,N_25261);
nand U26421 (N_26421,N_26077,N_25745);
xnor U26422 (N_26422,N_25644,N_26262);
xnor U26423 (N_26423,N_26270,N_25722);
or U26424 (N_26424,N_26170,N_26244);
or U26425 (N_26425,N_25758,N_25522);
or U26426 (N_26426,N_25853,N_25380);
or U26427 (N_26427,N_26356,N_26362);
xnor U26428 (N_26428,N_25550,N_25844);
nor U26429 (N_26429,N_26236,N_25378);
nand U26430 (N_26430,N_25415,N_26116);
and U26431 (N_26431,N_26312,N_26344);
or U26432 (N_26432,N_25970,N_25286);
nand U26433 (N_26433,N_26257,N_25934);
nand U26434 (N_26434,N_25417,N_26172);
nor U26435 (N_26435,N_26011,N_25306);
and U26436 (N_26436,N_25926,N_26215);
nor U26437 (N_26437,N_26180,N_25670);
nor U26438 (N_26438,N_25986,N_25775);
nor U26439 (N_26439,N_25251,N_25339);
and U26440 (N_26440,N_25792,N_25441);
nand U26441 (N_26441,N_25875,N_26297);
nor U26442 (N_26442,N_26001,N_25988);
or U26443 (N_26443,N_26377,N_25506);
or U26444 (N_26444,N_25655,N_26275);
or U26445 (N_26445,N_25410,N_26020);
xnor U26446 (N_26446,N_26027,N_25546);
nor U26447 (N_26447,N_25927,N_25692);
xnor U26448 (N_26448,N_26125,N_26237);
xnor U26449 (N_26449,N_25219,N_26056);
and U26450 (N_26450,N_25285,N_25297);
and U26451 (N_26451,N_25250,N_26325);
nor U26452 (N_26452,N_26383,N_25232);
nor U26453 (N_26453,N_25908,N_25987);
and U26454 (N_26454,N_25452,N_26251);
and U26455 (N_26455,N_25494,N_25742);
and U26456 (N_26456,N_25723,N_26289);
and U26457 (N_26457,N_26352,N_26053);
or U26458 (N_26458,N_26252,N_25815);
or U26459 (N_26459,N_25290,N_26296);
xor U26460 (N_26460,N_25230,N_25551);
nor U26461 (N_26461,N_25449,N_26290);
xor U26462 (N_26462,N_25467,N_25400);
nor U26463 (N_26463,N_26256,N_25289);
nand U26464 (N_26464,N_25423,N_25605);
or U26465 (N_26465,N_25253,N_25967);
and U26466 (N_26466,N_25740,N_25470);
nand U26467 (N_26467,N_25820,N_25450);
nor U26468 (N_26468,N_25572,N_25403);
xnor U26469 (N_26469,N_25554,N_25619);
nor U26470 (N_26470,N_26068,N_25733);
nand U26471 (N_26471,N_25870,N_26098);
and U26472 (N_26472,N_25440,N_25404);
xor U26473 (N_26473,N_26036,N_26299);
and U26474 (N_26474,N_25596,N_25992);
and U26475 (N_26475,N_26385,N_26047);
nor U26476 (N_26476,N_26305,N_25453);
nand U26477 (N_26477,N_25932,N_25952);
nand U26478 (N_26478,N_26375,N_26142);
and U26479 (N_26479,N_25531,N_26288);
nor U26480 (N_26480,N_26143,N_25951);
nor U26481 (N_26481,N_25746,N_25767);
or U26482 (N_26482,N_26196,N_25336);
nand U26483 (N_26483,N_25222,N_25834);
nand U26484 (N_26484,N_25255,N_26173);
nor U26485 (N_26485,N_25806,N_26364);
nor U26486 (N_26486,N_25977,N_25995);
nor U26487 (N_26487,N_26137,N_25846);
xnor U26488 (N_26488,N_25848,N_25840);
xor U26489 (N_26489,N_25744,N_26329);
nor U26490 (N_26490,N_25543,N_25203);
or U26491 (N_26491,N_25200,N_26024);
nand U26492 (N_26492,N_25625,N_25676);
and U26493 (N_26493,N_25728,N_25898);
nor U26494 (N_26494,N_25854,N_26348);
or U26495 (N_26495,N_26133,N_25502);
nand U26496 (N_26496,N_25482,N_25549);
or U26497 (N_26497,N_25401,N_25789);
xor U26498 (N_26498,N_25770,N_26023);
and U26499 (N_26499,N_25353,N_25749);
nand U26500 (N_26500,N_25771,N_26003);
nand U26501 (N_26501,N_25458,N_26310);
and U26502 (N_26502,N_25528,N_26057);
nand U26503 (N_26503,N_25617,N_26337);
nor U26504 (N_26504,N_25680,N_26219);
nand U26505 (N_26505,N_25371,N_25348);
xor U26506 (N_26506,N_25547,N_26387);
nand U26507 (N_26507,N_25968,N_25472);
or U26508 (N_26508,N_25313,N_25719);
and U26509 (N_26509,N_25924,N_25354);
or U26510 (N_26510,N_25239,N_26226);
and U26511 (N_26511,N_25471,N_25364);
xnor U26512 (N_26512,N_26086,N_26159);
nor U26513 (N_26513,N_25917,N_26330);
nand U26514 (N_26514,N_25727,N_25469);
and U26515 (N_26515,N_26171,N_25787);
nor U26516 (N_26516,N_25939,N_25704);
nand U26517 (N_26517,N_25838,N_26393);
nor U26518 (N_26518,N_25208,N_25713);
xor U26519 (N_26519,N_25931,N_25238);
nor U26520 (N_26520,N_25609,N_26005);
and U26521 (N_26521,N_26199,N_25212);
xnor U26522 (N_26522,N_25801,N_25517);
nand U26523 (N_26523,N_25539,N_25283);
and U26524 (N_26524,N_25669,N_25365);
nand U26525 (N_26525,N_25984,N_26102);
nor U26526 (N_26526,N_25635,N_25763);
nand U26527 (N_26527,N_26363,N_26082);
nor U26528 (N_26528,N_26368,N_26263);
xnor U26529 (N_26529,N_25529,N_25779);
or U26530 (N_26530,N_25485,N_25651);
and U26531 (N_26531,N_26333,N_26223);
or U26532 (N_26532,N_26146,N_25850);
and U26533 (N_26533,N_26324,N_25499);
nand U26534 (N_26534,N_25573,N_25249);
and U26535 (N_26535,N_26315,N_25795);
or U26536 (N_26536,N_25586,N_25310);
nor U26537 (N_26537,N_25929,N_25272);
xor U26538 (N_26538,N_25426,N_25366);
and U26539 (N_26539,N_26012,N_25533);
xnor U26540 (N_26540,N_25418,N_26370);
or U26541 (N_26541,N_25358,N_26323);
or U26542 (N_26542,N_25442,N_25759);
nor U26543 (N_26543,N_25439,N_25796);
xor U26544 (N_26544,N_25413,N_26260);
and U26545 (N_26545,N_26374,N_25750);
xnor U26546 (N_26546,N_25590,N_25591);
and U26547 (N_26547,N_25580,N_25414);
or U26548 (N_26548,N_25448,N_26188);
nor U26549 (N_26549,N_25925,N_25679);
and U26550 (N_26550,N_25468,N_26386);
and U26551 (N_26551,N_25715,N_25397);
nor U26552 (N_26552,N_25621,N_26074);
nand U26553 (N_26553,N_25457,N_25832);
xor U26554 (N_26554,N_25803,N_25646);
or U26555 (N_26555,N_26293,N_26115);
xor U26556 (N_26556,N_25774,N_25491);
or U26557 (N_26557,N_25693,N_25443);
and U26558 (N_26558,N_26093,N_25785);
nand U26559 (N_26559,N_25647,N_25303);
nand U26560 (N_26560,N_25891,N_25639);
nand U26561 (N_26561,N_25201,N_25691);
xnor U26562 (N_26562,N_26145,N_25548);
xor U26563 (N_26563,N_25629,N_25226);
nand U26564 (N_26564,N_25828,N_26126);
nor U26565 (N_26565,N_25961,N_25780);
or U26566 (N_26566,N_26064,N_25595);
nor U26567 (N_26567,N_26281,N_26050);
or U26568 (N_26568,N_25207,N_25507);
xor U26569 (N_26569,N_26000,N_26309);
and U26570 (N_26570,N_26378,N_25406);
xnor U26571 (N_26571,N_25399,N_25213);
nand U26572 (N_26572,N_25330,N_25957);
nand U26573 (N_26573,N_26351,N_25424);
xor U26574 (N_26574,N_25852,N_25390);
nand U26575 (N_26575,N_25786,N_25698);
and U26576 (N_26576,N_26062,N_25408);
nor U26577 (N_26577,N_25534,N_25508);
and U26578 (N_26578,N_26066,N_26306);
nand U26579 (N_26579,N_26092,N_26382);
xnor U26580 (N_26580,N_25275,N_26398);
or U26581 (N_26581,N_25949,N_26298);
nor U26582 (N_26582,N_26072,N_25429);
or U26583 (N_26583,N_25519,N_26080);
or U26584 (N_26584,N_26157,N_25907);
and U26585 (N_26585,N_26336,N_25363);
nand U26586 (N_26586,N_25849,N_25905);
and U26587 (N_26587,N_25826,N_25668);
xor U26588 (N_26588,N_25876,N_26063);
or U26589 (N_26589,N_25411,N_25524);
nor U26590 (N_26590,N_25976,N_25376);
xnor U26591 (N_26591,N_25794,N_25477);
nor U26592 (N_26592,N_25236,N_25612);
xnor U26593 (N_26593,N_25557,N_25257);
nor U26594 (N_26594,N_26155,N_25540);
nand U26595 (N_26595,N_26224,N_25483);
nand U26596 (N_26596,N_26111,N_25823);
or U26597 (N_26597,N_26217,N_25622);
nand U26598 (N_26598,N_26091,N_25765);
and U26599 (N_26599,N_26112,N_26141);
or U26600 (N_26600,N_25229,N_25950);
nor U26601 (N_26601,N_26350,N_25292);
and U26602 (N_26602,N_26273,N_25730);
and U26603 (N_26603,N_26345,N_25277);
nor U26604 (N_26604,N_26174,N_25456);
and U26605 (N_26605,N_26164,N_25460);
and U26606 (N_26606,N_25327,N_26354);
nand U26607 (N_26607,N_25465,N_26055);
nand U26608 (N_26608,N_25671,N_26235);
or U26609 (N_26609,N_25818,N_25493);
or U26610 (N_26610,N_25274,N_26104);
nand U26611 (N_26611,N_26274,N_25752);
nand U26612 (N_26612,N_25329,N_25293);
or U26613 (N_26613,N_25821,N_25210);
xor U26614 (N_26614,N_25420,N_25603);
or U26615 (N_26615,N_25464,N_25699);
or U26616 (N_26616,N_25802,N_26042);
nand U26617 (N_26617,N_25258,N_25824);
nor U26618 (N_26618,N_25707,N_25858);
xnor U26619 (N_26619,N_26109,N_26085);
xor U26620 (N_26620,N_25690,N_26208);
xnor U26621 (N_26621,N_25817,N_25735);
and U26622 (N_26622,N_26203,N_25663);
nor U26623 (N_26623,N_25247,N_26007);
xor U26624 (N_26624,N_26090,N_25355);
xnor U26625 (N_26625,N_26278,N_25489);
and U26626 (N_26626,N_26014,N_25511);
nor U26627 (N_26627,N_25703,N_25337);
nand U26628 (N_26628,N_25807,N_25545);
or U26629 (N_26629,N_25428,N_25665);
xor U26630 (N_26630,N_25438,N_25294);
xor U26631 (N_26631,N_25281,N_26234);
nor U26632 (N_26632,N_26120,N_25536);
or U26633 (N_26633,N_25566,N_26136);
or U26634 (N_26634,N_26338,N_25357);
nand U26635 (N_26635,N_25971,N_26051);
and U26636 (N_26636,N_26294,N_26328);
and U26637 (N_26637,N_25687,N_25835);
nor U26638 (N_26638,N_25433,N_25847);
or U26639 (N_26639,N_25737,N_25869);
and U26640 (N_26640,N_25656,N_25338);
and U26641 (N_26641,N_25711,N_26373);
or U26642 (N_26642,N_26206,N_26360);
xnor U26643 (N_26643,N_25445,N_25295);
and U26644 (N_26644,N_25955,N_25302);
and U26645 (N_26645,N_25963,N_25736);
and U26646 (N_26646,N_25667,N_26103);
and U26647 (N_26647,N_25326,N_25267);
xor U26648 (N_26648,N_25755,N_25553);
and U26649 (N_26649,N_25328,N_25799);
and U26650 (N_26650,N_26067,N_26240);
nand U26651 (N_26651,N_25761,N_25666);
or U26652 (N_26652,N_25892,N_26204);
xor U26653 (N_26653,N_26279,N_25215);
xor U26654 (N_26654,N_26127,N_26107);
or U26655 (N_26655,N_26213,N_26303);
nand U26656 (N_26656,N_25375,N_25351);
and U26657 (N_26657,N_25263,N_25718);
or U26658 (N_26658,N_25412,N_25659);
nand U26659 (N_26659,N_25855,N_26030);
xor U26660 (N_26660,N_25915,N_25822);
or U26661 (N_26661,N_25476,N_25756);
or U26662 (N_26662,N_25347,N_26031);
nand U26663 (N_26663,N_26140,N_26156);
and U26664 (N_26664,N_25396,N_25367);
nand U26665 (N_26665,N_25920,N_26061);
and U26666 (N_26666,N_26396,N_25863);
or U26667 (N_26667,N_25712,N_25897);
nor U26668 (N_26668,N_25217,N_26269);
nor U26669 (N_26669,N_26069,N_26008);
nor U26670 (N_26670,N_26372,N_26179);
nor U26671 (N_26671,N_26258,N_25562);
and U26672 (N_26672,N_26308,N_25696);
xor U26673 (N_26673,N_25938,N_25321);
nand U26674 (N_26674,N_25246,N_25672);
or U26675 (N_26675,N_26193,N_25317);
and U26676 (N_26676,N_25903,N_25416);
xor U26677 (N_26677,N_25487,N_26096);
and U26678 (N_26678,N_25709,N_25446);
nor U26679 (N_26679,N_26233,N_25322);
nand U26680 (N_26680,N_25579,N_26059);
or U26681 (N_26681,N_25587,N_25810);
nand U26682 (N_26682,N_25252,N_26052);
and U26683 (N_26683,N_25314,N_25993);
and U26684 (N_26684,N_26343,N_25387);
or U26685 (N_26685,N_25648,N_26198);
xor U26686 (N_26686,N_26191,N_25705);
nor U26687 (N_26687,N_25583,N_26158);
nor U26688 (N_26688,N_25325,N_25879);
nand U26689 (N_26689,N_25922,N_26124);
nand U26690 (N_26690,N_26004,N_26232);
nand U26691 (N_26691,N_25998,N_25643);
or U26692 (N_26692,N_25747,N_25444);
and U26693 (N_26693,N_26108,N_25262);
and U26694 (N_26694,N_26227,N_25486);
xnor U26695 (N_26695,N_26197,N_26039);
xor U26696 (N_26696,N_25362,N_26110);
or U26697 (N_26697,N_25377,N_25606);
xor U26698 (N_26698,N_25234,N_25636);
nand U26699 (N_26699,N_26094,N_25373);
xor U26700 (N_26700,N_26181,N_26081);
and U26701 (N_26701,N_25577,N_25532);
xor U26702 (N_26702,N_25899,N_25860);
and U26703 (N_26703,N_25425,N_26161);
or U26704 (N_26704,N_25784,N_26248);
nor U26705 (N_26705,N_26166,N_26033);
nor U26706 (N_26706,N_26218,N_25732);
nor U26707 (N_26707,N_25269,N_25216);
or U26708 (N_26708,N_26002,N_25650);
or U26709 (N_26709,N_25574,N_25983);
and U26710 (N_26710,N_25340,N_25883);
and U26711 (N_26711,N_25298,N_25356);
nor U26712 (N_26712,N_25607,N_25520);
nand U26713 (N_26713,N_25343,N_26332);
nor U26714 (N_26714,N_26169,N_25830);
xor U26715 (N_26715,N_26229,N_26040);
nor U26716 (N_26716,N_26349,N_25389);
or U26717 (N_26717,N_26015,N_26147);
xor U26718 (N_26718,N_26060,N_25500);
xnor U26719 (N_26719,N_25697,N_26316);
and U26720 (N_26720,N_25868,N_25381);
nand U26721 (N_26721,N_26201,N_26205);
xor U26722 (N_26722,N_25896,N_25515);
nand U26723 (N_26723,N_25563,N_25490);
and U26724 (N_26724,N_25827,N_25311);
nand U26725 (N_26725,N_25352,N_26250);
nand U26726 (N_26726,N_26361,N_26228);
or U26727 (N_26727,N_25972,N_26182);
xor U26728 (N_26728,N_25902,N_26300);
xor U26729 (N_26729,N_25565,N_25942);
nor U26730 (N_26730,N_26314,N_26178);
or U26731 (N_26731,N_25833,N_26302);
or U26732 (N_26732,N_25660,N_25268);
or U26733 (N_26733,N_25561,N_25716);
and U26734 (N_26734,N_25243,N_25335);
and U26735 (N_26735,N_26285,N_25836);
nor U26736 (N_26736,N_25649,N_26121);
xnor U26737 (N_26737,N_25652,N_25409);
xnor U26738 (N_26738,N_25632,N_25299);
nor U26739 (N_26739,N_25626,N_26376);
nor U26740 (N_26740,N_25701,N_26190);
nand U26741 (N_26741,N_25594,N_25382);
and U26742 (N_26742,N_26397,N_25913);
nand U26743 (N_26743,N_26335,N_25618);
nor U26744 (N_26744,N_25944,N_25997);
nor U26745 (N_26745,N_25978,N_25537);
or U26746 (N_26746,N_25941,N_25960);
xor U26747 (N_26747,N_25461,N_25323);
or U26748 (N_26748,N_25597,N_26177);
xnor U26749 (N_26749,N_25318,N_25804);
or U26750 (N_26750,N_25623,N_25361);
nand U26751 (N_26751,N_25296,N_25560);
or U26752 (N_26752,N_25615,N_26395);
xnor U26753 (N_26753,N_25598,N_25316);
and U26754 (N_26754,N_26019,N_26186);
nor U26755 (N_26755,N_25421,N_25884);
and U26756 (N_26756,N_25266,N_26192);
nor U26757 (N_26757,N_25739,N_25223);
nor U26758 (N_26758,N_26113,N_26148);
or U26759 (N_26759,N_25714,N_25874);
xor U26760 (N_26760,N_26117,N_25245);
and U26761 (N_26761,N_25738,N_25631);
nand U26762 (N_26762,N_25769,N_26207);
and U26763 (N_26763,N_25345,N_25569);
nand U26764 (N_26764,N_26097,N_25702);
or U26765 (N_26765,N_26313,N_25270);
nor U26766 (N_26766,N_26341,N_25783);
or U26767 (N_26767,N_26139,N_26399);
nor U26768 (N_26768,N_25990,N_25276);
and U26769 (N_26769,N_25599,N_25225);
or U26770 (N_26770,N_25819,N_25312);
nand U26771 (N_26771,N_25886,N_26183);
nor U26772 (N_26772,N_25535,N_25305);
nand U26773 (N_26773,N_26026,N_26021);
or U26774 (N_26774,N_25825,N_25965);
xnor U26775 (N_26775,N_25220,N_25684);
and U26776 (N_26776,N_25678,N_25558);
or U26777 (N_26777,N_26211,N_25265);
xor U26778 (N_26778,N_26046,N_25432);
nand U26779 (N_26779,N_26283,N_25206);
and U26780 (N_26780,N_25334,N_26163);
or U26781 (N_26781,N_25956,N_26175);
nand U26782 (N_26782,N_25492,N_26189);
nand U26783 (N_26783,N_25564,N_25495);
nor U26784 (N_26784,N_25708,N_26245);
nand U26785 (N_26785,N_25567,N_25205);
and U26786 (N_26786,N_25946,N_25989);
xnor U26787 (N_26787,N_26070,N_25478);
or U26788 (N_26788,N_26073,N_25673);
and U26789 (N_26789,N_26322,N_25556);
xnor U26790 (N_26790,N_25422,N_25505);
nor U26791 (N_26791,N_26267,N_26243);
nor U26792 (N_26792,N_25766,N_26134);
xor U26793 (N_26793,N_25451,N_25627);
and U26794 (N_26794,N_25405,N_26388);
nand U26795 (N_26795,N_25630,N_25264);
nand U26796 (N_26796,N_25278,N_25542);
nor U26797 (N_26797,N_26119,N_25857);
or U26798 (N_26798,N_25809,N_26165);
or U26799 (N_26799,N_25308,N_25805);
or U26800 (N_26800,N_25781,N_25510);
and U26801 (N_26801,N_25331,N_26167);
nor U26802 (N_26802,N_25991,N_25273);
nor U26803 (N_26803,N_25641,N_25657);
nor U26804 (N_26804,N_25773,N_26261);
xnor U26805 (N_26805,N_25231,N_25589);
and U26806 (N_26806,N_25282,N_25909);
xor U26807 (N_26807,N_25571,N_25741);
nand U26808 (N_26808,N_25751,N_25757);
nor U26809 (N_26809,N_25936,N_25209);
or U26810 (N_26810,N_25889,N_26038);
or U26811 (N_26811,N_26331,N_25582);
nand U26812 (N_26812,N_25611,N_26105);
nand U26813 (N_26813,N_25608,N_25935);
and U26814 (N_26814,N_25501,N_26230);
and U26815 (N_26815,N_26168,N_25918);
and U26816 (N_26816,N_26392,N_25873);
xnor U26817 (N_26817,N_26017,N_26129);
and U26818 (N_26818,N_26152,N_25241);
xor U26819 (N_26819,N_26216,N_25812);
xor U26820 (N_26820,N_26369,N_25394);
and U26821 (N_26821,N_25890,N_25981);
or U26822 (N_26822,N_26122,N_25504);
nand U26823 (N_26823,N_26123,N_25584);
nand U26824 (N_26824,N_25845,N_25513);
xnor U26825 (N_26825,N_26212,N_26225);
and U26826 (N_26826,N_25237,N_26282);
nand U26827 (N_26827,N_25385,N_25947);
and U26828 (N_26828,N_26150,N_26048);
xnor U26829 (N_26829,N_26284,N_26058);
or U26830 (N_26830,N_25975,N_26100);
nand U26831 (N_26831,N_25593,N_26380);
nor U26832 (N_26832,N_26037,N_25914);
xor U26833 (N_26833,N_25882,N_25674);
nand U26834 (N_26834,N_25284,N_25797);
and U26835 (N_26835,N_25710,N_26043);
and U26836 (N_26836,N_25475,N_25782);
xor U26837 (N_26837,N_25911,N_26153);
nand U26838 (N_26838,N_26162,N_25211);
and U26839 (N_26839,N_25653,N_25862);
nor U26840 (N_26840,N_25894,N_25342);
nor U26841 (N_26841,N_25228,N_25948);
and U26842 (N_26842,N_25633,N_25700);
and U26843 (N_26843,N_26118,N_25473);
xor U26844 (N_26844,N_25592,N_25530);
and U26845 (N_26845,N_25859,N_26287);
nor U26846 (N_26846,N_26187,N_25600);
nand U26847 (N_26847,N_25304,N_25431);
and U26848 (N_26848,N_25344,N_25260);
nand U26849 (N_26849,N_25793,N_25346);
and U26850 (N_26850,N_25829,N_25919);
xnor U26851 (N_26851,N_25658,N_25843);
xnor U26852 (N_26852,N_25570,N_25514);
nor U26853 (N_26853,N_25388,N_25224);
or U26854 (N_26854,N_25398,N_25333);
and U26855 (N_26855,N_26365,N_25434);
xor U26856 (N_26856,N_25259,N_25867);
xor U26857 (N_26857,N_25474,N_25837);
xor U26858 (N_26858,N_26160,N_26202);
nand U26859 (N_26859,N_25959,N_25402);
or U26860 (N_26860,N_25279,N_25865);
nand U26861 (N_26861,N_26304,N_25974);
and U26862 (N_26862,N_25242,N_25954);
xnor U26863 (N_26863,N_25620,N_25816);
xnor U26864 (N_26864,N_26280,N_25721);
xnor U26865 (N_26865,N_25720,N_26099);
xnor U26866 (N_26866,N_26200,N_25762);
nor U26867 (N_26867,N_26209,N_26013);
nor U26868 (N_26868,N_25760,N_26045);
nor U26869 (N_26869,N_25994,N_25880);
xnor U26870 (N_26870,N_25526,N_26366);
nor U26871 (N_26871,N_25628,N_25601);
xnor U26872 (N_26872,N_26106,N_25221);
nor U26873 (N_26873,N_26271,N_25729);
nor U26874 (N_26874,N_25895,N_25568);
nor U26875 (N_26875,N_26347,N_25734);
or U26876 (N_26876,N_26054,N_26089);
and U26877 (N_26877,N_25359,N_25419);
and U26878 (N_26878,N_26346,N_25204);
nand U26879 (N_26879,N_26384,N_26176);
nand U26880 (N_26880,N_26231,N_25407);
xor U26881 (N_26881,N_25945,N_25675);
xor U26882 (N_26882,N_25814,N_25662);
or U26883 (N_26883,N_25979,N_26041);
and U26884 (N_26884,N_26311,N_26101);
or U26885 (N_26885,N_25982,N_25753);
or U26886 (N_26886,N_25309,N_26044);
or U26887 (N_26887,N_25462,N_26138);
and U26888 (N_26888,N_26238,N_26154);
xnor U26889 (N_26889,N_25706,N_25393);
or U26890 (N_26890,N_26255,N_26131);
and U26891 (N_26891,N_26326,N_25904);
nor U26892 (N_26892,N_25498,N_25523);
and U26893 (N_26893,N_25369,N_25602);
nand U26894 (N_26894,N_25969,N_25372);
and U26895 (N_26895,N_26321,N_25370);
nand U26896 (N_26896,N_26355,N_25839);
or U26897 (N_26897,N_25808,N_26149);
and U26898 (N_26898,N_26242,N_25831);
or U26899 (N_26899,N_25427,N_26253);
or U26900 (N_26900,N_26214,N_26151);
or U26901 (N_26901,N_26381,N_26016);
or U26902 (N_26902,N_25463,N_25300);
and U26903 (N_26903,N_25613,N_26390);
xor U26904 (N_26904,N_25996,N_25480);
nor U26905 (N_26905,N_25768,N_26239);
and U26906 (N_26906,N_26185,N_25861);
nand U26907 (N_26907,N_25642,N_26035);
xnor U26908 (N_26908,N_25287,N_26087);
or U26909 (N_26909,N_25240,N_25368);
nor U26910 (N_26910,N_25616,N_26049);
xor U26911 (N_26911,N_26084,N_25466);
or U26912 (N_26912,N_25392,N_25731);
and U26913 (N_26913,N_25575,N_25754);
or U26914 (N_26914,N_26078,N_26320);
nand U26915 (N_26915,N_25777,N_25503);
nor U26916 (N_26916,N_25640,N_26249);
or U26917 (N_26917,N_26286,N_25588);
xor U26918 (N_26918,N_26259,N_25455);
and U26919 (N_26919,N_25685,N_25319);
and U26920 (N_26920,N_25881,N_25856);
and U26921 (N_26921,N_25689,N_25544);
nand U26922 (N_26922,N_26342,N_26071);
nand U26923 (N_26923,N_25256,N_25637);
and U26924 (N_26924,N_25447,N_26195);
xor U26925 (N_26925,N_25764,N_25686);
or U26926 (N_26926,N_26222,N_26319);
xnor U26927 (N_26927,N_25778,N_25906);
xnor U26928 (N_26928,N_25999,N_26277);
xnor U26929 (N_26929,N_25379,N_25349);
nand U26930 (N_26930,N_26028,N_25430);
nor U26931 (N_26931,N_25341,N_25943);
or U26932 (N_26932,N_25933,N_26065);
nor U26933 (N_26933,N_26327,N_26339);
xor U26934 (N_26934,N_25928,N_25921);
or U26935 (N_26935,N_25218,N_25435);
and U26936 (N_26936,N_25958,N_26268);
or U26937 (N_26937,N_26220,N_26276);
nor U26938 (N_26938,N_25604,N_25516);
nand U26939 (N_26939,N_26254,N_26353);
nand U26940 (N_26940,N_26247,N_25661);
xor U26941 (N_26941,N_25841,N_26083);
nand U26942 (N_26942,N_25743,N_26006);
or U26943 (N_26943,N_26135,N_26359);
nor U26944 (N_26944,N_25512,N_25985);
xor U26945 (N_26945,N_26367,N_25541);
nand U26946 (N_26946,N_26076,N_25454);
and U26947 (N_26947,N_26128,N_25866);
nand U26948 (N_26948,N_25227,N_25776);
and U26949 (N_26949,N_26301,N_25964);
and U26950 (N_26950,N_25552,N_25374);
nand U26951 (N_26951,N_25395,N_25581);
nand U26952 (N_26952,N_25271,N_25695);
xnor U26953 (N_26953,N_25638,N_25496);
nand U26954 (N_26954,N_25887,N_26194);
and U26955 (N_26955,N_25901,N_25910);
nand U26956 (N_26956,N_25788,N_25813);
and U26957 (N_26957,N_26318,N_26184);
and U26958 (N_26958,N_25654,N_25871);
nand U26959 (N_26959,N_25610,N_26130);
or U26960 (N_26960,N_25320,N_26371);
and U26961 (N_26961,N_25800,N_25851);
and U26962 (N_26962,N_25888,N_26291);
nand U26963 (N_26963,N_26025,N_25980);
or U26964 (N_26964,N_25893,N_26075);
xnor U26965 (N_26965,N_25798,N_26144);
or U26966 (N_26966,N_25962,N_26079);
nor U26967 (N_26967,N_26088,N_25688);
xnor U26968 (N_26968,N_25748,N_26391);
nand U26969 (N_26969,N_25645,N_25811);
xor U26970 (N_26970,N_26034,N_25291);
and U26971 (N_26971,N_25842,N_25360);
nor U26972 (N_26972,N_25878,N_26241);
and U26973 (N_26973,N_25288,N_25307);
and U26974 (N_26974,N_26295,N_25538);
xor U26975 (N_26975,N_26132,N_26264);
and U26976 (N_26976,N_25280,N_26009);
xor U26977 (N_26977,N_25940,N_26210);
xor U26978 (N_26978,N_25332,N_26029);
nand U26979 (N_26979,N_25391,N_25791);
nor U26980 (N_26980,N_25885,N_26357);
nor U26981 (N_26981,N_26340,N_25877);
xor U26982 (N_26982,N_25521,N_25953);
or U26983 (N_26983,N_25437,N_25725);
or U26984 (N_26984,N_25576,N_25664);
xnor U26985 (N_26985,N_26394,N_25254);
nor U26986 (N_26986,N_25235,N_25916);
xnor U26987 (N_26987,N_25479,N_25214);
xor U26988 (N_26988,N_26292,N_26022);
xnor U26989 (N_26989,N_25484,N_25525);
xnor U26990 (N_26990,N_26317,N_25585);
xor U26991 (N_26991,N_25634,N_25624);
nor U26992 (N_26992,N_25350,N_26221);
xor U26993 (N_26993,N_25694,N_25614);
nor U26994 (N_26994,N_25864,N_25559);
xor U26995 (N_26995,N_25248,N_25386);
and U26996 (N_26996,N_25724,N_25383);
or U26997 (N_26997,N_25527,N_26246);
and U26998 (N_26998,N_26358,N_25677);
xnor U26999 (N_26999,N_25202,N_25459);
nand U27000 (N_27000,N_25351,N_26087);
nand U27001 (N_27001,N_25448,N_25648);
or U27002 (N_27002,N_26349,N_26392);
or U27003 (N_27003,N_26264,N_25433);
nor U27004 (N_27004,N_25565,N_25307);
and U27005 (N_27005,N_25663,N_25743);
nor U27006 (N_27006,N_26250,N_25861);
xnor U27007 (N_27007,N_26117,N_26360);
nand U27008 (N_27008,N_25617,N_25593);
and U27009 (N_27009,N_25741,N_25409);
nand U27010 (N_27010,N_25566,N_26286);
or U27011 (N_27011,N_26186,N_25699);
or U27012 (N_27012,N_25663,N_25925);
and U27013 (N_27013,N_25249,N_26273);
nor U27014 (N_27014,N_26222,N_25475);
nand U27015 (N_27015,N_25465,N_25436);
or U27016 (N_27016,N_25501,N_25228);
xor U27017 (N_27017,N_25399,N_25652);
nor U27018 (N_27018,N_26395,N_25555);
xnor U27019 (N_27019,N_25525,N_25219);
or U27020 (N_27020,N_25732,N_25831);
xor U27021 (N_27021,N_25748,N_25391);
xor U27022 (N_27022,N_25767,N_25706);
nor U27023 (N_27023,N_25387,N_25495);
or U27024 (N_27024,N_25431,N_26204);
or U27025 (N_27025,N_26179,N_26007);
nor U27026 (N_27026,N_26244,N_25511);
nand U27027 (N_27027,N_25293,N_25767);
nand U27028 (N_27028,N_25973,N_25323);
xor U27029 (N_27029,N_25624,N_25436);
xor U27030 (N_27030,N_26099,N_26175);
nand U27031 (N_27031,N_25703,N_25345);
nand U27032 (N_27032,N_25636,N_25645);
xnor U27033 (N_27033,N_26371,N_26302);
nor U27034 (N_27034,N_25333,N_25990);
nor U27035 (N_27035,N_26099,N_26095);
nand U27036 (N_27036,N_25445,N_26354);
xor U27037 (N_27037,N_26257,N_25846);
nand U27038 (N_27038,N_25503,N_25360);
and U27039 (N_27039,N_26096,N_26177);
nand U27040 (N_27040,N_25398,N_25381);
and U27041 (N_27041,N_25997,N_26100);
nor U27042 (N_27042,N_26380,N_26221);
nor U27043 (N_27043,N_25711,N_25820);
nand U27044 (N_27044,N_25923,N_26367);
xnor U27045 (N_27045,N_26112,N_25300);
xor U27046 (N_27046,N_25740,N_25902);
xor U27047 (N_27047,N_26377,N_25815);
nand U27048 (N_27048,N_25306,N_26250);
and U27049 (N_27049,N_25297,N_25548);
and U27050 (N_27050,N_25974,N_25795);
nor U27051 (N_27051,N_26048,N_25659);
nor U27052 (N_27052,N_25392,N_25719);
or U27053 (N_27053,N_25216,N_25264);
xnor U27054 (N_27054,N_25861,N_25534);
and U27055 (N_27055,N_25641,N_25538);
and U27056 (N_27056,N_25776,N_26175);
nand U27057 (N_27057,N_26153,N_25711);
nor U27058 (N_27058,N_25401,N_26383);
xnor U27059 (N_27059,N_25790,N_26371);
nand U27060 (N_27060,N_25975,N_25858);
or U27061 (N_27061,N_25672,N_26282);
nor U27062 (N_27062,N_25599,N_26384);
and U27063 (N_27063,N_25522,N_25397);
nor U27064 (N_27064,N_25332,N_25743);
or U27065 (N_27065,N_25955,N_25791);
or U27066 (N_27066,N_26377,N_25493);
xor U27067 (N_27067,N_25439,N_25827);
or U27068 (N_27068,N_25768,N_25452);
or U27069 (N_27069,N_25474,N_26094);
xnor U27070 (N_27070,N_25851,N_25252);
nand U27071 (N_27071,N_26191,N_26377);
and U27072 (N_27072,N_26020,N_25631);
or U27073 (N_27073,N_25278,N_25597);
nand U27074 (N_27074,N_26147,N_25506);
nor U27075 (N_27075,N_25429,N_25241);
and U27076 (N_27076,N_25763,N_25654);
and U27077 (N_27077,N_25704,N_26184);
xor U27078 (N_27078,N_25948,N_25309);
xor U27079 (N_27079,N_25201,N_26301);
and U27080 (N_27080,N_26268,N_25626);
nor U27081 (N_27081,N_25979,N_25363);
xor U27082 (N_27082,N_25630,N_25288);
nor U27083 (N_27083,N_25377,N_25295);
xnor U27084 (N_27084,N_25240,N_26278);
nor U27085 (N_27085,N_26106,N_26092);
xor U27086 (N_27086,N_26261,N_26169);
nor U27087 (N_27087,N_25792,N_25296);
or U27088 (N_27088,N_25842,N_25815);
nand U27089 (N_27089,N_25910,N_25936);
and U27090 (N_27090,N_25979,N_26036);
nand U27091 (N_27091,N_26307,N_26217);
nor U27092 (N_27092,N_25341,N_25958);
xnor U27093 (N_27093,N_25524,N_26376);
xor U27094 (N_27094,N_25208,N_25587);
nor U27095 (N_27095,N_26096,N_25422);
and U27096 (N_27096,N_25371,N_26100);
or U27097 (N_27097,N_25567,N_25361);
nor U27098 (N_27098,N_25615,N_25656);
or U27099 (N_27099,N_25716,N_26190);
and U27100 (N_27100,N_25818,N_25774);
or U27101 (N_27101,N_25922,N_25755);
nor U27102 (N_27102,N_25727,N_25716);
nor U27103 (N_27103,N_25802,N_25897);
or U27104 (N_27104,N_26221,N_25643);
nor U27105 (N_27105,N_25377,N_26120);
or U27106 (N_27106,N_25656,N_25624);
nand U27107 (N_27107,N_26150,N_26140);
or U27108 (N_27108,N_25258,N_25710);
xnor U27109 (N_27109,N_25845,N_25887);
or U27110 (N_27110,N_25778,N_25400);
nand U27111 (N_27111,N_26214,N_26096);
xnor U27112 (N_27112,N_25569,N_25977);
or U27113 (N_27113,N_25958,N_26126);
nor U27114 (N_27114,N_26043,N_25553);
or U27115 (N_27115,N_26364,N_26120);
nand U27116 (N_27116,N_25385,N_26329);
or U27117 (N_27117,N_25494,N_25783);
xor U27118 (N_27118,N_26278,N_26298);
and U27119 (N_27119,N_25610,N_25461);
nand U27120 (N_27120,N_26260,N_25200);
or U27121 (N_27121,N_26310,N_25782);
xor U27122 (N_27122,N_26026,N_25795);
nand U27123 (N_27123,N_26333,N_25225);
nor U27124 (N_27124,N_25507,N_26202);
or U27125 (N_27125,N_26063,N_25480);
nand U27126 (N_27126,N_26014,N_25663);
nor U27127 (N_27127,N_25494,N_25364);
and U27128 (N_27128,N_25608,N_26018);
xnor U27129 (N_27129,N_26027,N_25395);
xnor U27130 (N_27130,N_26014,N_25964);
nand U27131 (N_27131,N_25273,N_25541);
and U27132 (N_27132,N_26107,N_25974);
or U27133 (N_27133,N_25609,N_25860);
xor U27134 (N_27134,N_25470,N_25973);
or U27135 (N_27135,N_26336,N_25639);
or U27136 (N_27136,N_26130,N_26069);
and U27137 (N_27137,N_25484,N_25502);
xor U27138 (N_27138,N_25655,N_25246);
and U27139 (N_27139,N_25710,N_25384);
nand U27140 (N_27140,N_25291,N_25433);
or U27141 (N_27141,N_25343,N_25616);
and U27142 (N_27142,N_26342,N_26001);
xnor U27143 (N_27143,N_25697,N_25921);
nor U27144 (N_27144,N_25690,N_25801);
or U27145 (N_27145,N_25855,N_26200);
and U27146 (N_27146,N_26388,N_25601);
xnor U27147 (N_27147,N_25255,N_25841);
and U27148 (N_27148,N_26313,N_26375);
or U27149 (N_27149,N_25438,N_25300);
nand U27150 (N_27150,N_26397,N_25327);
nor U27151 (N_27151,N_26207,N_25525);
or U27152 (N_27152,N_25837,N_25514);
nand U27153 (N_27153,N_25917,N_26270);
nor U27154 (N_27154,N_25782,N_25293);
xor U27155 (N_27155,N_25573,N_25387);
xor U27156 (N_27156,N_25946,N_26154);
nand U27157 (N_27157,N_26049,N_25591);
or U27158 (N_27158,N_26199,N_25792);
nand U27159 (N_27159,N_25580,N_26093);
nor U27160 (N_27160,N_25454,N_25865);
or U27161 (N_27161,N_25663,N_26234);
nand U27162 (N_27162,N_25762,N_26308);
xnor U27163 (N_27163,N_26073,N_26055);
nor U27164 (N_27164,N_25974,N_25727);
xnor U27165 (N_27165,N_26166,N_26041);
nor U27166 (N_27166,N_25592,N_26113);
nand U27167 (N_27167,N_25675,N_26363);
nor U27168 (N_27168,N_25885,N_25835);
nor U27169 (N_27169,N_25648,N_26171);
or U27170 (N_27170,N_25216,N_26043);
nor U27171 (N_27171,N_25616,N_26173);
nor U27172 (N_27172,N_26371,N_26200);
or U27173 (N_27173,N_25942,N_25863);
and U27174 (N_27174,N_26239,N_25367);
and U27175 (N_27175,N_26127,N_25987);
or U27176 (N_27176,N_25376,N_25517);
and U27177 (N_27177,N_25982,N_26313);
and U27178 (N_27178,N_26065,N_26027);
and U27179 (N_27179,N_26044,N_25265);
nand U27180 (N_27180,N_25304,N_25903);
nand U27181 (N_27181,N_25629,N_26328);
xnor U27182 (N_27182,N_26053,N_26010);
nand U27183 (N_27183,N_26209,N_25522);
xor U27184 (N_27184,N_26087,N_25920);
or U27185 (N_27185,N_25809,N_25857);
nor U27186 (N_27186,N_26278,N_25277);
or U27187 (N_27187,N_25726,N_25855);
or U27188 (N_27188,N_25297,N_26206);
or U27189 (N_27189,N_25465,N_25613);
nand U27190 (N_27190,N_26033,N_25957);
xnor U27191 (N_27191,N_25287,N_25306);
nor U27192 (N_27192,N_25213,N_26019);
nor U27193 (N_27193,N_26167,N_25989);
and U27194 (N_27194,N_26187,N_25920);
xnor U27195 (N_27195,N_26088,N_25700);
xor U27196 (N_27196,N_25686,N_25291);
nor U27197 (N_27197,N_26184,N_25537);
and U27198 (N_27198,N_25942,N_26288);
and U27199 (N_27199,N_25670,N_25203);
and U27200 (N_27200,N_25482,N_25664);
and U27201 (N_27201,N_25784,N_26053);
nand U27202 (N_27202,N_26086,N_26243);
nor U27203 (N_27203,N_25858,N_25351);
xor U27204 (N_27204,N_25853,N_25216);
nand U27205 (N_27205,N_25293,N_25559);
or U27206 (N_27206,N_26108,N_26083);
nand U27207 (N_27207,N_26131,N_25567);
nor U27208 (N_27208,N_26166,N_26141);
nor U27209 (N_27209,N_25499,N_25999);
nand U27210 (N_27210,N_25242,N_26276);
nand U27211 (N_27211,N_25496,N_26059);
xnor U27212 (N_27212,N_26237,N_26002);
nand U27213 (N_27213,N_26131,N_25867);
nand U27214 (N_27214,N_25383,N_25336);
nand U27215 (N_27215,N_26278,N_25391);
and U27216 (N_27216,N_25376,N_25234);
and U27217 (N_27217,N_25721,N_25448);
nand U27218 (N_27218,N_25669,N_25881);
or U27219 (N_27219,N_26288,N_25288);
or U27220 (N_27220,N_26247,N_25639);
and U27221 (N_27221,N_26390,N_26049);
or U27222 (N_27222,N_26180,N_25646);
or U27223 (N_27223,N_25369,N_26259);
nor U27224 (N_27224,N_25447,N_25669);
nor U27225 (N_27225,N_26122,N_25450);
nor U27226 (N_27226,N_25677,N_25430);
nor U27227 (N_27227,N_25466,N_25667);
nor U27228 (N_27228,N_25607,N_26045);
nor U27229 (N_27229,N_25939,N_25934);
nand U27230 (N_27230,N_25997,N_25423);
and U27231 (N_27231,N_26398,N_26380);
nor U27232 (N_27232,N_25852,N_25572);
or U27233 (N_27233,N_25861,N_25553);
and U27234 (N_27234,N_26233,N_25879);
nor U27235 (N_27235,N_25551,N_25343);
or U27236 (N_27236,N_25589,N_25319);
nand U27237 (N_27237,N_26103,N_25859);
and U27238 (N_27238,N_26323,N_25568);
and U27239 (N_27239,N_25844,N_26210);
or U27240 (N_27240,N_26336,N_25483);
nor U27241 (N_27241,N_25256,N_26094);
nor U27242 (N_27242,N_25220,N_25638);
nand U27243 (N_27243,N_25962,N_25818);
xnor U27244 (N_27244,N_25345,N_25437);
or U27245 (N_27245,N_25569,N_26060);
or U27246 (N_27246,N_25444,N_25352);
or U27247 (N_27247,N_25439,N_25732);
or U27248 (N_27248,N_26063,N_25246);
nand U27249 (N_27249,N_25925,N_26242);
xnor U27250 (N_27250,N_26361,N_25401);
and U27251 (N_27251,N_25212,N_26210);
or U27252 (N_27252,N_25273,N_26323);
or U27253 (N_27253,N_25640,N_25759);
or U27254 (N_27254,N_26311,N_25573);
or U27255 (N_27255,N_25898,N_25874);
xnor U27256 (N_27256,N_25847,N_25878);
or U27257 (N_27257,N_26375,N_26321);
nand U27258 (N_27258,N_26070,N_25281);
xnor U27259 (N_27259,N_25782,N_25319);
and U27260 (N_27260,N_26091,N_25798);
or U27261 (N_27261,N_25481,N_25283);
or U27262 (N_27262,N_25203,N_25490);
nand U27263 (N_27263,N_25566,N_26047);
nand U27264 (N_27264,N_26008,N_25654);
or U27265 (N_27265,N_25817,N_25217);
nor U27266 (N_27266,N_25516,N_26215);
or U27267 (N_27267,N_25645,N_25728);
and U27268 (N_27268,N_25316,N_26157);
or U27269 (N_27269,N_26068,N_25903);
xor U27270 (N_27270,N_25461,N_25878);
xnor U27271 (N_27271,N_25917,N_26092);
nand U27272 (N_27272,N_25744,N_25353);
xor U27273 (N_27273,N_25987,N_26337);
nand U27274 (N_27274,N_25376,N_26144);
and U27275 (N_27275,N_26179,N_26339);
xnor U27276 (N_27276,N_25746,N_26294);
nand U27277 (N_27277,N_26192,N_26240);
and U27278 (N_27278,N_25418,N_25413);
and U27279 (N_27279,N_25474,N_25946);
and U27280 (N_27280,N_25346,N_25662);
nand U27281 (N_27281,N_25205,N_25617);
xor U27282 (N_27282,N_25870,N_25790);
xnor U27283 (N_27283,N_26017,N_25461);
xor U27284 (N_27284,N_25699,N_26030);
and U27285 (N_27285,N_25943,N_25874);
nor U27286 (N_27286,N_25252,N_25605);
nand U27287 (N_27287,N_25707,N_25840);
xnor U27288 (N_27288,N_26237,N_25627);
or U27289 (N_27289,N_26274,N_25979);
or U27290 (N_27290,N_25308,N_25728);
and U27291 (N_27291,N_25265,N_26332);
xor U27292 (N_27292,N_26071,N_25571);
or U27293 (N_27293,N_26357,N_25442);
nor U27294 (N_27294,N_25578,N_26021);
nor U27295 (N_27295,N_25222,N_25637);
nor U27296 (N_27296,N_25515,N_26225);
xor U27297 (N_27297,N_26358,N_25758);
and U27298 (N_27298,N_26143,N_25324);
nand U27299 (N_27299,N_25872,N_25609);
and U27300 (N_27300,N_25658,N_25702);
nand U27301 (N_27301,N_26067,N_25948);
xnor U27302 (N_27302,N_25376,N_26167);
or U27303 (N_27303,N_26169,N_26224);
or U27304 (N_27304,N_25486,N_25293);
and U27305 (N_27305,N_25276,N_26215);
nor U27306 (N_27306,N_25584,N_26005);
nand U27307 (N_27307,N_26182,N_25515);
nand U27308 (N_27308,N_26246,N_25395);
and U27309 (N_27309,N_26269,N_25419);
xnor U27310 (N_27310,N_25893,N_26017);
nor U27311 (N_27311,N_25503,N_25651);
nand U27312 (N_27312,N_25703,N_25970);
nand U27313 (N_27313,N_25369,N_25490);
xnor U27314 (N_27314,N_25621,N_25829);
or U27315 (N_27315,N_25391,N_25908);
and U27316 (N_27316,N_25333,N_25929);
xnor U27317 (N_27317,N_25950,N_26200);
nor U27318 (N_27318,N_25825,N_25785);
nor U27319 (N_27319,N_25744,N_25952);
or U27320 (N_27320,N_26237,N_25436);
nor U27321 (N_27321,N_25595,N_25877);
nand U27322 (N_27322,N_26102,N_26034);
or U27323 (N_27323,N_26078,N_26394);
and U27324 (N_27324,N_25410,N_25637);
nand U27325 (N_27325,N_25530,N_25454);
nand U27326 (N_27326,N_26032,N_25997);
xnor U27327 (N_27327,N_25960,N_26254);
nor U27328 (N_27328,N_25771,N_26081);
nor U27329 (N_27329,N_25291,N_25493);
xor U27330 (N_27330,N_25838,N_26243);
or U27331 (N_27331,N_25529,N_25673);
xor U27332 (N_27332,N_25457,N_26314);
or U27333 (N_27333,N_25781,N_25708);
or U27334 (N_27334,N_25450,N_25525);
and U27335 (N_27335,N_25463,N_26171);
or U27336 (N_27336,N_25383,N_25257);
nor U27337 (N_27337,N_25989,N_25926);
xnor U27338 (N_27338,N_25236,N_26393);
nand U27339 (N_27339,N_25773,N_25592);
and U27340 (N_27340,N_26391,N_25369);
and U27341 (N_27341,N_25338,N_25974);
or U27342 (N_27342,N_26144,N_25474);
nor U27343 (N_27343,N_26221,N_25894);
nand U27344 (N_27344,N_26150,N_25528);
xor U27345 (N_27345,N_25676,N_25357);
or U27346 (N_27346,N_25881,N_25432);
nand U27347 (N_27347,N_26239,N_25457);
nor U27348 (N_27348,N_25874,N_25276);
and U27349 (N_27349,N_26163,N_25541);
xor U27350 (N_27350,N_26035,N_25372);
nand U27351 (N_27351,N_25609,N_26084);
and U27352 (N_27352,N_25516,N_25469);
or U27353 (N_27353,N_26265,N_25955);
and U27354 (N_27354,N_25281,N_26313);
or U27355 (N_27355,N_25859,N_25784);
nand U27356 (N_27356,N_26142,N_25853);
nand U27357 (N_27357,N_26267,N_25547);
nand U27358 (N_27358,N_25972,N_26135);
and U27359 (N_27359,N_25378,N_25344);
nor U27360 (N_27360,N_25960,N_25482);
nand U27361 (N_27361,N_25933,N_25522);
nand U27362 (N_27362,N_26294,N_25635);
and U27363 (N_27363,N_26307,N_25789);
nand U27364 (N_27364,N_26039,N_26006);
and U27365 (N_27365,N_25667,N_25869);
nor U27366 (N_27366,N_25881,N_26101);
nor U27367 (N_27367,N_25653,N_25272);
nor U27368 (N_27368,N_26225,N_26372);
or U27369 (N_27369,N_25399,N_26320);
and U27370 (N_27370,N_26194,N_26171);
nand U27371 (N_27371,N_25437,N_25294);
or U27372 (N_27372,N_25465,N_25552);
or U27373 (N_27373,N_25502,N_25799);
xnor U27374 (N_27374,N_25238,N_25880);
nor U27375 (N_27375,N_25955,N_26230);
or U27376 (N_27376,N_25549,N_26240);
and U27377 (N_27377,N_25657,N_25447);
nor U27378 (N_27378,N_25889,N_25983);
nor U27379 (N_27379,N_26372,N_25629);
and U27380 (N_27380,N_25996,N_25219);
nand U27381 (N_27381,N_26333,N_25437);
nor U27382 (N_27382,N_25371,N_25986);
nor U27383 (N_27383,N_25726,N_25792);
nand U27384 (N_27384,N_26216,N_25596);
nor U27385 (N_27385,N_25548,N_25486);
nor U27386 (N_27386,N_25361,N_25286);
xor U27387 (N_27387,N_25259,N_26216);
xnor U27388 (N_27388,N_25774,N_25585);
nor U27389 (N_27389,N_25499,N_25659);
nand U27390 (N_27390,N_26223,N_25457);
nor U27391 (N_27391,N_26022,N_25411);
and U27392 (N_27392,N_26304,N_25438);
xor U27393 (N_27393,N_25933,N_25248);
nand U27394 (N_27394,N_25319,N_26179);
or U27395 (N_27395,N_25940,N_25685);
nor U27396 (N_27396,N_25768,N_26368);
nand U27397 (N_27397,N_25865,N_25944);
or U27398 (N_27398,N_26239,N_25956);
nand U27399 (N_27399,N_25632,N_26022);
and U27400 (N_27400,N_25296,N_26389);
nor U27401 (N_27401,N_25334,N_26165);
xnor U27402 (N_27402,N_25453,N_26298);
and U27403 (N_27403,N_26044,N_25634);
and U27404 (N_27404,N_25940,N_25274);
nor U27405 (N_27405,N_25420,N_25948);
and U27406 (N_27406,N_25766,N_25549);
or U27407 (N_27407,N_25245,N_26312);
nor U27408 (N_27408,N_26353,N_25274);
nor U27409 (N_27409,N_25752,N_25865);
xor U27410 (N_27410,N_26186,N_25725);
nor U27411 (N_27411,N_25300,N_25873);
nor U27412 (N_27412,N_25587,N_26376);
and U27413 (N_27413,N_25341,N_25818);
xnor U27414 (N_27414,N_25704,N_26195);
or U27415 (N_27415,N_25383,N_25354);
nor U27416 (N_27416,N_25430,N_26048);
nor U27417 (N_27417,N_25536,N_26088);
nor U27418 (N_27418,N_25395,N_26382);
or U27419 (N_27419,N_25624,N_26218);
nand U27420 (N_27420,N_26246,N_26248);
nor U27421 (N_27421,N_25867,N_26347);
nand U27422 (N_27422,N_25959,N_25585);
nor U27423 (N_27423,N_25663,N_26132);
nand U27424 (N_27424,N_25557,N_25216);
nand U27425 (N_27425,N_25634,N_25492);
and U27426 (N_27426,N_26369,N_25891);
nand U27427 (N_27427,N_25841,N_25330);
or U27428 (N_27428,N_25642,N_26158);
and U27429 (N_27429,N_26241,N_25865);
nor U27430 (N_27430,N_25843,N_25908);
nand U27431 (N_27431,N_25414,N_25911);
and U27432 (N_27432,N_25818,N_26388);
xor U27433 (N_27433,N_25539,N_25942);
nand U27434 (N_27434,N_25355,N_25360);
xnor U27435 (N_27435,N_26068,N_26040);
and U27436 (N_27436,N_25226,N_26365);
or U27437 (N_27437,N_25923,N_26301);
nor U27438 (N_27438,N_25265,N_25254);
and U27439 (N_27439,N_25304,N_26017);
xnor U27440 (N_27440,N_26156,N_25919);
nand U27441 (N_27441,N_25284,N_25580);
xnor U27442 (N_27442,N_25588,N_25385);
xor U27443 (N_27443,N_25241,N_25897);
nand U27444 (N_27444,N_26050,N_25783);
nor U27445 (N_27445,N_25443,N_25743);
nor U27446 (N_27446,N_26299,N_25574);
or U27447 (N_27447,N_25279,N_25452);
nor U27448 (N_27448,N_25995,N_26046);
or U27449 (N_27449,N_25706,N_26135);
nor U27450 (N_27450,N_25235,N_25666);
nor U27451 (N_27451,N_26166,N_26217);
xnor U27452 (N_27452,N_26032,N_25496);
xnor U27453 (N_27453,N_26381,N_26332);
nor U27454 (N_27454,N_25799,N_26362);
nor U27455 (N_27455,N_25897,N_25620);
xor U27456 (N_27456,N_26184,N_25747);
and U27457 (N_27457,N_25218,N_26073);
nand U27458 (N_27458,N_25754,N_25365);
nand U27459 (N_27459,N_25955,N_25248);
nand U27460 (N_27460,N_26301,N_25676);
nor U27461 (N_27461,N_26305,N_26155);
nor U27462 (N_27462,N_26208,N_25870);
nor U27463 (N_27463,N_25305,N_25750);
nand U27464 (N_27464,N_25878,N_25409);
xor U27465 (N_27465,N_26074,N_25753);
xnor U27466 (N_27466,N_25514,N_25412);
nand U27467 (N_27467,N_25676,N_25385);
and U27468 (N_27468,N_25254,N_25294);
xnor U27469 (N_27469,N_25200,N_25444);
xor U27470 (N_27470,N_26196,N_25414);
nand U27471 (N_27471,N_25651,N_25683);
or U27472 (N_27472,N_25727,N_26397);
nor U27473 (N_27473,N_25685,N_25372);
or U27474 (N_27474,N_25597,N_26022);
nor U27475 (N_27475,N_25688,N_25573);
and U27476 (N_27476,N_26164,N_26211);
nor U27477 (N_27477,N_25552,N_26013);
and U27478 (N_27478,N_25849,N_26098);
or U27479 (N_27479,N_26076,N_25708);
and U27480 (N_27480,N_26371,N_25611);
or U27481 (N_27481,N_25293,N_26223);
xor U27482 (N_27482,N_25925,N_26255);
xor U27483 (N_27483,N_25929,N_25212);
nand U27484 (N_27484,N_26046,N_25787);
or U27485 (N_27485,N_25839,N_25520);
nor U27486 (N_27486,N_25810,N_26108);
nor U27487 (N_27487,N_26318,N_25383);
xnor U27488 (N_27488,N_25525,N_25813);
nor U27489 (N_27489,N_26064,N_25818);
nor U27490 (N_27490,N_25652,N_25251);
nand U27491 (N_27491,N_25953,N_26063);
nor U27492 (N_27492,N_26072,N_25506);
or U27493 (N_27493,N_25963,N_26248);
nand U27494 (N_27494,N_25922,N_26119);
or U27495 (N_27495,N_25906,N_25395);
nor U27496 (N_27496,N_25338,N_25841);
or U27497 (N_27497,N_25448,N_25994);
or U27498 (N_27498,N_26035,N_26014);
and U27499 (N_27499,N_26039,N_25261);
and U27500 (N_27500,N_26337,N_25253);
or U27501 (N_27501,N_25285,N_25506);
or U27502 (N_27502,N_25342,N_26309);
and U27503 (N_27503,N_25409,N_25954);
xnor U27504 (N_27504,N_25441,N_26200);
or U27505 (N_27505,N_25842,N_25669);
nand U27506 (N_27506,N_25760,N_25260);
nand U27507 (N_27507,N_26168,N_26131);
or U27508 (N_27508,N_25869,N_26089);
nor U27509 (N_27509,N_25759,N_25617);
xor U27510 (N_27510,N_26349,N_25466);
nand U27511 (N_27511,N_25513,N_25325);
or U27512 (N_27512,N_25941,N_25421);
nor U27513 (N_27513,N_26067,N_25705);
and U27514 (N_27514,N_26394,N_26268);
nand U27515 (N_27515,N_25332,N_25694);
and U27516 (N_27516,N_25419,N_26249);
or U27517 (N_27517,N_25569,N_25406);
and U27518 (N_27518,N_25384,N_25316);
xnor U27519 (N_27519,N_25946,N_26322);
or U27520 (N_27520,N_26119,N_25625);
nor U27521 (N_27521,N_25385,N_25783);
or U27522 (N_27522,N_26306,N_25965);
nor U27523 (N_27523,N_26191,N_26259);
nand U27524 (N_27524,N_25409,N_25388);
and U27525 (N_27525,N_25316,N_25580);
nand U27526 (N_27526,N_25737,N_25764);
nor U27527 (N_27527,N_25346,N_25755);
nor U27528 (N_27528,N_25406,N_26148);
nand U27529 (N_27529,N_25228,N_25322);
and U27530 (N_27530,N_25405,N_25588);
nor U27531 (N_27531,N_25648,N_25436);
or U27532 (N_27532,N_25392,N_26071);
xnor U27533 (N_27533,N_26196,N_25520);
xnor U27534 (N_27534,N_25774,N_25932);
nand U27535 (N_27535,N_25867,N_25575);
nor U27536 (N_27536,N_25229,N_25542);
nand U27537 (N_27537,N_25509,N_26054);
and U27538 (N_27538,N_26108,N_25828);
xnor U27539 (N_27539,N_25507,N_26293);
xnor U27540 (N_27540,N_26372,N_25833);
nand U27541 (N_27541,N_25286,N_25217);
nor U27542 (N_27542,N_25683,N_25993);
nor U27543 (N_27543,N_25411,N_25338);
or U27544 (N_27544,N_26029,N_26041);
and U27545 (N_27545,N_25857,N_25416);
nand U27546 (N_27546,N_25582,N_26137);
xnor U27547 (N_27547,N_25436,N_25801);
nand U27548 (N_27548,N_26046,N_25789);
and U27549 (N_27549,N_26098,N_26282);
nand U27550 (N_27550,N_25846,N_26101);
nand U27551 (N_27551,N_26131,N_26185);
nand U27552 (N_27552,N_26195,N_25220);
nor U27553 (N_27553,N_26045,N_25465);
xor U27554 (N_27554,N_25323,N_26328);
and U27555 (N_27555,N_26232,N_26197);
nand U27556 (N_27556,N_26013,N_25946);
nand U27557 (N_27557,N_26159,N_26073);
xnor U27558 (N_27558,N_26328,N_26122);
xnor U27559 (N_27559,N_25998,N_25693);
nand U27560 (N_27560,N_25357,N_26248);
nor U27561 (N_27561,N_25549,N_25243);
xor U27562 (N_27562,N_25794,N_25896);
xnor U27563 (N_27563,N_26221,N_25825);
or U27564 (N_27564,N_25304,N_25383);
or U27565 (N_27565,N_26240,N_26193);
and U27566 (N_27566,N_25618,N_25328);
nor U27567 (N_27567,N_26169,N_26113);
xnor U27568 (N_27568,N_25711,N_25529);
nor U27569 (N_27569,N_26011,N_25515);
and U27570 (N_27570,N_26392,N_26042);
nor U27571 (N_27571,N_25710,N_25565);
xnor U27572 (N_27572,N_26025,N_26147);
nor U27573 (N_27573,N_25380,N_25836);
xnor U27574 (N_27574,N_25629,N_25796);
or U27575 (N_27575,N_25418,N_25551);
nand U27576 (N_27576,N_25592,N_25393);
nand U27577 (N_27577,N_26057,N_25559);
nor U27578 (N_27578,N_25283,N_25795);
nand U27579 (N_27579,N_25755,N_26164);
nor U27580 (N_27580,N_26376,N_25964);
nor U27581 (N_27581,N_25551,N_25862);
nand U27582 (N_27582,N_25656,N_25996);
nand U27583 (N_27583,N_25611,N_25279);
nor U27584 (N_27584,N_25242,N_25881);
and U27585 (N_27585,N_25462,N_25610);
nand U27586 (N_27586,N_25736,N_26170);
nor U27587 (N_27587,N_25250,N_26134);
nand U27588 (N_27588,N_25424,N_25899);
nor U27589 (N_27589,N_26030,N_26352);
or U27590 (N_27590,N_26370,N_25310);
and U27591 (N_27591,N_25327,N_25939);
nand U27592 (N_27592,N_25262,N_25907);
or U27593 (N_27593,N_25372,N_25404);
or U27594 (N_27594,N_25212,N_25637);
and U27595 (N_27595,N_26048,N_25408);
xor U27596 (N_27596,N_26030,N_25714);
or U27597 (N_27597,N_25552,N_25654);
xnor U27598 (N_27598,N_25482,N_25364);
or U27599 (N_27599,N_26376,N_25599);
nor U27600 (N_27600,N_27302,N_27482);
or U27601 (N_27601,N_27594,N_26488);
or U27602 (N_27602,N_27458,N_27286);
nor U27603 (N_27603,N_26467,N_26857);
and U27604 (N_27604,N_26730,N_26418);
nor U27605 (N_27605,N_27124,N_27173);
or U27606 (N_27606,N_27100,N_27000);
nor U27607 (N_27607,N_27452,N_27434);
and U27608 (N_27608,N_27298,N_27512);
nor U27609 (N_27609,N_26670,N_26461);
and U27610 (N_27610,N_26469,N_27199);
xnor U27611 (N_27611,N_27561,N_27152);
nand U27612 (N_27612,N_27213,N_27033);
or U27613 (N_27613,N_27589,N_27459);
and U27614 (N_27614,N_27533,N_26801);
or U27615 (N_27615,N_27578,N_26546);
xnor U27616 (N_27616,N_27126,N_27523);
nor U27617 (N_27617,N_26421,N_26847);
and U27618 (N_27618,N_26692,N_27455);
xnor U27619 (N_27619,N_26594,N_27236);
or U27620 (N_27620,N_27392,N_27096);
nand U27621 (N_27621,N_26653,N_27117);
xor U27622 (N_27622,N_26654,N_26498);
and U27623 (N_27623,N_26870,N_27366);
or U27624 (N_27624,N_27277,N_26480);
xor U27625 (N_27625,N_27443,N_26604);
nand U27626 (N_27626,N_26973,N_27294);
nor U27627 (N_27627,N_26872,N_27131);
and U27628 (N_27628,N_26932,N_27371);
or U27629 (N_27629,N_27285,N_26699);
xnor U27630 (N_27630,N_26424,N_27116);
nand U27631 (N_27631,N_26922,N_27529);
nand U27632 (N_27632,N_27361,N_26404);
and U27633 (N_27633,N_27521,N_27164);
and U27634 (N_27634,N_26698,N_27179);
nand U27635 (N_27635,N_26769,N_26568);
xor U27636 (N_27636,N_26431,N_26737);
and U27637 (N_27637,N_26535,N_27065);
and U27638 (N_27638,N_27400,N_26852);
nand U27639 (N_27639,N_27522,N_27421);
nor U27640 (N_27640,N_26685,N_26448);
or U27641 (N_27641,N_26407,N_26758);
and U27642 (N_27642,N_26915,N_26950);
and U27643 (N_27643,N_27046,N_27225);
and U27644 (N_27644,N_27059,N_26457);
xnor U27645 (N_27645,N_27435,N_27386);
or U27646 (N_27646,N_26598,N_26601);
or U27647 (N_27647,N_27022,N_27147);
nor U27648 (N_27648,N_27471,N_26613);
xnor U27649 (N_27649,N_27241,N_26444);
and U27650 (N_27650,N_26731,N_27231);
and U27651 (N_27651,N_27258,N_26716);
and U27652 (N_27652,N_27234,N_27251);
or U27653 (N_27653,N_27353,N_27200);
or U27654 (N_27654,N_26638,N_27399);
or U27655 (N_27655,N_26612,N_26905);
xor U27656 (N_27656,N_27565,N_27429);
nor U27657 (N_27657,N_27584,N_26440);
or U27658 (N_27658,N_27190,N_26773);
nand U27659 (N_27659,N_27352,N_27516);
or U27660 (N_27660,N_27088,N_26865);
xor U27661 (N_27661,N_26624,N_27344);
xor U27662 (N_27662,N_26533,N_27507);
and U27663 (N_27663,N_27182,N_27020);
xnor U27664 (N_27664,N_27233,N_27550);
and U27665 (N_27665,N_27405,N_26800);
nor U27666 (N_27666,N_26539,N_27419);
and U27667 (N_27667,N_26635,N_26762);
and U27668 (N_27668,N_26789,N_26528);
nand U27669 (N_27669,N_27467,N_26400);
xor U27670 (N_27670,N_26556,N_27412);
xor U27671 (N_27671,N_27275,N_26435);
xnor U27672 (N_27672,N_26884,N_26833);
nand U27673 (N_27673,N_26927,N_27138);
nor U27674 (N_27674,N_27016,N_26593);
nor U27675 (N_27675,N_27239,N_26991);
nor U27676 (N_27676,N_27142,N_26456);
and U27677 (N_27677,N_27408,N_26896);
and U27678 (N_27678,N_26999,N_26881);
nand U27679 (N_27679,N_26590,N_27375);
nand U27680 (N_27680,N_26605,N_27268);
and U27681 (N_27681,N_26648,N_27252);
nand U27682 (N_27682,N_27163,N_27490);
or U27683 (N_27683,N_27276,N_26583);
or U27684 (N_27684,N_26840,N_27157);
xor U27685 (N_27685,N_26564,N_27536);
nand U27686 (N_27686,N_27290,N_26453);
xor U27687 (N_27687,N_26610,N_26671);
nand U27688 (N_27688,N_27169,N_27076);
and U27689 (N_27689,N_27530,N_26428);
nand U27690 (N_27690,N_26537,N_26581);
nand U27691 (N_27691,N_27359,N_27247);
or U27692 (N_27692,N_27488,N_26497);
nor U27693 (N_27693,N_26402,N_27205);
xnor U27694 (N_27694,N_27450,N_27288);
nor U27695 (N_27695,N_27278,N_27194);
xor U27696 (N_27696,N_26521,N_27107);
and U27697 (N_27697,N_26708,N_26628);
nand U27698 (N_27698,N_27071,N_26825);
and U27699 (N_27699,N_27201,N_27123);
and U27700 (N_27700,N_27072,N_26874);
and U27701 (N_27701,N_27017,N_26776);
nor U27702 (N_27702,N_26900,N_27040);
xnor U27703 (N_27703,N_26429,N_27484);
nand U27704 (N_27704,N_26458,N_27244);
or U27705 (N_27705,N_26783,N_26484);
and U27706 (N_27706,N_27178,N_26531);
xor U27707 (N_27707,N_27526,N_26586);
or U27708 (N_27708,N_26709,N_26935);
or U27709 (N_27709,N_26961,N_26771);
and U27710 (N_27710,N_27103,N_27240);
nand U27711 (N_27711,N_27214,N_26532);
nand U27712 (N_27712,N_27534,N_27365);
nor U27713 (N_27713,N_27451,N_26942);
or U27714 (N_27714,N_26982,N_26898);
and U27715 (N_27715,N_27255,N_27250);
nor U27716 (N_27716,N_27209,N_26412);
nor U27717 (N_27717,N_26686,N_27402);
xor U27718 (N_27718,N_27041,N_27099);
or U27719 (N_27719,N_27586,N_27326);
and U27720 (N_27720,N_26912,N_26891);
or U27721 (N_27721,N_27069,N_27215);
nand U27722 (N_27722,N_27281,N_26908);
and U27723 (N_27723,N_26669,N_27144);
nor U27724 (N_27724,N_27097,N_26784);
xnor U27725 (N_27725,N_27256,N_27028);
or U27726 (N_27726,N_27008,N_26423);
xnor U27727 (N_27727,N_26554,N_26615);
or U27728 (N_27728,N_27183,N_26657);
nor U27729 (N_27729,N_26466,N_27463);
and U27730 (N_27730,N_26965,N_26502);
and U27731 (N_27731,N_27414,N_26603);
nand U27732 (N_27732,N_26899,N_27440);
or U27733 (N_27733,N_27128,N_27035);
xor U27734 (N_27734,N_27356,N_26637);
nor U27735 (N_27735,N_26565,N_27551);
nor U27736 (N_27736,N_27563,N_26812);
or U27737 (N_27737,N_27162,N_27595);
and U27738 (N_27738,N_26880,N_27259);
xnor U27739 (N_27739,N_27038,N_26634);
and U27740 (N_27740,N_26658,N_27312);
or U27741 (N_27741,N_27360,N_27322);
xor U27742 (N_27742,N_26680,N_27120);
nand U27743 (N_27743,N_27474,N_26958);
or U27744 (N_27744,N_26482,N_26664);
nor U27745 (N_27745,N_26517,N_27125);
nor U27746 (N_27746,N_27525,N_26492);
xnor U27747 (N_27747,N_27106,N_26882);
nor U27748 (N_27748,N_27423,N_27427);
xor U27749 (N_27749,N_26577,N_26678);
or U27750 (N_27750,N_27397,N_27115);
and U27751 (N_27751,N_26726,N_26799);
and U27752 (N_27752,N_26572,N_27051);
nor U27753 (N_27753,N_27101,N_26767);
xnor U27754 (N_27754,N_27153,N_27570);
or U27755 (N_27755,N_26755,N_26720);
or U27756 (N_27756,N_27339,N_26975);
nand U27757 (N_27757,N_26761,N_26968);
nand U27758 (N_27758,N_27401,N_27052);
nor U27759 (N_27759,N_27195,N_27494);
or U27760 (N_27760,N_27393,N_27598);
and U27761 (N_27761,N_26756,N_27465);
nor U27762 (N_27762,N_27461,N_27379);
or U27763 (N_27763,N_27391,N_27568);
xnor U27764 (N_27764,N_26977,N_27282);
or U27765 (N_27765,N_26894,N_27222);
nor U27766 (N_27766,N_27394,N_27274);
nor U27767 (N_27767,N_27407,N_26729);
xnor U27768 (N_27768,N_27506,N_27567);
and U27769 (N_27769,N_27403,N_27166);
nand U27770 (N_27770,N_26401,N_26551);
xnor U27771 (N_27771,N_26588,N_27269);
xor U27772 (N_27772,N_26587,N_27289);
and U27773 (N_27773,N_27350,N_26614);
nand U27774 (N_27774,N_26795,N_27547);
nand U27775 (N_27775,N_26493,N_27495);
nor U27776 (N_27776,N_26510,N_27480);
nor U27777 (N_27777,N_27491,N_27068);
or U27778 (N_27778,N_26681,N_27347);
nand U27779 (N_27779,N_26934,N_26471);
and U27780 (N_27780,N_27420,N_27295);
nor U27781 (N_27781,N_27014,N_26794);
or U27782 (N_27782,N_26607,N_27457);
or U27783 (N_27783,N_26979,N_27082);
and U27784 (N_27784,N_26629,N_26623);
nand U27785 (N_27785,N_27160,N_27517);
xnor U27786 (N_27786,N_27515,N_26793);
nor U27787 (N_27787,N_27242,N_26739);
xor U27788 (N_27788,N_26682,N_26619);
xnor U27789 (N_27789,N_26580,N_26474);
and U27790 (N_27790,N_27029,N_27047);
xnor U27791 (N_27791,N_26436,N_27505);
or U27792 (N_27792,N_27221,N_26640);
nand U27793 (N_27793,N_27389,N_26974);
xor U27794 (N_27794,N_26509,N_26746);
nor U27795 (N_27795,N_27558,N_26515);
nand U27796 (N_27796,N_27409,N_27217);
nand U27797 (N_27797,N_26562,N_26547);
nand U27798 (N_27798,N_26516,N_27431);
nor U27799 (N_27799,N_26750,N_26489);
nand U27800 (N_27800,N_26585,N_26566);
xnor U27801 (N_27801,N_26426,N_27062);
nand U27802 (N_27802,N_27464,N_27304);
nand U27803 (N_27803,N_27532,N_26770);
nor U27804 (N_27804,N_26511,N_26449);
and U27805 (N_27805,N_27030,N_26764);
or U27806 (N_27806,N_26468,N_27470);
or U27807 (N_27807,N_26832,N_26477);
and U27808 (N_27808,N_27219,N_27202);
nor U27809 (N_27809,N_26751,N_27039);
nor U27810 (N_27810,N_27064,N_26667);
nand U27811 (N_27811,N_27486,N_27263);
and U27812 (N_27812,N_26911,N_27098);
nor U27813 (N_27813,N_27546,N_26494);
and U27814 (N_27814,N_26970,N_27541);
and U27815 (N_27815,N_26701,N_27332);
nand U27816 (N_27816,N_27118,N_26529);
and U27817 (N_27817,N_27406,N_26845);
nor U27818 (N_27818,N_27483,N_27024);
or U27819 (N_27819,N_26797,N_27271);
xor U27820 (N_27820,N_27143,N_27552);
xor U27821 (N_27821,N_26443,N_27264);
nand U27822 (N_27822,N_27333,N_27342);
nand U27823 (N_27823,N_26866,N_26867);
xor U27824 (N_27824,N_26486,N_27439);
and U27825 (N_27825,N_26842,N_26557);
xnor U27826 (N_27826,N_26919,N_26943);
and U27827 (N_27827,N_26879,N_26674);
and U27828 (N_27828,N_26707,N_26858);
nor U27829 (N_27829,N_26921,N_26676);
and U27830 (N_27830,N_26505,N_26419);
nand U27831 (N_27831,N_27127,N_26552);
and U27832 (N_27832,N_27500,N_26718);
nand U27833 (N_27833,N_26824,N_26633);
nor U27834 (N_27834,N_27318,N_26988);
xor U27835 (N_27835,N_27243,N_27133);
nor U27836 (N_27836,N_26883,N_26740);
and U27837 (N_27837,N_26976,N_27376);
xor U27838 (N_27838,N_26742,N_26822);
and U27839 (N_27839,N_27137,N_27254);
nor U27840 (N_27840,N_26673,N_26582);
xor U27841 (N_27841,N_26620,N_27001);
or U27842 (N_27842,N_27331,N_26768);
xor U27843 (N_27843,N_26441,N_27354);
and U27844 (N_27844,N_26567,N_27248);
xor U27845 (N_27845,N_26972,N_27167);
xnor U27846 (N_27846,N_27537,N_27575);
nand U27847 (N_27847,N_26873,N_26422);
nor U27848 (N_27848,N_26571,N_26438);
nor U27849 (N_27849,N_26575,N_27577);
or U27850 (N_27850,N_26630,N_26811);
and U27851 (N_27851,N_27544,N_26621);
or U27852 (N_27852,N_26661,N_27300);
nor U27853 (N_27853,N_27102,N_27426);
or U27854 (N_27854,N_26409,N_27003);
nand U27855 (N_27855,N_26893,N_27154);
and U27856 (N_27856,N_27324,N_26570);
and U27857 (N_27857,N_26616,N_26743);
nor U27858 (N_27858,N_26766,N_27364);
nor U27859 (N_27859,N_26775,N_26953);
nor U27860 (N_27860,N_27542,N_27105);
or U27861 (N_27861,N_27338,N_26948);
and U27862 (N_27862,N_26427,N_26817);
nor U27863 (N_27863,N_27398,N_27130);
nor U27864 (N_27864,N_27513,N_27438);
nand U27865 (N_27865,N_27155,N_26821);
or U27866 (N_27866,N_27260,N_27193);
nand U27867 (N_27867,N_26806,N_26536);
xor U27868 (N_27868,N_27496,N_26405);
and U27869 (N_27869,N_26753,N_27023);
and U27870 (N_27870,N_27079,N_27044);
nand U27871 (N_27871,N_26663,N_27572);
nand U27872 (N_27872,N_26446,N_27087);
nor U27873 (N_27873,N_27336,N_27587);
and U27874 (N_27874,N_26837,N_26668);
nand U27875 (N_27875,N_27114,N_27489);
xor U27876 (N_27876,N_26735,N_27381);
nor U27877 (N_27877,N_27232,N_26967);
and U27878 (N_27878,N_26864,N_27502);
nor U27879 (N_27879,N_26715,N_26732);
xor U27880 (N_27880,N_26717,N_26560);
or U27881 (N_27881,N_27206,N_27466);
or U27882 (N_27882,N_26534,N_27504);
nand U27883 (N_27883,N_27372,N_27599);
or U27884 (N_27884,N_26455,N_27368);
xnor U27885 (N_27885,N_26887,N_26785);
xor U27886 (N_27886,N_26597,N_26944);
nor U27887 (N_27887,N_26545,N_27367);
nor U27888 (N_27888,N_27313,N_26490);
nand U27889 (N_27889,N_27385,N_27067);
nand U27890 (N_27890,N_26595,N_26687);
nor U27891 (N_27891,N_27045,N_27210);
xnor U27892 (N_27892,N_26652,N_26544);
nand U27893 (N_27893,N_27272,N_26798);
and U27894 (N_27894,N_27237,N_27198);
nor U27895 (N_27895,N_27334,N_26917);
nor U27896 (N_27896,N_26826,N_26995);
or U27897 (N_27897,N_26719,N_27315);
nand U27898 (N_27898,N_26651,N_26949);
or U27899 (N_27899,N_26838,N_26705);
xnor U27900 (N_27900,N_26553,N_27299);
and U27901 (N_27901,N_27404,N_27086);
and U27902 (N_27902,N_27119,N_27493);
nor U27903 (N_27903,N_26589,N_26791);
nor U27904 (N_27904,N_26454,N_26814);
xnor U27905 (N_27905,N_27091,N_26907);
and U27906 (N_27906,N_26683,N_27306);
or U27907 (N_27907,N_27460,N_26877);
and U27908 (N_27908,N_26713,N_27485);
or U27909 (N_27909,N_26964,N_27170);
or U27910 (N_27910,N_26636,N_26856);
and U27911 (N_27911,N_27519,N_26895);
xnor U27912 (N_27912,N_27329,N_27009);
xnor U27913 (N_27913,N_26875,N_26839);
and U27914 (N_27914,N_27060,N_27284);
or U27915 (N_27915,N_26925,N_26733);
or U27916 (N_27916,N_27187,N_27050);
xnor U27917 (N_27917,N_26960,N_27015);
and U27918 (N_27918,N_26945,N_27553);
nand U27919 (N_27919,N_27596,N_26808);
and U27920 (N_27920,N_26573,N_26788);
nand U27921 (N_27921,N_27005,N_26527);
nor U27922 (N_27922,N_27080,N_26408);
xor U27923 (N_27923,N_27026,N_26631);
and U27924 (N_27924,N_27413,N_27535);
nand U27925 (N_27925,N_26696,N_27238);
or U27926 (N_27926,N_26955,N_27149);
nand U27927 (N_27927,N_27197,N_26869);
xor U27928 (N_27928,N_26650,N_27425);
nor U27929 (N_27929,N_27305,N_26714);
nor U27930 (N_27930,N_27564,N_27223);
nor U27931 (N_27931,N_26828,N_26659);
nand U27932 (N_27932,N_26989,N_27145);
or U27933 (N_27933,N_27063,N_27158);
or U27934 (N_27934,N_26809,N_27084);
nor U27935 (N_27935,N_26969,N_26844);
nand U27936 (N_27936,N_26871,N_26561);
or U27937 (N_27937,N_26748,N_26690);
and U27938 (N_27938,N_26853,N_27025);
nor U27939 (N_27939,N_27432,N_27327);
xnor U27940 (N_27940,N_27077,N_27311);
or U27941 (N_27941,N_27042,N_26816);
nand U27942 (N_27942,N_26888,N_26430);
xnor U27943 (N_27943,N_27321,N_27573);
or U27944 (N_27944,N_26574,N_26689);
or U27945 (N_27945,N_26656,N_26524);
nor U27946 (N_27946,N_27528,N_26928);
nor U27947 (N_27947,N_26736,N_27395);
nor U27948 (N_27948,N_27503,N_26956);
or U27949 (N_27949,N_26622,N_27351);
or U27950 (N_27950,N_26694,N_26823);
xor U27951 (N_27951,N_26897,N_27571);
and U27952 (N_27952,N_27176,N_26555);
nor U27953 (N_27953,N_26886,N_27058);
or U27954 (N_27954,N_26503,N_27235);
nor U27955 (N_27955,N_26706,N_26602);
xnor U27956 (N_27956,N_26963,N_26410);
or U27957 (N_27957,N_27262,N_26542);
and U27958 (N_27958,N_27560,N_27323);
nor U27959 (N_27959,N_27469,N_26578);
and U27960 (N_27960,N_26703,N_26728);
xor U27961 (N_27961,N_27473,N_26414);
xor U27962 (N_27962,N_27418,N_27283);
nand U27963 (N_27963,N_26849,N_27576);
xor U27964 (N_27964,N_26579,N_26757);
xnor U27965 (N_27965,N_27442,N_27267);
and U27966 (N_27966,N_27168,N_27031);
nand U27967 (N_27967,N_26752,N_26804);
or U27968 (N_27968,N_27172,N_26848);
nor U27969 (N_27969,N_27424,N_27095);
or U27970 (N_27970,N_27013,N_26712);
or U27971 (N_27971,N_27441,N_26485);
xor U27972 (N_27972,N_26513,N_27499);
xnor U27973 (N_27973,N_26843,N_27511);
nor U27974 (N_27974,N_27227,N_27390);
xnor U27975 (N_27975,N_26472,N_27061);
and U27976 (N_27976,N_26584,N_26987);
and U27977 (N_27977,N_26666,N_26876);
and U27978 (N_27978,N_26778,N_26786);
nor U27979 (N_27979,N_27348,N_27325);
nor U27980 (N_27980,N_27287,N_26951);
xor U27981 (N_27981,N_26452,N_27411);
xnor U27982 (N_27982,N_27369,N_27184);
or U27983 (N_27983,N_26906,N_26930);
nand U27984 (N_27984,N_26782,N_27510);
xor U27985 (N_27985,N_26918,N_26861);
nor U27986 (N_27986,N_26819,N_27543);
nor U27987 (N_27987,N_26836,N_27027);
and U27988 (N_27988,N_26672,N_26432);
nor U27989 (N_27989,N_27548,N_27316);
xnor U27990 (N_27990,N_26990,N_26941);
xnor U27991 (N_27991,N_27384,N_27557);
nor U27992 (N_27992,N_26563,N_26627);
or U27993 (N_27993,N_27265,N_27337);
and U27994 (N_27994,N_27134,N_26599);
or U27995 (N_27995,N_26914,N_27559);
nor U27996 (N_27996,N_27266,N_27230);
nor U27997 (N_27997,N_26924,N_26507);
or U27998 (N_27998,N_27310,N_26790);
xor U27999 (N_27999,N_26512,N_26998);
xor U28000 (N_28000,N_26996,N_27057);
and U28001 (N_28001,N_26754,N_26491);
or U28002 (N_28002,N_26992,N_27545);
nor U28003 (N_28003,N_27224,N_27446);
nor U28004 (N_28004,N_27211,N_26704);
nand U28005 (N_28005,N_26985,N_26618);
and U28006 (N_28006,N_27218,N_27509);
and U28007 (N_28007,N_27056,N_26643);
nand U28008 (N_28008,N_26966,N_26433);
nand U28009 (N_28009,N_26495,N_27301);
or U28010 (N_28010,N_26983,N_27083);
nand U28011 (N_28011,N_26500,N_27448);
nor U28012 (N_28012,N_26543,N_26462);
nor U28013 (N_28013,N_26781,N_27129);
and U28014 (N_28014,N_27380,N_27357);
nor U28015 (N_28015,N_26846,N_26765);
and U28016 (N_28016,N_27002,N_27109);
nor U28017 (N_28017,N_26530,N_26946);
or U28018 (N_28018,N_26611,N_26451);
nand U28019 (N_28019,N_27475,N_26892);
or U28020 (N_28020,N_27388,N_27518);
xor U28021 (N_28021,N_26541,N_26904);
xnor U28022 (N_28022,N_27019,N_26434);
and U28023 (N_28023,N_27345,N_26608);
or U28024 (N_28024,N_27593,N_26464);
and U28025 (N_28025,N_26600,N_26558);
nor U28026 (N_28026,N_26520,N_26450);
and U28027 (N_28027,N_26649,N_26501);
xor U28028 (N_28028,N_26487,N_27055);
or U28029 (N_28029,N_26576,N_26518);
nand U28030 (N_28030,N_27204,N_26916);
nand U28031 (N_28031,N_27588,N_27520);
nand U28032 (N_28032,N_26695,N_27387);
nor U28033 (N_28033,N_26660,N_27319);
nand U28034 (N_28034,N_27156,N_27280);
and U28035 (N_28035,N_26835,N_26508);
or U28036 (N_28036,N_27454,N_26878);
or U28037 (N_28037,N_26504,N_26459);
nand U28038 (N_28038,N_27362,N_27180);
nand U28039 (N_28039,N_26727,N_27341);
nor U28040 (N_28040,N_26665,N_26841);
or U28041 (N_28041,N_27444,N_27437);
nor U28042 (N_28042,N_26772,N_26747);
and U28043 (N_28043,N_27192,N_27349);
nand U28044 (N_28044,N_26475,N_27591);
or U28045 (N_28045,N_26763,N_27074);
nand U28046 (N_28046,N_26688,N_27292);
or U28047 (N_28047,N_26642,N_26724);
or U28048 (N_28048,N_26416,N_26851);
nor U28049 (N_28049,N_27228,N_26559);
nor U28050 (N_28050,N_27447,N_27108);
xor U28051 (N_28051,N_27508,N_26470);
nor U28052 (N_28052,N_26863,N_27245);
xor U28053 (N_28053,N_27492,N_27415);
nand U28054 (N_28054,N_27358,N_27478);
and U28055 (N_28055,N_26417,N_26465);
and U28056 (N_28056,N_27132,N_26437);
and U28057 (N_28057,N_26978,N_27580);
or U28058 (N_28058,N_26679,N_26700);
nand U28059 (N_28059,N_27073,N_27186);
nand U28060 (N_28060,N_27161,N_27497);
xor U28061 (N_28061,N_27273,N_27346);
and U28062 (N_28062,N_26954,N_26854);
and U28063 (N_28063,N_27212,N_26827);
nor U28064 (N_28064,N_26420,N_27297);
and U28065 (N_28065,N_26971,N_26933);
xnor U28066 (N_28066,N_26805,N_27246);
nand U28067 (N_28067,N_27092,N_27032);
nand U28068 (N_28068,N_27075,N_26749);
or U28069 (N_28069,N_27081,N_26994);
or U28070 (N_28070,N_26473,N_27396);
nand U28071 (N_28071,N_27150,N_27066);
and U28072 (N_28072,N_27151,N_27549);
nand U28073 (N_28073,N_27257,N_26818);
or U28074 (N_28074,N_27472,N_27481);
nand U28075 (N_28075,N_26980,N_26926);
nand U28076 (N_28076,N_26831,N_26759);
xnor U28077 (N_28077,N_26738,N_26403);
or U28078 (N_28078,N_27208,N_26890);
and U28079 (N_28079,N_26425,N_26862);
nand U28080 (N_28080,N_26939,N_27383);
or U28081 (N_28081,N_26721,N_26777);
or U28082 (N_28082,N_26675,N_26910);
or U28083 (N_28083,N_26929,N_26850);
nand U28084 (N_28084,N_27462,N_26885);
or U28085 (N_28085,N_27456,N_27279);
nor U28086 (N_28086,N_27514,N_26936);
nor U28087 (N_28087,N_27196,N_27216);
xor U28088 (N_28088,N_27307,N_26780);
nand U28089 (N_28089,N_27539,N_26646);
and U28090 (N_28090,N_27177,N_27185);
nand U28091 (N_28091,N_27078,N_27317);
and U28092 (N_28092,N_27007,N_26962);
or U28093 (N_28093,N_27363,N_26460);
nor U28094 (N_28094,N_26413,N_26802);
xor U28095 (N_28095,N_26957,N_26483);
xnor U28096 (N_28096,N_27468,N_27090);
and U28097 (N_28097,N_26984,N_26855);
nand U28098 (N_28098,N_26442,N_27012);
and U28099 (N_28099,N_26596,N_26986);
nand U28100 (N_28100,N_27527,N_27370);
nor U28101 (N_28101,N_26923,N_26496);
and U28102 (N_28102,N_27135,N_27165);
or U28103 (N_28103,N_27487,N_27270);
nor U28104 (N_28104,N_27094,N_27085);
or U28105 (N_28105,N_27328,N_26940);
xor U28106 (N_28106,N_27422,N_26645);
xor U28107 (N_28107,N_26445,N_27382);
xor U28108 (N_28108,N_26981,N_26815);
or U28109 (N_28109,N_26725,N_26523);
nor U28110 (N_28110,N_27181,N_27374);
nor U28111 (N_28111,N_27261,N_27556);
nand U28112 (N_28112,N_27036,N_27122);
and U28113 (N_28113,N_27189,N_27188);
xor U28114 (N_28114,N_26702,N_26909);
and U28115 (N_28115,N_27582,N_26813);
or U28116 (N_28116,N_27226,N_27428);
nor U28117 (N_28117,N_27476,N_26820);
or U28118 (N_28118,N_26463,N_27191);
xnor U28119 (N_28119,N_26774,N_26744);
xor U28120 (N_28120,N_26807,N_26830);
and U28121 (N_28121,N_27569,N_27378);
nor U28122 (N_28122,N_26525,N_27579);
nor U28123 (N_28123,N_27416,N_27340);
nand U28124 (N_28124,N_27111,N_27112);
nor U28125 (N_28125,N_27597,N_26760);
and U28126 (N_28126,N_27436,N_27498);
nand U28127 (N_28127,N_26889,N_27253);
nand U28128 (N_28128,N_26609,N_27291);
nand U28129 (N_28129,N_26641,N_26522);
nand U28130 (N_28130,N_26632,N_26903);
nor U28131 (N_28131,N_27034,N_27159);
and U28132 (N_28132,N_26506,N_27175);
xor U28133 (N_28133,N_27430,N_27110);
or U28134 (N_28134,N_26592,N_27320);
nand U28135 (N_28135,N_27053,N_26476);
or U28136 (N_28136,N_26796,N_26406);
xnor U28137 (N_28137,N_27136,N_26693);
nor U28138 (N_28138,N_27308,N_26745);
xor U28139 (N_28139,N_26859,N_27583);
or U28140 (N_28140,N_26734,N_26550);
or U28141 (N_28141,N_26415,N_26540);
and U28142 (N_28142,N_26792,N_26677);
nand U28143 (N_28143,N_26947,N_26519);
nor U28144 (N_28144,N_27574,N_26834);
or U28145 (N_28145,N_27174,N_27449);
nand U28146 (N_28146,N_27011,N_26868);
nand U28147 (N_28147,N_27140,N_26959);
nor U28148 (N_28148,N_27296,N_27229);
and U28149 (N_28149,N_26691,N_27540);
nand U28150 (N_28150,N_26993,N_26478);
xor U28151 (N_28151,N_26447,N_27141);
nor U28152 (N_28152,N_27538,N_26913);
xnor U28153 (N_28153,N_26779,N_27330);
and U28154 (N_28154,N_26549,N_26514);
and U28155 (N_28155,N_27343,N_26787);
or U28156 (N_28156,N_27021,N_27203);
nand U28157 (N_28157,N_26499,N_27146);
or U28158 (N_28158,N_27148,N_26526);
xor U28159 (N_28159,N_27335,N_26625);
xnor U28160 (N_28160,N_26684,N_27433);
or U28161 (N_28161,N_26860,N_27585);
and U28162 (N_28162,N_26829,N_27581);
and U28163 (N_28163,N_27048,N_26711);
and U28164 (N_28164,N_27453,N_27089);
xnor U28165 (N_28165,N_27037,N_27043);
and U28166 (N_28166,N_27093,N_27006);
nor U28167 (N_28167,N_26997,N_27314);
nand U28168 (N_28168,N_26803,N_27355);
nor U28169 (N_28169,N_27477,N_26655);
or U28170 (N_28170,N_26723,N_27377);
nand U28171 (N_28171,N_27410,N_27524);
nand U28172 (N_28172,N_26647,N_26548);
or U28173 (N_28173,N_26617,N_27054);
xnor U28174 (N_28174,N_26411,N_26538);
nand U28175 (N_28175,N_27139,N_26697);
xnor U28176 (N_28176,N_27113,N_27104);
and U28177 (N_28177,N_27479,N_26626);
or U28178 (N_28178,N_26952,N_27555);
or U28179 (N_28179,N_27049,N_26937);
and U28180 (N_28180,N_26481,N_27018);
nor U28181 (N_28181,N_27004,N_26902);
xor U28182 (N_28182,N_26479,N_26569);
or U28183 (N_28183,N_26606,N_27562);
nand U28184 (N_28184,N_26810,N_27592);
and U28185 (N_28185,N_27309,N_26662);
xnor U28186 (N_28186,N_27417,N_27566);
or U28187 (N_28187,N_26938,N_27220);
nand U28188 (N_28188,N_27445,N_27121);
nand U28189 (N_28189,N_26710,N_27171);
and U28190 (N_28190,N_26931,N_26722);
and U28191 (N_28191,N_27554,N_26741);
nand U28192 (N_28192,N_27010,N_27501);
and U28193 (N_28193,N_26439,N_27531);
xor U28194 (N_28194,N_26901,N_26639);
or U28195 (N_28195,N_27590,N_27303);
or U28196 (N_28196,N_27249,N_27373);
or U28197 (N_28197,N_27070,N_26920);
nor U28198 (N_28198,N_26591,N_27293);
nand U28199 (N_28199,N_27207,N_26644);
and U28200 (N_28200,N_27106,N_26870);
nor U28201 (N_28201,N_26487,N_27512);
or U28202 (N_28202,N_26402,N_26503);
xnor U28203 (N_28203,N_27004,N_27529);
nand U28204 (N_28204,N_27524,N_26838);
or U28205 (N_28205,N_27183,N_27581);
or U28206 (N_28206,N_26836,N_26525);
nor U28207 (N_28207,N_27189,N_26612);
nor U28208 (N_28208,N_26905,N_26869);
and U28209 (N_28209,N_26567,N_26575);
xnor U28210 (N_28210,N_27208,N_26480);
and U28211 (N_28211,N_27147,N_27355);
nand U28212 (N_28212,N_27424,N_27184);
nor U28213 (N_28213,N_27416,N_26664);
xor U28214 (N_28214,N_27487,N_27304);
xor U28215 (N_28215,N_27210,N_26683);
nand U28216 (N_28216,N_26579,N_27356);
or U28217 (N_28217,N_26440,N_26792);
nor U28218 (N_28218,N_26878,N_26763);
xnor U28219 (N_28219,N_26635,N_27069);
nor U28220 (N_28220,N_26967,N_27375);
nor U28221 (N_28221,N_27535,N_26862);
and U28222 (N_28222,N_27169,N_26578);
or U28223 (N_28223,N_26442,N_26856);
nand U28224 (N_28224,N_26764,N_26849);
or U28225 (N_28225,N_26977,N_27154);
nand U28226 (N_28226,N_26693,N_26843);
and U28227 (N_28227,N_27292,N_27341);
nand U28228 (N_28228,N_26574,N_27220);
and U28229 (N_28229,N_26625,N_27425);
nand U28230 (N_28230,N_27495,N_26609);
xnor U28231 (N_28231,N_27565,N_27037);
and U28232 (N_28232,N_26691,N_27538);
or U28233 (N_28233,N_26921,N_27484);
nor U28234 (N_28234,N_27051,N_27104);
xor U28235 (N_28235,N_26739,N_26737);
or U28236 (N_28236,N_27270,N_26959);
or U28237 (N_28237,N_26854,N_27324);
nand U28238 (N_28238,N_26542,N_26961);
xnor U28239 (N_28239,N_27441,N_26766);
nand U28240 (N_28240,N_27255,N_27146);
nor U28241 (N_28241,N_27111,N_26983);
xor U28242 (N_28242,N_26723,N_26662);
nand U28243 (N_28243,N_26558,N_27022);
nand U28244 (N_28244,N_26706,N_26827);
and U28245 (N_28245,N_27206,N_26644);
or U28246 (N_28246,N_27254,N_27208);
and U28247 (N_28247,N_26839,N_26760);
and U28248 (N_28248,N_27107,N_26719);
or U28249 (N_28249,N_26439,N_26422);
nor U28250 (N_28250,N_27131,N_26436);
nand U28251 (N_28251,N_26612,N_26497);
or U28252 (N_28252,N_26581,N_26843);
or U28253 (N_28253,N_26985,N_26683);
nor U28254 (N_28254,N_27043,N_26866);
nor U28255 (N_28255,N_27144,N_26722);
or U28256 (N_28256,N_26884,N_26675);
xnor U28257 (N_28257,N_26997,N_26457);
xnor U28258 (N_28258,N_26440,N_27237);
nor U28259 (N_28259,N_27597,N_27116);
nand U28260 (N_28260,N_26885,N_27230);
nand U28261 (N_28261,N_27107,N_26592);
and U28262 (N_28262,N_26985,N_27552);
nor U28263 (N_28263,N_27159,N_27204);
and U28264 (N_28264,N_27282,N_26443);
nand U28265 (N_28265,N_27386,N_27157);
and U28266 (N_28266,N_26604,N_26743);
or U28267 (N_28267,N_27381,N_26738);
and U28268 (N_28268,N_26707,N_27485);
xnor U28269 (N_28269,N_27421,N_26535);
nor U28270 (N_28270,N_26678,N_27330);
or U28271 (N_28271,N_26505,N_27221);
and U28272 (N_28272,N_26473,N_27350);
xor U28273 (N_28273,N_26474,N_27263);
nor U28274 (N_28274,N_27291,N_26762);
xor U28275 (N_28275,N_27107,N_27409);
and U28276 (N_28276,N_26940,N_27230);
and U28277 (N_28277,N_26661,N_27449);
xnor U28278 (N_28278,N_26562,N_26958);
or U28279 (N_28279,N_26991,N_27481);
nor U28280 (N_28280,N_27443,N_27472);
nor U28281 (N_28281,N_26685,N_27002);
nor U28282 (N_28282,N_27356,N_26890);
nand U28283 (N_28283,N_26546,N_26628);
and U28284 (N_28284,N_27179,N_27120);
nor U28285 (N_28285,N_27488,N_27510);
nor U28286 (N_28286,N_26490,N_26907);
and U28287 (N_28287,N_27025,N_27243);
xnor U28288 (N_28288,N_27460,N_26658);
nand U28289 (N_28289,N_26916,N_27019);
and U28290 (N_28290,N_26501,N_26668);
nand U28291 (N_28291,N_26455,N_27140);
or U28292 (N_28292,N_27323,N_27204);
and U28293 (N_28293,N_27007,N_27331);
nor U28294 (N_28294,N_27027,N_26905);
xor U28295 (N_28295,N_27232,N_26801);
nor U28296 (N_28296,N_26842,N_26630);
and U28297 (N_28297,N_27001,N_27525);
nor U28298 (N_28298,N_27005,N_27369);
xnor U28299 (N_28299,N_26467,N_26665);
and U28300 (N_28300,N_27408,N_26841);
nor U28301 (N_28301,N_26699,N_27015);
nor U28302 (N_28302,N_26997,N_27071);
and U28303 (N_28303,N_26948,N_27352);
nor U28304 (N_28304,N_26691,N_27185);
nor U28305 (N_28305,N_27222,N_26644);
nand U28306 (N_28306,N_26978,N_26944);
nand U28307 (N_28307,N_27390,N_26644);
and U28308 (N_28308,N_26777,N_27256);
nand U28309 (N_28309,N_26703,N_26556);
or U28310 (N_28310,N_26573,N_26896);
xor U28311 (N_28311,N_27008,N_27325);
xor U28312 (N_28312,N_26440,N_27311);
nand U28313 (N_28313,N_26886,N_27550);
or U28314 (N_28314,N_27472,N_26596);
nand U28315 (N_28315,N_26656,N_27564);
and U28316 (N_28316,N_27136,N_27391);
nand U28317 (N_28317,N_27109,N_27392);
or U28318 (N_28318,N_26909,N_27455);
xnor U28319 (N_28319,N_26883,N_26412);
nand U28320 (N_28320,N_27215,N_27406);
nand U28321 (N_28321,N_26438,N_26827);
nand U28322 (N_28322,N_27000,N_26455);
nor U28323 (N_28323,N_26808,N_27477);
or U28324 (N_28324,N_26903,N_27331);
xor U28325 (N_28325,N_26585,N_26489);
nand U28326 (N_28326,N_27487,N_26699);
nand U28327 (N_28327,N_26938,N_27456);
nand U28328 (N_28328,N_27529,N_26730);
or U28329 (N_28329,N_27402,N_26859);
and U28330 (N_28330,N_27416,N_26476);
xor U28331 (N_28331,N_27374,N_26944);
or U28332 (N_28332,N_27330,N_27456);
xor U28333 (N_28333,N_26796,N_27213);
nor U28334 (N_28334,N_26641,N_27182);
nand U28335 (N_28335,N_26838,N_26993);
nand U28336 (N_28336,N_26906,N_26464);
and U28337 (N_28337,N_27410,N_26647);
and U28338 (N_28338,N_27396,N_27407);
or U28339 (N_28339,N_26651,N_26472);
and U28340 (N_28340,N_27556,N_27044);
nor U28341 (N_28341,N_27384,N_26793);
nand U28342 (N_28342,N_27338,N_27100);
xnor U28343 (N_28343,N_27181,N_26541);
nand U28344 (N_28344,N_26451,N_26590);
and U28345 (N_28345,N_26519,N_27188);
xor U28346 (N_28346,N_26566,N_26875);
and U28347 (N_28347,N_26915,N_26584);
or U28348 (N_28348,N_27352,N_26427);
nand U28349 (N_28349,N_26999,N_27552);
nand U28350 (N_28350,N_26984,N_26514);
and U28351 (N_28351,N_26774,N_26650);
and U28352 (N_28352,N_26695,N_27398);
nor U28353 (N_28353,N_26425,N_26536);
nor U28354 (N_28354,N_26846,N_26866);
and U28355 (N_28355,N_26659,N_27438);
nor U28356 (N_28356,N_26474,N_26414);
xor U28357 (N_28357,N_26587,N_27389);
or U28358 (N_28358,N_26925,N_27340);
or U28359 (N_28359,N_27299,N_26497);
xnor U28360 (N_28360,N_27288,N_27397);
xor U28361 (N_28361,N_26676,N_27010);
nand U28362 (N_28362,N_26912,N_26827);
or U28363 (N_28363,N_27261,N_26535);
or U28364 (N_28364,N_27432,N_26463);
nand U28365 (N_28365,N_27135,N_27311);
nand U28366 (N_28366,N_27342,N_26779);
nor U28367 (N_28367,N_26576,N_26806);
nand U28368 (N_28368,N_27028,N_27140);
nor U28369 (N_28369,N_26539,N_26886);
and U28370 (N_28370,N_26901,N_27158);
or U28371 (N_28371,N_27351,N_27378);
and U28372 (N_28372,N_26570,N_27599);
or U28373 (N_28373,N_26538,N_27511);
xnor U28374 (N_28374,N_27252,N_27225);
nand U28375 (N_28375,N_27527,N_27154);
nand U28376 (N_28376,N_27326,N_27004);
xor U28377 (N_28377,N_27537,N_27338);
nor U28378 (N_28378,N_27591,N_27395);
or U28379 (N_28379,N_27203,N_27254);
nor U28380 (N_28380,N_27327,N_26562);
and U28381 (N_28381,N_27024,N_27018);
xnor U28382 (N_28382,N_26568,N_27347);
or U28383 (N_28383,N_26696,N_27095);
nor U28384 (N_28384,N_27037,N_27459);
nand U28385 (N_28385,N_26518,N_26925);
nand U28386 (N_28386,N_26870,N_26982);
nor U28387 (N_28387,N_27256,N_27517);
nor U28388 (N_28388,N_27352,N_26747);
xnor U28389 (N_28389,N_26667,N_26685);
nand U28390 (N_28390,N_27131,N_27454);
and U28391 (N_28391,N_26929,N_26640);
nand U28392 (N_28392,N_26570,N_27231);
nor U28393 (N_28393,N_27570,N_26510);
and U28394 (N_28394,N_26514,N_27110);
xor U28395 (N_28395,N_26473,N_26582);
xor U28396 (N_28396,N_27447,N_27254);
nand U28397 (N_28397,N_26776,N_26866);
or U28398 (N_28398,N_26515,N_27003);
or U28399 (N_28399,N_26848,N_27323);
or U28400 (N_28400,N_27461,N_26802);
and U28401 (N_28401,N_26609,N_27353);
nor U28402 (N_28402,N_26802,N_27290);
nand U28403 (N_28403,N_27294,N_26923);
nand U28404 (N_28404,N_27048,N_26895);
nor U28405 (N_28405,N_26876,N_26452);
xor U28406 (N_28406,N_27263,N_26964);
or U28407 (N_28407,N_26882,N_27516);
or U28408 (N_28408,N_26843,N_26859);
or U28409 (N_28409,N_27357,N_27081);
xnor U28410 (N_28410,N_26758,N_27197);
xnor U28411 (N_28411,N_27483,N_26580);
xnor U28412 (N_28412,N_26684,N_27212);
xor U28413 (N_28413,N_26874,N_27152);
and U28414 (N_28414,N_27449,N_26974);
nor U28415 (N_28415,N_26534,N_26496);
nor U28416 (N_28416,N_26574,N_27451);
nor U28417 (N_28417,N_27125,N_26603);
or U28418 (N_28418,N_26799,N_27367);
nand U28419 (N_28419,N_26615,N_26486);
nand U28420 (N_28420,N_26444,N_27152);
nand U28421 (N_28421,N_26493,N_27162);
nand U28422 (N_28422,N_26501,N_27512);
and U28423 (N_28423,N_27104,N_26536);
nor U28424 (N_28424,N_26505,N_27285);
nand U28425 (N_28425,N_27364,N_27424);
nand U28426 (N_28426,N_27551,N_27129);
and U28427 (N_28427,N_27033,N_27400);
nand U28428 (N_28428,N_26656,N_26608);
xor U28429 (N_28429,N_27212,N_27010);
and U28430 (N_28430,N_27487,N_27599);
nor U28431 (N_28431,N_27503,N_27283);
xor U28432 (N_28432,N_27476,N_26542);
xor U28433 (N_28433,N_26564,N_27240);
xnor U28434 (N_28434,N_27061,N_26409);
nand U28435 (N_28435,N_27234,N_27150);
xnor U28436 (N_28436,N_26521,N_27311);
nor U28437 (N_28437,N_26410,N_26728);
nand U28438 (N_28438,N_26488,N_27582);
xor U28439 (N_28439,N_26857,N_26722);
nor U28440 (N_28440,N_27039,N_27131);
and U28441 (N_28441,N_27489,N_26587);
or U28442 (N_28442,N_27452,N_27229);
nand U28443 (N_28443,N_26886,N_27118);
xnor U28444 (N_28444,N_26715,N_26424);
and U28445 (N_28445,N_27105,N_26955);
or U28446 (N_28446,N_27544,N_27400);
and U28447 (N_28447,N_27469,N_27464);
xnor U28448 (N_28448,N_27357,N_27053);
nor U28449 (N_28449,N_27151,N_26945);
and U28450 (N_28450,N_27281,N_26778);
and U28451 (N_28451,N_27188,N_26948);
xor U28452 (N_28452,N_27361,N_26628);
or U28453 (N_28453,N_27264,N_27479);
or U28454 (N_28454,N_26762,N_27076);
nor U28455 (N_28455,N_27195,N_27350);
nand U28456 (N_28456,N_27041,N_26787);
or U28457 (N_28457,N_26653,N_26598);
nor U28458 (N_28458,N_27398,N_27459);
and U28459 (N_28459,N_27472,N_26611);
nor U28460 (N_28460,N_26683,N_26919);
nor U28461 (N_28461,N_26843,N_26844);
nor U28462 (N_28462,N_26629,N_27378);
and U28463 (N_28463,N_26400,N_26926);
nand U28464 (N_28464,N_27305,N_27117);
nor U28465 (N_28465,N_26680,N_26991);
xnor U28466 (N_28466,N_26505,N_26940);
xnor U28467 (N_28467,N_27383,N_27291);
nand U28468 (N_28468,N_26956,N_26646);
and U28469 (N_28469,N_26528,N_26803);
nand U28470 (N_28470,N_27566,N_27333);
nor U28471 (N_28471,N_27519,N_26576);
xnor U28472 (N_28472,N_26805,N_26836);
and U28473 (N_28473,N_27182,N_26974);
or U28474 (N_28474,N_26757,N_26937);
and U28475 (N_28475,N_27255,N_26483);
and U28476 (N_28476,N_26456,N_26516);
nor U28477 (N_28477,N_26582,N_26512);
nand U28478 (N_28478,N_26781,N_26981);
nor U28479 (N_28479,N_27198,N_27300);
xor U28480 (N_28480,N_26948,N_26523);
and U28481 (N_28481,N_26758,N_27194);
xor U28482 (N_28482,N_27322,N_27195);
xor U28483 (N_28483,N_27041,N_26885);
nand U28484 (N_28484,N_26649,N_27156);
nor U28485 (N_28485,N_26523,N_27450);
nand U28486 (N_28486,N_26684,N_26563);
nor U28487 (N_28487,N_27015,N_27140);
nand U28488 (N_28488,N_26764,N_27147);
or U28489 (N_28489,N_27157,N_27292);
nand U28490 (N_28490,N_27388,N_26677);
nand U28491 (N_28491,N_27266,N_27026);
xnor U28492 (N_28492,N_27031,N_27327);
and U28493 (N_28493,N_27093,N_27162);
and U28494 (N_28494,N_26828,N_26897);
and U28495 (N_28495,N_26810,N_27071);
or U28496 (N_28496,N_26444,N_27314);
nand U28497 (N_28497,N_27249,N_26429);
xor U28498 (N_28498,N_27581,N_26425);
xor U28499 (N_28499,N_27503,N_27329);
xnor U28500 (N_28500,N_26457,N_27058);
and U28501 (N_28501,N_27380,N_27277);
nand U28502 (N_28502,N_27415,N_26899);
and U28503 (N_28503,N_26870,N_26817);
or U28504 (N_28504,N_26993,N_26678);
nand U28505 (N_28505,N_27271,N_27252);
or U28506 (N_28506,N_26934,N_26524);
or U28507 (N_28507,N_26867,N_26472);
nor U28508 (N_28508,N_27204,N_26564);
or U28509 (N_28509,N_26714,N_26477);
xnor U28510 (N_28510,N_27123,N_26878);
xnor U28511 (N_28511,N_27457,N_26936);
or U28512 (N_28512,N_26998,N_27284);
nand U28513 (N_28513,N_27373,N_27191);
or U28514 (N_28514,N_26810,N_27128);
or U28515 (N_28515,N_27418,N_27206);
nand U28516 (N_28516,N_27443,N_26670);
nand U28517 (N_28517,N_27220,N_27428);
nor U28518 (N_28518,N_27240,N_27124);
and U28519 (N_28519,N_26651,N_27081);
nand U28520 (N_28520,N_27495,N_27560);
or U28521 (N_28521,N_26632,N_26723);
nor U28522 (N_28522,N_26663,N_27227);
xor U28523 (N_28523,N_27278,N_26896);
nor U28524 (N_28524,N_27057,N_26640);
nand U28525 (N_28525,N_27538,N_27584);
or U28526 (N_28526,N_27540,N_27117);
or U28527 (N_28527,N_27408,N_26686);
and U28528 (N_28528,N_27259,N_26955);
nand U28529 (N_28529,N_26986,N_27418);
or U28530 (N_28530,N_26531,N_26956);
nor U28531 (N_28531,N_26904,N_27085);
nor U28532 (N_28532,N_26530,N_27479);
or U28533 (N_28533,N_26513,N_27079);
and U28534 (N_28534,N_27095,N_26479);
nand U28535 (N_28535,N_26874,N_26552);
nand U28536 (N_28536,N_27027,N_27408);
and U28537 (N_28537,N_27367,N_26549);
nand U28538 (N_28538,N_26860,N_26598);
nor U28539 (N_28539,N_26425,N_26725);
and U28540 (N_28540,N_26873,N_27389);
and U28541 (N_28541,N_26695,N_27367);
nor U28542 (N_28542,N_26786,N_26720);
nor U28543 (N_28543,N_27264,N_26599);
xnor U28544 (N_28544,N_26937,N_26767);
and U28545 (N_28545,N_27500,N_26653);
nand U28546 (N_28546,N_27307,N_26860);
xnor U28547 (N_28547,N_27539,N_26800);
nand U28548 (N_28548,N_27551,N_27409);
or U28549 (N_28549,N_26526,N_26811);
and U28550 (N_28550,N_27555,N_26706);
or U28551 (N_28551,N_26795,N_27149);
and U28552 (N_28552,N_26628,N_27345);
nand U28553 (N_28553,N_26643,N_27224);
and U28554 (N_28554,N_26648,N_26714);
and U28555 (N_28555,N_26508,N_26969);
nand U28556 (N_28556,N_27020,N_26521);
nor U28557 (N_28557,N_27106,N_27236);
nand U28558 (N_28558,N_27498,N_27112);
nor U28559 (N_28559,N_27463,N_26463);
xnor U28560 (N_28560,N_26946,N_27569);
and U28561 (N_28561,N_26719,N_26423);
xor U28562 (N_28562,N_27099,N_26966);
or U28563 (N_28563,N_27096,N_27112);
or U28564 (N_28564,N_26585,N_27105);
nand U28565 (N_28565,N_27561,N_27155);
nor U28566 (N_28566,N_27330,N_27216);
nand U28567 (N_28567,N_27574,N_27505);
and U28568 (N_28568,N_26460,N_26633);
and U28569 (N_28569,N_26762,N_27586);
nand U28570 (N_28570,N_27509,N_27283);
nor U28571 (N_28571,N_27316,N_26850);
nor U28572 (N_28572,N_27594,N_27583);
nand U28573 (N_28573,N_26496,N_26780);
nor U28574 (N_28574,N_26475,N_26815);
and U28575 (N_28575,N_26896,N_26492);
xnor U28576 (N_28576,N_26918,N_27301);
nand U28577 (N_28577,N_27425,N_27174);
and U28578 (N_28578,N_26763,N_27107);
or U28579 (N_28579,N_26734,N_27166);
nor U28580 (N_28580,N_26582,N_26671);
or U28581 (N_28581,N_26645,N_27294);
nor U28582 (N_28582,N_26470,N_26984);
or U28583 (N_28583,N_26562,N_27589);
xnor U28584 (N_28584,N_26922,N_26860);
or U28585 (N_28585,N_26458,N_26536);
nand U28586 (N_28586,N_26433,N_26783);
xnor U28587 (N_28587,N_27345,N_27185);
nand U28588 (N_28588,N_26440,N_26694);
and U28589 (N_28589,N_27392,N_26758);
nand U28590 (N_28590,N_26711,N_27404);
xor U28591 (N_28591,N_27050,N_27535);
xnor U28592 (N_28592,N_27474,N_27108);
nor U28593 (N_28593,N_26662,N_26888);
nor U28594 (N_28594,N_27166,N_27379);
xor U28595 (N_28595,N_26401,N_27258);
nand U28596 (N_28596,N_26866,N_26813);
nor U28597 (N_28597,N_26772,N_26660);
or U28598 (N_28598,N_27259,N_27526);
xnor U28599 (N_28599,N_26697,N_27042);
nor U28600 (N_28600,N_27293,N_27477);
nor U28601 (N_28601,N_26503,N_27198);
nor U28602 (N_28602,N_26863,N_27163);
nor U28603 (N_28603,N_27271,N_27184);
nand U28604 (N_28604,N_26604,N_27021);
nand U28605 (N_28605,N_26826,N_27591);
nor U28606 (N_28606,N_26742,N_27360);
or U28607 (N_28607,N_27461,N_27056);
or U28608 (N_28608,N_27436,N_26815);
xnor U28609 (N_28609,N_27174,N_26929);
xnor U28610 (N_28610,N_27586,N_27417);
nor U28611 (N_28611,N_27090,N_27524);
and U28612 (N_28612,N_26965,N_27136);
or U28613 (N_28613,N_27408,N_27058);
nand U28614 (N_28614,N_26939,N_26542);
xnor U28615 (N_28615,N_26606,N_26825);
and U28616 (N_28616,N_27141,N_27069);
or U28617 (N_28617,N_26563,N_26741);
and U28618 (N_28618,N_27097,N_27552);
or U28619 (N_28619,N_27107,N_26431);
nor U28620 (N_28620,N_27166,N_26639);
or U28621 (N_28621,N_26513,N_26414);
nor U28622 (N_28622,N_26941,N_27233);
or U28623 (N_28623,N_26511,N_27384);
nand U28624 (N_28624,N_27247,N_26704);
or U28625 (N_28625,N_26572,N_27462);
or U28626 (N_28626,N_27264,N_26775);
xor U28627 (N_28627,N_27254,N_26605);
nand U28628 (N_28628,N_26804,N_26533);
nor U28629 (N_28629,N_26819,N_26533);
nor U28630 (N_28630,N_26947,N_26443);
xnor U28631 (N_28631,N_26477,N_27367);
and U28632 (N_28632,N_26915,N_26972);
nand U28633 (N_28633,N_27116,N_27297);
or U28634 (N_28634,N_27161,N_26413);
or U28635 (N_28635,N_27431,N_26924);
xor U28636 (N_28636,N_26730,N_27452);
nor U28637 (N_28637,N_27412,N_26739);
or U28638 (N_28638,N_26434,N_26519);
or U28639 (N_28639,N_27328,N_26454);
nand U28640 (N_28640,N_26571,N_27249);
and U28641 (N_28641,N_27225,N_27080);
nand U28642 (N_28642,N_26526,N_27426);
xor U28643 (N_28643,N_27004,N_27462);
nor U28644 (N_28644,N_26729,N_26538);
nor U28645 (N_28645,N_26574,N_27225);
or U28646 (N_28646,N_27453,N_27120);
and U28647 (N_28647,N_27303,N_26740);
nand U28648 (N_28648,N_26850,N_26969);
nor U28649 (N_28649,N_26663,N_27460);
xor U28650 (N_28650,N_27014,N_26831);
or U28651 (N_28651,N_27267,N_26543);
nor U28652 (N_28652,N_26579,N_26823);
xnor U28653 (N_28653,N_26669,N_26982);
nand U28654 (N_28654,N_27363,N_26566);
and U28655 (N_28655,N_27057,N_26540);
and U28656 (N_28656,N_26660,N_27356);
xnor U28657 (N_28657,N_27263,N_27563);
nand U28658 (N_28658,N_27243,N_26611);
xnor U28659 (N_28659,N_26572,N_26960);
nand U28660 (N_28660,N_26638,N_26683);
nor U28661 (N_28661,N_27147,N_27357);
xor U28662 (N_28662,N_26707,N_27410);
or U28663 (N_28663,N_26872,N_27320);
nor U28664 (N_28664,N_26904,N_26625);
nor U28665 (N_28665,N_26814,N_26877);
xor U28666 (N_28666,N_26400,N_27242);
xnor U28667 (N_28667,N_27463,N_26953);
nor U28668 (N_28668,N_27020,N_26648);
and U28669 (N_28669,N_27262,N_26850);
and U28670 (N_28670,N_27118,N_26981);
or U28671 (N_28671,N_26452,N_27147);
xnor U28672 (N_28672,N_26522,N_26668);
xnor U28673 (N_28673,N_27428,N_27114);
nor U28674 (N_28674,N_26958,N_27122);
nand U28675 (N_28675,N_27566,N_26623);
and U28676 (N_28676,N_27582,N_27493);
or U28677 (N_28677,N_26941,N_27391);
nor U28678 (N_28678,N_26771,N_26736);
nor U28679 (N_28679,N_27055,N_26530);
nor U28680 (N_28680,N_26414,N_26727);
and U28681 (N_28681,N_26551,N_26552);
nor U28682 (N_28682,N_26429,N_26617);
and U28683 (N_28683,N_27364,N_27207);
nand U28684 (N_28684,N_27123,N_27397);
nand U28685 (N_28685,N_26569,N_27167);
nor U28686 (N_28686,N_27378,N_26854);
nand U28687 (N_28687,N_26860,N_27297);
nor U28688 (N_28688,N_26423,N_26535);
nor U28689 (N_28689,N_26500,N_26878);
nand U28690 (N_28690,N_26906,N_27195);
and U28691 (N_28691,N_26651,N_26505);
and U28692 (N_28692,N_26712,N_26822);
and U28693 (N_28693,N_26917,N_27495);
nand U28694 (N_28694,N_27247,N_27130);
nand U28695 (N_28695,N_26942,N_27593);
or U28696 (N_28696,N_27178,N_26687);
xor U28697 (N_28697,N_26479,N_26887);
nand U28698 (N_28698,N_27263,N_27506);
xor U28699 (N_28699,N_27005,N_27068);
nor U28700 (N_28700,N_26959,N_27217);
nand U28701 (N_28701,N_26411,N_26507);
or U28702 (N_28702,N_26830,N_27500);
nor U28703 (N_28703,N_27349,N_27198);
xnor U28704 (N_28704,N_27563,N_26571);
nor U28705 (N_28705,N_27420,N_27417);
xnor U28706 (N_28706,N_27047,N_26608);
or U28707 (N_28707,N_27027,N_27351);
or U28708 (N_28708,N_27511,N_26984);
xor U28709 (N_28709,N_26524,N_27152);
or U28710 (N_28710,N_26607,N_27573);
or U28711 (N_28711,N_26632,N_26782);
and U28712 (N_28712,N_26619,N_27220);
or U28713 (N_28713,N_27342,N_26934);
nor U28714 (N_28714,N_26782,N_27167);
xor U28715 (N_28715,N_26722,N_26505);
nor U28716 (N_28716,N_27570,N_27342);
xnor U28717 (N_28717,N_27278,N_26880);
nor U28718 (N_28718,N_27169,N_27082);
nand U28719 (N_28719,N_26818,N_27437);
and U28720 (N_28720,N_26937,N_27299);
and U28721 (N_28721,N_27382,N_26817);
and U28722 (N_28722,N_26516,N_27279);
nor U28723 (N_28723,N_27444,N_26655);
xor U28724 (N_28724,N_27552,N_27120);
nand U28725 (N_28725,N_26624,N_26699);
and U28726 (N_28726,N_26898,N_26649);
and U28727 (N_28727,N_26914,N_26516);
nand U28728 (N_28728,N_27564,N_26799);
or U28729 (N_28729,N_27563,N_26650);
nand U28730 (N_28730,N_27261,N_26413);
or U28731 (N_28731,N_27034,N_27256);
xnor U28732 (N_28732,N_26606,N_26900);
or U28733 (N_28733,N_27556,N_26897);
and U28734 (N_28734,N_27598,N_26687);
nand U28735 (N_28735,N_27155,N_27472);
nor U28736 (N_28736,N_26476,N_27127);
nor U28737 (N_28737,N_27528,N_27582);
xnor U28738 (N_28738,N_26792,N_26956);
nor U28739 (N_28739,N_27598,N_26992);
nand U28740 (N_28740,N_27063,N_27448);
nor U28741 (N_28741,N_27384,N_27428);
xor U28742 (N_28742,N_27490,N_26989);
and U28743 (N_28743,N_27458,N_27100);
and U28744 (N_28744,N_27068,N_26723);
nor U28745 (N_28745,N_26790,N_27338);
xnor U28746 (N_28746,N_27345,N_27228);
nand U28747 (N_28747,N_26655,N_27029);
and U28748 (N_28748,N_26741,N_26825);
or U28749 (N_28749,N_27420,N_26642);
nand U28750 (N_28750,N_26495,N_26933);
nor U28751 (N_28751,N_26823,N_27442);
or U28752 (N_28752,N_26851,N_26420);
nor U28753 (N_28753,N_26668,N_26528);
xor U28754 (N_28754,N_26805,N_26677);
nand U28755 (N_28755,N_27411,N_26737);
nand U28756 (N_28756,N_26905,N_27356);
nand U28757 (N_28757,N_26921,N_26630);
xnor U28758 (N_28758,N_26575,N_26920);
xor U28759 (N_28759,N_27235,N_26475);
or U28760 (N_28760,N_26778,N_27596);
xor U28761 (N_28761,N_26512,N_27257);
and U28762 (N_28762,N_27477,N_27010);
nand U28763 (N_28763,N_27552,N_27356);
xor U28764 (N_28764,N_27071,N_26746);
nor U28765 (N_28765,N_27407,N_27488);
xor U28766 (N_28766,N_26877,N_27378);
nor U28767 (N_28767,N_27098,N_27511);
and U28768 (N_28768,N_27195,N_26888);
and U28769 (N_28769,N_27052,N_27066);
xor U28770 (N_28770,N_26567,N_27130);
and U28771 (N_28771,N_26429,N_27385);
or U28772 (N_28772,N_26795,N_26942);
nand U28773 (N_28773,N_26644,N_27343);
nor U28774 (N_28774,N_26913,N_26956);
and U28775 (N_28775,N_27063,N_26496);
nor U28776 (N_28776,N_26805,N_26646);
xnor U28777 (N_28777,N_26719,N_27219);
xnor U28778 (N_28778,N_26462,N_27589);
nor U28779 (N_28779,N_26756,N_26691);
nand U28780 (N_28780,N_27202,N_26460);
or U28781 (N_28781,N_26577,N_27124);
and U28782 (N_28782,N_26891,N_26666);
nor U28783 (N_28783,N_27059,N_27111);
xnor U28784 (N_28784,N_27450,N_27340);
and U28785 (N_28785,N_27262,N_26917);
nand U28786 (N_28786,N_27477,N_26845);
and U28787 (N_28787,N_26473,N_27120);
or U28788 (N_28788,N_26858,N_27349);
and U28789 (N_28789,N_27078,N_27127);
nor U28790 (N_28790,N_26699,N_27033);
xnor U28791 (N_28791,N_26539,N_26666);
nor U28792 (N_28792,N_27082,N_27226);
nand U28793 (N_28793,N_26552,N_26911);
nand U28794 (N_28794,N_26636,N_26750);
nand U28795 (N_28795,N_27516,N_27495);
nand U28796 (N_28796,N_27599,N_26657);
and U28797 (N_28797,N_26758,N_27361);
and U28798 (N_28798,N_27555,N_26489);
and U28799 (N_28799,N_27520,N_26437);
nor U28800 (N_28800,N_28707,N_28768);
or U28801 (N_28801,N_28152,N_28581);
nand U28802 (N_28802,N_28374,N_28305);
nand U28803 (N_28803,N_27688,N_28040);
xnor U28804 (N_28804,N_28559,N_27672);
or U28805 (N_28805,N_28447,N_27864);
nor U28806 (N_28806,N_28520,N_28051);
and U28807 (N_28807,N_28649,N_27981);
and U28808 (N_28808,N_27654,N_28295);
xnor U28809 (N_28809,N_28771,N_28551);
xor U28810 (N_28810,N_28128,N_28290);
and U28811 (N_28811,N_28036,N_28723);
or U28812 (N_28812,N_28378,N_27953);
xnor U28813 (N_28813,N_27794,N_27648);
and U28814 (N_28814,N_27686,N_28348);
xor U28815 (N_28815,N_28709,N_27644);
nor U28816 (N_28816,N_27949,N_27865);
nor U28817 (N_28817,N_28079,N_28523);
or U28818 (N_28818,N_28435,N_27921);
or U28819 (N_28819,N_28364,N_28308);
nand U28820 (N_28820,N_28176,N_28461);
nor U28821 (N_28821,N_27725,N_28773);
and U28822 (N_28822,N_28181,N_28083);
and U28823 (N_28823,N_28517,N_27886);
nor U28824 (N_28824,N_27883,N_28798);
nand U28825 (N_28825,N_28651,N_28169);
and U28826 (N_28826,N_28380,N_28656);
nand U28827 (N_28827,N_27706,N_28668);
nand U28828 (N_28828,N_28449,N_28021);
nor U28829 (N_28829,N_27992,N_27980);
and U28830 (N_28830,N_27826,N_28667);
or U28831 (N_28831,N_28714,N_27782);
or U28832 (N_28832,N_27823,N_28319);
nor U28833 (N_28833,N_28587,N_28479);
nand U28834 (N_28834,N_28238,N_28410);
nand U28835 (N_28835,N_28278,N_27964);
xor U28836 (N_28836,N_27767,N_28680);
or U28837 (N_28837,N_28172,N_28562);
nor U28838 (N_28838,N_27973,N_28757);
nand U28839 (N_28839,N_28160,N_28043);
nor U28840 (N_28840,N_28637,N_28086);
and U28841 (N_28841,N_28750,N_28538);
xor U28842 (N_28842,N_28729,N_27754);
or U28843 (N_28843,N_27803,N_27907);
nor U28844 (N_28844,N_28735,N_28426);
or U28845 (N_28845,N_27674,N_28130);
or U28846 (N_28846,N_28499,N_27784);
or U28847 (N_28847,N_28591,N_28012);
xnor U28848 (N_28848,N_27749,N_28405);
xor U28849 (N_28849,N_28475,N_28793);
and U28850 (N_28850,N_28712,N_28498);
xnor U28851 (N_28851,N_28504,N_27763);
or U28852 (N_28852,N_27918,N_28217);
and U28853 (N_28853,N_28170,N_28417);
or U28854 (N_28854,N_27951,N_28783);
nand U28855 (N_28855,N_28749,N_28700);
xor U28856 (N_28856,N_28570,N_27994);
and U28857 (N_28857,N_28147,N_28187);
and U28858 (N_28858,N_27941,N_28137);
or U28859 (N_28859,N_28360,N_28366);
and U28860 (N_28860,N_27652,N_28001);
and U28861 (N_28861,N_28020,N_28324);
and U28862 (N_28862,N_28797,N_28382);
or U28863 (N_28863,N_28014,N_27770);
nand U28864 (N_28864,N_28180,N_28407);
and U28865 (N_28865,N_28546,N_28064);
and U28866 (N_28866,N_27666,N_28791);
or U28867 (N_28867,N_28090,N_28120);
nor U28868 (N_28868,N_27824,N_28486);
or U28869 (N_28869,N_27829,N_28450);
and U28870 (N_28870,N_28560,N_28048);
or U28871 (N_28871,N_28329,N_28286);
and U28872 (N_28872,N_28124,N_27958);
nor U28873 (N_28873,N_27894,N_28034);
nor U28874 (N_28874,N_28267,N_28182);
nand U28875 (N_28875,N_27868,N_28314);
nor U28876 (N_28876,N_28639,N_27866);
or U28877 (N_28877,N_28008,N_28775);
and U28878 (N_28878,N_28646,N_27881);
xnor U28879 (N_28879,N_27861,N_27825);
nor U28880 (N_28880,N_28701,N_28478);
and U28881 (N_28881,N_28188,N_27933);
nand U28882 (N_28882,N_28521,N_28703);
nand U28883 (N_28883,N_27735,N_28101);
nand U28884 (N_28884,N_28533,N_28658);
nor U28885 (N_28885,N_27668,N_27640);
nand U28886 (N_28886,N_28430,N_27885);
nor U28887 (N_28887,N_28746,N_28483);
or U28888 (N_28888,N_27968,N_28262);
nand U28889 (N_28889,N_28606,N_28281);
nand U28890 (N_28890,N_28399,N_28782);
or U28891 (N_28891,N_27955,N_28388);
and U28892 (N_28892,N_28194,N_28753);
nor U28893 (N_28893,N_27873,N_28009);
or U28894 (N_28894,N_28670,N_27743);
xor U28895 (N_28895,N_28654,N_28662);
nor U28896 (N_28896,N_28207,N_28223);
nand U28897 (N_28897,N_28443,N_27910);
nand U28898 (N_28898,N_27764,N_28344);
or U28899 (N_28899,N_28472,N_27775);
nand U28900 (N_28900,N_28027,N_28168);
nor U28901 (N_28901,N_28556,N_28770);
or U28902 (N_28902,N_28493,N_27840);
nor U28903 (N_28903,N_27732,N_28684);
or U28904 (N_28904,N_27830,N_27675);
and U28905 (N_28905,N_28257,N_28381);
and U28906 (N_28906,N_28738,N_28744);
and U28907 (N_28907,N_27948,N_27739);
xor U28908 (N_28908,N_28069,N_28126);
xnor U28909 (N_28909,N_27766,N_28370);
nand U28910 (N_28910,N_28296,N_28565);
and U28911 (N_28911,N_27720,N_28379);
nand U28912 (N_28912,N_28492,N_28537);
and U28913 (N_28913,N_28594,N_27999);
or U28914 (N_28914,N_28589,N_28511);
nand U28915 (N_28915,N_28588,N_27729);
or U28916 (N_28916,N_28136,N_27946);
nor U28917 (N_28917,N_28583,N_28740);
and U28918 (N_28918,N_28722,N_27718);
and U28919 (N_28919,N_28448,N_28299);
and U28920 (N_28920,N_27899,N_28110);
nand U28921 (N_28921,N_28728,N_28434);
nand U28922 (N_28922,N_28607,N_28731);
xor U28923 (N_28923,N_28481,N_28352);
or U28924 (N_28924,N_28664,N_28298);
or U28925 (N_28925,N_28484,N_28681);
xor U28926 (N_28926,N_27911,N_28055);
nand U28927 (N_28927,N_27726,N_28353);
or U28928 (N_28928,N_27925,N_27962);
or U28929 (N_28929,N_28491,N_28743);
nor U28930 (N_28930,N_27621,N_28028);
nor U28931 (N_28931,N_27659,N_27902);
xor U28932 (N_28932,N_28148,N_28432);
nor U28933 (N_28933,N_27934,N_28173);
or U28934 (N_28934,N_28569,N_27699);
nor U28935 (N_28935,N_28142,N_28088);
xnor U28936 (N_28936,N_27601,N_28074);
xor U28937 (N_28937,N_28760,N_28423);
and U28938 (N_28938,N_27929,N_27613);
and U28939 (N_28939,N_28463,N_27877);
and U28940 (N_28940,N_27855,N_28165);
nand U28941 (N_28941,N_28184,N_27920);
xnor U28942 (N_28942,N_28111,N_27893);
nor U28943 (N_28943,N_28421,N_28102);
nand U28944 (N_28944,N_27664,N_28433);
and U28945 (N_28945,N_28467,N_27858);
xnor U28946 (N_28946,N_28418,N_27738);
nor U28947 (N_28947,N_28376,N_27880);
nand U28948 (N_28948,N_27611,N_28362);
and U28949 (N_28949,N_28273,N_28208);
or U28950 (N_28950,N_28711,N_28203);
and U28951 (N_28951,N_28688,N_27627);
or U28952 (N_28952,N_28230,N_27737);
nand U28953 (N_28953,N_28320,N_28186);
and U28954 (N_28954,N_27786,N_27722);
nand U28955 (N_28955,N_28078,N_27744);
or U28956 (N_28956,N_28263,N_27930);
nand U28957 (N_28957,N_28465,N_28337);
or U28958 (N_28958,N_27944,N_28297);
nor U28959 (N_28959,N_28427,N_28250);
nand U28960 (N_28960,N_27814,N_28398);
xor U28961 (N_28961,N_28420,N_28747);
nand U28962 (N_28962,N_27891,N_28500);
nand U28963 (N_28963,N_27703,N_27787);
nand U28964 (N_28964,N_28211,N_28162);
nand U28965 (N_28965,N_28516,N_28438);
and U28966 (N_28966,N_28334,N_27645);
xor U28967 (N_28967,N_28220,N_28129);
xnor U28968 (N_28968,N_27671,N_28068);
or U28969 (N_28969,N_28392,N_27745);
and U28970 (N_28970,N_28387,N_27972);
and U28971 (N_28971,N_28592,N_28039);
nor U28972 (N_28972,N_28143,N_27616);
and U28973 (N_28973,N_28026,N_28779);
nor U28974 (N_28974,N_28045,N_28748);
and U28975 (N_28975,N_28144,N_28125);
or U28976 (N_28976,N_28140,N_28494);
xor U28977 (N_28977,N_27704,N_28118);
nand U28978 (N_28978,N_28510,N_28304);
nor U28979 (N_28979,N_28132,N_28041);
nor U28980 (N_28980,N_28071,N_28601);
and U28981 (N_28981,N_28248,N_27650);
nand U28982 (N_28982,N_28185,N_28215);
or U28983 (N_28983,N_27848,N_28620);
or U28984 (N_28984,N_28752,N_28503);
and U28985 (N_28985,N_28255,N_28786);
and U28986 (N_28986,N_28199,N_28054);
xor U28987 (N_28987,N_28710,N_28761);
or U28988 (N_28988,N_27982,N_28759);
and U28989 (N_28989,N_28695,N_27607);
and U28990 (N_28990,N_28726,N_28309);
or U28991 (N_28991,N_27698,N_27638);
or U28992 (N_28992,N_28471,N_28239);
xor U28993 (N_28993,N_28233,N_27727);
nand U28994 (N_28994,N_28369,N_27959);
and U28995 (N_28995,N_28704,N_28446);
nor U28996 (N_28996,N_28291,N_27987);
nor U28997 (N_28997,N_28554,N_28650);
or U28998 (N_28998,N_27736,N_28647);
and U28999 (N_28999,N_28502,N_27758);
and U29000 (N_29000,N_28536,N_28029);
nand U29001 (N_29001,N_27690,N_28466);
or U29002 (N_29002,N_28794,N_28696);
and U29003 (N_29003,N_28609,N_28076);
nand U29004 (N_29004,N_27771,N_28628);
xor U29005 (N_29005,N_27678,N_27854);
nor U29006 (N_29006,N_27708,N_27693);
or U29007 (N_29007,N_28718,N_28346);
nand U29008 (N_29008,N_27612,N_28699);
xnor U29009 (N_29009,N_28630,N_28631);
nor U29010 (N_29010,N_28105,N_27869);
nand U29011 (N_29011,N_27832,N_28285);
xor U29012 (N_29012,N_27609,N_28529);
nand U29013 (N_29013,N_27757,N_28350);
nor U29014 (N_29014,N_28519,N_28095);
nand U29015 (N_29015,N_27935,N_28416);
nand U29016 (N_29016,N_27783,N_28052);
xor U29017 (N_29017,N_28766,N_28580);
xnor U29018 (N_29018,N_28705,N_27651);
nor U29019 (N_29019,N_28719,N_28619);
or U29020 (N_29020,N_27924,N_27903);
or U29021 (N_29021,N_28657,N_28550);
and U29022 (N_29022,N_28400,N_27998);
nand U29023 (N_29023,N_28638,N_28539);
nand U29024 (N_29024,N_28279,N_28359);
xor U29025 (N_29025,N_28512,N_27643);
nor U29026 (N_29026,N_28505,N_27660);
xor U29027 (N_29027,N_28445,N_28401);
or U29028 (N_29028,N_28103,N_28356);
or U29029 (N_29029,N_27985,N_28236);
and U29030 (N_29030,N_28383,N_27694);
xnor U29031 (N_29031,N_27884,N_27802);
xnor U29032 (N_29032,N_28013,N_28145);
or U29033 (N_29033,N_27857,N_27871);
nor U29034 (N_29034,N_28301,N_28127);
nor U29035 (N_29035,N_27807,N_28623);
and U29036 (N_29036,N_27781,N_28155);
or U29037 (N_29037,N_28397,N_28477);
or U29038 (N_29038,N_27828,N_27821);
and U29039 (N_29039,N_27939,N_27801);
nand U29040 (N_29040,N_28600,N_28146);
and U29041 (N_29041,N_27870,N_27641);
and U29042 (N_29042,N_28235,N_28063);
or U29043 (N_29043,N_28338,N_28413);
nor U29044 (N_29044,N_27842,N_28572);
and U29045 (N_29045,N_28708,N_28582);
and U29046 (N_29046,N_27836,N_28070);
nor U29047 (N_29047,N_28240,N_28098);
and U29048 (N_29048,N_28683,N_28663);
or U29049 (N_29049,N_28178,N_28189);
or U29050 (N_29050,N_28056,N_28678);
nand U29051 (N_29051,N_28157,N_27841);
nand U29052 (N_29052,N_28367,N_28283);
xnor U29053 (N_29053,N_27620,N_27760);
nor U29054 (N_29054,N_28515,N_28597);
or U29055 (N_29055,N_27966,N_28799);
or U29056 (N_29056,N_28693,N_27707);
nor U29057 (N_29057,N_27993,N_27917);
nor U29058 (N_29058,N_27755,N_27751);
and U29059 (N_29059,N_28091,N_27629);
or U29060 (N_29060,N_28489,N_28200);
nand U29061 (N_29061,N_27734,N_28228);
xor U29062 (N_29062,N_28213,N_27681);
nand U29063 (N_29063,N_28293,N_28084);
or U29064 (N_29064,N_27833,N_28122);
nand U29065 (N_29065,N_28561,N_28059);
xor U29066 (N_29066,N_28037,N_27742);
nand U29067 (N_29067,N_28694,N_28602);
xnor U29068 (N_29068,N_28153,N_27665);
nand U29069 (N_29069,N_27740,N_27882);
nor U29070 (N_29070,N_28577,N_28300);
xnor U29071 (N_29071,N_28315,N_28612);
xor U29072 (N_29072,N_27909,N_27663);
nand U29073 (N_29073,N_28439,N_28024);
nand U29074 (N_29074,N_27713,N_27752);
or U29075 (N_29075,N_27624,N_28586);
nand U29076 (N_29076,N_28534,N_27990);
and U29077 (N_29077,N_27773,N_28393);
or U29078 (N_29078,N_27682,N_28487);
nor U29079 (N_29079,N_27667,N_28357);
and U29080 (N_29080,N_28596,N_28149);
and U29081 (N_29081,N_28751,N_27761);
and U29082 (N_29082,N_28373,N_28316);
xnor U29083 (N_29083,N_28764,N_27922);
xnor U29084 (N_29084,N_28307,N_28161);
xor U29085 (N_29085,N_28047,N_28196);
nand U29086 (N_29086,N_28218,N_28287);
nand U29087 (N_29087,N_28139,N_28568);
xnor U29088 (N_29088,N_27625,N_27916);
nor U29089 (N_29089,N_28573,N_28272);
xor U29090 (N_29090,N_27662,N_27863);
or U29091 (N_29091,N_28106,N_27721);
or U29092 (N_29092,N_27965,N_27862);
nor U29093 (N_29093,N_28222,N_28336);
nor U29094 (N_29094,N_27797,N_27605);
nand U29095 (N_29095,N_28289,N_28212);
xnor U29096 (N_29096,N_28038,N_28563);
nand U29097 (N_29097,N_27875,N_28627);
and U29098 (N_29098,N_28692,N_28624);
xnor U29099 (N_29099,N_28424,N_28555);
or U29100 (N_29100,N_28115,N_28073);
nor U29101 (N_29101,N_27931,N_28642);
nor U29102 (N_29102,N_28164,N_28677);
nand U29103 (N_29103,N_27631,N_28174);
and U29104 (N_29104,N_27859,N_27628);
or U29105 (N_29105,N_27655,N_28175);
xnor U29106 (N_29106,N_28395,N_28476);
nor U29107 (N_29107,N_28535,N_28109);
nand U29108 (N_29108,N_28672,N_27691);
and U29109 (N_29109,N_28116,N_28513);
nand U29110 (N_29110,N_28330,N_28274);
and U29111 (N_29111,N_27791,N_27632);
and U29112 (N_29112,N_28190,N_28616);
nand U29113 (N_29113,N_27653,N_28632);
xor U29114 (N_29114,N_28018,N_28525);
nand U29115 (N_29115,N_28322,N_28721);
and U29116 (N_29116,N_28249,N_28574);
nand U29117 (N_29117,N_28270,N_28227);
nor U29118 (N_29118,N_28016,N_27952);
nand U29119 (N_29119,N_28774,N_28386);
xor U29120 (N_29120,N_28275,N_27850);
xnor U29121 (N_29121,N_28345,N_27793);
or U29122 (N_29122,N_27780,N_27750);
or U29123 (N_29123,N_27677,N_28062);
xor U29124 (N_29124,N_28655,N_28527);
nor U29125 (N_29125,N_28765,N_28000);
nand U29126 (N_29126,N_27701,N_28545);
nand U29127 (N_29127,N_27856,N_28035);
or U29128 (N_29128,N_28404,N_28514);
nand U29129 (N_29129,N_28112,N_28371);
xor U29130 (N_29130,N_27622,N_28326);
nand U29131 (N_29131,N_27634,N_28675);
nor U29132 (N_29132,N_28615,N_28061);
and U29133 (N_29133,N_27969,N_28659);
nor U29134 (N_29134,N_27635,N_27756);
nand U29135 (N_29135,N_28634,N_28192);
or U29136 (N_29136,N_27905,N_28745);
nand U29137 (N_29137,N_28734,N_28724);
xnor U29138 (N_29138,N_28117,N_27615);
or U29139 (N_29139,N_28384,N_27687);
xor U29140 (N_29140,N_28781,N_28626);
or U29141 (N_29141,N_28576,N_28183);
nor U29142 (N_29142,N_27642,N_28567);
nor U29143 (N_29143,N_28480,N_28727);
nor U29144 (N_29144,N_28231,N_27895);
nand U29145 (N_29145,N_28593,N_28311);
and U29146 (N_29146,N_28134,N_28614);
or U29147 (N_29147,N_28221,N_28622);
xnor U29148 (N_29148,N_27847,N_28195);
nand U29149 (N_29149,N_28225,N_27904);
nand U29150 (N_29150,N_28737,N_28795);
xnor U29151 (N_29151,N_28328,N_27996);
and U29152 (N_29152,N_27817,N_28363);
nor U29153 (N_29153,N_27845,N_27741);
and U29154 (N_29154,N_28762,N_28259);
or U29155 (N_29155,N_27974,N_28666);
nor U29156 (N_29156,N_28394,N_28097);
xnor U29157 (N_29157,N_27805,N_28406);
and U29158 (N_29158,N_28197,N_28141);
or U29159 (N_29159,N_28495,N_27816);
and U29160 (N_29160,N_28444,N_28530);
xor U29161 (N_29161,N_28389,N_28458);
or U29162 (N_29162,N_28796,N_27988);
nand U29163 (N_29163,N_28457,N_28454);
nor U29164 (N_29164,N_27696,N_28264);
nand U29165 (N_29165,N_27683,N_28201);
nor U29166 (N_29166,N_28133,N_28518);
nor U29167 (N_29167,N_28096,N_28643);
nand U29168 (N_29168,N_27827,N_28396);
nor U29169 (N_29169,N_28093,N_28772);
and U29170 (N_29170,N_28682,N_28685);
xnor U29171 (N_29171,N_28460,N_28689);
xnor U29172 (N_29172,N_28686,N_27997);
xor U29173 (N_29173,N_28099,N_28540);
nor U29174 (N_29174,N_28224,N_28604);
nand U29175 (N_29175,N_28676,N_28113);
or U29176 (N_29176,N_27804,N_28302);
or U29177 (N_29177,N_28488,N_27710);
and U29178 (N_29178,N_28261,N_27623);
nor U29179 (N_29179,N_27717,N_28590);
nor U29180 (N_29180,N_28023,N_27957);
or U29181 (N_29181,N_27788,N_28661);
or U29182 (N_29182,N_28006,N_27890);
nor U29183 (N_29183,N_28720,N_28108);
or U29184 (N_29184,N_28121,N_28635);
or U29185 (N_29185,N_28339,N_28171);
nand U29186 (N_29186,N_27617,N_27711);
and U29187 (N_29187,N_28167,N_28022);
or U29188 (N_29188,N_28010,N_28792);
or U29189 (N_29189,N_28114,N_27932);
or U29190 (N_29190,N_28002,N_28241);
and U29191 (N_29191,N_28671,N_27689);
nor U29192 (N_29192,N_28653,N_28004);
or U29193 (N_29193,N_28754,N_28506);
nor U29194 (N_29194,N_28702,N_27908);
or U29195 (N_29195,N_27619,N_28209);
nand U29196 (N_29196,N_27614,N_28033);
xor U29197 (N_29197,N_27800,N_28310);
nor U29198 (N_29198,N_28072,N_28306);
and U29199 (N_29199,N_28608,N_28542);
and U29200 (N_29200,N_27942,N_28453);
or U29201 (N_29201,N_28541,N_27927);
nor U29202 (N_29202,N_28107,N_28159);
nand U29203 (N_29203,N_28049,N_28080);
and U29204 (N_29204,N_28377,N_28082);
nand U29205 (N_29205,N_27820,N_28216);
nand U29206 (N_29206,N_28564,N_27923);
nand U29207 (N_29207,N_28713,N_27796);
and U29208 (N_29208,N_28595,N_28053);
xor U29209 (N_29209,N_27647,N_28075);
nor U29210 (N_29210,N_28578,N_28354);
or U29211 (N_29211,N_28758,N_28214);
xnor U29212 (N_29212,N_28468,N_27971);
or U29213 (N_29213,N_27940,N_28733);
and U29214 (N_29214,N_28077,N_27600);
nand U29215 (N_29215,N_27810,N_28509);
and U29216 (N_29216,N_28408,N_28464);
xor U29217 (N_29217,N_28019,N_28790);
and U29218 (N_29218,N_28532,N_27731);
nand U29219 (N_29219,N_28585,N_27851);
and U29220 (N_29220,N_27785,N_27849);
or U29221 (N_29221,N_28349,N_27733);
and U29222 (N_29222,N_27919,N_28015);
and U29223 (N_29223,N_28251,N_27938);
or U29224 (N_29224,N_28046,N_27768);
and U29225 (N_29225,N_28252,N_28253);
xor U29226 (N_29226,N_28332,N_27913);
or U29227 (N_29227,N_28003,N_28469);
nor U29228 (N_29228,N_28697,N_28361);
and U29229 (N_29229,N_28456,N_27879);
and U29230 (N_29230,N_28007,N_28042);
nand U29231 (N_29231,N_28229,N_28769);
and U29232 (N_29232,N_28621,N_27852);
or U29233 (N_29233,N_28245,N_28548);
or U29234 (N_29234,N_28507,N_27936);
and U29235 (N_29235,N_27956,N_27748);
nand U29236 (N_29236,N_28531,N_28092);
and U29237 (N_29237,N_28219,N_28060);
nand U29238 (N_29238,N_28579,N_28232);
nand U29239 (N_29239,N_28280,N_28292);
nor U29240 (N_29240,N_28549,N_27986);
or U29241 (N_29241,N_28473,N_27692);
and U29242 (N_29242,N_28156,N_27837);
nor U29243 (N_29243,N_27639,N_28044);
and U29244 (N_29244,N_28005,N_28558);
nand U29245 (N_29245,N_28603,N_27716);
or U29246 (N_29246,N_28206,N_28669);
nand U29247 (N_29247,N_28584,N_28725);
xnor U29248 (N_29248,N_27937,N_28763);
xnor U29249 (N_29249,N_27657,N_27661);
and U29250 (N_29250,N_28690,N_28778);
or U29251 (N_29251,N_28266,N_28254);
nor U29252 (N_29252,N_27945,N_28025);
nor U29253 (N_29253,N_28547,N_27777);
xnor U29254 (N_29254,N_28409,N_28422);
nand U29255 (N_29255,N_28412,N_28347);
xor U29256 (N_29256,N_28459,N_28193);
nor U29257 (N_29257,N_28415,N_28303);
nand U29258 (N_29258,N_28462,N_27778);
and U29259 (N_29259,N_28429,N_27977);
nor U29260 (N_29260,N_28321,N_27790);
nor U29261 (N_29261,N_28313,N_28202);
nand U29262 (N_29262,N_28665,N_28276);
xor U29263 (N_29263,N_28644,N_28179);
nand U29264 (N_29264,N_28566,N_28526);
or U29265 (N_29265,N_27702,N_28247);
nor U29266 (N_29266,N_27960,N_28605);
xor U29267 (N_29267,N_28081,N_28094);
nor U29268 (N_29268,N_27914,N_28431);
nor U29269 (N_29269,N_28428,N_28150);
and U29270 (N_29270,N_28066,N_28244);
nor U29271 (N_29271,N_28440,N_28246);
or U29272 (N_29272,N_28104,N_27878);
nand U29273 (N_29273,N_27602,N_27943);
and U29274 (N_29274,N_27912,N_28123);
xnor U29275 (N_29275,N_27896,N_27714);
and U29276 (N_29276,N_28441,N_28451);
or U29277 (N_29277,N_28191,N_27926);
xnor U29278 (N_29278,N_28340,N_28177);
nor U29279 (N_29279,N_28617,N_27928);
nand U29280 (N_29280,N_28598,N_28557);
and U29281 (N_29281,N_28355,N_28335);
or U29282 (N_29282,N_28645,N_27844);
nor U29283 (N_29283,N_28327,N_27806);
or U29284 (N_29284,N_28470,N_27715);
nor U29285 (N_29285,N_28755,N_28282);
or U29286 (N_29286,N_28636,N_28089);
nor U29287 (N_29287,N_27915,N_28312);
xor U29288 (N_29288,N_27961,N_27947);
and U29289 (N_29289,N_28365,N_28402);
and U29290 (N_29290,N_28673,N_27892);
xor U29291 (N_29291,N_27676,N_28788);
nor U29292 (N_29292,N_28625,N_27670);
and U29293 (N_29293,N_27818,N_28776);
xnor U29294 (N_29294,N_28524,N_27963);
and U29295 (N_29295,N_28085,N_28343);
or U29296 (N_29296,N_28151,N_28785);
xnor U29297 (N_29297,N_28030,N_28732);
nor U29298 (N_29298,N_28698,N_28419);
or U29299 (N_29299,N_27889,N_28501);
nand U29300 (N_29300,N_27989,N_28391);
xnor U29301 (N_29301,N_28633,N_27637);
xnor U29302 (N_29302,N_28411,N_28767);
and U29303 (N_29303,N_28571,N_27728);
or U29304 (N_29304,N_27658,N_27809);
nand U29305 (N_29305,N_28242,N_28256);
nor U29306 (N_29306,N_28260,N_27712);
xor U29307 (N_29307,N_28351,N_28318);
nor U29308 (N_29308,N_27815,N_27603);
nand U29309 (N_29309,N_28067,N_27636);
xor U29310 (N_29310,N_28660,N_27970);
nand U29311 (N_29311,N_28135,N_27779);
and U29312 (N_29312,N_28425,N_28717);
and U29313 (N_29313,N_28553,N_27606);
nand U29314 (N_29314,N_28618,N_28648);
nor U29315 (N_29315,N_27610,N_27705);
nand U29316 (N_29316,N_27834,N_27684);
and U29317 (N_29317,N_28375,N_28131);
xor U29318 (N_29318,N_27774,N_27906);
and U29319 (N_29319,N_28730,N_28323);
xor U29320 (N_29320,N_27872,N_27604);
xnor U29321 (N_29321,N_28269,N_27630);
or U29322 (N_29322,N_27901,N_28204);
or U29323 (N_29323,N_28265,N_27843);
or U29324 (N_29324,N_28575,N_27976);
and U29325 (N_29325,N_28496,N_27975);
and U29326 (N_29326,N_27765,N_28237);
and U29327 (N_29327,N_27979,N_27789);
and U29328 (N_29328,N_27633,N_28100);
nand U29329 (N_29329,N_28599,N_27876);
nand U29330 (N_29330,N_28497,N_28358);
nor U29331 (N_29331,N_27798,N_28528);
xor U29332 (N_29332,N_28784,N_27888);
or U29333 (N_29333,N_27991,N_27673);
and U29334 (N_29334,N_27795,N_27983);
nor U29335 (N_29335,N_27769,N_28342);
xnor U29336 (N_29336,N_27867,N_27618);
and U29337 (N_29337,N_28706,N_28317);
and U29338 (N_29338,N_27900,N_27799);
and U29339 (N_29339,N_28158,N_28031);
xor U29340 (N_29340,N_28119,N_28271);
nand U29341 (N_29341,N_28437,N_27608);
and U29342 (N_29342,N_27759,N_28777);
or U29343 (N_29343,N_27709,N_27950);
xnor U29344 (N_29344,N_27719,N_27831);
nor U29345 (N_29345,N_28436,N_27838);
nor U29346 (N_29346,N_28032,N_28277);
xnor U29347 (N_29347,N_28687,N_27753);
or U29348 (N_29348,N_27649,N_27679);
nand U29349 (N_29349,N_28368,N_28742);
nor U29350 (N_29350,N_28163,N_28787);
nor U29351 (N_29351,N_28715,N_27724);
xnor U29352 (N_29352,N_27697,N_27874);
or U29353 (N_29353,N_27839,N_27792);
nand U29354 (N_29354,N_28325,N_28210);
or U29355 (N_29355,N_28294,N_27853);
nor U29356 (N_29356,N_28234,N_27897);
xor U29357 (N_29357,N_28610,N_28268);
xnor U29358 (N_29358,N_28205,N_28508);
or U29359 (N_29359,N_28455,N_27978);
and U29360 (N_29360,N_27898,N_28243);
nor U29361 (N_29361,N_27772,N_27819);
and U29362 (N_29362,N_28611,N_28679);
or U29363 (N_29363,N_28691,N_27626);
and U29364 (N_29364,N_28741,N_27746);
nor U29365 (N_29365,N_27812,N_28403);
nand U29366 (N_29366,N_28258,N_28017);
nor U29367 (N_29367,N_27776,N_27846);
nand U29368 (N_29368,N_27984,N_27656);
and U29369 (N_29369,N_27954,N_28442);
nor U29370 (N_29370,N_28485,N_28138);
nand U29371 (N_29371,N_28166,N_28736);
xnor U29372 (N_29372,N_28640,N_27730);
xnor U29373 (N_29373,N_27700,N_28198);
nand U29374 (N_29374,N_27762,N_28629);
xnor U29375 (N_29375,N_28490,N_28414);
xor U29376 (N_29376,N_28789,N_28543);
or U29377 (N_29377,N_28641,N_28522);
or U29378 (N_29378,N_28087,N_27835);
xor U29379 (N_29379,N_27669,N_28780);
or U29380 (N_29380,N_28739,N_27967);
nor U29381 (N_29381,N_28674,N_28552);
nor U29382 (N_29382,N_28390,N_27822);
nor U29383 (N_29383,N_28011,N_27685);
nand U29384 (N_29384,N_27860,N_28065);
xor U29385 (N_29385,N_28154,N_28050);
nand U29386 (N_29386,N_27723,N_27695);
or U29387 (N_29387,N_28284,N_27811);
or U29388 (N_29388,N_28057,N_27813);
xor U29389 (N_29389,N_28613,N_28474);
xor U29390 (N_29390,N_28226,N_28341);
or U29391 (N_29391,N_28372,N_28058);
nand U29392 (N_29392,N_27747,N_28333);
xor U29393 (N_29393,N_28331,N_27646);
and U29394 (N_29394,N_28482,N_28544);
and U29395 (N_29395,N_27995,N_28716);
nor U29396 (N_29396,N_27680,N_28756);
xor U29397 (N_29397,N_28288,N_27887);
nand U29398 (N_29398,N_28452,N_28652);
nand U29399 (N_29399,N_28385,N_27808);
nor U29400 (N_29400,N_28722,N_28224);
and U29401 (N_29401,N_27601,N_27777);
nand U29402 (N_29402,N_27847,N_28607);
nor U29403 (N_29403,N_28252,N_27671);
nand U29404 (N_29404,N_28128,N_27792);
nand U29405 (N_29405,N_27928,N_27777);
nand U29406 (N_29406,N_28620,N_28402);
xor U29407 (N_29407,N_28650,N_28603);
xor U29408 (N_29408,N_28440,N_28512);
nor U29409 (N_29409,N_27890,N_28415);
nand U29410 (N_29410,N_27943,N_28526);
nand U29411 (N_29411,N_28238,N_27881);
or U29412 (N_29412,N_28527,N_28411);
nand U29413 (N_29413,N_27721,N_28244);
and U29414 (N_29414,N_28556,N_28718);
or U29415 (N_29415,N_28403,N_28333);
and U29416 (N_29416,N_27687,N_27983);
or U29417 (N_29417,N_28053,N_28277);
or U29418 (N_29418,N_28376,N_28512);
nand U29419 (N_29419,N_27997,N_27963);
nor U29420 (N_29420,N_28142,N_27731);
nor U29421 (N_29421,N_28099,N_28596);
or U29422 (N_29422,N_27901,N_28069);
xor U29423 (N_29423,N_27779,N_28102);
xor U29424 (N_29424,N_27989,N_28776);
nor U29425 (N_29425,N_28483,N_28112);
or U29426 (N_29426,N_28551,N_28474);
or U29427 (N_29427,N_28568,N_28235);
xor U29428 (N_29428,N_28799,N_27887);
nor U29429 (N_29429,N_27858,N_27995);
xor U29430 (N_29430,N_27890,N_27843);
nor U29431 (N_29431,N_27999,N_28798);
or U29432 (N_29432,N_27638,N_28034);
or U29433 (N_29433,N_27781,N_28786);
xnor U29434 (N_29434,N_28214,N_27804);
xnor U29435 (N_29435,N_27669,N_28560);
or U29436 (N_29436,N_28388,N_28238);
and U29437 (N_29437,N_28309,N_28369);
and U29438 (N_29438,N_27652,N_28743);
or U29439 (N_29439,N_28154,N_27686);
xor U29440 (N_29440,N_27866,N_28147);
or U29441 (N_29441,N_28052,N_28636);
nand U29442 (N_29442,N_27965,N_28672);
or U29443 (N_29443,N_28331,N_27716);
and U29444 (N_29444,N_27639,N_28410);
nor U29445 (N_29445,N_27953,N_28297);
or U29446 (N_29446,N_27639,N_28476);
or U29447 (N_29447,N_28440,N_28411);
and U29448 (N_29448,N_28737,N_27983);
xnor U29449 (N_29449,N_28073,N_27691);
nor U29450 (N_29450,N_27739,N_28384);
nor U29451 (N_29451,N_27934,N_28690);
and U29452 (N_29452,N_27939,N_27892);
xnor U29453 (N_29453,N_28227,N_28398);
nor U29454 (N_29454,N_27820,N_28761);
nand U29455 (N_29455,N_28428,N_28661);
nand U29456 (N_29456,N_28767,N_28362);
nand U29457 (N_29457,N_27787,N_28714);
and U29458 (N_29458,N_27999,N_28024);
and U29459 (N_29459,N_27726,N_28070);
xor U29460 (N_29460,N_27673,N_28262);
or U29461 (N_29461,N_28628,N_28119);
xor U29462 (N_29462,N_27679,N_28362);
nand U29463 (N_29463,N_27955,N_28115);
nand U29464 (N_29464,N_28216,N_27790);
nand U29465 (N_29465,N_28329,N_27639);
nor U29466 (N_29466,N_27722,N_28658);
xnor U29467 (N_29467,N_27788,N_28012);
nor U29468 (N_29468,N_28143,N_28642);
or U29469 (N_29469,N_28380,N_28554);
nand U29470 (N_29470,N_28669,N_28135);
nor U29471 (N_29471,N_28630,N_28394);
xnor U29472 (N_29472,N_28034,N_28065);
nand U29473 (N_29473,N_27641,N_27826);
and U29474 (N_29474,N_28670,N_27619);
or U29475 (N_29475,N_28714,N_28169);
or U29476 (N_29476,N_27825,N_28108);
xor U29477 (N_29477,N_28549,N_28350);
and U29478 (N_29478,N_27673,N_27839);
nor U29479 (N_29479,N_27719,N_28138);
or U29480 (N_29480,N_27844,N_27602);
and U29481 (N_29481,N_28548,N_27750);
and U29482 (N_29482,N_28456,N_28720);
or U29483 (N_29483,N_27760,N_28628);
nand U29484 (N_29484,N_27694,N_27640);
nor U29485 (N_29485,N_28541,N_28152);
nor U29486 (N_29486,N_28503,N_28222);
and U29487 (N_29487,N_28217,N_27629);
xor U29488 (N_29488,N_28102,N_28532);
and U29489 (N_29489,N_28731,N_28554);
or U29490 (N_29490,N_27799,N_27767);
nor U29491 (N_29491,N_27764,N_27774);
xnor U29492 (N_29492,N_28024,N_28548);
xnor U29493 (N_29493,N_28319,N_27700);
xnor U29494 (N_29494,N_27933,N_27675);
xnor U29495 (N_29495,N_27687,N_28291);
xor U29496 (N_29496,N_28581,N_27848);
or U29497 (N_29497,N_28025,N_28776);
or U29498 (N_29498,N_27734,N_28793);
xnor U29499 (N_29499,N_27734,N_28380);
xnor U29500 (N_29500,N_27814,N_28393);
and U29501 (N_29501,N_28111,N_28581);
and U29502 (N_29502,N_27868,N_27640);
nand U29503 (N_29503,N_27717,N_28178);
xor U29504 (N_29504,N_27991,N_28274);
or U29505 (N_29505,N_28504,N_28473);
xnor U29506 (N_29506,N_27722,N_27605);
or U29507 (N_29507,N_28735,N_27921);
or U29508 (N_29508,N_28220,N_27632);
nand U29509 (N_29509,N_28365,N_28265);
nor U29510 (N_29510,N_28470,N_27901);
xor U29511 (N_29511,N_28771,N_27974);
xnor U29512 (N_29512,N_28697,N_27803);
nor U29513 (N_29513,N_28391,N_27844);
xnor U29514 (N_29514,N_28452,N_28325);
and U29515 (N_29515,N_27987,N_28521);
nor U29516 (N_29516,N_28306,N_28780);
and U29517 (N_29517,N_28127,N_28439);
or U29518 (N_29518,N_27611,N_27636);
nor U29519 (N_29519,N_28007,N_27685);
and U29520 (N_29520,N_27603,N_28161);
nand U29521 (N_29521,N_27875,N_28189);
and U29522 (N_29522,N_28657,N_27892);
xnor U29523 (N_29523,N_28586,N_28785);
xor U29524 (N_29524,N_28342,N_28701);
xnor U29525 (N_29525,N_28548,N_27798);
nand U29526 (N_29526,N_27906,N_28360);
nor U29527 (N_29527,N_28032,N_28417);
nor U29528 (N_29528,N_27852,N_28749);
nand U29529 (N_29529,N_27738,N_28627);
or U29530 (N_29530,N_28396,N_28254);
xor U29531 (N_29531,N_27930,N_27719);
nor U29532 (N_29532,N_27958,N_28142);
nand U29533 (N_29533,N_27654,N_28042);
or U29534 (N_29534,N_28534,N_28407);
xnor U29535 (N_29535,N_27835,N_28400);
and U29536 (N_29536,N_28609,N_28224);
nor U29537 (N_29537,N_28568,N_28273);
nor U29538 (N_29538,N_28419,N_28477);
or U29539 (N_29539,N_28469,N_28795);
and U29540 (N_29540,N_28479,N_28244);
nand U29541 (N_29541,N_28218,N_28308);
xnor U29542 (N_29542,N_27710,N_28193);
or U29543 (N_29543,N_27846,N_28484);
xor U29544 (N_29544,N_28209,N_27606);
or U29545 (N_29545,N_28174,N_27888);
and U29546 (N_29546,N_28124,N_27844);
and U29547 (N_29547,N_28405,N_28755);
or U29548 (N_29548,N_28734,N_27914);
nor U29549 (N_29549,N_28232,N_28482);
nand U29550 (N_29550,N_28585,N_28263);
or U29551 (N_29551,N_28091,N_28267);
nor U29552 (N_29552,N_27910,N_28003);
or U29553 (N_29553,N_27863,N_28765);
or U29554 (N_29554,N_28061,N_28323);
xnor U29555 (N_29555,N_27946,N_28442);
and U29556 (N_29556,N_28546,N_28764);
or U29557 (N_29557,N_28146,N_28018);
or U29558 (N_29558,N_27997,N_27606);
xor U29559 (N_29559,N_28117,N_27723);
or U29560 (N_29560,N_27999,N_28395);
and U29561 (N_29561,N_28259,N_28755);
nor U29562 (N_29562,N_28165,N_28148);
xnor U29563 (N_29563,N_28247,N_28049);
and U29564 (N_29564,N_28581,N_28585);
xnor U29565 (N_29565,N_28375,N_28735);
nand U29566 (N_29566,N_28757,N_27971);
or U29567 (N_29567,N_28475,N_28129);
nand U29568 (N_29568,N_28147,N_27785);
or U29569 (N_29569,N_28154,N_28100);
or U29570 (N_29570,N_27804,N_28720);
and U29571 (N_29571,N_28260,N_27871);
nand U29572 (N_29572,N_28596,N_28256);
nand U29573 (N_29573,N_27737,N_27942);
xor U29574 (N_29574,N_28066,N_27961);
or U29575 (N_29575,N_28600,N_28346);
and U29576 (N_29576,N_28239,N_28332);
or U29577 (N_29577,N_28247,N_27859);
nand U29578 (N_29578,N_28733,N_27909);
xnor U29579 (N_29579,N_28058,N_28289);
nor U29580 (N_29580,N_28178,N_28439);
nand U29581 (N_29581,N_28179,N_28342);
nor U29582 (N_29582,N_27983,N_28266);
nor U29583 (N_29583,N_28029,N_28614);
nor U29584 (N_29584,N_28181,N_28681);
and U29585 (N_29585,N_27944,N_28309);
nand U29586 (N_29586,N_28106,N_28486);
xnor U29587 (N_29587,N_28058,N_28127);
nand U29588 (N_29588,N_28638,N_28486);
xnor U29589 (N_29589,N_28475,N_27859);
nand U29590 (N_29590,N_28411,N_27755);
nand U29591 (N_29591,N_27795,N_28485);
nand U29592 (N_29592,N_28344,N_27867);
nand U29593 (N_29593,N_27940,N_27823);
and U29594 (N_29594,N_27956,N_28150);
or U29595 (N_29595,N_28712,N_28562);
nor U29596 (N_29596,N_28100,N_28231);
xnor U29597 (N_29597,N_28197,N_27793);
nor U29598 (N_29598,N_27726,N_27602);
or U29599 (N_29599,N_27993,N_28415);
nand U29600 (N_29600,N_28382,N_28024);
or U29601 (N_29601,N_28200,N_28468);
and U29602 (N_29602,N_28541,N_28123);
or U29603 (N_29603,N_28491,N_28597);
nand U29604 (N_29604,N_27603,N_28568);
and U29605 (N_29605,N_28254,N_28674);
and U29606 (N_29606,N_28073,N_28796);
nor U29607 (N_29607,N_28303,N_28006);
nand U29608 (N_29608,N_27747,N_28492);
nand U29609 (N_29609,N_28171,N_27856);
nand U29610 (N_29610,N_27601,N_27730);
xnor U29611 (N_29611,N_27847,N_28417);
and U29612 (N_29612,N_27750,N_28286);
xor U29613 (N_29613,N_27819,N_28248);
nand U29614 (N_29614,N_28640,N_28185);
xnor U29615 (N_29615,N_27682,N_28654);
and U29616 (N_29616,N_28787,N_28611);
nor U29617 (N_29617,N_28491,N_27715);
nor U29618 (N_29618,N_28642,N_28104);
nor U29619 (N_29619,N_28291,N_28355);
or U29620 (N_29620,N_28600,N_28151);
xor U29621 (N_29621,N_27904,N_28375);
xor U29622 (N_29622,N_28335,N_27997);
nor U29623 (N_29623,N_28620,N_28062);
nor U29624 (N_29624,N_28248,N_28367);
nor U29625 (N_29625,N_27601,N_28538);
nor U29626 (N_29626,N_28172,N_28270);
xnor U29627 (N_29627,N_28182,N_27899);
and U29628 (N_29628,N_28458,N_28519);
and U29629 (N_29629,N_28761,N_28348);
or U29630 (N_29630,N_28557,N_28036);
nor U29631 (N_29631,N_28397,N_28239);
and U29632 (N_29632,N_28597,N_28573);
nor U29633 (N_29633,N_28213,N_28598);
xor U29634 (N_29634,N_28218,N_28516);
or U29635 (N_29635,N_28769,N_28234);
xnor U29636 (N_29636,N_28711,N_28373);
nor U29637 (N_29637,N_27748,N_27712);
or U29638 (N_29638,N_28630,N_28497);
xor U29639 (N_29639,N_27801,N_28010);
nor U29640 (N_29640,N_28242,N_28364);
or U29641 (N_29641,N_28570,N_27857);
nor U29642 (N_29642,N_28711,N_28450);
and U29643 (N_29643,N_28262,N_28591);
or U29644 (N_29644,N_28724,N_28177);
xnor U29645 (N_29645,N_28619,N_28474);
and U29646 (N_29646,N_28747,N_27951);
xnor U29647 (N_29647,N_27916,N_28407);
and U29648 (N_29648,N_28170,N_28283);
nor U29649 (N_29649,N_28017,N_28365);
xnor U29650 (N_29650,N_27769,N_28151);
or U29651 (N_29651,N_28282,N_27710);
and U29652 (N_29652,N_28282,N_28576);
nand U29653 (N_29653,N_27988,N_27738);
or U29654 (N_29654,N_28037,N_28393);
and U29655 (N_29655,N_28662,N_28238);
xnor U29656 (N_29656,N_27751,N_27984);
nor U29657 (N_29657,N_28532,N_28602);
nand U29658 (N_29658,N_27924,N_28704);
nand U29659 (N_29659,N_28422,N_28651);
and U29660 (N_29660,N_28587,N_28156);
xor U29661 (N_29661,N_27882,N_28480);
xor U29662 (N_29662,N_28173,N_28527);
xnor U29663 (N_29663,N_28373,N_27602);
or U29664 (N_29664,N_28439,N_28175);
or U29665 (N_29665,N_27688,N_27797);
nand U29666 (N_29666,N_27640,N_28606);
nand U29667 (N_29667,N_27774,N_28264);
nor U29668 (N_29668,N_28010,N_27968);
nor U29669 (N_29669,N_28000,N_28045);
nor U29670 (N_29670,N_27786,N_28008);
or U29671 (N_29671,N_27921,N_28480);
xor U29672 (N_29672,N_27787,N_27685);
and U29673 (N_29673,N_27784,N_28113);
or U29674 (N_29674,N_28447,N_28588);
nand U29675 (N_29675,N_28038,N_28640);
and U29676 (N_29676,N_28457,N_27995);
nand U29677 (N_29677,N_27796,N_27953);
or U29678 (N_29678,N_28196,N_27862);
or U29679 (N_29679,N_28042,N_28178);
or U29680 (N_29680,N_27662,N_27982);
nor U29681 (N_29681,N_28653,N_27913);
nor U29682 (N_29682,N_28134,N_28776);
nor U29683 (N_29683,N_28265,N_28430);
nor U29684 (N_29684,N_28050,N_27658);
xor U29685 (N_29685,N_27620,N_28024);
nor U29686 (N_29686,N_28171,N_28479);
and U29687 (N_29687,N_28321,N_28341);
nand U29688 (N_29688,N_28340,N_27893);
nor U29689 (N_29689,N_27990,N_28343);
or U29690 (N_29690,N_28443,N_28056);
xnor U29691 (N_29691,N_28716,N_27802);
and U29692 (N_29692,N_27803,N_27615);
nor U29693 (N_29693,N_27689,N_28602);
xor U29694 (N_29694,N_28731,N_28128);
nor U29695 (N_29695,N_28051,N_27638);
or U29696 (N_29696,N_28026,N_28769);
xor U29697 (N_29697,N_27649,N_28320);
xor U29698 (N_29698,N_28112,N_28634);
or U29699 (N_29699,N_28029,N_28183);
xor U29700 (N_29700,N_27704,N_27698);
xnor U29701 (N_29701,N_27849,N_28250);
nor U29702 (N_29702,N_28111,N_28084);
nand U29703 (N_29703,N_28692,N_27930);
xor U29704 (N_29704,N_27925,N_28020);
nand U29705 (N_29705,N_28444,N_27946);
nor U29706 (N_29706,N_27741,N_27806);
nand U29707 (N_29707,N_28072,N_28523);
xnor U29708 (N_29708,N_27763,N_28621);
nand U29709 (N_29709,N_28505,N_28123);
nor U29710 (N_29710,N_28796,N_28382);
and U29711 (N_29711,N_27617,N_27830);
and U29712 (N_29712,N_27950,N_28145);
xor U29713 (N_29713,N_27733,N_28631);
xnor U29714 (N_29714,N_28726,N_27926);
nand U29715 (N_29715,N_28217,N_28505);
nor U29716 (N_29716,N_27689,N_27868);
xor U29717 (N_29717,N_28225,N_28679);
and U29718 (N_29718,N_27986,N_28504);
nor U29719 (N_29719,N_28522,N_27673);
or U29720 (N_29720,N_28747,N_28011);
nand U29721 (N_29721,N_28400,N_27842);
nand U29722 (N_29722,N_28331,N_28195);
nand U29723 (N_29723,N_27648,N_28285);
and U29724 (N_29724,N_28625,N_28093);
xor U29725 (N_29725,N_27699,N_27767);
nand U29726 (N_29726,N_28308,N_27734);
nor U29727 (N_29727,N_28223,N_28639);
nand U29728 (N_29728,N_28736,N_28023);
or U29729 (N_29729,N_28317,N_28537);
or U29730 (N_29730,N_27893,N_28710);
and U29731 (N_29731,N_28316,N_28656);
nand U29732 (N_29732,N_28718,N_28419);
and U29733 (N_29733,N_28404,N_27859);
nor U29734 (N_29734,N_27621,N_28793);
nor U29735 (N_29735,N_28581,N_28258);
or U29736 (N_29736,N_27929,N_28400);
or U29737 (N_29737,N_28365,N_28035);
nor U29738 (N_29738,N_28092,N_28716);
xnor U29739 (N_29739,N_27630,N_27732);
nand U29740 (N_29740,N_27761,N_27958);
xor U29741 (N_29741,N_28590,N_27890);
nand U29742 (N_29742,N_27968,N_27906);
nor U29743 (N_29743,N_27897,N_27979);
xnor U29744 (N_29744,N_28300,N_27961);
nand U29745 (N_29745,N_27820,N_28014);
xor U29746 (N_29746,N_28166,N_28313);
xnor U29747 (N_29747,N_28441,N_28220);
or U29748 (N_29748,N_28365,N_28514);
nand U29749 (N_29749,N_28271,N_27858);
or U29750 (N_29750,N_27863,N_28298);
nand U29751 (N_29751,N_28510,N_27687);
and U29752 (N_29752,N_27700,N_28741);
xor U29753 (N_29753,N_28225,N_27747);
nand U29754 (N_29754,N_28635,N_28427);
nor U29755 (N_29755,N_28290,N_27688);
and U29756 (N_29756,N_28522,N_28772);
or U29757 (N_29757,N_27895,N_28627);
nand U29758 (N_29758,N_28474,N_27603);
and U29759 (N_29759,N_28121,N_28325);
nand U29760 (N_29760,N_27981,N_28681);
xor U29761 (N_29761,N_28703,N_28283);
xnor U29762 (N_29762,N_28746,N_27692);
or U29763 (N_29763,N_28601,N_28659);
xnor U29764 (N_29764,N_28349,N_28079);
and U29765 (N_29765,N_28663,N_27600);
nor U29766 (N_29766,N_28534,N_28377);
xnor U29767 (N_29767,N_27849,N_28710);
or U29768 (N_29768,N_28662,N_28094);
and U29769 (N_29769,N_28513,N_28409);
xnor U29770 (N_29770,N_27940,N_27886);
nand U29771 (N_29771,N_28519,N_28115);
and U29772 (N_29772,N_28736,N_28419);
or U29773 (N_29773,N_28451,N_27614);
nor U29774 (N_29774,N_28542,N_28370);
and U29775 (N_29775,N_28589,N_28548);
nor U29776 (N_29776,N_28560,N_28686);
or U29777 (N_29777,N_27903,N_28529);
or U29778 (N_29778,N_27861,N_28043);
and U29779 (N_29779,N_27992,N_27785);
nor U29780 (N_29780,N_28248,N_28111);
nor U29781 (N_29781,N_27831,N_28534);
nand U29782 (N_29782,N_27980,N_28280);
xnor U29783 (N_29783,N_28504,N_28530);
nor U29784 (N_29784,N_28546,N_28249);
xnor U29785 (N_29785,N_28046,N_27821);
xnor U29786 (N_29786,N_27805,N_28298);
nand U29787 (N_29787,N_28166,N_28522);
nand U29788 (N_29788,N_28259,N_28340);
and U29789 (N_29789,N_28725,N_27614);
nand U29790 (N_29790,N_28536,N_28619);
and U29791 (N_29791,N_28478,N_27953);
and U29792 (N_29792,N_28367,N_27679);
or U29793 (N_29793,N_28501,N_28213);
nand U29794 (N_29794,N_27935,N_28730);
nor U29795 (N_29795,N_28579,N_28089);
nand U29796 (N_29796,N_28248,N_28016);
and U29797 (N_29797,N_28073,N_28501);
nor U29798 (N_29798,N_28705,N_27762);
or U29799 (N_29799,N_28034,N_27671);
and U29800 (N_29800,N_28122,N_27778);
nand U29801 (N_29801,N_28146,N_27832);
and U29802 (N_29802,N_28095,N_28588);
and U29803 (N_29803,N_27878,N_27849);
or U29804 (N_29804,N_27870,N_27634);
nand U29805 (N_29805,N_27652,N_27639);
xnor U29806 (N_29806,N_27677,N_28410);
and U29807 (N_29807,N_28525,N_28707);
xnor U29808 (N_29808,N_28786,N_28629);
xnor U29809 (N_29809,N_28106,N_27785);
nor U29810 (N_29810,N_28056,N_28354);
nor U29811 (N_29811,N_27851,N_28584);
and U29812 (N_29812,N_28741,N_28440);
xor U29813 (N_29813,N_28352,N_27821);
or U29814 (N_29814,N_28733,N_28102);
and U29815 (N_29815,N_28755,N_28280);
xor U29816 (N_29816,N_27862,N_28004);
or U29817 (N_29817,N_28751,N_28757);
nor U29818 (N_29818,N_28106,N_28179);
xor U29819 (N_29819,N_28225,N_28492);
nor U29820 (N_29820,N_27881,N_28367);
or U29821 (N_29821,N_28196,N_28148);
and U29822 (N_29822,N_27695,N_27911);
and U29823 (N_29823,N_27932,N_28420);
nand U29824 (N_29824,N_27902,N_28166);
xnor U29825 (N_29825,N_28029,N_28074);
xor U29826 (N_29826,N_28163,N_27703);
and U29827 (N_29827,N_27768,N_28202);
nand U29828 (N_29828,N_27694,N_28204);
xor U29829 (N_29829,N_28074,N_28730);
or U29830 (N_29830,N_28393,N_27739);
nor U29831 (N_29831,N_28009,N_28611);
or U29832 (N_29832,N_28408,N_28452);
and U29833 (N_29833,N_28422,N_28390);
nor U29834 (N_29834,N_28387,N_28544);
nand U29835 (N_29835,N_27965,N_27880);
xor U29836 (N_29836,N_28686,N_28708);
nor U29837 (N_29837,N_27993,N_28229);
or U29838 (N_29838,N_28340,N_28653);
and U29839 (N_29839,N_28709,N_28656);
nand U29840 (N_29840,N_28392,N_28316);
nor U29841 (N_29841,N_27944,N_28399);
nor U29842 (N_29842,N_27822,N_28763);
and U29843 (N_29843,N_28757,N_28464);
or U29844 (N_29844,N_28506,N_27660);
xor U29845 (N_29845,N_28048,N_28368);
or U29846 (N_29846,N_27687,N_28260);
and U29847 (N_29847,N_28095,N_28401);
nand U29848 (N_29848,N_27855,N_28573);
and U29849 (N_29849,N_28648,N_28727);
xor U29850 (N_29850,N_28785,N_27814);
nand U29851 (N_29851,N_28103,N_27660);
and U29852 (N_29852,N_28014,N_28302);
or U29853 (N_29853,N_28153,N_27728);
nor U29854 (N_29854,N_28492,N_27652);
nor U29855 (N_29855,N_27990,N_27799);
nand U29856 (N_29856,N_27958,N_28423);
nor U29857 (N_29857,N_27708,N_28476);
or U29858 (N_29858,N_28147,N_28785);
nand U29859 (N_29859,N_28771,N_28155);
xor U29860 (N_29860,N_27752,N_27957);
xnor U29861 (N_29861,N_28216,N_27989);
or U29862 (N_29862,N_28175,N_27928);
xnor U29863 (N_29863,N_28294,N_28589);
xor U29864 (N_29864,N_27622,N_28527);
nand U29865 (N_29865,N_27817,N_28517);
or U29866 (N_29866,N_28046,N_28078);
xor U29867 (N_29867,N_27674,N_27667);
nor U29868 (N_29868,N_27820,N_28091);
nor U29869 (N_29869,N_28732,N_27639);
xnor U29870 (N_29870,N_28048,N_28120);
xnor U29871 (N_29871,N_28692,N_27979);
or U29872 (N_29872,N_27868,N_27642);
or U29873 (N_29873,N_28083,N_27930);
xor U29874 (N_29874,N_28466,N_28441);
nand U29875 (N_29875,N_28148,N_28199);
and U29876 (N_29876,N_28696,N_28318);
and U29877 (N_29877,N_28422,N_28313);
xnor U29878 (N_29878,N_27655,N_28472);
nor U29879 (N_29879,N_28702,N_28449);
and U29880 (N_29880,N_28096,N_28269);
nand U29881 (N_29881,N_28648,N_28797);
or U29882 (N_29882,N_28710,N_28142);
and U29883 (N_29883,N_28660,N_28151);
nand U29884 (N_29884,N_27679,N_28480);
or U29885 (N_29885,N_28394,N_28486);
and U29886 (N_29886,N_28740,N_28177);
or U29887 (N_29887,N_28165,N_28082);
or U29888 (N_29888,N_28702,N_28219);
nor U29889 (N_29889,N_28560,N_27836);
xor U29890 (N_29890,N_28328,N_28427);
or U29891 (N_29891,N_28554,N_28708);
or U29892 (N_29892,N_28487,N_28450);
nor U29893 (N_29893,N_28692,N_27995);
xor U29894 (N_29894,N_27758,N_28102);
xnor U29895 (N_29895,N_27626,N_28696);
nand U29896 (N_29896,N_28567,N_28351);
xor U29897 (N_29897,N_27770,N_28322);
or U29898 (N_29898,N_28677,N_27602);
nand U29899 (N_29899,N_27665,N_28240);
nand U29900 (N_29900,N_28640,N_27989);
xnor U29901 (N_29901,N_27695,N_28167);
or U29902 (N_29902,N_28328,N_28601);
xnor U29903 (N_29903,N_27624,N_28781);
xor U29904 (N_29904,N_28490,N_28124);
xnor U29905 (N_29905,N_27709,N_28492);
and U29906 (N_29906,N_28557,N_28751);
and U29907 (N_29907,N_27838,N_28439);
and U29908 (N_29908,N_28393,N_28547);
xnor U29909 (N_29909,N_28407,N_28285);
and U29910 (N_29910,N_27628,N_27999);
xnor U29911 (N_29911,N_28322,N_28481);
xor U29912 (N_29912,N_27733,N_28694);
xnor U29913 (N_29913,N_28484,N_27690);
nor U29914 (N_29914,N_27956,N_28632);
or U29915 (N_29915,N_28119,N_28323);
nor U29916 (N_29916,N_28530,N_28094);
and U29917 (N_29917,N_28617,N_27640);
nor U29918 (N_29918,N_27665,N_27745);
xnor U29919 (N_29919,N_27716,N_28037);
nor U29920 (N_29920,N_27929,N_27964);
and U29921 (N_29921,N_28134,N_28726);
or U29922 (N_29922,N_28138,N_28578);
or U29923 (N_29923,N_28766,N_27878);
xnor U29924 (N_29924,N_28193,N_28742);
nor U29925 (N_29925,N_28502,N_28477);
nand U29926 (N_29926,N_28220,N_27837);
and U29927 (N_29927,N_27816,N_27790);
or U29928 (N_29928,N_28206,N_27786);
xor U29929 (N_29929,N_28181,N_27664);
xor U29930 (N_29930,N_28791,N_27884);
and U29931 (N_29931,N_27962,N_28542);
xor U29932 (N_29932,N_28249,N_28192);
or U29933 (N_29933,N_28433,N_28012);
xnor U29934 (N_29934,N_27734,N_28469);
and U29935 (N_29935,N_28024,N_28737);
nor U29936 (N_29936,N_28720,N_28579);
or U29937 (N_29937,N_28523,N_27779);
nor U29938 (N_29938,N_28114,N_27621);
xor U29939 (N_29939,N_27740,N_28225);
or U29940 (N_29940,N_27657,N_28478);
nor U29941 (N_29941,N_27635,N_27662);
nor U29942 (N_29942,N_28061,N_27627);
nand U29943 (N_29943,N_28142,N_27817);
nand U29944 (N_29944,N_27889,N_27965);
nor U29945 (N_29945,N_27841,N_28301);
xnor U29946 (N_29946,N_28318,N_28779);
xor U29947 (N_29947,N_28234,N_27624);
and U29948 (N_29948,N_28796,N_28395);
xnor U29949 (N_29949,N_28340,N_28508);
or U29950 (N_29950,N_28560,N_28144);
nor U29951 (N_29951,N_27639,N_28570);
xnor U29952 (N_29952,N_28338,N_28641);
nand U29953 (N_29953,N_28774,N_27845);
and U29954 (N_29954,N_28492,N_27666);
or U29955 (N_29955,N_28597,N_28104);
and U29956 (N_29956,N_28190,N_28106);
nor U29957 (N_29957,N_28081,N_27909);
xnor U29958 (N_29958,N_27811,N_28757);
nor U29959 (N_29959,N_28723,N_27762);
and U29960 (N_29960,N_28379,N_28116);
and U29961 (N_29961,N_28408,N_27903);
or U29962 (N_29962,N_28773,N_28157);
xor U29963 (N_29963,N_28796,N_28411);
and U29964 (N_29964,N_27995,N_28103);
xnor U29965 (N_29965,N_27954,N_27822);
or U29966 (N_29966,N_27828,N_28507);
nand U29967 (N_29967,N_27900,N_28337);
nor U29968 (N_29968,N_27699,N_28719);
nand U29969 (N_29969,N_28481,N_28502);
xnor U29970 (N_29970,N_28279,N_28726);
xnor U29971 (N_29971,N_27950,N_28517);
nor U29972 (N_29972,N_27894,N_28552);
xor U29973 (N_29973,N_28444,N_28092);
or U29974 (N_29974,N_27631,N_27619);
xor U29975 (N_29975,N_27912,N_28448);
nand U29976 (N_29976,N_27738,N_28796);
or U29977 (N_29977,N_27770,N_28403);
nor U29978 (N_29978,N_28530,N_28599);
xor U29979 (N_29979,N_27819,N_28379);
nor U29980 (N_29980,N_27831,N_28331);
nor U29981 (N_29981,N_27827,N_28278);
and U29982 (N_29982,N_28400,N_27999);
nor U29983 (N_29983,N_28077,N_28090);
nand U29984 (N_29984,N_28544,N_28420);
and U29985 (N_29985,N_28673,N_28497);
and U29986 (N_29986,N_27899,N_28321);
nand U29987 (N_29987,N_27670,N_28109);
nor U29988 (N_29988,N_27722,N_27858);
and U29989 (N_29989,N_28289,N_28446);
nand U29990 (N_29990,N_27633,N_28077);
xor U29991 (N_29991,N_28252,N_27695);
and U29992 (N_29992,N_28700,N_28643);
nand U29993 (N_29993,N_28199,N_27883);
and U29994 (N_29994,N_28529,N_28579);
nand U29995 (N_29995,N_27922,N_28515);
and U29996 (N_29996,N_27946,N_28435);
nor U29997 (N_29997,N_28093,N_27701);
and U29998 (N_29998,N_28594,N_28212);
nor U29999 (N_29999,N_28087,N_28323);
nor UO_0 (O_0,N_29146,N_29099);
or UO_1 (O_1,N_29728,N_28867);
nand UO_2 (O_2,N_29580,N_29677);
and UO_3 (O_3,N_29774,N_29762);
and UO_4 (O_4,N_28810,N_29595);
and UO_5 (O_5,N_29490,N_28801);
nand UO_6 (O_6,N_29711,N_29046);
nor UO_7 (O_7,N_29107,N_28819);
or UO_8 (O_8,N_29620,N_29212);
nand UO_9 (O_9,N_28901,N_29476);
nor UO_10 (O_10,N_29614,N_28870);
or UO_11 (O_11,N_29816,N_29308);
nand UO_12 (O_12,N_29373,N_28973);
xnor UO_13 (O_13,N_29819,N_29846);
nand UO_14 (O_14,N_29756,N_29842);
xnor UO_15 (O_15,N_29596,N_29760);
nand UO_16 (O_16,N_29541,N_29252);
nor UO_17 (O_17,N_29351,N_29489);
nand UO_18 (O_18,N_29321,N_29686);
xnor UO_19 (O_19,N_29072,N_29440);
nor UO_20 (O_20,N_28887,N_28827);
xnor UO_21 (O_21,N_29334,N_29158);
nand UO_22 (O_22,N_29181,N_29486);
nand UO_23 (O_23,N_29950,N_28895);
xnor UO_24 (O_24,N_29436,N_29818);
and UO_25 (O_25,N_28861,N_29162);
nor UO_26 (O_26,N_29178,N_29098);
nor UO_27 (O_27,N_29786,N_29716);
or UO_28 (O_28,N_29828,N_29791);
nor UO_29 (O_29,N_29908,N_29832);
xnor UO_30 (O_30,N_29001,N_29301);
nor UO_31 (O_31,N_29938,N_29992);
nor UO_32 (O_32,N_29244,N_29531);
or UO_33 (O_33,N_29803,N_29149);
and UO_34 (O_34,N_29282,N_29473);
or UO_35 (O_35,N_28982,N_29112);
xor UO_36 (O_36,N_29172,N_28990);
xnor UO_37 (O_37,N_29635,N_29763);
nor UO_38 (O_38,N_29539,N_29556);
nand UO_39 (O_39,N_29984,N_29312);
nor UO_40 (O_40,N_29398,N_29933);
nand UO_41 (O_41,N_29513,N_29815);
or UO_42 (O_42,N_29666,N_29429);
and UO_43 (O_43,N_29055,N_29148);
xor UO_44 (O_44,N_29338,N_28996);
xnor UO_45 (O_45,N_29788,N_29865);
xor UO_46 (O_46,N_29236,N_28800);
nor UO_47 (O_47,N_29289,N_28933);
or UO_48 (O_48,N_29066,N_28875);
or UO_49 (O_49,N_29889,N_29777);
or UO_50 (O_50,N_29372,N_29462);
nand UO_51 (O_51,N_28864,N_29696);
xnor UO_52 (O_52,N_29968,N_29384);
nor UO_53 (O_53,N_29250,N_29010);
and UO_54 (O_54,N_29195,N_29131);
and UO_55 (O_55,N_29016,N_29798);
or UO_56 (O_56,N_29434,N_29594);
nand UO_57 (O_57,N_29501,N_29703);
nand UO_58 (O_58,N_29985,N_29603);
nand UO_59 (O_59,N_29015,N_29492);
xor UO_60 (O_60,N_29358,N_28803);
nand UO_61 (O_61,N_29392,N_29515);
xnor UO_62 (O_62,N_29602,N_29408);
and UO_63 (O_63,N_29163,N_29026);
xnor UO_64 (O_64,N_28897,N_29088);
xnor UO_65 (O_65,N_29262,N_28838);
or UO_66 (O_66,N_29736,N_29826);
or UO_67 (O_67,N_29482,N_29038);
xor UO_68 (O_68,N_29197,N_29533);
and UO_69 (O_69,N_29022,N_29318);
and UO_70 (O_70,N_29977,N_29738);
nor UO_71 (O_71,N_29494,N_29847);
nor UO_72 (O_72,N_29712,N_29278);
and UO_73 (O_73,N_29560,N_29902);
xnor UO_74 (O_74,N_29709,N_29797);
or UO_75 (O_75,N_29306,N_28899);
nor UO_76 (O_76,N_28960,N_29412);
or UO_77 (O_77,N_29914,N_29379);
and UO_78 (O_78,N_29733,N_29461);
xnor UO_79 (O_79,N_29708,N_29781);
and UO_80 (O_80,N_29921,N_29545);
or UO_81 (O_81,N_29600,N_29309);
nor UO_82 (O_82,N_29617,N_29987);
xnor UO_83 (O_83,N_29287,N_29725);
or UO_84 (O_84,N_29844,N_29220);
or UO_85 (O_85,N_29405,N_28994);
nor UO_86 (O_86,N_29537,N_29215);
nand UO_87 (O_87,N_29458,N_28986);
nand UO_88 (O_88,N_29028,N_29518);
nor UO_89 (O_89,N_28863,N_29199);
nor UO_90 (O_90,N_29974,N_29477);
or UO_91 (O_91,N_28939,N_29587);
and UO_92 (O_92,N_29087,N_29772);
and UO_93 (O_93,N_29357,N_28891);
and UO_94 (O_94,N_29993,N_29530);
nand UO_95 (O_95,N_29588,N_29428);
xor UO_96 (O_96,N_28988,N_29549);
xnor UO_97 (O_97,N_28970,N_29647);
xnor UO_98 (O_98,N_29198,N_29936);
or UO_99 (O_99,N_29070,N_29657);
or UO_100 (O_100,N_29329,N_29852);
nor UO_101 (O_101,N_29117,N_29367);
or UO_102 (O_102,N_29827,N_29551);
nand UO_103 (O_103,N_29031,N_28886);
nand UO_104 (O_104,N_29285,N_29455);
xnor UO_105 (O_105,N_29930,N_29590);
or UO_106 (O_106,N_28911,N_29390);
and UO_107 (O_107,N_29391,N_28907);
nand UO_108 (O_108,N_29886,N_28916);
and UO_109 (O_109,N_29344,N_29266);
or UO_110 (O_110,N_29323,N_29809);
nor UO_111 (O_111,N_29354,N_29114);
xnor UO_112 (O_112,N_29267,N_29277);
or UO_113 (O_113,N_29151,N_29562);
or UO_114 (O_114,N_29194,N_29075);
nand UO_115 (O_115,N_28856,N_28993);
nand UO_116 (O_116,N_29260,N_29964);
nand UO_117 (O_117,N_29157,N_29479);
nand UO_118 (O_118,N_29810,N_28913);
xnor UO_119 (O_119,N_29626,N_28823);
xnor UO_120 (O_120,N_28807,N_29694);
or UO_121 (O_121,N_29341,N_28981);
xnor UO_122 (O_122,N_28919,N_28859);
or UO_123 (O_123,N_29645,N_29954);
nand UO_124 (O_124,N_29871,N_29128);
nand UO_125 (O_125,N_29167,N_29205);
and UO_126 (O_126,N_29256,N_29432);
or UO_127 (O_127,N_29928,N_29339);
nand UO_128 (O_128,N_28825,N_29792);
xor UO_129 (O_129,N_29129,N_29960);
xor UO_130 (O_130,N_29059,N_29700);
and UO_131 (O_131,N_29425,N_29823);
and UO_132 (O_132,N_29717,N_29385);
and UO_133 (O_133,N_29737,N_29891);
or UO_134 (O_134,N_29898,N_29693);
xnor UO_135 (O_135,N_29978,N_29648);
nand UO_136 (O_136,N_29729,N_29187);
nand UO_137 (O_137,N_29459,N_29275);
or UO_138 (O_138,N_29794,N_29142);
xor UO_139 (O_139,N_29526,N_29997);
and UO_140 (O_140,N_29121,N_29271);
and UO_141 (O_141,N_29221,N_29495);
and UO_142 (O_142,N_28975,N_29421);
and UO_143 (O_143,N_29170,N_29288);
nor UO_144 (O_144,N_29448,N_29965);
and UO_145 (O_145,N_29855,N_29862);
nor UO_146 (O_146,N_28942,N_29917);
xnor UO_147 (O_147,N_28900,N_29397);
nand UO_148 (O_148,N_29245,N_29858);
nand UO_149 (O_149,N_29957,N_29156);
nand UO_150 (O_150,N_29656,N_29018);
nand UO_151 (O_151,N_29643,N_29893);
nor UO_152 (O_152,N_29592,N_28987);
nand UO_153 (O_153,N_29060,N_29519);
nor UO_154 (O_154,N_29542,N_29290);
nor UO_155 (O_155,N_29672,N_29520);
xnor UO_156 (O_156,N_29269,N_29222);
and UO_157 (O_157,N_28883,N_28839);
xnor UO_158 (O_158,N_29330,N_29235);
nor UO_159 (O_159,N_29808,N_29332);
and UO_160 (O_160,N_29535,N_29238);
and UO_161 (O_161,N_29021,N_29231);
xnor UO_162 (O_162,N_29184,N_29140);
nand UO_163 (O_163,N_28815,N_29982);
nand UO_164 (O_164,N_29609,N_29120);
nand UO_165 (O_165,N_29399,N_29848);
xnor UO_166 (O_166,N_29211,N_29650);
and UO_167 (O_167,N_28881,N_29979);
or UO_168 (O_168,N_29710,N_28843);
and UO_169 (O_169,N_28834,N_29869);
or UO_170 (O_170,N_29715,N_29570);
or UO_171 (O_171,N_29942,N_29039);
or UO_172 (O_172,N_29906,N_29517);
and UO_173 (O_173,N_29940,N_29822);
or UO_174 (O_174,N_29365,N_29835);
nand UO_175 (O_175,N_29583,N_29634);
xnor UO_176 (O_176,N_29228,N_29663);
nand UO_177 (O_177,N_28860,N_29108);
xor UO_178 (O_178,N_29474,N_29757);
nand UO_179 (O_179,N_29564,N_28852);
xor UO_180 (O_180,N_28956,N_29057);
nand UO_181 (O_181,N_29868,N_29577);
nand UO_182 (O_182,N_29919,N_28824);
or UO_183 (O_183,N_28908,N_29347);
nor UO_184 (O_184,N_29403,N_28873);
nor UO_185 (O_185,N_29470,N_29090);
or UO_186 (O_186,N_29655,N_29543);
or UO_187 (O_187,N_29177,N_28917);
or UO_188 (O_188,N_29969,N_29825);
nor UO_189 (O_189,N_28826,N_29012);
nor UO_190 (O_190,N_28920,N_29785);
or UO_191 (O_191,N_29901,N_29553);
nor UO_192 (O_192,N_28948,N_29190);
and UO_193 (O_193,N_29446,N_29346);
and UO_194 (O_194,N_29613,N_29702);
nand UO_195 (O_195,N_29293,N_29261);
xor UO_196 (O_196,N_29444,N_29746);
xnor UO_197 (O_197,N_29472,N_29811);
xnor UO_198 (O_198,N_29004,N_29654);
nand UO_199 (O_199,N_28876,N_29775);
or UO_200 (O_200,N_29510,N_28931);
nand UO_201 (O_201,N_28905,N_29850);
xnor UO_202 (O_202,N_28952,N_29457);
and UO_203 (O_203,N_29604,N_29966);
nor UO_204 (O_204,N_29662,N_29935);
or UO_205 (O_205,N_29297,N_29524);
or UO_206 (O_206,N_29989,N_29179);
or UO_207 (O_207,N_29652,N_29233);
and UO_208 (O_208,N_29475,N_29814);
nor UO_209 (O_209,N_29761,N_29375);
or UO_210 (O_210,N_29735,N_29413);
nor UO_211 (O_211,N_29561,N_29801);
or UO_212 (O_212,N_29527,N_29749);
nand UO_213 (O_213,N_28806,N_29006);
xor UO_214 (O_214,N_29821,N_29103);
nand UO_215 (O_215,N_29368,N_29019);
nand UO_216 (O_216,N_28847,N_28822);
xor UO_217 (O_217,N_28928,N_29175);
and UO_218 (O_218,N_29741,N_29320);
nor UO_219 (O_219,N_29382,N_29183);
or UO_220 (O_220,N_29817,N_29130);
and UO_221 (O_221,N_29104,N_29764);
or UO_222 (O_222,N_29887,N_29606);
and UO_223 (O_223,N_29544,N_29364);
and UO_224 (O_224,N_29831,N_29029);
and UO_225 (O_225,N_29900,N_29314);
nand UO_226 (O_226,N_29214,N_29851);
nand UO_227 (O_227,N_29496,N_29094);
nand UO_228 (O_228,N_29624,N_29502);
and UO_229 (O_229,N_29962,N_29186);
xnor UO_230 (O_230,N_28945,N_29892);
nor UO_231 (O_231,N_29273,N_29020);
nor UO_232 (O_232,N_28885,N_29101);
xnor UO_233 (O_233,N_29873,N_29879);
nand UO_234 (O_234,N_29731,N_29953);
or UO_235 (O_235,N_29644,N_29356);
nand UO_236 (O_236,N_29213,N_29795);
and UO_237 (O_237,N_29065,N_29008);
nand UO_238 (O_238,N_28935,N_29150);
nand UO_239 (O_239,N_29699,N_28893);
nand UO_240 (O_240,N_29034,N_29443);
xor UO_241 (O_241,N_28850,N_29591);
nor UO_242 (O_242,N_29122,N_29174);
or UO_243 (O_243,N_29705,N_29598);
and UO_244 (O_244,N_29319,N_29529);
and UO_245 (O_245,N_29581,N_29695);
or UO_246 (O_246,N_29507,N_29866);
xor UO_247 (O_247,N_28951,N_29359);
nor UO_248 (O_248,N_29949,N_29052);
and UO_249 (O_249,N_29687,N_29441);
nor UO_250 (O_250,N_29109,N_29488);
nor UO_251 (O_251,N_28947,N_29878);
nor UO_252 (O_252,N_29833,N_28969);
nor UO_253 (O_253,N_29780,N_29000);
xnor UO_254 (O_254,N_29202,N_29264);
or UO_255 (O_255,N_29920,N_29281);
or UO_256 (O_256,N_29386,N_29134);
or UO_257 (O_257,N_29371,N_28929);
and UO_258 (O_258,N_29732,N_28912);
and UO_259 (O_259,N_29619,N_29680);
nor UO_260 (O_260,N_29996,N_28921);
and UO_261 (O_261,N_28940,N_29569);
xnor UO_262 (O_262,N_28836,N_28848);
nor UO_263 (O_263,N_29514,N_29904);
nor UO_264 (O_264,N_28927,N_29924);
and UO_265 (O_265,N_29983,N_29909);
or UO_266 (O_266,N_29929,N_29927);
or UO_267 (O_267,N_29417,N_29073);
xnor UO_268 (O_268,N_29916,N_29931);
nor UO_269 (O_269,N_28846,N_29779);
nand UO_270 (O_270,N_29383,N_28992);
and UO_271 (O_271,N_29415,N_29110);
nor UO_272 (O_272,N_29387,N_29802);
or UO_273 (O_273,N_29208,N_29546);
nor UO_274 (O_274,N_29509,N_29124);
and UO_275 (O_275,N_29947,N_29086);
xor UO_276 (O_276,N_29895,N_29324);
nor UO_277 (O_277,N_28936,N_29555);
and UO_278 (O_278,N_29582,N_29234);
nand UO_279 (O_279,N_29361,N_29721);
xnor UO_280 (O_280,N_29854,N_29912);
or UO_281 (O_281,N_28985,N_29951);
xor UO_282 (O_282,N_28957,N_29667);
xor UO_283 (O_283,N_29718,N_29678);
nor UO_284 (O_284,N_29601,N_29500);
or UO_285 (O_285,N_28914,N_28871);
and UO_286 (O_286,N_29279,N_29225);
nor UO_287 (O_287,N_29299,N_29505);
xor UO_288 (O_288,N_29229,N_29074);
nor UO_289 (O_289,N_29239,N_28889);
or UO_290 (O_290,N_28842,N_28878);
nand UO_291 (O_291,N_29210,N_29998);
and UO_292 (O_292,N_29925,N_29637);
and UO_293 (O_293,N_29830,N_29483);
nor UO_294 (O_294,N_29302,N_29952);
or UO_295 (O_295,N_29793,N_28857);
nand UO_296 (O_296,N_29433,N_28816);
and UO_297 (O_297,N_29240,N_29726);
and UO_298 (O_298,N_29438,N_29303);
and UO_299 (O_299,N_29013,N_29192);
nand UO_300 (O_300,N_28998,N_29783);
nand UO_301 (O_301,N_29430,N_29973);
nand UO_302 (O_302,N_29758,N_29536);
xnor UO_303 (O_303,N_29575,N_29599);
nand UO_304 (O_304,N_29431,N_29999);
nand UO_305 (O_305,N_29144,N_29911);
nor UO_306 (O_306,N_29525,N_29076);
xnor UO_307 (O_307,N_29316,N_29048);
xor UO_308 (O_308,N_29532,N_29932);
nand UO_309 (O_309,N_29340,N_29552);
xnor UO_310 (O_310,N_29706,N_29414);
or UO_311 (O_311,N_29880,N_29284);
or UO_312 (O_312,N_29342,N_28950);
xor UO_313 (O_313,N_29480,N_29054);
and UO_314 (O_314,N_29607,N_29493);
or UO_315 (O_315,N_29307,N_29169);
xor UO_316 (O_316,N_29789,N_29685);
xnor UO_317 (O_317,N_29300,N_28818);
xnor UO_318 (O_318,N_29946,N_28909);
nand UO_319 (O_319,N_29800,N_29478);
xor UO_320 (O_320,N_29463,N_29841);
nor UO_321 (O_321,N_29790,N_29298);
nor UO_322 (O_322,N_29196,N_29366);
and UO_323 (O_323,N_29755,N_29043);
or UO_324 (O_324,N_28851,N_29040);
xnor UO_325 (O_325,N_29032,N_29905);
xor UO_326 (O_326,N_29897,N_29396);
and UO_327 (O_327,N_29200,N_28923);
nand UO_328 (O_328,N_29102,N_29584);
nand UO_329 (O_329,N_29939,N_28967);
and UO_330 (O_330,N_29487,N_28844);
or UO_331 (O_331,N_29132,N_29115);
or UO_332 (O_332,N_29007,N_29166);
nand UO_333 (O_333,N_29631,N_29325);
xor UO_334 (O_334,N_29730,N_29137);
or UO_335 (O_335,N_29597,N_29870);
or UO_336 (O_336,N_29263,N_29464);
or UO_337 (O_337,N_29995,N_28946);
or UO_338 (O_338,N_29310,N_29388);
nand UO_339 (O_339,N_29812,N_29585);
and UO_340 (O_340,N_29503,N_28892);
or UO_341 (O_341,N_29498,N_29125);
nor UO_342 (O_342,N_29770,N_29119);
or UO_343 (O_343,N_29322,N_29744);
nand UO_344 (O_344,N_29750,N_28812);
nand UO_345 (O_345,N_29521,N_29305);
nor UO_346 (O_346,N_29380,N_29419);
nand UO_347 (O_347,N_29679,N_29171);
nor UO_348 (O_348,N_28965,N_29682);
xor UO_349 (O_349,N_29751,N_28963);
nand UO_350 (O_350,N_29216,N_28983);
xnor UO_351 (O_351,N_29217,N_29481);
and UO_352 (O_352,N_28829,N_28954);
xnor UO_353 (O_353,N_29037,N_29426);
xnor UO_354 (O_354,N_29247,N_29009);
and UO_355 (O_355,N_29834,N_29859);
nand UO_356 (O_356,N_29374,N_29990);
nand UO_357 (O_357,N_29050,N_28906);
nand UO_358 (O_358,N_29941,N_29230);
nand UO_359 (O_359,N_28837,N_29336);
and UO_360 (O_360,N_29056,N_29690);
nor UO_361 (O_361,N_29661,N_28971);
and UO_362 (O_362,N_29623,N_28968);
xor UO_363 (O_363,N_29625,N_29068);
or UO_364 (O_364,N_29218,N_29499);
or UO_365 (O_365,N_29024,N_29097);
nand UO_366 (O_366,N_28862,N_29437);
nor UO_367 (O_367,N_29402,N_29683);
and UO_368 (O_368,N_29722,N_29572);
or UO_369 (O_369,N_29899,N_29155);
or UO_370 (O_370,N_28880,N_28841);
nand UO_371 (O_371,N_29867,N_29460);
and UO_372 (O_372,N_29565,N_29512);
nor UO_373 (O_373,N_29427,N_28808);
or UO_374 (O_374,N_29720,N_29017);
or UO_375 (O_375,N_29265,N_28814);
nand UO_376 (O_376,N_29540,N_29424);
nor UO_377 (O_377,N_29274,N_28845);
and UO_378 (O_378,N_29471,N_29389);
nand UO_379 (O_379,N_28872,N_29159);
xnor UO_380 (O_380,N_29042,N_29566);
or UO_381 (O_381,N_29352,N_28910);
nand UO_382 (O_382,N_29804,N_29449);
nand UO_383 (O_383,N_29376,N_29910);
or UO_384 (O_384,N_29547,N_28953);
or UO_385 (O_385,N_29395,N_29669);
xor UO_386 (O_386,N_29106,N_29639);
nor UO_387 (O_387,N_29689,N_28868);
or UO_388 (O_388,N_29105,N_29608);
and UO_389 (O_389,N_29141,N_29116);
nor UO_390 (O_390,N_29857,N_28989);
or UO_391 (O_391,N_29051,N_28943);
or UO_392 (O_392,N_28958,N_28849);
nand UO_393 (O_393,N_29283,N_28811);
nor UO_394 (O_394,N_29630,N_29836);
nand UO_395 (O_395,N_29734,N_29853);
nand UO_396 (O_396,N_29280,N_29207);
xnor UO_397 (O_397,N_29664,N_29856);
nand UO_398 (O_398,N_29508,N_29956);
or UO_399 (O_399,N_28991,N_29069);
or UO_400 (O_400,N_29860,N_28894);
and UO_401 (O_401,N_29145,N_29615);
nor UO_402 (O_402,N_29123,N_29067);
nand UO_403 (O_403,N_29986,N_29410);
nand UO_404 (O_404,N_28884,N_29874);
or UO_405 (O_405,N_29994,N_29003);
xor UO_406 (O_406,N_29296,N_29885);
xnor UO_407 (O_407,N_29538,N_29988);
or UO_408 (O_408,N_29714,N_29154);
nor UO_409 (O_409,N_29232,N_28831);
nor UO_410 (O_410,N_29411,N_29922);
and UO_411 (O_411,N_29673,N_29084);
xor UO_412 (O_412,N_29681,N_29201);
xor UO_413 (O_413,N_29328,N_29743);
nand UO_414 (O_414,N_28853,N_29360);
or UO_415 (O_415,N_29511,N_29739);
nor UO_416 (O_416,N_28932,N_29863);
and UO_417 (O_417,N_29589,N_28938);
and UO_418 (O_418,N_29778,N_29618);
xor UO_419 (O_419,N_29972,N_29100);
xor UO_420 (O_420,N_29903,N_29317);
or UO_421 (O_421,N_29872,N_29058);
nor UO_422 (O_422,N_29467,N_29345);
xor UO_423 (O_423,N_29091,N_29333);
nor UO_424 (O_424,N_29085,N_29092);
xor UO_425 (O_425,N_29701,N_29369);
and UO_426 (O_426,N_28874,N_29049);
or UO_427 (O_427,N_29035,N_29571);
nor UO_428 (O_428,N_29971,N_29394);
nor UO_429 (O_429,N_28854,N_29041);
or UO_430 (O_430,N_29468,N_29724);
xnor UO_431 (O_431,N_29567,N_29133);
xnor UO_432 (O_432,N_29745,N_29161);
xor UO_433 (O_433,N_29829,N_29407);
or UO_434 (O_434,N_29504,N_29636);
nor UO_435 (O_435,N_28959,N_28964);
xor UO_436 (O_436,N_29295,N_29030);
or UO_437 (O_437,N_29651,N_29534);
or UO_438 (O_438,N_29135,N_29173);
or UO_439 (O_439,N_29767,N_29890);
nor UO_440 (O_440,N_29404,N_29023);
xnor UO_441 (O_441,N_29875,N_29451);
nor UO_442 (O_442,N_28877,N_29967);
or UO_443 (O_443,N_29136,N_29888);
xor UO_444 (O_444,N_29884,N_29079);
nand UO_445 (O_445,N_29840,N_29576);
nand UO_446 (O_446,N_29522,N_29688);
nor UO_447 (O_447,N_29423,N_28865);
or UO_448 (O_448,N_29189,N_29350);
or UO_449 (O_449,N_29506,N_29313);
nor UO_450 (O_450,N_28903,N_29053);
nand UO_451 (O_451,N_29629,N_29450);
nand UO_452 (O_452,N_29568,N_29698);
or UO_453 (O_453,N_29675,N_29627);
or UO_454 (O_454,N_29554,N_28995);
and UO_455 (O_455,N_29837,N_29268);
xnor UO_456 (O_456,N_29574,N_29061);
xor UO_457 (O_457,N_29241,N_29227);
and UO_458 (O_458,N_29557,N_29353);
xnor UO_459 (O_459,N_29578,N_28902);
and UO_460 (O_460,N_29160,N_29326);
nor UO_461 (O_461,N_29861,N_28821);
or UO_462 (O_462,N_29409,N_28925);
xor UO_463 (O_463,N_29484,N_29692);
nor UO_464 (O_464,N_29605,N_29782);
or UO_465 (O_465,N_29176,N_29913);
nor UO_466 (O_466,N_28896,N_29378);
nor UO_467 (O_467,N_29014,N_29945);
xor UO_468 (O_468,N_29077,N_29676);
nand UO_469 (O_469,N_28855,N_29027);
or UO_470 (O_470,N_29343,N_29838);
and UO_471 (O_471,N_29845,N_28924);
nor UO_472 (O_472,N_29418,N_28922);
nor UO_473 (O_473,N_29002,N_29454);
nand UO_474 (O_474,N_29168,N_29707);
and UO_475 (O_475,N_29658,N_29113);
nand UO_476 (O_476,N_29182,N_29401);
nand UO_477 (O_477,N_29528,N_28813);
or UO_478 (O_478,N_29980,N_28984);
xnor UO_479 (O_479,N_29628,N_29447);
and UO_480 (O_480,N_29991,N_28962);
xor UO_481 (O_481,N_29670,N_29704);
and UO_482 (O_482,N_28955,N_29025);
nor UO_483 (O_483,N_29491,N_29349);
or UO_484 (O_484,N_29078,N_29251);
nand UO_485 (O_485,N_29548,N_29671);
xnor UO_486 (O_486,N_29456,N_28830);
xnor UO_487 (O_487,N_29422,N_29713);
xor UO_488 (O_488,N_28835,N_29466);
or UO_489 (O_489,N_29082,N_28944);
and UO_490 (O_490,N_28974,N_29400);
or UO_491 (O_491,N_29523,N_29820);
and UO_492 (O_492,N_29337,N_28941);
nand UO_493 (O_493,N_29719,N_29573);
or UO_494 (O_494,N_29796,N_29640);
or UO_495 (O_495,N_29381,N_29579);
nor UO_496 (O_496,N_29766,N_29276);
nor UO_497 (O_497,N_29355,N_29754);
and UO_498 (O_498,N_29918,N_29616);
xnor UO_499 (O_499,N_29005,N_29944);
or UO_500 (O_500,N_29649,N_29806);
nor UO_501 (O_501,N_29420,N_28817);
nor UO_502 (O_502,N_28980,N_29416);
nor UO_503 (O_503,N_29242,N_29915);
and UO_504 (O_504,N_29219,N_29959);
nand UO_505 (O_505,N_29209,N_29748);
or UO_506 (O_506,N_29961,N_29249);
or UO_507 (O_507,N_29047,N_28961);
or UO_508 (O_508,N_29193,N_29272);
or UO_509 (O_509,N_29185,N_28972);
and UO_510 (O_510,N_28832,N_29062);
or UO_511 (O_511,N_28805,N_29180);
nor UO_512 (O_512,N_28997,N_28976);
nor UO_513 (O_513,N_28949,N_29246);
xnor UO_514 (O_514,N_29452,N_29291);
nand UO_515 (O_515,N_29882,N_29877);
xnor UO_516 (O_516,N_29611,N_29033);
and UO_517 (O_517,N_29976,N_29660);
xor UO_518 (O_518,N_29096,N_29363);
xnor UO_519 (O_519,N_28882,N_29485);
nor UO_520 (O_520,N_29586,N_29923);
or UO_521 (O_521,N_29784,N_29632);
and UO_522 (O_522,N_29612,N_29327);
nand UO_523 (O_523,N_29926,N_29093);
and UO_524 (O_524,N_29610,N_29362);
nor UO_525 (O_525,N_29638,N_29377);
nor UO_526 (O_526,N_28828,N_29805);
or UO_527 (O_527,N_29691,N_29152);
nand UO_528 (O_528,N_29453,N_29188);
xnor UO_529 (O_529,N_29907,N_29769);
and UO_530 (O_530,N_29622,N_28898);
nor UO_531 (O_531,N_29044,N_29089);
xnor UO_532 (O_532,N_29165,N_29684);
nor UO_533 (O_533,N_29143,N_28820);
and UO_534 (O_534,N_29445,N_29393);
nand UO_535 (O_535,N_28978,N_28809);
nand UO_536 (O_536,N_29081,N_28934);
and UO_537 (O_537,N_29593,N_28918);
nand UO_538 (O_538,N_29621,N_29011);
xnor UO_539 (O_539,N_29147,N_29080);
nand UO_540 (O_540,N_29226,N_29975);
nor UO_541 (O_541,N_29139,N_29191);
or UO_542 (O_542,N_28904,N_29727);
and UO_543 (O_543,N_29981,N_29071);
or UO_544 (O_544,N_29558,N_29697);
nor UO_545 (O_545,N_29752,N_28915);
and UO_546 (O_546,N_29559,N_29665);
or UO_547 (O_547,N_29937,N_29083);
nor UO_548 (O_548,N_29063,N_29864);
nor UO_549 (O_549,N_29894,N_29883);
or UO_550 (O_550,N_28804,N_29248);
and UO_551 (O_551,N_29331,N_29787);
nand UO_552 (O_552,N_29753,N_29668);
nand UO_553 (O_553,N_29292,N_29258);
xor UO_554 (O_554,N_29294,N_29253);
xor UO_555 (O_555,N_29768,N_29674);
and UO_556 (O_556,N_29127,N_29237);
nand UO_557 (O_557,N_29304,N_29934);
or UO_558 (O_558,N_29224,N_29659);
xnor UO_559 (O_559,N_28879,N_28930);
nor UO_560 (O_560,N_29435,N_28926);
nor UO_561 (O_561,N_29799,N_29203);
nand UO_562 (O_562,N_29311,N_29118);
nor UO_563 (O_563,N_29164,N_29439);
and UO_564 (O_564,N_29723,N_29286);
nor UO_565 (O_565,N_29896,N_29255);
xnor UO_566 (O_566,N_28840,N_29839);
or UO_567 (O_567,N_29653,N_29881);
nor UO_568 (O_568,N_29465,N_29641);
xnor UO_569 (O_569,N_29958,N_28937);
or UO_570 (O_570,N_29633,N_28802);
nand UO_571 (O_571,N_29095,N_28888);
and UO_572 (O_572,N_29064,N_29943);
nor UO_573 (O_573,N_28858,N_29642);
nor UO_574 (O_574,N_29849,N_29259);
nand UO_575 (O_575,N_28866,N_29824);
and UO_576 (O_576,N_28979,N_29563);
or UO_577 (O_577,N_29516,N_29963);
and UO_578 (O_578,N_29876,N_29111);
nand UO_579 (O_579,N_29765,N_28833);
nand UO_580 (O_580,N_29776,N_29469);
xor UO_581 (O_581,N_29206,N_29550);
and UO_582 (O_582,N_28977,N_29138);
nor UO_583 (O_583,N_29955,N_29270);
xor UO_584 (O_584,N_29257,N_29843);
xnor UO_585 (O_585,N_29970,N_29740);
nand UO_586 (O_586,N_29807,N_29646);
or UO_587 (O_587,N_28890,N_29497);
xnor UO_588 (O_588,N_29126,N_29204);
and UO_589 (O_589,N_29315,N_29045);
or UO_590 (O_590,N_29948,N_29153);
nand UO_591 (O_591,N_28869,N_29747);
and UO_592 (O_592,N_29773,N_29742);
nor UO_593 (O_593,N_29442,N_29036);
xor UO_594 (O_594,N_28966,N_29223);
or UO_595 (O_595,N_29759,N_29370);
or UO_596 (O_596,N_29406,N_29813);
nand UO_597 (O_597,N_29771,N_28999);
xnor UO_598 (O_598,N_29254,N_29335);
nand UO_599 (O_599,N_29348,N_29243);
and UO_600 (O_600,N_29498,N_28858);
and UO_601 (O_601,N_29741,N_29067);
or UO_602 (O_602,N_29592,N_29447);
and UO_603 (O_603,N_29401,N_29174);
and UO_604 (O_604,N_29829,N_29103);
or UO_605 (O_605,N_29737,N_29732);
or UO_606 (O_606,N_28956,N_28871);
and UO_607 (O_607,N_29687,N_28918);
nand UO_608 (O_608,N_29617,N_29241);
and UO_609 (O_609,N_29032,N_29438);
xor UO_610 (O_610,N_29643,N_29892);
nor UO_611 (O_611,N_29430,N_29741);
or UO_612 (O_612,N_29883,N_29734);
or UO_613 (O_613,N_29509,N_29722);
nor UO_614 (O_614,N_28882,N_29953);
and UO_615 (O_615,N_29396,N_29664);
nand UO_616 (O_616,N_29920,N_29829);
and UO_617 (O_617,N_28831,N_28905);
nand UO_618 (O_618,N_29286,N_29909);
nand UO_619 (O_619,N_29407,N_29782);
nor UO_620 (O_620,N_29516,N_29722);
xor UO_621 (O_621,N_29964,N_29095);
nand UO_622 (O_622,N_29775,N_29062);
nor UO_623 (O_623,N_29579,N_29340);
or UO_624 (O_624,N_29267,N_29045);
and UO_625 (O_625,N_29901,N_28950);
nand UO_626 (O_626,N_29186,N_29467);
and UO_627 (O_627,N_28977,N_29440);
xor UO_628 (O_628,N_29925,N_29450);
xor UO_629 (O_629,N_29896,N_28933);
nand UO_630 (O_630,N_29630,N_28947);
nor UO_631 (O_631,N_29601,N_29876);
nand UO_632 (O_632,N_29049,N_29339);
or UO_633 (O_633,N_28904,N_29652);
nor UO_634 (O_634,N_29857,N_28854);
and UO_635 (O_635,N_29623,N_29510);
nand UO_636 (O_636,N_29449,N_28921);
xnor UO_637 (O_637,N_29917,N_29453);
and UO_638 (O_638,N_29311,N_29089);
nand UO_639 (O_639,N_29284,N_29037);
and UO_640 (O_640,N_28844,N_29516);
and UO_641 (O_641,N_29868,N_29490);
and UO_642 (O_642,N_29584,N_29120);
nor UO_643 (O_643,N_29703,N_29872);
and UO_644 (O_644,N_29323,N_29867);
nor UO_645 (O_645,N_28879,N_29719);
and UO_646 (O_646,N_29966,N_29039);
xor UO_647 (O_647,N_29300,N_29050);
nor UO_648 (O_648,N_29074,N_29257);
or UO_649 (O_649,N_28902,N_28930);
or UO_650 (O_650,N_29329,N_28887);
and UO_651 (O_651,N_29146,N_29022);
xor UO_652 (O_652,N_29054,N_29194);
or UO_653 (O_653,N_28946,N_29152);
and UO_654 (O_654,N_28875,N_29271);
nand UO_655 (O_655,N_29760,N_29856);
xnor UO_656 (O_656,N_29474,N_29156);
or UO_657 (O_657,N_29152,N_29580);
nand UO_658 (O_658,N_29095,N_29768);
and UO_659 (O_659,N_29772,N_29533);
nor UO_660 (O_660,N_29588,N_29474);
xor UO_661 (O_661,N_29356,N_29573);
nand UO_662 (O_662,N_29101,N_29513);
xor UO_663 (O_663,N_29564,N_29663);
or UO_664 (O_664,N_29180,N_29920);
xnor UO_665 (O_665,N_29188,N_29910);
nand UO_666 (O_666,N_29430,N_28884);
or UO_667 (O_667,N_29554,N_28828);
nand UO_668 (O_668,N_29767,N_29422);
and UO_669 (O_669,N_29424,N_29267);
or UO_670 (O_670,N_28833,N_29626);
and UO_671 (O_671,N_29888,N_29306);
or UO_672 (O_672,N_29697,N_29071);
xnor UO_673 (O_673,N_28931,N_28916);
or UO_674 (O_674,N_29744,N_28807);
nand UO_675 (O_675,N_29213,N_29264);
and UO_676 (O_676,N_29261,N_29322);
nand UO_677 (O_677,N_29075,N_28813);
xor UO_678 (O_678,N_29966,N_28831);
and UO_679 (O_679,N_29554,N_29922);
and UO_680 (O_680,N_29081,N_28891);
or UO_681 (O_681,N_29855,N_29863);
nand UO_682 (O_682,N_29843,N_29770);
and UO_683 (O_683,N_29057,N_29469);
or UO_684 (O_684,N_29917,N_29933);
nor UO_685 (O_685,N_29737,N_29293);
nand UO_686 (O_686,N_29769,N_29356);
nor UO_687 (O_687,N_29277,N_29656);
nand UO_688 (O_688,N_29288,N_28826);
and UO_689 (O_689,N_29321,N_29471);
nand UO_690 (O_690,N_28920,N_28842);
nor UO_691 (O_691,N_28936,N_29207);
and UO_692 (O_692,N_29255,N_28877);
or UO_693 (O_693,N_29718,N_29318);
or UO_694 (O_694,N_29681,N_29532);
nand UO_695 (O_695,N_28967,N_29940);
nor UO_696 (O_696,N_29507,N_28890);
or UO_697 (O_697,N_28818,N_29608);
nor UO_698 (O_698,N_29154,N_28815);
nor UO_699 (O_699,N_29436,N_29175);
or UO_700 (O_700,N_29930,N_29427);
xor UO_701 (O_701,N_29201,N_29067);
and UO_702 (O_702,N_29230,N_29169);
or UO_703 (O_703,N_29884,N_29911);
nand UO_704 (O_704,N_28917,N_28906);
xnor UO_705 (O_705,N_29776,N_28986);
xnor UO_706 (O_706,N_29209,N_29802);
xor UO_707 (O_707,N_28829,N_29064);
nand UO_708 (O_708,N_29630,N_29063);
xnor UO_709 (O_709,N_28907,N_29733);
nor UO_710 (O_710,N_29491,N_29414);
nand UO_711 (O_711,N_29604,N_29162);
xnor UO_712 (O_712,N_28870,N_29059);
xnor UO_713 (O_713,N_29195,N_29246);
or UO_714 (O_714,N_28807,N_29083);
nand UO_715 (O_715,N_29926,N_29281);
xnor UO_716 (O_716,N_28976,N_28817);
or UO_717 (O_717,N_29720,N_29950);
nor UO_718 (O_718,N_29018,N_29665);
and UO_719 (O_719,N_29605,N_28961);
nand UO_720 (O_720,N_29479,N_29645);
xnor UO_721 (O_721,N_29623,N_29023);
nor UO_722 (O_722,N_28904,N_29271);
and UO_723 (O_723,N_29237,N_29204);
and UO_724 (O_724,N_28886,N_29569);
and UO_725 (O_725,N_29070,N_29444);
nor UO_726 (O_726,N_28851,N_29397);
nand UO_727 (O_727,N_29334,N_29384);
or UO_728 (O_728,N_29233,N_29664);
nor UO_729 (O_729,N_29346,N_29568);
xnor UO_730 (O_730,N_29671,N_29038);
or UO_731 (O_731,N_28854,N_29328);
and UO_732 (O_732,N_29591,N_29514);
or UO_733 (O_733,N_29276,N_29993);
nand UO_734 (O_734,N_29907,N_29710);
nand UO_735 (O_735,N_29246,N_29635);
xor UO_736 (O_736,N_29399,N_29823);
nand UO_737 (O_737,N_28877,N_29119);
nor UO_738 (O_738,N_29025,N_29933);
or UO_739 (O_739,N_29810,N_29507);
nand UO_740 (O_740,N_28914,N_28820);
or UO_741 (O_741,N_29929,N_29653);
nand UO_742 (O_742,N_29776,N_29374);
nand UO_743 (O_743,N_28805,N_29987);
or UO_744 (O_744,N_28972,N_29665);
nand UO_745 (O_745,N_28854,N_29546);
xor UO_746 (O_746,N_29108,N_29983);
xor UO_747 (O_747,N_29683,N_29255);
nand UO_748 (O_748,N_29460,N_29487);
nand UO_749 (O_749,N_29596,N_29181);
nand UO_750 (O_750,N_29341,N_29013);
xnor UO_751 (O_751,N_29913,N_29169);
and UO_752 (O_752,N_29906,N_29546);
nor UO_753 (O_753,N_29066,N_29417);
nor UO_754 (O_754,N_28909,N_29958);
nand UO_755 (O_755,N_29754,N_29053);
or UO_756 (O_756,N_29615,N_28985);
and UO_757 (O_757,N_29510,N_29856);
and UO_758 (O_758,N_29518,N_28933);
and UO_759 (O_759,N_29449,N_29972);
and UO_760 (O_760,N_29365,N_29496);
and UO_761 (O_761,N_29294,N_29243);
nand UO_762 (O_762,N_28855,N_29661);
and UO_763 (O_763,N_29458,N_29475);
nor UO_764 (O_764,N_28968,N_29604);
xnor UO_765 (O_765,N_29423,N_29730);
nor UO_766 (O_766,N_29765,N_29517);
nor UO_767 (O_767,N_28812,N_29391);
nor UO_768 (O_768,N_28845,N_29503);
nand UO_769 (O_769,N_29368,N_29958);
nand UO_770 (O_770,N_28939,N_28868);
or UO_771 (O_771,N_29310,N_29746);
nor UO_772 (O_772,N_29802,N_29902);
or UO_773 (O_773,N_29387,N_29117);
xor UO_774 (O_774,N_28831,N_29277);
and UO_775 (O_775,N_29285,N_28846);
xor UO_776 (O_776,N_29610,N_29155);
nand UO_777 (O_777,N_28934,N_28988);
nor UO_778 (O_778,N_29041,N_29270);
xor UO_779 (O_779,N_29501,N_29974);
nor UO_780 (O_780,N_29670,N_29787);
xor UO_781 (O_781,N_29230,N_28860);
nor UO_782 (O_782,N_29998,N_29235);
xnor UO_783 (O_783,N_29599,N_28868);
and UO_784 (O_784,N_29020,N_29503);
or UO_785 (O_785,N_29341,N_29474);
xor UO_786 (O_786,N_28942,N_28900);
xnor UO_787 (O_787,N_29107,N_28976);
or UO_788 (O_788,N_29909,N_28998);
xor UO_789 (O_789,N_29287,N_29060);
nand UO_790 (O_790,N_29099,N_29707);
xor UO_791 (O_791,N_28998,N_29362);
xor UO_792 (O_792,N_29067,N_29895);
nor UO_793 (O_793,N_28881,N_28862);
nand UO_794 (O_794,N_29840,N_29630);
nand UO_795 (O_795,N_29628,N_29727);
or UO_796 (O_796,N_29002,N_29764);
xnor UO_797 (O_797,N_29677,N_29383);
and UO_798 (O_798,N_29517,N_29137);
xor UO_799 (O_799,N_29807,N_29568);
xor UO_800 (O_800,N_29814,N_28854);
nor UO_801 (O_801,N_28963,N_29806);
and UO_802 (O_802,N_29790,N_28826);
xor UO_803 (O_803,N_29411,N_29869);
nor UO_804 (O_804,N_29775,N_29530);
and UO_805 (O_805,N_29193,N_29477);
and UO_806 (O_806,N_28962,N_29793);
nand UO_807 (O_807,N_29034,N_29781);
nand UO_808 (O_808,N_29666,N_29763);
and UO_809 (O_809,N_28871,N_29548);
nor UO_810 (O_810,N_29703,N_29100);
xnor UO_811 (O_811,N_29303,N_29288);
xnor UO_812 (O_812,N_29732,N_29781);
or UO_813 (O_813,N_29709,N_28891);
or UO_814 (O_814,N_29804,N_29753);
nor UO_815 (O_815,N_29090,N_28940);
nand UO_816 (O_816,N_29179,N_29484);
nor UO_817 (O_817,N_29174,N_29062);
xnor UO_818 (O_818,N_29454,N_29634);
nand UO_819 (O_819,N_29722,N_29607);
xor UO_820 (O_820,N_29784,N_29642);
nand UO_821 (O_821,N_29965,N_28974);
or UO_822 (O_822,N_29109,N_29228);
xor UO_823 (O_823,N_29855,N_29359);
or UO_824 (O_824,N_29579,N_29134);
nor UO_825 (O_825,N_29682,N_29580);
nor UO_826 (O_826,N_28932,N_29460);
nand UO_827 (O_827,N_29382,N_29805);
nor UO_828 (O_828,N_29909,N_29313);
nand UO_829 (O_829,N_28831,N_29909);
nor UO_830 (O_830,N_29194,N_29218);
or UO_831 (O_831,N_29277,N_29601);
or UO_832 (O_832,N_28927,N_28898);
xor UO_833 (O_833,N_29224,N_29389);
and UO_834 (O_834,N_29542,N_29587);
and UO_835 (O_835,N_29885,N_29154);
or UO_836 (O_836,N_29143,N_29912);
xnor UO_837 (O_837,N_29370,N_29503);
or UO_838 (O_838,N_29949,N_29712);
xnor UO_839 (O_839,N_28944,N_29423);
xor UO_840 (O_840,N_29129,N_29282);
nand UO_841 (O_841,N_29897,N_29846);
nand UO_842 (O_842,N_29558,N_29957);
nand UO_843 (O_843,N_28926,N_29699);
and UO_844 (O_844,N_29582,N_29997);
xnor UO_845 (O_845,N_29360,N_29909);
or UO_846 (O_846,N_28987,N_28981);
or UO_847 (O_847,N_29054,N_29706);
and UO_848 (O_848,N_29759,N_28809);
xnor UO_849 (O_849,N_29576,N_29448);
and UO_850 (O_850,N_29384,N_29440);
nand UO_851 (O_851,N_28890,N_29031);
xor UO_852 (O_852,N_29001,N_29297);
nand UO_853 (O_853,N_29656,N_29153);
xor UO_854 (O_854,N_29415,N_29221);
and UO_855 (O_855,N_29396,N_29022);
and UO_856 (O_856,N_29580,N_28986);
nor UO_857 (O_857,N_29786,N_29900);
nand UO_858 (O_858,N_29771,N_29669);
nand UO_859 (O_859,N_29465,N_28969);
xnor UO_860 (O_860,N_29975,N_29623);
and UO_861 (O_861,N_28941,N_28876);
or UO_862 (O_862,N_29627,N_29891);
nor UO_863 (O_863,N_29886,N_29475);
xnor UO_864 (O_864,N_29462,N_28911);
xnor UO_865 (O_865,N_29282,N_29046);
or UO_866 (O_866,N_29678,N_28895);
nor UO_867 (O_867,N_28899,N_29212);
or UO_868 (O_868,N_29602,N_29825);
xnor UO_869 (O_869,N_29028,N_29067);
nand UO_870 (O_870,N_28825,N_29235);
nor UO_871 (O_871,N_29643,N_29711);
nor UO_872 (O_872,N_28925,N_29003);
nor UO_873 (O_873,N_29865,N_29653);
and UO_874 (O_874,N_29627,N_28816);
or UO_875 (O_875,N_29085,N_29065);
nand UO_876 (O_876,N_29135,N_29709);
or UO_877 (O_877,N_29581,N_29242);
and UO_878 (O_878,N_29508,N_28971);
nand UO_879 (O_879,N_28983,N_28864);
xnor UO_880 (O_880,N_29288,N_29977);
nor UO_881 (O_881,N_28976,N_29726);
and UO_882 (O_882,N_28886,N_29670);
and UO_883 (O_883,N_29425,N_29178);
nand UO_884 (O_884,N_29379,N_29095);
xnor UO_885 (O_885,N_29648,N_29514);
or UO_886 (O_886,N_29155,N_29041);
nor UO_887 (O_887,N_28916,N_29461);
nor UO_888 (O_888,N_29039,N_29792);
or UO_889 (O_889,N_28846,N_29035);
nand UO_890 (O_890,N_29884,N_29514);
nand UO_891 (O_891,N_29538,N_29434);
nand UO_892 (O_892,N_29869,N_29752);
and UO_893 (O_893,N_29902,N_29362);
nand UO_894 (O_894,N_29270,N_29236);
or UO_895 (O_895,N_29262,N_29601);
and UO_896 (O_896,N_28992,N_29463);
nand UO_897 (O_897,N_29090,N_29897);
nand UO_898 (O_898,N_29905,N_28915);
xor UO_899 (O_899,N_28867,N_28812);
xnor UO_900 (O_900,N_29937,N_29645);
xor UO_901 (O_901,N_29325,N_29722);
xor UO_902 (O_902,N_29786,N_28897);
xor UO_903 (O_903,N_29021,N_29890);
nor UO_904 (O_904,N_29401,N_29467);
xnor UO_905 (O_905,N_29952,N_29695);
and UO_906 (O_906,N_29019,N_29466);
xnor UO_907 (O_907,N_29075,N_29449);
nand UO_908 (O_908,N_29646,N_29605);
xnor UO_909 (O_909,N_29815,N_29891);
nand UO_910 (O_910,N_29606,N_28988);
or UO_911 (O_911,N_28887,N_29198);
nor UO_912 (O_912,N_29251,N_28819);
nor UO_913 (O_913,N_29536,N_29648);
xor UO_914 (O_914,N_29375,N_29221);
and UO_915 (O_915,N_29071,N_28885);
nand UO_916 (O_916,N_29359,N_29924);
xor UO_917 (O_917,N_28988,N_29938);
and UO_918 (O_918,N_29245,N_29362);
and UO_919 (O_919,N_29098,N_29988);
or UO_920 (O_920,N_29861,N_29668);
and UO_921 (O_921,N_29052,N_29997);
and UO_922 (O_922,N_29009,N_29556);
nand UO_923 (O_923,N_28974,N_29615);
and UO_924 (O_924,N_29703,N_29818);
nor UO_925 (O_925,N_29953,N_29828);
and UO_926 (O_926,N_29893,N_29901);
or UO_927 (O_927,N_29700,N_28893);
and UO_928 (O_928,N_29366,N_29527);
nor UO_929 (O_929,N_29694,N_29711);
or UO_930 (O_930,N_29481,N_29927);
nand UO_931 (O_931,N_29113,N_28899);
nor UO_932 (O_932,N_29198,N_29452);
or UO_933 (O_933,N_29200,N_29189);
or UO_934 (O_934,N_29760,N_29461);
nand UO_935 (O_935,N_28897,N_28924);
nor UO_936 (O_936,N_29249,N_28868);
nor UO_937 (O_937,N_29981,N_29708);
xor UO_938 (O_938,N_29095,N_29145);
xnor UO_939 (O_939,N_29455,N_29079);
xor UO_940 (O_940,N_29945,N_29591);
and UO_941 (O_941,N_29802,N_29407);
xor UO_942 (O_942,N_29632,N_29082);
and UO_943 (O_943,N_28965,N_29424);
nand UO_944 (O_944,N_29159,N_29887);
xnor UO_945 (O_945,N_28944,N_29536);
and UO_946 (O_946,N_28833,N_29494);
or UO_947 (O_947,N_28906,N_29477);
nor UO_948 (O_948,N_29037,N_29036);
xnor UO_949 (O_949,N_28803,N_29690);
or UO_950 (O_950,N_29104,N_29475);
nand UO_951 (O_951,N_29893,N_28872);
nand UO_952 (O_952,N_29364,N_29795);
or UO_953 (O_953,N_28865,N_29597);
and UO_954 (O_954,N_29239,N_29051);
nor UO_955 (O_955,N_29533,N_29618);
and UO_956 (O_956,N_29108,N_28966);
nor UO_957 (O_957,N_29049,N_29449);
nor UO_958 (O_958,N_29868,N_29933);
or UO_959 (O_959,N_29731,N_29452);
nor UO_960 (O_960,N_29606,N_29699);
or UO_961 (O_961,N_29650,N_29631);
xnor UO_962 (O_962,N_29950,N_29265);
nand UO_963 (O_963,N_29409,N_29881);
nor UO_964 (O_964,N_29488,N_29470);
nor UO_965 (O_965,N_28997,N_28999);
xnor UO_966 (O_966,N_29585,N_29741);
or UO_967 (O_967,N_28813,N_28961);
nand UO_968 (O_968,N_29068,N_29720);
nor UO_969 (O_969,N_29000,N_29556);
or UO_970 (O_970,N_29195,N_29278);
and UO_971 (O_971,N_29576,N_29308);
nand UO_972 (O_972,N_28879,N_29454);
or UO_973 (O_973,N_28989,N_29085);
nand UO_974 (O_974,N_29960,N_29297);
xnor UO_975 (O_975,N_29998,N_29550);
and UO_976 (O_976,N_29587,N_29670);
nand UO_977 (O_977,N_29418,N_29454);
nand UO_978 (O_978,N_29308,N_28984);
and UO_979 (O_979,N_29401,N_29173);
and UO_980 (O_980,N_29412,N_29142);
nor UO_981 (O_981,N_28975,N_29314);
nand UO_982 (O_982,N_28828,N_29222);
nand UO_983 (O_983,N_28945,N_28981);
nor UO_984 (O_984,N_29437,N_29891);
nand UO_985 (O_985,N_29721,N_29616);
and UO_986 (O_986,N_29463,N_29324);
nor UO_987 (O_987,N_29627,N_29654);
nand UO_988 (O_988,N_29388,N_29248);
or UO_989 (O_989,N_29918,N_29425);
nand UO_990 (O_990,N_28931,N_29339);
nor UO_991 (O_991,N_29105,N_29983);
and UO_992 (O_992,N_29827,N_29977);
xor UO_993 (O_993,N_29992,N_28826);
and UO_994 (O_994,N_29041,N_29946);
or UO_995 (O_995,N_29739,N_29473);
and UO_996 (O_996,N_29416,N_29680);
or UO_997 (O_997,N_28891,N_28970);
xnor UO_998 (O_998,N_29869,N_29159);
nand UO_999 (O_999,N_29135,N_29868);
nor UO_1000 (O_1000,N_29682,N_29054);
xnor UO_1001 (O_1001,N_29605,N_29348);
nand UO_1002 (O_1002,N_29872,N_29319);
nand UO_1003 (O_1003,N_29584,N_28807);
nor UO_1004 (O_1004,N_28804,N_28969);
nand UO_1005 (O_1005,N_29419,N_28920);
and UO_1006 (O_1006,N_29484,N_29619);
and UO_1007 (O_1007,N_29847,N_29621);
xnor UO_1008 (O_1008,N_29720,N_29706);
and UO_1009 (O_1009,N_29252,N_28869);
nand UO_1010 (O_1010,N_28854,N_29984);
nand UO_1011 (O_1011,N_29289,N_29403);
and UO_1012 (O_1012,N_29754,N_29861);
xor UO_1013 (O_1013,N_29466,N_29725);
and UO_1014 (O_1014,N_29321,N_29730);
xor UO_1015 (O_1015,N_29542,N_29985);
and UO_1016 (O_1016,N_29354,N_29717);
nand UO_1017 (O_1017,N_29433,N_29424);
or UO_1018 (O_1018,N_29377,N_29174);
xor UO_1019 (O_1019,N_29032,N_29552);
xnor UO_1020 (O_1020,N_29851,N_29137);
nand UO_1021 (O_1021,N_29912,N_29976);
nand UO_1022 (O_1022,N_29244,N_29026);
xor UO_1023 (O_1023,N_29365,N_29301);
and UO_1024 (O_1024,N_29504,N_29943);
xnor UO_1025 (O_1025,N_29895,N_29758);
nand UO_1026 (O_1026,N_28984,N_29135);
nand UO_1027 (O_1027,N_29679,N_29996);
xor UO_1028 (O_1028,N_29327,N_28836);
or UO_1029 (O_1029,N_29242,N_29984);
nor UO_1030 (O_1030,N_29027,N_28939);
or UO_1031 (O_1031,N_29636,N_28871);
or UO_1032 (O_1032,N_29154,N_29217);
xnor UO_1033 (O_1033,N_29117,N_29491);
nor UO_1034 (O_1034,N_29402,N_29276);
nand UO_1035 (O_1035,N_28877,N_29863);
nand UO_1036 (O_1036,N_29031,N_29353);
or UO_1037 (O_1037,N_29216,N_28874);
nor UO_1038 (O_1038,N_29962,N_29742);
nor UO_1039 (O_1039,N_28969,N_29075);
xor UO_1040 (O_1040,N_29560,N_29077);
and UO_1041 (O_1041,N_28853,N_28918);
xnor UO_1042 (O_1042,N_29249,N_29055);
or UO_1043 (O_1043,N_29820,N_29072);
or UO_1044 (O_1044,N_29477,N_29983);
nor UO_1045 (O_1045,N_29881,N_29985);
nor UO_1046 (O_1046,N_29133,N_29636);
xor UO_1047 (O_1047,N_28862,N_28994);
nor UO_1048 (O_1048,N_28988,N_29505);
xor UO_1049 (O_1049,N_29464,N_29047);
and UO_1050 (O_1050,N_29516,N_28968);
nand UO_1051 (O_1051,N_29602,N_29859);
or UO_1052 (O_1052,N_29769,N_29740);
xor UO_1053 (O_1053,N_29825,N_28836);
nand UO_1054 (O_1054,N_29367,N_28800);
nor UO_1055 (O_1055,N_29665,N_29358);
nand UO_1056 (O_1056,N_29315,N_29734);
nor UO_1057 (O_1057,N_29281,N_29228);
or UO_1058 (O_1058,N_29816,N_28932);
nand UO_1059 (O_1059,N_29716,N_29185);
nand UO_1060 (O_1060,N_29406,N_29051);
xor UO_1061 (O_1061,N_29427,N_29215);
nor UO_1062 (O_1062,N_29934,N_28920);
xor UO_1063 (O_1063,N_29226,N_29323);
xnor UO_1064 (O_1064,N_28918,N_28996);
or UO_1065 (O_1065,N_29555,N_29535);
xor UO_1066 (O_1066,N_29096,N_29326);
or UO_1067 (O_1067,N_29965,N_29508);
nor UO_1068 (O_1068,N_29564,N_29131);
and UO_1069 (O_1069,N_29934,N_29172);
and UO_1070 (O_1070,N_29184,N_29434);
nor UO_1071 (O_1071,N_29886,N_29971);
nor UO_1072 (O_1072,N_29037,N_29886);
or UO_1073 (O_1073,N_28987,N_29538);
nand UO_1074 (O_1074,N_28914,N_29379);
nand UO_1075 (O_1075,N_29402,N_29560);
or UO_1076 (O_1076,N_29041,N_28851);
xnor UO_1077 (O_1077,N_29554,N_28896);
xor UO_1078 (O_1078,N_28887,N_29685);
nor UO_1079 (O_1079,N_29903,N_29141);
nor UO_1080 (O_1080,N_29813,N_29696);
and UO_1081 (O_1081,N_28831,N_29279);
xor UO_1082 (O_1082,N_29005,N_29333);
xnor UO_1083 (O_1083,N_29170,N_28971);
nand UO_1084 (O_1084,N_29164,N_29946);
and UO_1085 (O_1085,N_29424,N_29434);
or UO_1086 (O_1086,N_29926,N_29395);
nand UO_1087 (O_1087,N_29509,N_28986);
nand UO_1088 (O_1088,N_29973,N_29010);
and UO_1089 (O_1089,N_28921,N_28884);
nand UO_1090 (O_1090,N_28891,N_29981);
or UO_1091 (O_1091,N_29762,N_29689);
nand UO_1092 (O_1092,N_29666,N_29097);
nand UO_1093 (O_1093,N_29021,N_29804);
and UO_1094 (O_1094,N_29872,N_28956);
nand UO_1095 (O_1095,N_29037,N_29446);
xnor UO_1096 (O_1096,N_29792,N_29680);
and UO_1097 (O_1097,N_29979,N_29328);
nor UO_1098 (O_1098,N_29234,N_28916);
nand UO_1099 (O_1099,N_29388,N_29626);
nor UO_1100 (O_1100,N_29301,N_29792);
and UO_1101 (O_1101,N_29090,N_29676);
xnor UO_1102 (O_1102,N_28978,N_29562);
xnor UO_1103 (O_1103,N_29291,N_29703);
xor UO_1104 (O_1104,N_29571,N_28829);
xor UO_1105 (O_1105,N_29654,N_29132);
nand UO_1106 (O_1106,N_29420,N_28888);
and UO_1107 (O_1107,N_29512,N_29774);
or UO_1108 (O_1108,N_29163,N_29975);
nor UO_1109 (O_1109,N_29173,N_29704);
xnor UO_1110 (O_1110,N_29867,N_29341);
and UO_1111 (O_1111,N_28822,N_29445);
and UO_1112 (O_1112,N_29766,N_28879);
nand UO_1113 (O_1113,N_29296,N_29237);
nor UO_1114 (O_1114,N_29720,N_28988);
nor UO_1115 (O_1115,N_29287,N_29975);
nor UO_1116 (O_1116,N_29123,N_29758);
or UO_1117 (O_1117,N_29899,N_29363);
or UO_1118 (O_1118,N_28946,N_29752);
nor UO_1119 (O_1119,N_29321,N_29297);
xor UO_1120 (O_1120,N_29039,N_28811);
or UO_1121 (O_1121,N_29805,N_29201);
nor UO_1122 (O_1122,N_29838,N_29439);
and UO_1123 (O_1123,N_29721,N_29043);
and UO_1124 (O_1124,N_29852,N_29020);
nand UO_1125 (O_1125,N_29245,N_29633);
nand UO_1126 (O_1126,N_28921,N_29821);
xnor UO_1127 (O_1127,N_29261,N_29964);
and UO_1128 (O_1128,N_29118,N_29370);
xnor UO_1129 (O_1129,N_29403,N_29958);
nor UO_1130 (O_1130,N_29920,N_28929);
and UO_1131 (O_1131,N_29874,N_29883);
xor UO_1132 (O_1132,N_29751,N_28830);
and UO_1133 (O_1133,N_29468,N_29332);
nand UO_1134 (O_1134,N_29272,N_29354);
xnor UO_1135 (O_1135,N_29935,N_29928);
nand UO_1136 (O_1136,N_29663,N_29336);
and UO_1137 (O_1137,N_29894,N_28970);
xnor UO_1138 (O_1138,N_29412,N_28909);
and UO_1139 (O_1139,N_28802,N_29858);
or UO_1140 (O_1140,N_29728,N_29903);
and UO_1141 (O_1141,N_28863,N_29468);
nor UO_1142 (O_1142,N_29987,N_29244);
or UO_1143 (O_1143,N_29745,N_29264);
xor UO_1144 (O_1144,N_29528,N_29158);
xor UO_1145 (O_1145,N_29513,N_29271);
nor UO_1146 (O_1146,N_29035,N_29738);
and UO_1147 (O_1147,N_28945,N_29631);
nand UO_1148 (O_1148,N_28870,N_28895);
xnor UO_1149 (O_1149,N_29596,N_29778);
xnor UO_1150 (O_1150,N_28879,N_29547);
nand UO_1151 (O_1151,N_29644,N_28935);
nand UO_1152 (O_1152,N_29183,N_29908);
xnor UO_1153 (O_1153,N_29628,N_29664);
or UO_1154 (O_1154,N_29113,N_28844);
xnor UO_1155 (O_1155,N_28825,N_29299);
xor UO_1156 (O_1156,N_29239,N_29711);
and UO_1157 (O_1157,N_29648,N_29073);
nand UO_1158 (O_1158,N_29601,N_29440);
nor UO_1159 (O_1159,N_29809,N_29902);
nor UO_1160 (O_1160,N_29241,N_29216);
and UO_1161 (O_1161,N_29255,N_29189);
and UO_1162 (O_1162,N_28836,N_29004);
nor UO_1163 (O_1163,N_29510,N_29802);
nand UO_1164 (O_1164,N_29040,N_28965);
nand UO_1165 (O_1165,N_28945,N_29520);
and UO_1166 (O_1166,N_29709,N_29103);
and UO_1167 (O_1167,N_29853,N_28965);
nor UO_1168 (O_1168,N_29214,N_29471);
nor UO_1169 (O_1169,N_29501,N_28814);
nor UO_1170 (O_1170,N_29709,N_28840);
xnor UO_1171 (O_1171,N_29765,N_29192);
or UO_1172 (O_1172,N_29600,N_29165);
or UO_1173 (O_1173,N_29617,N_29593);
nand UO_1174 (O_1174,N_29322,N_28907);
or UO_1175 (O_1175,N_29031,N_29213);
or UO_1176 (O_1176,N_29033,N_29646);
xor UO_1177 (O_1177,N_29239,N_29742);
and UO_1178 (O_1178,N_29181,N_29733);
xor UO_1179 (O_1179,N_29187,N_28806);
and UO_1180 (O_1180,N_29149,N_29132);
nand UO_1181 (O_1181,N_29887,N_29829);
or UO_1182 (O_1182,N_29703,N_29491);
or UO_1183 (O_1183,N_29513,N_29701);
nand UO_1184 (O_1184,N_29460,N_28990);
xor UO_1185 (O_1185,N_29555,N_29385);
xnor UO_1186 (O_1186,N_29403,N_29575);
or UO_1187 (O_1187,N_29197,N_29441);
and UO_1188 (O_1188,N_28922,N_29651);
nand UO_1189 (O_1189,N_28977,N_29063);
nor UO_1190 (O_1190,N_29077,N_28945);
or UO_1191 (O_1191,N_29257,N_28857);
or UO_1192 (O_1192,N_29998,N_29104);
or UO_1193 (O_1193,N_29133,N_29458);
nand UO_1194 (O_1194,N_28848,N_29869);
nand UO_1195 (O_1195,N_29830,N_29912);
and UO_1196 (O_1196,N_29335,N_29385);
or UO_1197 (O_1197,N_29173,N_29051);
nor UO_1198 (O_1198,N_29971,N_28852);
xnor UO_1199 (O_1199,N_29122,N_29899);
nor UO_1200 (O_1200,N_29594,N_29623);
nor UO_1201 (O_1201,N_29746,N_29605);
nor UO_1202 (O_1202,N_29844,N_29804);
nand UO_1203 (O_1203,N_29229,N_29980);
nand UO_1204 (O_1204,N_29117,N_28870);
xnor UO_1205 (O_1205,N_29586,N_29538);
nor UO_1206 (O_1206,N_29728,N_29687);
nor UO_1207 (O_1207,N_29130,N_29013);
or UO_1208 (O_1208,N_29312,N_29362);
and UO_1209 (O_1209,N_29645,N_29414);
nand UO_1210 (O_1210,N_28823,N_29828);
nor UO_1211 (O_1211,N_29621,N_29688);
and UO_1212 (O_1212,N_28940,N_29528);
or UO_1213 (O_1213,N_29649,N_29645);
nor UO_1214 (O_1214,N_29413,N_29675);
and UO_1215 (O_1215,N_29654,N_29503);
and UO_1216 (O_1216,N_29831,N_29752);
nor UO_1217 (O_1217,N_29243,N_29803);
xnor UO_1218 (O_1218,N_29092,N_29565);
or UO_1219 (O_1219,N_28983,N_29868);
nand UO_1220 (O_1220,N_28903,N_29849);
xnor UO_1221 (O_1221,N_29800,N_29704);
xor UO_1222 (O_1222,N_29456,N_28877);
nor UO_1223 (O_1223,N_29997,N_29763);
and UO_1224 (O_1224,N_29562,N_28992);
nor UO_1225 (O_1225,N_29344,N_28890);
nand UO_1226 (O_1226,N_29170,N_29262);
nor UO_1227 (O_1227,N_29652,N_29309);
or UO_1228 (O_1228,N_29596,N_29626);
or UO_1229 (O_1229,N_29780,N_29927);
and UO_1230 (O_1230,N_29266,N_29185);
nand UO_1231 (O_1231,N_29093,N_29046);
or UO_1232 (O_1232,N_29612,N_29908);
xnor UO_1233 (O_1233,N_29694,N_29974);
nand UO_1234 (O_1234,N_29570,N_29483);
nor UO_1235 (O_1235,N_29496,N_29638);
nand UO_1236 (O_1236,N_29068,N_29713);
nor UO_1237 (O_1237,N_29387,N_29877);
xnor UO_1238 (O_1238,N_29098,N_29934);
nor UO_1239 (O_1239,N_29605,N_29157);
and UO_1240 (O_1240,N_29634,N_29388);
or UO_1241 (O_1241,N_28861,N_28891);
or UO_1242 (O_1242,N_29897,N_29610);
nor UO_1243 (O_1243,N_28891,N_29581);
nor UO_1244 (O_1244,N_29902,N_29095);
and UO_1245 (O_1245,N_28861,N_29083);
and UO_1246 (O_1246,N_28960,N_29991);
or UO_1247 (O_1247,N_29954,N_29230);
nor UO_1248 (O_1248,N_29887,N_29589);
nor UO_1249 (O_1249,N_29113,N_29778);
nor UO_1250 (O_1250,N_29263,N_29619);
and UO_1251 (O_1251,N_29922,N_28844);
xnor UO_1252 (O_1252,N_28900,N_29826);
nor UO_1253 (O_1253,N_29759,N_28859);
nor UO_1254 (O_1254,N_29231,N_29254);
xnor UO_1255 (O_1255,N_28825,N_29333);
nor UO_1256 (O_1256,N_29976,N_29088);
or UO_1257 (O_1257,N_29507,N_29008);
nand UO_1258 (O_1258,N_29596,N_29839);
and UO_1259 (O_1259,N_29594,N_29352);
nand UO_1260 (O_1260,N_29194,N_28921);
nand UO_1261 (O_1261,N_29066,N_29378);
or UO_1262 (O_1262,N_29115,N_29175);
nor UO_1263 (O_1263,N_29220,N_29488);
and UO_1264 (O_1264,N_28816,N_28859);
and UO_1265 (O_1265,N_29585,N_29045);
nor UO_1266 (O_1266,N_29138,N_29818);
nand UO_1267 (O_1267,N_28983,N_29003);
and UO_1268 (O_1268,N_29588,N_29010);
nor UO_1269 (O_1269,N_29297,N_29293);
and UO_1270 (O_1270,N_29171,N_29910);
and UO_1271 (O_1271,N_29355,N_29247);
and UO_1272 (O_1272,N_29218,N_29847);
and UO_1273 (O_1273,N_29561,N_28841);
nand UO_1274 (O_1274,N_29989,N_29316);
and UO_1275 (O_1275,N_29789,N_29101);
and UO_1276 (O_1276,N_29930,N_28992);
and UO_1277 (O_1277,N_29909,N_29389);
or UO_1278 (O_1278,N_28802,N_28989);
nand UO_1279 (O_1279,N_29720,N_29719);
nor UO_1280 (O_1280,N_29350,N_29471);
and UO_1281 (O_1281,N_29944,N_29191);
xnor UO_1282 (O_1282,N_29039,N_28916);
and UO_1283 (O_1283,N_28954,N_29295);
xnor UO_1284 (O_1284,N_29047,N_29370);
or UO_1285 (O_1285,N_28823,N_29485);
nor UO_1286 (O_1286,N_29896,N_29065);
or UO_1287 (O_1287,N_29552,N_29922);
and UO_1288 (O_1288,N_29624,N_29173);
and UO_1289 (O_1289,N_29597,N_29831);
and UO_1290 (O_1290,N_28832,N_29394);
nand UO_1291 (O_1291,N_29683,N_29026);
xnor UO_1292 (O_1292,N_29561,N_29030);
xnor UO_1293 (O_1293,N_29963,N_29785);
or UO_1294 (O_1294,N_29196,N_29958);
or UO_1295 (O_1295,N_29366,N_29628);
or UO_1296 (O_1296,N_29054,N_28823);
nor UO_1297 (O_1297,N_29257,N_29584);
or UO_1298 (O_1298,N_29780,N_29943);
xor UO_1299 (O_1299,N_29121,N_29153);
nor UO_1300 (O_1300,N_29859,N_29451);
and UO_1301 (O_1301,N_29505,N_28838);
nand UO_1302 (O_1302,N_29602,N_28800);
or UO_1303 (O_1303,N_29344,N_29861);
nand UO_1304 (O_1304,N_29911,N_29916);
or UO_1305 (O_1305,N_29450,N_29421);
nand UO_1306 (O_1306,N_29031,N_28854);
nand UO_1307 (O_1307,N_29554,N_29679);
xnor UO_1308 (O_1308,N_29625,N_29139);
and UO_1309 (O_1309,N_29051,N_29515);
or UO_1310 (O_1310,N_29835,N_29879);
or UO_1311 (O_1311,N_28958,N_29289);
or UO_1312 (O_1312,N_29089,N_29013);
or UO_1313 (O_1313,N_29568,N_29064);
nor UO_1314 (O_1314,N_29028,N_29826);
and UO_1315 (O_1315,N_29879,N_29758);
nand UO_1316 (O_1316,N_29973,N_29975);
and UO_1317 (O_1317,N_29930,N_29816);
nand UO_1318 (O_1318,N_28874,N_29365);
nor UO_1319 (O_1319,N_29044,N_29041);
and UO_1320 (O_1320,N_29530,N_29383);
or UO_1321 (O_1321,N_28873,N_29665);
or UO_1322 (O_1322,N_28934,N_29561);
xnor UO_1323 (O_1323,N_29690,N_29935);
or UO_1324 (O_1324,N_29548,N_29498);
nand UO_1325 (O_1325,N_29533,N_29957);
nand UO_1326 (O_1326,N_28963,N_29405);
xor UO_1327 (O_1327,N_29278,N_29486);
and UO_1328 (O_1328,N_28969,N_28888);
xor UO_1329 (O_1329,N_29000,N_29191);
nor UO_1330 (O_1330,N_29258,N_29102);
nor UO_1331 (O_1331,N_29786,N_28963);
or UO_1332 (O_1332,N_29844,N_29786);
xor UO_1333 (O_1333,N_29600,N_29533);
xor UO_1334 (O_1334,N_29111,N_28904);
xnor UO_1335 (O_1335,N_29766,N_28844);
and UO_1336 (O_1336,N_29898,N_29555);
nand UO_1337 (O_1337,N_29322,N_29336);
or UO_1338 (O_1338,N_29284,N_29573);
xor UO_1339 (O_1339,N_29552,N_28812);
and UO_1340 (O_1340,N_29477,N_29219);
and UO_1341 (O_1341,N_29700,N_29788);
or UO_1342 (O_1342,N_29649,N_29625);
nor UO_1343 (O_1343,N_28951,N_29790);
xnor UO_1344 (O_1344,N_29363,N_29115);
nand UO_1345 (O_1345,N_29675,N_29861);
nand UO_1346 (O_1346,N_29114,N_29522);
or UO_1347 (O_1347,N_29101,N_28985);
nand UO_1348 (O_1348,N_29674,N_29806);
nor UO_1349 (O_1349,N_29254,N_28856);
nor UO_1350 (O_1350,N_28902,N_28985);
xnor UO_1351 (O_1351,N_28929,N_29850);
nand UO_1352 (O_1352,N_29310,N_29050);
nand UO_1353 (O_1353,N_29011,N_29086);
xnor UO_1354 (O_1354,N_29290,N_28817);
xor UO_1355 (O_1355,N_29034,N_28879);
or UO_1356 (O_1356,N_29417,N_29231);
xor UO_1357 (O_1357,N_29396,N_29592);
xor UO_1358 (O_1358,N_29861,N_29798);
and UO_1359 (O_1359,N_29748,N_29489);
and UO_1360 (O_1360,N_29419,N_28828);
nand UO_1361 (O_1361,N_29317,N_29800);
or UO_1362 (O_1362,N_29820,N_28991);
xor UO_1363 (O_1363,N_29933,N_29987);
or UO_1364 (O_1364,N_29431,N_29962);
or UO_1365 (O_1365,N_29171,N_29157);
or UO_1366 (O_1366,N_29646,N_29015);
xor UO_1367 (O_1367,N_29341,N_29010);
nor UO_1368 (O_1368,N_29490,N_29983);
or UO_1369 (O_1369,N_29664,N_29549);
or UO_1370 (O_1370,N_29583,N_29234);
xnor UO_1371 (O_1371,N_29934,N_29721);
and UO_1372 (O_1372,N_29720,N_28823);
nand UO_1373 (O_1373,N_29950,N_29538);
or UO_1374 (O_1374,N_29456,N_29960);
nor UO_1375 (O_1375,N_29653,N_28937);
or UO_1376 (O_1376,N_29754,N_29230);
nand UO_1377 (O_1377,N_29093,N_29095);
xnor UO_1378 (O_1378,N_29502,N_29533);
nor UO_1379 (O_1379,N_28857,N_29283);
xnor UO_1380 (O_1380,N_29941,N_29011);
nor UO_1381 (O_1381,N_29553,N_29276);
nand UO_1382 (O_1382,N_29049,N_29967);
nor UO_1383 (O_1383,N_29399,N_29152);
nand UO_1384 (O_1384,N_29114,N_29083);
nor UO_1385 (O_1385,N_29783,N_29978);
and UO_1386 (O_1386,N_29868,N_28810);
xnor UO_1387 (O_1387,N_29073,N_29596);
and UO_1388 (O_1388,N_28948,N_29166);
nor UO_1389 (O_1389,N_29653,N_29534);
nor UO_1390 (O_1390,N_29260,N_29054);
nand UO_1391 (O_1391,N_29857,N_29333);
nand UO_1392 (O_1392,N_29010,N_28809);
and UO_1393 (O_1393,N_29611,N_29104);
and UO_1394 (O_1394,N_29208,N_29752);
or UO_1395 (O_1395,N_29310,N_29108);
nand UO_1396 (O_1396,N_29462,N_29937);
nor UO_1397 (O_1397,N_28815,N_29679);
or UO_1398 (O_1398,N_29691,N_29305);
or UO_1399 (O_1399,N_29271,N_29076);
xnor UO_1400 (O_1400,N_28997,N_29796);
or UO_1401 (O_1401,N_29290,N_29998);
xnor UO_1402 (O_1402,N_29416,N_29926);
and UO_1403 (O_1403,N_29088,N_29008);
or UO_1404 (O_1404,N_28899,N_29599);
or UO_1405 (O_1405,N_29814,N_29958);
xor UO_1406 (O_1406,N_29520,N_29452);
or UO_1407 (O_1407,N_28878,N_29881);
or UO_1408 (O_1408,N_29685,N_28959);
xnor UO_1409 (O_1409,N_29923,N_29232);
nor UO_1410 (O_1410,N_29664,N_29068);
nor UO_1411 (O_1411,N_28892,N_28916);
and UO_1412 (O_1412,N_29771,N_29674);
xor UO_1413 (O_1413,N_29434,N_29603);
xnor UO_1414 (O_1414,N_29112,N_29854);
nor UO_1415 (O_1415,N_29861,N_29118);
xnor UO_1416 (O_1416,N_29592,N_29310);
xnor UO_1417 (O_1417,N_29155,N_28998);
xnor UO_1418 (O_1418,N_28952,N_29734);
xnor UO_1419 (O_1419,N_29990,N_29480);
and UO_1420 (O_1420,N_29697,N_29628);
and UO_1421 (O_1421,N_28863,N_29220);
xnor UO_1422 (O_1422,N_29116,N_29761);
nor UO_1423 (O_1423,N_28924,N_28980);
and UO_1424 (O_1424,N_28858,N_29003);
and UO_1425 (O_1425,N_29663,N_28931);
nor UO_1426 (O_1426,N_29931,N_29342);
nor UO_1427 (O_1427,N_29448,N_29435);
nand UO_1428 (O_1428,N_28960,N_29827);
nand UO_1429 (O_1429,N_29462,N_29911);
xor UO_1430 (O_1430,N_29211,N_29748);
and UO_1431 (O_1431,N_29615,N_29642);
or UO_1432 (O_1432,N_29488,N_29161);
or UO_1433 (O_1433,N_29615,N_29653);
and UO_1434 (O_1434,N_29123,N_29342);
xnor UO_1435 (O_1435,N_29796,N_29609);
and UO_1436 (O_1436,N_29415,N_29280);
or UO_1437 (O_1437,N_29884,N_29522);
xnor UO_1438 (O_1438,N_29485,N_29159);
xor UO_1439 (O_1439,N_28890,N_29480);
or UO_1440 (O_1440,N_28864,N_29928);
nor UO_1441 (O_1441,N_29247,N_29248);
xor UO_1442 (O_1442,N_29481,N_28848);
or UO_1443 (O_1443,N_29843,N_29444);
nor UO_1444 (O_1444,N_29915,N_28964);
nand UO_1445 (O_1445,N_29833,N_29720);
or UO_1446 (O_1446,N_29837,N_28866);
xnor UO_1447 (O_1447,N_29519,N_28988);
nand UO_1448 (O_1448,N_29691,N_29469);
nor UO_1449 (O_1449,N_28829,N_29009);
and UO_1450 (O_1450,N_29610,N_29165);
and UO_1451 (O_1451,N_28873,N_29087);
and UO_1452 (O_1452,N_29523,N_29276);
or UO_1453 (O_1453,N_29063,N_29778);
or UO_1454 (O_1454,N_29586,N_29924);
nor UO_1455 (O_1455,N_29773,N_29804);
or UO_1456 (O_1456,N_28899,N_29742);
and UO_1457 (O_1457,N_28900,N_29785);
and UO_1458 (O_1458,N_29447,N_29920);
nor UO_1459 (O_1459,N_29333,N_29454);
and UO_1460 (O_1460,N_29309,N_29784);
nand UO_1461 (O_1461,N_28829,N_29537);
xnor UO_1462 (O_1462,N_28812,N_29163);
nor UO_1463 (O_1463,N_29908,N_29990);
xor UO_1464 (O_1464,N_28901,N_29829);
nand UO_1465 (O_1465,N_29959,N_29483);
nand UO_1466 (O_1466,N_29474,N_29177);
and UO_1467 (O_1467,N_29198,N_29925);
and UO_1468 (O_1468,N_29279,N_29762);
or UO_1469 (O_1469,N_29300,N_28993);
nor UO_1470 (O_1470,N_29206,N_29454);
nor UO_1471 (O_1471,N_29973,N_29878);
nand UO_1472 (O_1472,N_29510,N_29353);
nand UO_1473 (O_1473,N_29310,N_29952);
xnor UO_1474 (O_1474,N_29940,N_29668);
or UO_1475 (O_1475,N_29126,N_29063);
and UO_1476 (O_1476,N_29295,N_29185);
or UO_1477 (O_1477,N_29211,N_29619);
or UO_1478 (O_1478,N_29317,N_28884);
nor UO_1479 (O_1479,N_29333,N_28867);
and UO_1480 (O_1480,N_29727,N_29630);
or UO_1481 (O_1481,N_29027,N_29161);
xor UO_1482 (O_1482,N_29045,N_28882);
and UO_1483 (O_1483,N_29066,N_29517);
and UO_1484 (O_1484,N_29246,N_28989);
and UO_1485 (O_1485,N_29340,N_28924);
xnor UO_1486 (O_1486,N_29718,N_29466);
nor UO_1487 (O_1487,N_29824,N_28870);
or UO_1488 (O_1488,N_29482,N_29304);
and UO_1489 (O_1489,N_29077,N_29456);
or UO_1490 (O_1490,N_29094,N_29490);
nor UO_1491 (O_1491,N_29417,N_29727);
and UO_1492 (O_1492,N_28866,N_29683);
or UO_1493 (O_1493,N_29154,N_29570);
xnor UO_1494 (O_1494,N_28942,N_29234);
nor UO_1495 (O_1495,N_29786,N_29184);
and UO_1496 (O_1496,N_29682,N_29598);
or UO_1497 (O_1497,N_29570,N_28950);
and UO_1498 (O_1498,N_28954,N_29568);
xor UO_1499 (O_1499,N_29686,N_29805);
or UO_1500 (O_1500,N_29579,N_29260);
xnor UO_1501 (O_1501,N_29733,N_29594);
or UO_1502 (O_1502,N_29967,N_29968);
nand UO_1503 (O_1503,N_28983,N_29447);
or UO_1504 (O_1504,N_29168,N_29767);
nand UO_1505 (O_1505,N_29165,N_29659);
nand UO_1506 (O_1506,N_28968,N_28936);
xnor UO_1507 (O_1507,N_29125,N_29740);
or UO_1508 (O_1508,N_28851,N_28974);
or UO_1509 (O_1509,N_29096,N_29274);
nand UO_1510 (O_1510,N_28905,N_29604);
and UO_1511 (O_1511,N_28880,N_28817);
nand UO_1512 (O_1512,N_29647,N_29453);
nor UO_1513 (O_1513,N_29159,N_29933);
xnor UO_1514 (O_1514,N_29400,N_28833);
nor UO_1515 (O_1515,N_29653,N_29096);
or UO_1516 (O_1516,N_29155,N_29567);
xnor UO_1517 (O_1517,N_29377,N_29161);
nand UO_1518 (O_1518,N_28838,N_29602);
and UO_1519 (O_1519,N_29738,N_29847);
nand UO_1520 (O_1520,N_29952,N_29820);
nand UO_1521 (O_1521,N_29249,N_29614);
or UO_1522 (O_1522,N_29776,N_28853);
or UO_1523 (O_1523,N_28979,N_29040);
or UO_1524 (O_1524,N_29300,N_29493);
xnor UO_1525 (O_1525,N_29581,N_28940);
xnor UO_1526 (O_1526,N_28979,N_29684);
or UO_1527 (O_1527,N_29349,N_28809);
xor UO_1528 (O_1528,N_29931,N_28940);
and UO_1529 (O_1529,N_29061,N_28975);
nand UO_1530 (O_1530,N_29508,N_29437);
nand UO_1531 (O_1531,N_29008,N_29127);
and UO_1532 (O_1532,N_29626,N_29691);
nand UO_1533 (O_1533,N_29471,N_29424);
and UO_1534 (O_1534,N_28994,N_29045);
nor UO_1535 (O_1535,N_29712,N_29516);
xnor UO_1536 (O_1536,N_29568,N_29453);
or UO_1537 (O_1537,N_29036,N_29065);
or UO_1538 (O_1538,N_29282,N_29258);
or UO_1539 (O_1539,N_28900,N_29254);
xor UO_1540 (O_1540,N_29935,N_28887);
and UO_1541 (O_1541,N_29815,N_29830);
or UO_1542 (O_1542,N_29778,N_29763);
or UO_1543 (O_1543,N_29896,N_29808);
nand UO_1544 (O_1544,N_29059,N_29940);
xnor UO_1545 (O_1545,N_29387,N_29235);
or UO_1546 (O_1546,N_29963,N_29433);
or UO_1547 (O_1547,N_29023,N_28866);
and UO_1548 (O_1548,N_29338,N_29162);
nor UO_1549 (O_1549,N_29557,N_29400);
xnor UO_1550 (O_1550,N_29654,N_29482);
nand UO_1551 (O_1551,N_29617,N_29279);
xnor UO_1552 (O_1552,N_28922,N_29128);
nor UO_1553 (O_1553,N_28891,N_28905);
or UO_1554 (O_1554,N_29158,N_29116);
or UO_1555 (O_1555,N_29075,N_28924);
or UO_1556 (O_1556,N_29178,N_29703);
or UO_1557 (O_1557,N_29400,N_29802);
nand UO_1558 (O_1558,N_29343,N_29555);
nand UO_1559 (O_1559,N_28826,N_28946);
and UO_1560 (O_1560,N_28989,N_29680);
nor UO_1561 (O_1561,N_29514,N_29682);
nand UO_1562 (O_1562,N_29513,N_28910);
or UO_1563 (O_1563,N_29768,N_28801);
nor UO_1564 (O_1564,N_29264,N_29956);
nand UO_1565 (O_1565,N_29059,N_29342);
and UO_1566 (O_1566,N_29688,N_29086);
and UO_1567 (O_1567,N_28881,N_29657);
or UO_1568 (O_1568,N_29474,N_29685);
xor UO_1569 (O_1569,N_29104,N_29113);
xor UO_1570 (O_1570,N_29781,N_29307);
and UO_1571 (O_1571,N_29855,N_29141);
nand UO_1572 (O_1572,N_29773,N_29952);
xor UO_1573 (O_1573,N_29173,N_28821);
or UO_1574 (O_1574,N_29556,N_29177);
and UO_1575 (O_1575,N_29029,N_29980);
nor UO_1576 (O_1576,N_29338,N_29055);
and UO_1577 (O_1577,N_29571,N_29118);
nand UO_1578 (O_1578,N_29406,N_29350);
nand UO_1579 (O_1579,N_29729,N_29612);
xor UO_1580 (O_1580,N_28956,N_29381);
nand UO_1581 (O_1581,N_29767,N_29900);
or UO_1582 (O_1582,N_29708,N_29812);
xor UO_1583 (O_1583,N_29985,N_29394);
or UO_1584 (O_1584,N_29014,N_29636);
nand UO_1585 (O_1585,N_29455,N_29519);
xor UO_1586 (O_1586,N_28822,N_29061);
or UO_1587 (O_1587,N_28880,N_29785);
or UO_1588 (O_1588,N_29577,N_29948);
and UO_1589 (O_1589,N_29972,N_29906);
nand UO_1590 (O_1590,N_28885,N_29727);
nor UO_1591 (O_1591,N_29531,N_28994);
and UO_1592 (O_1592,N_29799,N_29968);
and UO_1593 (O_1593,N_29466,N_29302);
nand UO_1594 (O_1594,N_28984,N_28979);
nor UO_1595 (O_1595,N_29164,N_29829);
xnor UO_1596 (O_1596,N_29794,N_28947);
xnor UO_1597 (O_1597,N_29440,N_28926);
nor UO_1598 (O_1598,N_29340,N_29278);
and UO_1599 (O_1599,N_29588,N_29590);
or UO_1600 (O_1600,N_29692,N_29433);
or UO_1601 (O_1601,N_29319,N_29927);
xnor UO_1602 (O_1602,N_29581,N_28982);
xor UO_1603 (O_1603,N_29618,N_28800);
nand UO_1604 (O_1604,N_29918,N_29545);
nor UO_1605 (O_1605,N_29269,N_28857);
xnor UO_1606 (O_1606,N_29684,N_29824);
xor UO_1607 (O_1607,N_29698,N_29432);
and UO_1608 (O_1608,N_28988,N_28936);
and UO_1609 (O_1609,N_29336,N_29525);
xnor UO_1610 (O_1610,N_29272,N_28808);
nor UO_1611 (O_1611,N_29405,N_29245);
or UO_1612 (O_1612,N_29482,N_29193);
nand UO_1613 (O_1613,N_29364,N_28894);
or UO_1614 (O_1614,N_28807,N_29877);
or UO_1615 (O_1615,N_28846,N_28965);
nor UO_1616 (O_1616,N_29540,N_29117);
and UO_1617 (O_1617,N_29370,N_28845);
nand UO_1618 (O_1618,N_29645,N_29237);
or UO_1619 (O_1619,N_29425,N_28980);
nor UO_1620 (O_1620,N_28809,N_29043);
nor UO_1621 (O_1621,N_29340,N_29398);
nand UO_1622 (O_1622,N_29228,N_29725);
and UO_1623 (O_1623,N_29423,N_28931);
nor UO_1624 (O_1624,N_29979,N_29135);
nor UO_1625 (O_1625,N_28886,N_29618);
xnor UO_1626 (O_1626,N_29554,N_28818);
nand UO_1627 (O_1627,N_29793,N_29613);
nand UO_1628 (O_1628,N_29052,N_29057);
or UO_1629 (O_1629,N_28989,N_29828);
or UO_1630 (O_1630,N_28907,N_29382);
xnor UO_1631 (O_1631,N_29965,N_29196);
nand UO_1632 (O_1632,N_29355,N_29083);
nand UO_1633 (O_1633,N_29621,N_28898);
or UO_1634 (O_1634,N_29320,N_29381);
xnor UO_1635 (O_1635,N_29529,N_29430);
xnor UO_1636 (O_1636,N_29253,N_28974);
nor UO_1637 (O_1637,N_29788,N_29224);
nor UO_1638 (O_1638,N_28949,N_29179);
or UO_1639 (O_1639,N_29912,N_29190);
and UO_1640 (O_1640,N_29280,N_29800);
and UO_1641 (O_1641,N_29860,N_29362);
or UO_1642 (O_1642,N_29757,N_29573);
and UO_1643 (O_1643,N_29290,N_29171);
xor UO_1644 (O_1644,N_29065,N_29685);
or UO_1645 (O_1645,N_29241,N_29122);
nor UO_1646 (O_1646,N_29804,N_29018);
nor UO_1647 (O_1647,N_29693,N_29638);
and UO_1648 (O_1648,N_29354,N_28993);
nand UO_1649 (O_1649,N_29171,N_29678);
xnor UO_1650 (O_1650,N_29661,N_29749);
xnor UO_1651 (O_1651,N_29385,N_29663);
nand UO_1652 (O_1652,N_29818,N_29201);
and UO_1653 (O_1653,N_29353,N_29928);
and UO_1654 (O_1654,N_29102,N_28969);
nor UO_1655 (O_1655,N_29267,N_29502);
nand UO_1656 (O_1656,N_29985,N_29377);
nand UO_1657 (O_1657,N_28822,N_29102);
xnor UO_1658 (O_1658,N_29878,N_28895);
and UO_1659 (O_1659,N_29856,N_29345);
nor UO_1660 (O_1660,N_29320,N_29159);
nand UO_1661 (O_1661,N_28894,N_29962);
or UO_1662 (O_1662,N_28954,N_29223);
nor UO_1663 (O_1663,N_29998,N_29689);
and UO_1664 (O_1664,N_29273,N_28837);
nor UO_1665 (O_1665,N_29960,N_29391);
nand UO_1666 (O_1666,N_29301,N_28874);
nand UO_1667 (O_1667,N_29388,N_29829);
nand UO_1668 (O_1668,N_29420,N_29017);
nor UO_1669 (O_1669,N_29913,N_29255);
nor UO_1670 (O_1670,N_29158,N_29704);
xor UO_1671 (O_1671,N_29639,N_29687);
and UO_1672 (O_1672,N_28920,N_29495);
or UO_1673 (O_1673,N_29786,N_28939);
nand UO_1674 (O_1674,N_28860,N_29845);
nor UO_1675 (O_1675,N_29164,N_28964);
or UO_1676 (O_1676,N_29023,N_29906);
nor UO_1677 (O_1677,N_28958,N_29281);
xor UO_1678 (O_1678,N_29981,N_29951);
nor UO_1679 (O_1679,N_29885,N_29908);
xor UO_1680 (O_1680,N_29501,N_28820);
and UO_1681 (O_1681,N_29643,N_29194);
or UO_1682 (O_1682,N_29173,N_28841);
nand UO_1683 (O_1683,N_29969,N_28955);
nand UO_1684 (O_1684,N_28857,N_29615);
and UO_1685 (O_1685,N_29019,N_29654);
nor UO_1686 (O_1686,N_29905,N_29399);
nand UO_1687 (O_1687,N_29045,N_29645);
or UO_1688 (O_1688,N_29973,N_29381);
nand UO_1689 (O_1689,N_29602,N_28851);
nand UO_1690 (O_1690,N_29880,N_28981);
or UO_1691 (O_1691,N_29524,N_29211);
nor UO_1692 (O_1692,N_28871,N_29306);
and UO_1693 (O_1693,N_29961,N_29451);
nor UO_1694 (O_1694,N_29158,N_29046);
nor UO_1695 (O_1695,N_29010,N_29353);
nor UO_1696 (O_1696,N_29215,N_29918);
or UO_1697 (O_1697,N_29613,N_29504);
nor UO_1698 (O_1698,N_28936,N_29134);
xnor UO_1699 (O_1699,N_29111,N_29202);
nand UO_1700 (O_1700,N_29501,N_29687);
xor UO_1701 (O_1701,N_29864,N_29882);
and UO_1702 (O_1702,N_29204,N_29987);
and UO_1703 (O_1703,N_29837,N_29348);
nor UO_1704 (O_1704,N_29675,N_29672);
and UO_1705 (O_1705,N_29028,N_29356);
and UO_1706 (O_1706,N_29494,N_29933);
or UO_1707 (O_1707,N_29862,N_29192);
xnor UO_1708 (O_1708,N_28991,N_29763);
nand UO_1709 (O_1709,N_28995,N_29071);
and UO_1710 (O_1710,N_29066,N_29564);
and UO_1711 (O_1711,N_29591,N_28914);
nor UO_1712 (O_1712,N_29613,N_28899);
nand UO_1713 (O_1713,N_29529,N_29022);
nor UO_1714 (O_1714,N_29544,N_29012);
nor UO_1715 (O_1715,N_28838,N_28997);
nand UO_1716 (O_1716,N_29424,N_29831);
nand UO_1717 (O_1717,N_29696,N_29901);
and UO_1718 (O_1718,N_29192,N_28857);
and UO_1719 (O_1719,N_29903,N_29268);
xor UO_1720 (O_1720,N_29500,N_29360);
xor UO_1721 (O_1721,N_28961,N_29905);
nand UO_1722 (O_1722,N_28862,N_29329);
and UO_1723 (O_1723,N_29420,N_29541);
xor UO_1724 (O_1724,N_28917,N_29271);
nor UO_1725 (O_1725,N_29978,N_29620);
nand UO_1726 (O_1726,N_29098,N_29011);
and UO_1727 (O_1727,N_29556,N_29783);
xor UO_1728 (O_1728,N_29425,N_29139);
or UO_1729 (O_1729,N_29572,N_29064);
nor UO_1730 (O_1730,N_28914,N_29066);
or UO_1731 (O_1731,N_29210,N_29409);
and UO_1732 (O_1732,N_29477,N_29369);
nor UO_1733 (O_1733,N_29260,N_29197);
nand UO_1734 (O_1734,N_29215,N_29279);
nand UO_1735 (O_1735,N_29688,N_29473);
and UO_1736 (O_1736,N_29688,N_29357);
or UO_1737 (O_1737,N_29356,N_29944);
or UO_1738 (O_1738,N_28884,N_29739);
or UO_1739 (O_1739,N_29256,N_29957);
nand UO_1740 (O_1740,N_29289,N_29199);
nor UO_1741 (O_1741,N_28908,N_29416);
and UO_1742 (O_1742,N_28846,N_28861);
and UO_1743 (O_1743,N_29277,N_29748);
nand UO_1744 (O_1744,N_29273,N_28820);
nand UO_1745 (O_1745,N_29579,N_29801);
nand UO_1746 (O_1746,N_29651,N_28803);
nand UO_1747 (O_1747,N_29278,N_29459);
or UO_1748 (O_1748,N_29635,N_29888);
nand UO_1749 (O_1749,N_28988,N_28989);
or UO_1750 (O_1750,N_29644,N_29275);
nand UO_1751 (O_1751,N_29375,N_29518);
nor UO_1752 (O_1752,N_29310,N_29931);
or UO_1753 (O_1753,N_29778,N_28906);
and UO_1754 (O_1754,N_29316,N_29958);
or UO_1755 (O_1755,N_29483,N_28931);
and UO_1756 (O_1756,N_29807,N_29865);
nand UO_1757 (O_1757,N_29765,N_29504);
xnor UO_1758 (O_1758,N_29777,N_29832);
nor UO_1759 (O_1759,N_29956,N_28973);
xnor UO_1760 (O_1760,N_29725,N_29254);
nor UO_1761 (O_1761,N_29386,N_28975);
and UO_1762 (O_1762,N_29992,N_29711);
or UO_1763 (O_1763,N_29661,N_29662);
or UO_1764 (O_1764,N_29617,N_29950);
nor UO_1765 (O_1765,N_29404,N_28838);
nor UO_1766 (O_1766,N_29718,N_29773);
nand UO_1767 (O_1767,N_29246,N_29780);
nand UO_1768 (O_1768,N_28865,N_28978);
nand UO_1769 (O_1769,N_29372,N_29566);
nor UO_1770 (O_1770,N_29972,N_29221);
nor UO_1771 (O_1771,N_29839,N_29385);
nand UO_1772 (O_1772,N_29954,N_29488);
nand UO_1773 (O_1773,N_28872,N_29618);
nor UO_1774 (O_1774,N_29100,N_29848);
xor UO_1775 (O_1775,N_29161,N_29740);
nor UO_1776 (O_1776,N_29031,N_29101);
nor UO_1777 (O_1777,N_29520,N_29113);
and UO_1778 (O_1778,N_29051,N_29391);
and UO_1779 (O_1779,N_29749,N_29924);
nor UO_1780 (O_1780,N_29649,N_29413);
nand UO_1781 (O_1781,N_29733,N_29443);
xor UO_1782 (O_1782,N_29509,N_28928);
and UO_1783 (O_1783,N_28922,N_29797);
nand UO_1784 (O_1784,N_28883,N_29690);
nand UO_1785 (O_1785,N_28830,N_29578);
xnor UO_1786 (O_1786,N_29294,N_29042);
and UO_1787 (O_1787,N_28967,N_29565);
or UO_1788 (O_1788,N_29401,N_29278);
nand UO_1789 (O_1789,N_29349,N_29197);
nand UO_1790 (O_1790,N_29714,N_29773);
or UO_1791 (O_1791,N_28904,N_29020);
and UO_1792 (O_1792,N_29297,N_28800);
xor UO_1793 (O_1793,N_29883,N_29163);
or UO_1794 (O_1794,N_28831,N_29960);
or UO_1795 (O_1795,N_29347,N_28925);
nor UO_1796 (O_1796,N_29796,N_29544);
nor UO_1797 (O_1797,N_29262,N_29218);
xnor UO_1798 (O_1798,N_29188,N_29382);
and UO_1799 (O_1799,N_28908,N_29072);
nand UO_1800 (O_1800,N_29960,N_29822);
nor UO_1801 (O_1801,N_29796,N_29409);
or UO_1802 (O_1802,N_29684,N_29227);
nand UO_1803 (O_1803,N_29534,N_29788);
or UO_1804 (O_1804,N_29045,N_29775);
nor UO_1805 (O_1805,N_28800,N_29750);
and UO_1806 (O_1806,N_29279,N_29239);
nand UO_1807 (O_1807,N_29850,N_29801);
xnor UO_1808 (O_1808,N_29706,N_29223);
nor UO_1809 (O_1809,N_29377,N_29984);
or UO_1810 (O_1810,N_28847,N_29407);
or UO_1811 (O_1811,N_29229,N_28991);
and UO_1812 (O_1812,N_28879,N_29561);
nor UO_1813 (O_1813,N_29606,N_29222);
xnor UO_1814 (O_1814,N_29870,N_29157);
or UO_1815 (O_1815,N_29264,N_29883);
and UO_1816 (O_1816,N_29848,N_29028);
or UO_1817 (O_1817,N_29327,N_29759);
nand UO_1818 (O_1818,N_29886,N_28917);
or UO_1819 (O_1819,N_29173,N_29019);
and UO_1820 (O_1820,N_29605,N_29807);
and UO_1821 (O_1821,N_29289,N_29829);
nor UO_1822 (O_1822,N_29752,N_29790);
nand UO_1823 (O_1823,N_29076,N_28814);
and UO_1824 (O_1824,N_29753,N_29203);
xor UO_1825 (O_1825,N_29756,N_29618);
and UO_1826 (O_1826,N_29894,N_29364);
and UO_1827 (O_1827,N_29888,N_29556);
or UO_1828 (O_1828,N_29866,N_29712);
xor UO_1829 (O_1829,N_28806,N_29914);
and UO_1830 (O_1830,N_28938,N_29999);
nand UO_1831 (O_1831,N_29580,N_29177);
nor UO_1832 (O_1832,N_29730,N_29865);
nand UO_1833 (O_1833,N_29748,N_29596);
or UO_1834 (O_1834,N_29196,N_29134);
nor UO_1835 (O_1835,N_29393,N_29851);
nand UO_1836 (O_1836,N_28828,N_29944);
nand UO_1837 (O_1837,N_28935,N_29932);
and UO_1838 (O_1838,N_29576,N_28965);
and UO_1839 (O_1839,N_29994,N_28903);
xor UO_1840 (O_1840,N_29387,N_29441);
nand UO_1841 (O_1841,N_28996,N_29979);
and UO_1842 (O_1842,N_29405,N_29866);
xnor UO_1843 (O_1843,N_29211,N_29889);
or UO_1844 (O_1844,N_29511,N_29572);
xor UO_1845 (O_1845,N_29369,N_28961);
and UO_1846 (O_1846,N_29849,N_29002);
or UO_1847 (O_1847,N_29022,N_29832);
nor UO_1848 (O_1848,N_28834,N_28806);
xnor UO_1849 (O_1849,N_28806,N_28862);
or UO_1850 (O_1850,N_29261,N_29641);
xor UO_1851 (O_1851,N_29680,N_29458);
nand UO_1852 (O_1852,N_29279,N_29786);
or UO_1853 (O_1853,N_29074,N_29606);
nand UO_1854 (O_1854,N_29316,N_29085);
nand UO_1855 (O_1855,N_29601,N_29589);
or UO_1856 (O_1856,N_29844,N_29672);
nand UO_1857 (O_1857,N_29749,N_29699);
nor UO_1858 (O_1858,N_29805,N_29442);
and UO_1859 (O_1859,N_29947,N_29889);
nor UO_1860 (O_1860,N_29971,N_29025);
xnor UO_1861 (O_1861,N_29744,N_29798);
nor UO_1862 (O_1862,N_29555,N_29483);
nor UO_1863 (O_1863,N_29166,N_29325);
and UO_1864 (O_1864,N_29828,N_29420);
or UO_1865 (O_1865,N_29802,N_29941);
nand UO_1866 (O_1866,N_29720,N_29147);
or UO_1867 (O_1867,N_29893,N_28874);
or UO_1868 (O_1868,N_29438,N_29614);
and UO_1869 (O_1869,N_29279,N_28902);
or UO_1870 (O_1870,N_29311,N_28856);
nor UO_1871 (O_1871,N_29521,N_29184);
nand UO_1872 (O_1872,N_29024,N_29668);
nor UO_1873 (O_1873,N_29530,N_29698);
nor UO_1874 (O_1874,N_29183,N_29367);
xor UO_1875 (O_1875,N_29783,N_29077);
xnor UO_1876 (O_1876,N_29298,N_29813);
or UO_1877 (O_1877,N_29369,N_29124);
or UO_1878 (O_1878,N_29312,N_29170);
nor UO_1879 (O_1879,N_29844,N_28902);
nor UO_1880 (O_1880,N_29754,N_29147);
and UO_1881 (O_1881,N_29723,N_29610);
and UO_1882 (O_1882,N_28844,N_29469);
nand UO_1883 (O_1883,N_29452,N_29119);
or UO_1884 (O_1884,N_29105,N_29407);
and UO_1885 (O_1885,N_29204,N_28907);
xor UO_1886 (O_1886,N_28947,N_29560);
or UO_1887 (O_1887,N_29939,N_29440);
or UO_1888 (O_1888,N_28824,N_29522);
or UO_1889 (O_1889,N_29709,N_29782);
nand UO_1890 (O_1890,N_28803,N_28903);
xor UO_1891 (O_1891,N_29644,N_28839);
nand UO_1892 (O_1892,N_29528,N_29702);
nor UO_1893 (O_1893,N_29452,N_29825);
nor UO_1894 (O_1894,N_29502,N_28999);
or UO_1895 (O_1895,N_28974,N_29106);
nand UO_1896 (O_1896,N_29396,N_29764);
nor UO_1897 (O_1897,N_29487,N_29604);
or UO_1898 (O_1898,N_29373,N_29609);
nand UO_1899 (O_1899,N_29628,N_29097);
xor UO_1900 (O_1900,N_29158,N_29346);
and UO_1901 (O_1901,N_29803,N_29720);
nor UO_1902 (O_1902,N_29987,N_28849);
or UO_1903 (O_1903,N_29600,N_28803);
xnor UO_1904 (O_1904,N_29692,N_29269);
nand UO_1905 (O_1905,N_29200,N_29078);
nand UO_1906 (O_1906,N_29810,N_29179);
nor UO_1907 (O_1907,N_28882,N_28851);
nand UO_1908 (O_1908,N_29930,N_29135);
nand UO_1909 (O_1909,N_29171,N_29487);
nor UO_1910 (O_1910,N_29319,N_28916);
nor UO_1911 (O_1911,N_29699,N_29851);
xnor UO_1912 (O_1912,N_29739,N_28925);
or UO_1913 (O_1913,N_29769,N_28890);
or UO_1914 (O_1914,N_29365,N_29335);
xnor UO_1915 (O_1915,N_28930,N_28808);
nor UO_1916 (O_1916,N_29789,N_28823);
nor UO_1917 (O_1917,N_29742,N_28832);
nor UO_1918 (O_1918,N_29714,N_29537);
nand UO_1919 (O_1919,N_29420,N_29101);
and UO_1920 (O_1920,N_29033,N_29360);
nand UO_1921 (O_1921,N_29088,N_29946);
and UO_1922 (O_1922,N_29270,N_29820);
and UO_1923 (O_1923,N_29314,N_29204);
nor UO_1924 (O_1924,N_28965,N_29414);
xnor UO_1925 (O_1925,N_29041,N_29249);
nor UO_1926 (O_1926,N_29605,N_29774);
and UO_1927 (O_1927,N_28947,N_29959);
or UO_1928 (O_1928,N_29130,N_29126);
and UO_1929 (O_1929,N_29474,N_29762);
nor UO_1930 (O_1930,N_29959,N_29597);
xnor UO_1931 (O_1931,N_29391,N_29767);
and UO_1932 (O_1932,N_29292,N_29373);
and UO_1933 (O_1933,N_29229,N_29726);
nand UO_1934 (O_1934,N_29651,N_29058);
or UO_1935 (O_1935,N_29229,N_29827);
nand UO_1936 (O_1936,N_29179,N_29097);
and UO_1937 (O_1937,N_29089,N_29290);
or UO_1938 (O_1938,N_29767,N_29454);
nor UO_1939 (O_1939,N_29467,N_29622);
nor UO_1940 (O_1940,N_29462,N_29468);
xnor UO_1941 (O_1941,N_29939,N_29530);
nand UO_1942 (O_1942,N_29345,N_29521);
or UO_1943 (O_1943,N_28935,N_29191);
and UO_1944 (O_1944,N_29533,N_29515);
nor UO_1945 (O_1945,N_29751,N_29736);
nand UO_1946 (O_1946,N_28801,N_29707);
nand UO_1947 (O_1947,N_29192,N_29127);
nor UO_1948 (O_1948,N_28926,N_29328);
nor UO_1949 (O_1949,N_29789,N_28843);
and UO_1950 (O_1950,N_29055,N_29305);
nor UO_1951 (O_1951,N_29946,N_29585);
and UO_1952 (O_1952,N_29094,N_29182);
or UO_1953 (O_1953,N_29107,N_29590);
nor UO_1954 (O_1954,N_29304,N_29825);
nand UO_1955 (O_1955,N_29589,N_29783);
or UO_1956 (O_1956,N_29622,N_29911);
and UO_1957 (O_1957,N_29780,N_29784);
and UO_1958 (O_1958,N_29853,N_29724);
nand UO_1959 (O_1959,N_29159,N_28910);
nor UO_1960 (O_1960,N_29784,N_29022);
nor UO_1961 (O_1961,N_29634,N_29925);
and UO_1962 (O_1962,N_29506,N_28897);
xor UO_1963 (O_1963,N_29321,N_28898);
xor UO_1964 (O_1964,N_29248,N_29693);
and UO_1965 (O_1965,N_29483,N_29608);
nand UO_1966 (O_1966,N_29692,N_29700);
xor UO_1967 (O_1967,N_28894,N_28938);
nor UO_1968 (O_1968,N_29548,N_29915);
xor UO_1969 (O_1969,N_29477,N_29854);
and UO_1970 (O_1970,N_29078,N_28817);
xor UO_1971 (O_1971,N_29063,N_29593);
xor UO_1972 (O_1972,N_29721,N_29259);
nand UO_1973 (O_1973,N_29825,N_29055);
nand UO_1974 (O_1974,N_29685,N_29436);
nor UO_1975 (O_1975,N_29994,N_29218);
nor UO_1976 (O_1976,N_29231,N_29341);
nor UO_1977 (O_1977,N_29060,N_28990);
nor UO_1978 (O_1978,N_29529,N_29649);
and UO_1979 (O_1979,N_29455,N_29151);
nor UO_1980 (O_1980,N_29304,N_28805);
xor UO_1981 (O_1981,N_29224,N_29698);
nor UO_1982 (O_1982,N_29333,N_29777);
xor UO_1983 (O_1983,N_29397,N_29266);
nand UO_1984 (O_1984,N_29177,N_28827);
or UO_1985 (O_1985,N_29341,N_29233);
or UO_1986 (O_1986,N_29902,N_29477);
xor UO_1987 (O_1987,N_29853,N_29682);
and UO_1988 (O_1988,N_29918,N_29694);
xnor UO_1989 (O_1989,N_28913,N_29335);
or UO_1990 (O_1990,N_28903,N_28994);
nor UO_1991 (O_1991,N_29223,N_29976);
nor UO_1992 (O_1992,N_29386,N_29722);
nor UO_1993 (O_1993,N_29534,N_28808);
or UO_1994 (O_1994,N_28879,N_28871);
nand UO_1995 (O_1995,N_29845,N_29856);
nor UO_1996 (O_1996,N_29007,N_28942);
nor UO_1997 (O_1997,N_29435,N_29174);
and UO_1998 (O_1998,N_29673,N_28826);
or UO_1999 (O_1999,N_29049,N_29777);
xnor UO_2000 (O_2000,N_29231,N_29568);
or UO_2001 (O_2001,N_29666,N_29256);
nor UO_2002 (O_2002,N_29456,N_29788);
and UO_2003 (O_2003,N_29700,N_29972);
nand UO_2004 (O_2004,N_29107,N_29958);
nand UO_2005 (O_2005,N_29534,N_28984);
nor UO_2006 (O_2006,N_29969,N_29124);
or UO_2007 (O_2007,N_29705,N_29430);
xor UO_2008 (O_2008,N_29916,N_28825);
and UO_2009 (O_2009,N_29936,N_29130);
or UO_2010 (O_2010,N_29835,N_28895);
nor UO_2011 (O_2011,N_29876,N_29079);
and UO_2012 (O_2012,N_29986,N_28895);
nor UO_2013 (O_2013,N_29218,N_29965);
and UO_2014 (O_2014,N_29023,N_29861);
or UO_2015 (O_2015,N_28927,N_28840);
xor UO_2016 (O_2016,N_28995,N_29182);
xor UO_2017 (O_2017,N_29662,N_29637);
or UO_2018 (O_2018,N_28870,N_29446);
nand UO_2019 (O_2019,N_29175,N_29391);
nand UO_2020 (O_2020,N_29808,N_29437);
nand UO_2021 (O_2021,N_29902,N_28969);
and UO_2022 (O_2022,N_29390,N_29258);
xnor UO_2023 (O_2023,N_28905,N_29186);
nor UO_2024 (O_2024,N_29389,N_29956);
xnor UO_2025 (O_2025,N_29790,N_29370);
and UO_2026 (O_2026,N_29149,N_28929);
and UO_2027 (O_2027,N_29175,N_28881);
or UO_2028 (O_2028,N_29217,N_29843);
or UO_2029 (O_2029,N_29911,N_28826);
nand UO_2030 (O_2030,N_29703,N_29656);
nor UO_2031 (O_2031,N_29655,N_28854);
xor UO_2032 (O_2032,N_29217,N_29126);
and UO_2033 (O_2033,N_29522,N_29008);
xnor UO_2034 (O_2034,N_29890,N_29110);
or UO_2035 (O_2035,N_28936,N_29944);
xnor UO_2036 (O_2036,N_29552,N_29174);
or UO_2037 (O_2037,N_29159,N_29885);
and UO_2038 (O_2038,N_29768,N_29624);
or UO_2039 (O_2039,N_29140,N_29314);
nand UO_2040 (O_2040,N_29512,N_29272);
and UO_2041 (O_2041,N_29760,N_29667);
nand UO_2042 (O_2042,N_29417,N_28916);
nor UO_2043 (O_2043,N_29920,N_29665);
and UO_2044 (O_2044,N_29798,N_29071);
nor UO_2045 (O_2045,N_28939,N_29568);
or UO_2046 (O_2046,N_29579,N_29531);
nor UO_2047 (O_2047,N_29526,N_29582);
xor UO_2048 (O_2048,N_29465,N_29019);
or UO_2049 (O_2049,N_28941,N_29340);
xor UO_2050 (O_2050,N_29690,N_29481);
xor UO_2051 (O_2051,N_28912,N_29351);
nand UO_2052 (O_2052,N_29869,N_29391);
or UO_2053 (O_2053,N_29419,N_29038);
and UO_2054 (O_2054,N_29140,N_29053);
nand UO_2055 (O_2055,N_29160,N_29763);
xnor UO_2056 (O_2056,N_29457,N_29095);
nor UO_2057 (O_2057,N_28814,N_29271);
or UO_2058 (O_2058,N_29676,N_29687);
nand UO_2059 (O_2059,N_29751,N_29931);
and UO_2060 (O_2060,N_29232,N_29686);
nor UO_2061 (O_2061,N_29406,N_29696);
nand UO_2062 (O_2062,N_29839,N_29376);
nand UO_2063 (O_2063,N_29579,N_29176);
and UO_2064 (O_2064,N_28991,N_29253);
or UO_2065 (O_2065,N_29818,N_29131);
or UO_2066 (O_2066,N_29164,N_29202);
nand UO_2067 (O_2067,N_28826,N_29890);
nor UO_2068 (O_2068,N_29971,N_28984);
and UO_2069 (O_2069,N_29402,N_29445);
nor UO_2070 (O_2070,N_28957,N_29265);
and UO_2071 (O_2071,N_29502,N_29777);
and UO_2072 (O_2072,N_29400,N_29448);
xnor UO_2073 (O_2073,N_29893,N_29342);
and UO_2074 (O_2074,N_28834,N_29271);
nand UO_2075 (O_2075,N_28804,N_29662);
nor UO_2076 (O_2076,N_29926,N_28899);
xnor UO_2077 (O_2077,N_29523,N_29675);
and UO_2078 (O_2078,N_29396,N_29437);
and UO_2079 (O_2079,N_29498,N_29869);
or UO_2080 (O_2080,N_29981,N_29048);
and UO_2081 (O_2081,N_29127,N_29848);
or UO_2082 (O_2082,N_29730,N_29389);
and UO_2083 (O_2083,N_29628,N_29520);
and UO_2084 (O_2084,N_29191,N_28930);
or UO_2085 (O_2085,N_29345,N_29984);
and UO_2086 (O_2086,N_29332,N_29709);
nand UO_2087 (O_2087,N_29453,N_29379);
and UO_2088 (O_2088,N_28983,N_29803);
xor UO_2089 (O_2089,N_28854,N_28841);
or UO_2090 (O_2090,N_28995,N_29576);
and UO_2091 (O_2091,N_29179,N_29542);
nor UO_2092 (O_2092,N_29869,N_29168);
nor UO_2093 (O_2093,N_29181,N_29212);
nand UO_2094 (O_2094,N_29628,N_29561);
or UO_2095 (O_2095,N_28940,N_28936);
and UO_2096 (O_2096,N_29292,N_29291);
xnor UO_2097 (O_2097,N_28804,N_29142);
xnor UO_2098 (O_2098,N_29278,N_29532);
xor UO_2099 (O_2099,N_29333,N_29367);
nand UO_2100 (O_2100,N_29161,N_29319);
xnor UO_2101 (O_2101,N_29158,N_28853);
nand UO_2102 (O_2102,N_29273,N_29499);
nand UO_2103 (O_2103,N_29894,N_29206);
or UO_2104 (O_2104,N_29457,N_29369);
xor UO_2105 (O_2105,N_29220,N_29013);
nor UO_2106 (O_2106,N_29491,N_29070);
or UO_2107 (O_2107,N_28857,N_29559);
or UO_2108 (O_2108,N_29729,N_29394);
nor UO_2109 (O_2109,N_29863,N_29361);
nor UO_2110 (O_2110,N_29835,N_29801);
nand UO_2111 (O_2111,N_29534,N_29413);
and UO_2112 (O_2112,N_29357,N_28865);
and UO_2113 (O_2113,N_29399,N_29334);
and UO_2114 (O_2114,N_28991,N_29720);
nor UO_2115 (O_2115,N_29648,N_29116);
nor UO_2116 (O_2116,N_29744,N_29072);
xor UO_2117 (O_2117,N_29550,N_29235);
or UO_2118 (O_2118,N_29951,N_29089);
nand UO_2119 (O_2119,N_29549,N_29859);
nor UO_2120 (O_2120,N_29768,N_28857);
and UO_2121 (O_2121,N_29078,N_29484);
and UO_2122 (O_2122,N_29348,N_28935);
nor UO_2123 (O_2123,N_29920,N_28862);
nand UO_2124 (O_2124,N_29988,N_29711);
or UO_2125 (O_2125,N_29649,N_29058);
nand UO_2126 (O_2126,N_29736,N_29356);
xnor UO_2127 (O_2127,N_29127,N_29949);
nand UO_2128 (O_2128,N_29566,N_29110);
xnor UO_2129 (O_2129,N_29501,N_29261);
and UO_2130 (O_2130,N_29983,N_29717);
or UO_2131 (O_2131,N_29390,N_29909);
xor UO_2132 (O_2132,N_29218,N_29278);
nor UO_2133 (O_2133,N_29368,N_29792);
nand UO_2134 (O_2134,N_28992,N_28939);
and UO_2135 (O_2135,N_28839,N_28956);
xor UO_2136 (O_2136,N_29678,N_29661);
nor UO_2137 (O_2137,N_29565,N_29527);
nor UO_2138 (O_2138,N_28934,N_29810);
nor UO_2139 (O_2139,N_29287,N_29303);
or UO_2140 (O_2140,N_29508,N_29805);
nor UO_2141 (O_2141,N_29229,N_29358);
nor UO_2142 (O_2142,N_29205,N_29578);
xnor UO_2143 (O_2143,N_29545,N_29947);
or UO_2144 (O_2144,N_29699,N_29170);
xor UO_2145 (O_2145,N_29542,N_28910);
xor UO_2146 (O_2146,N_29790,N_28982);
xor UO_2147 (O_2147,N_29176,N_29476);
xnor UO_2148 (O_2148,N_29491,N_29734);
nand UO_2149 (O_2149,N_29209,N_29784);
nand UO_2150 (O_2150,N_29070,N_29398);
nor UO_2151 (O_2151,N_29050,N_29461);
xnor UO_2152 (O_2152,N_29907,N_29448);
xnor UO_2153 (O_2153,N_29991,N_29130);
nand UO_2154 (O_2154,N_29272,N_29078);
xnor UO_2155 (O_2155,N_29726,N_29452);
and UO_2156 (O_2156,N_29246,N_29412);
and UO_2157 (O_2157,N_29396,N_29746);
nand UO_2158 (O_2158,N_29599,N_28844);
xnor UO_2159 (O_2159,N_29545,N_29570);
xnor UO_2160 (O_2160,N_28976,N_29908);
nor UO_2161 (O_2161,N_29773,N_29281);
nor UO_2162 (O_2162,N_29564,N_29656);
nand UO_2163 (O_2163,N_28973,N_28870);
and UO_2164 (O_2164,N_29360,N_29724);
and UO_2165 (O_2165,N_29512,N_29463);
nor UO_2166 (O_2166,N_29481,N_29014);
xor UO_2167 (O_2167,N_28818,N_28978);
nor UO_2168 (O_2168,N_29324,N_28880);
nand UO_2169 (O_2169,N_29885,N_28822);
and UO_2170 (O_2170,N_28835,N_29968);
nor UO_2171 (O_2171,N_29171,N_29886);
or UO_2172 (O_2172,N_29566,N_29301);
xnor UO_2173 (O_2173,N_29814,N_29119);
nand UO_2174 (O_2174,N_29189,N_29880);
or UO_2175 (O_2175,N_29259,N_29419);
nor UO_2176 (O_2176,N_29983,N_29178);
xnor UO_2177 (O_2177,N_29004,N_29615);
xor UO_2178 (O_2178,N_29684,N_29168);
nand UO_2179 (O_2179,N_28910,N_29669);
xnor UO_2180 (O_2180,N_29807,N_29235);
and UO_2181 (O_2181,N_29772,N_29472);
or UO_2182 (O_2182,N_29791,N_28823);
xnor UO_2183 (O_2183,N_28953,N_29299);
and UO_2184 (O_2184,N_29383,N_29614);
nor UO_2185 (O_2185,N_29722,N_29478);
and UO_2186 (O_2186,N_29422,N_28860);
nor UO_2187 (O_2187,N_29502,N_29271);
and UO_2188 (O_2188,N_29665,N_29485);
nor UO_2189 (O_2189,N_28860,N_28892);
or UO_2190 (O_2190,N_29453,N_29964);
or UO_2191 (O_2191,N_29855,N_29580);
or UO_2192 (O_2192,N_29351,N_29570);
and UO_2193 (O_2193,N_28927,N_29750);
and UO_2194 (O_2194,N_28839,N_29494);
or UO_2195 (O_2195,N_29806,N_29719);
nor UO_2196 (O_2196,N_29426,N_29836);
or UO_2197 (O_2197,N_29777,N_29354);
xnor UO_2198 (O_2198,N_29405,N_29909);
nand UO_2199 (O_2199,N_29237,N_29993);
nor UO_2200 (O_2200,N_28831,N_29832);
and UO_2201 (O_2201,N_29326,N_29818);
or UO_2202 (O_2202,N_29608,N_29980);
or UO_2203 (O_2203,N_29661,N_29206);
nor UO_2204 (O_2204,N_29225,N_29461);
and UO_2205 (O_2205,N_29888,N_29649);
nand UO_2206 (O_2206,N_28957,N_29719);
xnor UO_2207 (O_2207,N_29501,N_29679);
and UO_2208 (O_2208,N_29657,N_29753);
nor UO_2209 (O_2209,N_29915,N_29169);
or UO_2210 (O_2210,N_29053,N_29893);
and UO_2211 (O_2211,N_29006,N_29982);
nor UO_2212 (O_2212,N_29708,N_29078);
nor UO_2213 (O_2213,N_29941,N_29553);
nor UO_2214 (O_2214,N_28949,N_29585);
or UO_2215 (O_2215,N_29465,N_29989);
or UO_2216 (O_2216,N_29200,N_29389);
xor UO_2217 (O_2217,N_28942,N_29288);
nor UO_2218 (O_2218,N_28969,N_29845);
nand UO_2219 (O_2219,N_29308,N_29593);
nand UO_2220 (O_2220,N_28824,N_29155);
nor UO_2221 (O_2221,N_29161,N_29414);
nand UO_2222 (O_2222,N_28874,N_29422);
nor UO_2223 (O_2223,N_29284,N_29877);
and UO_2224 (O_2224,N_29012,N_29216);
and UO_2225 (O_2225,N_29763,N_28825);
nand UO_2226 (O_2226,N_29211,N_29128);
xnor UO_2227 (O_2227,N_29471,N_29560);
or UO_2228 (O_2228,N_29455,N_29592);
nor UO_2229 (O_2229,N_29042,N_29062);
nand UO_2230 (O_2230,N_29449,N_29530);
nand UO_2231 (O_2231,N_29727,N_29582);
and UO_2232 (O_2232,N_28999,N_29762);
or UO_2233 (O_2233,N_29659,N_29678);
or UO_2234 (O_2234,N_29452,N_29026);
nor UO_2235 (O_2235,N_29961,N_29939);
or UO_2236 (O_2236,N_29480,N_28925);
and UO_2237 (O_2237,N_29547,N_29204);
nor UO_2238 (O_2238,N_28897,N_29010);
nor UO_2239 (O_2239,N_29841,N_28806);
xor UO_2240 (O_2240,N_29517,N_29582);
and UO_2241 (O_2241,N_29426,N_29444);
or UO_2242 (O_2242,N_29021,N_29053);
nor UO_2243 (O_2243,N_29130,N_29402);
nor UO_2244 (O_2244,N_29097,N_28971);
nor UO_2245 (O_2245,N_29507,N_29481);
or UO_2246 (O_2246,N_29428,N_29101);
or UO_2247 (O_2247,N_29921,N_29944);
xor UO_2248 (O_2248,N_29354,N_29279);
and UO_2249 (O_2249,N_29397,N_28984);
nand UO_2250 (O_2250,N_29750,N_28819);
nor UO_2251 (O_2251,N_29856,N_28878);
nor UO_2252 (O_2252,N_29187,N_29917);
xnor UO_2253 (O_2253,N_29003,N_29241);
nand UO_2254 (O_2254,N_29894,N_29967);
and UO_2255 (O_2255,N_28877,N_29857);
nor UO_2256 (O_2256,N_29362,N_29395);
xor UO_2257 (O_2257,N_29047,N_29278);
nor UO_2258 (O_2258,N_29222,N_29028);
xor UO_2259 (O_2259,N_29731,N_29781);
and UO_2260 (O_2260,N_29408,N_29994);
xnor UO_2261 (O_2261,N_29672,N_29493);
xor UO_2262 (O_2262,N_29372,N_29412);
and UO_2263 (O_2263,N_29103,N_29231);
and UO_2264 (O_2264,N_29976,N_28964);
or UO_2265 (O_2265,N_29730,N_29641);
xnor UO_2266 (O_2266,N_28984,N_29522);
and UO_2267 (O_2267,N_29476,N_29516);
and UO_2268 (O_2268,N_29279,N_29480);
nand UO_2269 (O_2269,N_29662,N_28819);
xnor UO_2270 (O_2270,N_28861,N_29621);
xor UO_2271 (O_2271,N_29621,N_29790);
and UO_2272 (O_2272,N_28886,N_29107);
xor UO_2273 (O_2273,N_29001,N_29807);
and UO_2274 (O_2274,N_28933,N_28903);
and UO_2275 (O_2275,N_29116,N_29458);
and UO_2276 (O_2276,N_29561,N_29594);
or UO_2277 (O_2277,N_28955,N_29358);
xor UO_2278 (O_2278,N_29422,N_29815);
and UO_2279 (O_2279,N_29936,N_29744);
nor UO_2280 (O_2280,N_29702,N_29424);
or UO_2281 (O_2281,N_29623,N_29712);
or UO_2282 (O_2282,N_28950,N_28987);
nor UO_2283 (O_2283,N_29905,N_29364);
nor UO_2284 (O_2284,N_29131,N_29055);
and UO_2285 (O_2285,N_29107,N_29843);
nor UO_2286 (O_2286,N_29272,N_29460);
xor UO_2287 (O_2287,N_29244,N_28812);
and UO_2288 (O_2288,N_29652,N_29613);
and UO_2289 (O_2289,N_29544,N_28860);
and UO_2290 (O_2290,N_28842,N_29180);
or UO_2291 (O_2291,N_29584,N_29440);
or UO_2292 (O_2292,N_29987,N_29982);
nor UO_2293 (O_2293,N_29256,N_29715);
and UO_2294 (O_2294,N_29922,N_29295);
and UO_2295 (O_2295,N_29832,N_29863);
nor UO_2296 (O_2296,N_29602,N_29143);
xnor UO_2297 (O_2297,N_29438,N_28983);
nand UO_2298 (O_2298,N_29418,N_29925);
or UO_2299 (O_2299,N_29271,N_28935);
and UO_2300 (O_2300,N_29667,N_29596);
and UO_2301 (O_2301,N_29724,N_28971);
xor UO_2302 (O_2302,N_28966,N_29927);
xor UO_2303 (O_2303,N_29517,N_29340);
nor UO_2304 (O_2304,N_29454,N_29712);
or UO_2305 (O_2305,N_29987,N_29095);
nor UO_2306 (O_2306,N_29711,N_29692);
or UO_2307 (O_2307,N_29261,N_29256);
xnor UO_2308 (O_2308,N_29692,N_29494);
nor UO_2309 (O_2309,N_28910,N_28962);
nand UO_2310 (O_2310,N_29693,N_29469);
nand UO_2311 (O_2311,N_28870,N_29622);
nand UO_2312 (O_2312,N_28821,N_29706);
xnor UO_2313 (O_2313,N_29428,N_29073);
and UO_2314 (O_2314,N_29569,N_29114);
xor UO_2315 (O_2315,N_29119,N_28968);
nand UO_2316 (O_2316,N_29248,N_29267);
or UO_2317 (O_2317,N_28933,N_29799);
xor UO_2318 (O_2318,N_29946,N_29797);
or UO_2319 (O_2319,N_29082,N_29299);
xnor UO_2320 (O_2320,N_29088,N_29265);
nand UO_2321 (O_2321,N_29562,N_29797);
nand UO_2322 (O_2322,N_29780,N_29205);
nor UO_2323 (O_2323,N_29054,N_29908);
nor UO_2324 (O_2324,N_29563,N_29752);
nand UO_2325 (O_2325,N_29214,N_29496);
or UO_2326 (O_2326,N_29677,N_28813);
nor UO_2327 (O_2327,N_29476,N_29948);
nor UO_2328 (O_2328,N_29633,N_29891);
nand UO_2329 (O_2329,N_29779,N_29868);
nor UO_2330 (O_2330,N_29513,N_29889);
and UO_2331 (O_2331,N_28988,N_29617);
and UO_2332 (O_2332,N_29653,N_29994);
or UO_2333 (O_2333,N_29971,N_29070);
nand UO_2334 (O_2334,N_29021,N_29540);
nor UO_2335 (O_2335,N_29894,N_29919);
nor UO_2336 (O_2336,N_29707,N_29517);
nand UO_2337 (O_2337,N_29927,N_29055);
nor UO_2338 (O_2338,N_29121,N_29057);
nor UO_2339 (O_2339,N_28810,N_29781);
or UO_2340 (O_2340,N_29416,N_29660);
xor UO_2341 (O_2341,N_29849,N_28926);
and UO_2342 (O_2342,N_29849,N_28923);
or UO_2343 (O_2343,N_29308,N_29986);
and UO_2344 (O_2344,N_29118,N_29451);
xor UO_2345 (O_2345,N_29342,N_29843);
nor UO_2346 (O_2346,N_29041,N_29354);
nor UO_2347 (O_2347,N_29739,N_29922);
or UO_2348 (O_2348,N_29704,N_29098);
nand UO_2349 (O_2349,N_29649,N_29553);
nand UO_2350 (O_2350,N_29712,N_28930);
or UO_2351 (O_2351,N_29076,N_29485);
and UO_2352 (O_2352,N_29117,N_29005);
nand UO_2353 (O_2353,N_28916,N_28974);
and UO_2354 (O_2354,N_28836,N_29189);
xnor UO_2355 (O_2355,N_29124,N_29117);
nor UO_2356 (O_2356,N_29336,N_28829);
nand UO_2357 (O_2357,N_29605,N_29566);
nand UO_2358 (O_2358,N_28997,N_29475);
or UO_2359 (O_2359,N_29142,N_29189);
nor UO_2360 (O_2360,N_29193,N_28957);
nor UO_2361 (O_2361,N_29890,N_29719);
nor UO_2362 (O_2362,N_29547,N_29620);
and UO_2363 (O_2363,N_29651,N_29561);
and UO_2364 (O_2364,N_29464,N_28886);
nor UO_2365 (O_2365,N_29210,N_28963);
xnor UO_2366 (O_2366,N_29161,N_29967);
or UO_2367 (O_2367,N_29577,N_29669);
nand UO_2368 (O_2368,N_29339,N_29110);
nor UO_2369 (O_2369,N_29171,N_29271);
xnor UO_2370 (O_2370,N_29187,N_28904);
or UO_2371 (O_2371,N_29635,N_29027);
or UO_2372 (O_2372,N_29190,N_29657);
nand UO_2373 (O_2373,N_29767,N_29316);
nor UO_2374 (O_2374,N_28932,N_29185);
and UO_2375 (O_2375,N_29059,N_29446);
nor UO_2376 (O_2376,N_29740,N_29287);
nor UO_2377 (O_2377,N_29914,N_29773);
xor UO_2378 (O_2378,N_29592,N_29843);
nand UO_2379 (O_2379,N_29338,N_29454);
nand UO_2380 (O_2380,N_29331,N_29683);
nor UO_2381 (O_2381,N_28954,N_29370);
nor UO_2382 (O_2382,N_29423,N_29502);
nor UO_2383 (O_2383,N_29990,N_29685);
nor UO_2384 (O_2384,N_29141,N_29578);
and UO_2385 (O_2385,N_29141,N_29825);
nand UO_2386 (O_2386,N_29279,N_28976);
xor UO_2387 (O_2387,N_29658,N_29403);
nand UO_2388 (O_2388,N_29124,N_29870);
and UO_2389 (O_2389,N_29722,N_29952);
or UO_2390 (O_2390,N_29786,N_29734);
nor UO_2391 (O_2391,N_29401,N_29553);
nand UO_2392 (O_2392,N_29611,N_29640);
xor UO_2393 (O_2393,N_29095,N_29789);
or UO_2394 (O_2394,N_29057,N_29487);
nor UO_2395 (O_2395,N_28999,N_29507);
or UO_2396 (O_2396,N_29854,N_29546);
xnor UO_2397 (O_2397,N_29033,N_29265);
nand UO_2398 (O_2398,N_29110,N_29535);
xnor UO_2399 (O_2399,N_29916,N_29074);
xor UO_2400 (O_2400,N_28940,N_29384);
or UO_2401 (O_2401,N_29796,N_29025);
nor UO_2402 (O_2402,N_29947,N_29059);
nand UO_2403 (O_2403,N_29904,N_29924);
and UO_2404 (O_2404,N_29326,N_29730);
or UO_2405 (O_2405,N_29818,N_29037);
and UO_2406 (O_2406,N_29670,N_29963);
nor UO_2407 (O_2407,N_29840,N_29681);
nand UO_2408 (O_2408,N_29816,N_29771);
or UO_2409 (O_2409,N_29904,N_29990);
and UO_2410 (O_2410,N_28986,N_29042);
xor UO_2411 (O_2411,N_29827,N_29570);
and UO_2412 (O_2412,N_28880,N_28981);
or UO_2413 (O_2413,N_29134,N_29153);
and UO_2414 (O_2414,N_29699,N_29897);
and UO_2415 (O_2415,N_29948,N_29565);
and UO_2416 (O_2416,N_29744,N_29728);
or UO_2417 (O_2417,N_29518,N_29193);
xnor UO_2418 (O_2418,N_29474,N_29947);
nand UO_2419 (O_2419,N_29966,N_29897);
and UO_2420 (O_2420,N_29887,N_29503);
xor UO_2421 (O_2421,N_29968,N_29865);
xor UO_2422 (O_2422,N_29819,N_29667);
nor UO_2423 (O_2423,N_29881,N_29868);
xnor UO_2424 (O_2424,N_29500,N_29451);
and UO_2425 (O_2425,N_29666,N_29230);
xnor UO_2426 (O_2426,N_28810,N_28960);
nor UO_2427 (O_2427,N_28980,N_29604);
xor UO_2428 (O_2428,N_29241,N_29948);
and UO_2429 (O_2429,N_29170,N_29396);
xnor UO_2430 (O_2430,N_29772,N_29465);
or UO_2431 (O_2431,N_29819,N_29577);
nor UO_2432 (O_2432,N_29072,N_29688);
nand UO_2433 (O_2433,N_28834,N_29583);
and UO_2434 (O_2434,N_28932,N_29320);
nor UO_2435 (O_2435,N_29114,N_29402);
or UO_2436 (O_2436,N_28903,N_29298);
nor UO_2437 (O_2437,N_29672,N_29034);
nand UO_2438 (O_2438,N_28973,N_29872);
xor UO_2439 (O_2439,N_29486,N_29543);
nand UO_2440 (O_2440,N_29101,N_29163);
xor UO_2441 (O_2441,N_29451,N_29082);
nand UO_2442 (O_2442,N_29001,N_29914);
xnor UO_2443 (O_2443,N_29630,N_29669);
xor UO_2444 (O_2444,N_29547,N_29697);
or UO_2445 (O_2445,N_29578,N_29812);
nand UO_2446 (O_2446,N_29448,N_29731);
xnor UO_2447 (O_2447,N_28903,N_29146);
and UO_2448 (O_2448,N_29697,N_29031);
nor UO_2449 (O_2449,N_29072,N_28965);
xor UO_2450 (O_2450,N_29700,N_28985);
xor UO_2451 (O_2451,N_29348,N_28994);
nand UO_2452 (O_2452,N_29523,N_29980);
nand UO_2453 (O_2453,N_29506,N_29639);
xor UO_2454 (O_2454,N_29404,N_29929);
and UO_2455 (O_2455,N_29687,N_29249);
or UO_2456 (O_2456,N_29965,N_29947);
xnor UO_2457 (O_2457,N_29257,N_29057);
nor UO_2458 (O_2458,N_29568,N_29206);
or UO_2459 (O_2459,N_29090,N_29906);
nand UO_2460 (O_2460,N_29713,N_29007);
and UO_2461 (O_2461,N_29378,N_29949);
or UO_2462 (O_2462,N_29031,N_29910);
and UO_2463 (O_2463,N_29103,N_29653);
and UO_2464 (O_2464,N_29368,N_29873);
xor UO_2465 (O_2465,N_29633,N_28877);
nor UO_2466 (O_2466,N_29986,N_29437);
nor UO_2467 (O_2467,N_29221,N_29808);
and UO_2468 (O_2468,N_28978,N_29057);
or UO_2469 (O_2469,N_29417,N_29070);
or UO_2470 (O_2470,N_29028,N_29924);
nor UO_2471 (O_2471,N_29802,N_28809);
and UO_2472 (O_2472,N_28822,N_29343);
or UO_2473 (O_2473,N_29022,N_29468);
or UO_2474 (O_2474,N_29786,N_28877);
and UO_2475 (O_2475,N_29837,N_29648);
nor UO_2476 (O_2476,N_29120,N_28806);
and UO_2477 (O_2477,N_29440,N_29703);
nor UO_2478 (O_2478,N_29196,N_29237);
or UO_2479 (O_2479,N_28996,N_29705);
nor UO_2480 (O_2480,N_29632,N_29805);
or UO_2481 (O_2481,N_29206,N_29458);
and UO_2482 (O_2482,N_29048,N_29533);
nand UO_2483 (O_2483,N_29891,N_29408);
xnor UO_2484 (O_2484,N_29318,N_29243);
and UO_2485 (O_2485,N_29204,N_29445);
or UO_2486 (O_2486,N_29394,N_29539);
nand UO_2487 (O_2487,N_29346,N_29071);
and UO_2488 (O_2488,N_29740,N_29898);
and UO_2489 (O_2489,N_29645,N_29007);
or UO_2490 (O_2490,N_29280,N_29130);
nand UO_2491 (O_2491,N_28994,N_29607);
nor UO_2492 (O_2492,N_29265,N_28868);
or UO_2493 (O_2493,N_29435,N_29842);
and UO_2494 (O_2494,N_29204,N_29097);
and UO_2495 (O_2495,N_29913,N_28935);
nor UO_2496 (O_2496,N_29184,N_29869);
xor UO_2497 (O_2497,N_29275,N_29065);
and UO_2498 (O_2498,N_29518,N_29917);
and UO_2499 (O_2499,N_29146,N_29365);
nor UO_2500 (O_2500,N_29749,N_29114);
and UO_2501 (O_2501,N_29832,N_29134);
and UO_2502 (O_2502,N_29565,N_29836);
nor UO_2503 (O_2503,N_29001,N_29135);
nand UO_2504 (O_2504,N_29483,N_29389);
nor UO_2505 (O_2505,N_28861,N_29274);
and UO_2506 (O_2506,N_29727,N_28859);
nor UO_2507 (O_2507,N_29370,N_29815);
or UO_2508 (O_2508,N_29315,N_29656);
nor UO_2509 (O_2509,N_29198,N_29962);
nor UO_2510 (O_2510,N_29575,N_29788);
nand UO_2511 (O_2511,N_29624,N_29296);
nor UO_2512 (O_2512,N_28817,N_29776);
or UO_2513 (O_2513,N_29029,N_29808);
or UO_2514 (O_2514,N_29619,N_29790);
or UO_2515 (O_2515,N_29548,N_29698);
or UO_2516 (O_2516,N_29522,N_28803);
or UO_2517 (O_2517,N_28873,N_29992);
nor UO_2518 (O_2518,N_29915,N_29278);
nor UO_2519 (O_2519,N_29173,N_29435);
nor UO_2520 (O_2520,N_29701,N_29423);
or UO_2521 (O_2521,N_28881,N_29176);
and UO_2522 (O_2522,N_28933,N_29464);
nand UO_2523 (O_2523,N_29524,N_29613);
nor UO_2524 (O_2524,N_29956,N_29826);
xor UO_2525 (O_2525,N_29325,N_28806);
nand UO_2526 (O_2526,N_29241,N_29558);
xnor UO_2527 (O_2527,N_28969,N_28958);
xnor UO_2528 (O_2528,N_28858,N_29566);
and UO_2529 (O_2529,N_29175,N_29794);
nand UO_2530 (O_2530,N_28876,N_29425);
nand UO_2531 (O_2531,N_29741,N_29322);
nand UO_2532 (O_2532,N_29052,N_29216);
xnor UO_2533 (O_2533,N_29802,N_29697);
or UO_2534 (O_2534,N_29650,N_29326);
nand UO_2535 (O_2535,N_29780,N_29546);
or UO_2536 (O_2536,N_28931,N_29114);
xnor UO_2537 (O_2537,N_28809,N_29972);
xnor UO_2538 (O_2538,N_29029,N_29729);
nor UO_2539 (O_2539,N_29711,N_28971);
or UO_2540 (O_2540,N_29952,N_29284);
or UO_2541 (O_2541,N_29770,N_29952);
nor UO_2542 (O_2542,N_29147,N_29406);
nand UO_2543 (O_2543,N_29966,N_29769);
nand UO_2544 (O_2544,N_29491,N_29394);
xnor UO_2545 (O_2545,N_29049,N_29027);
or UO_2546 (O_2546,N_29253,N_29446);
or UO_2547 (O_2547,N_28977,N_29052);
nand UO_2548 (O_2548,N_29040,N_29960);
nand UO_2549 (O_2549,N_29788,N_29222);
and UO_2550 (O_2550,N_28936,N_29651);
nor UO_2551 (O_2551,N_29798,N_29356);
or UO_2552 (O_2552,N_29026,N_29681);
nor UO_2553 (O_2553,N_28974,N_28803);
or UO_2554 (O_2554,N_29637,N_28832);
nor UO_2555 (O_2555,N_29483,N_29698);
xor UO_2556 (O_2556,N_29147,N_29669);
xor UO_2557 (O_2557,N_29673,N_29211);
xnor UO_2558 (O_2558,N_29112,N_29702);
or UO_2559 (O_2559,N_29142,N_29725);
xnor UO_2560 (O_2560,N_28805,N_29884);
nor UO_2561 (O_2561,N_29124,N_29428);
nor UO_2562 (O_2562,N_29606,N_29549);
xor UO_2563 (O_2563,N_29309,N_29164);
xor UO_2564 (O_2564,N_29454,N_29655);
nand UO_2565 (O_2565,N_29714,N_29632);
and UO_2566 (O_2566,N_28857,N_28832);
nand UO_2567 (O_2567,N_29487,N_29166);
nand UO_2568 (O_2568,N_29400,N_29333);
xnor UO_2569 (O_2569,N_28826,N_29333);
and UO_2570 (O_2570,N_28873,N_29484);
or UO_2571 (O_2571,N_29202,N_29679);
and UO_2572 (O_2572,N_28917,N_29811);
xnor UO_2573 (O_2573,N_29706,N_29986);
nor UO_2574 (O_2574,N_29902,N_29561);
xnor UO_2575 (O_2575,N_29840,N_29108);
nor UO_2576 (O_2576,N_29077,N_29264);
or UO_2577 (O_2577,N_29872,N_29372);
nor UO_2578 (O_2578,N_29707,N_29243);
and UO_2579 (O_2579,N_29443,N_29160);
nor UO_2580 (O_2580,N_29584,N_28966);
xor UO_2581 (O_2581,N_29459,N_29570);
nand UO_2582 (O_2582,N_29376,N_29761);
or UO_2583 (O_2583,N_28852,N_28886);
nand UO_2584 (O_2584,N_29953,N_28810);
and UO_2585 (O_2585,N_28849,N_29409);
and UO_2586 (O_2586,N_29059,N_28933);
nand UO_2587 (O_2587,N_29201,N_29665);
or UO_2588 (O_2588,N_29193,N_28881);
nand UO_2589 (O_2589,N_29740,N_29934);
or UO_2590 (O_2590,N_29159,N_29582);
nand UO_2591 (O_2591,N_29519,N_29074);
nor UO_2592 (O_2592,N_29616,N_29897);
nand UO_2593 (O_2593,N_29556,N_29401);
or UO_2594 (O_2594,N_29825,N_29948);
nor UO_2595 (O_2595,N_29669,N_29862);
or UO_2596 (O_2596,N_29201,N_29197);
nand UO_2597 (O_2597,N_29618,N_28838);
nor UO_2598 (O_2598,N_28989,N_29258);
xnor UO_2599 (O_2599,N_29977,N_29676);
xor UO_2600 (O_2600,N_28955,N_28939);
xnor UO_2601 (O_2601,N_29206,N_29141);
xnor UO_2602 (O_2602,N_28810,N_29837);
nand UO_2603 (O_2603,N_28951,N_29310);
and UO_2604 (O_2604,N_29954,N_29566);
and UO_2605 (O_2605,N_29715,N_29628);
or UO_2606 (O_2606,N_29416,N_29670);
xor UO_2607 (O_2607,N_29991,N_29183);
nor UO_2608 (O_2608,N_29923,N_29961);
nand UO_2609 (O_2609,N_29396,N_29138);
nand UO_2610 (O_2610,N_29309,N_29258);
and UO_2611 (O_2611,N_29714,N_29492);
nand UO_2612 (O_2612,N_29576,N_28912);
and UO_2613 (O_2613,N_29277,N_29892);
and UO_2614 (O_2614,N_28945,N_28961);
xnor UO_2615 (O_2615,N_29374,N_29137);
and UO_2616 (O_2616,N_29779,N_29062);
and UO_2617 (O_2617,N_29682,N_29423);
xnor UO_2618 (O_2618,N_29522,N_29337);
and UO_2619 (O_2619,N_29069,N_29802);
and UO_2620 (O_2620,N_28814,N_29376);
nand UO_2621 (O_2621,N_28850,N_29859);
and UO_2622 (O_2622,N_29722,N_29939);
nand UO_2623 (O_2623,N_29194,N_29392);
and UO_2624 (O_2624,N_29673,N_29153);
nor UO_2625 (O_2625,N_29071,N_29429);
and UO_2626 (O_2626,N_29207,N_29346);
xnor UO_2627 (O_2627,N_29436,N_29472);
nand UO_2628 (O_2628,N_29543,N_29051);
nand UO_2629 (O_2629,N_29380,N_29624);
and UO_2630 (O_2630,N_29625,N_28920);
xnor UO_2631 (O_2631,N_29584,N_28833);
nor UO_2632 (O_2632,N_29926,N_29555);
nor UO_2633 (O_2633,N_28961,N_29320);
nor UO_2634 (O_2634,N_29765,N_28841);
nand UO_2635 (O_2635,N_29750,N_29569);
nand UO_2636 (O_2636,N_28874,N_29861);
nand UO_2637 (O_2637,N_29048,N_29828);
nand UO_2638 (O_2638,N_29648,N_29398);
and UO_2639 (O_2639,N_29620,N_29483);
xor UO_2640 (O_2640,N_29362,N_29835);
nand UO_2641 (O_2641,N_29433,N_29262);
nor UO_2642 (O_2642,N_29453,N_29431);
and UO_2643 (O_2643,N_29557,N_28835);
xnor UO_2644 (O_2644,N_28981,N_29487);
or UO_2645 (O_2645,N_29547,N_29230);
or UO_2646 (O_2646,N_29064,N_29880);
nor UO_2647 (O_2647,N_28852,N_29915);
or UO_2648 (O_2648,N_29281,N_29645);
nand UO_2649 (O_2649,N_28910,N_29787);
and UO_2650 (O_2650,N_29606,N_28826);
xor UO_2651 (O_2651,N_29015,N_28982);
xnor UO_2652 (O_2652,N_28989,N_29472);
or UO_2653 (O_2653,N_29935,N_29703);
nor UO_2654 (O_2654,N_29921,N_29842);
nor UO_2655 (O_2655,N_29385,N_29336);
and UO_2656 (O_2656,N_29594,N_28866);
nor UO_2657 (O_2657,N_29269,N_29828);
xor UO_2658 (O_2658,N_29418,N_29709);
nand UO_2659 (O_2659,N_29161,N_29411);
nor UO_2660 (O_2660,N_29455,N_28839);
nand UO_2661 (O_2661,N_28960,N_29844);
xor UO_2662 (O_2662,N_29130,N_29436);
or UO_2663 (O_2663,N_29757,N_29537);
or UO_2664 (O_2664,N_29511,N_29964);
nor UO_2665 (O_2665,N_29711,N_29466);
nand UO_2666 (O_2666,N_29163,N_29761);
nand UO_2667 (O_2667,N_29433,N_28879);
and UO_2668 (O_2668,N_29893,N_29170);
xnor UO_2669 (O_2669,N_29167,N_29686);
xor UO_2670 (O_2670,N_28937,N_29759);
xor UO_2671 (O_2671,N_28991,N_29727);
nor UO_2672 (O_2672,N_28871,N_29909);
nand UO_2673 (O_2673,N_29496,N_29436);
nor UO_2674 (O_2674,N_29993,N_28939);
or UO_2675 (O_2675,N_29504,N_29816);
nor UO_2676 (O_2676,N_29451,N_29719);
and UO_2677 (O_2677,N_29152,N_29651);
xor UO_2678 (O_2678,N_29902,N_29543);
and UO_2679 (O_2679,N_29935,N_28877);
or UO_2680 (O_2680,N_29557,N_29842);
xnor UO_2681 (O_2681,N_29190,N_28956);
or UO_2682 (O_2682,N_29973,N_29391);
or UO_2683 (O_2683,N_29988,N_29753);
and UO_2684 (O_2684,N_29188,N_28899);
xor UO_2685 (O_2685,N_29685,N_29089);
nand UO_2686 (O_2686,N_29972,N_29594);
xnor UO_2687 (O_2687,N_29368,N_29901);
nand UO_2688 (O_2688,N_29034,N_29047);
or UO_2689 (O_2689,N_29376,N_28870);
xor UO_2690 (O_2690,N_28987,N_29418);
and UO_2691 (O_2691,N_29377,N_28965);
xor UO_2692 (O_2692,N_29102,N_29893);
xnor UO_2693 (O_2693,N_29421,N_29012);
nand UO_2694 (O_2694,N_29183,N_29787);
and UO_2695 (O_2695,N_29242,N_29924);
or UO_2696 (O_2696,N_29809,N_29289);
and UO_2697 (O_2697,N_29148,N_28923);
xnor UO_2698 (O_2698,N_29998,N_29856);
and UO_2699 (O_2699,N_29660,N_29988);
or UO_2700 (O_2700,N_29963,N_29774);
xor UO_2701 (O_2701,N_29918,N_29877);
and UO_2702 (O_2702,N_28924,N_29192);
xor UO_2703 (O_2703,N_29979,N_28877);
and UO_2704 (O_2704,N_28818,N_28885);
nand UO_2705 (O_2705,N_29443,N_29977);
xor UO_2706 (O_2706,N_28801,N_28820);
and UO_2707 (O_2707,N_28924,N_29959);
nor UO_2708 (O_2708,N_28940,N_29050);
xnor UO_2709 (O_2709,N_29134,N_29809);
and UO_2710 (O_2710,N_29970,N_29403);
nand UO_2711 (O_2711,N_29658,N_29919);
and UO_2712 (O_2712,N_29208,N_29696);
or UO_2713 (O_2713,N_29103,N_29532);
nor UO_2714 (O_2714,N_29305,N_29423);
nand UO_2715 (O_2715,N_29150,N_29250);
and UO_2716 (O_2716,N_29389,N_29173);
xor UO_2717 (O_2717,N_29332,N_29913);
nand UO_2718 (O_2718,N_29477,N_29830);
nand UO_2719 (O_2719,N_29079,N_29796);
nor UO_2720 (O_2720,N_29536,N_29406);
nand UO_2721 (O_2721,N_29530,N_29725);
xnor UO_2722 (O_2722,N_29793,N_29753);
nand UO_2723 (O_2723,N_29416,N_29531);
and UO_2724 (O_2724,N_29000,N_29953);
xor UO_2725 (O_2725,N_29223,N_29449);
or UO_2726 (O_2726,N_29095,N_29088);
and UO_2727 (O_2727,N_29538,N_29348);
and UO_2728 (O_2728,N_29662,N_29270);
nand UO_2729 (O_2729,N_29284,N_29113);
and UO_2730 (O_2730,N_28967,N_29936);
nor UO_2731 (O_2731,N_29663,N_29810);
nor UO_2732 (O_2732,N_29994,N_29959);
or UO_2733 (O_2733,N_29689,N_29259);
nand UO_2734 (O_2734,N_29964,N_28899);
xnor UO_2735 (O_2735,N_29891,N_29230);
nor UO_2736 (O_2736,N_28820,N_29824);
nand UO_2737 (O_2737,N_29736,N_29690);
xnor UO_2738 (O_2738,N_28861,N_29030);
or UO_2739 (O_2739,N_29075,N_29702);
and UO_2740 (O_2740,N_29363,N_29472);
and UO_2741 (O_2741,N_28860,N_29438);
and UO_2742 (O_2742,N_29008,N_29001);
nor UO_2743 (O_2743,N_29633,N_28837);
xnor UO_2744 (O_2744,N_29947,N_29012);
and UO_2745 (O_2745,N_29276,N_28842);
nor UO_2746 (O_2746,N_29679,N_29819);
xnor UO_2747 (O_2747,N_29404,N_29011);
nor UO_2748 (O_2748,N_29261,N_28924);
nor UO_2749 (O_2749,N_29880,N_29870);
nand UO_2750 (O_2750,N_29660,N_29278);
nor UO_2751 (O_2751,N_29652,N_29663);
xor UO_2752 (O_2752,N_29099,N_29590);
nand UO_2753 (O_2753,N_29870,N_29773);
nor UO_2754 (O_2754,N_29540,N_29811);
nand UO_2755 (O_2755,N_28851,N_29276);
nor UO_2756 (O_2756,N_29000,N_29236);
nor UO_2757 (O_2757,N_29551,N_28958);
nor UO_2758 (O_2758,N_29225,N_29961);
nor UO_2759 (O_2759,N_28968,N_29553);
nor UO_2760 (O_2760,N_29190,N_29592);
or UO_2761 (O_2761,N_29036,N_29800);
nand UO_2762 (O_2762,N_29725,N_29675);
and UO_2763 (O_2763,N_29807,N_29741);
and UO_2764 (O_2764,N_29368,N_29278);
nand UO_2765 (O_2765,N_29147,N_29244);
nor UO_2766 (O_2766,N_29914,N_29970);
xnor UO_2767 (O_2767,N_29167,N_28844);
nor UO_2768 (O_2768,N_28818,N_28881);
xnor UO_2769 (O_2769,N_29612,N_29190);
xnor UO_2770 (O_2770,N_29930,N_29879);
xnor UO_2771 (O_2771,N_29568,N_29784);
nand UO_2772 (O_2772,N_29264,N_29526);
or UO_2773 (O_2773,N_29678,N_29184);
xnor UO_2774 (O_2774,N_29700,N_29767);
nand UO_2775 (O_2775,N_29133,N_29527);
nor UO_2776 (O_2776,N_28912,N_28904);
nand UO_2777 (O_2777,N_29292,N_29189);
nand UO_2778 (O_2778,N_29587,N_29681);
nor UO_2779 (O_2779,N_29901,N_29695);
nand UO_2780 (O_2780,N_29787,N_29028);
or UO_2781 (O_2781,N_29834,N_29727);
xnor UO_2782 (O_2782,N_29261,N_28845);
and UO_2783 (O_2783,N_29680,N_28954);
and UO_2784 (O_2784,N_29044,N_29702);
or UO_2785 (O_2785,N_29955,N_29359);
nor UO_2786 (O_2786,N_28852,N_29310);
xnor UO_2787 (O_2787,N_29509,N_29039);
nor UO_2788 (O_2788,N_29550,N_29011);
nor UO_2789 (O_2789,N_29921,N_29406);
and UO_2790 (O_2790,N_29449,N_29151);
or UO_2791 (O_2791,N_28841,N_29585);
nor UO_2792 (O_2792,N_29974,N_28999);
xor UO_2793 (O_2793,N_29345,N_29645);
and UO_2794 (O_2794,N_29281,N_29759);
or UO_2795 (O_2795,N_29403,N_29551);
and UO_2796 (O_2796,N_29141,N_29582);
or UO_2797 (O_2797,N_29689,N_29271);
nor UO_2798 (O_2798,N_28966,N_29873);
nand UO_2799 (O_2799,N_29421,N_29298);
nor UO_2800 (O_2800,N_29055,N_29423);
or UO_2801 (O_2801,N_29549,N_28943);
or UO_2802 (O_2802,N_29092,N_29047);
nand UO_2803 (O_2803,N_29627,N_29200);
nor UO_2804 (O_2804,N_29462,N_29874);
nand UO_2805 (O_2805,N_29406,N_28821);
xnor UO_2806 (O_2806,N_28806,N_29599);
or UO_2807 (O_2807,N_28888,N_29568);
xor UO_2808 (O_2808,N_29729,N_29014);
xor UO_2809 (O_2809,N_29748,N_28840);
and UO_2810 (O_2810,N_29423,N_29567);
or UO_2811 (O_2811,N_29031,N_29727);
nand UO_2812 (O_2812,N_29237,N_29359);
and UO_2813 (O_2813,N_29107,N_29459);
nor UO_2814 (O_2814,N_29162,N_28851);
nand UO_2815 (O_2815,N_29849,N_29992);
and UO_2816 (O_2816,N_29715,N_29156);
nand UO_2817 (O_2817,N_29925,N_29555);
or UO_2818 (O_2818,N_29508,N_28881);
nor UO_2819 (O_2819,N_29113,N_29728);
or UO_2820 (O_2820,N_29179,N_29394);
and UO_2821 (O_2821,N_29900,N_29096);
nand UO_2822 (O_2822,N_29583,N_29810);
and UO_2823 (O_2823,N_29471,N_29026);
nand UO_2824 (O_2824,N_28982,N_29320);
nand UO_2825 (O_2825,N_29243,N_29518);
xnor UO_2826 (O_2826,N_29312,N_29537);
or UO_2827 (O_2827,N_29904,N_28937);
nor UO_2828 (O_2828,N_29772,N_29676);
and UO_2829 (O_2829,N_29169,N_29676);
nand UO_2830 (O_2830,N_29348,N_28826);
and UO_2831 (O_2831,N_28883,N_29369);
and UO_2832 (O_2832,N_29832,N_29125);
nor UO_2833 (O_2833,N_29218,N_29848);
nand UO_2834 (O_2834,N_28911,N_29003);
or UO_2835 (O_2835,N_29415,N_29091);
xor UO_2836 (O_2836,N_29780,N_29811);
nand UO_2837 (O_2837,N_29625,N_29720);
nand UO_2838 (O_2838,N_29022,N_29551);
nor UO_2839 (O_2839,N_29497,N_29322);
nand UO_2840 (O_2840,N_29725,N_29172);
and UO_2841 (O_2841,N_28885,N_29729);
nand UO_2842 (O_2842,N_29941,N_29731);
or UO_2843 (O_2843,N_29827,N_29822);
nor UO_2844 (O_2844,N_29843,N_29605);
and UO_2845 (O_2845,N_28847,N_29814);
and UO_2846 (O_2846,N_29633,N_29710);
and UO_2847 (O_2847,N_28997,N_29410);
nand UO_2848 (O_2848,N_29368,N_29154);
and UO_2849 (O_2849,N_29407,N_29667);
and UO_2850 (O_2850,N_29573,N_29686);
and UO_2851 (O_2851,N_28894,N_29376);
and UO_2852 (O_2852,N_29444,N_28901);
nand UO_2853 (O_2853,N_29341,N_29140);
or UO_2854 (O_2854,N_29723,N_29753);
or UO_2855 (O_2855,N_29135,N_29348);
xor UO_2856 (O_2856,N_29015,N_29193);
and UO_2857 (O_2857,N_29962,N_29269);
xor UO_2858 (O_2858,N_29762,N_29362);
and UO_2859 (O_2859,N_29678,N_29348);
xor UO_2860 (O_2860,N_29287,N_29251);
nand UO_2861 (O_2861,N_29565,N_29274);
nor UO_2862 (O_2862,N_29076,N_29598);
nor UO_2863 (O_2863,N_29148,N_29625);
and UO_2864 (O_2864,N_28927,N_29910);
nor UO_2865 (O_2865,N_29460,N_28823);
nand UO_2866 (O_2866,N_29549,N_29174);
nand UO_2867 (O_2867,N_29867,N_29199);
xnor UO_2868 (O_2868,N_29089,N_28931);
and UO_2869 (O_2869,N_29818,N_29249);
or UO_2870 (O_2870,N_28812,N_29395);
nand UO_2871 (O_2871,N_29709,N_28892);
nor UO_2872 (O_2872,N_29739,N_29887);
and UO_2873 (O_2873,N_29227,N_29244);
nor UO_2874 (O_2874,N_29886,N_29638);
nand UO_2875 (O_2875,N_29626,N_29867);
nand UO_2876 (O_2876,N_29886,N_29313);
xnor UO_2877 (O_2877,N_29818,N_28932);
xnor UO_2878 (O_2878,N_29690,N_29403);
nand UO_2879 (O_2879,N_28949,N_29870);
nand UO_2880 (O_2880,N_28931,N_29675);
and UO_2881 (O_2881,N_29945,N_29242);
xnor UO_2882 (O_2882,N_28890,N_29668);
nand UO_2883 (O_2883,N_29760,N_28863);
nand UO_2884 (O_2884,N_29131,N_29435);
xor UO_2885 (O_2885,N_29922,N_29178);
xor UO_2886 (O_2886,N_29138,N_29910);
nor UO_2887 (O_2887,N_29637,N_29433);
xor UO_2888 (O_2888,N_29406,N_29949);
and UO_2889 (O_2889,N_28821,N_29218);
nor UO_2890 (O_2890,N_29516,N_29592);
nor UO_2891 (O_2891,N_29494,N_29472);
and UO_2892 (O_2892,N_29201,N_28931);
or UO_2893 (O_2893,N_29123,N_28824);
xor UO_2894 (O_2894,N_29914,N_29377);
nand UO_2895 (O_2895,N_29750,N_29104);
and UO_2896 (O_2896,N_29053,N_29911);
xor UO_2897 (O_2897,N_29196,N_29204);
nand UO_2898 (O_2898,N_29280,N_28906);
or UO_2899 (O_2899,N_29464,N_29503);
and UO_2900 (O_2900,N_29601,N_29659);
nor UO_2901 (O_2901,N_29912,N_28979);
xnor UO_2902 (O_2902,N_29962,N_29680);
nor UO_2903 (O_2903,N_28835,N_29994);
nor UO_2904 (O_2904,N_29288,N_29755);
nand UO_2905 (O_2905,N_29668,N_29212);
and UO_2906 (O_2906,N_29417,N_29349);
and UO_2907 (O_2907,N_29848,N_28840);
or UO_2908 (O_2908,N_29071,N_29086);
and UO_2909 (O_2909,N_29050,N_28823);
nand UO_2910 (O_2910,N_29124,N_29354);
and UO_2911 (O_2911,N_29143,N_29940);
nor UO_2912 (O_2912,N_29188,N_29943);
nand UO_2913 (O_2913,N_28952,N_28814);
and UO_2914 (O_2914,N_29036,N_29614);
and UO_2915 (O_2915,N_29547,N_29857);
nor UO_2916 (O_2916,N_29509,N_29328);
and UO_2917 (O_2917,N_29524,N_29690);
nor UO_2918 (O_2918,N_29211,N_29155);
and UO_2919 (O_2919,N_28884,N_29892);
nor UO_2920 (O_2920,N_29712,N_29956);
or UO_2921 (O_2921,N_29374,N_29830);
and UO_2922 (O_2922,N_29527,N_29509);
nand UO_2923 (O_2923,N_29203,N_29797);
xnor UO_2924 (O_2924,N_28855,N_29355);
xor UO_2925 (O_2925,N_29991,N_29684);
nand UO_2926 (O_2926,N_29484,N_29921);
nor UO_2927 (O_2927,N_29496,N_29885);
nor UO_2928 (O_2928,N_29186,N_29625);
nand UO_2929 (O_2929,N_29941,N_29232);
nor UO_2930 (O_2930,N_29253,N_29433);
or UO_2931 (O_2931,N_29039,N_28909);
xnor UO_2932 (O_2932,N_29479,N_29012);
xor UO_2933 (O_2933,N_29736,N_29649);
or UO_2934 (O_2934,N_28945,N_29445);
and UO_2935 (O_2935,N_28995,N_29026);
nand UO_2936 (O_2936,N_29687,N_29812);
nand UO_2937 (O_2937,N_28968,N_28932);
nor UO_2938 (O_2938,N_29596,N_29154);
and UO_2939 (O_2939,N_29402,N_28913);
nand UO_2940 (O_2940,N_28822,N_29350);
and UO_2941 (O_2941,N_29936,N_29248);
or UO_2942 (O_2942,N_29824,N_29375);
and UO_2943 (O_2943,N_29438,N_28989);
nand UO_2944 (O_2944,N_29993,N_29866);
xor UO_2945 (O_2945,N_29534,N_29871);
xnor UO_2946 (O_2946,N_29572,N_28992);
nor UO_2947 (O_2947,N_29006,N_28846);
xnor UO_2948 (O_2948,N_28874,N_29671);
nand UO_2949 (O_2949,N_29704,N_29457);
and UO_2950 (O_2950,N_29943,N_28948);
and UO_2951 (O_2951,N_29552,N_29012);
xor UO_2952 (O_2952,N_29524,N_29330);
nor UO_2953 (O_2953,N_29087,N_29311);
xor UO_2954 (O_2954,N_28872,N_29278);
and UO_2955 (O_2955,N_29319,N_29671);
and UO_2956 (O_2956,N_29886,N_28841);
and UO_2957 (O_2957,N_29112,N_29840);
or UO_2958 (O_2958,N_29887,N_29598);
nor UO_2959 (O_2959,N_29587,N_29862);
xnor UO_2960 (O_2960,N_28918,N_28861);
or UO_2961 (O_2961,N_29868,N_29973);
and UO_2962 (O_2962,N_29603,N_29363);
nand UO_2963 (O_2963,N_29335,N_29662);
xor UO_2964 (O_2964,N_29274,N_29868);
and UO_2965 (O_2965,N_29240,N_29226);
or UO_2966 (O_2966,N_29878,N_29636);
and UO_2967 (O_2967,N_29904,N_29834);
and UO_2968 (O_2968,N_29470,N_29535);
xnor UO_2969 (O_2969,N_29526,N_29581);
xnor UO_2970 (O_2970,N_29646,N_28922);
xor UO_2971 (O_2971,N_29016,N_29044);
nand UO_2972 (O_2972,N_28803,N_29087);
or UO_2973 (O_2973,N_28889,N_29826);
nor UO_2974 (O_2974,N_29701,N_29729);
nor UO_2975 (O_2975,N_29714,N_29439);
xor UO_2976 (O_2976,N_28809,N_28904);
nor UO_2977 (O_2977,N_29776,N_29839);
or UO_2978 (O_2978,N_29464,N_28848);
nor UO_2979 (O_2979,N_29169,N_29948);
or UO_2980 (O_2980,N_29280,N_29513);
nor UO_2981 (O_2981,N_29876,N_29472);
and UO_2982 (O_2982,N_29277,N_29335);
nor UO_2983 (O_2983,N_28967,N_28964);
or UO_2984 (O_2984,N_29767,N_29735);
xnor UO_2985 (O_2985,N_28900,N_28989);
and UO_2986 (O_2986,N_28895,N_29728);
xnor UO_2987 (O_2987,N_29195,N_29797);
nor UO_2988 (O_2988,N_28953,N_29387);
or UO_2989 (O_2989,N_29545,N_29810);
or UO_2990 (O_2990,N_29637,N_29666);
nor UO_2991 (O_2991,N_29062,N_29054);
and UO_2992 (O_2992,N_29871,N_29385);
nor UO_2993 (O_2993,N_28914,N_28992);
and UO_2994 (O_2994,N_29637,N_28860);
nor UO_2995 (O_2995,N_29011,N_29403);
or UO_2996 (O_2996,N_28966,N_28856);
nand UO_2997 (O_2997,N_29284,N_29727);
xor UO_2998 (O_2998,N_29887,N_29998);
xor UO_2999 (O_2999,N_28921,N_29056);
nor UO_3000 (O_3000,N_28902,N_29229);
nand UO_3001 (O_3001,N_29971,N_29928);
and UO_3002 (O_3002,N_29516,N_28972);
or UO_3003 (O_3003,N_29473,N_29174);
nand UO_3004 (O_3004,N_29256,N_28842);
and UO_3005 (O_3005,N_29728,N_29425);
nand UO_3006 (O_3006,N_29294,N_28994);
nand UO_3007 (O_3007,N_29724,N_29146);
nor UO_3008 (O_3008,N_29814,N_29514);
xnor UO_3009 (O_3009,N_29564,N_29821);
or UO_3010 (O_3010,N_29618,N_29380);
xor UO_3011 (O_3011,N_29643,N_28992);
nor UO_3012 (O_3012,N_29464,N_28805);
and UO_3013 (O_3013,N_29196,N_28857);
and UO_3014 (O_3014,N_29791,N_29840);
xnor UO_3015 (O_3015,N_29300,N_29530);
or UO_3016 (O_3016,N_29652,N_29676);
or UO_3017 (O_3017,N_29703,N_29774);
and UO_3018 (O_3018,N_28871,N_29486);
and UO_3019 (O_3019,N_29446,N_29274);
and UO_3020 (O_3020,N_29221,N_29386);
nor UO_3021 (O_3021,N_29130,N_28949);
and UO_3022 (O_3022,N_29027,N_28851);
and UO_3023 (O_3023,N_29419,N_29274);
nand UO_3024 (O_3024,N_29882,N_29238);
and UO_3025 (O_3025,N_29532,N_29805);
and UO_3026 (O_3026,N_29749,N_29161);
nor UO_3027 (O_3027,N_29489,N_28982);
and UO_3028 (O_3028,N_28890,N_29602);
xor UO_3029 (O_3029,N_29592,N_29533);
or UO_3030 (O_3030,N_29105,N_29460);
nor UO_3031 (O_3031,N_29863,N_29157);
and UO_3032 (O_3032,N_28840,N_29996);
or UO_3033 (O_3033,N_29713,N_29400);
or UO_3034 (O_3034,N_29134,N_29678);
nand UO_3035 (O_3035,N_29416,N_29937);
or UO_3036 (O_3036,N_29635,N_29540);
or UO_3037 (O_3037,N_29041,N_29560);
xnor UO_3038 (O_3038,N_29862,N_29677);
xnor UO_3039 (O_3039,N_28920,N_29887);
or UO_3040 (O_3040,N_29372,N_29714);
xor UO_3041 (O_3041,N_28886,N_29332);
and UO_3042 (O_3042,N_29219,N_29073);
nand UO_3043 (O_3043,N_29993,N_28999);
and UO_3044 (O_3044,N_29810,N_29235);
nor UO_3045 (O_3045,N_29005,N_29332);
nand UO_3046 (O_3046,N_29002,N_28878);
nand UO_3047 (O_3047,N_29107,N_29962);
and UO_3048 (O_3048,N_28997,N_29732);
and UO_3049 (O_3049,N_29641,N_29036);
or UO_3050 (O_3050,N_29459,N_29989);
xnor UO_3051 (O_3051,N_29693,N_29438);
xnor UO_3052 (O_3052,N_29001,N_29366);
and UO_3053 (O_3053,N_29816,N_29391);
nor UO_3054 (O_3054,N_29417,N_29291);
and UO_3055 (O_3055,N_29596,N_29440);
xnor UO_3056 (O_3056,N_29930,N_29323);
xnor UO_3057 (O_3057,N_29992,N_29422);
nand UO_3058 (O_3058,N_28924,N_28977);
or UO_3059 (O_3059,N_29440,N_29076);
or UO_3060 (O_3060,N_29404,N_29248);
and UO_3061 (O_3061,N_29978,N_29575);
and UO_3062 (O_3062,N_28955,N_29973);
or UO_3063 (O_3063,N_29218,N_29267);
and UO_3064 (O_3064,N_29122,N_29388);
xnor UO_3065 (O_3065,N_29555,N_29048);
or UO_3066 (O_3066,N_29612,N_28928);
nor UO_3067 (O_3067,N_28972,N_29103);
nor UO_3068 (O_3068,N_29243,N_28955);
nand UO_3069 (O_3069,N_29390,N_28886);
nor UO_3070 (O_3070,N_29476,N_29214);
or UO_3071 (O_3071,N_29156,N_28846);
xnor UO_3072 (O_3072,N_29945,N_28850);
xnor UO_3073 (O_3073,N_29564,N_29017);
xnor UO_3074 (O_3074,N_29908,N_29062);
nor UO_3075 (O_3075,N_29593,N_29481);
nor UO_3076 (O_3076,N_28850,N_29585);
xnor UO_3077 (O_3077,N_29243,N_29098);
nand UO_3078 (O_3078,N_29740,N_29517);
or UO_3079 (O_3079,N_29783,N_29186);
or UO_3080 (O_3080,N_29451,N_28947);
nor UO_3081 (O_3081,N_29089,N_29259);
or UO_3082 (O_3082,N_29121,N_29285);
nand UO_3083 (O_3083,N_29669,N_29684);
nor UO_3084 (O_3084,N_29882,N_29310);
nor UO_3085 (O_3085,N_29516,N_29781);
nand UO_3086 (O_3086,N_29201,N_29927);
or UO_3087 (O_3087,N_29046,N_29665);
and UO_3088 (O_3088,N_28829,N_29437);
and UO_3089 (O_3089,N_28950,N_29757);
nor UO_3090 (O_3090,N_29699,N_29423);
or UO_3091 (O_3091,N_29085,N_29990);
nand UO_3092 (O_3092,N_28950,N_29430);
nor UO_3093 (O_3093,N_29684,N_29721);
xnor UO_3094 (O_3094,N_29440,N_28846);
or UO_3095 (O_3095,N_29572,N_29826);
xor UO_3096 (O_3096,N_28800,N_29987);
and UO_3097 (O_3097,N_28929,N_28847);
xnor UO_3098 (O_3098,N_29007,N_29772);
and UO_3099 (O_3099,N_29795,N_29586);
nand UO_3100 (O_3100,N_28816,N_29991);
and UO_3101 (O_3101,N_29683,N_29408);
and UO_3102 (O_3102,N_29255,N_29167);
xor UO_3103 (O_3103,N_29036,N_29246);
nor UO_3104 (O_3104,N_29716,N_29086);
nor UO_3105 (O_3105,N_29828,N_29790);
xor UO_3106 (O_3106,N_28835,N_29285);
and UO_3107 (O_3107,N_29506,N_29992);
xnor UO_3108 (O_3108,N_29545,N_29943);
and UO_3109 (O_3109,N_29164,N_29827);
nor UO_3110 (O_3110,N_29572,N_29172);
nand UO_3111 (O_3111,N_29567,N_29784);
or UO_3112 (O_3112,N_29167,N_29773);
xnor UO_3113 (O_3113,N_28885,N_29483);
xnor UO_3114 (O_3114,N_29358,N_28888);
xor UO_3115 (O_3115,N_29853,N_29310);
nand UO_3116 (O_3116,N_29526,N_29147);
or UO_3117 (O_3117,N_29460,N_29289);
or UO_3118 (O_3118,N_29354,N_29017);
xor UO_3119 (O_3119,N_29758,N_29617);
nor UO_3120 (O_3120,N_29789,N_28935);
and UO_3121 (O_3121,N_28808,N_29910);
xor UO_3122 (O_3122,N_29035,N_29377);
or UO_3123 (O_3123,N_29021,N_29918);
nand UO_3124 (O_3124,N_29954,N_28873);
nand UO_3125 (O_3125,N_29821,N_28857);
nand UO_3126 (O_3126,N_29042,N_29983);
and UO_3127 (O_3127,N_29542,N_29081);
nand UO_3128 (O_3128,N_29044,N_29227);
xnor UO_3129 (O_3129,N_29111,N_29139);
nor UO_3130 (O_3130,N_29483,N_29691);
xnor UO_3131 (O_3131,N_29868,N_29827);
xor UO_3132 (O_3132,N_29068,N_28851);
nand UO_3133 (O_3133,N_28950,N_29822);
or UO_3134 (O_3134,N_28866,N_29671);
or UO_3135 (O_3135,N_29884,N_28821);
nand UO_3136 (O_3136,N_28966,N_28817);
or UO_3137 (O_3137,N_29856,N_29291);
xnor UO_3138 (O_3138,N_29341,N_29547);
and UO_3139 (O_3139,N_29957,N_29204);
xor UO_3140 (O_3140,N_29783,N_28979);
or UO_3141 (O_3141,N_28838,N_29869);
or UO_3142 (O_3142,N_28923,N_29477);
and UO_3143 (O_3143,N_29406,N_29368);
nand UO_3144 (O_3144,N_29593,N_29766);
and UO_3145 (O_3145,N_29287,N_29775);
nor UO_3146 (O_3146,N_29883,N_28868);
or UO_3147 (O_3147,N_29564,N_29966);
or UO_3148 (O_3148,N_29683,N_29231);
nand UO_3149 (O_3149,N_28923,N_29499);
or UO_3150 (O_3150,N_29624,N_29276);
nand UO_3151 (O_3151,N_29525,N_29418);
xor UO_3152 (O_3152,N_29038,N_28929);
or UO_3153 (O_3153,N_29024,N_28990);
nor UO_3154 (O_3154,N_29729,N_29182);
nand UO_3155 (O_3155,N_29792,N_29273);
xor UO_3156 (O_3156,N_28832,N_29951);
xnor UO_3157 (O_3157,N_29489,N_29467);
nor UO_3158 (O_3158,N_29271,N_28883);
and UO_3159 (O_3159,N_29338,N_29943);
nor UO_3160 (O_3160,N_29368,N_29859);
or UO_3161 (O_3161,N_29385,N_29485);
nand UO_3162 (O_3162,N_29905,N_29177);
nor UO_3163 (O_3163,N_29494,N_29105);
nand UO_3164 (O_3164,N_29283,N_28825);
nand UO_3165 (O_3165,N_29955,N_29186);
nand UO_3166 (O_3166,N_29486,N_29506);
nand UO_3167 (O_3167,N_29387,N_29742);
xnor UO_3168 (O_3168,N_28801,N_29514);
and UO_3169 (O_3169,N_28939,N_29709);
and UO_3170 (O_3170,N_29706,N_29966);
nor UO_3171 (O_3171,N_29332,N_29383);
and UO_3172 (O_3172,N_29713,N_29578);
nand UO_3173 (O_3173,N_28884,N_29490);
nor UO_3174 (O_3174,N_29668,N_28897);
nor UO_3175 (O_3175,N_29041,N_29515);
xor UO_3176 (O_3176,N_29254,N_29638);
and UO_3177 (O_3177,N_28974,N_29929);
xor UO_3178 (O_3178,N_29553,N_28862);
and UO_3179 (O_3179,N_29622,N_29642);
nor UO_3180 (O_3180,N_29575,N_28809);
nand UO_3181 (O_3181,N_29303,N_29913);
nand UO_3182 (O_3182,N_29786,N_29326);
nor UO_3183 (O_3183,N_29870,N_29123);
nand UO_3184 (O_3184,N_29441,N_28884);
xnor UO_3185 (O_3185,N_29400,N_29609);
xnor UO_3186 (O_3186,N_29881,N_29148);
nor UO_3187 (O_3187,N_29177,N_29985);
or UO_3188 (O_3188,N_28826,N_29866);
nand UO_3189 (O_3189,N_29001,N_28817);
nand UO_3190 (O_3190,N_29070,N_29644);
or UO_3191 (O_3191,N_28886,N_29767);
nand UO_3192 (O_3192,N_29470,N_29385);
xor UO_3193 (O_3193,N_29781,N_29919);
nand UO_3194 (O_3194,N_29507,N_28987);
or UO_3195 (O_3195,N_29264,N_29351);
nand UO_3196 (O_3196,N_28850,N_29919);
nand UO_3197 (O_3197,N_28832,N_28878);
nor UO_3198 (O_3198,N_28906,N_29440);
nor UO_3199 (O_3199,N_29002,N_29400);
nor UO_3200 (O_3200,N_29610,N_29096);
nor UO_3201 (O_3201,N_28959,N_29945);
and UO_3202 (O_3202,N_29002,N_29240);
nor UO_3203 (O_3203,N_29176,N_29381);
xor UO_3204 (O_3204,N_29846,N_29168);
xor UO_3205 (O_3205,N_29540,N_29517);
or UO_3206 (O_3206,N_29035,N_28885);
xor UO_3207 (O_3207,N_29860,N_29316);
and UO_3208 (O_3208,N_29885,N_29610);
nand UO_3209 (O_3209,N_29131,N_28862);
nor UO_3210 (O_3210,N_29666,N_29625);
xor UO_3211 (O_3211,N_29287,N_29185);
and UO_3212 (O_3212,N_29343,N_29432);
and UO_3213 (O_3213,N_29683,N_28956);
xnor UO_3214 (O_3214,N_29662,N_29655);
nand UO_3215 (O_3215,N_29353,N_29585);
xnor UO_3216 (O_3216,N_29041,N_29829);
nand UO_3217 (O_3217,N_29436,N_29224);
or UO_3218 (O_3218,N_29468,N_29403);
nand UO_3219 (O_3219,N_28807,N_29763);
nand UO_3220 (O_3220,N_29861,N_29653);
and UO_3221 (O_3221,N_29575,N_29642);
nand UO_3222 (O_3222,N_29785,N_29614);
xor UO_3223 (O_3223,N_29927,N_29955);
xor UO_3224 (O_3224,N_29322,N_29113);
xor UO_3225 (O_3225,N_29945,N_29383);
xor UO_3226 (O_3226,N_29922,N_29310);
xor UO_3227 (O_3227,N_28971,N_29147);
nand UO_3228 (O_3228,N_29545,N_29132);
and UO_3229 (O_3229,N_29669,N_29330);
and UO_3230 (O_3230,N_29176,N_29432);
or UO_3231 (O_3231,N_29192,N_29369);
or UO_3232 (O_3232,N_29598,N_29396);
and UO_3233 (O_3233,N_29663,N_29966);
nor UO_3234 (O_3234,N_29583,N_29018);
nand UO_3235 (O_3235,N_29102,N_29964);
nor UO_3236 (O_3236,N_29678,N_29255);
nand UO_3237 (O_3237,N_29595,N_29262);
nor UO_3238 (O_3238,N_29175,N_29460);
or UO_3239 (O_3239,N_29736,N_29509);
xnor UO_3240 (O_3240,N_29265,N_29841);
nand UO_3241 (O_3241,N_29923,N_29010);
or UO_3242 (O_3242,N_29971,N_29055);
and UO_3243 (O_3243,N_29916,N_29310);
xor UO_3244 (O_3244,N_29034,N_29067);
xor UO_3245 (O_3245,N_29929,N_28830);
and UO_3246 (O_3246,N_28940,N_28953);
or UO_3247 (O_3247,N_29391,N_29596);
nor UO_3248 (O_3248,N_28888,N_29438);
or UO_3249 (O_3249,N_28885,N_29322);
and UO_3250 (O_3250,N_29661,N_28947);
and UO_3251 (O_3251,N_29650,N_29726);
and UO_3252 (O_3252,N_29089,N_29397);
nand UO_3253 (O_3253,N_28804,N_29289);
or UO_3254 (O_3254,N_28994,N_29074);
nand UO_3255 (O_3255,N_29481,N_29060);
nand UO_3256 (O_3256,N_29564,N_29927);
or UO_3257 (O_3257,N_29157,N_29086);
nor UO_3258 (O_3258,N_28803,N_29678);
nor UO_3259 (O_3259,N_29567,N_29461);
and UO_3260 (O_3260,N_29968,N_29579);
nor UO_3261 (O_3261,N_29914,N_29599);
nor UO_3262 (O_3262,N_29695,N_29440);
nor UO_3263 (O_3263,N_29142,N_29017);
nand UO_3264 (O_3264,N_29033,N_29866);
xnor UO_3265 (O_3265,N_29132,N_29501);
nand UO_3266 (O_3266,N_29347,N_29503);
and UO_3267 (O_3267,N_28977,N_29126);
xnor UO_3268 (O_3268,N_29419,N_29257);
nand UO_3269 (O_3269,N_29702,N_29571);
and UO_3270 (O_3270,N_28819,N_29855);
xor UO_3271 (O_3271,N_28956,N_29196);
nor UO_3272 (O_3272,N_29263,N_29903);
nand UO_3273 (O_3273,N_29671,N_29050);
nand UO_3274 (O_3274,N_28965,N_29595);
or UO_3275 (O_3275,N_29457,N_29991);
and UO_3276 (O_3276,N_28811,N_28984);
and UO_3277 (O_3277,N_29889,N_29836);
and UO_3278 (O_3278,N_29770,N_29210);
nor UO_3279 (O_3279,N_29278,N_28885);
or UO_3280 (O_3280,N_29654,N_29796);
or UO_3281 (O_3281,N_29076,N_29934);
xnor UO_3282 (O_3282,N_29078,N_29522);
or UO_3283 (O_3283,N_29788,N_29721);
and UO_3284 (O_3284,N_29336,N_29316);
xnor UO_3285 (O_3285,N_28942,N_29817);
nand UO_3286 (O_3286,N_29083,N_29103);
xor UO_3287 (O_3287,N_28960,N_28935);
or UO_3288 (O_3288,N_29434,N_29126);
nor UO_3289 (O_3289,N_29438,N_29086);
or UO_3290 (O_3290,N_29010,N_29143);
xor UO_3291 (O_3291,N_29100,N_29493);
or UO_3292 (O_3292,N_29163,N_29521);
or UO_3293 (O_3293,N_29451,N_29873);
and UO_3294 (O_3294,N_28924,N_29600);
and UO_3295 (O_3295,N_29606,N_29998);
nand UO_3296 (O_3296,N_28967,N_29002);
nand UO_3297 (O_3297,N_29278,N_28807);
or UO_3298 (O_3298,N_29861,N_29989);
or UO_3299 (O_3299,N_29860,N_29072);
nand UO_3300 (O_3300,N_29896,N_29162);
and UO_3301 (O_3301,N_29874,N_29833);
nand UO_3302 (O_3302,N_29951,N_29647);
nand UO_3303 (O_3303,N_28935,N_29379);
nor UO_3304 (O_3304,N_29067,N_28830);
xor UO_3305 (O_3305,N_29524,N_29241);
and UO_3306 (O_3306,N_29893,N_29989);
nor UO_3307 (O_3307,N_29015,N_29110);
nand UO_3308 (O_3308,N_28944,N_29113);
xnor UO_3309 (O_3309,N_29253,N_29945);
or UO_3310 (O_3310,N_29170,N_29250);
xor UO_3311 (O_3311,N_29782,N_29724);
nand UO_3312 (O_3312,N_29476,N_29808);
or UO_3313 (O_3313,N_29848,N_29080);
xnor UO_3314 (O_3314,N_29054,N_29986);
and UO_3315 (O_3315,N_29274,N_29166);
or UO_3316 (O_3316,N_29546,N_29563);
and UO_3317 (O_3317,N_29156,N_29451);
nor UO_3318 (O_3318,N_28822,N_29888);
nand UO_3319 (O_3319,N_28891,N_29862);
and UO_3320 (O_3320,N_29110,N_29776);
nor UO_3321 (O_3321,N_29421,N_29063);
and UO_3322 (O_3322,N_29500,N_29508);
nor UO_3323 (O_3323,N_28827,N_29377);
nor UO_3324 (O_3324,N_28884,N_29605);
or UO_3325 (O_3325,N_29887,N_29197);
nand UO_3326 (O_3326,N_29739,N_29200);
and UO_3327 (O_3327,N_29317,N_28812);
and UO_3328 (O_3328,N_29530,N_29066);
and UO_3329 (O_3329,N_29023,N_29373);
and UO_3330 (O_3330,N_28810,N_29096);
and UO_3331 (O_3331,N_29727,N_29294);
nand UO_3332 (O_3332,N_29373,N_29630);
or UO_3333 (O_3333,N_29509,N_29448);
xor UO_3334 (O_3334,N_29579,N_29219);
and UO_3335 (O_3335,N_28899,N_29723);
or UO_3336 (O_3336,N_29246,N_29975);
nor UO_3337 (O_3337,N_29298,N_29734);
nand UO_3338 (O_3338,N_29245,N_29134);
and UO_3339 (O_3339,N_29461,N_29282);
xor UO_3340 (O_3340,N_29554,N_28932);
xor UO_3341 (O_3341,N_29831,N_29955);
and UO_3342 (O_3342,N_29703,N_28825);
or UO_3343 (O_3343,N_29719,N_28896);
xnor UO_3344 (O_3344,N_29917,N_29158);
xnor UO_3345 (O_3345,N_29061,N_29225);
xor UO_3346 (O_3346,N_29734,N_29067);
or UO_3347 (O_3347,N_29706,N_29861);
nand UO_3348 (O_3348,N_29081,N_29571);
nor UO_3349 (O_3349,N_29051,N_29500);
nand UO_3350 (O_3350,N_29058,N_29135);
nor UO_3351 (O_3351,N_29687,N_28860);
xnor UO_3352 (O_3352,N_29903,N_29672);
xnor UO_3353 (O_3353,N_29381,N_29972);
nor UO_3354 (O_3354,N_29953,N_29518);
or UO_3355 (O_3355,N_28814,N_29459);
and UO_3356 (O_3356,N_29425,N_29248);
or UO_3357 (O_3357,N_28820,N_29892);
or UO_3358 (O_3358,N_29405,N_29561);
xnor UO_3359 (O_3359,N_29071,N_29781);
nor UO_3360 (O_3360,N_29055,N_29430);
or UO_3361 (O_3361,N_29819,N_29828);
xnor UO_3362 (O_3362,N_29151,N_28822);
nor UO_3363 (O_3363,N_29515,N_28856);
nand UO_3364 (O_3364,N_29484,N_29251);
nand UO_3365 (O_3365,N_29764,N_29946);
nand UO_3366 (O_3366,N_29632,N_29428);
nor UO_3367 (O_3367,N_28940,N_29015);
xor UO_3368 (O_3368,N_29401,N_29322);
and UO_3369 (O_3369,N_29704,N_29689);
and UO_3370 (O_3370,N_29435,N_29124);
xor UO_3371 (O_3371,N_29454,N_28862);
nand UO_3372 (O_3372,N_29599,N_29550);
or UO_3373 (O_3373,N_28846,N_29866);
nand UO_3374 (O_3374,N_29481,N_29563);
and UO_3375 (O_3375,N_28889,N_29883);
nor UO_3376 (O_3376,N_28964,N_28850);
xnor UO_3377 (O_3377,N_29523,N_29465);
or UO_3378 (O_3378,N_29793,N_29071);
xor UO_3379 (O_3379,N_29802,N_28941);
xnor UO_3380 (O_3380,N_28830,N_29692);
or UO_3381 (O_3381,N_29736,N_29241);
xnor UO_3382 (O_3382,N_29489,N_29049);
nor UO_3383 (O_3383,N_29692,N_28954);
and UO_3384 (O_3384,N_29828,N_29529);
or UO_3385 (O_3385,N_28955,N_29023);
or UO_3386 (O_3386,N_29613,N_29276);
nor UO_3387 (O_3387,N_28900,N_29789);
and UO_3388 (O_3388,N_29377,N_29681);
nor UO_3389 (O_3389,N_29685,N_29512);
nand UO_3390 (O_3390,N_29841,N_29588);
nor UO_3391 (O_3391,N_29409,N_29370);
and UO_3392 (O_3392,N_29973,N_29081);
and UO_3393 (O_3393,N_28887,N_29176);
nand UO_3394 (O_3394,N_29989,N_29539);
xor UO_3395 (O_3395,N_28877,N_29342);
or UO_3396 (O_3396,N_29130,N_29517);
xnor UO_3397 (O_3397,N_28944,N_28878);
or UO_3398 (O_3398,N_29964,N_29210);
nand UO_3399 (O_3399,N_28802,N_29189);
and UO_3400 (O_3400,N_29358,N_29957);
xnor UO_3401 (O_3401,N_29988,N_29691);
or UO_3402 (O_3402,N_29978,N_29408);
nand UO_3403 (O_3403,N_28814,N_29611);
nor UO_3404 (O_3404,N_29778,N_29153);
and UO_3405 (O_3405,N_29900,N_29040);
or UO_3406 (O_3406,N_29820,N_29067);
nor UO_3407 (O_3407,N_28935,N_29756);
nand UO_3408 (O_3408,N_29664,N_29679);
nand UO_3409 (O_3409,N_29823,N_29407);
or UO_3410 (O_3410,N_28918,N_28967);
nand UO_3411 (O_3411,N_29046,N_29735);
nand UO_3412 (O_3412,N_29395,N_28868);
nor UO_3413 (O_3413,N_29954,N_29703);
nand UO_3414 (O_3414,N_29494,N_29806);
nand UO_3415 (O_3415,N_29021,N_29543);
nor UO_3416 (O_3416,N_29234,N_29303);
or UO_3417 (O_3417,N_29397,N_29927);
nor UO_3418 (O_3418,N_29019,N_29967);
nor UO_3419 (O_3419,N_29434,N_29464);
nand UO_3420 (O_3420,N_29650,N_29137);
and UO_3421 (O_3421,N_29405,N_29827);
or UO_3422 (O_3422,N_29594,N_29556);
or UO_3423 (O_3423,N_29066,N_29212);
xnor UO_3424 (O_3424,N_29898,N_28881);
or UO_3425 (O_3425,N_29909,N_29677);
xnor UO_3426 (O_3426,N_29953,N_29557);
nand UO_3427 (O_3427,N_29087,N_29634);
nand UO_3428 (O_3428,N_29389,N_28940);
nor UO_3429 (O_3429,N_29150,N_29643);
nor UO_3430 (O_3430,N_29742,N_29252);
or UO_3431 (O_3431,N_29462,N_29222);
xnor UO_3432 (O_3432,N_29065,N_28850);
nor UO_3433 (O_3433,N_29214,N_29294);
nor UO_3434 (O_3434,N_28981,N_29925);
nand UO_3435 (O_3435,N_29843,N_29710);
xor UO_3436 (O_3436,N_29769,N_29400);
nand UO_3437 (O_3437,N_28865,N_29607);
nor UO_3438 (O_3438,N_28860,N_29154);
or UO_3439 (O_3439,N_29348,N_29680);
or UO_3440 (O_3440,N_29713,N_29299);
nand UO_3441 (O_3441,N_29357,N_29703);
nand UO_3442 (O_3442,N_29361,N_28880);
nor UO_3443 (O_3443,N_28892,N_28835);
nand UO_3444 (O_3444,N_28898,N_29594);
xor UO_3445 (O_3445,N_29862,N_29107);
xor UO_3446 (O_3446,N_29323,N_29396);
xnor UO_3447 (O_3447,N_29449,N_29978);
or UO_3448 (O_3448,N_29781,N_29343);
or UO_3449 (O_3449,N_29363,N_29536);
or UO_3450 (O_3450,N_29385,N_29315);
and UO_3451 (O_3451,N_29724,N_29316);
nor UO_3452 (O_3452,N_29666,N_29597);
nand UO_3453 (O_3453,N_29041,N_29734);
nor UO_3454 (O_3454,N_29168,N_29487);
nor UO_3455 (O_3455,N_29996,N_29495);
nor UO_3456 (O_3456,N_29787,N_29850);
or UO_3457 (O_3457,N_29703,N_28874);
and UO_3458 (O_3458,N_29056,N_29963);
nand UO_3459 (O_3459,N_29425,N_28902);
xor UO_3460 (O_3460,N_29735,N_29968);
xnor UO_3461 (O_3461,N_29120,N_29968);
nand UO_3462 (O_3462,N_29284,N_29186);
nand UO_3463 (O_3463,N_29678,N_28939);
nor UO_3464 (O_3464,N_28961,N_29888);
xor UO_3465 (O_3465,N_29608,N_29631);
and UO_3466 (O_3466,N_28822,N_29669);
and UO_3467 (O_3467,N_28945,N_29884);
nand UO_3468 (O_3468,N_28983,N_29973);
or UO_3469 (O_3469,N_29215,N_29116);
xor UO_3470 (O_3470,N_28865,N_29390);
or UO_3471 (O_3471,N_29818,N_29081);
nor UO_3472 (O_3472,N_29568,N_29801);
nand UO_3473 (O_3473,N_29844,N_29733);
nor UO_3474 (O_3474,N_28844,N_28942);
xor UO_3475 (O_3475,N_29571,N_29012);
and UO_3476 (O_3476,N_29031,N_29424);
or UO_3477 (O_3477,N_29618,N_29811);
nand UO_3478 (O_3478,N_29652,N_28898);
nor UO_3479 (O_3479,N_28949,N_28856);
and UO_3480 (O_3480,N_29215,N_29463);
and UO_3481 (O_3481,N_29468,N_29014);
and UO_3482 (O_3482,N_29126,N_29808);
and UO_3483 (O_3483,N_29548,N_28977);
and UO_3484 (O_3484,N_29252,N_28923);
nand UO_3485 (O_3485,N_28859,N_29757);
nand UO_3486 (O_3486,N_28994,N_29040);
xnor UO_3487 (O_3487,N_29848,N_29448);
nand UO_3488 (O_3488,N_29903,N_29481);
and UO_3489 (O_3489,N_29828,N_28986);
and UO_3490 (O_3490,N_29663,N_29421);
nor UO_3491 (O_3491,N_28822,N_29864);
or UO_3492 (O_3492,N_29857,N_28848);
nor UO_3493 (O_3493,N_29815,N_29794);
nand UO_3494 (O_3494,N_29185,N_28933);
or UO_3495 (O_3495,N_28816,N_29282);
nor UO_3496 (O_3496,N_29094,N_29070);
xnor UO_3497 (O_3497,N_29262,N_29472);
nand UO_3498 (O_3498,N_29461,N_29867);
nand UO_3499 (O_3499,N_29783,N_29644);
endmodule