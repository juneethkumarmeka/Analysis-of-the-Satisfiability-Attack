module basic_1000_10000_1500_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_426,In_744);
nand U1 (N_1,In_55,In_781);
nor U2 (N_2,In_284,In_899);
and U3 (N_3,In_699,In_446);
nor U4 (N_4,In_346,In_754);
or U5 (N_5,In_871,In_670);
and U6 (N_6,In_339,In_789);
nor U7 (N_7,In_958,In_610);
nand U8 (N_8,In_255,In_440);
or U9 (N_9,In_896,In_413);
and U10 (N_10,In_411,In_712);
or U11 (N_11,In_756,In_315);
nand U12 (N_12,In_246,In_589);
or U13 (N_13,In_567,In_456);
nand U14 (N_14,In_115,In_476);
nor U15 (N_15,In_356,In_907);
nand U16 (N_16,In_412,In_340);
or U17 (N_17,In_29,In_478);
nor U18 (N_18,In_70,In_777);
nand U19 (N_19,In_10,In_89);
and U20 (N_20,In_92,In_441);
nand U21 (N_21,In_759,In_853);
and U22 (N_22,In_883,In_435);
nand U23 (N_23,In_1,In_826);
nor U24 (N_24,In_725,In_336);
or U25 (N_25,In_602,In_144);
nor U26 (N_26,In_214,In_547);
and U27 (N_27,In_4,In_893);
nand U28 (N_28,In_205,In_686);
or U29 (N_29,In_731,In_785);
or U30 (N_30,In_50,In_382);
nor U31 (N_31,In_981,In_180);
nor U32 (N_32,In_943,In_778);
nand U33 (N_33,In_287,In_911);
nand U34 (N_34,In_835,In_854);
nor U35 (N_35,In_424,In_662);
or U36 (N_36,In_692,In_519);
nor U37 (N_37,In_836,In_822);
xnor U38 (N_38,In_88,In_949);
nand U39 (N_39,In_128,In_698);
and U40 (N_40,In_261,In_782);
nand U41 (N_41,In_733,In_251);
or U42 (N_42,In_280,In_809);
and U43 (N_43,In_528,In_347);
and U44 (N_44,In_929,In_245);
and U45 (N_45,In_930,In_653);
or U46 (N_46,In_950,In_217);
nor U47 (N_47,In_565,In_114);
or U48 (N_48,In_8,In_860);
or U49 (N_49,In_450,In_558);
or U50 (N_50,In_700,In_104);
and U51 (N_51,In_442,In_574);
xnor U52 (N_52,In_223,In_649);
nor U53 (N_53,In_44,In_397);
nor U54 (N_54,In_269,In_617);
nand U55 (N_55,In_975,In_242);
nand U56 (N_56,In_608,In_869);
nand U57 (N_57,In_443,In_827);
and U58 (N_58,In_609,In_654);
nand U59 (N_59,In_579,In_38);
xnor U60 (N_60,In_576,In_429);
nand U61 (N_61,In_120,In_906);
or U62 (N_62,In_961,In_679);
or U63 (N_63,In_655,In_297);
nand U64 (N_64,In_239,In_454);
and U65 (N_65,In_630,In_518);
nor U66 (N_66,In_714,In_695);
nand U67 (N_67,In_267,In_509);
and U68 (N_68,In_228,In_514);
nand U69 (N_69,In_867,In_345);
and U70 (N_70,In_438,In_858);
and U71 (N_71,In_485,In_362);
or U72 (N_72,In_365,In_36);
and U73 (N_73,In_274,In_475);
or U74 (N_74,In_585,In_783);
or U75 (N_75,In_322,In_933);
or U76 (N_76,In_618,In_647);
nor U77 (N_77,In_290,In_221);
nand U78 (N_78,In_760,In_53);
and U79 (N_79,In_934,In_195);
or U80 (N_80,In_371,In_999);
nor U81 (N_81,In_821,In_806);
nand U82 (N_82,In_86,In_743);
xor U83 (N_83,In_123,In_747);
or U84 (N_84,In_801,In_220);
or U85 (N_85,In_148,In_741);
nor U86 (N_86,In_13,In_265);
nand U87 (N_87,In_517,In_661);
nand U88 (N_88,In_249,In_582);
xor U89 (N_89,In_663,In_2);
nor U90 (N_90,In_542,In_421);
or U91 (N_91,In_166,In_885);
nor U92 (N_92,In_215,In_384);
nor U93 (N_93,In_229,In_256);
nand U94 (N_94,In_570,In_562);
and U95 (N_95,In_73,In_40);
nor U96 (N_96,In_449,In_761);
nor U97 (N_97,In_24,In_736);
nor U98 (N_98,In_738,In_804);
nand U99 (N_99,In_82,In_259);
and U100 (N_100,In_203,In_786);
nor U101 (N_101,In_49,In_717);
and U102 (N_102,In_814,In_237);
xor U103 (N_103,In_489,In_665);
and U104 (N_104,In_206,In_524);
or U105 (N_105,In_468,In_726);
nor U106 (N_106,In_427,In_829);
xnor U107 (N_107,In_176,In_664);
nor U108 (N_108,In_138,In_409);
nor U109 (N_109,In_728,In_320);
nand U110 (N_110,In_296,In_982);
nand U111 (N_111,In_666,In_291);
nor U112 (N_112,In_130,In_191);
nor U113 (N_113,In_887,In_85);
or U114 (N_114,In_26,In_812);
xnor U115 (N_115,In_964,In_878);
nand U116 (N_116,In_306,In_299);
and U117 (N_117,In_75,In_625);
or U118 (N_118,In_637,In_6);
or U119 (N_119,In_233,In_58);
nor U120 (N_120,In_57,In_54);
nand U121 (N_121,In_861,In_658);
and U122 (N_122,In_374,In_11);
nand U123 (N_123,In_67,In_156);
nor U124 (N_124,In_210,In_711);
and U125 (N_125,In_335,In_369);
nor U126 (N_126,In_399,In_522);
nor U127 (N_127,In_243,In_897);
or U128 (N_128,In_250,In_834);
xor U129 (N_129,In_419,In_710);
xor U130 (N_130,In_707,In_83);
and U131 (N_131,In_702,In_61);
and U132 (N_132,In_740,In_616);
or U133 (N_133,In_72,In_453);
xor U134 (N_134,In_311,In_690);
or U135 (N_135,In_671,In_175);
or U136 (N_136,In_76,In_687);
or U137 (N_137,In_940,In_23);
nor U138 (N_138,In_792,In_207);
nand U139 (N_139,In_987,In_605);
nor U140 (N_140,In_656,In_624);
nor U141 (N_141,In_795,In_776);
nor U142 (N_142,In_500,In_392);
and U143 (N_143,In_141,In_640);
nand U144 (N_144,In_373,In_969);
nor U145 (N_145,In_723,In_404);
nor U146 (N_146,In_877,In_62);
or U147 (N_147,In_462,In_437);
nor U148 (N_148,In_937,In_847);
or U149 (N_149,In_729,In_708);
nand U150 (N_150,In_739,In_995);
nor U151 (N_151,In_414,In_200);
nor U152 (N_152,In_888,In_416);
or U153 (N_153,In_954,In_660);
nand U154 (N_154,In_116,In_641);
xnor U155 (N_155,In_722,In_455);
nand U156 (N_156,In_842,In_719);
xnor U157 (N_157,In_534,In_587);
nor U158 (N_158,In_946,In_535);
nand U159 (N_159,In_241,In_721);
nand U160 (N_160,In_967,In_797);
nor U161 (N_161,In_387,In_828);
nor U162 (N_162,In_63,In_359);
nor U163 (N_163,In_257,In_963);
or U164 (N_164,In_160,In_928);
or U165 (N_165,In_881,In_368);
and U166 (N_166,In_18,In_650);
xnor U167 (N_167,In_216,In_941);
xor U168 (N_168,In_155,In_140);
and U169 (N_169,In_876,In_80);
nor U170 (N_170,In_499,In_919);
or U171 (N_171,In_389,In_715);
or U172 (N_172,In_56,In_282);
nand U173 (N_173,In_95,In_504);
or U174 (N_174,In_332,In_613);
and U175 (N_175,In_927,In_596);
nor U176 (N_176,In_774,In_109);
nor U177 (N_177,In_799,In_263);
or U178 (N_178,In_457,In_966);
nand U179 (N_179,In_298,In_451);
or U180 (N_180,In_681,In_218);
and U181 (N_181,In_396,In_619);
or U182 (N_182,In_187,In_669);
and U183 (N_183,In_198,In_595);
xnor U184 (N_184,In_601,In_846);
or U185 (N_185,In_60,In_16);
or U186 (N_186,In_43,In_150);
and U187 (N_187,In_763,In_945);
and U188 (N_188,In_341,In_693);
and U189 (N_189,In_0,In_9);
or U190 (N_190,In_568,In_922);
nor U191 (N_191,In_573,In_460);
nand U192 (N_192,In_372,In_734);
or U193 (N_193,In_172,In_467);
and U194 (N_194,In_968,In_764);
nand U195 (N_195,In_872,In_793);
nor U196 (N_196,In_64,In_353);
or U197 (N_197,In_90,In_386);
nor U198 (N_198,In_401,In_701);
nor U199 (N_199,In_349,In_973);
or U200 (N_200,In_807,In_262);
nand U201 (N_201,In_645,In_874);
and U202 (N_202,In_163,In_525);
nor U203 (N_203,In_182,In_638);
nor U204 (N_204,In_244,In_926);
nand U205 (N_205,In_361,In_121);
and U206 (N_206,In_886,In_375);
nor U207 (N_207,In_979,In_931);
and U208 (N_208,In_976,In_915);
nand U209 (N_209,In_612,In_580);
or U210 (N_210,In_755,In_985);
xnor U211 (N_211,In_321,In_838);
nand U212 (N_212,In_902,In_490);
or U213 (N_213,In_330,In_864);
nor U214 (N_214,In_21,In_66);
and U215 (N_215,In_683,In_192);
nor U216 (N_216,In_342,In_790);
or U217 (N_217,In_972,In_100);
nand U218 (N_218,In_498,In_91);
xnor U219 (N_219,In_94,In_594);
xor U220 (N_220,In_136,In_477);
and U221 (N_221,In_491,In_367);
nor U222 (N_222,In_993,In_572);
nor U223 (N_223,In_481,In_788);
nor U224 (N_224,In_96,In_178);
nor U225 (N_225,In_168,In_318);
and U226 (N_226,In_938,In_407);
nor U227 (N_227,In_844,In_448);
nor U228 (N_228,In_190,In_988);
and U229 (N_229,In_627,In_204);
or U230 (N_230,In_420,In_151);
and U231 (N_231,In_74,In_388);
nor U232 (N_232,In_366,In_541);
or U233 (N_233,In_808,In_537);
or U234 (N_234,In_270,In_980);
nor U235 (N_235,In_415,In_157);
nand U236 (N_236,In_604,In_352);
nand U237 (N_237,In_620,In_286);
and U238 (N_238,In_557,In_532);
or U239 (N_239,In_87,In_227);
or U240 (N_240,In_3,In_402);
nand U241 (N_241,In_276,In_135);
nor U242 (N_242,In_14,In_873);
and U243 (N_243,In_521,In_564);
and U244 (N_244,In_948,In_264);
nand U245 (N_245,In_631,In_971);
nand U246 (N_246,In_780,In_493);
nand U247 (N_247,In_944,In_132);
nand U248 (N_248,In_566,In_615);
nand U249 (N_249,In_628,In_300);
nand U250 (N_250,In_578,In_603);
nor U251 (N_251,In_762,In_169);
and U252 (N_252,In_561,In_830);
xor U253 (N_253,In_600,In_184);
nand U254 (N_254,In_395,In_939);
nand U255 (N_255,In_817,In_212);
nand U256 (N_256,In_716,In_870);
and U257 (N_257,In_730,In_905);
or U258 (N_258,In_355,In_46);
nor U259 (N_259,In_328,In_513);
or U260 (N_260,In_431,In_819);
or U261 (N_261,In_879,In_235);
and U262 (N_262,In_678,In_597);
and U263 (N_263,In_354,In_784);
nand U264 (N_264,In_598,In_550);
and U265 (N_265,In_219,In_868);
nand U266 (N_266,In_901,In_78);
nand U267 (N_267,In_381,In_465);
nor U268 (N_268,In_677,In_188);
and U269 (N_269,In_832,In_520);
and U270 (N_270,In_805,In_294);
nand U271 (N_271,In_735,In_569);
nor U272 (N_272,In_20,In_125);
and U273 (N_273,In_252,In_614);
or U274 (N_274,In_752,In_179);
nand U275 (N_275,In_28,In_277);
or U276 (N_276,In_553,In_432);
xor U277 (N_277,In_746,In_380);
nor U278 (N_278,In_751,In_588);
nand U279 (N_279,In_545,In_142);
nand U280 (N_280,In_644,In_105);
nor U281 (N_281,In_494,In_845);
and U282 (N_282,In_12,In_273);
nor U283 (N_283,In_5,In_921);
xnor U284 (N_284,In_894,In_145);
or U285 (N_285,In_770,In_279);
nand U286 (N_286,In_430,In_225);
and U287 (N_287,In_326,In_508);
nand U288 (N_288,In_471,In_301);
nor U289 (N_289,In_19,In_757);
and U290 (N_290,In_304,In_882);
nor U291 (N_291,In_484,In_25);
and U292 (N_292,In_33,In_316);
and U293 (N_293,In_652,In_393);
and U294 (N_294,In_952,In_487);
and U295 (N_295,In_555,In_331);
or U296 (N_296,In_935,In_815);
and U297 (N_297,In_254,In_523);
nor U298 (N_298,In_463,In_197);
or U299 (N_299,In_32,In_22);
and U300 (N_300,In_593,In_611);
xnor U301 (N_301,In_676,In_434);
or U302 (N_302,In_970,In_942);
and U303 (N_303,In_153,In_93);
nor U304 (N_304,In_636,In_394);
xnor U305 (N_305,In_101,In_164);
nand U306 (N_306,In_583,In_856);
and U307 (N_307,In_540,In_621);
xnor U308 (N_308,In_486,In_680);
nand U309 (N_309,In_848,In_802);
xor U310 (N_310,In_556,In_173);
or U311 (N_311,In_41,In_283);
or U312 (N_312,In_497,In_425);
xor U313 (N_313,In_996,In_492);
and U314 (N_314,In_503,In_98);
or U315 (N_315,In_586,In_266);
xor U316 (N_316,In_167,In_324);
nor U317 (N_317,In_839,In_183);
or U318 (N_318,In_480,In_916);
nand U319 (N_319,In_236,In_956);
xor U320 (N_320,In_840,In_272);
and U321 (N_321,In_947,In_193);
nor U322 (N_322,In_312,In_674);
and U323 (N_323,In_862,In_202);
nand U324 (N_324,In_131,In_559);
nor U325 (N_325,In_400,In_81);
or U326 (N_326,In_170,In_127);
nor U327 (N_327,In_348,In_526);
nor U328 (N_328,In_516,In_231);
nor U329 (N_329,In_232,In_48);
xnor U330 (N_330,In_599,In_955);
or U331 (N_331,In_360,In_459);
nand U332 (N_332,In_97,In_303);
or U333 (N_333,In_452,In_831);
and U334 (N_334,In_289,In_194);
nand U335 (N_335,In_753,In_122);
or U336 (N_336,In_994,In_103);
nand U337 (N_337,In_657,In_633);
or U338 (N_338,In_811,In_124);
nand U339 (N_339,In_119,In_208);
nor U340 (N_340,In_507,In_936);
nor U341 (N_341,In_659,In_334);
nor U342 (N_342,In_960,In_779);
nor U343 (N_343,In_646,In_724);
nor U344 (N_344,In_923,In_410);
nand U345 (N_345,In_495,In_473);
xnor U346 (N_346,In_152,In_196);
or U347 (N_347,In_803,In_112);
nand U348 (N_348,In_458,In_248);
and U349 (N_349,In_201,In_281);
and U350 (N_350,In_479,In_977);
and U351 (N_351,In_989,In_466);
nor U352 (N_352,In_767,In_531);
nand U353 (N_353,In_506,In_745);
xor U354 (N_354,In_909,In_482);
and U355 (N_355,In_765,In_704);
or U356 (N_356,In_533,In_816);
or U357 (N_357,In_99,In_865);
and U358 (N_358,In_47,In_713);
nor U359 (N_359,In_496,In_626);
nor U360 (N_360,In_15,In_833);
nor U361 (N_361,In_813,In_161);
nor U362 (N_362,In_824,In_643);
nor U363 (N_363,In_775,In_732);
nand U364 (N_364,In_880,In_823);
and U365 (N_365,In_351,In_45);
and U366 (N_366,In_749,In_398);
or U367 (N_367,In_313,In_635);
and U368 (N_368,In_709,In_383);
and U369 (N_369,In_162,In_910);
and U370 (N_370,In_691,In_293);
nand U371 (N_371,In_852,In_841);
and U372 (N_372,In_222,In_863);
nor U373 (N_373,In_800,In_837);
and U374 (N_374,In_791,In_978);
or U375 (N_375,In_998,In_908);
nand U376 (N_376,In_849,In_850);
and U377 (N_377,In_787,In_689);
nor U378 (N_378,In_623,In_469);
nand U379 (N_379,In_773,In_651);
and U380 (N_380,In_549,In_370);
nand U381 (N_381,In_913,In_990);
nand U382 (N_382,In_914,In_209);
nor U383 (N_383,In_953,In_539);
and U384 (N_384,In_357,In_69);
and U385 (N_385,In_551,In_672);
nand U386 (N_386,In_439,In_584);
xnor U387 (N_387,In_7,In_333);
or U388 (N_388,In_607,In_720);
or U389 (N_389,In_859,In_511);
xnor U390 (N_390,In_510,In_17);
nor U391 (N_391,In_900,In_472);
nor U392 (N_392,In_238,In_308);
or U393 (N_393,In_983,In_117);
and U394 (N_394,In_932,In_35);
nor U395 (N_395,In_158,In_234);
nor U396 (N_396,In_102,In_275);
and U397 (N_397,In_185,In_378);
and U398 (N_398,In_984,In_675);
nand U399 (N_399,In_697,In_563);
and U400 (N_400,In_959,In_685);
or U401 (N_401,In_632,In_329);
nor U402 (N_402,In_177,In_884);
nor U403 (N_403,In_727,In_338);
and U404 (N_404,In_577,In_159);
and U405 (N_405,In_673,In_997);
or U406 (N_406,In_474,In_766);
or U407 (N_407,In_376,In_917);
xor U408 (N_408,In_552,In_337);
and U409 (N_409,In_924,In_149);
nor U410 (N_410,In_891,In_171);
and U411 (N_411,In_364,In_667);
nand U412 (N_412,In_642,In_718);
nand U413 (N_413,In_146,In_260);
nand U414 (N_414,In_591,In_464);
or U415 (N_415,In_307,In_895);
and U416 (N_416,In_696,In_211);
xnor U417 (N_417,In_505,In_818);
nand U418 (N_418,In_34,In_820);
nand U419 (N_419,In_288,In_343);
nand U420 (N_420,In_113,In_768);
or U421 (N_421,In_42,In_889);
xor U422 (N_422,In_189,In_278);
or U423 (N_423,In_560,In_769);
or U424 (N_424,In_634,In_546);
nor U425 (N_425,In_592,In_390);
or U426 (N_426,In_344,In_461);
nand U427 (N_427,In_137,In_240);
or U428 (N_428,In_403,In_133);
nor U429 (N_429,In_575,In_737);
or U430 (N_430,In_309,In_962);
nor U431 (N_431,In_554,In_772);
nor U432 (N_432,In_428,In_536);
and U433 (N_433,In_501,In_951);
nand U434 (N_434,In_258,In_110);
nand U435 (N_435,In_143,In_268);
nand U436 (N_436,In_302,In_684);
nor U437 (N_437,In_857,In_295);
nand U438 (N_438,In_904,In_918);
nor U439 (N_439,In_543,In_213);
and U440 (N_440,In_181,In_571);
nand U441 (N_441,In_377,In_538);
nor U442 (N_442,In_323,In_111);
and U443 (N_443,In_758,In_855);
nor U444 (N_444,In_706,In_292);
nand U445 (N_445,In_639,In_317);
and U446 (N_446,In_798,In_447);
or U447 (N_447,In_974,In_39);
and U448 (N_448,In_59,In_920);
xnor U449 (N_449,In_51,In_385);
nor U450 (N_450,In_77,In_925);
nand U451 (N_451,In_31,In_705);
and U452 (N_452,In_530,In_310);
nor U453 (N_453,In_992,In_129);
or U454 (N_454,In_502,In_694);
or U455 (N_455,In_165,In_890);
nand U456 (N_456,In_512,In_668);
xor U457 (N_457,In_417,In_866);
nor U458 (N_458,In_405,In_688);
xnor U459 (N_459,In_418,In_892);
or U460 (N_460,In_629,In_30);
nand U461 (N_461,In_406,In_898);
nand U462 (N_462,In_358,In_957);
nor U463 (N_463,In_796,In_107);
nand U464 (N_464,In_544,In_325);
nor U465 (N_465,In_147,In_703);
nor U466 (N_466,In_682,In_581);
or U467 (N_467,In_27,In_379);
and U468 (N_468,In_986,In_154);
and U469 (N_469,In_445,In_199);
xnor U470 (N_470,In_68,In_285);
nand U471 (N_471,In_139,In_84);
nand U472 (N_472,In_875,In_118);
nor U473 (N_473,In_327,In_37);
and U474 (N_474,In_483,In_851);
nor U475 (N_475,In_606,In_810);
nor U476 (N_476,In_912,In_363);
nand U477 (N_477,In_965,In_79);
or U478 (N_478,In_319,In_305);
and U479 (N_479,In_843,In_529);
nand U480 (N_480,In_314,In_903);
and U481 (N_481,In_186,In_134);
nor U482 (N_482,In_224,In_648);
xnor U483 (N_483,In_436,In_174);
xnor U484 (N_484,In_350,In_423);
or U485 (N_485,In_748,In_271);
and U486 (N_486,In_230,In_391);
and U487 (N_487,In_65,In_590);
nand U488 (N_488,In_253,In_433);
and U489 (N_489,In_771,In_488);
xnor U490 (N_490,In_71,In_515);
nand U491 (N_491,In_408,In_750);
nor U492 (N_492,In_991,In_226);
and U493 (N_493,In_527,In_548);
nor U494 (N_494,In_247,In_422);
or U495 (N_495,In_825,In_622);
or U496 (N_496,In_794,In_106);
nand U497 (N_497,In_108,In_742);
or U498 (N_498,In_126,In_444);
or U499 (N_499,In_52,In_470);
or U500 (N_500,In_411,In_642);
nand U501 (N_501,In_438,In_115);
or U502 (N_502,In_103,In_482);
and U503 (N_503,In_132,In_407);
or U504 (N_504,In_648,In_897);
nor U505 (N_505,In_47,In_286);
or U506 (N_506,In_659,In_540);
nor U507 (N_507,In_724,In_976);
nor U508 (N_508,In_295,In_793);
and U509 (N_509,In_943,In_283);
or U510 (N_510,In_912,In_756);
nand U511 (N_511,In_631,In_305);
nor U512 (N_512,In_581,In_133);
xor U513 (N_513,In_799,In_526);
nand U514 (N_514,In_316,In_879);
and U515 (N_515,In_554,In_6);
nor U516 (N_516,In_723,In_708);
and U517 (N_517,In_28,In_990);
nand U518 (N_518,In_543,In_246);
nand U519 (N_519,In_674,In_790);
and U520 (N_520,In_633,In_938);
and U521 (N_521,In_845,In_514);
or U522 (N_522,In_716,In_424);
or U523 (N_523,In_570,In_171);
and U524 (N_524,In_419,In_810);
or U525 (N_525,In_70,In_127);
and U526 (N_526,In_542,In_481);
nor U527 (N_527,In_444,In_681);
nand U528 (N_528,In_396,In_852);
xor U529 (N_529,In_780,In_641);
and U530 (N_530,In_76,In_619);
nand U531 (N_531,In_332,In_219);
nor U532 (N_532,In_161,In_719);
or U533 (N_533,In_524,In_576);
nand U534 (N_534,In_5,In_79);
nor U535 (N_535,In_515,In_339);
nand U536 (N_536,In_934,In_121);
nand U537 (N_537,In_84,In_347);
xor U538 (N_538,In_819,In_710);
and U539 (N_539,In_659,In_864);
and U540 (N_540,In_756,In_243);
nor U541 (N_541,In_416,In_374);
nand U542 (N_542,In_814,In_221);
xor U543 (N_543,In_980,In_422);
and U544 (N_544,In_770,In_998);
and U545 (N_545,In_338,In_527);
nand U546 (N_546,In_2,In_924);
nand U547 (N_547,In_429,In_788);
nand U548 (N_548,In_346,In_576);
xnor U549 (N_549,In_854,In_628);
nor U550 (N_550,In_431,In_364);
and U551 (N_551,In_919,In_887);
xnor U552 (N_552,In_442,In_516);
and U553 (N_553,In_127,In_928);
nand U554 (N_554,In_435,In_881);
nand U555 (N_555,In_353,In_247);
and U556 (N_556,In_806,In_191);
xor U557 (N_557,In_523,In_974);
or U558 (N_558,In_640,In_906);
nand U559 (N_559,In_807,In_111);
xor U560 (N_560,In_356,In_568);
nor U561 (N_561,In_534,In_988);
and U562 (N_562,In_231,In_502);
and U563 (N_563,In_286,In_910);
and U564 (N_564,In_597,In_92);
or U565 (N_565,In_709,In_952);
nand U566 (N_566,In_316,In_696);
or U567 (N_567,In_442,In_844);
or U568 (N_568,In_542,In_948);
xnor U569 (N_569,In_839,In_705);
or U570 (N_570,In_112,In_463);
and U571 (N_571,In_837,In_494);
or U572 (N_572,In_494,In_429);
or U573 (N_573,In_552,In_199);
xor U574 (N_574,In_952,In_394);
xor U575 (N_575,In_468,In_270);
and U576 (N_576,In_747,In_301);
and U577 (N_577,In_297,In_531);
or U578 (N_578,In_688,In_747);
nor U579 (N_579,In_356,In_259);
nand U580 (N_580,In_946,In_577);
and U581 (N_581,In_430,In_259);
xor U582 (N_582,In_253,In_502);
nor U583 (N_583,In_987,In_256);
or U584 (N_584,In_267,In_749);
nor U585 (N_585,In_883,In_158);
nand U586 (N_586,In_761,In_955);
or U587 (N_587,In_377,In_191);
and U588 (N_588,In_320,In_913);
nand U589 (N_589,In_219,In_211);
and U590 (N_590,In_875,In_241);
nor U591 (N_591,In_868,In_594);
or U592 (N_592,In_410,In_809);
and U593 (N_593,In_645,In_653);
nor U594 (N_594,In_817,In_77);
nand U595 (N_595,In_398,In_420);
or U596 (N_596,In_722,In_273);
and U597 (N_597,In_737,In_967);
nor U598 (N_598,In_650,In_595);
nand U599 (N_599,In_978,In_671);
or U600 (N_600,In_840,In_521);
or U601 (N_601,In_164,In_749);
and U602 (N_602,In_479,In_720);
xor U603 (N_603,In_628,In_622);
or U604 (N_604,In_649,In_465);
nand U605 (N_605,In_700,In_563);
xor U606 (N_606,In_446,In_415);
or U607 (N_607,In_770,In_683);
and U608 (N_608,In_810,In_74);
xor U609 (N_609,In_560,In_814);
nor U610 (N_610,In_587,In_487);
nand U611 (N_611,In_957,In_924);
nand U612 (N_612,In_173,In_706);
or U613 (N_613,In_759,In_685);
and U614 (N_614,In_804,In_92);
nand U615 (N_615,In_321,In_57);
nor U616 (N_616,In_83,In_872);
nor U617 (N_617,In_781,In_134);
nand U618 (N_618,In_481,In_350);
nor U619 (N_619,In_941,In_900);
and U620 (N_620,In_827,In_813);
and U621 (N_621,In_329,In_507);
nand U622 (N_622,In_148,In_565);
nand U623 (N_623,In_76,In_895);
and U624 (N_624,In_84,In_202);
nor U625 (N_625,In_143,In_769);
and U626 (N_626,In_168,In_502);
or U627 (N_627,In_742,In_976);
or U628 (N_628,In_773,In_902);
nor U629 (N_629,In_911,In_920);
xnor U630 (N_630,In_251,In_718);
nand U631 (N_631,In_670,In_663);
and U632 (N_632,In_236,In_731);
and U633 (N_633,In_883,In_670);
nor U634 (N_634,In_520,In_181);
xor U635 (N_635,In_248,In_833);
nor U636 (N_636,In_778,In_802);
nor U637 (N_637,In_641,In_81);
nor U638 (N_638,In_997,In_146);
nand U639 (N_639,In_812,In_433);
xnor U640 (N_640,In_945,In_492);
or U641 (N_641,In_469,In_748);
nand U642 (N_642,In_895,In_985);
nand U643 (N_643,In_512,In_398);
and U644 (N_644,In_295,In_468);
or U645 (N_645,In_24,In_562);
or U646 (N_646,In_543,In_390);
or U647 (N_647,In_457,In_166);
or U648 (N_648,In_980,In_707);
and U649 (N_649,In_528,In_472);
nand U650 (N_650,In_109,In_46);
and U651 (N_651,In_291,In_9);
nor U652 (N_652,In_272,In_470);
and U653 (N_653,In_186,In_699);
or U654 (N_654,In_733,In_61);
xnor U655 (N_655,In_116,In_692);
and U656 (N_656,In_749,In_184);
and U657 (N_657,In_966,In_305);
xnor U658 (N_658,In_191,In_477);
nand U659 (N_659,In_561,In_942);
nor U660 (N_660,In_818,In_543);
or U661 (N_661,In_65,In_556);
nor U662 (N_662,In_947,In_231);
xor U663 (N_663,In_694,In_561);
or U664 (N_664,In_672,In_510);
or U665 (N_665,In_586,In_478);
and U666 (N_666,In_933,In_451);
nand U667 (N_667,In_146,In_701);
and U668 (N_668,In_499,In_268);
nor U669 (N_669,In_285,In_963);
and U670 (N_670,In_577,In_490);
and U671 (N_671,In_128,In_487);
nand U672 (N_672,In_710,In_100);
nand U673 (N_673,In_658,In_474);
nor U674 (N_674,In_68,In_721);
xnor U675 (N_675,In_591,In_462);
nor U676 (N_676,In_323,In_552);
or U677 (N_677,In_296,In_235);
nand U678 (N_678,In_231,In_959);
nand U679 (N_679,In_818,In_145);
or U680 (N_680,In_159,In_983);
nor U681 (N_681,In_351,In_758);
and U682 (N_682,In_841,In_935);
xor U683 (N_683,In_453,In_841);
or U684 (N_684,In_986,In_54);
or U685 (N_685,In_382,In_75);
nand U686 (N_686,In_498,In_581);
nor U687 (N_687,In_622,In_875);
nand U688 (N_688,In_142,In_699);
or U689 (N_689,In_540,In_709);
or U690 (N_690,In_177,In_648);
or U691 (N_691,In_855,In_111);
and U692 (N_692,In_523,In_37);
and U693 (N_693,In_897,In_789);
nor U694 (N_694,In_801,In_831);
nor U695 (N_695,In_885,In_886);
or U696 (N_696,In_562,In_120);
and U697 (N_697,In_148,In_451);
nor U698 (N_698,In_242,In_549);
and U699 (N_699,In_557,In_39);
or U700 (N_700,In_577,In_336);
xor U701 (N_701,In_188,In_928);
nand U702 (N_702,In_476,In_973);
or U703 (N_703,In_559,In_488);
nand U704 (N_704,In_987,In_568);
xnor U705 (N_705,In_874,In_984);
or U706 (N_706,In_996,In_885);
or U707 (N_707,In_159,In_549);
nand U708 (N_708,In_305,In_357);
nand U709 (N_709,In_854,In_127);
or U710 (N_710,In_869,In_405);
and U711 (N_711,In_384,In_727);
nor U712 (N_712,In_430,In_174);
and U713 (N_713,In_464,In_318);
or U714 (N_714,In_588,In_282);
and U715 (N_715,In_747,In_506);
nor U716 (N_716,In_243,In_142);
and U717 (N_717,In_350,In_65);
nor U718 (N_718,In_258,In_249);
nor U719 (N_719,In_335,In_551);
and U720 (N_720,In_588,In_67);
nand U721 (N_721,In_644,In_82);
or U722 (N_722,In_401,In_252);
and U723 (N_723,In_309,In_954);
xor U724 (N_724,In_548,In_204);
nand U725 (N_725,In_928,In_238);
nor U726 (N_726,In_830,In_693);
nor U727 (N_727,In_223,In_688);
nor U728 (N_728,In_827,In_890);
nor U729 (N_729,In_495,In_973);
or U730 (N_730,In_46,In_527);
nor U731 (N_731,In_523,In_166);
nor U732 (N_732,In_838,In_882);
or U733 (N_733,In_273,In_70);
nor U734 (N_734,In_133,In_499);
nor U735 (N_735,In_275,In_33);
or U736 (N_736,In_391,In_521);
nand U737 (N_737,In_972,In_348);
nor U738 (N_738,In_575,In_489);
or U739 (N_739,In_936,In_176);
and U740 (N_740,In_331,In_645);
nor U741 (N_741,In_144,In_62);
or U742 (N_742,In_158,In_101);
or U743 (N_743,In_741,In_597);
nor U744 (N_744,In_501,In_238);
nor U745 (N_745,In_793,In_670);
xor U746 (N_746,In_756,In_35);
or U747 (N_747,In_986,In_915);
nand U748 (N_748,In_465,In_964);
or U749 (N_749,In_453,In_110);
nor U750 (N_750,In_238,In_239);
and U751 (N_751,In_988,In_859);
nand U752 (N_752,In_459,In_239);
nand U753 (N_753,In_382,In_168);
or U754 (N_754,In_750,In_281);
and U755 (N_755,In_322,In_819);
nand U756 (N_756,In_579,In_960);
nor U757 (N_757,In_168,In_341);
or U758 (N_758,In_280,In_135);
nor U759 (N_759,In_320,In_856);
nand U760 (N_760,In_912,In_354);
nand U761 (N_761,In_125,In_276);
nand U762 (N_762,In_23,In_956);
or U763 (N_763,In_371,In_38);
nand U764 (N_764,In_928,In_196);
or U765 (N_765,In_315,In_659);
nor U766 (N_766,In_369,In_447);
or U767 (N_767,In_833,In_171);
nand U768 (N_768,In_488,In_534);
xor U769 (N_769,In_936,In_906);
nand U770 (N_770,In_425,In_32);
nor U771 (N_771,In_277,In_804);
nor U772 (N_772,In_863,In_172);
nand U773 (N_773,In_15,In_168);
or U774 (N_774,In_274,In_658);
nand U775 (N_775,In_68,In_779);
or U776 (N_776,In_790,In_41);
xor U777 (N_777,In_176,In_726);
nor U778 (N_778,In_173,In_309);
nand U779 (N_779,In_736,In_731);
or U780 (N_780,In_893,In_199);
nor U781 (N_781,In_215,In_273);
nor U782 (N_782,In_763,In_901);
or U783 (N_783,In_493,In_813);
and U784 (N_784,In_992,In_878);
and U785 (N_785,In_353,In_82);
xor U786 (N_786,In_775,In_912);
nor U787 (N_787,In_925,In_705);
nand U788 (N_788,In_8,In_144);
and U789 (N_789,In_288,In_743);
and U790 (N_790,In_789,In_445);
and U791 (N_791,In_959,In_936);
nor U792 (N_792,In_930,In_211);
nand U793 (N_793,In_936,In_764);
and U794 (N_794,In_716,In_616);
and U795 (N_795,In_345,In_488);
nor U796 (N_796,In_801,In_167);
nand U797 (N_797,In_241,In_568);
and U798 (N_798,In_320,In_379);
nand U799 (N_799,In_280,In_158);
nor U800 (N_800,In_135,In_878);
nor U801 (N_801,In_962,In_333);
or U802 (N_802,In_240,In_711);
nand U803 (N_803,In_474,In_767);
and U804 (N_804,In_224,In_44);
nor U805 (N_805,In_895,In_296);
nor U806 (N_806,In_389,In_317);
nor U807 (N_807,In_256,In_227);
xnor U808 (N_808,In_707,In_123);
nand U809 (N_809,In_48,In_394);
or U810 (N_810,In_67,In_164);
nor U811 (N_811,In_748,In_875);
and U812 (N_812,In_408,In_336);
nand U813 (N_813,In_636,In_752);
nor U814 (N_814,In_569,In_172);
nand U815 (N_815,In_363,In_67);
nor U816 (N_816,In_429,In_64);
nand U817 (N_817,In_331,In_532);
nor U818 (N_818,In_199,In_219);
and U819 (N_819,In_237,In_205);
nand U820 (N_820,In_507,In_77);
and U821 (N_821,In_377,In_481);
nand U822 (N_822,In_972,In_279);
or U823 (N_823,In_667,In_840);
or U824 (N_824,In_607,In_742);
or U825 (N_825,In_404,In_177);
or U826 (N_826,In_417,In_82);
and U827 (N_827,In_165,In_120);
nand U828 (N_828,In_885,In_612);
nand U829 (N_829,In_332,In_148);
nor U830 (N_830,In_342,In_219);
and U831 (N_831,In_631,In_827);
nor U832 (N_832,In_486,In_66);
nor U833 (N_833,In_147,In_755);
nor U834 (N_834,In_966,In_85);
and U835 (N_835,In_896,In_316);
nand U836 (N_836,In_846,In_477);
nor U837 (N_837,In_424,In_940);
nand U838 (N_838,In_22,In_604);
and U839 (N_839,In_956,In_671);
or U840 (N_840,In_781,In_306);
nor U841 (N_841,In_111,In_40);
nand U842 (N_842,In_238,In_233);
nand U843 (N_843,In_624,In_662);
and U844 (N_844,In_272,In_435);
nor U845 (N_845,In_362,In_671);
nand U846 (N_846,In_388,In_951);
xor U847 (N_847,In_313,In_451);
or U848 (N_848,In_393,In_677);
nand U849 (N_849,In_454,In_466);
or U850 (N_850,In_651,In_631);
or U851 (N_851,In_157,In_924);
nand U852 (N_852,In_917,In_477);
or U853 (N_853,In_879,In_145);
nor U854 (N_854,In_578,In_186);
nand U855 (N_855,In_506,In_640);
xor U856 (N_856,In_768,In_172);
or U857 (N_857,In_10,In_247);
xor U858 (N_858,In_870,In_764);
and U859 (N_859,In_20,In_994);
nor U860 (N_860,In_937,In_795);
or U861 (N_861,In_699,In_436);
nand U862 (N_862,In_690,In_414);
xor U863 (N_863,In_203,In_915);
or U864 (N_864,In_730,In_95);
or U865 (N_865,In_851,In_659);
nand U866 (N_866,In_190,In_888);
nand U867 (N_867,In_589,In_796);
or U868 (N_868,In_761,In_573);
and U869 (N_869,In_994,In_593);
and U870 (N_870,In_481,In_968);
nor U871 (N_871,In_927,In_249);
xnor U872 (N_872,In_676,In_409);
nor U873 (N_873,In_718,In_135);
or U874 (N_874,In_42,In_759);
nand U875 (N_875,In_728,In_723);
nand U876 (N_876,In_46,In_100);
and U877 (N_877,In_272,In_93);
nand U878 (N_878,In_616,In_204);
nor U879 (N_879,In_774,In_776);
and U880 (N_880,In_300,In_430);
xor U881 (N_881,In_766,In_311);
nor U882 (N_882,In_721,In_737);
nor U883 (N_883,In_349,In_444);
or U884 (N_884,In_919,In_443);
nor U885 (N_885,In_709,In_934);
nor U886 (N_886,In_766,In_486);
and U887 (N_887,In_188,In_997);
nand U888 (N_888,In_700,In_930);
and U889 (N_889,In_102,In_825);
nor U890 (N_890,In_497,In_339);
and U891 (N_891,In_42,In_437);
xor U892 (N_892,In_561,In_473);
nor U893 (N_893,In_710,In_341);
or U894 (N_894,In_399,In_403);
and U895 (N_895,In_43,In_805);
xnor U896 (N_896,In_908,In_645);
xnor U897 (N_897,In_570,In_105);
nand U898 (N_898,In_570,In_520);
or U899 (N_899,In_345,In_853);
and U900 (N_900,In_235,In_250);
and U901 (N_901,In_604,In_379);
and U902 (N_902,In_92,In_188);
or U903 (N_903,In_383,In_864);
nand U904 (N_904,In_352,In_856);
nand U905 (N_905,In_239,In_484);
and U906 (N_906,In_388,In_315);
or U907 (N_907,In_378,In_352);
nand U908 (N_908,In_687,In_69);
nand U909 (N_909,In_368,In_849);
nor U910 (N_910,In_951,In_950);
or U911 (N_911,In_720,In_586);
nor U912 (N_912,In_535,In_669);
nand U913 (N_913,In_159,In_195);
or U914 (N_914,In_533,In_729);
and U915 (N_915,In_54,In_522);
or U916 (N_916,In_492,In_518);
or U917 (N_917,In_338,In_30);
nand U918 (N_918,In_924,In_488);
nor U919 (N_919,In_820,In_644);
nor U920 (N_920,In_724,In_375);
or U921 (N_921,In_34,In_997);
xnor U922 (N_922,In_313,In_398);
and U923 (N_923,In_84,In_789);
or U924 (N_924,In_561,In_322);
xor U925 (N_925,In_770,In_927);
nor U926 (N_926,In_279,In_529);
and U927 (N_927,In_854,In_118);
nor U928 (N_928,In_917,In_530);
xor U929 (N_929,In_462,In_485);
nand U930 (N_930,In_33,In_926);
nor U931 (N_931,In_593,In_524);
nand U932 (N_932,In_769,In_274);
nand U933 (N_933,In_337,In_455);
or U934 (N_934,In_887,In_251);
xnor U935 (N_935,In_478,In_724);
xor U936 (N_936,In_970,In_242);
and U937 (N_937,In_970,In_914);
nand U938 (N_938,In_259,In_555);
and U939 (N_939,In_403,In_153);
and U940 (N_940,In_675,In_468);
nor U941 (N_941,In_963,In_238);
nor U942 (N_942,In_682,In_826);
or U943 (N_943,In_49,In_650);
xnor U944 (N_944,In_351,In_882);
nand U945 (N_945,In_567,In_803);
nand U946 (N_946,In_519,In_72);
or U947 (N_947,In_874,In_761);
and U948 (N_948,In_533,In_427);
or U949 (N_949,In_189,In_100);
nand U950 (N_950,In_380,In_609);
nand U951 (N_951,In_20,In_840);
nor U952 (N_952,In_584,In_985);
and U953 (N_953,In_371,In_325);
nand U954 (N_954,In_208,In_345);
and U955 (N_955,In_372,In_52);
nand U956 (N_956,In_736,In_664);
nand U957 (N_957,In_145,In_677);
xnor U958 (N_958,In_86,In_132);
nor U959 (N_959,In_311,In_888);
nor U960 (N_960,In_667,In_809);
xor U961 (N_961,In_827,In_975);
nand U962 (N_962,In_480,In_227);
nor U963 (N_963,In_498,In_460);
nand U964 (N_964,In_533,In_596);
nor U965 (N_965,In_546,In_117);
or U966 (N_966,In_166,In_305);
nand U967 (N_967,In_537,In_656);
or U968 (N_968,In_982,In_49);
nor U969 (N_969,In_593,In_529);
or U970 (N_970,In_50,In_798);
nor U971 (N_971,In_797,In_30);
xnor U972 (N_972,In_895,In_125);
and U973 (N_973,In_212,In_269);
nand U974 (N_974,In_330,In_149);
or U975 (N_975,In_114,In_298);
or U976 (N_976,In_822,In_72);
xor U977 (N_977,In_223,In_844);
and U978 (N_978,In_982,In_11);
and U979 (N_979,In_849,In_907);
nand U980 (N_980,In_226,In_386);
nor U981 (N_981,In_433,In_466);
nor U982 (N_982,In_790,In_917);
or U983 (N_983,In_67,In_842);
and U984 (N_984,In_0,In_477);
or U985 (N_985,In_287,In_807);
nand U986 (N_986,In_940,In_439);
nor U987 (N_987,In_40,In_139);
or U988 (N_988,In_288,In_275);
and U989 (N_989,In_721,In_23);
and U990 (N_990,In_472,In_91);
or U991 (N_991,In_771,In_282);
xor U992 (N_992,In_873,In_350);
and U993 (N_993,In_558,In_145);
nand U994 (N_994,In_377,In_929);
nor U995 (N_995,In_745,In_43);
or U996 (N_996,In_750,In_494);
nand U997 (N_997,In_357,In_395);
and U998 (N_998,In_435,In_562);
nor U999 (N_999,In_789,In_590);
nor U1000 (N_1000,N_701,N_230);
nand U1001 (N_1001,N_780,N_914);
nand U1002 (N_1002,N_948,N_294);
nand U1003 (N_1003,N_631,N_165);
nand U1004 (N_1004,N_476,N_343);
nand U1005 (N_1005,N_710,N_619);
and U1006 (N_1006,N_10,N_439);
or U1007 (N_1007,N_273,N_980);
nand U1008 (N_1008,N_496,N_953);
nand U1009 (N_1009,N_829,N_920);
nand U1010 (N_1010,N_360,N_212);
and U1011 (N_1011,N_451,N_804);
or U1012 (N_1012,N_909,N_383);
or U1013 (N_1013,N_21,N_602);
nor U1014 (N_1014,N_70,N_595);
and U1015 (N_1015,N_785,N_364);
and U1016 (N_1016,N_621,N_510);
or U1017 (N_1017,N_659,N_239);
and U1018 (N_1018,N_961,N_340);
nor U1019 (N_1019,N_292,N_579);
or U1020 (N_1020,N_247,N_818);
nand U1021 (N_1021,N_404,N_492);
nor U1022 (N_1022,N_306,N_23);
nand U1023 (N_1023,N_204,N_880);
nand U1024 (N_1024,N_994,N_288);
or U1025 (N_1025,N_267,N_97);
xnor U1026 (N_1026,N_215,N_935);
nand U1027 (N_1027,N_145,N_666);
nand U1028 (N_1028,N_128,N_169);
nor U1029 (N_1029,N_740,N_896);
nand U1030 (N_1030,N_946,N_125);
nand U1031 (N_1031,N_535,N_851);
and U1032 (N_1032,N_121,N_782);
xor U1033 (N_1033,N_558,N_521);
nor U1034 (N_1034,N_585,N_205);
or U1035 (N_1035,N_14,N_49);
nand U1036 (N_1036,N_362,N_466);
xnor U1037 (N_1037,N_922,N_51);
and U1038 (N_1038,N_485,N_684);
and U1039 (N_1039,N_155,N_40);
or U1040 (N_1040,N_99,N_741);
or U1041 (N_1041,N_412,N_794);
or U1042 (N_1042,N_130,N_675);
nand U1043 (N_1043,N_414,N_736);
or U1044 (N_1044,N_458,N_94);
and U1045 (N_1045,N_256,N_930);
and U1046 (N_1046,N_877,N_136);
and U1047 (N_1047,N_416,N_725);
nor U1048 (N_1048,N_559,N_885);
or U1049 (N_1049,N_777,N_583);
nand U1050 (N_1050,N_609,N_366);
and U1051 (N_1051,N_652,N_942);
nand U1052 (N_1052,N_223,N_275);
nand U1053 (N_1053,N_76,N_891);
nand U1054 (N_1054,N_398,N_623);
and U1055 (N_1055,N_539,N_351);
and U1056 (N_1056,N_95,N_866);
or U1057 (N_1057,N_194,N_798);
nand U1058 (N_1058,N_327,N_810);
or U1059 (N_1059,N_557,N_981);
nor U1060 (N_1060,N_937,N_706);
nand U1061 (N_1061,N_775,N_724);
nand U1062 (N_1062,N_816,N_435);
nand U1063 (N_1063,N_511,N_24);
nand U1064 (N_1064,N_887,N_839);
or U1065 (N_1065,N_831,N_111);
nand U1066 (N_1066,N_897,N_6);
and U1067 (N_1067,N_620,N_911);
or U1068 (N_1068,N_770,N_312);
xnor U1069 (N_1069,N_187,N_386);
nand U1070 (N_1070,N_960,N_175);
nor U1071 (N_1071,N_949,N_957);
nor U1072 (N_1072,N_367,N_170);
nand U1073 (N_1073,N_532,N_389);
nor U1074 (N_1074,N_803,N_952);
or U1075 (N_1075,N_923,N_191);
nand U1076 (N_1076,N_749,N_462);
nor U1077 (N_1077,N_148,N_436);
and U1078 (N_1078,N_913,N_682);
or U1079 (N_1079,N_235,N_625);
and U1080 (N_1080,N_931,N_464);
or U1081 (N_1081,N_184,N_192);
nor U1082 (N_1082,N_475,N_197);
nor U1083 (N_1083,N_255,N_159);
and U1084 (N_1084,N_743,N_497);
xnor U1085 (N_1085,N_124,N_453);
nor U1086 (N_1086,N_153,N_939);
or U1087 (N_1087,N_938,N_80);
nand U1088 (N_1088,N_392,N_632);
or U1089 (N_1089,N_728,N_556);
nor U1090 (N_1090,N_189,N_567);
or U1091 (N_1091,N_339,N_468);
nand U1092 (N_1092,N_713,N_237);
nor U1093 (N_1093,N_448,N_699);
nor U1094 (N_1094,N_719,N_457);
or U1095 (N_1095,N_31,N_59);
nand U1096 (N_1096,N_742,N_424);
nand U1097 (N_1097,N_917,N_940);
xnor U1098 (N_1098,N_797,N_307);
or U1099 (N_1099,N_924,N_830);
xnor U1100 (N_1100,N_562,N_86);
or U1101 (N_1101,N_951,N_657);
xnor U1102 (N_1102,N_899,N_36);
nor U1103 (N_1103,N_745,N_397);
or U1104 (N_1104,N_598,N_519);
and U1105 (N_1105,N_926,N_3);
and U1106 (N_1106,N_119,N_310);
nor U1107 (N_1107,N_872,N_808);
xnor U1108 (N_1108,N_102,N_615);
nand U1109 (N_1109,N_57,N_517);
nand U1110 (N_1110,N_892,N_863);
and U1111 (N_1111,N_206,N_857);
or U1112 (N_1112,N_847,N_495);
nor U1113 (N_1113,N_591,N_918);
xor U1114 (N_1114,N_336,N_429);
nor U1115 (N_1115,N_744,N_382);
nand U1116 (N_1116,N_201,N_802);
nand U1117 (N_1117,N_42,N_793);
nor U1118 (N_1118,N_18,N_972);
nor U1119 (N_1119,N_482,N_131);
nor U1120 (N_1120,N_748,N_985);
nor U1121 (N_1121,N_779,N_586);
nand U1122 (N_1122,N_478,N_754);
nand U1123 (N_1123,N_947,N_842);
nor U1124 (N_1124,N_238,N_305);
xor U1125 (N_1125,N_322,N_762);
or U1126 (N_1126,N_614,N_552);
nor U1127 (N_1127,N_297,N_873);
and U1128 (N_1128,N_37,N_442);
nand U1129 (N_1129,N_489,N_444);
or U1130 (N_1130,N_520,N_893);
nor U1131 (N_1131,N_443,N_222);
nor U1132 (N_1132,N_551,N_253);
and U1133 (N_1133,N_231,N_582);
nor U1134 (N_1134,N_164,N_574);
xnor U1135 (N_1135,N_848,N_450);
nor U1136 (N_1136,N_229,N_859);
nor U1137 (N_1137,N_565,N_499);
nor U1138 (N_1138,N_525,N_261);
nor U1139 (N_1139,N_642,N_648);
xnor U1140 (N_1140,N_507,N_549);
and U1141 (N_1141,N_195,N_162);
or U1142 (N_1142,N_796,N_638);
nor U1143 (N_1143,N_167,N_67);
or U1144 (N_1144,N_705,N_157);
nand U1145 (N_1145,N_19,N_954);
and U1146 (N_1146,N_732,N_72);
nand U1147 (N_1147,N_225,N_266);
xor U1148 (N_1148,N_203,N_393);
or U1149 (N_1149,N_168,N_597);
nand U1150 (N_1150,N_143,N_245);
and U1151 (N_1151,N_656,N_426);
or U1152 (N_1152,N_965,N_427);
and U1153 (N_1153,N_672,N_932);
nand U1154 (N_1154,N_140,N_811);
and U1155 (N_1155,N_304,N_64);
nor U1156 (N_1156,N_228,N_678);
nand U1157 (N_1157,N_976,N_88);
or U1158 (N_1158,N_950,N_871);
nand U1159 (N_1159,N_771,N_359);
nor U1160 (N_1160,N_856,N_285);
nor U1161 (N_1161,N_193,N_141);
nor U1162 (N_1162,N_760,N_372);
or U1163 (N_1163,N_934,N_303);
and U1164 (N_1164,N_368,N_828);
nor U1165 (N_1165,N_555,N_680);
or U1166 (N_1166,N_628,N_983);
nor U1167 (N_1167,N_577,N_5);
or U1168 (N_1168,N_433,N_461);
nand U1169 (N_1169,N_884,N_469);
and U1170 (N_1170,N_211,N_467);
nand U1171 (N_1171,N_272,N_606);
xnor U1172 (N_1172,N_258,N_216);
or U1173 (N_1173,N_68,N_110);
nand U1174 (N_1174,N_737,N_773);
nand U1175 (N_1175,N_116,N_480);
or U1176 (N_1176,N_487,N_459);
and U1177 (N_1177,N_969,N_408);
xnor U1178 (N_1178,N_115,N_146);
xnor U1179 (N_1179,N_694,N_751);
nand U1180 (N_1180,N_276,N_217);
nand U1181 (N_1181,N_731,N_271);
and U1182 (N_1182,N_721,N_455);
nand U1183 (N_1183,N_346,N_668);
xnor U1184 (N_1184,N_895,N_317);
and U1185 (N_1185,N_208,N_463);
or U1186 (N_1186,N_149,N_575);
and U1187 (N_1187,N_844,N_415);
nand U1188 (N_1188,N_66,N_755);
and U1189 (N_1189,N_975,N_686);
or U1190 (N_1190,N_270,N_542);
nand U1191 (N_1191,N_837,N_257);
and U1192 (N_1192,N_83,N_827);
nor U1193 (N_1193,N_333,N_547);
and U1194 (N_1194,N_612,N_502);
and U1195 (N_1195,N_423,N_38);
and U1196 (N_1196,N_908,N_987);
and U1197 (N_1197,N_881,N_815);
nand U1198 (N_1198,N_279,N_323);
or U1199 (N_1199,N_113,N_945);
or U1200 (N_1200,N_864,N_784);
and U1201 (N_1201,N_4,N_207);
and U1202 (N_1202,N_405,N_471);
nor U1203 (N_1203,N_63,N_377);
xor U1204 (N_1204,N_107,N_243);
or U1205 (N_1205,N_479,N_603);
nor U1206 (N_1206,N_409,N_27);
nor U1207 (N_1207,N_387,N_826);
or U1208 (N_1208,N_910,N_993);
nor U1209 (N_1209,N_792,N_825);
nand U1210 (N_1210,N_630,N_548);
nor U1211 (N_1211,N_654,N_852);
nor U1212 (N_1212,N_500,N_538);
or U1213 (N_1213,N_202,N_353);
nor U1214 (N_1214,N_596,N_388);
nor U1215 (N_1215,N_580,N_966);
nor U1216 (N_1216,N_639,N_308);
xnor U1217 (N_1217,N_707,N_379);
and U1218 (N_1218,N_447,N_540);
or U1219 (N_1219,N_61,N_139);
or U1220 (N_1220,N_399,N_999);
or U1221 (N_1221,N_89,N_26);
xnor U1222 (N_1222,N_287,N_209);
nor U1223 (N_1223,N_677,N_268);
and U1224 (N_1224,N_514,N_841);
nand U1225 (N_1225,N_233,N_868);
nand U1226 (N_1226,N_144,N_190);
nor U1227 (N_1227,N_365,N_901);
or U1228 (N_1228,N_753,N_299);
and U1229 (N_1229,N_325,N_309);
xor U1230 (N_1230,N_440,N_823);
nand U1231 (N_1231,N_791,N_992);
nor U1232 (N_1232,N_867,N_902);
xnor U1233 (N_1233,N_905,N_927);
or U1234 (N_1234,N_33,N_356);
nand U1235 (N_1235,N_79,N_958);
or U1236 (N_1236,N_154,N_262);
or U1237 (N_1237,N_996,N_236);
xnor U1238 (N_1238,N_60,N_401);
xnor U1239 (N_1239,N_198,N_363);
xnor U1240 (N_1240,N_284,N_522);
nand U1241 (N_1241,N_681,N_93);
and U1242 (N_1242,N_104,N_173);
nor U1243 (N_1243,N_759,N_85);
or U1244 (N_1244,N_127,N_296);
or U1245 (N_1245,N_508,N_278);
nand U1246 (N_1246,N_7,N_509);
and U1247 (N_1247,N_894,N_550);
or U1248 (N_1248,N_670,N_177);
nand U1249 (N_1249,N_814,N_313);
or U1250 (N_1250,N_150,N_71);
or U1251 (N_1251,N_69,N_103);
and U1252 (N_1252,N_528,N_730);
nor U1253 (N_1253,N_766,N_413);
or U1254 (N_1254,N_50,N_286);
or U1255 (N_1255,N_249,N_536);
or U1256 (N_1256,N_347,N_955);
nor U1257 (N_1257,N_75,N_788);
xor U1258 (N_1258,N_20,N_530);
xnor U1259 (N_1259,N_274,N_460);
xor U1260 (N_1260,N_15,N_977);
and U1261 (N_1261,N_778,N_676);
xor U1262 (N_1262,N_219,N_32);
nor U1263 (N_1263,N_795,N_456);
nand U1264 (N_1264,N_515,N_758);
xor U1265 (N_1265,N_358,N_490);
and U1266 (N_1266,N_703,N_991);
xor U1267 (N_1267,N_526,N_473);
nor U1268 (N_1268,N_915,N_962);
and U1269 (N_1269,N_665,N_137);
xor U1270 (N_1270,N_645,N_700);
or U1271 (N_1271,N_156,N_772);
nand U1272 (N_1272,N_318,N_348);
nor U1273 (N_1273,N_371,N_428);
nand U1274 (N_1274,N_878,N_335);
and U1275 (N_1275,N_717,N_739);
nor U1276 (N_1276,N_504,N_834);
nor U1277 (N_1277,N_430,N_820);
nor U1278 (N_1278,N_722,N_662);
nand U1279 (N_1279,N_432,N_316);
or U1280 (N_1280,N_481,N_13);
or U1281 (N_1281,N_990,N_17);
or U1282 (N_1282,N_45,N_250);
or U1283 (N_1283,N_344,N_929);
and U1284 (N_1284,N_324,N_311);
and U1285 (N_1285,N_874,N_576);
and U1286 (N_1286,N_98,N_352);
nand U1287 (N_1287,N_840,N_617);
nor U1288 (N_1288,N_338,N_232);
nor U1289 (N_1289,N_767,N_384);
or U1290 (N_1290,N_587,N_817);
xnor U1291 (N_1291,N_112,N_369);
nand U1292 (N_1292,N_373,N_964);
and U1293 (N_1293,N_84,N_410);
nand U1294 (N_1294,N_805,N_315);
or U1295 (N_1295,N_634,N_769);
nor U1296 (N_1296,N_968,N_2);
nand U1297 (N_1297,N_166,N_858);
or U1298 (N_1298,N_698,N_936);
nand U1299 (N_1299,N_246,N_210);
nand U1300 (N_1300,N_445,N_752);
and U1301 (N_1301,N_252,N_746);
nor U1302 (N_1302,N_807,N_761);
nand U1303 (N_1303,N_763,N_970);
or U1304 (N_1304,N_643,N_692);
xnor U1305 (N_1305,N_875,N_855);
or U1306 (N_1306,N_337,N_669);
or U1307 (N_1307,N_251,N_180);
and U1308 (N_1308,N_16,N_685);
nor U1309 (N_1309,N_293,N_503);
nand U1310 (N_1310,N_849,N_123);
and U1311 (N_1311,N_378,N_738);
or U1312 (N_1312,N_610,N_158);
nand U1313 (N_1313,N_400,N_571);
or U1314 (N_1314,N_101,N_330);
nor U1315 (N_1315,N_683,N_394);
xnor U1316 (N_1316,N_854,N_697);
and U1317 (N_1317,N_133,N_53);
and U1318 (N_1318,N_860,N_30);
nor U1319 (N_1319,N_882,N_513);
or U1320 (N_1320,N_693,N_454);
or U1321 (N_1321,N_709,N_501);
nor U1322 (N_1322,N_269,N_819);
nand U1323 (N_1323,N_906,N_302);
nor U1324 (N_1324,N_765,N_789);
and U1325 (N_1325,N_824,N_712);
xor U1326 (N_1326,N_786,N_474);
or U1327 (N_1327,N_90,N_39);
xnor U1328 (N_1328,N_512,N_385);
nor U1329 (N_1329,N_374,N_114);
xor U1330 (N_1330,N_812,N_100);
or U1331 (N_1331,N_376,N_543);
nand U1332 (N_1332,N_117,N_518);
nand U1333 (N_1333,N_56,N_91);
xor U1334 (N_1334,N_822,N_890);
nor U1335 (N_1335,N_733,N_281);
nand U1336 (N_1336,N_853,N_653);
nand U1337 (N_1337,N_47,N_605);
and U1338 (N_1338,N_221,N_544);
nand U1339 (N_1339,N_919,N_613);
nand U1340 (N_1340,N_626,N_241);
nor U1341 (N_1341,N_572,N_437);
nor U1342 (N_1342,N_264,N_527);
and U1343 (N_1343,N_58,N_298);
nand U1344 (N_1344,N_29,N_718);
nor U1345 (N_1345,N_182,N_265);
or U1346 (N_1346,N_226,N_646);
nor U1347 (N_1347,N_644,N_488);
nor U1348 (N_1348,N_498,N_341);
nor U1349 (N_1349,N_912,N_879);
and U1350 (N_1350,N_688,N_46);
xor U1351 (N_1351,N_702,N_865);
or U1352 (N_1352,N_664,N_118);
nand U1353 (N_1353,N_869,N_838);
nor U1354 (N_1354,N_34,N_982);
nor U1355 (N_1355,N_406,N_928);
xor U1356 (N_1356,N_714,N_781);
or U1357 (N_1357,N_986,N_77);
and U1358 (N_1358,N_870,N_592);
or U1359 (N_1359,N_647,N_650);
nand U1360 (N_1360,N_402,N_581);
nand U1361 (N_1361,N_845,N_199);
xor U1362 (N_1362,N_846,N_533);
nand U1363 (N_1363,N_534,N_81);
nand U1364 (N_1364,N_998,N_354);
nor U1365 (N_1365,N_244,N_438);
nor U1366 (N_1366,N_799,N_196);
nand U1367 (N_1367,N_301,N_833);
xnor U1368 (N_1368,N_505,N_641);
or U1369 (N_1369,N_135,N_801);
nor U1370 (N_1370,N_989,N_573);
nor U1371 (N_1371,N_390,N_523);
nor U1372 (N_1372,N_350,N_974);
nand U1373 (N_1373,N_661,N_78);
nor U1374 (N_1374,N_898,N_734);
xnor U1375 (N_1375,N_959,N_28);
and U1376 (N_1376,N_283,N_48);
or U1377 (N_1377,N_524,N_419);
nor U1378 (N_1378,N_944,N_422);
nand U1379 (N_1379,N_564,N_396);
nand U1380 (N_1380,N_560,N_151);
nand U1381 (N_1381,N_1,N_941);
nand U1382 (N_1382,N_674,N_254);
or U1383 (N_1383,N_493,N_978);
nand U1384 (N_1384,N_622,N_291);
or U1385 (N_1385,N_821,N_345);
and U1386 (N_1386,N_616,N_420);
nand U1387 (N_1387,N_431,N_349);
nor U1388 (N_1388,N_715,N_806);
and U1389 (N_1389,N_174,N_783);
and U1390 (N_1390,N_618,N_9);
or U1391 (N_1391,N_134,N_843);
or U1392 (N_1392,N_636,N_608);
nand U1393 (N_1393,N_716,N_43);
nor U1394 (N_1394,N_142,N_470);
or U1395 (N_1395,N_220,N_326);
and U1396 (N_1396,N_234,N_465);
nor U1397 (N_1397,N_750,N_494);
nor U1398 (N_1398,N_321,N_65);
nand U1399 (N_1399,N_590,N_280);
nand U1400 (N_1400,N_188,N_679);
nand U1401 (N_1401,N_629,N_263);
nor U1402 (N_1402,N_183,N_375);
or U1403 (N_1403,N_704,N_214);
and U1404 (N_1404,N_607,N_54);
nand U1405 (N_1405,N_747,N_129);
and U1406 (N_1406,N_649,N_132);
and U1407 (N_1407,N_655,N_836);
and U1408 (N_1408,N_178,N_355);
nand U1409 (N_1409,N_570,N_813);
nand U1410 (N_1410,N_282,N_850);
nand U1411 (N_1411,N_667,N_411);
and U1412 (N_1412,N_635,N_599);
nor U1413 (N_1413,N_147,N_391);
or U1414 (N_1414,N_35,N_963);
nand U1415 (N_1415,N_691,N_441);
and U1416 (N_1416,N_900,N_764);
or U1417 (N_1417,N_988,N_888);
nor U1418 (N_1418,N_862,N_483);
nor U1419 (N_1419,N_171,N_593);
and U1420 (N_1420,N_624,N_248);
nand U1421 (N_1421,N_651,N_861);
or U1422 (N_1422,N_589,N_627);
or U1423 (N_1423,N_96,N_105);
xor U1424 (N_1424,N_477,N_907);
nand U1425 (N_1425,N_213,N_290);
nor U1426 (N_1426,N_452,N_109);
xor U1427 (N_1427,N_711,N_44);
and U1428 (N_1428,N_395,N_726);
and U1429 (N_1429,N_240,N_163);
or U1430 (N_1430,N_545,N_588);
nor U1431 (N_1431,N_277,N_637);
nor U1432 (N_1432,N_916,N_876);
nand U1433 (N_1433,N_832,N_563);
and U1434 (N_1434,N_92,N_809);
nor U1435 (N_1435,N_708,N_152);
or U1436 (N_1436,N_995,N_126);
nor U1437 (N_1437,N_600,N_361);
nor U1438 (N_1438,N_224,N_611);
nand U1439 (N_1439,N_800,N_529);
or U1440 (N_1440,N_295,N_835);
nand U1441 (N_1441,N_673,N_578);
and U1442 (N_1442,N_74,N_314);
xor U1443 (N_1443,N_242,N_889);
xor U1444 (N_1444,N_55,N_484);
xnor U1445 (N_1445,N_200,N_735);
xor U1446 (N_1446,N_179,N_122);
and U1447 (N_1447,N_62,N_903);
xor U1448 (N_1448,N_106,N_289);
nand U1449 (N_1449,N_604,N_160);
and U1450 (N_1450,N_449,N_138);
nor U1451 (N_1451,N_120,N_569);
or U1452 (N_1452,N_633,N_331);
and U1453 (N_1453,N_328,N_554);
xnor U1454 (N_1454,N_421,N_260);
and U1455 (N_1455,N_566,N_12);
nor U1456 (N_1456,N_407,N_768);
or U1457 (N_1457,N_594,N_660);
nor U1458 (N_1458,N_52,N_486);
or U1459 (N_1459,N_108,N_546);
and U1460 (N_1460,N_921,N_663);
nor U1461 (N_1461,N_756,N_185);
and U1462 (N_1462,N_434,N_687);
xor U1463 (N_1463,N_329,N_601);
nand U1464 (N_1464,N_227,N_997);
and U1465 (N_1465,N_541,N_774);
nor U1466 (N_1466,N_357,N_658);
and U1467 (N_1467,N_640,N_506);
and U1468 (N_1468,N_787,N_973);
nand U1469 (N_1469,N_933,N_790);
xor U1470 (N_1470,N_181,N_380);
nand U1471 (N_1471,N_417,N_883);
or U1472 (N_1472,N_568,N_332);
nor U1473 (N_1473,N_979,N_690);
or U1474 (N_1474,N_729,N_320);
nor U1475 (N_1475,N_11,N_967);
xnor U1476 (N_1476,N_472,N_561);
or U1477 (N_1477,N_381,N_516);
nand U1478 (N_1478,N_87,N_531);
nor U1479 (N_1479,N_41,N_319);
nor U1480 (N_1480,N_696,N_537);
nor U1481 (N_1481,N_904,N_418);
and U1482 (N_1482,N_776,N_720);
nor U1483 (N_1483,N_25,N_886);
nand U1484 (N_1484,N_723,N_218);
nor U1485 (N_1485,N_943,N_334);
or U1486 (N_1486,N_553,N_446);
nand U1487 (N_1487,N_971,N_176);
or U1488 (N_1488,N_956,N_186);
nor U1489 (N_1489,N_22,N_73);
nand U1490 (N_1490,N_172,N_342);
nor U1491 (N_1491,N_370,N_425);
nand U1492 (N_1492,N_491,N_695);
and U1493 (N_1493,N_82,N_925);
and U1494 (N_1494,N_161,N_727);
nand U1495 (N_1495,N_584,N_8);
or U1496 (N_1496,N_671,N_300);
nand U1497 (N_1497,N_259,N_403);
nor U1498 (N_1498,N_984,N_0);
xor U1499 (N_1499,N_689,N_757);
nor U1500 (N_1500,N_26,N_39);
nor U1501 (N_1501,N_702,N_674);
and U1502 (N_1502,N_300,N_884);
or U1503 (N_1503,N_186,N_738);
xor U1504 (N_1504,N_114,N_164);
nor U1505 (N_1505,N_339,N_632);
and U1506 (N_1506,N_740,N_291);
nand U1507 (N_1507,N_467,N_798);
xnor U1508 (N_1508,N_165,N_787);
nand U1509 (N_1509,N_330,N_477);
or U1510 (N_1510,N_442,N_716);
nand U1511 (N_1511,N_473,N_558);
nand U1512 (N_1512,N_855,N_554);
xor U1513 (N_1513,N_953,N_723);
and U1514 (N_1514,N_510,N_181);
nor U1515 (N_1515,N_588,N_189);
and U1516 (N_1516,N_28,N_771);
and U1517 (N_1517,N_860,N_333);
nor U1518 (N_1518,N_221,N_812);
or U1519 (N_1519,N_805,N_423);
and U1520 (N_1520,N_69,N_311);
xnor U1521 (N_1521,N_513,N_225);
nand U1522 (N_1522,N_484,N_619);
xnor U1523 (N_1523,N_181,N_784);
nand U1524 (N_1524,N_303,N_719);
nand U1525 (N_1525,N_30,N_744);
and U1526 (N_1526,N_209,N_117);
and U1527 (N_1527,N_436,N_107);
or U1528 (N_1528,N_100,N_962);
and U1529 (N_1529,N_649,N_143);
or U1530 (N_1530,N_637,N_222);
and U1531 (N_1531,N_967,N_431);
nand U1532 (N_1532,N_5,N_17);
and U1533 (N_1533,N_277,N_752);
nor U1534 (N_1534,N_383,N_86);
nor U1535 (N_1535,N_942,N_122);
and U1536 (N_1536,N_24,N_212);
nor U1537 (N_1537,N_93,N_75);
nor U1538 (N_1538,N_54,N_520);
nand U1539 (N_1539,N_297,N_484);
and U1540 (N_1540,N_497,N_977);
nor U1541 (N_1541,N_301,N_645);
or U1542 (N_1542,N_209,N_829);
nand U1543 (N_1543,N_622,N_663);
nand U1544 (N_1544,N_746,N_765);
xnor U1545 (N_1545,N_120,N_817);
nand U1546 (N_1546,N_40,N_84);
or U1547 (N_1547,N_336,N_553);
and U1548 (N_1548,N_320,N_777);
or U1549 (N_1549,N_580,N_581);
nor U1550 (N_1550,N_166,N_372);
xnor U1551 (N_1551,N_682,N_700);
or U1552 (N_1552,N_753,N_463);
and U1553 (N_1553,N_793,N_648);
or U1554 (N_1554,N_482,N_906);
nor U1555 (N_1555,N_585,N_939);
or U1556 (N_1556,N_850,N_202);
xnor U1557 (N_1557,N_83,N_766);
and U1558 (N_1558,N_40,N_759);
and U1559 (N_1559,N_968,N_730);
nand U1560 (N_1560,N_610,N_369);
nand U1561 (N_1561,N_116,N_597);
nand U1562 (N_1562,N_852,N_593);
nor U1563 (N_1563,N_532,N_385);
nor U1564 (N_1564,N_544,N_413);
and U1565 (N_1565,N_205,N_887);
and U1566 (N_1566,N_611,N_319);
and U1567 (N_1567,N_804,N_532);
nand U1568 (N_1568,N_796,N_121);
or U1569 (N_1569,N_56,N_278);
or U1570 (N_1570,N_437,N_232);
or U1571 (N_1571,N_248,N_371);
nor U1572 (N_1572,N_894,N_947);
nand U1573 (N_1573,N_944,N_366);
and U1574 (N_1574,N_659,N_770);
nor U1575 (N_1575,N_70,N_854);
and U1576 (N_1576,N_418,N_387);
nand U1577 (N_1577,N_497,N_618);
nor U1578 (N_1578,N_331,N_899);
nor U1579 (N_1579,N_850,N_586);
or U1580 (N_1580,N_798,N_499);
and U1581 (N_1581,N_135,N_990);
or U1582 (N_1582,N_436,N_864);
nor U1583 (N_1583,N_396,N_405);
nor U1584 (N_1584,N_967,N_792);
nor U1585 (N_1585,N_674,N_539);
and U1586 (N_1586,N_759,N_373);
nand U1587 (N_1587,N_532,N_152);
or U1588 (N_1588,N_813,N_294);
and U1589 (N_1589,N_636,N_221);
nor U1590 (N_1590,N_353,N_784);
nand U1591 (N_1591,N_364,N_801);
nor U1592 (N_1592,N_240,N_576);
nor U1593 (N_1593,N_948,N_852);
nand U1594 (N_1594,N_50,N_308);
nand U1595 (N_1595,N_841,N_223);
and U1596 (N_1596,N_366,N_456);
nor U1597 (N_1597,N_152,N_563);
and U1598 (N_1598,N_882,N_381);
and U1599 (N_1599,N_278,N_868);
and U1600 (N_1600,N_17,N_559);
xnor U1601 (N_1601,N_779,N_28);
nand U1602 (N_1602,N_476,N_770);
and U1603 (N_1603,N_509,N_573);
and U1604 (N_1604,N_399,N_844);
xor U1605 (N_1605,N_112,N_8);
nor U1606 (N_1606,N_450,N_679);
nor U1607 (N_1607,N_378,N_32);
nand U1608 (N_1608,N_942,N_81);
xnor U1609 (N_1609,N_212,N_69);
or U1610 (N_1610,N_848,N_496);
nor U1611 (N_1611,N_902,N_51);
or U1612 (N_1612,N_869,N_984);
or U1613 (N_1613,N_336,N_12);
or U1614 (N_1614,N_792,N_353);
or U1615 (N_1615,N_275,N_957);
and U1616 (N_1616,N_798,N_282);
nor U1617 (N_1617,N_387,N_285);
or U1618 (N_1618,N_588,N_989);
or U1619 (N_1619,N_607,N_284);
and U1620 (N_1620,N_57,N_966);
nor U1621 (N_1621,N_183,N_765);
nor U1622 (N_1622,N_795,N_812);
nor U1623 (N_1623,N_89,N_203);
xor U1624 (N_1624,N_506,N_91);
nand U1625 (N_1625,N_462,N_289);
or U1626 (N_1626,N_191,N_150);
or U1627 (N_1627,N_776,N_996);
nor U1628 (N_1628,N_373,N_109);
or U1629 (N_1629,N_368,N_426);
nand U1630 (N_1630,N_561,N_577);
nor U1631 (N_1631,N_126,N_975);
nand U1632 (N_1632,N_445,N_834);
xnor U1633 (N_1633,N_549,N_343);
or U1634 (N_1634,N_362,N_752);
or U1635 (N_1635,N_987,N_303);
or U1636 (N_1636,N_661,N_978);
nor U1637 (N_1637,N_196,N_946);
and U1638 (N_1638,N_47,N_777);
and U1639 (N_1639,N_401,N_567);
and U1640 (N_1640,N_419,N_570);
nand U1641 (N_1641,N_293,N_434);
and U1642 (N_1642,N_111,N_157);
and U1643 (N_1643,N_285,N_267);
or U1644 (N_1644,N_880,N_864);
nand U1645 (N_1645,N_731,N_100);
nand U1646 (N_1646,N_147,N_493);
nand U1647 (N_1647,N_295,N_330);
nor U1648 (N_1648,N_114,N_55);
or U1649 (N_1649,N_931,N_160);
xor U1650 (N_1650,N_427,N_736);
or U1651 (N_1651,N_241,N_283);
nor U1652 (N_1652,N_543,N_511);
nor U1653 (N_1653,N_414,N_137);
nor U1654 (N_1654,N_737,N_263);
or U1655 (N_1655,N_162,N_995);
nand U1656 (N_1656,N_160,N_801);
xnor U1657 (N_1657,N_388,N_828);
nor U1658 (N_1658,N_931,N_749);
and U1659 (N_1659,N_638,N_64);
or U1660 (N_1660,N_98,N_185);
or U1661 (N_1661,N_898,N_61);
or U1662 (N_1662,N_567,N_62);
and U1663 (N_1663,N_783,N_484);
xor U1664 (N_1664,N_537,N_94);
xor U1665 (N_1665,N_297,N_643);
nor U1666 (N_1666,N_564,N_555);
and U1667 (N_1667,N_717,N_323);
nand U1668 (N_1668,N_276,N_675);
or U1669 (N_1669,N_217,N_770);
and U1670 (N_1670,N_163,N_868);
or U1671 (N_1671,N_197,N_522);
nor U1672 (N_1672,N_501,N_31);
and U1673 (N_1673,N_682,N_939);
nand U1674 (N_1674,N_849,N_356);
or U1675 (N_1675,N_695,N_251);
nand U1676 (N_1676,N_794,N_945);
or U1677 (N_1677,N_988,N_696);
nor U1678 (N_1678,N_84,N_322);
and U1679 (N_1679,N_23,N_662);
nor U1680 (N_1680,N_624,N_625);
xnor U1681 (N_1681,N_449,N_64);
and U1682 (N_1682,N_125,N_404);
xnor U1683 (N_1683,N_523,N_308);
nor U1684 (N_1684,N_719,N_864);
nor U1685 (N_1685,N_703,N_511);
nand U1686 (N_1686,N_552,N_550);
or U1687 (N_1687,N_202,N_583);
and U1688 (N_1688,N_845,N_582);
or U1689 (N_1689,N_995,N_697);
nand U1690 (N_1690,N_193,N_119);
nor U1691 (N_1691,N_88,N_654);
or U1692 (N_1692,N_770,N_567);
nand U1693 (N_1693,N_968,N_703);
nand U1694 (N_1694,N_677,N_384);
nor U1695 (N_1695,N_27,N_938);
nand U1696 (N_1696,N_672,N_387);
nor U1697 (N_1697,N_197,N_78);
or U1698 (N_1698,N_180,N_261);
or U1699 (N_1699,N_698,N_802);
xnor U1700 (N_1700,N_132,N_344);
or U1701 (N_1701,N_889,N_351);
nand U1702 (N_1702,N_284,N_625);
and U1703 (N_1703,N_956,N_1);
or U1704 (N_1704,N_702,N_696);
nand U1705 (N_1705,N_868,N_817);
xor U1706 (N_1706,N_177,N_208);
and U1707 (N_1707,N_860,N_90);
nand U1708 (N_1708,N_31,N_766);
nor U1709 (N_1709,N_520,N_424);
or U1710 (N_1710,N_219,N_338);
xnor U1711 (N_1711,N_374,N_302);
nor U1712 (N_1712,N_710,N_792);
and U1713 (N_1713,N_7,N_991);
and U1714 (N_1714,N_59,N_233);
or U1715 (N_1715,N_359,N_599);
nor U1716 (N_1716,N_459,N_520);
xor U1717 (N_1717,N_291,N_176);
nand U1718 (N_1718,N_293,N_107);
and U1719 (N_1719,N_621,N_537);
or U1720 (N_1720,N_558,N_784);
xor U1721 (N_1721,N_792,N_764);
or U1722 (N_1722,N_167,N_721);
xnor U1723 (N_1723,N_486,N_743);
nand U1724 (N_1724,N_359,N_903);
nor U1725 (N_1725,N_844,N_710);
xor U1726 (N_1726,N_555,N_614);
nand U1727 (N_1727,N_389,N_896);
or U1728 (N_1728,N_510,N_137);
and U1729 (N_1729,N_320,N_820);
nor U1730 (N_1730,N_791,N_325);
and U1731 (N_1731,N_427,N_295);
nand U1732 (N_1732,N_19,N_344);
nor U1733 (N_1733,N_251,N_758);
and U1734 (N_1734,N_103,N_967);
nand U1735 (N_1735,N_488,N_743);
or U1736 (N_1736,N_719,N_680);
nor U1737 (N_1737,N_296,N_114);
or U1738 (N_1738,N_761,N_196);
and U1739 (N_1739,N_160,N_273);
nand U1740 (N_1740,N_92,N_798);
xnor U1741 (N_1741,N_1,N_164);
xnor U1742 (N_1742,N_369,N_142);
nand U1743 (N_1743,N_940,N_102);
nor U1744 (N_1744,N_487,N_657);
or U1745 (N_1745,N_821,N_216);
and U1746 (N_1746,N_217,N_673);
nand U1747 (N_1747,N_42,N_391);
xor U1748 (N_1748,N_73,N_146);
nand U1749 (N_1749,N_235,N_368);
nor U1750 (N_1750,N_219,N_314);
and U1751 (N_1751,N_651,N_533);
and U1752 (N_1752,N_434,N_666);
nor U1753 (N_1753,N_169,N_656);
nand U1754 (N_1754,N_562,N_131);
nor U1755 (N_1755,N_469,N_813);
and U1756 (N_1756,N_588,N_548);
nor U1757 (N_1757,N_186,N_226);
or U1758 (N_1758,N_701,N_699);
nand U1759 (N_1759,N_919,N_184);
nand U1760 (N_1760,N_656,N_354);
or U1761 (N_1761,N_965,N_294);
and U1762 (N_1762,N_949,N_53);
and U1763 (N_1763,N_374,N_20);
nor U1764 (N_1764,N_341,N_309);
and U1765 (N_1765,N_607,N_726);
or U1766 (N_1766,N_812,N_178);
nor U1767 (N_1767,N_247,N_44);
nor U1768 (N_1768,N_966,N_127);
nor U1769 (N_1769,N_569,N_615);
nor U1770 (N_1770,N_919,N_476);
xor U1771 (N_1771,N_360,N_892);
nand U1772 (N_1772,N_124,N_309);
and U1773 (N_1773,N_3,N_643);
xnor U1774 (N_1774,N_426,N_940);
nand U1775 (N_1775,N_112,N_184);
nand U1776 (N_1776,N_964,N_189);
nor U1777 (N_1777,N_0,N_272);
and U1778 (N_1778,N_381,N_687);
or U1779 (N_1779,N_429,N_350);
nor U1780 (N_1780,N_413,N_207);
or U1781 (N_1781,N_115,N_242);
nor U1782 (N_1782,N_37,N_589);
and U1783 (N_1783,N_253,N_256);
or U1784 (N_1784,N_543,N_851);
nand U1785 (N_1785,N_465,N_2);
nor U1786 (N_1786,N_63,N_497);
nand U1787 (N_1787,N_235,N_950);
and U1788 (N_1788,N_57,N_59);
or U1789 (N_1789,N_1,N_281);
or U1790 (N_1790,N_155,N_363);
nor U1791 (N_1791,N_401,N_114);
or U1792 (N_1792,N_811,N_130);
or U1793 (N_1793,N_493,N_80);
nand U1794 (N_1794,N_984,N_786);
nand U1795 (N_1795,N_72,N_457);
or U1796 (N_1796,N_66,N_652);
or U1797 (N_1797,N_517,N_246);
or U1798 (N_1798,N_960,N_222);
and U1799 (N_1799,N_551,N_561);
and U1800 (N_1800,N_283,N_505);
and U1801 (N_1801,N_351,N_961);
or U1802 (N_1802,N_784,N_459);
or U1803 (N_1803,N_594,N_960);
or U1804 (N_1804,N_714,N_88);
nand U1805 (N_1805,N_986,N_496);
nand U1806 (N_1806,N_983,N_893);
nor U1807 (N_1807,N_196,N_676);
nand U1808 (N_1808,N_753,N_820);
and U1809 (N_1809,N_149,N_422);
nor U1810 (N_1810,N_38,N_480);
nor U1811 (N_1811,N_858,N_568);
nand U1812 (N_1812,N_319,N_202);
nor U1813 (N_1813,N_399,N_170);
or U1814 (N_1814,N_361,N_344);
and U1815 (N_1815,N_530,N_624);
and U1816 (N_1816,N_749,N_866);
xnor U1817 (N_1817,N_224,N_853);
nor U1818 (N_1818,N_40,N_172);
xnor U1819 (N_1819,N_208,N_693);
and U1820 (N_1820,N_74,N_120);
nand U1821 (N_1821,N_481,N_563);
and U1822 (N_1822,N_950,N_287);
and U1823 (N_1823,N_530,N_973);
nand U1824 (N_1824,N_206,N_549);
nor U1825 (N_1825,N_851,N_635);
or U1826 (N_1826,N_142,N_693);
or U1827 (N_1827,N_210,N_684);
or U1828 (N_1828,N_325,N_221);
xnor U1829 (N_1829,N_619,N_463);
or U1830 (N_1830,N_767,N_906);
nand U1831 (N_1831,N_900,N_747);
nor U1832 (N_1832,N_28,N_47);
nand U1833 (N_1833,N_17,N_78);
or U1834 (N_1834,N_836,N_753);
nor U1835 (N_1835,N_306,N_856);
xnor U1836 (N_1836,N_616,N_715);
xnor U1837 (N_1837,N_347,N_17);
and U1838 (N_1838,N_930,N_376);
or U1839 (N_1839,N_447,N_801);
nor U1840 (N_1840,N_108,N_116);
and U1841 (N_1841,N_30,N_798);
nor U1842 (N_1842,N_546,N_790);
and U1843 (N_1843,N_128,N_308);
or U1844 (N_1844,N_859,N_261);
or U1845 (N_1845,N_664,N_936);
nand U1846 (N_1846,N_415,N_480);
and U1847 (N_1847,N_740,N_534);
nor U1848 (N_1848,N_763,N_746);
and U1849 (N_1849,N_175,N_570);
or U1850 (N_1850,N_423,N_900);
nand U1851 (N_1851,N_357,N_90);
nor U1852 (N_1852,N_295,N_378);
nand U1853 (N_1853,N_217,N_83);
nand U1854 (N_1854,N_408,N_615);
and U1855 (N_1855,N_663,N_931);
nor U1856 (N_1856,N_137,N_15);
or U1857 (N_1857,N_905,N_344);
nor U1858 (N_1858,N_333,N_141);
nor U1859 (N_1859,N_424,N_973);
or U1860 (N_1860,N_784,N_502);
nor U1861 (N_1861,N_395,N_146);
or U1862 (N_1862,N_27,N_853);
xnor U1863 (N_1863,N_504,N_790);
and U1864 (N_1864,N_203,N_629);
or U1865 (N_1865,N_758,N_493);
nor U1866 (N_1866,N_240,N_217);
nand U1867 (N_1867,N_240,N_69);
xnor U1868 (N_1868,N_239,N_781);
nand U1869 (N_1869,N_328,N_0);
or U1870 (N_1870,N_53,N_994);
nor U1871 (N_1871,N_187,N_62);
xnor U1872 (N_1872,N_53,N_967);
nor U1873 (N_1873,N_8,N_249);
nor U1874 (N_1874,N_673,N_730);
or U1875 (N_1875,N_574,N_317);
or U1876 (N_1876,N_680,N_232);
nand U1877 (N_1877,N_242,N_149);
and U1878 (N_1878,N_668,N_418);
or U1879 (N_1879,N_868,N_624);
xor U1880 (N_1880,N_161,N_208);
nand U1881 (N_1881,N_532,N_901);
or U1882 (N_1882,N_407,N_266);
or U1883 (N_1883,N_526,N_492);
or U1884 (N_1884,N_75,N_526);
and U1885 (N_1885,N_866,N_660);
nor U1886 (N_1886,N_835,N_737);
nand U1887 (N_1887,N_968,N_183);
nand U1888 (N_1888,N_866,N_802);
nand U1889 (N_1889,N_7,N_193);
nor U1890 (N_1890,N_113,N_471);
or U1891 (N_1891,N_676,N_613);
nand U1892 (N_1892,N_772,N_998);
nor U1893 (N_1893,N_355,N_169);
and U1894 (N_1894,N_6,N_423);
nand U1895 (N_1895,N_93,N_328);
nand U1896 (N_1896,N_923,N_38);
or U1897 (N_1897,N_160,N_428);
nand U1898 (N_1898,N_452,N_169);
nand U1899 (N_1899,N_684,N_345);
and U1900 (N_1900,N_419,N_731);
and U1901 (N_1901,N_427,N_465);
nor U1902 (N_1902,N_437,N_434);
nand U1903 (N_1903,N_761,N_419);
xnor U1904 (N_1904,N_872,N_430);
xor U1905 (N_1905,N_815,N_181);
or U1906 (N_1906,N_192,N_98);
nand U1907 (N_1907,N_386,N_909);
nand U1908 (N_1908,N_620,N_44);
xor U1909 (N_1909,N_281,N_435);
xnor U1910 (N_1910,N_418,N_311);
and U1911 (N_1911,N_314,N_414);
nor U1912 (N_1912,N_916,N_777);
or U1913 (N_1913,N_199,N_694);
nor U1914 (N_1914,N_125,N_111);
xor U1915 (N_1915,N_302,N_746);
or U1916 (N_1916,N_805,N_880);
xor U1917 (N_1917,N_872,N_383);
nand U1918 (N_1918,N_290,N_995);
nor U1919 (N_1919,N_985,N_9);
nand U1920 (N_1920,N_232,N_296);
or U1921 (N_1921,N_79,N_990);
nor U1922 (N_1922,N_711,N_851);
nor U1923 (N_1923,N_949,N_216);
or U1924 (N_1924,N_574,N_652);
or U1925 (N_1925,N_268,N_615);
nand U1926 (N_1926,N_270,N_115);
nor U1927 (N_1927,N_708,N_727);
or U1928 (N_1928,N_517,N_854);
and U1929 (N_1929,N_912,N_362);
or U1930 (N_1930,N_319,N_690);
and U1931 (N_1931,N_270,N_311);
nand U1932 (N_1932,N_692,N_841);
and U1933 (N_1933,N_206,N_967);
or U1934 (N_1934,N_705,N_815);
xor U1935 (N_1935,N_427,N_196);
and U1936 (N_1936,N_855,N_473);
nor U1937 (N_1937,N_303,N_229);
and U1938 (N_1938,N_443,N_603);
nand U1939 (N_1939,N_628,N_340);
nand U1940 (N_1940,N_125,N_712);
and U1941 (N_1941,N_489,N_209);
nor U1942 (N_1942,N_75,N_674);
nor U1943 (N_1943,N_13,N_835);
or U1944 (N_1944,N_989,N_577);
xor U1945 (N_1945,N_476,N_316);
or U1946 (N_1946,N_658,N_67);
nor U1947 (N_1947,N_558,N_444);
or U1948 (N_1948,N_639,N_89);
or U1949 (N_1949,N_798,N_705);
nor U1950 (N_1950,N_126,N_236);
xnor U1951 (N_1951,N_124,N_120);
nor U1952 (N_1952,N_807,N_909);
and U1953 (N_1953,N_894,N_327);
nand U1954 (N_1954,N_892,N_273);
nor U1955 (N_1955,N_258,N_145);
nor U1956 (N_1956,N_79,N_694);
or U1957 (N_1957,N_845,N_325);
and U1958 (N_1958,N_475,N_190);
or U1959 (N_1959,N_982,N_722);
nand U1960 (N_1960,N_728,N_515);
or U1961 (N_1961,N_984,N_22);
nand U1962 (N_1962,N_406,N_614);
or U1963 (N_1963,N_539,N_16);
nand U1964 (N_1964,N_414,N_473);
and U1965 (N_1965,N_292,N_420);
and U1966 (N_1966,N_700,N_598);
nor U1967 (N_1967,N_356,N_959);
nor U1968 (N_1968,N_118,N_724);
nand U1969 (N_1969,N_590,N_73);
or U1970 (N_1970,N_66,N_203);
and U1971 (N_1971,N_397,N_980);
nor U1972 (N_1972,N_675,N_847);
nor U1973 (N_1973,N_387,N_147);
or U1974 (N_1974,N_968,N_709);
and U1975 (N_1975,N_794,N_982);
or U1976 (N_1976,N_152,N_570);
nor U1977 (N_1977,N_980,N_368);
nor U1978 (N_1978,N_577,N_235);
or U1979 (N_1979,N_506,N_851);
nand U1980 (N_1980,N_156,N_552);
nand U1981 (N_1981,N_470,N_432);
or U1982 (N_1982,N_577,N_174);
nor U1983 (N_1983,N_57,N_226);
nand U1984 (N_1984,N_60,N_80);
and U1985 (N_1985,N_90,N_468);
nand U1986 (N_1986,N_285,N_229);
nor U1987 (N_1987,N_57,N_760);
or U1988 (N_1988,N_402,N_299);
nand U1989 (N_1989,N_404,N_214);
xnor U1990 (N_1990,N_446,N_137);
xnor U1991 (N_1991,N_683,N_483);
nand U1992 (N_1992,N_660,N_813);
xor U1993 (N_1993,N_308,N_585);
and U1994 (N_1994,N_578,N_916);
xor U1995 (N_1995,N_904,N_716);
nand U1996 (N_1996,N_461,N_401);
nand U1997 (N_1997,N_531,N_209);
nor U1998 (N_1998,N_150,N_558);
nor U1999 (N_1999,N_427,N_488);
or U2000 (N_2000,N_1883,N_1029);
and U2001 (N_2001,N_1367,N_1688);
nand U2002 (N_2002,N_1739,N_1473);
or U2003 (N_2003,N_1487,N_1421);
nand U2004 (N_2004,N_1162,N_1842);
nor U2005 (N_2005,N_1881,N_1951);
or U2006 (N_2006,N_1348,N_1661);
and U2007 (N_2007,N_1787,N_1003);
xor U2008 (N_2008,N_1685,N_1146);
nor U2009 (N_2009,N_1167,N_1806);
nand U2010 (N_2010,N_1343,N_1605);
nor U2011 (N_2011,N_1975,N_1347);
nand U2012 (N_2012,N_1648,N_1283);
or U2013 (N_2013,N_1838,N_1490);
and U2014 (N_2014,N_1371,N_1115);
xor U2015 (N_2015,N_1668,N_1135);
nor U2016 (N_2016,N_1525,N_1043);
or U2017 (N_2017,N_1982,N_1464);
xor U2018 (N_2018,N_1048,N_1608);
or U2019 (N_2019,N_1789,N_1878);
nand U2020 (N_2020,N_1887,N_1895);
nand U2021 (N_2021,N_1234,N_1851);
and U2022 (N_2022,N_1216,N_1528);
and U2023 (N_2023,N_1164,N_1751);
nand U2024 (N_2024,N_1529,N_1932);
nand U2025 (N_2025,N_1736,N_1361);
nor U2026 (N_2026,N_1405,N_1433);
and U2027 (N_2027,N_1839,N_1402);
nand U2028 (N_2028,N_1293,N_1779);
and U2029 (N_2029,N_1626,N_1259);
xor U2030 (N_2030,N_1733,N_1209);
nand U2031 (N_2031,N_1847,N_1854);
or U2032 (N_2032,N_1319,N_1694);
or U2033 (N_2033,N_1239,N_1340);
and U2034 (N_2034,N_1019,N_1336);
nor U2035 (N_2035,N_1142,N_1993);
nand U2036 (N_2036,N_1501,N_1756);
or U2037 (N_2037,N_1709,N_1317);
nand U2038 (N_2038,N_1510,N_1168);
and U2039 (N_2039,N_1492,N_1531);
nor U2040 (N_2040,N_1075,N_1084);
or U2041 (N_2041,N_1395,N_1765);
and U2042 (N_2042,N_1461,N_1800);
nor U2043 (N_2043,N_1231,N_1355);
or U2044 (N_2044,N_1938,N_1737);
and U2045 (N_2045,N_1623,N_1536);
nor U2046 (N_2046,N_1578,N_1248);
nor U2047 (N_2047,N_1811,N_1260);
xor U2048 (N_2048,N_1426,N_1675);
nor U2049 (N_2049,N_1962,N_1474);
or U2050 (N_2050,N_1724,N_1449);
and U2051 (N_2051,N_1049,N_1273);
or U2052 (N_2052,N_1123,N_1390);
or U2053 (N_2053,N_1140,N_1611);
nand U2054 (N_2054,N_1151,N_1750);
or U2055 (N_2055,N_1870,N_1296);
nand U2056 (N_2056,N_1833,N_1483);
or U2057 (N_2057,N_1555,N_1440);
nand U2058 (N_2058,N_1022,N_1882);
xor U2059 (N_2059,N_1398,N_1324);
nor U2060 (N_2060,N_1908,N_1238);
nand U2061 (N_2061,N_1144,N_1108);
nand U2062 (N_2062,N_1557,N_1481);
or U2063 (N_2063,N_1337,N_1120);
and U2064 (N_2064,N_1934,N_1314);
and U2065 (N_2065,N_1432,N_1969);
and U2066 (N_2066,N_1808,N_1069);
or U2067 (N_2067,N_1233,N_1393);
nor U2068 (N_2068,N_1752,N_1153);
nor U2069 (N_2069,N_1727,N_1587);
nor U2070 (N_2070,N_1715,N_1015);
nor U2071 (N_2071,N_1793,N_1147);
xor U2072 (N_2072,N_1594,N_1313);
nor U2073 (N_2073,N_1845,N_1877);
nand U2074 (N_2074,N_1519,N_1760);
and U2075 (N_2075,N_1219,N_1307);
xor U2076 (N_2076,N_1287,N_1482);
nand U2077 (N_2077,N_1170,N_1024);
and U2078 (N_2078,N_1601,N_1182);
and U2079 (N_2079,N_1013,N_1628);
nand U2080 (N_2080,N_1974,N_1226);
xnor U2081 (N_2081,N_1602,N_1740);
nand U2082 (N_2082,N_1844,N_1677);
nor U2083 (N_2083,N_1191,N_1921);
nand U2084 (N_2084,N_1837,N_1965);
or U2085 (N_2085,N_1571,N_1448);
or U2086 (N_2086,N_1849,N_1082);
nor U2087 (N_2087,N_1865,N_1673);
or U2088 (N_2088,N_1949,N_1918);
or U2089 (N_2089,N_1547,N_1128);
or U2090 (N_2090,N_1420,N_1880);
and U2091 (N_2091,N_1505,N_1796);
or U2092 (N_2092,N_1526,N_1667);
nand U2093 (N_2093,N_1696,N_1595);
nand U2094 (N_2094,N_1972,N_1381);
or U2095 (N_2095,N_1286,N_1753);
and U2096 (N_2096,N_1879,N_1744);
nor U2097 (N_2097,N_1979,N_1443);
or U2098 (N_2098,N_1901,N_1925);
and U2099 (N_2099,N_1928,N_1585);
and U2100 (N_2100,N_1590,N_1141);
and U2101 (N_2101,N_1615,N_1558);
xnor U2102 (N_2102,N_1459,N_1358);
nand U2103 (N_2103,N_1859,N_1717);
nand U2104 (N_2104,N_1251,N_1772);
and U2105 (N_2105,N_1775,N_1954);
and U2106 (N_2106,N_1624,N_1645);
nor U2107 (N_2107,N_1068,N_1155);
or U2108 (N_2108,N_1955,N_1281);
and U2109 (N_2109,N_1995,N_1549);
nor U2110 (N_2110,N_1388,N_1994);
nand U2111 (N_2111,N_1984,N_1256);
nor U2112 (N_2112,N_1726,N_1771);
nand U2113 (N_2113,N_1897,N_1607);
and U2114 (N_2114,N_1657,N_1819);
nor U2115 (N_2115,N_1521,N_1695);
nand U2116 (N_2116,N_1349,N_1679);
nand U2117 (N_2117,N_1697,N_1438);
nand U2118 (N_2118,N_1264,N_1091);
nor U2119 (N_2119,N_1241,N_1812);
and U2120 (N_2120,N_1655,N_1758);
nand U2121 (N_2121,N_1941,N_1570);
or U2122 (N_2122,N_1574,N_1647);
and U2123 (N_2123,N_1412,N_1825);
nand U2124 (N_2124,N_1020,N_1242);
nor U2125 (N_2125,N_1189,N_1814);
xnor U2126 (N_2126,N_1397,N_1413);
and U2127 (N_2127,N_1614,N_1391);
and U2128 (N_2128,N_1504,N_1052);
nor U2129 (N_2129,N_1406,N_1818);
or U2130 (N_2130,N_1143,N_1940);
or U2131 (N_2131,N_1042,N_1738);
or U2132 (N_2132,N_1408,N_1550);
or U2133 (N_2133,N_1996,N_1923);
nand U2134 (N_2134,N_1165,N_1205);
nor U2135 (N_2135,N_1554,N_1915);
nor U2136 (N_2136,N_1236,N_1279);
and U2137 (N_2137,N_1471,N_1725);
and U2138 (N_2138,N_1537,N_1705);
nand U2139 (N_2139,N_1781,N_1272);
nor U2140 (N_2140,N_1097,N_1890);
and U2141 (N_2141,N_1630,N_1342);
xor U2142 (N_2142,N_1593,N_1576);
nand U2143 (N_2143,N_1306,N_1861);
nor U2144 (N_2144,N_1060,N_1245);
and U2145 (N_2145,N_1442,N_1992);
nor U2146 (N_2146,N_1354,N_1382);
nor U2147 (N_2147,N_1129,N_1439);
nand U2148 (N_2148,N_1184,N_1201);
nor U2149 (N_2149,N_1327,N_1429);
or U2150 (N_2150,N_1517,N_1889);
and U2151 (N_2151,N_1058,N_1700);
nand U2152 (N_2152,N_1683,N_1004);
or U2153 (N_2153,N_1916,N_1088);
or U2154 (N_2154,N_1553,N_1090);
nor U2155 (N_2155,N_1672,N_1378);
or U2156 (N_2156,N_1435,N_1425);
nand U2157 (N_2157,N_1821,N_1629);
nor U2158 (N_2158,N_1404,N_1308);
xnor U2159 (N_2159,N_1360,N_1055);
or U2160 (N_2160,N_1855,N_1112);
nand U2161 (N_2161,N_1802,N_1565);
or U2162 (N_2162,N_1431,N_1912);
nor U2163 (N_2163,N_1476,N_1546);
nand U2164 (N_2164,N_1947,N_1805);
or U2165 (N_2165,N_1017,N_1458);
xnor U2166 (N_2166,N_1479,N_1176);
nor U2167 (N_2167,N_1285,N_1809);
or U2168 (N_2168,N_1621,N_1706);
or U2169 (N_2169,N_1244,N_1970);
nand U2170 (N_2170,N_1664,N_1935);
and U2171 (N_2171,N_1180,N_1930);
nand U2172 (N_2172,N_1310,N_1542);
or U2173 (N_2173,N_1380,N_1376);
and U2174 (N_2174,N_1640,N_1454);
nand U2175 (N_2175,N_1896,N_1261);
or U2176 (N_2176,N_1530,N_1902);
nand U2177 (N_2177,N_1061,N_1552);
and U2178 (N_2178,N_1037,N_1514);
xnor U2179 (N_2179,N_1633,N_1400);
nor U2180 (N_2180,N_1929,N_1289);
nor U2181 (N_2181,N_1823,N_1888);
and U2182 (N_2182,N_1669,N_1062);
and U2183 (N_2183,N_1864,N_1522);
and U2184 (N_2184,N_1172,N_1866);
or U2185 (N_2185,N_1116,N_1145);
and U2186 (N_2186,N_1315,N_1338);
nor U2187 (N_2187,N_1704,N_1952);
and U2188 (N_2188,N_1192,N_1494);
and U2189 (N_2189,N_1462,N_1794);
nor U2190 (N_2190,N_1009,N_1227);
or U2191 (N_2191,N_1689,N_1292);
or U2192 (N_2192,N_1228,N_1436);
or U2193 (N_2193,N_1222,N_1268);
and U2194 (N_2194,N_1790,N_1067);
and U2195 (N_2195,N_1240,N_1920);
nor U2196 (N_2196,N_1508,N_1687);
or U2197 (N_2197,N_1444,N_1910);
or U2198 (N_2198,N_1121,N_1712);
or U2199 (N_2199,N_1945,N_1783);
or U2200 (N_2200,N_1913,N_1497);
or U2201 (N_2201,N_1803,N_1111);
nor U2202 (N_2202,N_1356,N_1014);
or U2203 (N_2203,N_1654,N_1316);
nor U2204 (N_2204,N_1196,N_1956);
nor U2205 (N_2205,N_1339,N_1914);
xnor U2206 (N_2206,N_1034,N_1099);
or U2207 (N_2207,N_1755,N_1869);
or U2208 (N_2208,N_1345,N_1187);
nand U2209 (N_2209,N_1843,N_1110);
nor U2210 (N_2210,N_1350,N_1074);
or U2211 (N_2211,N_1702,N_1502);
and U2212 (N_2212,N_1506,N_1560);
or U2213 (N_2213,N_1489,N_1991);
nand U2214 (N_2214,N_1046,N_1225);
xor U2215 (N_2215,N_1987,N_1266);
xor U2216 (N_2216,N_1967,N_1942);
nor U2217 (N_2217,N_1538,N_1762);
xor U2218 (N_2218,N_1416,N_1212);
nor U2219 (N_2219,N_1032,N_1224);
nand U2220 (N_2220,N_1711,N_1002);
nand U2221 (N_2221,N_1617,N_1276);
nand U2222 (N_2222,N_1853,N_1229);
nand U2223 (N_2223,N_1036,N_1562);
nand U2224 (N_2224,N_1159,N_1769);
or U2225 (N_2225,N_1714,N_1832);
or U2226 (N_2226,N_1114,N_1499);
xnor U2227 (N_2227,N_1858,N_1173);
and U2228 (N_2228,N_1214,N_1957);
nand U2229 (N_2229,N_1682,N_1723);
or U2230 (N_2230,N_1437,N_1076);
nand U2231 (N_2231,N_1252,N_1978);
nor U2232 (N_2232,N_1516,N_1813);
or U2233 (N_2233,N_1867,N_1101);
nor U2234 (N_2234,N_1953,N_1038);
nor U2235 (N_2235,N_1950,N_1312);
and U2236 (N_2236,N_1986,N_1094);
or U2237 (N_2237,N_1177,N_1399);
nand U2238 (N_2238,N_1963,N_1797);
nand U2239 (N_2239,N_1917,N_1690);
xnor U2240 (N_2240,N_1323,N_1884);
nand U2241 (N_2241,N_1417,N_1840);
nand U2242 (N_2242,N_1761,N_1362);
nor U2243 (N_2243,N_1495,N_1670);
nor U2244 (N_2244,N_1188,N_1335);
and U2245 (N_2245,N_1302,N_1721);
nor U2246 (N_2246,N_1044,N_1290);
nor U2247 (N_2247,N_1100,N_1305);
or U2248 (N_2248,N_1665,N_1613);
and U2249 (N_2249,N_1215,N_1749);
nor U2250 (N_2250,N_1053,N_1127);
or U2251 (N_2251,N_1871,N_1211);
nor U2252 (N_2252,N_1786,N_1671);
nor U2253 (N_2253,N_1103,N_1894);
or U2254 (N_2254,N_1001,N_1485);
nor U2255 (N_2255,N_1007,N_1078);
or U2256 (N_2256,N_1588,N_1788);
and U2257 (N_2257,N_1325,N_1493);
nand U2258 (N_2258,N_1810,N_1085);
xnor U2259 (N_2259,N_1124,N_1270);
nand U2260 (N_2260,N_1057,N_1424);
or U2261 (N_2261,N_1937,N_1575);
xor U2262 (N_2262,N_1973,N_1401);
or U2263 (N_2263,N_1041,N_1269);
nand U2264 (N_2264,N_1518,N_1332);
nor U2265 (N_2265,N_1206,N_1634);
xor U2266 (N_2266,N_1079,N_1543);
and U2267 (N_2267,N_1523,N_1604);
and U2268 (N_2268,N_1780,N_1262);
xnor U2269 (N_2269,N_1568,N_1455);
nor U2270 (N_2270,N_1208,N_1357);
or U2271 (N_2271,N_1692,N_1389);
nand U2272 (N_2272,N_1300,N_1359);
or U2273 (N_2273,N_1784,N_1072);
or U2274 (N_2274,N_1830,N_1743);
nand U2275 (N_2275,N_1311,N_1409);
nor U2276 (N_2276,N_1403,N_1383);
and U2277 (N_2277,N_1841,N_1021);
or U2278 (N_2278,N_1230,N_1713);
or U2279 (N_2279,N_1109,N_1478);
nand U2280 (N_2280,N_1081,N_1632);
nand U2281 (N_2281,N_1924,N_1544);
nor U2282 (N_2282,N_1469,N_1175);
or U2283 (N_2283,N_1720,N_1453);
nor U2284 (N_2284,N_1137,N_1083);
and U2285 (N_2285,N_1396,N_1451);
nor U2286 (N_2286,N_1581,N_1559);
or U2287 (N_2287,N_1092,N_1370);
or U2288 (N_2288,N_1681,N_1500);
xnor U2289 (N_2289,N_1735,N_1710);
xnor U2290 (N_2290,N_1777,N_1322);
nand U2291 (N_2291,N_1834,N_1318);
or U2292 (N_2292,N_1567,N_1520);
nand U2293 (N_2293,N_1663,N_1785);
or U2294 (N_2294,N_1641,N_1643);
and U2295 (N_2295,N_1152,N_1597);
or U2296 (N_2296,N_1139,N_1977);
xor U2297 (N_2297,N_1030,N_1158);
nor U2298 (N_2298,N_1829,N_1028);
nand U2299 (N_2299,N_1271,N_1330);
nor U2300 (N_2300,N_1255,N_1445);
xnor U2301 (N_2301,N_1816,N_1618);
and U2302 (N_2302,N_1759,N_1911);
or U2303 (N_2303,N_1535,N_1457);
nand U2304 (N_2304,N_1131,N_1768);
and U2305 (N_2305,N_1122,N_1958);
or U2306 (N_2306,N_1463,N_1250);
or U2307 (N_2307,N_1616,N_1394);
or U2308 (N_2308,N_1874,N_1686);
and U2309 (N_2309,N_1512,N_1798);
or U2310 (N_2310,N_1693,N_1698);
nand U2311 (N_2311,N_1876,N_1297);
nor U2312 (N_2312,N_1441,N_1792);
nor U2313 (N_2313,N_1625,N_1352);
nand U2314 (N_2314,N_1579,N_1148);
nor U2315 (N_2315,N_1232,N_1638);
and U2316 (N_2316,N_1366,N_1598);
nand U2317 (N_2317,N_1275,N_1080);
nand U2318 (N_2318,N_1922,N_1025);
nand U2319 (N_2319,N_1875,N_1363);
nor U2320 (N_2320,N_1527,N_1507);
and U2321 (N_2321,N_1386,N_1906);
nand U2322 (N_2322,N_1171,N_1334);
nor U2323 (N_2323,N_1933,N_1178);
nor U2324 (N_2324,N_1368,N_1005);
or U2325 (N_2325,N_1278,N_1646);
or U2326 (N_2326,N_1770,N_1249);
nor U2327 (N_2327,N_1364,N_1660);
or U2328 (N_2328,N_1631,N_1353);
xnor U2329 (N_2329,N_1873,N_1610);
xnor U2330 (N_2330,N_1541,N_1008);
or U2331 (N_2331,N_1218,N_1096);
and U2332 (N_2332,N_1235,N_1862);
nand U2333 (N_2333,N_1943,N_1221);
xnor U2334 (N_2334,N_1427,N_1320);
or U2335 (N_2335,N_1534,N_1466);
nand U2336 (N_2336,N_1545,N_1154);
xnor U2337 (N_2337,N_1946,N_1635);
or U2338 (N_2338,N_1467,N_1460);
and U2339 (N_2339,N_1596,N_1748);
nor U2340 (N_2340,N_1138,N_1680);
and U2341 (N_2341,N_1846,N_1826);
or U2342 (N_2342,N_1649,N_1220);
nand U2343 (N_2343,N_1326,N_1484);
nand U2344 (N_2344,N_1095,N_1971);
and U2345 (N_2345,N_1333,N_1385);
or U2346 (N_2346,N_1113,N_1513);
or U2347 (N_2347,N_1985,N_1179);
nand U2348 (N_2348,N_1288,N_1377);
xor U2349 (N_2349,N_1026,N_1998);
nand U2350 (N_2350,N_1045,N_1701);
nor U2351 (N_2351,N_1540,N_1098);
nor U2352 (N_2352,N_1868,N_1572);
or U2353 (N_2353,N_1470,N_1757);
or U2354 (N_2354,N_1265,N_1966);
nor U2355 (N_2355,N_1125,N_1166);
and U2356 (N_2356,N_1656,N_1609);
and U2357 (N_2357,N_1691,N_1509);
or U2358 (N_2358,N_1282,N_1822);
nor U2359 (N_2359,N_1659,N_1927);
nor U2360 (N_2360,N_1134,N_1939);
and U2361 (N_2361,N_1132,N_1160);
xnor U2362 (N_2362,N_1071,N_1856);
nor U2363 (N_2363,N_1899,N_1447);
and U2364 (N_2364,N_1186,N_1213);
nand U2365 (N_2365,N_1989,N_1253);
nor U2366 (N_2366,N_1488,N_1919);
and U2367 (N_2367,N_1056,N_1741);
nor U2368 (N_2368,N_1886,N_1551);
xor U2369 (N_2369,N_1199,N_1716);
and U2370 (N_2370,N_1351,N_1157);
xnor U2371 (N_2371,N_1718,N_1133);
or U2372 (N_2372,N_1223,N_1892);
nand U2373 (N_2373,N_1309,N_1722);
xnor U2374 (N_2374,N_1303,N_1666);
and U2375 (N_2375,N_1407,N_1106);
and U2376 (N_2376,N_1480,N_1582);
nand U2377 (N_2377,N_1468,N_1642);
nand U2378 (N_2378,N_1936,N_1622);
or U2379 (N_2379,N_1532,N_1782);
nand U2380 (N_2380,N_1369,N_1263);
nor U2381 (N_2381,N_1118,N_1047);
or U2382 (N_2382,N_1411,N_1990);
nor U2383 (N_2383,N_1331,N_1104);
and U2384 (N_2384,N_1754,N_1277);
nand U2385 (N_2385,N_1893,N_1776);
nand U2386 (N_2386,N_1745,N_1294);
and U2387 (N_2387,N_1763,N_1006);
nand U2388 (N_2388,N_1795,N_1600);
and U2389 (N_2389,N_1372,N_1872);
nand U2390 (N_2390,N_1446,N_1831);
nor U2391 (N_2391,N_1746,N_1577);
and U2392 (N_2392,N_1018,N_1729);
and U2393 (N_2393,N_1496,N_1243);
nand U2394 (N_2394,N_1848,N_1774);
nand U2395 (N_2395,N_1707,N_1027);
nand U2396 (N_2396,N_1742,N_1773);
and U2397 (N_2397,N_1299,N_1384);
or U2398 (N_2398,N_1533,N_1503);
and U2399 (N_2399,N_1850,N_1824);
xnor U2400 (N_2400,N_1346,N_1387);
nand U2401 (N_2401,N_1764,N_1548);
or U2402 (N_2402,N_1612,N_1237);
nand U2403 (N_2403,N_1857,N_1375);
nor U2404 (N_2404,N_1373,N_1475);
or U2405 (N_2405,N_1040,N_1012);
xnor U2406 (N_2406,N_1039,N_1524);
nor U2407 (N_2407,N_1301,N_1247);
nor U2408 (N_2408,N_1183,N_1556);
nor U2409 (N_2409,N_1905,N_1246);
nand U2410 (N_2410,N_1093,N_1107);
or U2411 (N_2411,N_1653,N_1434);
xor U2412 (N_2412,N_1817,N_1365);
nor U2413 (N_2413,N_1456,N_1898);
nand U2414 (N_2414,N_1778,N_1258);
and U2415 (N_2415,N_1515,N_1684);
xnor U2416 (N_2416,N_1591,N_1731);
and U2417 (N_2417,N_1931,N_1011);
xor U2418 (N_2418,N_1010,N_1035);
nor U2419 (N_2419,N_1070,N_1730);
and U2420 (N_2420,N_1728,N_1584);
and U2421 (N_2421,N_1804,N_1900);
nand U2422 (N_2422,N_1163,N_1328);
nor U2423 (N_2423,N_1592,N_1988);
nor U2424 (N_2424,N_1298,N_1117);
nor U2425 (N_2425,N_1767,N_1202);
nand U2426 (N_2426,N_1280,N_1603);
nor U2427 (N_2427,N_1102,N_1291);
nor U2428 (N_2428,N_1891,N_1274);
nand U2429 (N_2429,N_1295,N_1708);
and U2430 (N_2430,N_1051,N_1959);
or U2431 (N_2431,N_1065,N_1486);
nand U2432 (N_2432,N_1566,N_1828);
nand U2433 (N_2433,N_1948,N_1119);
or U2434 (N_2434,N_1637,N_1619);
nand U2435 (N_2435,N_1827,N_1392);
xor U2436 (N_2436,N_1586,N_1089);
xor U2437 (N_2437,N_1747,N_1732);
nand U2438 (N_2438,N_1968,N_1699);
and U2439 (N_2439,N_1836,N_1204);
nand U2440 (N_2440,N_1639,N_1200);
nor U2441 (N_2441,N_1606,N_1086);
nand U2442 (N_2442,N_1428,N_1379);
nor U2443 (N_2443,N_1063,N_1498);
or U2444 (N_2444,N_1059,N_1304);
nor U2445 (N_2445,N_1860,N_1105);
or U2446 (N_2446,N_1341,N_1169);
and U2447 (N_2447,N_1820,N_1410);
nand U2448 (N_2448,N_1193,N_1734);
nand U2449 (N_2449,N_1197,N_1419);
or U2450 (N_2450,N_1997,N_1799);
or U2451 (N_2451,N_1976,N_1511);
and U2452 (N_2452,N_1909,N_1257);
nor U2453 (N_2453,N_1964,N_1644);
nor U2454 (N_2454,N_1980,N_1885);
or U2455 (N_2455,N_1652,N_1580);
nor U2456 (N_2456,N_1194,N_1589);
or U2457 (N_2457,N_1620,N_1491);
and U2458 (N_2458,N_1422,N_1033);
nand U2459 (N_2459,N_1791,N_1329);
or U2460 (N_2460,N_1801,N_1073);
or U2461 (N_2461,N_1863,N_1423);
nor U2462 (N_2462,N_1150,N_1835);
or U2463 (N_2463,N_1766,N_1161);
and U2464 (N_2464,N_1210,N_1926);
xor U2465 (N_2465,N_1676,N_1207);
nor U2466 (N_2466,N_1573,N_1198);
or U2467 (N_2467,N_1452,N_1126);
and U2468 (N_2468,N_1136,N_1903);
and U2469 (N_2469,N_1130,N_1662);
nand U2470 (N_2470,N_1156,N_1627);
nand U2471 (N_2471,N_1983,N_1658);
and U2472 (N_2472,N_1719,N_1174);
nor U2473 (N_2473,N_1430,N_1583);
nor U2474 (N_2474,N_1195,N_1374);
nand U2475 (N_2475,N_1344,N_1472);
or U2476 (N_2476,N_1650,N_1981);
and U2477 (N_2477,N_1050,N_1852);
and U2478 (N_2478,N_1087,N_1703);
and U2479 (N_2479,N_1149,N_1031);
xor U2480 (N_2480,N_1000,N_1181);
and U2481 (N_2481,N_1054,N_1321);
nor U2482 (N_2482,N_1064,N_1267);
nand U2483 (N_2483,N_1465,N_1999);
nor U2484 (N_2484,N_1561,N_1217);
or U2485 (N_2485,N_1418,N_1185);
nor U2486 (N_2486,N_1284,N_1807);
nor U2487 (N_2487,N_1636,N_1651);
and U2488 (N_2488,N_1960,N_1904);
or U2489 (N_2489,N_1944,N_1674);
or U2490 (N_2490,N_1477,N_1077);
and U2491 (N_2491,N_1678,N_1016);
xnor U2492 (N_2492,N_1414,N_1450);
nor U2493 (N_2493,N_1815,N_1563);
or U2494 (N_2494,N_1023,N_1539);
nand U2495 (N_2495,N_1907,N_1066);
xor U2496 (N_2496,N_1564,N_1190);
or U2497 (N_2497,N_1415,N_1599);
or U2498 (N_2498,N_1569,N_1254);
nor U2499 (N_2499,N_1961,N_1203);
and U2500 (N_2500,N_1162,N_1025);
xor U2501 (N_2501,N_1532,N_1296);
nor U2502 (N_2502,N_1034,N_1281);
or U2503 (N_2503,N_1823,N_1231);
or U2504 (N_2504,N_1242,N_1820);
nor U2505 (N_2505,N_1957,N_1318);
and U2506 (N_2506,N_1587,N_1398);
nor U2507 (N_2507,N_1387,N_1949);
and U2508 (N_2508,N_1359,N_1978);
and U2509 (N_2509,N_1368,N_1611);
nor U2510 (N_2510,N_1472,N_1636);
or U2511 (N_2511,N_1118,N_1574);
or U2512 (N_2512,N_1012,N_1257);
nor U2513 (N_2513,N_1721,N_1651);
and U2514 (N_2514,N_1674,N_1832);
nor U2515 (N_2515,N_1769,N_1790);
nor U2516 (N_2516,N_1735,N_1262);
nor U2517 (N_2517,N_1300,N_1571);
or U2518 (N_2518,N_1165,N_1423);
nor U2519 (N_2519,N_1092,N_1956);
nor U2520 (N_2520,N_1952,N_1098);
or U2521 (N_2521,N_1554,N_1897);
nand U2522 (N_2522,N_1635,N_1135);
or U2523 (N_2523,N_1663,N_1526);
xor U2524 (N_2524,N_1886,N_1841);
and U2525 (N_2525,N_1024,N_1153);
xnor U2526 (N_2526,N_1183,N_1855);
nand U2527 (N_2527,N_1912,N_1806);
xnor U2528 (N_2528,N_1343,N_1568);
and U2529 (N_2529,N_1572,N_1257);
xor U2530 (N_2530,N_1655,N_1407);
nand U2531 (N_2531,N_1717,N_1276);
and U2532 (N_2532,N_1550,N_1281);
and U2533 (N_2533,N_1370,N_1126);
or U2534 (N_2534,N_1417,N_1431);
and U2535 (N_2535,N_1013,N_1862);
nor U2536 (N_2536,N_1466,N_1373);
nand U2537 (N_2537,N_1190,N_1131);
or U2538 (N_2538,N_1513,N_1246);
and U2539 (N_2539,N_1390,N_1423);
nor U2540 (N_2540,N_1770,N_1163);
xor U2541 (N_2541,N_1468,N_1572);
nand U2542 (N_2542,N_1356,N_1288);
or U2543 (N_2543,N_1083,N_1232);
xor U2544 (N_2544,N_1247,N_1499);
xnor U2545 (N_2545,N_1669,N_1988);
nand U2546 (N_2546,N_1623,N_1741);
or U2547 (N_2547,N_1075,N_1506);
and U2548 (N_2548,N_1789,N_1689);
nand U2549 (N_2549,N_1615,N_1691);
and U2550 (N_2550,N_1546,N_1992);
xor U2551 (N_2551,N_1469,N_1872);
nor U2552 (N_2552,N_1776,N_1829);
nor U2553 (N_2553,N_1486,N_1115);
or U2554 (N_2554,N_1459,N_1445);
nand U2555 (N_2555,N_1612,N_1574);
nor U2556 (N_2556,N_1402,N_1182);
nor U2557 (N_2557,N_1849,N_1398);
and U2558 (N_2558,N_1252,N_1572);
nand U2559 (N_2559,N_1137,N_1853);
nand U2560 (N_2560,N_1234,N_1129);
nand U2561 (N_2561,N_1108,N_1837);
or U2562 (N_2562,N_1369,N_1386);
nor U2563 (N_2563,N_1612,N_1183);
nand U2564 (N_2564,N_1332,N_1607);
or U2565 (N_2565,N_1681,N_1057);
or U2566 (N_2566,N_1749,N_1180);
and U2567 (N_2567,N_1889,N_1950);
and U2568 (N_2568,N_1909,N_1356);
or U2569 (N_2569,N_1945,N_1163);
nand U2570 (N_2570,N_1123,N_1355);
nand U2571 (N_2571,N_1791,N_1221);
or U2572 (N_2572,N_1180,N_1914);
nand U2573 (N_2573,N_1939,N_1283);
and U2574 (N_2574,N_1560,N_1055);
nand U2575 (N_2575,N_1434,N_1760);
and U2576 (N_2576,N_1230,N_1354);
nor U2577 (N_2577,N_1096,N_1522);
nor U2578 (N_2578,N_1966,N_1773);
or U2579 (N_2579,N_1671,N_1575);
or U2580 (N_2580,N_1441,N_1963);
nor U2581 (N_2581,N_1210,N_1200);
or U2582 (N_2582,N_1020,N_1803);
and U2583 (N_2583,N_1117,N_1811);
nor U2584 (N_2584,N_1511,N_1182);
or U2585 (N_2585,N_1170,N_1494);
and U2586 (N_2586,N_1249,N_1274);
nor U2587 (N_2587,N_1096,N_1455);
xor U2588 (N_2588,N_1798,N_1373);
or U2589 (N_2589,N_1675,N_1390);
nor U2590 (N_2590,N_1566,N_1577);
and U2591 (N_2591,N_1880,N_1566);
or U2592 (N_2592,N_1805,N_1702);
or U2593 (N_2593,N_1941,N_1534);
or U2594 (N_2594,N_1939,N_1494);
nor U2595 (N_2595,N_1608,N_1637);
nand U2596 (N_2596,N_1781,N_1767);
and U2597 (N_2597,N_1097,N_1044);
nor U2598 (N_2598,N_1087,N_1935);
nand U2599 (N_2599,N_1122,N_1957);
nand U2600 (N_2600,N_1564,N_1393);
xnor U2601 (N_2601,N_1225,N_1753);
xnor U2602 (N_2602,N_1998,N_1810);
nand U2603 (N_2603,N_1356,N_1262);
or U2604 (N_2604,N_1570,N_1252);
nand U2605 (N_2605,N_1539,N_1767);
or U2606 (N_2606,N_1033,N_1359);
nand U2607 (N_2607,N_1749,N_1891);
and U2608 (N_2608,N_1960,N_1517);
nor U2609 (N_2609,N_1310,N_1421);
and U2610 (N_2610,N_1412,N_1512);
or U2611 (N_2611,N_1642,N_1021);
or U2612 (N_2612,N_1340,N_1430);
or U2613 (N_2613,N_1466,N_1904);
nor U2614 (N_2614,N_1355,N_1804);
and U2615 (N_2615,N_1435,N_1533);
or U2616 (N_2616,N_1944,N_1191);
nor U2617 (N_2617,N_1302,N_1732);
or U2618 (N_2618,N_1664,N_1708);
and U2619 (N_2619,N_1051,N_1768);
and U2620 (N_2620,N_1079,N_1223);
or U2621 (N_2621,N_1219,N_1531);
and U2622 (N_2622,N_1224,N_1659);
nand U2623 (N_2623,N_1858,N_1924);
and U2624 (N_2624,N_1799,N_1687);
and U2625 (N_2625,N_1201,N_1387);
nor U2626 (N_2626,N_1846,N_1122);
nand U2627 (N_2627,N_1147,N_1771);
or U2628 (N_2628,N_1819,N_1711);
nand U2629 (N_2629,N_1802,N_1904);
nand U2630 (N_2630,N_1361,N_1005);
or U2631 (N_2631,N_1037,N_1401);
nor U2632 (N_2632,N_1070,N_1540);
xnor U2633 (N_2633,N_1082,N_1074);
or U2634 (N_2634,N_1563,N_1687);
xor U2635 (N_2635,N_1785,N_1425);
nand U2636 (N_2636,N_1948,N_1894);
and U2637 (N_2637,N_1231,N_1892);
or U2638 (N_2638,N_1739,N_1837);
and U2639 (N_2639,N_1785,N_1056);
and U2640 (N_2640,N_1726,N_1245);
and U2641 (N_2641,N_1440,N_1760);
nand U2642 (N_2642,N_1307,N_1243);
xnor U2643 (N_2643,N_1783,N_1765);
or U2644 (N_2644,N_1651,N_1446);
nand U2645 (N_2645,N_1488,N_1816);
or U2646 (N_2646,N_1491,N_1456);
or U2647 (N_2647,N_1417,N_1723);
nor U2648 (N_2648,N_1171,N_1451);
or U2649 (N_2649,N_1835,N_1284);
nor U2650 (N_2650,N_1979,N_1300);
nand U2651 (N_2651,N_1517,N_1154);
nand U2652 (N_2652,N_1839,N_1339);
or U2653 (N_2653,N_1381,N_1729);
xnor U2654 (N_2654,N_1181,N_1515);
nand U2655 (N_2655,N_1611,N_1487);
and U2656 (N_2656,N_1060,N_1562);
nand U2657 (N_2657,N_1619,N_1612);
xor U2658 (N_2658,N_1976,N_1723);
xnor U2659 (N_2659,N_1824,N_1375);
or U2660 (N_2660,N_1229,N_1993);
nand U2661 (N_2661,N_1635,N_1698);
nand U2662 (N_2662,N_1234,N_1569);
or U2663 (N_2663,N_1225,N_1713);
and U2664 (N_2664,N_1775,N_1317);
or U2665 (N_2665,N_1394,N_1038);
nor U2666 (N_2666,N_1989,N_1136);
and U2667 (N_2667,N_1560,N_1602);
nor U2668 (N_2668,N_1429,N_1597);
xor U2669 (N_2669,N_1448,N_1907);
or U2670 (N_2670,N_1465,N_1059);
nor U2671 (N_2671,N_1988,N_1063);
or U2672 (N_2672,N_1709,N_1550);
and U2673 (N_2673,N_1470,N_1553);
and U2674 (N_2674,N_1578,N_1090);
nor U2675 (N_2675,N_1635,N_1122);
and U2676 (N_2676,N_1323,N_1441);
and U2677 (N_2677,N_1091,N_1743);
or U2678 (N_2678,N_1004,N_1332);
and U2679 (N_2679,N_1430,N_1664);
nand U2680 (N_2680,N_1591,N_1509);
and U2681 (N_2681,N_1965,N_1990);
nor U2682 (N_2682,N_1548,N_1948);
nand U2683 (N_2683,N_1763,N_1689);
nand U2684 (N_2684,N_1845,N_1703);
xor U2685 (N_2685,N_1824,N_1184);
nor U2686 (N_2686,N_1442,N_1885);
and U2687 (N_2687,N_1684,N_1359);
nand U2688 (N_2688,N_1015,N_1554);
or U2689 (N_2689,N_1039,N_1178);
or U2690 (N_2690,N_1424,N_1860);
or U2691 (N_2691,N_1311,N_1328);
nor U2692 (N_2692,N_1061,N_1129);
and U2693 (N_2693,N_1039,N_1047);
or U2694 (N_2694,N_1333,N_1097);
or U2695 (N_2695,N_1111,N_1083);
nor U2696 (N_2696,N_1699,N_1959);
and U2697 (N_2697,N_1509,N_1150);
nor U2698 (N_2698,N_1604,N_1866);
or U2699 (N_2699,N_1416,N_1373);
and U2700 (N_2700,N_1095,N_1358);
or U2701 (N_2701,N_1857,N_1927);
or U2702 (N_2702,N_1677,N_1899);
and U2703 (N_2703,N_1155,N_1072);
and U2704 (N_2704,N_1743,N_1461);
and U2705 (N_2705,N_1637,N_1520);
or U2706 (N_2706,N_1246,N_1356);
nor U2707 (N_2707,N_1563,N_1705);
or U2708 (N_2708,N_1917,N_1555);
or U2709 (N_2709,N_1368,N_1892);
or U2710 (N_2710,N_1690,N_1419);
nor U2711 (N_2711,N_1958,N_1702);
and U2712 (N_2712,N_1585,N_1661);
nor U2713 (N_2713,N_1691,N_1566);
nand U2714 (N_2714,N_1704,N_1466);
nand U2715 (N_2715,N_1332,N_1673);
nand U2716 (N_2716,N_1323,N_1216);
nand U2717 (N_2717,N_1375,N_1671);
or U2718 (N_2718,N_1655,N_1632);
nand U2719 (N_2719,N_1366,N_1114);
or U2720 (N_2720,N_1104,N_1427);
or U2721 (N_2721,N_1595,N_1020);
nor U2722 (N_2722,N_1184,N_1677);
nor U2723 (N_2723,N_1504,N_1929);
and U2724 (N_2724,N_1938,N_1238);
nor U2725 (N_2725,N_1156,N_1310);
or U2726 (N_2726,N_1230,N_1155);
or U2727 (N_2727,N_1813,N_1732);
nor U2728 (N_2728,N_1290,N_1631);
or U2729 (N_2729,N_1357,N_1496);
nor U2730 (N_2730,N_1485,N_1871);
and U2731 (N_2731,N_1665,N_1501);
nor U2732 (N_2732,N_1415,N_1817);
xor U2733 (N_2733,N_1615,N_1066);
or U2734 (N_2734,N_1308,N_1579);
nor U2735 (N_2735,N_1084,N_1653);
and U2736 (N_2736,N_1290,N_1487);
or U2737 (N_2737,N_1897,N_1390);
or U2738 (N_2738,N_1628,N_1495);
or U2739 (N_2739,N_1405,N_1574);
nand U2740 (N_2740,N_1711,N_1089);
and U2741 (N_2741,N_1303,N_1558);
nand U2742 (N_2742,N_1274,N_1750);
and U2743 (N_2743,N_1565,N_1855);
nor U2744 (N_2744,N_1535,N_1097);
and U2745 (N_2745,N_1748,N_1269);
and U2746 (N_2746,N_1478,N_1352);
nand U2747 (N_2747,N_1094,N_1893);
or U2748 (N_2748,N_1537,N_1870);
xnor U2749 (N_2749,N_1894,N_1990);
nor U2750 (N_2750,N_1781,N_1442);
xnor U2751 (N_2751,N_1315,N_1238);
nand U2752 (N_2752,N_1696,N_1600);
and U2753 (N_2753,N_1465,N_1508);
or U2754 (N_2754,N_1747,N_1355);
or U2755 (N_2755,N_1103,N_1509);
nand U2756 (N_2756,N_1201,N_1004);
nor U2757 (N_2757,N_1536,N_1576);
nor U2758 (N_2758,N_1039,N_1966);
nor U2759 (N_2759,N_1352,N_1883);
nand U2760 (N_2760,N_1079,N_1191);
or U2761 (N_2761,N_1642,N_1909);
and U2762 (N_2762,N_1902,N_1078);
nor U2763 (N_2763,N_1251,N_1509);
nor U2764 (N_2764,N_1573,N_1342);
xor U2765 (N_2765,N_1769,N_1892);
nor U2766 (N_2766,N_1287,N_1500);
nor U2767 (N_2767,N_1271,N_1457);
nor U2768 (N_2768,N_1398,N_1500);
nand U2769 (N_2769,N_1816,N_1371);
and U2770 (N_2770,N_1541,N_1641);
nor U2771 (N_2771,N_1202,N_1813);
xor U2772 (N_2772,N_1260,N_1707);
and U2773 (N_2773,N_1928,N_1119);
nand U2774 (N_2774,N_1699,N_1375);
nand U2775 (N_2775,N_1175,N_1698);
nor U2776 (N_2776,N_1054,N_1705);
nor U2777 (N_2777,N_1992,N_1618);
nand U2778 (N_2778,N_1501,N_1221);
nand U2779 (N_2779,N_1477,N_1640);
or U2780 (N_2780,N_1391,N_1871);
or U2781 (N_2781,N_1268,N_1310);
xor U2782 (N_2782,N_1293,N_1292);
nand U2783 (N_2783,N_1394,N_1757);
and U2784 (N_2784,N_1467,N_1606);
and U2785 (N_2785,N_1006,N_1124);
and U2786 (N_2786,N_1160,N_1834);
or U2787 (N_2787,N_1790,N_1841);
nand U2788 (N_2788,N_1548,N_1632);
nor U2789 (N_2789,N_1408,N_1509);
xnor U2790 (N_2790,N_1474,N_1133);
nor U2791 (N_2791,N_1175,N_1495);
nor U2792 (N_2792,N_1724,N_1580);
nor U2793 (N_2793,N_1277,N_1304);
and U2794 (N_2794,N_1033,N_1361);
and U2795 (N_2795,N_1760,N_1483);
or U2796 (N_2796,N_1447,N_1880);
nand U2797 (N_2797,N_1272,N_1366);
and U2798 (N_2798,N_1364,N_1203);
nand U2799 (N_2799,N_1331,N_1621);
nor U2800 (N_2800,N_1479,N_1288);
nand U2801 (N_2801,N_1551,N_1188);
and U2802 (N_2802,N_1428,N_1073);
nand U2803 (N_2803,N_1110,N_1535);
xnor U2804 (N_2804,N_1572,N_1674);
or U2805 (N_2805,N_1659,N_1525);
and U2806 (N_2806,N_1710,N_1099);
or U2807 (N_2807,N_1374,N_1193);
nand U2808 (N_2808,N_1235,N_1452);
and U2809 (N_2809,N_1791,N_1059);
nor U2810 (N_2810,N_1158,N_1389);
nor U2811 (N_2811,N_1706,N_1786);
and U2812 (N_2812,N_1500,N_1966);
or U2813 (N_2813,N_1326,N_1173);
and U2814 (N_2814,N_1642,N_1864);
or U2815 (N_2815,N_1984,N_1493);
and U2816 (N_2816,N_1034,N_1800);
nor U2817 (N_2817,N_1077,N_1311);
and U2818 (N_2818,N_1258,N_1093);
nor U2819 (N_2819,N_1024,N_1999);
xnor U2820 (N_2820,N_1482,N_1919);
xnor U2821 (N_2821,N_1180,N_1776);
or U2822 (N_2822,N_1509,N_1320);
nand U2823 (N_2823,N_1415,N_1589);
or U2824 (N_2824,N_1136,N_1128);
nor U2825 (N_2825,N_1480,N_1813);
or U2826 (N_2826,N_1109,N_1543);
nor U2827 (N_2827,N_1409,N_1724);
and U2828 (N_2828,N_1444,N_1387);
or U2829 (N_2829,N_1664,N_1301);
or U2830 (N_2830,N_1138,N_1699);
or U2831 (N_2831,N_1464,N_1081);
and U2832 (N_2832,N_1272,N_1782);
nand U2833 (N_2833,N_1438,N_1506);
and U2834 (N_2834,N_1691,N_1037);
and U2835 (N_2835,N_1264,N_1796);
nor U2836 (N_2836,N_1149,N_1451);
or U2837 (N_2837,N_1517,N_1122);
nor U2838 (N_2838,N_1763,N_1408);
nand U2839 (N_2839,N_1500,N_1636);
nand U2840 (N_2840,N_1757,N_1363);
nand U2841 (N_2841,N_1179,N_1940);
nor U2842 (N_2842,N_1695,N_1623);
nor U2843 (N_2843,N_1146,N_1027);
nor U2844 (N_2844,N_1570,N_1212);
nand U2845 (N_2845,N_1776,N_1258);
nor U2846 (N_2846,N_1611,N_1919);
or U2847 (N_2847,N_1987,N_1523);
nor U2848 (N_2848,N_1781,N_1416);
and U2849 (N_2849,N_1080,N_1607);
nor U2850 (N_2850,N_1762,N_1664);
nor U2851 (N_2851,N_1314,N_1725);
nand U2852 (N_2852,N_1383,N_1146);
nand U2853 (N_2853,N_1663,N_1738);
nand U2854 (N_2854,N_1894,N_1253);
and U2855 (N_2855,N_1520,N_1236);
nand U2856 (N_2856,N_1348,N_1090);
or U2857 (N_2857,N_1249,N_1892);
xnor U2858 (N_2858,N_1243,N_1148);
nand U2859 (N_2859,N_1743,N_1654);
nor U2860 (N_2860,N_1905,N_1038);
nor U2861 (N_2861,N_1778,N_1330);
nor U2862 (N_2862,N_1366,N_1894);
and U2863 (N_2863,N_1753,N_1718);
and U2864 (N_2864,N_1686,N_1700);
or U2865 (N_2865,N_1451,N_1586);
nor U2866 (N_2866,N_1732,N_1750);
or U2867 (N_2867,N_1319,N_1349);
and U2868 (N_2868,N_1802,N_1995);
nor U2869 (N_2869,N_1363,N_1141);
or U2870 (N_2870,N_1731,N_1982);
nand U2871 (N_2871,N_1352,N_1096);
nor U2872 (N_2872,N_1629,N_1639);
and U2873 (N_2873,N_1560,N_1811);
nand U2874 (N_2874,N_1590,N_1085);
and U2875 (N_2875,N_1148,N_1824);
nor U2876 (N_2876,N_1657,N_1971);
or U2877 (N_2877,N_1220,N_1748);
nor U2878 (N_2878,N_1493,N_1332);
and U2879 (N_2879,N_1385,N_1683);
and U2880 (N_2880,N_1086,N_1533);
or U2881 (N_2881,N_1171,N_1665);
xor U2882 (N_2882,N_1440,N_1651);
xnor U2883 (N_2883,N_1371,N_1570);
or U2884 (N_2884,N_1289,N_1669);
and U2885 (N_2885,N_1632,N_1139);
and U2886 (N_2886,N_1513,N_1674);
nand U2887 (N_2887,N_1399,N_1056);
nand U2888 (N_2888,N_1590,N_1214);
and U2889 (N_2889,N_1771,N_1611);
nand U2890 (N_2890,N_1635,N_1717);
and U2891 (N_2891,N_1582,N_1253);
and U2892 (N_2892,N_1315,N_1739);
xnor U2893 (N_2893,N_1813,N_1898);
or U2894 (N_2894,N_1165,N_1453);
and U2895 (N_2895,N_1563,N_1467);
nand U2896 (N_2896,N_1642,N_1831);
xnor U2897 (N_2897,N_1830,N_1386);
nand U2898 (N_2898,N_1423,N_1777);
nor U2899 (N_2899,N_1916,N_1944);
or U2900 (N_2900,N_1880,N_1464);
nor U2901 (N_2901,N_1957,N_1857);
nor U2902 (N_2902,N_1621,N_1556);
nand U2903 (N_2903,N_1642,N_1160);
nand U2904 (N_2904,N_1794,N_1171);
or U2905 (N_2905,N_1117,N_1587);
nand U2906 (N_2906,N_1615,N_1583);
and U2907 (N_2907,N_1791,N_1353);
and U2908 (N_2908,N_1738,N_1846);
or U2909 (N_2909,N_1915,N_1745);
nand U2910 (N_2910,N_1594,N_1543);
nand U2911 (N_2911,N_1360,N_1757);
and U2912 (N_2912,N_1478,N_1308);
or U2913 (N_2913,N_1176,N_1951);
nand U2914 (N_2914,N_1783,N_1292);
or U2915 (N_2915,N_1454,N_1410);
or U2916 (N_2916,N_1100,N_1910);
or U2917 (N_2917,N_1934,N_1469);
or U2918 (N_2918,N_1357,N_1507);
or U2919 (N_2919,N_1063,N_1890);
and U2920 (N_2920,N_1589,N_1161);
nor U2921 (N_2921,N_1905,N_1371);
nor U2922 (N_2922,N_1333,N_1076);
nor U2923 (N_2923,N_1211,N_1585);
and U2924 (N_2924,N_1353,N_1005);
nor U2925 (N_2925,N_1075,N_1426);
and U2926 (N_2926,N_1742,N_1139);
nand U2927 (N_2927,N_1810,N_1407);
nand U2928 (N_2928,N_1918,N_1140);
or U2929 (N_2929,N_1734,N_1382);
nor U2930 (N_2930,N_1123,N_1070);
and U2931 (N_2931,N_1505,N_1167);
nand U2932 (N_2932,N_1226,N_1369);
and U2933 (N_2933,N_1730,N_1766);
or U2934 (N_2934,N_1156,N_1628);
and U2935 (N_2935,N_1761,N_1293);
nand U2936 (N_2936,N_1311,N_1441);
nor U2937 (N_2937,N_1487,N_1191);
nand U2938 (N_2938,N_1799,N_1456);
or U2939 (N_2939,N_1825,N_1996);
xor U2940 (N_2940,N_1073,N_1699);
xnor U2941 (N_2941,N_1455,N_1584);
nand U2942 (N_2942,N_1060,N_1595);
nor U2943 (N_2943,N_1607,N_1193);
xor U2944 (N_2944,N_1699,N_1597);
nand U2945 (N_2945,N_1807,N_1699);
or U2946 (N_2946,N_1569,N_1095);
or U2947 (N_2947,N_1368,N_1897);
or U2948 (N_2948,N_1840,N_1032);
or U2949 (N_2949,N_1983,N_1797);
or U2950 (N_2950,N_1815,N_1790);
or U2951 (N_2951,N_1633,N_1361);
nor U2952 (N_2952,N_1391,N_1170);
nor U2953 (N_2953,N_1067,N_1966);
nor U2954 (N_2954,N_1520,N_1603);
nand U2955 (N_2955,N_1341,N_1144);
and U2956 (N_2956,N_1076,N_1017);
nor U2957 (N_2957,N_1564,N_1412);
and U2958 (N_2958,N_1317,N_1305);
and U2959 (N_2959,N_1948,N_1685);
nand U2960 (N_2960,N_1028,N_1749);
or U2961 (N_2961,N_1138,N_1207);
nand U2962 (N_2962,N_1341,N_1505);
nor U2963 (N_2963,N_1673,N_1618);
or U2964 (N_2964,N_1627,N_1980);
nor U2965 (N_2965,N_1877,N_1444);
or U2966 (N_2966,N_1978,N_1850);
nor U2967 (N_2967,N_1157,N_1464);
nand U2968 (N_2968,N_1113,N_1142);
nand U2969 (N_2969,N_1446,N_1205);
nor U2970 (N_2970,N_1874,N_1323);
xnor U2971 (N_2971,N_1723,N_1969);
or U2972 (N_2972,N_1259,N_1430);
nand U2973 (N_2973,N_1461,N_1370);
nand U2974 (N_2974,N_1329,N_1088);
nor U2975 (N_2975,N_1606,N_1949);
nor U2976 (N_2976,N_1849,N_1930);
nand U2977 (N_2977,N_1953,N_1334);
xor U2978 (N_2978,N_1368,N_1404);
and U2979 (N_2979,N_1625,N_1618);
xnor U2980 (N_2980,N_1714,N_1870);
or U2981 (N_2981,N_1168,N_1056);
and U2982 (N_2982,N_1412,N_1706);
and U2983 (N_2983,N_1336,N_1973);
nor U2984 (N_2984,N_1827,N_1186);
nand U2985 (N_2985,N_1758,N_1886);
or U2986 (N_2986,N_1955,N_1950);
nand U2987 (N_2987,N_1091,N_1223);
nor U2988 (N_2988,N_1086,N_1335);
and U2989 (N_2989,N_1835,N_1450);
nor U2990 (N_2990,N_1988,N_1966);
nor U2991 (N_2991,N_1605,N_1706);
and U2992 (N_2992,N_1001,N_1672);
nor U2993 (N_2993,N_1742,N_1503);
xor U2994 (N_2994,N_1411,N_1172);
and U2995 (N_2995,N_1293,N_1194);
nor U2996 (N_2996,N_1038,N_1599);
xor U2997 (N_2997,N_1129,N_1898);
or U2998 (N_2998,N_1658,N_1376);
or U2999 (N_2999,N_1033,N_1383);
and U3000 (N_3000,N_2333,N_2340);
xnor U3001 (N_3001,N_2433,N_2204);
and U3002 (N_3002,N_2580,N_2299);
nand U3003 (N_3003,N_2217,N_2496);
or U3004 (N_3004,N_2110,N_2952);
nor U3005 (N_3005,N_2756,N_2783);
nand U3006 (N_3006,N_2965,N_2505);
nor U3007 (N_3007,N_2855,N_2524);
and U3008 (N_3008,N_2130,N_2193);
nor U3009 (N_3009,N_2406,N_2487);
nand U3010 (N_3010,N_2999,N_2611);
or U3011 (N_3011,N_2605,N_2891);
and U3012 (N_3012,N_2219,N_2454);
nor U3013 (N_3013,N_2561,N_2187);
nand U3014 (N_3014,N_2818,N_2283);
or U3015 (N_3015,N_2323,N_2362);
and U3016 (N_3016,N_2774,N_2922);
xnor U3017 (N_3017,N_2511,N_2736);
xnor U3018 (N_3018,N_2240,N_2490);
and U3019 (N_3019,N_2596,N_2215);
nand U3020 (N_3020,N_2290,N_2878);
or U3021 (N_3021,N_2152,N_2989);
nand U3022 (N_3022,N_2755,N_2390);
and U3023 (N_3023,N_2781,N_2024);
or U3024 (N_3024,N_2759,N_2932);
or U3025 (N_3025,N_2788,N_2334);
or U3026 (N_3026,N_2730,N_2654);
or U3027 (N_3027,N_2369,N_2313);
nand U3028 (N_3028,N_2363,N_2615);
xnor U3029 (N_3029,N_2548,N_2230);
or U3030 (N_3030,N_2728,N_2255);
or U3031 (N_3031,N_2798,N_2396);
nor U3032 (N_3032,N_2639,N_2311);
or U3033 (N_3033,N_2913,N_2695);
or U3034 (N_3034,N_2661,N_2448);
or U3035 (N_3035,N_2810,N_2655);
nand U3036 (N_3036,N_2321,N_2983);
nor U3037 (N_3037,N_2384,N_2974);
nor U3038 (N_3038,N_2813,N_2287);
or U3039 (N_3039,N_2149,N_2565);
and U3040 (N_3040,N_2468,N_2729);
nand U3041 (N_3041,N_2156,N_2610);
nand U3042 (N_3042,N_2971,N_2439);
nor U3043 (N_3043,N_2318,N_2038);
or U3044 (N_3044,N_2725,N_2459);
and U3045 (N_3045,N_2009,N_2282);
nor U3046 (N_3046,N_2638,N_2484);
and U3047 (N_3047,N_2183,N_2114);
nor U3048 (N_3048,N_2748,N_2811);
and U3049 (N_3049,N_2857,N_2420);
nor U3050 (N_3050,N_2234,N_2864);
nor U3051 (N_3051,N_2735,N_2395);
and U3052 (N_3052,N_2276,N_2249);
nand U3053 (N_3053,N_2049,N_2734);
nor U3054 (N_3054,N_2260,N_2348);
and U3055 (N_3055,N_2602,N_2414);
nor U3056 (N_3056,N_2645,N_2691);
nor U3057 (N_3057,N_2270,N_2520);
or U3058 (N_3058,N_2324,N_2224);
nand U3059 (N_3059,N_2918,N_2630);
and U3060 (N_3060,N_2707,N_2651);
nor U3061 (N_3061,N_2447,N_2048);
and U3062 (N_3062,N_2692,N_2238);
xnor U3063 (N_3063,N_2435,N_2591);
nand U3064 (N_3064,N_2208,N_2832);
or U3065 (N_3065,N_2241,N_2477);
nor U3066 (N_3066,N_2292,N_2214);
nand U3067 (N_3067,N_2417,N_2162);
nand U3068 (N_3068,N_2163,N_2557);
xor U3069 (N_3069,N_2760,N_2405);
and U3070 (N_3070,N_2688,N_2223);
nor U3071 (N_3071,N_2118,N_2476);
and U3072 (N_3072,N_2942,N_2551);
xor U3073 (N_3073,N_2198,N_2212);
and U3074 (N_3074,N_2455,N_2665);
or U3075 (N_3075,N_2286,N_2978);
or U3076 (N_3076,N_2745,N_2039);
and U3077 (N_3077,N_2573,N_2957);
and U3078 (N_3078,N_2350,N_2153);
nor U3079 (N_3079,N_2571,N_2155);
nand U3080 (N_3080,N_2002,N_2308);
and U3081 (N_3081,N_2806,N_2180);
or U3082 (N_3082,N_2034,N_2397);
nor U3083 (N_3083,N_2025,N_2101);
nand U3084 (N_3084,N_2257,N_2938);
or U3085 (N_3085,N_2947,N_2589);
nand U3086 (N_3086,N_2252,N_2139);
or U3087 (N_3087,N_2194,N_2841);
or U3088 (N_3088,N_2694,N_2815);
or U3089 (N_3089,N_2227,N_2124);
and U3090 (N_3090,N_2233,N_2457);
or U3091 (N_3091,N_2613,N_2222);
and U3092 (N_3092,N_2086,N_2686);
nor U3093 (N_3093,N_2393,N_2077);
nand U3094 (N_3094,N_2545,N_2320);
and U3095 (N_3095,N_2181,N_2663);
nor U3096 (N_3096,N_2933,N_2081);
nor U3097 (N_3097,N_2951,N_2840);
and U3098 (N_3098,N_2606,N_2154);
and U3099 (N_3099,N_2418,N_2791);
and U3100 (N_3100,N_2043,N_2868);
nor U3101 (N_3101,N_2880,N_2724);
nand U3102 (N_3102,N_2403,N_2342);
and U3103 (N_3103,N_2770,N_2738);
nand U3104 (N_3104,N_2078,N_2926);
and U3105 (N_3105,N_2923,N_2536);
nand U3106 (N_3106,N_2553,N_2068);
nand U3107 (N_3107,N_2570,N_2178);
nor U3108 (N_3108,N_2901,N_2629);
nor U3109 (N_3109,N_2102,N_2479);
nand U3110 (N_3110,N_2030,N_2205);
or U3111 (N_3111,N_2834,N_2460);
nand U3112 (N_3112,N_2528,N_2097);
nand U3113 (N_3113,N_2507,N_2305);
nor U3114 (N_3114,N_2055,N_2751);
nand U3115 (N_3115,N_2683,N_2035);
or U3116 (N_3116,N_2358,N_2601);
nor U3117 (N_3117,N_2415,N_2137);
or U3118 (N_3118,N_2191,N_2175);
nand U3119 (N_3119,N_2593,N_2157);
nor U3120 (N_3120,N_2353,N_2842);
or U3121 (N_3121,N_2091,N_2514);
xnor U3122 (N_3122,N_2005,N_2243);
nand U3123 (N_3123,N_2543,N_2731);
xor U3124 (N_3124,N_2170,N_2660);
or U3125 (N_3125,N_2560,N_2873);
nand U3126 (N_3126,N_2141,N_2753);
nor U3127 (N_3127,N_2497,N_2453);
nand U3128 (N_3128,N_2116,N_2014);
nor U3129 (N_3129,N_2885,N_2402);
or U3130 (N_3130,N_2295,N_2595);
or U3131 (N_3131,N_2360,N_2160);
and U3132 (N_3132,N_2517,N_2940);
nor U3133 (N_3133,N_2145,N_2177);
nand U3134 (N_3134,N_2858,N_2909);
nor U3135 (N_3135,N_2657,N_2888);
nand U3136 (N_3136,N_2159,N_2247);
nor U3137 (N_3137,N_2349,N_2833);
or U3138 (N_3138,N_2112,N_2277);
and U3139 (N_3139,N_2054,N_2166);
and U3140 (N_3140,N_2658,N_2000);
nand U3141 (N_3141,N_2341,N_2111);
xnor U3142 (N_3142,N_2310,N_2072);
or U3143 (N_3143,N_2019,N_2931);
nand U3144 (N_3144,N_2144,N_2196);
nor U3145 (N_3145,N_2003,N_2452);
nor U3146 (N_3146,N_2211,N_2343);
nor U3147 (N_3147,N_2192,N_2911);
nand U3148 (N_3148,N_2807,N_2047);
or U3149 (N_3149,N_2365,N_2073);
and U3150 (N_3150,N_2960,N_2328);
and U3151 (N_3151,N_2764,N_2887);
xnor U3152 (N_3152,N_2104,N_2347);
nor U3153 (N_3153,N_2702,N_2203);
and U3154 (N_3154,N_2377,N_2776);
nor U3155 (N_3155,N_2714,N_2797);
and U3156 (N_3156,N_2441,N_2622);
nand U3157 (N_3157,N_2673,N_2209);
nor U3158 (N_3158,N_2268,N_2248);
nor U3159 (N_3159,N_2837,N_2962);
nor U3160 (N_3160,N_2389,N_2977);
nor U3161 (N_3161,N_2905,N_2552);
or U3162 (N_3162,N_2941,N_2500);
xor U3163 (N_3163,N_2172,N_2325);
or U3164 (N_3164,N_2147,N_2699);
or U3165 (N_3165,N_2134,N_2850);
or U3166 (N_3166,N_2562,N_2555);
and U3167 (N_3167,N_2998,N_2317);
or U3168 (N_3168,N_2356,N_2188);
nor U3169 (N_3169,N_2762,N_2904);
and U3170 (N_3170,N_2994,N_2564);
nand U3171 (N_3171,N_2074,N_2142);
or U3172 (N_3172,N_2822,N_2438);
or U3173 (N_3173,N_2127,N_2096);
and U3174 (N_3174,N_2437,N_2509);
nor U3175 (N_3175,N_2012,N_2493);
nand U3176 (N_3176,N_2063,N_2411);
and U3177 (N_3177,N_2800,N_2330);
nand U3178 (N_3178,N_2794,N_2603);
xor U3179 (N_3179,N_2119,N_2006);
nand U3180 (N_3180,N_2523,N_2625);
nand U3181 (N_3181,N_2836,N_2817);
and U3182 (N_3182,N_2890,N_2632);
nand U3183 (N_3183,N_2371,N_2559);
nor U3184 (N_3184,N_2291,N_2863);
xor U3185 (N_3185,N_2083,N_2143);
nor U3186 (N_3186,N_2387,N_2768);
nand U3187 (N_3187,N_2620,N_2367);
nor U3188 (N_3188,N_2637,N_2823);
and U3189 (N_3189,N_2779,N_2169);
nor U3190 (N_3190,N_2424,N_2053);
or U3191 (N_3191,N_2279,N_2975);
nand U3192 (N_3192,N_2407,N_2567);
nand U3193 (N_3193,N_2264,N_2802);
nand U3194 (N_3194,N_2754,N_2984);
nand U3195 (N_3195,N_2314,N_2618);
and U3196 (N_3196,N_2251,N_2907);
or U3197 (N_3197,N_2769,N_2289);
nor U3198 (N_3198,N_2288,N_2865);
nand U3199 (N_3199,N_2973,N_2838);
and U3200 (N_3200,N_2261,N_2161);
nor U3201 (N_3201,N_2015,N_2094);
and U3202 (N_3202,N_2716,N_2004);
nor U3203 (N_3203,N_2210,N_2506);
nand U3204 (N_3204,N_2352,N_2385);
nand U3205 (N_3205,N_2700,N_2107);
nand U3206 (N_3206,N_2782,N_2828);
or U3207 (N_3207,N_2380,N_2711);
or U3208 (N_3208,N_2001,N_2016);
nand U3209 (N_3209,N_2515,N_2168);
or U3210 (N_3210,N_2540,N_2480);
and U3211 (N_3211,N_2098,N_2633);
or U3212 (N_3212,N_2426,N_2703);
nand U3213 (N_3213,N_2967,N_2920);
nand U3214 (N_3214,N_2258,N_2184);
or U3215 (N_3215,N_2451,N_2237);
or U3216 (N_3216,N_2848,N_2301);
xnor U3217 (N_3217,N_2586,N_2440);
nor U3218 (N_3218,N_2267,N_2747);
nand U3219 (N_3219,N_2988,N_2982);
nand U3220 (N_3220,N_2616,N_2554);
nand U3221 (N_3221,N_2943,N_2588);
or U3222 (N_3222,N_2895,N_2336);
or U3223 (N_3223,N_2445,N_2882);
and U3224 (N_3224,N_2599,N_2062);
or U3225 (N_3225,N_2067,N_2190);
or U3226 (N_3226,N_2950,N_2028);
nor U3227 (N_3227,N_2302,N_2082);
nand U3228 (N_3228,N_2372,N_2563);
nor U3229 (N_3229,N_2446,N_2976);
or U3230 (N_3230,N_2093,N_2835);
nor U3231 (N_3231,N_2912,N_2158);
or U3232 (N_3232,N_2547,N_2549);
or U3233 (N_3233,N_2337,N_2011);
nand U3234 (N_3234,N_2626,N_2100);
or U3235 (N_3235,N_2767,N_2641);
or U3236 (N_3236,N_2874,N_2737);
or U3237 (N_3237,N_2409,N_2359);
and U3238 (N_3238,N_2908,N_2609);
and U3239 (N_3239,N_2594,N_2659);
nand U3240 (N_3240,N_2566,N_2164);
or U3241 (N_3241,N_2787,N_2690);
nor U3242 (N_3242,N_2572,N_2539);
nor U3243 (N_3243,N_2766,N_2826);
nor U3244 (N_3244,N_2122,N_2262);
nand U3245 (N_3245,N_2478,N_2103);
nand U3246 (N_3246,N_2869,N_2274);
or U3247 (N_3247,N_2825,N_2176);
and U3248 (N_3248,N_2532,N_2743);
nor U3249 (N_3249,N_2600,N_2550);
or U3250 (N_3250,N_2051,N_2805);
xnor U3251 (N_3251,N_2167,N_2881);
nand U3252 (N_3252,N_2883,N_2579);
and U3253 (N_3253,N_2450,N_2546);
nor U3254 (N_3254,N_2023,N_2482);
nor U3255 (N_3255,N_2099,N_2085);
nor U3256 (N_3256,N_2354,N_2064);
and U3257 (N_3257,N_2758,N_2036);
xor U3258 (N_3258,N_2900,N_2293);
or U3259 (N_3259,N_2026,N_2309);
and U3260 (N_3260,N_2510,N_2542);
nand U3261 (N_3261,N_2682,N_2432);
nand U3262 (N_3262,N_2401,N_2374);
xor U3263 (N_3263,N_2990,N_2979);
or U3264 (N_3264,N_2698,N_2419);
nand U3265 (N_3265,N_2796,N_2461);
xor U3266 (N_3266,N_2079,N_2200);
nor U3267 (N_3267,N_2526,N_2525);
nand U3268 (N_3268,N_2467,N_2592);
or U3269 (N_3269,N_2568,N_2186);
nand U3270 (N_3270,N_2242,N_2919);
xnor U3271 (N_3271,N_2521,N_2117);
xor U3272 (N_3272,N_2648,N_2008);
and U3273 (N_3273,N_2392,N_2429);
nand U3274 (N_3274,N_2173,N_2533);
xnor U3275 (N_3275,N_2206,N_2899);
and U3276 (N_3276,N_2494,N_2430);
nor U3277 (N_3277,N_2884,N_2229);
nor U3278 (N_3278,N_2017,N_2705);
or U3279 (N_3279,N_2379,N_2558);
and U3280 (N_3280,N_2361,N_2772);
nor U3281 (N_3281,N_2031,N_2061);
or U3282 (N_3282,N_2236,N_2272);
and U3283 (N_3283,N_2959,N_2676);
and U3284 (N_3284,N_2582,N_2851);
nor U3285 (N_3285,N_2284,N_2860);
and U3286 (N_3286,N_2125,N_2421);
or U3287 (N_3287,N_2653,N_2803);
nand U3288 (N_3288,N_2980,N_2503);
nor U3289 (N_3289,N_2844,N_2488);
or U3290 (N_3290,N_2373,N_2351);
or U3291 (N_3291,N_2221,N_2627);
and U3292 (N_3292,N_2831,N_2256);
or U3293 (N_3293,N_2816,N_2076);
xnor U3294 (N_3294,N_2715,N_2778);
xnor U3295 (N_3295,N_2761,N_2721);
xnor U3296 (N_3296,N_2041,N_2875);
and U3297 (N_3297,N_2671,N_2642);
nand U3298 (N_3298,N_2140,N_2464);
nand U3299 (N_3299,N_2070,N_2171);
and U3300 (N_3300,N_2687,N_2033);
and U3301 (N_3301,N_2040,N_2133);
nand U3302 (N_3302,N_2696,N_2538);
nor U3303 (N_3303,N_2710,N_2502);
nand U3304 (N_3304,N_2329,N_2604);
nand U3305 (N_3305,N_2271,N_2677);
nor U3306 (N_3306,N_2801,N_2893);
or U3307 (N_3307,N_2966,N_2531);
or U3308 (N_3308,N_2646,N_2916);
or U3309 (N_3309,N_2213,N_2120);
nand U3310 (N_3310,N_2266,N_2216);
and U3311 (N_3311,N_2492,N_2644);
nand U3312 (N_3312,N_2150,N_2471);
nor U3313 (N_3313,N_2821,N_2956);
nor U3314 (N_3314,N_2253,N_2953);
or U3315 (N_3315,N_2332,N_2892);
nor U3316 (N_3316,N_2945,N_2013);
nor U3317 (N_3317,N_2534,N_2958);
xor U3318 (N_3318,N_2537,N_2583);
nor U3319 (N_3319,N_2667,N_2465);
or U3320 (N_3320,N_2631,N_2466);
or U3321 (N_3321,N_2335,N_2784);
nor U3322 (N_3322,N_2576,N_2856);
xnor U3323 (N_3323,N_2829,N_2719);
nor U3324 (N_3324,N_2643,N_2022);
or U3325 (N_3325,N_2723,N_2740);
nand U3326 (N_3326,N_2870,N_2458);
nand U3327 (N_3327,N_2244,N_2148);
or U3328 (N_3328,N_2556,N_2640);
nand U3329 (N_3329,N_2614,N_2628);
nor U3330 (N_3330,N_2634,N_2469);
nand U3331 (N_3331,N_2273,N_2578);
nor U3332 (N_3332,N_2339,N_2780);
or U3333 (N_3333,N_2199,N_2431);
nand U3334 (N_3334,N_2512,N_2220);
nor U3335 (N_3335,N_2704,N_2092);
nand U3336 (N_3336,N_2894,N_2027);
and U3337 (N_3337,N_2131,N_2095);
nor U3338 (N_3338,N_2297,N_2486);
nand U3339 (N_3339,N_2872,N_2058);
or U3340 (N_3340,N_2612,N_2044);
or U3341 (N_3341,N_2750,N_2886);
and U3342 (N_3342,N_2970,N_2852);
nor U3343 (N_3343,N_2434,N_2239);
nand U3344 (N_3344,N_2773,N_2535);
xor U3345 (N_3345,N_2914,N_2927);
nand U3346 (N_3346,N_2129,N_2059);
or U3347 (N_3347,N_2775,N_2830);
nand U3348 (N_3348,N_2410,N_2381);
nand U3349 (N_3349,N_2843,N_2896);
and U3350 (N_3350,N_2151,N_2992);
nor U3351 (N_3351,N_2281,N_2635);
nor U3352 (N_3352,N_2808,N_2935);
nor U3353 (N_3353,N_2697,N_2052);
and U3354 (N_3354,N_2518,N_2996);
nor U3355 (N_3355,N_2732,N_2386);
nor U3356 (N_3356,N_2189,N_2981);
or U3357 (N_3357,N_2793,N_2877);
or U3358 (N_3358,N_2060,N_2720);
nor U3359 (N_3359,N_2179,N_2944);
or U3360 (N_3360,N_2581,N_2777);
nand U3361 (N_3361,N_2809,N_2861);
or U3362 (N_3362,N_2814,N_2423);
and U3363 (N_3363,N_2057,N_2598);
nor U3364 (N_3364,N_2513,N_2394);
or U3365 (N_3365,N_2669,N_2444);
or U3366 (N_3366,N_2066,N_2527);
and U3367 (N_3367,N_2936,N_2785);
nand U3368 (N_3368,N_2544,N_2934);
or U3369 (N_3369,N_2495,N_2115);
and U3370 (N_3370,N_2121,N_2706);
nand U3371 (N_3371,N_2508,N_2463);
and U3372 (N_3372,N_2250,N_2853);
nand U3373 (N_3373,N_2991,N_2607);
nand U3374 (N_3374,N_2866,N_2427);
nand U3375 (N_3375,N_2278,N_2968);
or U3376 (N_3376,N_2742,N_2307);
or U3377 (N_3377,N_2300,N_2712);
or U3378 (N_3378,N_2929,N_2504);
and U3379 (N_3379,N_2235,N_2298);
or U3380 (N_3380,N_2498,N_2174);
and U3381 (N_3381,N_2416,N_2584);
or U3382 (N_3382,N_2889,N_2898);
and U3383 (N_3383,N_2069,N_2917);
or U3384 (N_3384,N_2915,N_2867);
nor U3385 (N_3385,N_2925,N_2846);
xor U3386 (N_3386,N_2485,N_2827);
or U3387 (N_3387,N_2961,N_2046);
or U3388 (N_3388,N_2790,N_2428);
and U3389 (N_3389,N_2042,N_2182);
nor U3390 (N_3390,N_2516,N_2819);
and U3391 (N_3391,N_2995,N_2408);
nand U3392 (N_3392,N_2792,N_2456);
or U3393 (N_3393,N_2226,N_2368);
nand U3394 (N_3394,N_2483,N_2871);
or U3395 (N_3395,N_2804,N_2799);
xor U3396 (N_3396,N_2263,N_2577);
and U3397 (N_3397,N_2949,N_2765);
and U3398 (N_3398,N_2443,N_2294);
and U3399 (N_3399,N_2327,N_2388);
and U3400 (N_3400,N_2338,N_2656);
nand U3401 (N_3401,N_2985,N_2664);
or U3402 (N_3402,N_2109,N_2201);
nand U3403 (N_3403,N_2954,N_2930);
nor U3404 (N_3404,N_2231,N_2075);
nand U3405 (N_3405,N_2436,N_2071);
and U3406 (N_3406,N_2621,N_2280);
and U3407 (N_3407,N_2364,N_2541);
nor U3408 (N_3408,N_2680,N_2128);
or U3409 (N_3409,N_2624,N_2963);
nor U3410 (N_3410,N_2202,N_2662);
nor U3411 (N_3411,N_2845,N_2106);
nor U3412 (N_3412,N_2259,N_2275);
nor U3413 (N_3413,N_2713,N_2474);
or U3414 (N_3414,N_2499,N_2399);
and U3415 (N_3415,N_2820,N_2400);
xor U3416 (N_3416,N_2897,N_2910);
nand U3417 (N_3417,N_2739,N_2032);
nor U3418 (N_3418,N_2597,N_2425);
nor U3419 (N_3419,N_2617,N_2123);
nor U3420 (N_3420,N_2587,N_2473);
and U3421 (N_3421,N_2376,N_2303);
nor U3422 (N_3422,N_2398,N_2529);
or U3423 (N_3423,N_2717,N_2470);
and U3424 (N_3424,N_2530,N_2197);
and U3425 (N_3425,N_2928,N_2679);
nor U3426 (N_3426,N_2246,N_2903);
or U3427 (N_3427,N_2489,N_2969);
nor U3428 (N_3428,N_2590,N_2746);
nor U3429 (N_3429,N_2413,N_2678);
or U3430 (N_3430,N_2007,N_2849);
and U3431 (N_3431,N_2757,N_2939);
and U3432 (N_3432,N_2685,N_2449);
nand U3433 (N_3433,N_2986,N_2859);
nor U3434 (N_3434,N_2113,N_2056);
and U3435 (N_3435,N_2304,N_2422);
or U3436 (N_3436,N_2647,N_2741);
or U3437 (N_3437,N_2225,N_2574);
nor U3438 (N_3438,N_2285,N_2650);
or U3439 (N_3439,N_2357,N_2331);
or U3440 (N_3440,N_2383,N_2854);
nor U3441 (N_3441,N_2050,N_2652);
and U3442 (N_3442,N_2708,N_2668);
and U3443 (N_3443,N_2136,N_2232);
nand U3444 (N_3444,N_2195,N_2087);
xnor U3445 (N_3445,N_2733,N_2404);
and U3446 (N_3446,N_2245,N_2619);
and U3447 (N_3447,N_2752,N_2839);
and U3448 (N_3448,N_2672,N_2824);
and U3449 (N_3449,N_2876,N_2472);
nor U3450 (N_3450,N_2020,N_2569);
or U3451 (N_3451,N_2375,N_2021);
nand U3452 (N_3452,N_2481,N_2987);
nor U3453 (N_3453,N_2089,N_2316);
or U3454 (N_3454,N_2378,N_2722);
nor U3455 (N_3455,N_2847,N_2366);
xor U3456 (N_3456,N_2649,N_2132);
nor U3457 (N_3457,N_2218,N_2675);
and U3458 (N_3458,N_2997,N_2090);
nor U3459 (N_3459,N_2344,N_2108);
and U3460 (N_3460,N_2522,N_2391);
nor U3461 (N_3461,N_2010,N_2906);
or U3462 (N_3462,N_2902,N_2269);
nor U3463 (N_3463,N_2585,N_2382);
or U3464 (N_3464,N_2322,N_2045);
and U3465 (N_3465,N_2955,N_2126);
nor U3466 (N_3466,N_2862,N_2519);
nor U3467 (N_3467,N_2972,N_2088);
nor U3468 (N_3468,N_2623,N_2674);
and U3469 (N_3469,N_2345,N_2146);
or U3470 (N_3470,N_2254,N_2771);
nor U3471 (N_3471,N_2789,N_2946);
or U3472 (N_3472,N_2105,N_2312);
nor U3473 (N_3473,N_2666,N_2185);
and U3474 (N_3474,N_2786,N_2744);
nor U3475 (N_3475,N_2749,N_2462);
or U3476 (N_3476,N_2681,N_2924);
nand U3477 (N_3477,N_2937,N_2763);
nor U3478 (N_3478,N_2475,N_2709);
and U3479 (N_3479,N_2306,N_2636);
xor U3480 (N_3480,N_2689,N_2207);
nand U3481 (N_3481,N_2412,N_2948);
or U3482 (N_3482,N_2135,N_2296);
nand U3483 (N_3483,N_2355,N_2265);
nor U3484 (N_3484,N_2080,N_2084);
nand U3485 (N_3485,N_2501,N_2491);
and U3486 (N_3486,N_2684,N_2346);
nor U3487 (N_3487,N_2037,N_2608);
nor U3488 (N_3488,N_2018,N_2921);
or U3489 (N_3489,N_2326,N_2993);
xnor U3490 (N_3490,N_2315,N_2718);
nor U3491 (N_3491,N_2575,N_2795);
or U3492 (N_3492,N_2228,N_2812);
or U3493 (N_3493,N_2701,N_2693);
xnor U3494 (N_3494,N_2065,N_2165);
and U3495 (N_3495,N_2442,N_2370);
nand U3496 (N_3496,N_2319,N_2727);
or U3497 (N_3497,N_2879,N_2964);
nand U3498 (N_3498,N_2670,N_2029);
or U3499 (N_3499,N_2138,N_2726);
and U3500 (N_3500,N_2333,N_2160);
or U3501 (N_3501,N_2073,N_2704);
nand U3502 (N_3502,N_2744,N_2223);
nor U3503 (N_3503,N_2309,N_2909);
nor U3504 (N_3504,N_2490,N_2533);
nand U3505 (N_3505,N_2119,N_2881);
nor U3506 (N_3506,N_2397,N_2872);
nand U3507 (N_3507,N_2849,N_2842);
nor U3508 (N_3508,N_2279,N_2177);
nor U3509 (N_3509,N_2029,N_2602);
nor U3510 (N_3510,N_2121,N_2259);
nand U3511 (N_3511,N_2928,N_2540);
nand U3512 (N_3512,N_2670,N_2147);
and U3513 (N_3513,N_2928,N_2189);
and U3514 (N_3514,N_2755,N_2571);
or U3515 (N_3515,N_2520,N_2089);
and U3516 (N_3516,N_2696,N_2609);
nand U3517 (N_3517,N_2828,N_2876);
and U3518 (N_3518,N_2795,N_2833);
or U3519 (N_3519,N_2051,N_2946);
nand U3520 (N_3520,N_2251,N_2531);
and U3521 (N_3521,N_2410,N_2271);
nand U3522 (N_3522,N_2034,N_2667);
and U3523 (N_3523,N_2058,N_2387);
xor U3524 (N_3524,N_2940,N_2867);
or U3525 (N_3525,N_2859,N_2553);
nand U3526 (N_3526,N_2398,N_2720);
xor U3527 (N_3527,N_2183,N_2225);
or U3528 (N_3528,N_2920,N_2375);
nor U3529 (N_3529,N_2876,N_2432);
nand U3530 (N_3530,N_2642,N_2576);
or U3531 (N_3531,N_2331,N_2912);
or U3532 (N_3532,N_2850,N_2208);
or U3533 (N_3533,N_2523,N_2522);
and U3534 (N_3534,N_2313,N_2408);
xnor U3535 (N_3535,N_2882,N_2818);
nor U3536 (N_3536,N_2044,N_2617);
nand U3537 (N_3537,N_2950,N_2965);
nor U3538 (N_3538,N_2760,N_2767);
nor U3539 (N_3539,N_2360,N_2158);
or U3540 (N_3540,N_2068,N_2471);
and U3541 (N_3541,N_2828,N_2619);
nand U3542 (N_3542,N_2505,N_2665);
or U3543 (N_3543,N_2581,N_2378);
and U3544 (N_3544,N_2823,N_2026);
and U3545 (N_3545,N_2304,N_2267);
or U3546 (N_3546,N_2949,N_2809);
or U3547 (N_3547,N_2460,N_2358);
and U3548 (N_3548,N_2189,N_2711);
or U3549 (N_3549,N_2504,N_2717);
xnor U3550 (N_3550,N_2921,N_2408);
nand U3551 (N_3551,N_2829,N_2388);
or U3552 (N_3552,N_2445,N_2999);
and U3553 (N_3553,N_2885,N_2771);
and U3554 (N_3554,N_2804,N_2249);
nor U3555 (N_3555,N_2339,N_2316);
nand U3556 (N_3556,N_2803,N_2446);
nor U3557 (N_3557,N_2067,N_2668);
or U3558 (N_3558,N_2284,N_2345);
xnor U3559 (N_3559,N_2520,N_2260);
or U3560 (N_3560,N_2245,N_2613);
nand U3561 (N_3561,N_2552,N_2885);
nor U3562 (N_3562,N_2899,N_2999);
or U3563 (N_3563,N_2552,N_2115);
or U3564 (N_3564,N_2135,N_2326);
and U3565 (N_3565,N_2213,N_2945);
and U3566 (N_3566,N_2687,N_2902);
and U3567 (N_3567,N_2843,N_2684);
and U3568 (N_3568,N_2159,N_2697);
nor U3569 (N_3569,N_2141,N_2802);
nand U3570 (N_3570,N_2718,N_2028);
nor U3571 (N_3571,N_2065,N_2117);
or U3572 (N_3572,N_2877,N_2253);
and U3573 (N_3573,N_2381,N_2592);
and U3574 (N_3574,N_2758,N_2746);
or U3575 (N_3575,N_2942,N_2202);
nor U3576 (N_3576,N_2763,N_2867);
nor U3577 (N_3577,N_2982,N_2606);
nor U3578 (N_3578,N_2813,N_2791);
or U3579 (N_3579,N_2771,N_2630);
nor U3580 (N_3580,N_2013,N_2931);
nand U3581 (N_3581,N_2777,N_2287);
nand U3582 (N_3582,N_2496,N_2001);
nand U3583 (N_3583,N_2010,N_2299);
or U3584 (N_3584,N_2571,N_2003);
and U3585 (N_3585,N_2627,N_2805);
nor U3586 (N_3586,N_2940,N_2096);
and U3587 (N_3587,N_2730,N_2864);
xor U3588 (N_3588,N_2945,N_2138);
xor U3589 (N_3589,N_2026,N_2102);
and U3590 (N_3590,N_2158,N_2536);
xor U3591 (N_3591,N_2175,N_2791);
nor U3592 (N_3592,N_2604,N_2559);
nand U3593 (N_3593,N_2957,N_2498);
xor U3594 (N_3594,N_2031,N_2974);
nand U3595 (N_3595,N_2143,N_2481);
xnor U3596 (N_3596,N_2074,N_2909);
nand U3597 (N_3597,N_2546,N_2244);
nand U3598 (N_3598,N_2350,N_2322);
nand U3599 (N_3599,N_2127,N_2068);
and U3600 (N_3600,N_2678,N_2417);
nand U3601 (N_3601,N_2899,N_2253);
and U3602 (N_3602,N_2478,N_2557);
and U3603 (N_3603,N_2851,N_2341);
or U3604 (N_3604,N_2208,N_2645);
nand U3605 (N_3605,N_2028,N_2119);
or U3606 (N_3606,N_2815,N_2686);
nand U3607 (N_3607,N_2105,N_2805);
and U3608 (N_3608,N_2455,N_2557);
nand U3609 (N_3609,N_2376,N_2392);
nor U3610 (N_3610,N_2718,N_2890);
nor U3611 (N_3611,N_2447,N_2464);
or U3612 (N_3612,N_2343,N_2700);
and U3613 (N_3613,N_2032,N_2828);
nor U3614 (N_3614,N_2252,N_2372);
nor U3615 (N_3615,N_2842,N_2214);
nand U3616 (N_3616,N_2825,N_2906);
xnor U3617 (N_3617,N_2330,N_2567);
and U3618 (N_3618,N_2628,N_2789);
nor U3619 (N_3619,N_2231,N_2334);
or U3620 (N_3620,N_2017,N_2522);
or U3621 (N_3621,N_2991,N_2008);
xor U3622 (N_3622,N_2053,N_2264);
or U3623 (N_3623,N_2754,N_2233);
nor U3624 (N_3624,N_2169,N_2402);
or U3625 (N_3625,N_2268,N_2063);
or U3626 (N_3626,N_2314,N_2121);
nand U3627 (N_3627,N_2714,N_2659);
or U3628 (N_3628,N_2126,N_2510);
or U3629 (N_3629,N_2089,N_2932);
nor U3630 (N_3630,N_2426,N_2483);
nor U3631 (N_3631,N_2696,N_2224);
nor U3632 (N_3632,N_2938,N_2998);
xnor U3633 (N_3633,N_2869,N_2014);
and U3634 (N_3634,N_2512,N_2676);
and U3635 (N_3635,N_2917,N_2360);
and U3636 (N_3636,N_2962,N_2930);
nand U3637 (N_3637,N_2601,N_2116);
or U3638 (N_3638,N_2097,N_2428);
nor U3639 (N_3639,N_2277,N_2233);
nand U3640 (N_3640,N_2187,N_2593);
and U3641 (N_3641,N_2738,N_2700);
nor U3642 (N_3642,N_2916,N_2236);
or U3643 (N_3643,N_2225,N_2546);
nor U3644 (N_3644,N_2496,N_2556);
nand U3645 (N_3645,N_2609,N_2125);
nand U3646 (N_3646,N_2739,N_2514);
nand U3647 (N_3647,N_2034,N_2788);
nand U3648 (N_3648,N_2330,N_2344);
nand U3649 (N_3649,N_2246,N_2131);
and U3650 (N_3650,N_2039,N_2223);
nand U3651 (N_3651,N_2919,N_2264);
and U3652 (N_3652,N_2856,N_2627);
and U3653 (N_3653,N_2987,N_2583);
and U3654 (N_3654,N_2445,N_2600);
or U3655 (N_3655,N_2417,N_2412);
nand U3656 (N_3656,N_2736,N_2871);
and U3657 (N_3657,N_2616,N_2378);
xnor U3658 (N_3658,N_2139,N_2525);
nand U3659 (N_3659,N_2065,N_2297);
nand U3660 (N_3660,N_2118,N_2319);
nor U3661 (N_3661,N_2103,N_2570);
or U3662 (N_3662,N_2519,N_2964);
or U3663 (N_3663,N_2935,N_2151);
nor U3664 (N_3664,N_2029,N_2821);
or U3665 (N_3665,N_2316,N_2298);
nor U3666 (N_3666,N_2341,N_2205);
xnor U3667 (N_3667,N_2152,N_2979);
and U3668 (N_3668,N_2562,N_2750);
nand U3669 (N_3669,N_2323,N_2749);
nor U3670 (N_3670,N_2877,N_2999);
nor U3671 (N_3671,N_2058,N_2229);
or U3672 (N_3672,N_2131,N_2424);
and U3673 (N_3673,N_2508,N_2654);
nor U3674 (N_3674,N_2962,N_2487);
nand U3675 (N_3675,N_2437,N_2349);
nand U3676 (N_3676,N_2765,N_2943);
or U3677 (N_3677,N_2340,N_2290);
nor U3678 (N_3678,N_2408,N_2160);
or U3679 (N_3679,N_2689,N_2812);
and U3680 (N_3680,N_2059,N_2421);
or U3681 (N_3681,N_2976,N_2583);
xnor U3682 (N_3682,N_2454,N_2946);
or U3683 (N_3683,N_2027,N_2853);
nor U3684 (N_3684,N_2293,N_2523);
or U3685 (N_3685,N_2404,N_2693);
xor U3686 (N_3686,N_2050,N_2053);
nand U3687 (N_3687,N_2255,N_2252);
nand U3688 (N_3688,N_2107,N_2748);
nand U3689 (N_3689,N_2129,N_2071);
and U3690 (N_3690,N_2524,N_2780);
and U3691 (N_3691,N_2424,N_2343);
and U3692 (N_3692,N_2364,N_2930);
nand U3693 (N_3693,N_2219,N_2142);
nand U3694 (N_3694,N_2588,N_2297);
or U3695 (N_3695,N_2830,N_2297);
or U3696 (N_3696,N_2968,N_2085);
nor U3697 (N_3697,N_2599,N_2009);
nand U3698 (N_3698,N_2696,N_2860);
nand U3699 (N_3699,N_2924,N_2236);
nor U3700 (N_3700,N_2067,N_2523);
xnor U3701 (N_3701,N_2313,N_2620);
and U3702 (N_3702,N_2922,N_2986);
nand U3703 (N_3703,N_2408,N_2449);
nand U3704 (N_3704,N_2337,N_2402);
nand U3705 (N_3705,N_2858,N_2764);
nor U3706 (N_3706,N_2803,N_2017);
and U3707 (N_3707,N_2003,N_2442);
and U3708 (N_3708,N_2723,N_2837);
or U3709 (N_3709,N_2922,N_2195);
nand U3710 (N_3710,N_2233,N_2674);
and U3711 (N_3711,N_2993,N_2783);
nor U3712 (N_3712,N_2418,N_2152);
nand U3713 (N_3713,N_2527,N_2480);
xnor U3714 (N_3714,N_2896,N_2761);
xnor U3715 (N_3715,N_2525,N_2392);
nand U3716 (N_3716,N_2068,N_2724);
or U3717 (N_3717,N_2707,N_2199);
nor U3718 (N_3718,N_2983,N_2725);
or U3719 (N_3719,N_2888,N_2561);
nor U3720 (N_3720,N_2582,N_2111);
or U3721 (N_3721,N_2605,N_2030);
nand U3722 (N_3722,N_2137,N_2539);
nand U3723 (N_3723,N_2172,N_2830);
nand U3724 (N_3724,N_2189,N_2485);
nor U3725 (N_3725,N_2435,N_2354);
xnor U3726 (N_3726,N_2672,N_2478);
and U3727 (N_3727,N_2270,N_2028);
and U3728 (N_3728,N_2447,N_2131);
nor U3729 (N_3729,N_2363,N_2470);
nand U3730 (N_3730,N_2115,N_2055);
or U3731 (N_3731,N_2902,N_2653);
nor U3732 (N_3732,N_2308,N_2347);
xor U3733 (N_3733,N_2138,N_2831);
or U3734 (N_3734,N_2132,N_2128);
nor U3735 (N_3735,N_2934,N_2433);
or U3736 (N_3736,N_2820,N_2803);
xnor U3737 (N_3737,N_2198,N_2656);
and U3738 (N_3738,N_2249,N_2988);
or U3739 (N_3739,N_2493,N_2771);
or U3740 (N_3740,N_2122,N_2090);
nand U3741 (N_3741,N_2552,N_2689);
nor U3742 (N_3742,N_2119,N_2732);
or U3743 (N_3743,N_2621,N_2916);
nor U3744 (N_3744,N_2934,N_2348);
nor U3745 (N_3745,N_2653,N_2112);
and U3746 (N_3746,N_2644,N_2704);
nand U3747 (N_3747,N_2448,N_2457);
nand U3748 (N_3748,N_2925,N_2430);
xnor U3749 (N_3749,N_2217,N_2510);
nor U3750 (N_3750,N_2834,N_2887);
nand U3751 (N_3751,N_2878,N_2170);
and U3752 (N_3752,N_2289,N_2073);
and U3753 (N_3753,N_2695,N_2322);
nor U3754 (N_3754,N_2153,N_2374);
nand U3755 (N_3755,N_2182,N_2699);
or U3756 (N_3756,N_2105,N_2038);
xnor U3757 (N_3757,N_2528,N_2575);
nor U3758 (N_3758,N_2773,N_2246);
nand U3759 (N_3759,N_2647,N_2115);
nor U3760 (N_3760,N_2424,N_2734);
nor U3761 (N_3761,N_2487,N_2760);
nand U3762 (N_3762,N_2551,N_2237);
and U3763 (N_3763,N_2834,N_2199);
and U3764 (N_3764,N_2416,N_2618);
and U3765 (N_3765,N_2690,N_2150);
and U3766 (N_3766,N_2650,N_2588);
nor U3767 (N_3767,N_2166,N_2481);
and U3768 (N_3768,N_2422,N_2638);
nand U3769 (N_3769,N_2515,N_2506);
nand U3770 (N_3770,N_2409,N_2089);
xnor U3771 (N_3771,N_2787,N_2339);
or U3772 (N_3772,N_2673,N_2129);
nor U3773 (N_3773,N_2818,N_2432);
nand U3774 (N_3774,N_2061,N_2196);
and U3775 (N_3775,N_2262,N_2604);
nand U3776 (N_3776,N_2639,N_2846);
nor U3777 (N_3777,N_2452,N_2967);
and U3778 (N_3778,N_2925,N_2197);
or U3779 (N_3779,N_2351,N_2816);
nand U3780 (N_3780,N_2356,N_2099);
nor U3781 (N_3781,N_2740,N_2843);
xor U3782 (N_3782,N_2701,N_2579);
and U3783 (N_3783,N_2759,N_2467);
and U3784 (N_3784,N_2493,N_2679);
or U3785 (N_3785,N_2914,N_2658);
nor U3786 (N_3786,N_2718,N_2267);
nand U3787 (N_3787,N_2712,N_2491);
or U3788 (N_3788,N_2296,N_2823);
nor U3789 (N_3789,N_2608,N_2242);
nor U3790 (N_3790,N_2154,N_2128);
or U3791 (N_3791,N_2827,N_2717);
or U3792 (N_3792,N_2307,N_2759);
nand U3793 (N_3793,N_2025,N_2775);
and U3794 (N_3794,N_2992,N_2406);
nand U3795 (N_3795,N_2505,N_2409);
and U3796 (N_3796,N_2821,N_2414);
xor U3797 (N_3797,N_2897,N_2325);
nand U3798 (N_3798,N_2614,N_2988);
or U3799 (N_3799,N_2647,N_2979);
and U3800 (N_3800,N_2467,N_2531);
or U3801 (N_3801,N_2333,N_2707);
and U3802 (N_3802,N_2248,N_2394);
and U3803 (N_3803,N_2637,N_2225);
nor U3804 (N_3804,N_2877,N_2198);
xor U3805 (N_3805,N_2388,N_2101);
xor U3806 (N_3806,N_2156,N_2459);
and U3807 (N_3807,N_2956,N_2649);
or U3808 (N_3808,N_2148,N_2585);
nor U3809 (N_3809,N_2228,N_2477);
and U3810 (N_3810,N_2596,N_2442);
nand U3811 (N_3811,N_2790,N_2161);
or U3812 (N_3812,N_2584,N_2299);
nor U3813 (N_3813,N_2148,N_2267);
nand U3814 (N_3814,N_2506,N_2054);
or U3815 (N_3815,N_2302,N_2032);
and U3816 (N_3816,N_2682,N_2047);
or U3817 (N_3817,N_2313,N_2993);
or U3818 (N_3818,N_2901,N_2516);
or U3819 (N_3819,N_2226,N_2750);
nand U3820 (N_3820,N_2365,N_2023);
nand U3821 (N_3821,N_2814,N_2802);
nor U3822 (N_3822,N_2350,N_2707);
nand U3823 (N_3823,N_2634,N_2123);
and U3824 (N_3824,N_2599,N_2353);
and U3825 (N_3825,N_2628,N_2848);
nor U3826 (N_3826,N_2827,N_2478);
nor U3827 (N_3827,N_2809,N_2677);
and U3828 (N_3828,N_2792,N_2695);
nand U3829 (N_3829,N_2239,N_2588);
and U3830 (N_3830,N_2907,N_2836);
nand U3831 (N_3831,N_2459,N_2871);
nand U3832 (N_3832,N_2981,N_2056);
or U3833 (N_3833,N_2086,N_2286);
nand U3834 (N_3834,N_2564,N_2864);
xor U3835 (N_3835,N_2551,N_2031);
nand U3836 (N_3836,N_2593,N_2479);
or U3837 (N_3837,N_2443,N_2381);
xnor U3838 (N_3838,N_2284,N_2506);
or U3839 (N_3839,N_2999,N_2369);
nand U3840 (N_3840,N_2652,N_2480);
nor U3841 (N_3841,N_2534,N_2811);
or U3842 (N_3842,N_2875,N_2140);
or U3843 (N_3843,N_2860,N_2070);
nand U3844 (N_3844,N_2418,N_2618);
or U3845 (N_3845,N_2850,N_2265);
xor U3846 (N_3846,N_2277,N_2482);
nor U3847 (N_3847,N_2364,N_2816);
nor U3848 (N_3848,N_2796,N_2985);
xor U3849 (N_3849,N_2831,N_2988);
or U3850 (N_3850,N_2573,N_2592);
or U3851 (N_3851,N_2404,N_2541);
nand U3852 (N_3852,N_2451,N_2947);
or U3853 (N_3853,N_2757,N_2605);
nor U3854 (N_3854,N_2272,N_2944);
nor U3855 (N_3855,N_2973,N_2166);
nor U3856 (N_3856,N_2336,N_2051);
and U3857 (N_3857,N_2277,N_2993);
nor U3858 (N_3858,N_2560,N_2053);
xnor U3859 (N_3859,N_2382,N_2773);
nor U3860 (N_3860,N_2918,N_2606);
xor U3861 (N_3861,N_2962,N_2892);
nand U3862 (N_3862,N_2246,N_2348);
nand U3863 (N_3863,N_2179,N_2497);
nand U3864 (N_3864,N_2190,N_2761);
and U3865 (N_3865,N_2639,N_2838);
nand U3866 (N_3866,N_2946,N_2028);
or U3867 (N_3867,N_2248,N_2082);
or U3868 (N_3868,N_2295,N_2855);
or U3869 (N_3869,N_2779,N_2381);
nand U3870 (N_3870,N_2577,N_2830);
or U3871 (N_3871,N_2893,N_2698);
or U3872 (N_3872,N_2494,N_2632);
xor U3873 (N_3873,N_2574,N_2330);
nor U3874 (N_3874,N_2956,N_2527);
or U3875 (N_3875,N_2043,N_2732);
nand U3876 (N_3876,N_2884,N_2236);
nor U3877 (N_3877,N_2730,N_2567);
xor U3878 (N_3878,N_2760,N_2979);
and U3879 (N_3879,N_2212,N_2813);
nand U3880 (N_3880,N_2460,N_2444);
or U3881 (N_3881,N_2323,N_2348);
nor U3882 (N_3882,N_2713,N_2490);
xor U3883 (N_3883,N_2234,N_2338);
nand U3884 (N_3884,N_2559,N_2359);
and U3885 (N_3885,N_2114,N_2467);
nand U3886 (N_3886,N_2103,N_2012);
nor U3887 (N_3887,N_2832,N_2355);
nor U3888 (N_3888,N_2928,N_2191);
xnor U3889 (N_3889,N_2128,N_2166);
or U3890 (N_3890,N_2909,N_2644);
nor U3891 (N_3891,N_2524,N_2671);
nor U3892 (N_3892,N_2550,N_2112);
nand U3893 (N_3893,N_2713,N_2472);
or U3894 (N_3894,N_2644,N_2147);
nand U3895 (N_3895,N_2543,N_2011);
or U3896 (N_3896,N_2730,N_2336);
or U3897 (N_3897,N_2429,N_2578);
and U3898 (N_3898,N_2044,N_2344);
nand U3899 (N_3899,N_2264,N_2078);
xnor U3900 (N_3900,N_2229,N_2938);
nor U3901 (N_3901,N_2906,N_2282);
and U3902 (N_3902,N_2048,N_2664);
nand U3903 (N_3903,N_2424,N_2503);
or U3904 (N_3904,N_2401,N_2784);
or U3905 (N_3905,N_2146,N_2419);
or U3906 (N_3906,N_2875,N_2630);
or U3907 (N_3907,N_2349,N_2934);
nor U3908 (N_3908,N_2621,N_2927);
nor U3909 (N_3909,N_2607,N_2199);
or U3910 (N_3910,N_2949,N_2834);
or U3911 (N_3911,N_2504,N_2973);
nor U3912 (N_3912,N_2998,N_2427);
or U3913 (N_3913,N_2961,N_2557);
or U3914 (N_3914,N_2458,N_2801);
nand U3915 (N_3915,N_2322,N_2803);
nor U3916 (N_3916,N_2082,N_2959);
nor U3917 (N_3917,N_2291,N_2073);
xnor U3918 (N_3918,N_2887,N_2948);
or U3919 (N_3919,N_2602,N_2798);
and U3920 (N_3920,N_2447,N_2794);
nor U3921 (N_3921,N_2742,N_2644);
nor U3922 (N_3922,N_2810,N_2145);
nand U3923 (N_3923,N_2812,N_2817);
or U3924 (N_3924,N_2620,N_2676);
and U3925 (N_3925,N_2260,N_2529);
or U3926 (N_3926,N_2118,N_2022);
nand U3927 (N_3927,N_2839,N_2384);
and U3928 (N_3928,N_2838,N_2728);
nand U3929 (N_3929,N_2082,N_2716);
or U3930 (N_3930,N_2488,N_2726);
and U3931 (N_3931,N_2181,N_2233);
nand U3932 (N_3932,N_2478,N_2070);
nand U3933 (N_3933,N_2373,N_2633);
nor U3934 (N_3934,N_2214,N_2863);
nand U3935 (N_3935,N_2656,N_2027);
nand U3936 (N_3936,N_2986,N_2085);
or U3937 (N_3937,N_2678,N_2103);
nand U3938 (N_3938,N_2764,N_2398);
xor U3939 (N_3939,N_2597,N_2403);
or U3940 (N_3940,N_2744,N_2991);
nor U3941 (N_3941,N_2612,N_2940);
nand U3942 (N_3942,N_2017,N_2537);
xor U3943 (N_3943,N_2671,N_2886);
nand U3944 (N_3944,N_2898,N_2672);
and U3945 (N_3945,N_2063,N_2671);
nand U3946 (N_3946,N_2080,N_2930);
and U3947 (N_3947,N_2179,N_2514);
nor U3948 (N_3948,N_2391,N_2109);
nor U3949 (N_3949,N_2978,N_2403);
xor U3950 (N_3950,N_2179,N_2695);
and U3951 (N_3951,N_2074,N_2914);
nand U3952 (N_3952,N_2377,N_2589);
nand U3953 (N_3953,N_2567,N_2488);
nand U3954 (N_3954,N_2638,N_2739);
or U3955 (N_3955,N_2152,N_2568);
or U3956 (N_3956,N_2768,N_2802);
nand U3957 (N_3957,N_2423,N_2761);
nand U3958 (N_3958,N_2431,N_2810);
or U3959 (N_3959,N_2263,N_2934);
or U3960 (N_3960,N_2444,N_2096);
nand U3961 (N_3961,N_2394,N_2358);
nand U3962 (N_3962,N_2261,N_2536);
and U3963 (N_3963,N_2746,N_2261);
and U3964 (N_3964,N_2278,N_2554);
and U3965 (N_3965,N_2128,N_2538);
nand U3966 (N_3966,N_2199,N_2838);
and U3967 (N_3967,N_2492,N_2158);
and U3968 (N_3968,N_2757,N_2634);
nand U3969 (N_3969,N_2083,N_2583);
nand U3970 (N_3970,N_2361,N_2760);
nor U3971 (N_3971,N_2662,N_2579);
and U3972 (N_3972,N_2506,N_2064);
and U3973 (N_3973,N_2483,N_2669);
and U3974 (N_3974,N_2067,N_2899);
and U3975 (N_3975,N_2510,N_2079);
nand U3976 (N_3976,N_2785,N_2935);
nand U3977 (N_3977,N_2581,N_2194);
nor U3978 (N_3978,N_2875,N_2691);
or U3979 (N_3979,N_2862,N_2204);
and U3980 (N_3980,N_2520,N_2804);
or U3981 (N_3981,N_2880,N_2804);
nor U3982 (N_3982,N_2831,N_2273);
nor U3983 (N_3983,N_2263,N_2634);
nand U3984 (N_3984,N_2085,N_2661);
nor U3985 (N_3985,N_2358,N_2207);
nor U3986 (N_3986,N_2141,N_2067);
nand U3987 (N_3987,N_2640,N_2091);
or U3988 (N_3988,N_2788,N_2697);
nor U3989 (N_3989,N_2158,N_2517);
xnor U3990 (N_3990,N_2555,N_2531);
or U3991 (N_3991,N_2020,N_2464);
and U3992 (N_3992,N_2547,N_2034);
nor U3993 (N_3993,N_2210,N_2765);
nand U3994 (N_3994,N_2112,N_2075);
nor U3995 (N_3995,N_2108,N_2226);
nand U3996 (N_3996,N_2835,N_2859);
and U3997 (N_3997,N_2785,N_2205);
xor U3998 (N_3998,N_2186,N_2440);
nor U3999 (N_3999,N_2548,N_2847);
nor U4000 (N_4000,N_3329,N_3325);
and U4001 (N_4001,N_3159,N_3455);
nor U4002 (N_4002,N_3569,N_3151);
nor U4003 (N_4003,N_3383,N_3533);
and U4004 (N_4004,N_3520,N_3235);
or U4005 (N_4005,N_3759,N_3493);
or U4006 (N_4006,N_3084,N_3788);
and U4007 (N_4007,N_3993,N_3295);
nand U4008 (N_4008,N_3089,N_3584);
and U4009 (N_4009,N_3248,N_3983);
nor U4010 (N_4010,N_3179,N_3884);
nor U4011 (N_4011,N_3800,N_3036);
nand U4012 (N_4012,N_3504,N_3103);
or U4013 (N_4013,N_3540,N_3515);
nand U4014 (N_4014,N_3136,N_3738);
nand U4015 (N_4015,N_3698,N_3213);
and U4016 (N_4016,N_3463,N_3686);
nor U4017 (N_4017,N_3385,N_3966);
or U4018 (N_4018,N_3557,N_3953);
nor U4019 (N_4019,N_3960,N_3560);
nor U4020 (N_4020,N_3491,N_3715);
nor U4021 (N_4021,N_3739,N_3886);
nand U4022 (N_4022,N_3361,N_3796);
nor U4023 (N_4023,N_3845,N_3681);
xnor U4024 (N_4024,N_3651,N_3776);
nor U4025 (N_4025,N_3967,N_3790);
nor U4026 (N_4026,N_3995,N_3287);
nor U4027 (N_4027,N_3674,N_3128);
nand U4028 (N_4028,N_3895,N_3032);
or U4029 (N_4029,N_3158,N_3414);
and U4030 (N_4030,N_3180,N_3453);
or U4031 (N_4031,N_3372,N_3530);
and U4032 (N_4032,N_3044,N_3870);
nor U4033 (N_4033,N_3989,N_3605);
nor U4034 (N_4034,N_3598,N_3402);
nor U4035 (N_4035,N_3801,N_3577);
nor U4036 (N_4036,N_3282,N_3363);
nand U4037 (N_4037,N_3052,N_3269);
nor U4038 (N_4038,N_3413,N_3003);
nand U4039 (N_4039,N_3452,N_3568);
and U4040 (N_4040,N_3571,N_3029);
or U4041 (N_4041,N_3318,N_3147);
or U4042 (N_4042,N_3410,N_3204);
and U4043 (N_4043,N_3654,N_3205);
xnor U4044 (N_4044,N_3711,N_3604);
or U4045 (N_4045,N_3538,N_3426);
nand U4046 (N_4046,N_3603,N_3623);
or U4047 (N_4047,N_3648,N_3547);
or U4048 (N_4048,N_3169,N_3767);
or U4049 (N_4049,N_3545,N_3197);
nor U4050 (N_4050,N_3659,N_3497);
and U4051 (N_4051,N_3411,N_3108);
and U4052 (N_4052,N_3885,N_3183);
xor U4053 (N_4053,N_3041,N_3375);
nor U4054 (N_4054,N_3883,N_3393);
and U4055 (N_4055,N_3358,N_3717);
and U4056 (N_4056,N_3233,N_3071);
or U4057 (N_4057,N_3498,N_3432);
nand U4058 (N_4058,N_3521,N_3792);
nand U4059 (N_4059,N_3002,N_3823);
nand U4060 (N_4060,N_3900,N_3735);
nor U4061 (N_4061,N_3203,N_3035);
nand U4062 (N_4062,N_3665,N_3317);
xnor U4063 (N_4063,N_3890,N_3555);
and U4064 (N_4064,N_3579,N_3914);
and U4065 (N_4065,N_3333,N_3502);
nor U4066 (N_4066,N_3763,N_3892);
or U4067 (N_4067,N_3795,N_3457);
nand U4068 (N_4068,N_3961,N_3246);
nor U4069 (N_4069,N_3947,N_3118);
and U4070 (N_4070,N_3524,N_3042);
nor U4071 (N_4071,N_3285,N_3311);
and U4072 (N_4072,N_3682,N_3423);
nor U4073 (N_4073,N_3572,N_3722);
nor U4074 (N_4074,N_3589,N_3458);
and U4075 (N_4075,N_3219,N_3748);
or U4076 (N_4076,N_3775,N_3630);
nor U4077 (N_4077,N_3543,N_3783);
nand U4078 (N_4078,N_3011,N_3805);
and U4079 (N_4079,N_3825,N_3643);
nor U4080 (N_4080,N_3242,N_3652);
and U4081 (N_4081,N_3326,N_3370);
and U4082 (N_4082,N_3069,N_3184);
nor U4083 (N_4083,N_3461,N_3534);
or U4084 (N_4084,N_3818,N_3086);
nor U4085 (N_4085,N_3516,N_3239);
and U4086 (N_4086,N_3119,N_3033);
nand U4087 (N_4087,N_3274,N_3847);
nor U4088 (N_4088,N_3428,N_3951);
and U4089 (N_4089,N_3580,N_3403);
and U4090 (N_4090,N_3250,N_3996);
or U4091 (N_4091,N_3125,N_3418);
nor U4092 (N_4092,N_3039,N_3396);
nand U4093 (N_4093,N_3244,N_3709);
nor U4094 (N_4094,N_3142,N_3982);
and U4095 (N_4095,N_3309,N_3321);
or U4096 (N_4096,N_3487,N_3808);
nor U4097 (N_4097,N_3171,N_3310);
nor U4098 (N_4098,N_3078,N_3669);
nand U4099 (N_4099,N_3240,N_3561);
nor U4100 (N_4100,N_3658,N_3588);
and U4101 (N_4101,N_3905,N_3469);
nand U4102 (N_4102,N_3211,N_3009);
nor U4103 (N_4103,N_3189,N_3936);
and U4104 (N_4104,N_3680,N_3859);
nand U4105 (N_4105,N_3111,N_3077);
and U4106 (N_4106,N_3021,N_3693);
or U4107 (N_4107,N_3950,N_3852);
nand U4108 (N_4108,N_3956,N_3830);
or U4109 (N_4109,N_3733,N_3121);
xor U4110 (N_4110,N_3388,N_3273);
and U4111 (N_4111,N_3175,N_3924);
nor U4112 (N_4112,N_3196,N_3050);
nor U4113 (N_4113,N_3632,N_3997);
xnor U4114 (N_4114,N_3292,N_3344);
and U4115 (N_4115,N_3064,N_3208);
nand U4116 (N_4116,N_3312,N_3695);
or U4117 (N_4117,N_3758,N_3928);
and U4118 (N_4118,N_3929,N_3869);
nand U4119 (N_4119,N_3839,N_3153);
or U4120 (N_4120,N_3278,N_3575);
nand U4121 (N_4121,N_3721,N_3148);
nor U4122 (N_4122,N_3080,N_3815);
xor U4123 (N_4123,N_3440,N_3958);
nor U4124 (N_4124,N_3744,N_3489);
nor U4125 (N_4125,N_3880,N_3000);
and U4126 (N_4126,N_3416,N_3083);
and U4127 (N_4127,N_3764,N_3412);
nand U4128 (N_4128,N_3434,N_3262);
nand U4129 (N_4129,N_3467,N_3096);
nand U4130 (N_4130,N_3952,N_3694);
nand U4131 (N_4131,N_3139,N_3846);
and U4132 (N_4132,N_3821,N_3523);
nor U4133 (N_4133,N_3451,N_3220);
and U4134 (N_4134,N_3065,N_3867);
or U4135 (N_4135,N_3713,N_3356);
nand U4136 (N_4136,N_3802,N_3728);
or U4137 (N_4137,N_3186,N_3712);
or U4138 (N_4138,N_3727,N_3488);
or U4139 (N_4139,N_3877,N_3746);
xor U4140 (N_4140,N_3229,N_3117);
and U4141 (N_4141,N_3275,N_3324);
nand U4142 (N_4142,N_3822,N_3480);
and U4143 (N_4143,N_3703,N_3760);
nor U4144 (N_4144,N_3930,N_3368);
nand U4145 (N_4145,N_3509,N_3181);
nor U4146 (N_4146,N_3798,N_3201);
and U4147 (N_4147,N_3062,N_3627);
nand U4148 (N_4148,N_3610,N_3191);
nand U4149 (N_4149,N_3789,N_3657);
nor U4150 (N_4150,N_3499,N_3305);
or U4151 (N_4151,N_3655,N_3421);
nor U4152 (N_4152,N_3200,N_3948);
xor U4153 (N_4153,N_3550,N_3761);
or U4154 (N_4154,N_3770,N_3519);
nand U4155 (N_4155,N_3168,N_3109);
or U4156 (N_4156,N_3095,N_3602);
nand U4157 (N_4157,N_3970,N_3227);
and U4158 (N_4158,N_3409,N_3553);
and U4159 (N_4159,N_3261,N_3897);
nor U4160 (N_4160,N_3353,N_3638);
and U4161 (N_4161,N_3126,N_3018);
or U4162 (N_4162,N_3307,N_3620);
nand U4163 (N_4163,N_3391,N_3146);
nor U4164 (N_4164,N_3070,N_3755);
nor U4165 (N_4165,N_3536,N_3558);
or U4166 (N_4166,N_3718,N_3056);
nor U4167 (N_4167,N_3639,N_3696);
or U4168 (N_4168,N_3829,N_3150);
or U4169 (N_4169,N_3909,N_3689);
nand U4170 (N_4170,N_3592,N_3981);
and U4171 (N_4171,N_3864,N_3286);
nor U4172 (N_4172,N_3591,N_3915);
and U4173 (N_4173,N_3962,N_3088);
nand U4174 (N_4174,N_3851,N_3230);
and U4175 (N_4175,N_3094,N_3397);
nand U4176 (N_4176,N_3228,N_3855);
or U4177 (N_4177,N_3366,N_3124);
or U4178 (N_4178,N_3898,N_3221);
or U4179 (N_4179,N_3833,N_3621);
or U4180 (N_4180,N_3820,N_3777);
and U4181 (N_4181,N_3300,N_3678);
and U4182 (N_4182,N_3145,N_3023);
nand U4183 (N_4183,N_3209,N_3773);
nand U4184 (N_4184,N_3048,N_3247);
or U4185 (N_4185,N_3214,N_3192);
or U4186 (N_4186,N_3386,N_3743);
xnor U4187 (N_4187,N_3031,N_3600);
nor U4188 (N_4188,N_3918,N_3508);
nor U4189 (N_4189,N_3774,N_3236);
nand U4190 (N_4190,N_3185,N_3231);
nand U4191 (N_4191,N_3435,N_3010);
and U4192 (N_4192,N_3384,N_3445);
nand U4193 (N_4193,N_3026,N_3263);
and U4194 (N_4194,N_3133,N_3719);
xnor U4195 (N_4195,N_3336,N_3155);
nand U4196 (N_4196,N_3373,N_3296);
or U4197 (N_4197,N_3264,N_3762);
and U4198 (N_4198,N_3587,N_3038);
nand U4199 (N_4199,N_3157,N_3490);
and U4200 (N_4200,N_3645,N_3351);
or U4201 (N_4201,N_3433,N_3673);
or U4202 (N_4202,N_3955,N_3076);
and U4203 (N_4203,N_3249,N_3215);
and U4204 (N_4204,N_3943,N_3430);
and U4205 (N_4205,N_3653,N_3978);
and U4206 (N_4206,N_3985,N_3838);
xor U4207 (N_4207,N_3268,N_3170);
or U4208 (N_4208,N_3857,N_3615);
nor U4209 (N_4209,N_3848,N_3398);
nand U4210 (N_4210,N_3628,N_3597);
and U4211 (N_4211,N_3283,N_3465);
nor U4212 (N_4212,N_3258,N_3299);
and U4213 (N_4213,N_3656,N_3327);
nor U4214 (N_4214,N_3710,N_3888);
xnor U4215 (N_4215,N_3097,N_3431);
nand U4216 (N_4216,N_3644,N_3688);
or U4217 (N_4217,N_3834,N_3772);
or U4218 (N_4218,N_3872,N_3700);
xor U4219 (N_4219,N_3475,N_3182);
nand U4220 (N_4220,N_3899,N_3135);
or U4221 (N_4221,N_3276,N_3176);
nor U4222 (N_4222,N_3944,N_3616);
nand U4223 (N_4223,N_3706,N_3741);
nor U4224 (N_4224,N_3672,N_3716);
nand U4225 (N_4225,N_3562,N_3359);
and U4226 (N_4226,N_3861,N_3771);
nand U4227 (N_4227,N_3190,N_3174);
and U4228 (N_4228,N_3259,N_3456);
or U4229 (N_4229,N_3570,N_3692);
xnor U4230 (N_4230,N_3766,N_3875);
nor U4231 (N_4231,N_3871,N_3389);
and U4232 (N_4232,N_3690,N_3328);
nor U4233 (N_4233,N_3866,N_3750);
nand U4234 (N_4234,N_3751,N_3510);
or U4235 (N_4235,N_3163,N_3816);
xnor U4236 (N_4236,N_3315,N_3040);
and U4237 (N_4237,N_3544,N_3606);
and U4238 (N_4238,N_3532,N_3392);
nand U4239 (N_4239,N_3290,N_3154);
and U4240 (N_4240,N_3850,N_3302);
nand U4241 (N_4241,N_3232,N_3152);
nor U4242 (N_4242,N_3559,N_3980);
nand U4243 (N_4243,N_3210,N_3277);
nand U4244 (N_4244,N_3140,N_3008);
xnor U4245 (N_4245,N_3831,N_3723);
xor U4246 (N_4246,N_3454,N_3194);
xor U4247 (N_4247,N_3974,N_3664);
or U4248 (N_4248,N_3786,N_3685);
and U4249 (N_4249,N_3496,N_3666);
nor U4250 (N_4250,N_3484,N_3293);
xor U4251 (N_4251,N_3986,N_3217);
xor U4252 (N_4252,N_3676,N_3503);
and U4253 (N_4253,N_3068,N_3406);
or U4254 (N_4254,N_3090,N_3992);
and U4255 (N_4255,N_3531,N_3522);
and U4256 (N_4256,N_3878,N_3099);
nand U4257 (N_4257,N_3791,N_3034);
xor U4258 (N_4258,N_3752,N_3724);
xnor U4259 (N_4259,N_3260,N_3253);
nand U4260 (N_4260,N_3072,N_3518);
xor U4261 (N_4261,N_3408,N_3517);
nand U4262 (N_4262,N_3505,N_3374);
and U4263 (N_4263,N_3622,N_3267);
nand U4264 (N_4264,N_3225,N_3684);
and U4265 (N_4265,N_3173,N_3471);
or U4266 (N_4266,N_3799,N_3566);
nand U4267 (N_4267,N_3853,N_3889);
or U4268 (N_4268,N_3882,N_3486);
or U4269 (N_4269,N_3856,N_3495);
nor U4270 (N_4270,N_3049,N_3891);
and U4271 (N_4271,N_3976,N_3782);
nand U4272 (N_4272,N_3301,N_3443);
xnor U4273 (N_4273,N_3542,N_3641);
nand U4274 (N_4274,N_3964,N_3779);
nor U4275 (N_4275,N_3514,N_3378);
and U4276 (N_4276,N_3345,N_3707);
or U4277 (N_4277,N_3459,N_3051);
nor U4278 (N_4278,N_3593,N_3313);
or U4279 (N_4279,N_3991,N_3731);
nand U4280 (N_4280,N_3166,N_3331);
xor U4281 (N_4281,N_3102,N_3687);
xor U4282 (N_4282,N_3691,N_3279);
nor U4283 (N_4283,N_3780,N_3007);
nor U4284 (N_4284,N_3187,N_3060);
nor U4285 (N_4285,N_3478,N_3994);
nor U4286 (N_4286,N_3357,N_3949);
and U4287 (N_4287,N_3303,N_3234);
nand U4288 (N_4288,N_3946,N_3424);
nand U4289 (N_4289,N_3419,N_3968);
nand U4290 (N_4290,N_3649,N_3811);
nor U4291 (N_4291,N_3226,N_3223);
or U4292 (N_4292,N_3107,N_3362);
and U4293 (N_4293,N_3784,N_3507);
nor U4294 (N_4294,N_3061,N_3708);
nand U4295 (N_4295,N_3873,N_3827);
nand U4296 (N_4296,N_3195,N_3549);
nor U4297 (N_4297,N_3617,N_3144);
and U4298 (N_4298,N_3104,N_3063);
and U4299 (N_4299,N_3699,N_3913);
nand U4300 (N_4300,N_3626,N_3400);
or U4301 (N_4301,N_3965,N_3939);
or U4302 (N_4302,N_3245,N_3025);
or U4303 (N_4303,N_3573,N_3216);
nor U4304 (N_4304,N_3998,N_3266);
xor U4305 (N_4305,N_3280,N_3595);
and U4306 (N_4306,N_3016,N_3932);
nor U4307 (N_4307,N_3807,N_3156);
nand U4308 (N_4308,N_3165,N_3319);
nor U4309 (N_4309,N_3954,N_3093);
and U4310 (N_4310,N_3841,N_3394);
and U4311 (N_4311,N_3134,N_3270);
nand U4312 (N_4312,N_3485,N_3500);
nand U4313 (N_4313,N_3619,N_3537);
nand U4314 (N_4314,N_3646,N_3323);
and U4315 (N_4315,N_3826,N_3824);
or U4316 (N_4316,N_3346,N_3612);
nand U4317 (N_4317,N_3129,N_3481);
nor U4318 (N_4318,N_3565,N_3222);
nor U4319 (N_4319,N_3896,N_3395);
and U4320 (N_4320,N_3637,N_3552);
nand U4321 (N_4321,N_3979,N_3339);
xnor U4322 (N_4322,N_3390,N_3251);
or U4323 (N_4323,N_3112,N_3629);
and U4324 (N_4324,N_3901,N_3564);
nor U4325 (N_4325,N_3675,N_3714);
nor U4326 (N_4326,N_3320,N_3427);
or U4327 (N_4327,N_3106,N_3447);
nand U4328 (N_4328,N_3868,N_3046);
nor U4329 (N_4329,N_3161,N_3330);
or U4330 (N_4330,N_3768,N_3574);
or U4331 (N_4331,N_3030,N_3919);
and U4332 (N_4332,N_3705,N_3417);
and U4333 (N_4333,N_3405,N_3081);
or U4334 (N_4334,N_3043,N_3482);
or U4335 (N_4335,N_3670,N_3683);
nor U4336 (N_4336,N_3137,N_3742);
or U4337 (N_4337,N_3726,N_3843);
xnor U4338 (N_4338,N_3702,N_3466);
nor U4339 (N_4339,N_3057,N_3661);
or U4340 (N_4340,N_3350,N_3840);
and U4341 (N_4341,N_3399,N_3047);
or U4342 (N_4342,N_3757,N_3100);
nand U4343 (N_4343,N_3460,N_3835);
and U4344 (N_4344,N_3272,N_3291);
and U4345 (N_4345,N_3740,N_3662);
nor U4346 (N_4346,N_3624,N_3828);
nand U4347 (N_4347,N_3576,N_3407);
and U4348 (N_4348,N_3611,N_3854);
nand U4349 (N_4349,N_3631,N_3640);
and U4350 (N_4350,N_3338,N_3581);
or U4351 (N_4351,N_3131,N_3349);
and U4352 (N_4352,N_3341,N_3304);
or U4353 (N_4353,N_3202,N_3472);
and U4354 (N_4354,N_3091,N_3923);
or U4355 (N_4355,N_3663,N_3288);
xor U4356 (N_4356,N_3005,N_3468);
and U4357 (N_4357,N_3720,N_3364);
or U4358 (N_4358,N_3198,N_3073);
and U4359 (N_4359,N_3024,N_3959);
nor U4360 (N_4360,N_3590,N_3441);
nor U4361 (N_4361,N_3667,N_3376);
or U4362 (N_4362,N_3793,N_3206);
nand U4363 (N_4363,N_3887,N_3725);
nor U4364 (N_4364,N_3127,N_3167);
and U4365 (N_4365,N_3483,N_3382);
or U4366 (N_4366,N_3902,N_3092);
nand U4367 (N_4367,N_3701,N_3563);
nor U4368 (N_4368,N_3753,N_3252);
nand U4369 (N_4369,N_3449,N_3477);
or U4370 (N_4370,N_3237,N_3922);
or U4371 (N_4371,N_3066,N_3613);
nor U4372 (N_4372,N_3347,N_3844);
and U4373 (N_4373,N_3511,N_3963);
nor U4374 (N_4374,N_3907,N_3355);
nor U4375 (N_4375,N_3474,N_3238);
nand U4376 (N_4376,N_3438,N_3284);
nand U4377 (N_4377,N_3614,N_3837);
nor U4378 (N_4378,N_3436,N_3212);
or U4379 (N_4379,N_3990,N_3585);
and U4380 (N_4380,N_3243,N_3367);
xnor U4381 (N_4381,N_3404,N_3813);
or U4382 (N_4382,N_3972,N_3879);
and U4383 (N_4383,N_3446,N_3401);
nor U4384 (N_4384,N_3164,N_3874);
nor U4385 (N_4385,N_3933,N_3420);
nand U4386 (N_4386,N_3527,N_3945);
nand U4387 (N_4387,N_3360,N_3437);
or U4388 (N_4388,N_3819,N_3218);
and U4389 (N_4389,N_3984,N_3832);
nand U4390 (N_4390,N_3849,N_3754);
and U4391 (N_4391,N_3594,N_3113);
nand U4392 (N_4392,N_3730,N_3794);
and U4393 (N_4393,N_3987,N_3925);
or U4394 (N_4394,N_3999,N_3015);
nor U4395 (N_4395,N_3006,N_3634);
and U4396 (N_4396,N_3917,N_3817);
nor U4397 (N_4397,N_3425,N_3546);
nor U4398 (N_4398,N_3354,N_3098);
nand U4399 (N_4399,N_3904,N_3609);
and U4400 (N_4400,N_3797,N_3814);
and U4401 (N_4401,N_3123,N_3941);
and U4402 (N_4402,N_3858,N_3747);
or U4403 (N_4403,N_3756,N_3462);
nor U4404 (N_4404,N_3059,N_3860);
nand U4405 (N_4405,N_3749,N_3316);
or U4406 (N_4406,N_3027,N_3241);
and U4407 (N_4407,N_3105,N_3865);
nand U4408 (N_4408,N_3037,N_3054);
and U4409 (N_4409,N_3938,N_3255);
and U4410 (N_4410,N_3314,N_3074);
or U4411 (N_4411,N_3380,N_3308);
nand U4412 (N_4412,N_3650,N_3732);
nand U4413 (N_4413,N_3332,N_3342);
and U4414 (N_4414,N_3541,N_3582);
and U4415 (N_4415,N_3803,N_3479);
nor U4416 (N_4416,N_3668,N_3642);
or U4417 (N_4417,N_3337,N_3058);
and U4418 (N_4418,N_3188,N_3528);
nor U4419 (N_4419,N_3130,N_3371);
nand U4420 (N_4420,N_3671,N_3492);
or U4421 (N_4421,N_3556,N_3608);
and U4422 (N_4422,N_3906,N_3138);
nor U4423 (N_4423,N_3271,N_3975);
or U4424 (N_4424,N_3931,N_3122);
and U4425 (N_4425,N_3607,N_3470);
nand U4426 (N_4426,N_3734,N_3893);
nor U4427 (N_4427,N_3087,N_3110);
nor U4428 (N_4428,N_3306,N_3625);
nand U4429 (N_4429,N_3551,N_3578);
and U4430 (N_4430,N_3017,N_3529);
and U4431 (N_4431,N_3369,N_3132);
and U4432 (N_4432,N_3012,N_3004);
nand U4433 (N_4433,N_3114,N_3804);
nand U4434 (N_4434,N_3476,N_3067);
nor U4435 (N_4435,N_3014,N_3298);
nand U4436 (N_4436,N_3281,N_3876);
nand U4437 (N_4437,N_3494,N_3916);
nor U4438 (N_4438,N_3920,N_3903);
or U4439 (N_4439,N_3082,N_3935);
nor U4440 (N_4440,N_3199,N_3526);
nor U4441 (N_4441,N_3448,N_3862);
and U4442 (N_4442,N_3019,N_3352);
nand U4443 (N_4443,N_3973,N_3377);
and U4444 (N_4444,N_3806,N_3075);
nor U4445 (N_4445,N_3335,N_3809);
nor U4446 (N_4446,N_3737,N_3116);
nand U4447 (N_4447,N_3921,N_3178);
and U4448 (N_4448,N_3863,N_3697);
or U4449 (N_4449,N_3745,N_3765);
or U4450 (N_4450,N_3842,N_3365);
or U4451 (N_4451,N_3387,N_3535);
and U4452 (N_4452,N_3415,N_3787);
xor U4453 (N_4453,N_3177,N_3442);
and U4454 (N_4454,N_3894,N_3957);
nor U4455 (N_4455,N_3971,N_3439);
xor U4456 (N_4456,N_3506,N_3115);
nand U4457 (N_4457,N_3020,N_3567);
nand U4458 (N_4458,N_3729,N_3207);
or U4459 (N_4459,N_3473,N_3289);
nand U4460 (N_4460,N_3660,N_3736);
nor U4461 (N_4461,N_3265,N_3149);
nor U4462 (N_4462,N_3704,N_3444);
or U4463 (N_4463,N_3769,N_3926);
and U4464 (N_4464,N_3079,N_3586);
nand U4465 (N_4465,N_3969,N_3379);
nand U4466 (N_4466,N_3781,N_3172);
or U4467 (N_4467,N_3257,N_3910);
nor U4468 (N_4468,N_3785,N_3635);
nor U4469 (N_4469,N_3778,N_3633);
xnor U4470 (N_4470,N_3677,N_3934);
nand U4471 (N_4471,N_3085,N_3422);
nand U4472 (N_4472,N_3120,N_3001);
nor U4473 (N_4473,N_3141,N_3977);
nand U4474 (N_4474,N_3927,N_3583);
nand U4475 (N_4475,N_3881,N_3294);
xnor U4476 (N_4476,N_3340,N_3636);
and U4477 (N_4477,N_3908,N_3450);
nand U4478 (N_4478,N_3940,N_3937);
or U4479 (N_4479,N_3912,N_3512);
and U4480 (N_4480,N_3322,N_3464);
or U4481 (N_4481,N_3836,N_3053);
nand U4482 (N_4482,N_3022,N_3942);
nand U4483 (N_4483,N_3548,N_3055);
nand U4484 (N_4484,N_3554,N_3911);
nand U4485 (N_4485,N_3193,N_3045);
nand U4486 (N_4486,N_3596,N_3143);
nor U4487 (N_4487,N_3348,N_3297);
and U4488 (N_4488,N_3429,N_3334);
xnor U4489 (N_4489,N_3513,N_3028);
or U4490 (N_4490,N_3256,N_3381);
nand U4491 (N_4491,N_3647,N_3343);
and U4492 (N_4492,N_3525,N_3160);
nand U4493 (N_4493,N_3162,N_3812);
and U4494 (N_4494,N_3254,N_3013);
or U4495 (N_4495,N_3599,N_3224);
and U4496 (N_4496,N_3539,N_3601);
or U4497 (N_4497,N_3618,N_3810);
nand U4498 (N_4498,N_3679,N_3501);
or U4499 (N_4499,N_3988,N_3101);
xor U4500 (N_4500,N_3698,N_3167);
and U4501 (N_4501,N_3779,N_3067);
nand U4502 (N_4502,N_3585,N_3536);
nor U4503 (N_4503,N_3070,N_3232);
or U4504 (N_4504,N_3817,N_3610);
nand U4505 (N_4505,N_3756,N_3147);
nand U4506 (N_4506,N_3776,N_3710);
or U4507 (N_4507,N_3759,N_3498);
or U4508 (N_4508,N_3054,N_3466);
and U4509 (N_4509,N_3089,N_3037);
nand U4510 (N_4510,N_3169,N_3437);
or U4511 (N_4511,N_3174,N_3860);
or U4512 (N_4512,N_3009,N_3943);
xor U4513 (N_4513,N_3360,N_3025);
xor U4514 (N_4514,N_3016,N_3436);
nand U4515 (N_4515,N_3854,N_3831);
or U4516 (N_4516,N_3890,N_3644);
nand U4517 (N_4517,N_3349,N_3460);
and U4518 (N_4518,N_3008,N_3242);
nand U4519 (N_4519,N_3747,N_3438);
nand U4520 (N_4520,N_3986,N_3928);
xor U4521 (N_4521,N_3102,N_3520);
and U4522 (N_4522,N_3475,N_3768);
or U4523 (N_4523,N_3315,N_3834);
or U4524 (N_4524,N_3561,N_3832);
xnor U4525 (N_4525,N_3818,N_3110);
or U4526 (N_4526,N_3977,N_3640);
nand U4527 (N_4527,N_3709,N_3377);
and U4528 (N_4528,N_3394,N_3039);
nor U4529 (N_4529,N_3880,N_3784);
and U4530 (N_4530,N_3621,N_3236);
nor U4531 (N_4531,N_3746,N_3014);
nand U4532 (N_4532,N_3403,N_3646);
xor U4533 (N_4533,N_3540,N_3575);
or U4534 (N_4534,N_3022,N_3213);
nor U4535 (N_4535,N_3772,N_3964);
or U4536 (N_4536,N_3354,N_3966);
nand U4537 (N_4537,N_3962,N_3118);
nand U4538 (N_4538,N_3174,N_3351);
nand U4539 (N_4539,N_3183,N_3471);
nor U4540 (N_4540,N_3778,N_3963);
nand U4541 (N_4541,N_3378,N_3557);
and U4542 (N_4542,N_3302,N_3389);
or U4543 (N_4543,N_3211,N_3944);
nand U4544 (N_4544,N_3535,N_3653);
or U4545 (N_4545,N_3493,N_3295);
nor U4546 (N_4546,N_3801,N_3827);
or U4547 (N_4547,N_3778,N_3035);
nor U4548 (N_4548,N_3728,N_3893);
xor U4549 (N_4549,N_3793,N_3501);
nor U4550 (N_4550,N_3887,N_3930);
nand U4551 (N_4551,N_3020,N_3891);
and U4552 (N_4552,N_3293,N_3099);
nand U4553 (N_4553,N_3667,N_3492);
and U4554 (N_4554,N_3017,N_3436);
nand U4555 (N_4555,N_3713,N_3700);
and U4556 (N_4556,N_3978,N_3696);
nand U4557 (N_4557,N_3909,N_3476);
and U4558 (N_4558,N_3439,N_3804);
or U4559 (N_4559,N_3400,N_3195);
xnor U4560 (N_4560,N_3164,N_3877);
or U4561 (N_4561,N_3020,N_3222);
or U4562 (N_4562,N_3571,N_3866);
nand U4563 (N_4563,N_3052,N_3600);
or U4564 (N_4564,N_3990,N_3154);
and U4565 (N_4565,N_3709,N_3688);
nand U4566 (N_4566,N_3072,N_3111);
or U4567 (N_4567,N_3768,N_3160);
nand U4568 (N_4568,N_3371,N_3078);
nor U4569 (N_4569,N_3343,N_3517);
and U4570 (N_4570,N_3252,N_3342);
nand U4571 (N_4571,N_3578,N_3164);
xor U4572 (N_4572,N_3911,N_3835);
and U4573 (N_4573,N_3196,N_3329);
nand U4574 (N_4574,N_3728,N_3493);
xor U4575 (N_4575,N_3919,N_3697);
nor U4576 (N_4576,N_3996,N_3696);
nor U4577 (N_4577,N_3829,N_3105);
and U4578 (N_4578,N_3927,N_3874);
and U4579 (N_4579,N_3326,N_3073);
nor U4580 (N_4580,N_3332,N_3367);
nor U4581 (N_4581,N_3430,N_3012);
nand U4582 (N_4582,N_3845,N_3871);
or U4583 (N_4583,N_3781,N_3908);
or U4584 (N_4584,N_3889,N_3477);
and U4585 (N_4585,N_3272,N_3005);
nor U4586 (N_4586,N_3902,N_3164);
xor U4587 (N_4587,N_3599,N_3297);
xnor U4588 (N_4588,N_3714,N_3594);
or U4589 (N_4589,N_3925,N_3581);
or U4590 (N_4590,N_3170,N_3414);
and U4591 (N_4591,N_3788,N_3154);
and U4592 (N_4592,N_3038,N_3552);
and U4593 (N_4593,N_3857,N_3522);
and U4594 (N_4594,N_3694,N_3621);
and U4595 (N_4595,N_3733,N_3552);
and U4596 (N_4596,N_3367,N_3019);
or U4597 (N_4597,N_3678,N_3558);
or U4598 (N_4598,N_3939,N_3224);
or U4599 (N_4599,N_3312,N_3333);
and U4600 (N_4600,N_3575,N_3082);
and U4601 (N_4601,N_3277,N_3888);
nor U4602 (N_4602,N_3603,N_3136);
and U4603 (N_4603,N_3952,N_3079);
xor U4604 (N_4604,N_3056,N_3861);
nor U4605 (N_4605,N_3716,N_3344);
and U4606 (N_4606,N_3753,N_3805);
nor U4607 (N_4607,N_3668,N_3149);
nor U4608 (N_4608,N_3499,N_3241);
and U4609 (N_4609,N_3718,N_3431);
nand U4610 (N_4610,N_3221,N_3058);
nor U4611 (N_4611,N_3355,N_3567);
nand U4612 (N_4612,N_3050,N_3469);
or U4613 (N_4613,N_3789,N_3763);
and U4614 (N_4614,N_3921,N_3007);
and U4615 (N_4615,N_3257,N_3362);
nand U4616 (N_4616,N_3634,N_3341);
nor U4617 (N_4617,N_3711,N_3149);
nor U4618 (N_4618,N_3449,N_3277);
nor U4619 (N_4619,N_3159,N_3969);
nor U4620 (N_4620,N_3628,N_3517);
or U4621 (N_4621,N_3460,N_3906);
and U4622 (N_4622,N_3382,N_3566);
and U4623 (N_4623,N_3578,N_3518);
nand U4624 (N_4624,N_3504,N_3827);
xnor U4625 (N_4625,N_3035,N_3962);
and U4626 (N_4626,N_3691,N_3509);
or U4627 (N_4627,N_3653,N_3493);
or U4628 (N_4628,N_3266,N_3552);
nor U4629 (N_4629,N_3168,N_3463);
nand U4630 (N_4630,N_3178,N_3116);
or U4631 (N_4631,N_3231,N_3273);
nand U4632 (N_4632,N_3521,N_3074);
or U4633 (N_4633,N_3914,N_3537);
or U4634 (N_4634,N_3085,N_3273);
and U4635 (N_4635,N_3492,N_3622);
nor U4636 (N_4636,N_3909,N_3159);
xor U4637 (N_4637,N_3321,N_3012);
nor U4638 (N_4638,N_3819,N_3844);
nor U4639 (N_4639,N_3883,N_3958);
or U4640 (N_4640,N_3875,N_3034);
xnor U4641 (N_4641,N_3048,N_3378);
nand U4642 (N_4642,N_3709,N_3486);
xor U4643 (N_4643,N_3948,N_3097);
or U4644 (N_4644,N_3561,N_3254);
nand U4645 (N_4645,N_3269,N_3652);
nand U4646 (N_4646,N_3345,N_3041);
nand U4647 (N_4647,N_3797,N_3287);
or U4648 (N_4648,N_3710,N_3521);
xor U4649 (N_4649,N_3631,N_3772);
or U4650 (N_4650,N_3566,N_3092);
and U4651 (N_4651,N_3333,N_3265);
nor U4652 (N_4652,N_3511,N_3528);
and U4653 (N_4653,N_3124,N_3290);
nand U4654 (N_4654,N_3013,N_3815);
nand U4655 (N_4655,N_3935,N_3793);
xor U4656 (N_4656,N_3396,N_3958);
nor U4657 (N_4657,N_3579,N_3619);
or U4658 (N_4658,N_3099,N_3929);
or U4659 (N_4659,N_3009,N_3648);
nand U4660 (N_4660,N_3864,N_3494);
nor U4661 (N_4661,N_3074,N_3595);
nand U4662 (N_4662,N_3834,N_3313);
nor U4663 (N_4663,N_3635,N_3520);
nor U4664 (N_4664,N_3199,N_3701);
or U4665 (N_4665,N_3377,N_3606);
nand U4666 (N_4666,N_3928,N_3627);
xnor U4667 (N_4667,N_3287,N_3982);
nor U4668 (N_4668,N_3198,N_3350);
nand U4669 (N_4669,N_3217,N_3150);
or U4670 (N_4670,N_3426,N_3629);
xor U4671 (N_4671,N_3481,N_3468);
xnor U4672 (N_4672,N_3663,N_3865);
xnor U4673 (N_4673,N_3967,N_3642);
nand U4674 (N_4674,N_3627,N_3990);
xnor U4675 (N_4675,N_3213,N_3696);
nor U4676 (N_4676,N_3850,N_3190);
or U4677 (N_4677,N_3641,N_3602);
nand U4678 (N_4678,N_3404,N_3069);
and U4679 (N_4679,N_3129,N_3244);
xor U4680 (N_4680,N_3799,N_3716);
or U4681 (N_4681,N_3117,N_3107);
nand U4682 (N_4682,N_3823,N_3745);
nor U4683 (N_4683,N_3393,N_3784);
xor U4684 (N_4684,N_3967,N_3356);
and U4685 (N_4685,N_3451,N_3535);
nand U4686 (N_4686,N_3822,N_3697);
nand U4687 (N_4687,N_3140,N_3854);
or U4688 (N_4688,N_3979,N_3667);
nand U4689 (N_4689,N_3340,N_3472);
or U4690 (N_4690,N_3706,N_3716);
or U4691 (N_4691,N_3081,N_3635);
nor U4692 (N_4692,N_3683,N_3819);
xor U4693 (N_4693,N_3428,N_3276);
nor U4694 (N_4694,N_3971,N_3156);
nor U4695 (N_4695,N_3165,N_3914);
xor U4696 (N_4696,N_3028,N_3766);
xor U4697 (N_4697,N_3759,N_3365);
or U4698 (N_4698,N_3041,N_3530);
or U4699 (N_4699,N_3434,N_3143);
and U4700 (N_4700,N_3996,N_3786);
nand U4701 (N_4701,N_3165,N_3541);
xor U4702 (N_4702,N_3301,N_3320);
and U4703 (N_4703,N_3471,N_3533);
or U4704 (N_4704,N_3424,N_3118);
nand U4705 (N_4705,N_3980,N_3823);
nand U4706 (N_4706,N_3415,N_3602);
nand U4707 (N_4707,N_3256,N_3755);
nor U4708 (N_4708,N_3422,N_3821);
and U4709 (N_4709,N_3112,N_3792);
nand U4710 (N_4710,N_3892,N_3865);
nor U4711 (N_4711,N_3120,N_3497);
nor U4712 (N_4712,N_3668,N_3228);
nor U4713 (N_4713,N_3022,N_3331);
nand U4714 (N_4714,N_3303,N_3634);
nor U4715 (N_4715,N_3092,N_3057);
nand U4716 (N_4716,N_3798,N_3032);
or U4717 (N_4717,N_3669,N_3443);
nor U4718 (N_4718,N_3215,N_3943);
nand U4719 (N_4719,N_3665,N_3068);
nand U4720 (N_4720,N_3199,N_3016);
xor U4721 (N_4721,N_3126,N_3596);
or U4722 (N_4722,N_3357,N_3981);
and U4723 (N_4723,N_3545,N_3444);
and U4724 (N_4724,N_3745,N_3283);
and U4725 (N_4725,N_3436,N_3662);
and U4726 (N_4726,N_3252,N_3771);
and U4727 (N_4727,N_3825,N_3706);
nand U4728 (N_4728,N_3462,N_3862);
nor U4729 (N_4729,N_3284,N_3092);
nor U4730 (N_4730,N_3260,N_3943);
or U4731 (N_4731,N_3448,N_3379);
or U4732 (N_4732,N_3475,N_3942);
nand U4733 (N_4733,N_3987,N_3919);
nand U4734 (N_4734,N_3141,N_3612);
nor U4735 (N_4735,N_3578,N_3947);
or U4736 (N_4736,N_3370,N_3638);
and U4737 (N_4737,N_3333,N_3247);
xor U4738 (N_4738,N_3511,N_3914);
nand U4739 (N_4739,N_3862,N_3509);
nand U4740 (N_4740,N_3784,N_3161);
nand U4741 (N_4741,N_3558,N_3423);
nand U4742 (N_4742,N_3284,N_3659);
nor U4743 (N_4743,N_3123,N_3033);
and U4744 (N_4744,N_3300,N_3028);
nand U4745 (N_4745,N_3272,N_3768);
or U4746 (N_4746,N_3219,N_3349);
nor U4747 (N_4747,N_3885,N_3681);
or U4748 (N_4748,N_3639,N_3454);
nor U4749 (N_4749,N_3198,N_3232);
nand U4750 (N_4750,N_3461,N_3653);
nor U4751 (N_4751,N_3013,N_3128);
or U4752 (N_4752,N_3655,N_3203);
xor U4753 (N_4753,N_3412,N_3033);
or U4754 (N_4754,N_3709,N_3323);
and U4755 (N_4755,N_3865,N_3684);
nor U4756 (N_4756,N_3872,N_3026);
nor U4757 (N_4757,N_3147,N_3419);
nor U4758 (N_4758,N_3923,N_3981);
or U4759 (N_4759,N_3839,N_3630);
and U4760 (N_4760,N_3701,N_3289);
or U4761 (N_4761,N_3866,N_3453);
nor U4762 (N_4762,N_3921,N_3013);
nor U4763 (N_4763,N_3289,N_3919);
or U4764 (N_4764,N_3380,N_3628);
nor U4765 (N_4765,N_3697,N_3535);
nor U4766 (N_4766,N_3208,N_3770);
or U4767 (N_4767,N_3121,N_3385);
and U4768 (N_4768,N_3518,N_3887);
and U4769 (N_4769,N_3175,N_3527);
or U4770 (N_4770,N_3079,N_3529);
nand U4771 (N_4771,N_3448,N_3497);
xor U4772 (N_4772,N_3591,N_3300);
nor U4773 (N_4773,N_3552,N_3904);
nand U4774 (N_4774,N_3663,N_3421);
or U4775 (N_4775,N_3832,N_3728);
nand U4776 (N_4776,N_3236,N_3847);
or U4777 (N_4777,N_3094,N_3050);
nand U4778 (N_4778,N_3951,N_3658);
nor U4779 (N_4779,N_3136,N_3865);
nand U4780 (N_4780,N_3526,N_3160);
nand U4781 (N_4781,N_3784,N_3611);
xnor U4782 (N_4782,N_3088,N_3489);
nor U4783 (N_4783,N_3896,N_3527);
nand U4784 (N_4784,N_3765,N_3424);
nor U4785 (N_4785,N_3019,N_3419);
nand U4786 (N_4786,N_3054,N_3083);
or U4787 (N_4787,N_3525,N_3814);
nand U4788 (N_4788,N_3873,N_3815);
or U4789 (N_4789,N_3073,N_3313);
or U4790 (N_4790,N_3566,N_3142);
xnor U4791 (N_4791,N_3001,N_3945);
nor U4792 (N_4792,N_3113,N_3245);
xnor U4793 (N_4793,N_3317,N_3454);
or U4794 (N_4794,N_3281,N_3985);
nor U4795 (N_4795,N_3506,N_3368);
nor U4796 (N_4796,N_3170,N_3095);
nor U4797 (N_4797,N_3899,N_3826);
and U4798 (N_4798,N_3337,N_3586);
or U4799 (N_4799,N_3320,N_3025);
nand U4800 (N_4800,N_3708,N_3179);
nand U4801 (N_4801,N_3468,N_3164);
nor U4802 (N_4802,N_3539,N_3566);
or U4803 (N_4803,N_3173,N_3040);
nand U4804 (N_4804,N_3878,N_3265);
and U4805 (N_4805,N_3221,N_3709);
and U4806 (N_4806,N_3330,N_3440);
or U4807 (N_4807,N_3411,N_3322);
or U4808 (N_4808,N_3885,N_3008);
and U4809 (N_4809,N_3663,N_3324);
and U4810 (N_4810,N_3275,N_3212);
and U4811 (N_4811,N_3993,N_3315);
or U4812 (N_4812,N_3205,N_3542);
xnor U4813 (N_4813,N_3470,N_3432);
nand U4814 (N_4814,N_3386,N_3725);
nor U4815 (N_4815,N_3427,N_3599);
and U4816 (N_4816,N_3029,N_3759);
nand U4817 (N_4817,N_3083,N_3033);
or U4818 (N_4818,N_3947,N_3768);
or U4819 (N_4819,N_3042,N_3615);
nand U4820 (N_4820,N_3098,N_3032);
and U4821 (N_4821,N_3450,N_3304);
nand U4822 (N_4822,N_3193,N_3935);
and U4823 (N_4823,N_3098,N_3075);
nor U4824 (N_4824,N_3851,N_3247);
nand U4825 (N_4825,N_3837,N_3668);
xnor U4826 (N_4826,N_3858,N_3599);
nand U4827 (N_4827,N_3742,N_3556);
and U4828 (N_4828,N_3002,N_3635);
nand U4829 (N_4829,N_3949,N_3502);
nor U4830 (N_4830,N_3391,N_3303);
and U4831 (N_4831,N_3216,N_3316);
nor U4832 (N_4832,N_3577,N_3586);
and U4833 (N_4833,N_3217,N_3121);
or U4834 (N_4834,N_3567,N_3315);
nor U4835 (N_4835,N_3803,N_3792);
and U4836 (N_4836,N_3512,N_3997);
nand U4837 (N_4837,N_3313,N_3163);
or U4838 (N_4838,N_3389,N_3488);
nor U4839 (N_4839,N_3258,N_3645);
nand U4840 (N_4840,N_3559,N_3891);
or U4841 (N_4841,N_3996,N_3524);
nand U4842 (N_4842,N_3609,N_3883);
and U4843 (N_4843,N_3928,N_3541);
and U4844 (N_4844,N_3789,N_3455);
nand U4845 (N_4845,N_3330,N_3980);
and U4846 (N_4846,N_3480,N_3932);
nand U4847 (N_4847,N_3676,N_3545);
nand U4848 (N_4848,N_3787,N_3892);
and U4849 (N_4849,N_3580,N_3180);
xnor U4850 (N_4850,N_3484,N_3926);
nand U4851 (N_4851,N_3561,N_3100);
xor U4852 (N_4852,N_3219,N_3913);
nor U4853 (N_4853,N_3536,N_3911);
nand U4854 (N_4854,N_3274,N_3509);
nand U4855 (N_4855,N_3719,N_3299);
xnor U4856 (N_4856,N_3545,N_3852);
nor U4857 (N_4857,N_3859,N_3409);
nand U4858 (N_4858,N_3884,N_3381);
nor U4859 (N_4859,N_3428,N_3423);
and U4860 (N_4860,N_3015,N_3953);
nor U4861 (N_4861,N_3146,N_3128);
and U4862 (N_4862,N_3520,N_3527);
and U4863 (N_4863,N_3348,N_3691);
nand U4864 (N_4864,N_3954,N_3229);
nor U4865 (N_4865,N_3754,N_3341);
and U4866 (N_4866,N_3244,N_3937);
xnor U4867 (N_4867,N_3028,N_3850);
xnor U4868 (N_4868,N_3255,N_3459);
nand U4869 (N_4869,N_3109,N_3964);
nor U4870 (N_4870,N_3538,N_3071);
or U4871 (N_4871,N_3766,N_3213);
or U4872 (N_4872,N_3972,N_3394);
nand U4873 (N_4873,N_3611,N_3106);
or U4874 (N_4874,N_3114,N_3646);
and U4875 (N_4875,N_3238,N_3442);
nand U4876 (N_4876,N_3417,N_3804);
or U4877 (N_4877,N_3611,N_3750);
nand U4878 (N_4878,N_3286,N_3294);
nand U4879 (N_4879,N_3359,N_3334);
nand U4880 (N_4880,N_3127,N_3735);
and U4881 (N_4881,N_3806,N_3413);
nand U4882 (N_4882,N_3463,N_3900);
or U4883 (N_4883,N_3765,N_3730);
and U4884 (N_4884,N_3366,N_3276);
and U4885 (N_4885,N_3621,N_3875);
and U4886 (N_4886,N_3311,N_3213);
or U4887 (N_4887,N_3691,N_3979);
and U4888 (N_4888,N_3615,N_3351);
nor U4889 (N_4889,N_3713,N_3099);
nor U4890 (N_4890,N_3026,N_3907);
nand U4891 (N_4891,N_3333,N_3262);
nor U4892 (N_4892,N_3507,N_3329);
nor U4893 (N_4893,N_3779,N_3276);
and U4894 (N_4894,N_3213,N_3627);
or U4895 (N_4895,N_3136,N_3470);
or U4896 (N_4896,N_3577,N_3596);
or U4897 (N_4897,N_3181,N_3798);
or U4898 (N_4898,N_3212,N_3691);
nor U4899 (N_4899,N_3618,N_3258);
nor U4900 (N_4900,N_3759,N_3240);
nand U4901 (N_4901,N_3039,N_3307);
and U4902 (N_4902,N_3414,N_3791);
nor U4903 (N_4903,N_3672,N_3010);
nand U4904 (N_4904,N_3353,N_3025);
nor U4905 (N_4905,N_3553,N_3233);
nor U4906 (N_4906,N_3474,N_3948);
and U4907 (N_4907,N_3726,N_3523);
or U4908 (N_4908,N_3676,N_3196);
nor U4909 (N_4909,N_3255,N_3854);
nand U4910 (N_4910,N_3107,N_3751);
nand U4911 (N_4911,N_3689,N_3050);
nand U4912 (N_4912,N_3211,N_3515);
nor U4913 (N_4913,N_3533,N_3688);
or U4914 (N_4914,N_3145,N_3006);
nor U4915 (N_4915,N_3746,N_3307);
and U4916 (N_4916,N_3270,N_3567);
or U4917 (N_4917,N_3014,N_3458);
xor U4918 (N_4918,N_3124,N_3817);
nand U4919 (N_4919,N_3965,N_3154);
nor U4920 (N_4920,N_3369,N_3379);
nor U4921 (N_4921,N_3531,N_3737);
and U4922 (N_4922,N_3250,N_3407);
nand U4923 (N_4923,N_3850,N_3243);
nand U4924 (N_4924,N_3811,N_3986);
nand U4925 (N_4925,N_3250,N_3472);
nand U4926 (N_4926,N_3327,N_3772);
and U4927 (N_4927,N_3385,N_3618);
nor U4928 (N_4928,N_3375,N_3545);
nand U4929 (N_4929,N_3499,N_3610);
nand U4930 (N_4930,N_3896,N_3064);
nand U4931 (N_4931,N_3726,N_3594);
and U4932 (N_4932,N_3982,N_3849);
nand U4933 (N_4933,N_3311,N_3664);
or U4934 (N_4934,N_3470,N_3190);
nor U4935 (N_4935,N_3184,N_3775);
nand U4936 (N_4936,N_3744,N_3772);
nor U4937 (N_4937,N_3206,N_3029);
nand U4938 (N_4938,N_3016,N_3032);
nor U4939 (N_4939,N_3472,N_3379);
and U4940 (N_4940,N_3228,N_3384);
nor U4941 (N_4941,N_3777,N_3406);
nand U4942 (N_4942,N_3264,N_3962);
nor U4943 (N_4943,N_3846,N_3556);
nand U4944 (N_4944,N_3092,N_3777);
nand U4945 (N_4945,N_3263,N_3591);
nor U4946 (N_4946,N_3700,N_3555);
nand U4947 (N_4947,N_3974,N_3854);
xnor U4948 (N_4948,N_3881,N_3687);
or U4949 (N_4949,N_3467,N_3590);
xnor U4950 (N_4950,N_3858,N_3268);
and U4951 (N_4951,N_3921,N_3395);
and U4952 (N_4952,N_3100,N_3754);
and U4953 (N_4953,N_3884,N_3793);
or U4954 (N_4954,N_3682,N_3817);
nand U4955 (N_4955,N_3272,N_3353);
nor U4956 (N_4956,N_3825,N_3798);
and U4957 (N_4957,N_3114,N_3682);
or U4958 (N_4958,N_3454,N_3042);
nand U4959 (N_4959,N_3647,N_3774);
nor U4960 (N_4960,N_3415,N_3230);
nor U4961 (N_4961,N_3404,N_3519);
nor U4962 (N_4962,N_3315,N_3251);
xnor U4963 (N_4963,N_3679,N_3652);
nor U4964 (N_4964,N_3854,N_3126);
and U4965 (N_4965,N_3642,N_3942);
nor U4966 (N_4966,N_3835,N_3315);
nor U4967 (N_4967,N_3506,N_3451);
nor U4968 (N_4968,N_3425,N_3130);
nor U4969 (N_4969,N_3460,N_3562);
and U4970 (N_4970,N_3547,N_3834);
or U4971 (N_4971,N_3002,N_3883);
and U4972 (N_4972,N_3619,N_3289);
xnor U4973 (N_4973,N_3319,N_3789);
and U4974 (N_4974,N_3004,N_3725);
and U4975 (N_4975,N_3794,N_3072);
nor U4976 (N_4976,N_3557,N_3448);
and U4977 (N_4977,N_3572,N_3442);
nor U4978 (N_4978,N_3508,N_3783);
nor U4979 (N_4979,N_3878,N_3548);
xor U4980 (N_4980,N_3430,N_3543);
or U4981 (N_4981,N_3528,N_3748);
and U4982 (N_4982,N_3659,N_3095);
and U4983 (N_4983,N_3638,N_3840);
and U4984 (N_4984,N_3627,N_3466);
nor U4985 (N_4985,N_3779,N_3789);
nand U4986 (N_4986,N_3854,N_3918);
nor U4987 (N_4987,N_3491,N_3722);
and U4988 (N_4988,N_3846,N_3169);
or U4989 (N_4989,N_3212,N_3453);
xor U4990 (N_4990,N_3233,N_3697);
xor U4991 (N_4991,N_3313,N_3640);
nand U4992 (N_4992,N_3349,N_3261);
and U4993 (N_4993,N_3590,N_3493);
nor U4994 (N_4994,N_3397,N_3251);
or U4995 (N_4995,N_3751,N_3363);
nor U4996 (N_4996,N_3543,N_3313);
or U4997 (N_4997,N_3524,N_3731);
and U4998 (N_4998,N_3567,N_3913);
nand U4999 (N_4999,N_3235,N_3567);
or U5000 (N_5000,N_4597,N_4742);
nand U5001 (N_5001,N_4646,N_4239);
nor U5002 (N_5002,N_4483,N_4756);
xnor U5003 (N_5003,N_4576,N_4023);
or U5004 (N_5004,N_4031,N_4780);
nor U5005 (N_5005,N_4809,N_4220);
or U5006 (N_5006,N_4366,N_4301);
nor U5007 (N_5007,N_4029,N_4424);
or U5008 (N_5008,N_4464,N_4553);
xor U5009 (N_5009,N_4984,N_4952);
nand U5010 (N_5010,N_4787,N_4891);
nand U5011 (N_5011,N_4371,N_4907);
or U5012 (N_5012,N_4234,N_4453);
xnor U5013 (N_5013,N_4916,N_4449);
and U5014 (N_5014,N_4428,N_4688);
or U5015 (N_5015,N_4647,N_4425);
nand U5016 (N_5016,N_4141,N_4888);
xor U5017 (N_5017,N_4030,N_4755);
nand U5018 (N_5018,N_4667,N_4716);
nand U5019 (N_5019,N_4648,N_4185);
and U5020 (N_5020,N_4217,N_4108);
and U5021 (N_5021,N_4462,N_4434);
nand U5022 (N_5022,N_4624,N_4327);
and U5023 (N_5023,N_4680,N_4718);
or U5024 (N_5024,N_4993,N_4207);
nor U5025 (N_5025,N_4033,N_4825);
nand U5026 (N_5026,N_4697,N_4078);
or U5027 (N_5027,N_4244,N_4886);
and U5028 (N_5028,N_4728,N_4457);
and U5029 (N_5029,N_4087,N_4757);
nor U5030 (N_5030,N_4972,N_4329);
and U5031 (N_5031,N_4067,N_4016);
nor U5032 (N_5032,N_4867,N_4089);
and U5033 (N_5033,N_4395,N_4843);
and U5034 (N_5034,N_4403,N_4857);
nand U5035 (N_5035,N_4130,N_4817);
nand U5036 (N_5036,N_4397,N_4662);
nor U5037 (N_5037,N_4213,N_4171);
nand U5038 (N_5038,N_4512,N_4791);
or U5039 (N_5039,N_4333,N_4987);
nor U5040 (N_5040,N_4992,N_4900);
nor U5041 (N_5041,N_4518,N_4298);
and U5042 (N_5042,N_4111,N_4883);
nor U5043 (N_5043,N_4710,N_4632);
and U5044 (N_5044,N_4418,N_4775);
nand U5045 (N_5045,N_4488,N_4516);
or U5046 (N_5046,N_4440,N_4915);
or U5047 (N_5047,N_4392,N_4898);
nand U5048 (N_5048,N_4194,N_4102);
nor U5049 (N_5049,N_4943,N_4572);
or U5050 (N_5050,N_4228,N_4508);
and U5051 (N_5051,N_4426,N_4567);
xor U5052 (N_5052,N_4681,N_4538);
or U5053 (N_5053,N_4455,N_4798);
xnor U5054 (N_5054,N_4138,N_4838);
nor U5055 (N_5055,N_4153,N_4621);
and U5056 (N_5056,N_4677,N_4314);
xnor U5057 (N_5057,N_4629,N_4924);
nand U5058 (N_5058,N_4357,N_4316);
nor U5059 (N_5059,N_4676,N_4476);
and U5060 (N_5060,N_4570,N_4223);
or U5061 (N_5061,N_4154,N_4054);
and U5062 (N_5062,N_4837,N_4671);
nand U5063 (N_5063,N_4747,N_4580);
nand U5064 (N_5064,N_4431,N_4152);
nand U5065 (N_5065,N_4276,N_4783);
nand U5066 (N_5066,N_4880,N_4986);
nor U5067 (N_5067,N_4255,N_4715);
nand U5068 (N_5068,N_4432,N_4699);
nand U5069 (N_5069,N_4170,N_4313);
or U5070 (N_5070,N_4399,N_4912);
nand U5071 (N_5071,N_4723,N_4807);
or U5072 (N_5072,N_4147,N_4132);
xor U5073 (N_5073,N_4413,N_4534);
nor U5074 (N_5074,N_4633,N_4811);
or U5075 (N_5075,N_4969,N_4705);
xnor U5076 (N_5076,N_4332,N_4919);
nor U5077 (N_5077,N_4639,N_4539);
nor U5078 (N_5078,N_4674,N_4012);
and U5079 (N_5079,N_4139,N_4335);
nand U5080 (N_5080,N_4252,N_4872);
or U5081 (N_5081,N_4182,N_4010);
nand U5082 (N_5082,N_4394,N_4473);
or U5083 (N_5083,N_4577,N_4061);
nand U5084 (N_5084,N_4794,N_4272);
nand U5085 (N_5085,N_4180,N_4211);
or U5086 (N_5086,N_4804,N_4035);
nor U5087 (N_5087,N_4582,N_4007);
or U5088 (N_5088,N_4616,N_4364);
nand U5089 (N_5089,N_4446,N_4941);
and U5090 (N_5090,N_4748,N_4469);
nand U5091 (N_5091,N_4776,N_4527);
and U5092 (N_5092,N_4528,N_4732);
nand U5093 (N_5093,N_4878,N_4140);
and U5094 (N_5094,N_4810,N_4247);
xnor U5095 (N_5095,N_4549,N_4183);
nand U5096 (N_5096,N_4300,N_4053);
nand U5097 (N_5097,N_4841,N_4753);
xnor U5098 (N_5098,N_4558,N_4369);
nand U5099 (N_5099,N_4655,N_4853);
nor U5100 (N_5100,N_4261,N_4556);
or U5101 (N_5101,N_4450,N_4096);
xor U5102 (N_5102,N_4926,N_4103);
xnor U5103 (N_5103,N_4965,N_4229);
nand U5104 (N_5104,N_4289,N_4610);
or U5105 (N_5105,N_4977,N_4295);
and U5106 (N_5106,N_4828,N_4186);
or U5107 (N_5107,N_4782,N_4842);
or U5108 (N_5108,N_4873,N_4573);
and U5109 (N_5109,N_4487,N_4443);
nand U5110 (N_5110,N_4378,N_4064);
or U5111 (N_5111,N_4981,N_4870);
nand U5112 (N_5112,N_4197,N_4649);
or U5113 (N_5113,N_4059,N_4806);
and U5114 (N_5114,N_4419,N_4686);
and U5115 (N_5115,N_4945,N_4998);
nand U5116 (N_5116,N_4060,N_4687);
xnor U5117 (N_5117,N_4899,N_4179);
and U5118 (N_5118,N_4934,N_4693);
nand U5119 (N_5119,N_4133,N_4859);
nor U5120 (N_5120,N_4684,N_4833);
xor U5121 (N_5121,N_4043,N_4526);
and U5122 (N_5122,N_4956,N_4156);
or U5123 (N_5123,N_4374,N_4409);
xnor U5124 (N_5124,N_4122,N_4422);
or U5125 (N_5125,N_4190,N_4381);
nor U5126 (N_5126,N_4675,N_4321);
or U5127 (N_5127,N_4968,N_4772);
or U5128 (N_5128,N_4702,N_4134);
and U5129 (N_5129,N_4442,N_4513);
or U5130 (N_5130,N_4013,N_4124);
nor U5131 (N_5131,N_4540,N_4068);
and U5132 (N_5132,N_4215,N_4493);
and U5133 (N_5133,N_4692,N_4701);
nand U5134 (N_5134,N_4104,N_4020);
nand U5135 (N_5135,N_4018,N_4354);
and U5136 (N_5136,N_4600,N_4596);
nand U5137 (N_5137,N_4401,N_4522);
and U5138 (N_5138,N_4254,N_4191);
nor U5139 (N_5139,N_4066,N_4939);
and U5140 (N_5140,N_4725,N_4002);
and U5141 (N_5141,N_4942,N_4338);
nand U5142 (N_5142,N_4330,N_4658);
nand U5143 (N_5143,N_4612,N_4601);
xor U5144 (N_5144,N_4051,N_4468);
xor U5145 (N_5145,N_4997,N_4331);
and U5146 (N_5146,N_4865,N_4232);
or U5147 (N_5147,N_4174,N_4887);
and U5148 (N_5148,N_4014,N_4685);
or U5149 (N_5149,N_4816,N_4669);
or U5150 (N_5150,N_4226,N_4980);
nor U5151 (N_5151,N_4547,N_4277);
nand U5152 (N_5152,N_4781,N_4949);
nand U5153 (N_5153,N_4559,N_4773);
nor U5154 (N_5154,N_4387,N_4678);
nor U5155 (N_5155,N_4283,N_4441);
nand U5156 (N_5156,N_4412,N_4963);
xor U5157 (N_5157,N_4703,N_4454);
or U5158 (N_5158,N_4990,N_4737);
or U5159 (N_5159,N_4599,N_4375);
nand U5160 (N_5160,N_4188,N_4829);
nand U5161 (N_5161,N_4082,N_4415);
nor U5162 (N_5162,N_4734,N_4714);
xor U5163 (N_5163,N_4458,N_4480);
xnor U5164 (N_5164,N_4263,N_4172);
and U5165 (N_5165,N_4322,N_4097);
and U5166 (N_5166,N_4584,N_4417);
nand U5167 (N_5167,N_4935,N_4490);
nand U5168 (N_5168,N_4187,N_4447);
and U5169 (N_5169,N_4511,N_4819);
and U5170 (N_5170,N_4115,N_4323);
nor U5171 (N_5171,N_4799,N_4861);
nand U5172 (N_5172,N_4712,N_4523);
or U5173 (N_5173,N_4666,N_4668);
and U5174 (N_5174,N_4940,N_4448);
nand U5175 (N_5175,N_4709,N_4656);
nor U5176 (N_5176,N_4165,N_4879);
and U5177 (N_5177,N_4000,N_4383);
nor U5178 (N_5178,N_4200,N_4273);
and U5179 (N_5179,N_4202,N_4920);
nor U5180 (N_5180,N_4292,N_4854);
nor U5181 (N_5181,N_4763,N_4199);
nor U5182 (N_5182,N_4585,N_4264);
and U5183 (N_5183,N_4575,N_4947);
nand U5184 (N_5184,N_4721,N_4856);
nand U5185 (N_5185,N_4896,N_4386);
xnor U5186 (N_5186,N_4988,N_4151);
and U5187 (N_5187,N_4451,N_4146);
and U5188 (N_5188,N_4039,N_4914);
and U5189 (N_5189,N_4076,N_4274);
or U5190 (N_5190,N_4683,N_4958);
nor U5191 (N_5191,N_4543,N_4209);
nor U5192 (N_5192,N_4704,N_4533);
nand U5193 (N_5193,N_4877,N_4938);
nor U5194 (N_5194,N_4037,N_4406);
nor U5195 (N_5195,N_4964,N_4665);
nand U5196 (N_5196,N_4243,N_4358);
or U5197 (N_5197,N_4155,N_4805);
nand U5198 (N_5198,N_4863,N_4173);
or U5199 (N_5199,N_4435,N_4720);
nand U5200 (N_5200,N_4628,N_4587);
xor U5201 (N_5201,N_4225,N_4249);
or U5202 (N_5202,N_4614,N_4080);
xnor U5203 (N_5203,N_4933,N_4074);
and U5204 (N_5204,N_4778,N_4373);
or U5205 (N_5205,N_4796,N_4869);
nand U5206 (N_5206,N_4175,N_4670);
and U5207 (N_5207,N_4660,N_4477);
nand U5208 (N_5208,N_4803,N_4478);
nand U5209 (N_5209,N_4083,N_4430);
nand U5210 (N_5210,N_4168,N_4785);
and U5211 (N_5211,N_4400,N_4729);
xnor U5212 (N_5212,N_4334,N_4315);
and U5213 (N_5213,N_4296,N_4063);
and U5214 (N_5214,N_4218,N_4834);
xnor U5215 (N_5215,N_4765,N_4137);
or U5216 (N_5216,N_4749,N_4966);
nor U5217 (N_5217,N_4895,N_4216);
nor U5218 (N_5218,N_4456,N_4820);
or U5219 (N_5219,N_4631,N_4881);
nand U5220 (N_5220,N_4005,N_4348);
nand U5221 (N_5221,N_4911,N_4241);
nand U5222 (N_5222,N_4495,N_4944);
nand U5223 (N_5223,N_4619,N_4248);
nor U5224 (N_5224,N_4630,N_4497);
or U5225 (N_5225,N_4706,N_4991);
or U5226 (N_5226,N_4955,N_4306);
nor U5227 (N_5227,N_4983,N_4740);
nand U5228 (N_5228,N_4555,N_4048);
nand U5229 (N_5229,N_4491,N_4390);
nand U5230 (N_5230,N_4563,N_4098);
nor U5231 (N_5231,N_4741,N_4717);
nor U5232 (N_5232,N_4767,N_4653);
and U5233 (N_5233,N_4069,N_4815);
nand U5234 (N_5234,N_4470,N_4282);
or U5235 (N_5235,N_4620,N_4318);
or U5236 (N_5236,N_4618,N_4024);
and U5237 (N_5237,N_4541,N_4135);
nor U5238 (N_5238,N_4797,N_4384);
nand U5239 (N_5239,N_4548,N_4546);
or U5240 (N_5240,N_4404,N_4251);
and U5241 (N_5241,N_4342,N_4351);
or U5242 (N_5242,N_4303,N_4858);
nand U5243 (N_5243,N_4913,N_4123);
nor U5244 (N_5244,N_4245,N_4967);
and U5245 (N_5245,N_4844,N_4376);
and U5246 (N_5246,N_4071,N_4627);
and U5247 (N_5247,N_4117,N_4113);
nand U5248 (N_5248,N_4906,N_4542);
nand U5249 (N_5249,N_4324,N_4948);
and U5250 (N_5250,N_4496,N_4554);
and U5251 (N_5251,N_4738,N_4144);
and U5252 (N_5252,N_4501,N_4890);
nand U5253 (N_5253,N_4161,N_4481);
and U5254 (N_5254,N_4637,N_4408);
nor U5255 (N_5255,N_4520,N_4379);
xnor U5256 (N_5256,N_4826,N_4617);
nor U5257 (N_5257,N_4325,N_4485);
or U5258 (N_5258,N_4270,N_4673);
nand U5259 (N_5259,N_4405,N_4855);
or U5260 (N_5260,N_4730,N_4482);
xnor U5261 (N_5261,N_4903,N_4586);
and U5262 (N_5262,N_4463,N_4615);
xnor U5263 (N_5263,N_4836,N_4875);
or U5264 (N_5264,N_4242,N_4902);
or U5265 (N_5265,N_4046,N_4847);
nor U5266 (N_5266,N_4982,N_4659);
nand U5267 (N_5267,N_4792,N_4827);
nand U5268 (N_5268,N_4143,N_4831);
xnor U5269 (N_5269,N_4347,N_4885);
or U5270 (N_5270,N_4205,N_4057);
nor U5271 (N_5271,N_4100,N_4294);
nor U5272 (N_5272,N_4259,N_4305);
or U5273 (N_5273,N_4689,N_4360);
and U5274 (N_5274,N_4085,N_4230);
nor U5275 (N_5275,N_4908,N_4128);
nand U5276 (N_5276,N_4075,N_4265);
nor U5277 (N_5277,N_4937,N_4638);
nand U5278 (N_5278,N_4727,N_4592);
nor U5279 (N_5279,N_4044,N_4840);
xor U5280 (N_5280,N_4994,N_4429);
nand U5281 (N_5281,N_4336,N_4866);
and U5282 (N_5282,N_4045,N_4946);
and U5283 (N_5283,N_4893,N_4250);
or U5284 (N_5284,N_4724,N_4286);
nand U5285 (N_5285,N_4041,N_4433);
or U5286 (N_5286,N_4974,N_4606);
nand U5287 (N_5287,N_4176,N_4472);
nand U5288 (N_5288,N_4396,N_4636);
nand U5289 (N_5289,N_4641,N_4850);
nor U5290 (N_5290,N_4049,N_4568);
nor U5291 (N_5291,N_4127,N_4735);
xor U5292 (N_5292,N_4611,N_4163);
nor U5293 (N_5293,N_4852,N_4500);
nand U5294 (N_5294,N_4367,N_4136);
or U5295 (N_5295,N_4790,N_4504);
nor U5296 (N_5296,N_4736,N_4452);
or U5297 (N_5297,N_4605,N_4643);
nor U5298 (N_5298,N_4445,N_4311);
or U5299 (N_5299,N_4973,N_4793);
xor U5300 (N_5300,N_4608,N_4622);
xor U5301 (N_5301,N_4438,N_4407);
and U5302 (N_5302,N_4388,N_4106);
and U5303 (N_5303,N_4253,N_4698);
or U5304 (N_5304,N_4589,N_4028);
and U5305 (N_5305,N_4789,N_4832);
or U5306 (N_5306,N_4918,N_4722);
xor U5307 (N_5307,N_4164,N_4101);
nor U5308 (N_5308,N_4532,N_4091);
nand U5309 (N_5309,N_4588,N_4571);
nor U5310 (N_5310,N_4564,N_4203);
or U5311 (N_5311,N_4084,N_4328);
nor U5312 (N_5312,N_4711,N_4466);
nand U5313 (N_5313,N_4953,N_4874);
or U5314 (N_5314,N_4979,N_4644);
and U5315 (N_5315,N_4436,N_4650);
nand U5316 (N_5316,N_4079,N_4719);
nor U5317 (N_5317,N_4235,N_4411);
and U5318 (N_5318,N_4224,N_4439);
nor U5319 (N_5319,N_4356,N_4222);
or U5320 (N_5320,N_4011,N_4524);
nor U5321 (N_5321,N_4707,N_4499);
nor U5322 (N_5322,N_4679,N_4593);
or U5323 (N_5323,N_4281,N_4365);
nand U5324 (N_5324,N_4774,N_4484);
or U5325 (N_5325,N_4999,N_4486);
and U5326 (N_5326,N_4768,N_4744);
and U5327 (N_5327,N_4110,N_4525);
nand U5328 (N_5328,N_4090,N_4910);
and U5329 (N_5329,N_4739,N_4363);
nand U5330 (N_5330,N_4019,N_4343);
nand U5331 (N_5331,N_4726,N_4795);
or U5332 (N_5332,N_4420,N_4788);
nor U5333 (N_5333,N_4536,N_4960);
and U5334 (N_5334,N_4579,N_4006);
or U5335 (N_5335,N_4801,N_4905);
nor U5336 (N_5336,N_4494,N_4131);
xnor U5337 (N_5337,N_4003,N_4625);
or U5338 (N_5338,N_4193,N_4713);
nand U5339 (N_5339,N_4545,N_4754);
and U5340 (N_5340,N_4813,N_4672);
nand U5341 (N_5341,N_4818,N_4385);
and U5342 (N_5342,N_4377,N_4574);
xor U5343 (N_5343,N_4654,N_4056);
or U5344 (N_5344,N_4690,N_4962);
and U5345 (N_5345,N_4498,N_4609);
nand U5346 (N_5346,N_4519,N_4931);
xor U5347 (N_5347,N_4970,N_4510);
and U5348 (N_5348,N_4393,N_4923);
or U5349 (N_5349,N_4214,N_4317);
nor U5350 (N_5350,N_4897,N_4359);
nor U5351 (N_5351,N_4055,N_4975);
nor U5352 (N_5352,N_4460,N_4635);
nor U5353 (N_5353,N_4350,N_4752);
or U5354 (N_5354,N_4927,N_4846);
xor U5355 (N_5355,N_4746,N_4760);
or U5356 (N_5356,N_4959,N_4038);
nand U5357 (N_5357,N_4864,N_4604);
nor U5358 (N_5358,N_4645,N_4380);
and U5359 (N_5359,N_4278,N_4557);
nand U5360 (N_5360,N_4894,N_4502);
or U5361 (N_5361,N_4786,N_4086);
nor U5362 (N_5362,N_4427,N_4109);
nand U5363 (N_5363,N_4800,N_4204);
nand U5364 (N_5364,N_4015,N_4731);
or U5365 (N_5365,N_4664,N_4227);
nor U5366 (N_5366,N_4114,N_4070);
nor U5367 (N_5367,N_4126,N_4021);
or U5368 (N_5368,N_4762,N_4565);
and U5369 (N_5369,N_4107,N_4237);
and U5370 (N_5370,N_4437,N_4093);
nor U5371 (N_5371,N_4507,N_4177);
nand U5372 (N_5372,N_4238,N_4651);
and U5373 (N_5373,N_4634,N_4416);
nand U5374 (N_5374,N_4036,N_4279);
nor U5375 (N_5375,N_4047,N_4062);
or U5376 (N_5376,N_4544,N_4976);
nor U5377 (N_5377,N_4184,N_4262);
and U5378 (N_5378,N_4052,N_4266);
nand U5379 (N_5379,N_4240,N_4909);
and U5380 (N_5380,N_4954,N_4779);
and U5381 (N_5381,N_4149,N_4219);
xnor U5382 (N_5382,N_4602,N_4862);
nor U5383 (N_5383,N_4368,N_4623);
nor U5384 (N_5384,N_4304,N_4830);
and U5385 (N_5385,N_4663,N_4148);
or U5386 (N_5386,N_4471,N_4771);
and U5387 (N_5387,N_4824,N_4694);
and U5388 (N_5388,N_4751,N_4529);
nand U5389 (N_5389,N_4201,N_4370);
or U5390 (N_5390,N_4178,N_4092);
and U5391 (N_5391,N_4917,N_4743);
nor U5392 (N_5392,N_4196,N_4515);
xnor U5393 (N_5393,N_4121,N_4221);
and U5394 (N_5394,N_4352,N_4822);
nand U5395 (N_5395,N_4835,N_4299);
nor U5396 (N_5396,N_4157,N_4319);
and U5397 (N_5397,N_4034,N_4192);
nor U5398 (N_5398,N_4882,N_4506);
nand U5399 (N_5399,N_4361,N_4957);
nand U5400 (N_5400,N_4246,N_4509);
nor U5401 (N_5401,N_4355,N_4167);
nand U5402 (N_5402,N_4026,N_4088);
xnor U5403 (N_5403,N_4236,N_4022);
or U5404 (N_5404,N_4868,N_4372);
nor U5405 (N_5405,N_4904,N_4849);
nor U5406 (N_5406,N_4339,N_4142);
nand U5407 (N_5407,N_4581,N_4072);
or U5408 (N_5408,N_4695,N_4065);
nand U5409 (N_5409,N_4901,N_4337);
nand U5410 (N_5410,N_4613,N_4421);
and U5411 (N_5411,N_4349,N_4821);
and U5412 (N_5412,N_4884,N_4233);
and U5413 (N_5413,N_4257,N_4591);
xnor U5414 (N_5414,N_4040,N_4118);
nor U5415 (N_5415,N_4465,N_4008);
xor U5416 (N_5416,N_4297,N_4308);
nand U5417 (N_5417,N_4626,N_4761);
xnor U5418 (N_5418,N_4708,N_4640);
nand U5419 (N_5419,N_4733,N_4770);
and U5420 (N_5420,N_4661,N_4961);
and U5421 (N_5421,N_4551,N_4745);
nand U5422 (N_5422,N_4206,N_4461);
nand U5423 (N_5423,N_4258,N_4150);
nor U5424 (N_5424,N_4459,N_4848);
or U5425 (N_5425,N_4985,N_4081);
and U5426 (N_5426,N_4530,N_4537);
nor U5427 (N_5427,N_4758,N_4391);
and U5428 (N_5428,N_4777,N_4845);
xor U5429 (N_5429,N_4603,N_4607);
or U5430 (N_5430,N_4851,N_4814);
or U5431 (N_5431,N_4802,N_4489);
or U5432 (N_5432,N_4578,N_4932);
nand U5433 (N_5433,N_4700,N_4169);
nand U5434 (N_5434,N_4657,N_4989);
nor U5435 (N_5435,N_4212,N_4921);
nor U5436 (N_5436,N_4479,N_4922);
or U5437 (N_5437,N_4531,N_4210);
xor U5438 (N_5438,N_4058,N_4764);
nor U5439 (N_5439,N_4889,N_4004);
nor U5440 (N_5440,N_4808,N_4839);
and U5441 (N_5441,N_4256,N_4208);
nand U5442 (N_5442,N_4492,N_4340);
and U5443 (N_5443,N_4326,N_4269);
and U5444 (N_5444,N_4162,N_4198);
or U5445 (N_5445,N_4503,N_4017);
or U5446 (N_5446,N_4181,N_4535);
or U5447 (N_5447,N_4474,N_4562);
or U5448 (N_5448,N_4996,N_4583);
nand U5449 (N_5449,N_4892,N_4231);
and U5450 (N_5450,N_4561,N_4290);
nor U5451 (N_5451,N_4001,N_4929);
nor U5452 (N_5452,N_4590,N_4159);
nand U5453 (N_5453,N_4260,N_4341);
and U5454 (N_5454,N_4050,N_4280);
and U5455 (N_5455,N_4288,N_4950);
and U5456 (N_5456,N_4569,N_4099);
nand U5457 (N_5457,N_4598,N_4271);
or U5458 (N_5458,N_4009,N_4309);
nor U5459 (N_5459,N_4812,N_4467);
nor U5460 (N_5460,N_4951,N_4195);
or U5461 (N_5461,N_4287,N_4166);
xnor U5462 (N_5462,N_4346,N_4129);
or U5463 (N_5463,N_4095,N_4766);
and U5464 (N_5464,N_4691,N_4302);
nor U5465 (N_5465,N_4310,N_4312);
and U5466 (N_5466,N_4284,N_4769);
or U5467 (N_5467,N_4145,N_4925);
nor U5468 (N_5468,N_4860,N_4560);
and U5469 (N_5469,N_4119,N_4032);
nand U5470 (N_5470,N_4042,N_4094);
and U5471 (N_5471,N_4025,N_4402);
xnor U5472 (N_5472,N_4936,N_4594);
nor U5473 (N_5473,N_4759,N_4410);
nor U5474 (N_5474,N_4125,N_4414);
nand U5475 (N_5475,N_4112,N_4160);
nand U5476 (N_5476,N_4784,N_4475);
or U5477 (N_5477,N_4105,N_4871);
or U5478 (N_5478,N_4978,N_4514);
nand U5479 (N_5479,N_4398,N_4293);
and U5480 (N_5480,N_4505,N_4876);
xnor U5481 (N_5481,N_4696,N_4267);
or U5482 (N_5482,N_4750,N_4189);
and U5483 (N_5483,N_4823,N_4275);
nand U5484 (N_5484,N_4995,N_4073);
nand U5485 (N_5485,N_4566,N_4027);
nand U5486 (N_5486,N_4344,N_4077);
nand U5487 (N_5487,N_4971,N_4389);
nor U5488 (N_5488,N_4120,N_4517);
nor U5489 (N_5489,N_4595,N_4291);
xnor U5490 (N_5490,N_4423,N_4652);
nand U5491 (N_5491,N_4521,N_4552);
or U5492 (N_5492,N_4158,N_4285);
and U5493 (N_5493,N_4353,N_4642);
and U5494 (N_5494,N_4682,N_4444);
nor U5495 (N_5495,N_4928,N_4362);
nor U5496 (N_5496,N_4307,N_4930);
and U5497 (N_5497,N_4268,N_4550);
nor U5498 (N_5498,N_4320,N_4382);
nor U5499 (N_5499,N_4345,N_4116);
xnor U5500 (N_5500,N_4933,N_4338);
xnor U5501 (N_5501,N_4383,N_4253);
or U5502 (N_5502,N_4493,N_4437);
nand U5503 (N_5503,N_4755,N_4716);
and U5504 (N_5504,N_4784,N_4722);
nand U5505 (N_5505,N_4097,N_4861);
nand U5506 (N_5506,N_4342,N_4803);
nand U5507 (N_5507,N_4158,N_4045);
and U5508 (N_5508,N_4972,N_4092);
nand U5509 (N_5509,N_4650,N_4373);
nand U5510 (N_5510,N_4346,N_4737);
or U5511 (N_5511,N_4321,N_4233);
nor U5512 (N_5512,N_4179,N_4108);
and U5513 (N_5513,N_4996,N_4918);
xnor U5514 (N_5514,N_4934,N_4098);
nand U5515 (N_5515,N_4839,N_4635);
and U5516 (N_5516,N_4568,N_4583);
nand U5517 (N_5517,N_4095,N_4612);
or U5518 (N_5518,N_4727,N_4695);
nor U5519 (N_5519,N_4012,N_4810);
nand U5520 (N_5520,N_4085,N_4343);
and U5521 (N_5521,N_4153,N_4070);
nor U5522 (N_5522,N_4417,N_4142);
nor U5523 (N_5523,N_4501,N_4621);
nor U5524 (N_5524,N_4092,N_4171);
nor U5525 (N_5525,N_4801,N_4142);
xor U5526 (N_5526,N_4764,N_4215);
nor U5527 (N_5527,N_4088,N_4442);
nor U5528 (N_5528,N_4828,N_4581);
nor U5529 (N_5529,N_4615,N_4600);
xor U5530 (N_5530,N_4420,N_4456);
nor U5531 (N_5531,N_4477,N_4278);
nand U5532 (N_5532,N_4315,N_4936);
or U5533 (N_5533,N_4552,N_4205);
nand U5534 (N_5534,N_4480,N_4211);
nor U5535 (N_5535,N_4774,N_4422);
and U5536 (N_5536,N_4763,N_4211);
and U5537 (N_5537,N_4502,N_4299);
nand U5538 (N_5538,N_4231,N_4825);
or U5539 (N_5539,N_4981,N_4971);
xor U5540 (N_5540,N_4282,N_4915);
nand U5541 (N_5541,N_4782,N_4549);
nor U5542 (N_5542,N_4479,N_4916);
nor U5543 (N_5543,N_4355,N_4035);
nand U5544 (N_5544,N_4323,N_4254);
nor U5545 (N_5545,N_4370,N_4908);
nor U5546 (N_5546,N_4552,N_4615);
nor U5547 (N_5547,N_4677,N_4799);
and U5548 (N_5548,N_4754,N_4219);
xnor U5549 (N_5549,N_4912,N_4592);
xor U5550 (N_5550,N_4562,N_4437);
nand U5551 (N_5551,N_4363,N_4710);
nand U5552 (N_5552,N_4806,N_4787);
or U5553 (N_5553,N_4346,N_4009);
and U5554 (N_5554,N_4307,N_4195);
and U5555 (N_5555,N_4305,N_4819);
or U5556 (N_5556,N_4546,N_4472);
nor U5557 (N_5557,N_4650,N_4045);
nand U5558 (N_5558,N_4199,N_4156);
nor U5559 (N_5559,N_4005,N_4665);
nor U5560 (N_5560,N_4228,N_4791);
nand U5561 (N_5561,N_4740,N_4793);
nor U5562 (N_5562,N_4886,N_4415);
or U5563 (N_5563,N_4995,N_4435);
and U5564 (N_5564,N_4281,N_4850);
nand U5565 (N_5565,N_4960,N_4694);
nand U5566 (N_5566,N_4850,N_4258);
or U5567 (N_5567,N_4568,N_4253);
or U5568 (N_5568,N_4882,N_4377);
and U5569 (N_5569,N_4808,N_4448);
or U5570 (N_5570,N_4215,N_4321);
or U5571 (N_5571,N_4247,N_4075);
and U5572 (N_5572,N_4216,N_4133);
nor U5573 (N_5573,N_4654,N_4587);
nand U5574 (N_5574,N_4222,N_4774);
and U5575 (N_5575,N_4024,N_4390);
nor U5576 (N_5576,N_4564,N_4083);
and U5577 (N_5577,N_4665,N_4362);
nand U5578 (N_5578,N_4601,N_4425);
and U5579 (N_5579,N_4147,N_4825);
nor U5580 (N_5580,N_4094,N_4370);
nor U5581 (N_5581,N_4566,N_4154);
nand U5582 (N_5582,N_4601,N_4002);
and U5583 (N_5583,N_4417,N_4283);
nor U5584 (N_5584,N_4258,N_4636);
and U5585 (N_5585,N_4154,N_4702);
nand U5586 (N_5586,N_4726,N_4487);
or U5587 (N_5587,N_4785,N_4349);
xor U5588 (N_5588,N_4467,N_4410);
nor U5589 (N_5589,N_4364,N_4594);
nand U5590 (N_5590,N_4315,N_4773);
or U5591 (N_5591,N_4174,N_4878);
xnor U5592 (N_5592,N_4533,N_4587);
and U5593 (N_5593,N_4021,N_4641);
xnor U5594 (N_5594,N_4923,N_4351);
nor U5595 (N_5595,N_4496,N_4786);
nor U5596 (N_5596,N_4397,N_4449);
and U5597 (N_5597,N_4659,N_4420);
and U5598 (N_5598,N_4598,N_4034);
nor U5599 (N_5599,N_4213,N_4503);
and U5600 (N_5600,N_4844,N_4087);
nor U5601 (N_5601,N_4558,N_4131);
and U5602 (N_5602,N_4965,N_4074);
xnor U5603 (N_5603,N_4617,N_4454);
and U5604 (N_5604,N_4481,N_4215);
and U5605 (N_5605,N_4118,N_4668);
xor U5606 (N_5606,N_4335,N_4243);
or U5607 (N_5607,N_4686,N_4463);
and U5608 (N_5608,N_4135,N_4429);
nor U5609 (N_5609,N_4423,N_4898);
nor U5610 (N_5610,N_4733,N_4737);
nor U5611 (N_5611,N_4457,N_4115);
nor U5612 (N_5612,N_4730,N_4219);
nor U5613 (N_5613,N_4668,N_4788);
xor U5614 (N_5614,N_4384,N_4855);
nor U5615 (N_5615,N_4232,N_4191);
and U5616 (N_5616,N_4045,N_4907);
or U5617 (N_5617,N_4301,N_4428);
xnor U5618 (N_5618,N_4261,N_4121);
xor U5619 (N_5619,N_4737,N_4579);
nand U5620 (N_5620,N_4144,N_4996);
and U5621 (N_5621,N_4665,N_4372);
or U5622 (N_5622,N_4028,N_4385);
xnor U5623 (N_5623,N_4136,N_4685);
or U5624 (N_5624,N_4861,N_4489);
nand U5625 (N_5625,N_4450,N_4263);
xor U5626 (N_5626,N_4210,N_4224);
and U5627 (N_5627,N_4600,N_4717);
and U5628 (N_5628,N_4207,N_4543);
or U5629 (N_5629,N_4586,N_4056);
or U5630 (N_5630,N_4679,N_4267);
nor U5631 (N_5631,N_4383,N_4900);
nor U5632 (N_5632,N_4339,N_4075);
or U5633 (N_5633,N_4208,N_4999);
nor U5634 (N_5634,N_4211,N_4273);
or U5635 (N_5635,N_4828,N_4639);
nand U5636 (N_5636,N_4891,N_4472);
nor U5637 (N_5637,N_4346,N_4414);
nand U5638 (N_5638,N_4407,N_4886);
or U5639 (N_5639,N_4125,N_4837);
xnor U5640 (N_5640,N_4134,N_4755);
nand U5641 (N_5641,N_4533,N_4032);
nand U5642 (N_5642,N_4226,N_4519);
or U5643 (N_5643,N_4379,N_4741);
or U5644 (N_5644,N_4859,N_4509);
and U5645 (N_5645,N_4836,N_4857);
and U5646 (N_5646,N_4378,N_4581);
and U5647 (N_5647,N_4742,N_4927);
and U5648 (N_5648,N_4579,N_4674);
nand U5649 (N_5649,N_4597,N_4569);
nand U5650 (N_5650,N_4251,N_4179);
nor U5651 (N_5651,N_4935,N_4919);
and U5652 (N_5652,N_4194,N_4017);
and U5653 (N_5653,N_4742,N_4365);
nor U5654 (N_5654,N_4913,N_4257);
nand U5655 (N_5655,N_4136,N_4239);
xnor U5656 (N_5656,N_4331,N_4657);
nor U5657 (N_5657,N_4644,N_4425);
nand U5658 (N_5658,N_4154,N_4387);
or U5659 (N_5659,N_4086,N_4349);
nor U5660 (N_5660,N_4175,N_4766);
and U5661 (N_5661,N_4714,N_4267);
and U5662 (N_5662,N_4689,N_4024);
or U5663 (N_5663,N_4968,N_4003);
and U5664 (N_5664,N_4426,N_4856);
nand U5665 (N_5665,N_4287,N_4051);
nand U5666 (N_5666,N_4010,N_4899);
nor U5667 (N_5667,N_4964,N_4776);
or U5668 (N_5668,N_4963,N_4095);
and U5669 (N_5669,N_4380,N_4560);
nand U5670 (N_5670,N_4174,N_4468);
or U5671 (N_5671,N_4683,N_4166);
xnor U5672 (N_5672,N_4312,N_4648);
xor U5673 (N_5673,N_4755,N_4630);
nor U5674 (N_5674,N_4156,N_4092);
nor U5675 (N_5675,N_4400,N_4634);
nor U5676 (N_5676,N_4514,N_4170);
xnor U5677 (N_5677,N_4615,N_4058);
or U5678 (N_5678,N_4296,N_4660);
or U5679 (N_5679,N_4586,N_4330);
or U5680 (N_5680,N_4668,N_4545);
nand U5681 (N_5681,N_4138,N_4098);
xnor U5682 (N_5682,N_4828,N_4179);
nor U5683 (N_5683,N_4248,N_4269);
or U5684 (N_5684,N_4177,N_4673);
or U5685 (N_5685,N_4592,N_4882);
nand U5686 (N_5686,N_4570,N_4599);
nor U5687 (N_5687,N_4447,N_4368);
xor U5688 (N_5688,N_4201,N_4491);
and U5689 (N_5689,N_4758,N_4857);
or U5690 (N_5690,N_4692,N_4909);
xnor U5691 (N_5691,N_4691,N_4592);
nand U5692 (N_5692,N_4207,N_4216);
nor U5693 (N_5693,N_4853,N_4490);
nor U5694 (N_5694,N_4498,N_4416);
or U5695 (N_5695,N_4476,N_4255);
nor U5696 (N_5696,N_4041,N_4330);
nand U5697 (N_5697,N_4034,N_4198);
or U5698 (N_5698,N_4592,N_4553);
xnor U5699 (N_5699,N_4605,N_4165);
nor U5700 (N_5700,N_4738,N_4866);
nor U5701 (N_5701,N_4504,N_4915);
or U5702 (N_5702,N_4598,N_4611);
and U5703 (N_5703,N_4337,N_4749);
nand U5704 (N_5704,N_4016,N_4191);
and U5705 (N_5705,N_4083,N_4986);
and U5706 (N_5706,N_4549,N_4239);
or U5707 (N_5707,N_4462,N_4837);
or U5708 (N_5708,N_4830,N_4804);
or U5709 (N_5709,N_4782,N_4711);
xor U5710 (N_5710,N_4320,N_4483);
or U5711 (N_5711,N_4813,N_4606);
or U5712 (N_5712,N_4194,N_4300);
xnor U5713 (N_5713,N_4777,N_4909);
nand U5714 (N_5714,N_4452,N_4929);
and U5715 (N_5715,N_4661,N_4973);
and U5716 (N_5716,N_4444,N_4867);
or U5717 (N_5717,N_4068,N_4191);
xor U5718 (N_5718,N_4530,N_4497);
or U5719 (N_5719,N_4563,N_4833);
and U5720 (N_5720,N_4191,N_4085);
nand U5721 (N_5721,N_4582,N_4618);
and U5722 (N_5722,N_4130,N_4306);
nor U5723 (N_5723,N_4900,N_4377);
xor U5724 (N_5724,N_4388,N_4499);
or U5725 (N_5725,N_4908,N_4489);
nor U5726 (N_5726,N_4877,N_4435);
and U5727 (N_5727,N_4713,N_4921);
nand U5728 (N_5728,N_4988,N_4964);
or U5729 (N_5729,N_4099,N_4896);
and U5730 (N_5730,N_4641,N_4668);
nand U5731 (N_5731,N_4981,N_4384);
xor U5732 (N_5732,N_4274,N_4159);
xnor U5733 (N_5733,N_4110,N_4681);
or U5734 (N_5734,N_4621,N_4882);
and U5735 (N_5735,N_4716,N_4182);
xor U5736 (N_5736,N_4882,N_4108);
xnor U5737 (N_5737,N_4978,N_4153);
and U5738 (N_5738,N_4972,N_4968);
nor U5739 (N_5739,N_4338,N_4199);
nand U5740 (N_5740,N_4462,N_4365);
nand U5741 (N_5741,N_4662,N_4081);
nand U5742 (N_5742,N_4880,N_4064);
and U5743 (N_5743,N_4416,N_4924);
nand U5744 (N_5744,N_4690,N_4175);
nor U5745 (N_5745,N_4784,N_4170);
nand U5746 (N_5746,N_4375,N_4347);
and U5747 (N_5747,N_4146,N_4774);
nor U5748 (N_5748,N_4263,N_4260);
nand U5749 (N_5749,N_4976,N_4293);
nor U5750 (N_5750,N_4219,N_4502);
nand U5751 (N_5751,N_4287,N_4552);
or U5752 (N_5752,N_4877,N_4803);
or U5753 (N_5753,N_4786,N_4899);
and U5754 (N_5754,N_4206,N_4245);
nor U5755 (N_5755,N_4823,N_4195);
xor U5756 (N_5756,N_4217,N_4483);
nand U5757 (N_5757,N_4771,N_4583);
or U5758 (N_5758,N_4431,N_4561);
or U5759 (N_5759,N_4024,N_4971);
nor U5760 (N_5760,N_4916,N_4496);
and U5761 (N_5761,N_4673,N_4256);
nand U5762 (N_5762,N_4776,N_4768);
nor U5763 (N_5763,N_4831,N_4244);
nand U5764 (N_5764,N_4153,N_4398);
nand U5765 (N_5765,N_4653,N_4746);
xnor U5766 (N_5766,N_4447,N_4012);
or U5767 (N_5767,N_4460,N_4244);
nand U5768 (N_5768,N_4246,N_4377);
or U5769 (N_5769,N_4187,N_4536);
or U5770 (N_5770,N_4527,N_4150);
nand U5771 (N_5771,N_4542,N_4624);
nor U5772 (N_5772,N_4206,N_4049);
and U5773 (N_5773,N_4103,N_4090);
or U5774 (N_5774,N_4507,N_4132);
nor U5775 (N_5775,N_4412,N_4193);
and U5776 (N_5776,N_4795,N_4973);
nor U5777 (N_5777,N_4896,N_4737);
or U5778 (N_5778,N_4237,N_4665);
nor U5779 (N_5779,N_4155,N_4472);
nand U5780 (N_5780,N_4262,N_4369);
xnor U5781 (N_5781,N_4525,N_4801);
or U5782 (N_5782,N_4422,N_4184);
and U5783 (N_5783,N_4632,N_4982);
nand U5784 (N_5784,N_4550,N_4063);
xnor U5785 (N_5785,N_4728,N_4936);
or U5786 (N_5786,N_4597,N_4324);
nand U5787 (N_5787,N_4078,N_4393);
xnor U5788 (N_5788,N_4101,N_4477);
or U5789 (N_5789,N_4083,N_4196);
nor U5790 (N_5790,N_4345,N_4654);
nand U5791 (N_5791,N_4873,N_4552);
or U5792 (N_5792,N_4315,N_4031);
or U5793 (N_5793,N_4308,N_4541);
xnor U5794 (N_5794,N_4401,N_4760);
nor U5795 (N_5795,N_4748,N_4453);
nand U5796 (N_5796,N_4396,N_4534);
or U5797 (N_5797,N_4280,N_4370);
or U5798 (N_5798,N_4543,N_4762);
and U5799 (N_5799,N_4572,N_4908);
or U5800 (N_5800,N_4535,N_4577);
nor U5801 (N_5801,N_4824,N_4064);
nand U5802 (N_5802,N_4595,N_4304);
and U5803 (N_5803,N_4542,N_4240);
and U5804 (N_5804,N_4524,N_4221);
and U5805 (N_5805,N_4161,N_4863);
nand U5806 (N_5806,N_4912,N_4819);
xor U5807 (N_5807,N_4117,N_4532);
nand U5808 (N_5808,N_4465,N_4944);
or U5809 (N_5809,N_4730,N_4574);
nor U5810 (N_5810,N_4489,N_4027);
or U5811 (N_5811,N_4882,N_4261);
xor U5812 (N_5812,N_4279,N_4525);
nand U5813 (N_5813,N_4427,N_4386);
and U5814 (N_5814,N_4215,N_4571);
or U5815 (N_5815,N_4482,N_4807);
nor U5816 (N_5816,N_4809,N_4389);
nor U5817 (N_5817,N_4210,N_4564);
nand U5818 (N_5818,N_4696,N_4844);
nand U5819 (N_5819,N_4919,N_4676);
nor U5820 (N_5820,N_4103,N_4143);
or U5821 (N_5821,N_4997,N_4144);
or U5822 (N_5822,N_4601,N_4826);
or U5823 (N_5823,N_4308,N_4139);
or U5824 (N_5824,N_4861,N_4184);
or U5825 (N_5825,N_4297,N_4975);
or U5826 (N_5826,N_4246,N_4325);
and U5827 (N_5827,N_4404,N_4516);
and U5828 (N_5828,N_4689,N_4828);
and U5829 (N_5829,N_4227,N_4167);
and U5830 (N_5830,N_4049,N_4275);
nor U5831 (N_5831,N_4722,N_4882);
nor U5832 (N_5832,N_4476,N_4021);
and U5833 (N_5833,N_4187,N_4987);
and U5834 (N_5834,N_4312,N_4652);
nor U5835 (N_5835,N_4902,N_4133);
nor U5836 (N_5836,N_4463,N_4688);
and U5837 (N_5837,N_4384,N_4951);
nand U5838 (N_5838,N_4684,N_4964);
nor U5839 (N_5839,N_4461,N_4254);
or U5840 (N_5840,N_4267,N_4155);
nand U5841 (N_5841,N_4186,N_4491);
or U5842 (N_5842,N_4700,N_4282);
or U5843 (N_5843,N_4803,N_4585);
and U5844 (N_5844,N_4086,N_4815);
xnor U5845 (N_5845,N_4116,N_4386);
or U5846 (N_5846,N_4738,N_4092);
and U5847 (N_5847,N_4536,N_4244);
and U5848 (N_5848,N_4770,N_4464);
nor U5849 (N_5849,N_4441,N_4118);
or U5850 (N_5850,N_4792,N_4135);
and U5851 (N_5851,N_4817,N_4066);
xor U5852 (N_5852,N_4744,N_4319);
nand U5853 (N_5853,N_4544,N_4372);
xor U5854 (N_5854,N_4553,N_4545);
and U5855 (N_5855,N_4056,N_4306);
nand U5856 (N_5856,N_4830,N_4582);
or U5857 (N_5857,N_4763,N_4010);
nand U5858 (N_5858,N_4316,N_4387);
nand U5859 (N_5859,N_4728,N_4510);
and U5860 (N_5860,N_4695,N_4210);
nor U5861 (N_5861,N_4262,N_4230);
and U5862 (N_5862,N_4860,N_4879);
and U5863 (N_5863,N_4643,N_4150);
nand U5864 (N_5864,N_4986,N_4724);
nand U5865 (N_5865,N_4556,N_4576);
nand U5866 (N_5866,N_4283,N_4521);
nand U5867 (N_5867,N_4604,N_4062);
nor U5868 (N_5868,N_4387,N_4869);
xnor U5869 (N_5869,N_4247,N_4987);
xor U5870 (N_5870,N_4938,N_4563);
and U5871 (N_5871,N_4013,N_4349);
and U5872 (N_5872,N_4733,N_4848);
nor U5873 (N_5873,N_4829,N_4685);
nand U5874 (N_5874,N_4980,N_4371);
and U5875 (N_5875,N_4610,N_4008);
nand U5876 (N_5876,N_4898,N_4185);
nand U5877 (N_5877,N_4195,N_4551);
or U5878 (N_5878,N_4190,N_4285);
or U5879 (N_5879,N_4250,N_4588);
and U5880 (N_5880,N_4027,N_4945);
or U5881 (N_5881,N_4759,N_4014);
nor U5882 (N_5882,N_4387,N_4192);
xnor U5883 (N_5883,N_4598,N_4325);
and U5884 (N_5884,N_4918,N_4260);
or U5885 (N_5885,N_4347,N_4255);
and U5886 (N_5886,N_4609,N_4046);
and U5887 (N_5887,N_4957,N_4637);
or U5888 (N_5888,N_4415,N_4406);
and U5889 (N_5889,N_4942,N_4819);
and U5890 (N_5890,N_4859,N_4246);
or U5891 (N_5891,N_4273,N_4298);
or U5892 (N_5892,N_4910,N_4017);
xnor U5893 (N_5893,N_4171,N_4389);
nand U5894 (N_5894,N_4795,N_4404);
or U5895 (N_5895,N_4796,N_4150);
xor U5896 (N_5896,N_4664,N_4456);
and U5897 (N_5897,N_4202,N_4819);
and U5898 (N_5898,N_4539,N_4109);
xor U5899 (N_5899,N_4305,N_4525);
nand U5900 (N_5900,N_4399,N_4214);
nand U5901 (N_5901,N_4858,N_4710);
nand U5902 (N_5902,N_4700,N_4401);
nand U5903 (N_5903,N_4991,N_4545);
and U5904 (N_5904,N_4870,N_4101);
and U5905 (N_5905,N_4719,N_4959);
nor U5906 (N_5906,N_4843,N_4722);
or U5907 (N_5907,N_4065,N_4006);
or U5908 (N_5908,N_4331,N_4589);
nor U5909 (N_5909,N_4207,N_4080);
nand U5910 (N_5910,N_4378,N_4430);
nand U5911 (N_5911,N_4992,N_4235);
and U5912 (N_5912,N_4470,N_4404);
or U5913 (N_5913,N_4745,N_4751);
and U5914 (N_5914,N_4527,N_4687);
nand U5915 (N_5915,N_4858,N_4243);
xor U5916 (N_5916,N_4305,N_4965);
and U5917 (N_5917,N_4420,N_4280);
or U5918 (N_5918,N_4814,N_4917);
nand U5919 (N_5919,N_4992,N_4319);
and U5920 (N_5920,N_4743,N_4697);
and U5921 (N_5921,N_4649,N_4063);
nand U5922 (N_5922,N_4614,N_4142);
nor U5923 (N_5923,N_4043,N_4848);
nor U5924 (N_5924,N_4608,N_4555);
and U5925 (N_5925,N_4043,N_4176);
or U5926 (N_5926,N_4720,N_4867);
or U5927 (N_5927,N_4667,N_4421);
nor U5928 (N_5928,N_4514,N_4235);
xnor U5929 (N_5929,N_4423,N_4114);
or U5930 (N_5930,N_4806,N_4437);
or U5931 (N_5931,N_4614,N_4873);
xnor U5932 (N_5932,N_4467,N_4557);
nand U5933 (N_5933,N_4199,N_4398);
or U5934 (N_5934,N_4563,N_4945);
and U5935 (N_5935,N_4358,N_4206);
and U5936 (N_5936,N_4802,N_4892);
xnor U5937 (N_5937,N_4820,N_4631);
nor U5938 (N_5938,N_4586,N_4874);
and U5939 (N_5939,N_4578,N_4539);
or U5940 (N_5940,N_4784,N_4497);
or U5941 (N_5941,N_4137,N_4541);
nand U5942 (N_5942,N_4703,N_4315);
nor U5943 (N_5943,N_4764,N_4042);
nor U5944 (N_5944,N_4600,N_4773);
nor U5945 (N_5945,N_4049,N_4358);
nand U5946 (N_5946,N_4227,N_4502);
or U5947 (N_5947,N_4783,N_4941);
nor U5948 (N_5948,N_4317,N_4627);
nand U5949 (N_5949,N_4764,N_4795);
nor U5950 (N_5950,N_4855,N_4654);
xnor U5951 (N_5951,N_4110,N_4717);
and U5952 (N_5952,N_4037,N_4891);
nand U5953 (N_5953,N_4771,N_4169);
or U5954 (N_5954,N_4940,N_4100);
nor U5955 (N_5955,N_4342,N_4053);
nor U5956 (N_5956,N_4185,N_4153);
or U5957 (N_5957,N_4686,N_4848);
and U5958 (N_5958,N_4773,N_4624);
and U5959 (N_5959,N_4270,N_4376);
nand U5960 (N_5960,N_4976,N_4511);
xnor U5961 (N_5961,N_4676,N_4856);
nor U5962 (N_5962,N_4188,N_4017);
and U5963 (N_5963,N_4749,N_4092);
and U5964 (N_5964,N_4443,N_4213);
or U5965 (N_5965,N_4437,N_4038);
and U5966 (N_5966,N_4168,N_4717);
and U5967 (N_5967,N_4512,N_4530);
nand U5968 (N_5968,N_4872,N_4634);
and U5969 (N_5969,N_4354,N_4898);
xnor U5970 (N_5970,N_4278,N_4392);
and U5971 (N_5971,N_4256,N_4402);
nor U5972 (N_5972,N_4708,N_4887);
xnor U5973 (N_5973,N_4329,N_4413);
nand U5974 (N_5974,N_4712,N_4420);
or U5975 (N_5975,N_4836,N_4271);
nor U5976 (N_5976,N_4426,N_4547);
nor U5977 (N_5977,N_4055,N_4812);
nand U5978 (N_5978,N_4281,N_4173);
nor U5979 (N_5979,N_4917,N_4678);
nand U5980 (N_5980,N_4309,N_4545);
or U5981 (N_5981,N_4479,N_4978);
nor U5982 (N_5982,N_4628,N_4627);
and U5983 (N_5983,N_4575,N_4963);
nor U5984 (N_5984,N_4687,N_4264);
or U5985 (N_5985,N_4801,N_4554);
nor U5986 (N_5986,N_4712,N_4153);
or U5987 (N_5987,N_4300,N_4485);
nand U5988 (N_5988,N_4594,N_4671);
nand U5989 (N_5989,N_4132,N_4342);
or U5990 (N_5990,N_4441,N_4110);
nand U5991 (N_5991,N_4805,N_4625);
and U5992 (N_5992,N_4267,N_4028);
nor U5993 (N_5993,N_4241,N_4155);
nor U5994 (N_5994,N_4680,N_4454);
nor U5995 (N_5995,N_4623,N_4385);
nand U5996 (N_5996,N_4318,N_4978);
nand U5997 (N_5997,N_4323,N_4851);
or U5998 (N_5998,N_4275,N_4699);
nand U5999 (N_5999,N_4214,N_4748);
nand U6000 (N_6000,N_5154,N_5872);
xnor U6001 (N_6001,N_5662,N_5783);
nand U6002 (N_6002,N_5284,N_5216);
nand U6003 (N_6003,N_5102,N_5003);
or U6004 (N_6004,N_5565,N_5130);
xnor U6005 (N_6005,N_5789,N_5695);
xnor U6006 (N_6006,N_5489,N_5016);
or U6007 (N_6007,N_5204,N_5366);
nor U6008 (N_6008,N_5183,N_5397);
or U6009 (N_6009,N_5038,N_5959);
and U6010 (N_6010,N_5206,N_5004);
or U6011 (N_6011,N_5466,N_5920);
xor U6012 (N_6012,N_5054,N_5069);
nor U6013 (N_6013,N_5833,N_5879);
nor U6014 (N_6014,N_5231,N_5376);
nand U6015 (N_6015,N_5954,N_5190);
or U6016 (N_6016,N_5581,N_5125);
nor U6017 (N_6017,N_5659,N_5498);
or U6018 (N_6018,N_5573,N_5707);
xnor U6019 (N_6019,N_5388,N_5664);
nor U6020 (N_6020,N_5624,N_5324);
xor U6021 (N_6021,N_5785,N_5224);
xnor U6022 (N_6022,N_5264,N_5274);
and U6023 (N_6023,N_5962,N_5219);
nor U6024 (N_6024,N_5876,N_5652);
nor U6025 (N_6025,N_5122,N_5586);
or U6026 (N_6026,N_5481,N_5764);
nand U6027 (N_6027,N_5591,N_5223);
and U6028 (N_6028,N_5618,N_5487);
nor U6029 (N_6029,N_5492,N_5916);
nand U6030 (N_6030,N_5716,N_5305);
or U6031 (N_6031,N_5890,N_5436);
nand U6032 (N_6032,N_5454,N_5060);
or U6033 (N_6033,N_5243,N_5734);
and U6034 (N_6034,N_5234,N_5170);
and U6035 (N_6035,N_5812,N_5157);
or U6036 (N_6036,N_5275,N_5021);
nand U6037 (N_6037,N_5596,N_5367);
and U6038 (N_6038,N_5158,N_5490);
xor U6039 (N_6039,N_5052,N_5497);
or U6040 (N_6040,N_5688,N_5176);
nand U6041 (N_6041,N_5855,N_5257);
nand U6042 (N_6042,N_5718,N_5251);
nor U6043 (N_6043,N_5296,N_5336);
nand U6044 (N_6044,N_5164,N_5646);
nor U6045 (N_6045,N_5484,N_5922);
nand U6046 (N_6046,N_5899,N_5988);
nor U6047 (N_6047,N_5273,N_5051);
or U6048 (N_6048,N_5373,N_5555);
nor U6049 (N_6049,N_5720,N_5094);
or U6050 (N_6050,N_5647,N_5001);
or U6051 (N_6051,N_5831,N_5897);
and U6052 (N_6052,N_5518,N_5491);
nand U6053 (N_6053,N_5469,N_5149);
nand U6054 (N_6054,N_5196,N_5532);
or U6055 (N_6055,N_5145,N_5961);
and U6056 (N_6056,N_5625,N_5299);
or U6057 (N_6057,N_5358,N_5008);
or U6058 (N_6058,N_5749,N_5545);
and U6059 (N_6059,N_5293,N_5445);
and U6060 (N_6060,N_5369,N_5352);
and U6061 (N_6061,N_5632,N_5623);
nor U6062 (N_6062,N_5665,N_5280);
and U6063 (N_6063,N_5761,N_5056);
and U6064 (N_6064,N_5282,N_5870);
nand U6065 (N_6065,N_5576,N_5285);
nand U6066 (N_6066,N_5807,N_5998);
and U6067 (N_6067,N_5730,N_5560);
xnor U6068 (N_6068,N_5171,N_5858);
nand U6069 (N_6069,N_5245,N_5111);
nor U6070 (N_6070,N_5940,N_5236);
nor U6071 (N_6071,N_5078,N_5594);
and U6072 (N_6072,N_5743,N_5391);
and U6073 (N_6073,N_5146,N_5648);
or U6074 (N_6074,N_5522,N_5809);
nor U6075 (N_6075,N_5086,N_5902);
or U6076 (N_6076,N_5419,N_5825);
and U6077 (N_6077,N_5744,N_5690);
or U6078 (N_6078,N_5992,N_5929);
or U6079 (N_6079,N_5974,N_5815);
nor U6080 (N_6080,N_5393,N_5141);
or U6081 (N_6081,N_5026,N_5898);
nor U6082 (N_6082,N_5649,N_5830);
xnor U6083 (N_6083,N_5200,N_5944);
and U6084 (N_6084,N_5042,N_5950);
or U6085 (N_6085,N_5503,N_5975);
or U6086 (N_6086,N_5455,N_5029);
nor U6087 (N_6087,N_5258,N_5344);
nand U6088 (N_6088,N_5033,N_5242);
nor U6089 (N_6089,N_5933,N_5129);
nor U6090 (N_6090,N_5509,N_5381);
and U6091 (N_6091,N_5605,N_5856);
or U6092 (N_6092,N_5639,N_5750);
or U6093 (N_6093,N_5349,N_5763);
nor U6094 (N_6094,N_5109,N_5568);
and U6095 (N_6095,N_5453,N_5713);
nor U6096 (N_6096,N_5112,N_5414);
or U6097 (N_6097,N_5116,N_5207);
xor U6098 (N_6098,N_5980,N_5816);
or U6099 (N_6099,N_5229,N_5579);
and U6100 (N_6100,N_5602,N_5409);
nand U6101 (N_6101,N_5525,N_5607);
or U6102 (N_6102,N_5092,N_5240);
xnor U6103 (N_6103,N_5262,N_5569);
nand U6104 (N_6104,N_5776,N_5850);
or U6105 (N_6105,N_5524,N_5353);
or U6106 (N_6106,N_5127,N_5045);
nor U6107 (N_6107,N_5502,N_5194);
xnor U6108 (N_6108,N_5197,N_5089);
nand U6109 (N_6109,N_5418,N_5844);
nor U6110 (N_6110,N_5059,N_5631);
nand U6111 (N_6111,N_5198,N_5926);
nand U6112 (N_6112,N_5660,N_5612);
nand U6113 (N_6113,N_5722,N_5517);
nor U6114 (N_6114,N_5805,N_5860);
and U6115 (N_6115,N_5173,N_5803);
or U6116 (N_6116,N_5259,N_5931);
and U6117 (N_6117,N_5727,N_5055);
or U6118 (N_6118,N_5709,N_5433);
nor U6119 (N_6119,N_5082,N_5239);
and U6120 (N_6120,N_5629,N_5679);
nor U6121 (N_6121,N_5510,N_5210);
or U6122 (N_6122,N_5601,N_5226);
or U6123 (N_6123,N_5057,N_5272);
nand U6124 (N_6124,N_5883,N_5717);
and U6125 (N_6125,N_5759,N_5006);
nand U6126 (N_6126,N_5392,N_5277);
or U6127 (N_6127,N_5339,N_5348);
nand U6128 (N_6128,N_5838,N_5984);
and U6129 (N_6129,N_5420,N_5681);
nor U6130 (N_6130,N_5018,N_5731);
and U6131 (N_6131,N_5979,N_5768);
or U6132 (N_6132,N_5495,N_5777);
and U6133 (N_6133,N_5312,N_5758);
nor U6134 (N_6134,N_5614,N_5286);
or U6135 (N_6135,N_5009,N_5824);
and U6136 (N_6136,N_5175,N_5686);
nand U6137 (N_6137,N_5435,N_5477);
or U6138 (N_6138,N_5804,N_5185);
xnor U6139 (N_6139,N_5249,N_5449);
nor U6140 (N_6140,N_5041,N_5637);
or U6141 (N_6141,N_5209,N_5039);
nor U6142 (N_6142,N_5620,N_5889);
or U6143 (N_6143,N_5482,N_5235);
or U6144 (N_6144,N_5827,N_5553);
and U6145 (N_6145,N_5737,N_5972);
nor U6146 (N_6146,N_5582,N_5745);
or U6147 (N_6147,N_5499,N_5557);
nor U6148 (N_6148,N_5085,N_5372);
nand U6149 (N_6149,N_5031,N_5203);
nor U6150 (N_6150,N_5252,N_5480);
and U6151 (N_6151,N_5301,N_5548);
xor U6152 (N_6152,N_5746,N_5182);
and U6153 (N_6153,N_5460,N_5297);
or U6154 (N_6154,N_5027,N_5053);
or U6155 (N_6155,N_5314,N_5318);
and U6156 (N_6156,N_5007,N_5539);
nor U6157 (N_6157,N_5327,N_5893);
or U6158 (N_6158,N_5762,N_5871);
and U6159 (N_6159,N_5609,N_5911);
xnor U6160 (N_6160,N_5329,N_5636);
nor U6161 (N_6161,N_5124,N_5521);
nand U6162 (N_6162,N_5541,N_5395);
nor U6163 (N_6163,N_5426,N_5775);
nor U6164 (N_6164,N_5658,N_5120);
nor U6165 (N_6165,N_5494,N_5861);
nand U6166 (N_6166,N_5799,N_5507);
nor U6167 (N_6167,N_5696,N_5315);
nor U6168 (N_6168,N_5993,N_5685);
xor U6169 (N_6169,N_5306,N_5705);
nand U6170 (N_6170,N_5653,N_5673);
nor U6171 (N_6171,N_5332,N_5968);
or U6172 (N_6172,N_5802,N_5338);
and U6173 (N_6173,N_5757,N_5266);
nand U6174 (N_6174,N_5523,N_5990);
nor U6175 (N_6175,N_5921,N_5583);
xor U6176 (N_6176,N_5852,N_5733);
and U6177 (N_6177,N_5951,N_5821);
or U6178 (N_6178,N_5295,N_5794);
nand U6179 (N_6179,N_5706,N_5997);
or U6180 (N_6180,N_5364,N_5989);
and U6181 (N_6181,N_5829,N_5140);
nand U6182 (N_6182,N_5135,N_5389);
nand U6183 (N_6183,N_5702,N_5865);
or U6184 (N_6184,N_5192,N_5177);
nand U6185 (N_6185,N_5062,N_5778);
nand U6186 (N_6186,N_5148,N_5347);
or U6187 (N_6187,N_5361,N_5368);
or U6188 (N_6188,N_5782,N_5735);
nand U6189 (N_6189,N_5691,N_5398);
nand U6190 (N_6190,N_5611,N_5843);
nand U6191 (N_6191,N_5093,N_5096);
nor U6192 (N_6192,N_5310,N_5715);
nand U6193 (N_6193,N_5379,N_5956);
xnor U6194 (N_6194,N_5810,N_5996);
or U6195 (N_6195,N_5533,N_5211);
and U6196 (N_6196,N_5544,N_5982);
nand U6197 (N_6197,N_5084,N_5873);
nand U6198 (N_6198,N_5694,N_5857);
nor U6199 (N_6199,N_5698,N_5047);
nand U6200 (N_6200,N_5374,N_5070);
or U6201 (N_6201,N_5322,N_5946);
nor U6202 (N_6202,N_5342,N_5121);
or U6203 (N_6203,N_5708,N_5986);
nor U6204 (N_6204,N_5114,N_5650);
xor U6205 (N_6205,N_5848,N_5808);
nand U6206 (N_6206,N_5193,N_5437);
nand U6207 (N_6207,N_5676,N_5215);
nor U6208 (N_6208,N_5942,N_5447);
or U6209 (N_6209,N_5640,N_5836);
nand U6210 (N_6210,N_5065,N_5105);
xor U6211 (N_6211,N_5377,N_5519);
nand U6212 (N_6212,N_5323,N_5534);
nor U6213 (N_6213,N_5080,N_5895);
nand U6214 (N_6214,N_5955,N_5790);
nand U6215 (N_6215,N_5365,N_5474);
nand U6216 (N_6216,N_5244,N_5813);
nand U6217 (N_6217,N_5464,N_5630);
nand U6218 (N_6218,N_5471,N_5947);
and U6219 (N_6219,N_5739,N_5877);
nand U6220 (N_6220,N_5504,N_5119);
nor U6221 (N_6221,N_5167,N_5030);
or U6222 (N_6222,N_5963,N_5050);
nor U6223 (N_6223,N_5232,N_5723);
and U6224 (N_6224,N_5567,N_5958);
nor U6225 (N_6225,N_5115,N_5303);
nand U6226 (N_6226,N_5136,N_5287);
and U6227 (N_6227,N_5422,N_5246);
nor U6228 (N_6228,N_5725,N_5627);
or U6229 (N_6229,N_5866,N_5796);
xnor U6230 (N_6230,N_5408,N_5985);
nand U6231 (N_6231,N_5994,N_5320);
or U6232 (N_6232,N_5655,N_5868);
nor U6233 (N_6233,N_5819,N_5128);
nand U6234 (N_6234,N_5036,N_5307);
and U6235 (N_6235,N_5936,N_5514);
and U6236 (N_6236,N_5046,N_5401);
or U6237 (N_6237,N_5896,N_5237);
or U6238 (N_6238,N_5867,N_5847);
and U6239 (N_6239,N_5987,N_5081);
or U6240 (N_6240,N_5106,N_5025);
and U6241 (N_6241,N_5180,N_5642);
or U6242 (N_6242,N_5270,N_5820);
nand U6243 (N_6243,N_5666,N_5091);
nor U6244 (N_6244,N_5766,N_5832);
or U6245 (N_6245,N_5400,N_5184);
or U6246 (N_6246,N_5276,N_5924);
and U6247 (N_6247,N_5538,N_5587);
xor U6248 (N_6248,N_5948,N_5438);
or U6249 (N_6249,N_5585,N_5360);
and U6250 (N_6250,N_5588,N_5371);
nor U6251 (N_6251,N_5462,N_5095);
and U6252 (N_6252,N_5859,N_5387);
or U6253 (N_6253,N_5359,N_5887);
or U6254 (N_6254,N_5779,N_5268);
and U6255 (N_6255,N_5619,N_5754);
nand U6256 (N_6256,N_5279,N_5467);
nand U6257 (N_6257,N_5869,N_5147);
nor U6258 (N_6258,N_5385,N_5542);
and U6259 (N_6259,N_5227,N_5826);
nor U6260 (N_6260,N_5978,N_5651);
or U6261 (N_6261,N_5319,N_5927);
nor U6262 (N_6262,N_5903,N_5769);
nand U6263 (N_6263,N_5577,N_5317);
nand U6264 (N_6264,N_5104,N_5732);
nand U6265 (N_6265,N_5891,N_5719);
nand U6266 (N_6266,N_5930,N_5174);
or U6267 (N_6267,N_5298,N_5513);
nand U6268 (N_6268,N_5615,N_5788);
nand U6269 (N_6269,N_5846,N_5780);
nand U6270 (N_6270,N_5325,N_5465);
nor U6271 (N_6271,N_5034,N_5668);
or U6272 (N_6272,N_5547,N_5151);
or U6273 (N_6273,N_5726,N_5399);
nand U6274 (N_6274,N_5281,N_5269);
and U6275 (N_6275,N_5603,N_5983);
or U6276 (N_6276,N_5440,N_5335);
xor U6277 (N_6277,N_5217,N_5017);
xnor U6278 (N_6278,N_5915,N_5058);
nor U6279 (N_6279,N_5434,N_5443);
nor U6280 (N_6280,N_5431,N_5580);
xor U6281 (N_6281,N_5977,N_5291);
nor U6282 (N_6282,N_5981,N_5256);
nand U6283 (N_6283,N_5238,N_5678);
xnor U6284 (N_6284,N_5496,N_5839);
xor U6285 (N_6285,N_5500,N_5202);
and U6286 (N_6286,N_5067,N_5172);
and U6287 (N_6287,N_5066,N_5014);
xor U6288 (N_6288,N_5132,N_5461);
and U6289 (N_6289,N_5967,N_5863);
nor U6290 (N_6290,N_5571,N_5995);
and U6291 (N_6291,N_5905,N_5561);
nand U6292 (N_6292,N_5772,N_5015);
nor U6293 (N_6293,N_5073,N_5787);
nor U6294 (N_6294,N_5765,N_5040);
nand U6295 (N_6295,N_5597,N_5241);
or U6296 (N_6296,N_5090,N_5308);
nand U6297 (N_6297,N_5456,N_5378);
and U6298 (N_6298,N_5535,N_5024);
and U6299 (N_6299,N_5446,N_5670);
or U6300 (N_6300,N_5355,N_5792);
nand U6301 (N_6301,N_5061,N_5901);
nor U6302 (N_6302,N_5386,N_5134);
and U6303 (N_6303,N_5851,N_5753);
and U6304 (N_6304,N_5250,N_5405);
nor U6305 (N_6305,N_5689,N_5537);
nor U6306 (N_6306,N_5801,N_5774);
and U6307 (N_6307,N_5283,N_5222);
or U6308 (N_6308,N_5156,N_5598);
nor U6309 (N_6309,N_5012,N_5728);
and U6310 (N_6310,N_5600,N_5949);
nor U6311 (N_6311,N_5321,N_5101);
or U6312 (N_6312,N_5442,N_5404);
nor U6313 (N_6313,N_5515,N_5593);
nor U6314 (N_6314,N_5110,N_5674);
xor U6315 (N_6315,N_5700,N_5526);
or U6316 (N_6316,N_5751,N_5729);
nand U6317 (N_6317,N_5468,N_5072);
or U6318 (N_6318,N_5412,N_5806);
or U6319 (N_6319,N_5189,N_5699);
nand U6320 (N_6320,N_5205,N_5362);
or U6321 (N_6321,N_5928,N_5075);
xnor U6322 (N_6322,N_5218,N_5278);
and U6323 (N_6323,N_5097,N_5022);
nor U6324 (N_6324,N_5786,N_5107);
and U6325 (N_6325,N_5589,N_5396);
nor U6326 (N_6326,N_5656,N_5667);
nor U6327 (N_6327,N_5828,N_5552);
nand U6328 (N_6328,N_5212,N_5350);
or U6329 (N_6329,N_5126,N_5516);
nand U6330 (N_6330,N_5773,N_5575);
and U6331 (N_6331,N_5874,N_5152);
and U6332 (N_6332,N_5578,N_5584);
nand U6333 (N_6333,N_5939,N_5721);
nand U6334 (N_6334,N_5188,N_5740);
or U6335 (N_6335,N_5351,N_5260);
nand U6336 (N_6336,N_5439,N_5049);
nor U6337 (N_6337,N_5800,N_5595);
or U6338 (N_6338,N_5613,N_5248);
nand U6339 (N_6339,N_5363,N_5520);
nand U6340 (N_6340,N_5160,N_5937);
and U6341 (N_6341,N_5934,N_5019);
nand U6342 (N_6342,N_5448,N_5459);
or U6343 (N_6343,N_5900,N_5292);
nor U6344 (N_6344,N_5311,N_5752);
nor U6345 (N_6345,N_5341,N_5912);
and U6346 (N_6346,N_5976,N_5225);
and U6347 (N_6347,N_5020,N_5626);
nor U6348 (N_6348,N_5087,N_5823);
nor U6349 (N_6349,N_5452,N_5079);
and U6350 (N_6350,N_5470,N_5076);
and U6351 (N_6351,N_5634,N_5501);
and U6352 (N_6352,N_5406,N_5736);
nand U6353 (N_6353,N_5923,N_5488);
and U6354 (N_6354,N_5458,N_5330);
nand U6355 (N_6355,N_5131,N_5165);
and U6356 (N_6356,N_5044,N_5845);
nand U6357 (N_6357,N_5913,N_5904);
xnor U6358 (N_6358,N_5621,N_5849);
xor U6359 (N_6359,N_5558,N_5403);
xnor U6360 (N_6360,N_5712,N_5328);
nand U6361 (N_6361,N_5635,N_5068);
xnor U6362 (N_6362,N_5383,N_5064);
nand U6363 (N_6363,N_5380,N_5617);
and U6364 (N_6364,N_5610,N_5384);
nand U6365 (N_6365,N_5233,N_5531);
nor U6366 (N_6366,N_5755,N_5063);
or U6367 (N_6367,N_5424,N_5407);
nand U6368 (N_6368,N_5088,N_5028);
nand U6369 (N_6369,N_5168,N_5410);
nor U6370 (N_6370,N_5290,N_5162);
nor U6371 (N_6371,N_5313,N_5247);
or U6372 (N_6372,N_5797,N_5117);
and U6373 (N_6373,N_5337,N_5756);
or U6374 (N_6374,N_5304,N_5529);
nor U6375 (N_6375,N_5214,N_5427);
nand U6376 (N_6376,N_5892,N_5113);
nand U6377 (N_6377,N_5043,N_5854);
and U6378 (N_6378,N_5770,N_5817);
or U6379 (N_6379,N_5142,N_5345);
and U6380 (N_6380,N_5166,N_5375);
nor U6381 (N_6381,N_5346,N_5098);
and U6382 (N_6382,N_5894,N_5687);
nand U6383 (N_6383,N_5703,N_5738);
xnor U6384 (N_6384,N_5853,N_5528);
nor U6385 (N_6385,N_5118,N_5748);
nor U6386 (N_6386,N_5506,N_5952);
nor U6387 (N_6387,N_5032,N_5508);
and U6388 (N_6388,N_5953,N_5382);
nand U6389 (N_6389,N_5463,N_5261);
or U6390 (N_6390,N_5444,N_5253);
nor U6391 (N_6391,N_5159,N_5144);
and U6392 (N_6392,N_5178,N_5133);
nor U6393 (N_6393,N_5562,N_5143);
or U6394 (N_6394,N_5862,N_5415);
xor U6395 (N_6395,N_5566,N_5294);
or U6396 (N_6396,N_5724,N_5878);
or U6397 (N_6397,N_5483,N_5841);
nand U6398 (N_6398,N_5633,N_5965);
or U6399 (N_6399,N_5622,N_5475);
or U6400 (N_6400,N_5645,N_5155);
nor U6401 (N_6401,N_5010,N_5302);
or U6402 (N_6402,N_5512,N_5935);
nand U6403 (N_6403,N_5333,N_5331);
and U6404 (N_6404,N_5563,N_5885);
xnor U6405 (N_6405,N_5334,N_5875);
and U6406 (N_6406,N_5457,N_5536);
nand U6407 (N_6407,N_5864,N_5478);
or U6408 (N_6408,N_5000,N_5590);
nor U6409 (N_6409,N_5908,N_5811);
nor U6410 (N_6410,N_5417,N_5035);
nand U6411 (N_6411,N_5964,N_5966);
and U6412 (N_6412,N_5394,N_5886);
or U6413 (N_6413,N_5781,N_5880);
or U6414 (N_6414,N_5187,N_5914);
nor U6415 (N_6415,N_5451,N_5628);
or U6416 (N_6416,N_5201,N_5657);
nor U6417 (N_6417,N_5071,N_5932);
and U6418 (N_6418,N_5429,N_5814);
nor U6419 (N_6419,N_5263,N_5559);
nor U6420 (N_6420,N_5680,N_5220);
nor U6421 (N_6421,N_5641,N_5199);
or U6422 (N_6422,N_5300,N_5711);
nor U6423 (N_6423,N_5551,N_5005);
nor U6424 (N_6424,N_5479,N_5357);
or U6425 (N_6425,N_5818,N_5710);
nand U6426 (N_6426,N_5161,N_5549);
or U6427 (N_6427,N_5099,N_5530);
nand U6428 (N_6428,N_5999,N_5704);
or U6429 (N_6429,N_5693,N_5473);
nor U6430 (N_6430,N_5390,N_5682);
nor U6431 (N_6431,N_5230,N_5960);
and U6432 (N_6432,N_5697,N_5784);
nor U6433 (N_6433,N_5074,N_5543);
nor U6434 (N_6434,N_5572,N_5969);
nor U6435 (N_6435,N_5011,N_5925);
or U6436 (N_6436,N_5606,N_5023);
or U6437 (N_6437,N_5604,N_5592);
nand U6438 (N_6438,N_5123,N_5326);
and U6439 (N_6439,N_5970,N_5430);
or U6440 (N_6440,N_5195,N_5910);
nand U6441 (N_6441,N_5265,N_5644);
nor U6442 (N_6442,N_5413,N_5485);
or U6443 (N_6443,N_5556,N_5669);
nand U6444 (N_6444,N_5881,N_5540);
xnor U6445 (N_6445,N_5416,N_5441);
or U6446 (N_6446,N_5137,N_5791);
and U6447 (N_6447,N_5684,N_5472);
and U6448 (N_6448,N_5882,N_5991);
or U6449 (N_6449,N_5511,N_5767);
or U6450 (N_6450,N_5554,N_5048);
nor U6451 (N_6451,N_5271,N_5747);
xnor U6452 (N_6452,N_5428,N_5677);
nand U6453 (N_6453,N_5425,N_5077);
xor U6454 (N_6454,N_5888,N_5169);
nand U6455 (N_6455,N_5255,N_5840);
and U6456 (N_6456,N_5599,N_5343);
nor U6457 (N_6457,N_5316,N_5103);
nor U6458 (N_6458,N_5683,N_5638);
or U6459 (N_6459,N_5153,N_5692);
nor U6460 (N_6460,N_5957,N_5909);
nor U6461 (N_6461,N_5083,N_5795);
nand U6462 (N_6462,N_5945,N_5798);
or U6463 (N_6463,N_5837,N_5505);
nand U6464 (N_6464,N_5191,N_5714);
nand U6465 (N_6465,N_5493,N_5643);
nand U6466 (N_6466,N_5108,N_5163);
and U6467 (N_6467,N_5918,N_5267);
nand U6468 (N_6468,N_5884,N_5186);
and U6469 (N_6469,N_5834,N_5661);
nor U6470 (N_6470,N_5675,N_5971);
nor U6471 (N_6471,N_5917,N_5179);
nor U6472 (N_6472,N_5221,N_5100);
and U6473 (N_6473,N_5208,N_5037);
nand U6474 (N_6474,N_5421,N_5476);
and U6475 (N_6475,N_5370,N_5150);
or U6476 (N_6476,N_5228,N_5411);
xnor U6477 (N_6477,N_5943,N_5432);
nor U6478 (N_6478,N_5907,N_5760);
or U6479 (N_6479,N_5973,N_5616);
nor U6480 (N_6480,N_5574,N_5423);
xor U6481 (N_6481,N_5289,N_5288);
xor U6482 (N_6482,N_5906,N_5486);
nor U6483 (N_6483,N_5254,N_5938);
nand U6484 (N_6484,N_5822,N_5013);
nand U6485 (N_6485,N_5138,N_5356);
nor U6486 (N_6486,N_5663,N_5701);
or U6487 (N_6487,N_5654,N_5002);
and U6488 (N_6488,N_5213,N_5181);
nand U6489 (N_6489,N_5742,N_5309);
nand U6490 (N_6490,N_5671,N_5835);
or U6491 (N_6491,N_5771,N_5842);
xnor U6492 (N_6492,N_5741,N_5450);
and U6493 (N_6493,N_5139,N_5793);
nor U6494 (N_6494,N_5546,N_5564);
and U6495 (N_6495,N_5570,N_5527);
or U6496 (N_6496,N_5340,N_5354);
and U6497 (N_6497,N_5941,N_5672);
or U6498 (N_6498,N_5402,N_5919);
and U6499 (N_6499,N_5550,N_5608);
and U6500 (N_6500,N_5413,N_5280);
nor U6501 (N_6501,N_5387,N_5475);
nor U6502 (N_6502,N_5188,N_5355);
nand U6503 (N_6503,N_5764,N_5414);
and U6504 (N_6504,N_5980,N_5337);
nand U6505 (N_6505,N_5423,N_5624);
nor U6506 (N_6506,N_5139,N_5847);
nor U6507 (N_6507,N_5409,N_5174);
nand U6508 (N_6508,N_5034,N_5518);
nand U6509 (N_6509,N_5832,N_5164);
or U6510 (N_6510,N_5757,N_5646);
xor U6511 (N_6511,N_5592,N_5389);
and U6512 (N_6512,N_5159,N_5511);
and U6513 (N_6513,N_5474,N_5394);
nor U6514 (N_6514,N_5067,N_5288);
or U6515 (N_6515,N_5182,N_5281);
and U6516 (N_6516,N_5825,N_5571);
nand U6517 (N_6517,N_5550,N_5479);
and U6518 (N_6518,N_5761,N_5751);
nand U6519 (N_6519,N_5088,N_5684);
or U6520 (N_6520,N_5511,N_5488);
xnor U6521 (N_6521,N_5436,N_5220);
or U6522 (N_6522,N_5079,N_5666);
xnor U6523 (N_6523,N_5823,N_5523);
or U6524 (N_6524,N_5437,N_5105);
or U6525 (N_6525,N_5387,N_5512);
nor U6526 (N_6526,N_5257,N_5854);
nor U6527 (N_6527,N_5080,N_5432);
and U6528 (N_6528,N_5862,N_5504);
nand U6529 (N_6529,N_5709,N_5159);
nand U6530 (N_6530,N_5494,N_5701);
nand U6531 (N_6531,N_5109,N_5867);
xnor U6532 (N_6532,N_5636,N_5343);
nand U6533 (N_6533,N_5751,N_5146);
nand U6534 (N_6534,N_5454,N_5957);
or U6535 (N_6535,N_5949,N_5635);
or U6536 (N_6536,N_5940,N_5531);
and U6537 (N_6537,N_5448,N_5413);
xor U6538 (N_6538,N_5678,N_5673);
nor U6539 (N_6539,N_5934,N_5588);
nand U6540 (N_6540,N_5604,N_5127);
nor U6541 (N_6541,N_5063,N_5303);
and U6542 (N_6542,N_5416,N_5074);
xor U6543 (N_6543,N_5869,N_5930);
nor U6544 (N_6544,N_5457,N_5616);
nand U6545 (N_6545,N_5483,N_5967);
and U6546 (N_6546,N_5374,N_5001);
nand U6547 (N_6547,N_5376,N_5902);
nand U6548 (N_6548,N_5612,N_5318);
or U6549 (N_6549,N_5506,N_5169);
nand U6550 (N_6550,N_5119,N_5472);
xor U6551 (N_6551,N_5285,N_5939);
nand U6552 (N_6552,N_5793,N_5907);
and U6553 (N_6553,N_5007,N_5669);
nand U6554 (N_6554,N_5680,N_5008);
xnor U6555 (N_6555,N_5028,N_5626);
nand U6556 (N_6556,N_5016,N_5189);
nand U6557 (N_6557,N_5518,N_5707);
and U6558 (N_6558,N_5449,N_5082);
xor U6559 (N_6559,N_5375,N_5558);
nand U6560 (N_6560,N_5796,N_5966);
nor U6561 (N_6561,N_5058,N_5274);
nor U6562 (N_6562,N_5431,N_5931);
nand U6563 (N_6563,N_5081,N_5167);
nand U6564 (N_6564,N_5507,N_5529);
and U6565 (N_6565,N_5438,N_5235);
nand U6566 (N_6566,N_5542,N_5237);
nor U6567 (N_6567,N_5699,N_5907);
xor U6568 (N_6568,N_5692,N_5575);
or U6569 (N_6569,N_5165,N_5334);
and U6570 (N_6570,N_5582,N_5741);
nand U6571 (N_6571,N_5152,N_5877);
and U6572 (N_6572,N_5504,N_5572);
and U6573 (N_6573,N_5378,N_5120);
nand U6574 (N_6574,N_5840,N_5974);
nand U6575 (N_6575,N_5866,N_5629);
or U6576 (N_6576,N_5358,N_5097);
or U6577 (N_6577,N_5126,N_5981);
or U6578 (N_6578,N_5928,N_5852);
nor U6579 (N_6579,N_5615,N_5849);
or U6580 (N_6580,N_5242,N_5214);
and U6581 (N_6581,N_5107,N_5678);
or U6582 (N_6582,N_5309,N_5785);
nand U6583 (N_6583,N_5447,N_5590);
nor U6584 (N_6584,N_5641,N_5791);
and U6585 (N_6585,N_5434,N_5127);
or U6586 (N_6586,N_5796,N_5202);
and U6587 (N_6587,N_5606,N_5309);
nand U6588 (N_6588,N_5732,N_5479);
or U6589 (N_6589,N_5524,N_5681);
and U6590 (N_6590,N_5374,N_5877);
and U6591 (N_6591,N_5581,N_5620);
xor U6592 (N_6592,N_5365,N_5123);
or U6593 (N_6593,N_5091,N_5391);
xor U6594 (N_6594,N_5196,N_5134);
or U6595 (N_6595,N_5266,N_5301);
nand U6596 (N_6596,N_5439,N_5947);
and U6597 (N_6597,N_5525,N_5039);
nor U6598 (N_6598,N_5526,N_5359);
nand U6599 (N_6599,N_5561,N_5516);
nor U6600 (N_6600,N_5298,N_5330);
nor U6601 (N_6601,N_5300,N_5297);
nor U6602 (N_6602,N_5632,N_5857);
or U6603 (N_6603,N_5974,N_5577);
or U6604 (N_6604,N_5122,N_5240);
and U6605 (N_6605,N_5605,N_5088);
or U6606 (N_6606,N_5980,N_5052);
and U6607 (N_6607,N_5321,N_5081);
or U6608 (N_6608,N_5452,N_5480);
nand U6609 (N_6609,N_5696,N_5671);
nand U6610 (N_6610,N_5276,N_5748);
or U6611 (N_6611,N_5707,N_5465);
xnor U6612 (N_6612,N_5374,N_5936);
nand U6613 (N_6613,N_5949,N_5550);
nand U6614 (N_6614,N_5552,N_5684);
xor U6615 (N_6615,N_5051,N_5335);
nand U6616 (N_6616,N_5172,N_5755);
nor U6617 (N_6617,N_5961,N_5673);
nor U6618 (N_6618,N_5231,N_5340);
or U6619 (N_6619,N_5199,N_5782);
nand U6620 (N_6620,N_5216,N_5122);
nand U6621 (N_6621,N_5778,N_5389);
xor U6622 (N_6622,N_5937,N_5024);
or U6623 (N_6623,N_5302,N_5159);
nand U6624 (N_6624,N_5460,N_5842);
nor U6625 (N_6625,N_5306,N_5374);
nor U6626 (N_6626,N_5746,N_5335);
or U6627 (N_6627,N_5281,N_5849);
xnor U6628 (N_6628,N_5456,N_5661);
and U6629 (N_6629,N_5584,N_5577);
or U6630 (N_6630,N_5211,N_5066);
or U6631 (N_6631,N_5131,N_5217);
and U6632 (N_6632,N_5521,N_5942);
xnor U6633 (N_6633,N_5690,N_5706);
nand U6634 (N_6634,N_5200,N_5434);
nand U6635 (N_6635,N_5644,N_5772);
nor U6636 (N_6636,N_5613,N_5992);
or U6637 (N_6637,N_5579,N_5407);
and U6638 (N_6638,N_5841,N_5371);
or U6639 (N_6639,N_5423,N_5614);
nand U6640 (N_6640,N_5407,N_5255);
and U6641 (N_6641,N_5532,N_5339);
nand U6642 (N_6642,N_5630,N_5472);
or U6643 (N_6643,N_5051,N_5610);
nand U6644 (N_6644,N_5443,N_5361);
nor U6645 (N_6645,N_5224,N_5910);
nand U6646 (N_6646,N_5519,N_5184);
and U6647 (N_6647,N_5607,N_5237);
and U6648 (N_6648,N_5042,N_5050);
or U6649 (N_6649,N_5588,N_5563);
xor U6650 (N_6650,N_5209,N_5333);
or U6651 (N_6651,N_5600,N_5208);
and U6652 (N_6652,N_5143,N_5053);
nand U6653 (N_6653,N_5782,N_5423);
and U6654 (N_6654,N_5292,N_5296);
and U6655 (N_6655,N_5785,N_5450);
nor U6656 (N_6656,N_5331,N_5134);
nand U6657 (N_6657,N_5195,N_5365);
or U6658 (N_6658,N_5611,N_5572);
or U6659 (N_6659,N_5121,N_5156);
nand U6660 (N_6660,N_5397,N_5539);
nand U6661 (N_6661,N_5862,N_5032);
nor U6662 (N_6662,N_5239,N_5974);
or U6663 (N_6663,N_5207,N_5829);
nor U6664 (N_6664,N_5466,N_5911);
nor U6665 (N_6665,N_5847,N_5158);
and U6666 (N_6666,N_5898,N_5069);
and U6667 (N_6667,N_5549,N_5233);
xor U6668 (N_6668,N_5688,N_5624);
nor U6669 (N_6669,N_5003,N_5491);
or U6670 (N_6670,N_5186,N_5609);
nor U6671 (N_6671,N_5551,N_5775);
nand U6672 (N_6672,N_5286,N_5333);
nand U6673 (N_6673,N_5391,N_5448);
xor U6674 (N_6674,N_5695,N_5341);
or U6675 (N_6675,N_5360,N_5438);
xnor U6676 (N_6676,N_5867,N_5794);
nor U6677 (N_6677,N_5835,N_5712);
and U6678 (N_6678,N_5593,N_5087);
nor U6679 (N_6679,N_5446,N_5161);
and U6680 (N_6680,N_5807,N_5599);
nand U6681 (N_6681,N_5912,N_5181);
or U6682 (N_6682,N_5980,N_5797);
xor U6683 (N_6683,N_5545,N_5038);
and U6684 (N_6684,N_5876,N_5056);
nor U6685 (N_6685,N_5343,N_5640);
nand U6686 (N_6686,N_5684,N_5553);
nor U6687 (N_6687,N_5384,N_5363);
or U6688 (N_6688,N_5477,N_5156);
nand U6689 (N_6689,N_5895,N_5534);
xnor U6690 (N_6690,N_5940,N_5933);
or U6691 (N_6691,N_5775,N_5214);
nand U6692 (N_6692,N_5962,N_5539);
nand U6693 (N_6693,N_5685,N_5733);
and U6694 (N_6694,N_5482,N_5484);
xor U6695 (N_6695,N_5666,N_5089);
or U6696 (N_6696,N_5813,N_5105);
or U6697 (N_6697,N_5983,N_5436);
nand U6698 (N_6698,N_5021,N_5267);
xor U6699 (N_6699,N_5834,N_5483);
xor U6700 (N_6700,N_5710,N_5974);
nor U6701 (N_6701,N_5625,N_5186);
nand U6702 (N_6702,N_5514,N_5117);
or U6703 (N_6703,N_5189,N_5993);
nor U6704 (N_6704,N_5461,N_5517);
nor U6705 (N_6705,N_5275,N_5807);
and U6706 (N_6706,N_5903,N_5473);
and U6707 (N_6707,N_5000,N_5706);
and U6708 (N_6708,N_5881,N_5926);
or U6709 (N_6709,N_5819,N_5758);
nand U6710 (N_6710,N_5996,N_5524);
and U6711 (N_6711,N_5471,N_5336);
and U6712 (N_6712,N_5147,N_5050);
or U6713 (N_6713,N_5825,N_5367);
nor U6714 (N_6714,N_5324,N_5545);
nor U6715 (N_6715,N_5970,N_5350);
nor U6716 (N_6716,N_5891,N_5517);
xor U6717 (N_6717,N_5233,N_5037);
and U6718 (N_6718,N_5820,N_5052);
and U6719 (N_6719,N_5504,N_5839);
and U6720 (N_6720,N_5636,N_5395);
or U6721 (N_6721,N_5888,N_5826);
or U6722 (N_6722,N_5207,N_5602);
nor U6723 (N_6723,N_5524,N_5554);
or U6724 (N_6724,N_5392,N_5709);
nand U6725 (N_6725,N_5102,N_5710);
nand U6726 (N_6726,N_5741,N_5632);
and U6727 (N_6727,N_5694,N_5165);
nor U6728 (N_6728,N_5661,N_5316);
and U6729 (N_6729,N_5640,N_5307);
nor U6730 (N_6730,N_5100,N_5726);
nand U6731 (N_6731,N_5479,N_5061);
nand U6732 (N_6732,N_5006,N_5038);
xnor U6733 (N_6733,N_5005,N_5390);
nand U6734 (N_6734,N_5089,N_5579);
or U6735 (N_6735,N_5336,N_5330);
or U6736 (N_6736,N_5774,N_5495);
nor U6737 (N_6737,N_5427,N_5451);
or U6738 (N_6738,N_5953,N_5669);
and U6739 (N_6739,N_5165,N_5516);
nand U6740 (N_6740,N_5391,N_5231);
or U6741 (N_6741,N_5617,N_5210);
nor U6742 (N_6742,N_5385,N_5080);
and U6743 (N_6743,N_5128,N_5968);
nand U6744 (N_6744,N_5220,N_5118);
and U6745 (N_6745,N_5061,N_5011);
or U6746 (N_6746,N_5058,N_5528);
or U6747 (N_6747,N_5806,N_5980);
xor U6748 (N_6748,N_5212,N_5346);
or U6749 (N_6749,N_5720,N_5405);
or U6750 (N_6750,N_5475,N_5601);
and U6751 (N_6751,N_5766,N_5146);
or U6752 (N_6752,N_5396,N_5155);
or U6753 (N_6753,N_5112,N_5413);
nand U6754 (N_6754,N_5451,N_5016);
xor U6755 (N_6755,N_5007,N_5591);
or U6756 (N_6756,N_5137,N_5882);
nor U6757 (N_6757,N_5005,N_5107);
and U6758 (N_6758,N_5671,N_5131);
nor U6759 (N_6759,N_5360,N_5003);
nand U6760 (N_6760,N_5388,N_5602);
or U6761 (N_6761,N_5910,N_5207);
nand U6762 (N_6762,N_5154,N_5428);
nor U6763 (N_6763,N_5638,N_5808);
or U6764 (N_6764,N_5021,N_5473);
and U6765 (N_6765,N_5939,N_5872);
and U6766 (N_6766,N_5729,N_5400);
and U6767 (N_6767,N_5275,N_5693);
nand U6768 (N_6768,N_5454,N_5414);
and U6769 (N_6769,N_5876,N_5519);
nor U6770 (N_6770,N_5726,N_5302);
nand U6771 (N_6771,N_5007,N_5458);
nand U6772 (N_6772,N_5971,N_5088);
nand U6773 (N_6773,N_5454,N_5580);
or U6774 (N_6774,N_5302,N_5540);
or U6775 (N_6775,N_5993,N_5759);
nor U6776 (N_6776,N_5194,N_5579);
nand U6777 (N_6777,N_5715,N_5085);
or U6778 (N_6778,N_5971,N_5589);
and U6779 (N_6779,N_5821,N_5748);
nor U6780 (N_6780,N_5191,N_5981);
nand U6781 (N_6781,N_5462,N_5130);
nor U6782 (N_6782,N_5556,N_5097);
xor U6783 (N_6783,N_5620,N_5186);
or U6784 (N_6784,N_5222,N_5289);
nand U6785 (N_6785,N_5760,N_5851);
and U6786 (N_6786,N_5811,N_5661);
nor U6787 (N_6787,N_5939,N_5525);
or U6788 (N_6788,N_5640,N_5098);
nand U6789 (N_6789,N_5402,N_5666);
or U6790 (N_6790,N_5254,N_5409);
nand U6791 (N_6791,N_5001,N_5297);
nand U6792 (N_6792,N_5624,N_5978);
nand U6793 (N_6793,N_5466,N_5873);
nand U6794 (N_6794,N_5433,N_5601);
or U6795 (N_6795,N_5211,N_5496);
nand U6796 (N_6796,N_5166,N_5588);
or U6797 (N_6797,N_5994,N_5939);
nand U6798 (N_6798,N_5519,N_5058);
nor U6799 (N_6799,N_5872,N_5825);
or U6800 (N_6800,N_5065,N_5602);
or U6801 (N_6801,N_5335,N_5605);
nand U6802 (N_6802,N_5253,N_5248);
or U6803 (N_6803,N_5188,N_5899);
or U6804 (N_6804,N_5529,N_5516);
and U6805 (N_6805,N_5877,N_5652);
nor U6806 (N_6806,N_5198,N_5662);
and U6807 (N_6807,N_5209,N_5947);
nand U6808 (N_6808,N_5900,N_5655);
and U6809 (N_6809,N_5510,N_5983);
or U6810 (N_6810,N_5387,N_5746);
nor U6811 (N_6811,N_5525,N_5084);
and U6812 (N_6812,N_5380,N_5726);
and U6813 (N_6813,N_5288,N_5688);
or U6814 (N_6814,N_5077,N_5179);
or U6815 (N_6815,N_5118,N_5683);
nand U6816 (N_6816,N_5437,N_5196);
or U6817 (N_6817,N_5953,N_5004);
nand U6818 (N_6818,N_5600,N_5730);
and U6819 (N_6819,N_5524,N_5270);
nor U6820 (N_6820,N_5597,N_5628);
nand U6821 (N_6821,N_5593,N_5432);
nor U6822 (N_6822,N_5761,N_5981);
nor U6823 (N_6823,N_5964,N_5610);
and U6824 (N_6824,N_5524,N_5352);
xnor U6825 (N_6825,N_5657,N_5017);
xor U6826 (N_6826,N_5281,N_5549);
nand U6827 (N_6827,N_5646,N_5593);
and U6828 (N_6828,N_5609,N_5763);
or U6829 (N_6829,N_5689,N_5815);
nor U6830 (N_6830,N_5622,N_5252);
nor U6831 (N_6831,N_5604,N_5693);
or U6832 (N_6832,N_5658,N_5113);
nand U6833 (N_6833,N_5430,N_5516);
nand U6834 (N_6834,N_5390,N_5200);
nor U6835 (N_6835,N_5852,N_5110);
and U6836 (N_6836,N_5016,N_5506);
or U6837 (N_6837,N_5664,N_5905);
and U6838 (N_6838,N_5267,N_5938);
or U6839 (N_6839,N_5987,N_5066);
xnor U6840 (N_6840,N_5826,N_5914);
or U6841 (N_6841,N_5905,N_5966);
nor U6842 (N_6842,N_5780,N_5462);
nor U6843 (N_6843,N_5357,N_5844);
and U6844 (N_6844,N_5954,N_5276);
nand U6845 (N_6845,N_5441,N_5253);
nor U6846 (N_6846,N_5949,N_5753);
nor U6847 (N_6847,N_5454,N_5199);
nand U6848 (N_6848,N_5290,N_5967);
nor U6849 (N_6849,N_5489,N_5111);
or U6850 (N_6850,N_5358,N_5721);
or U6851 (N_6851,N_5632,N_5123);
and U6852 (N_6852,N_5735,N_5019);
or U6853 (N_6853,N_5057,N_5841);
and U6854 (N_6854,N_5366,N_5738);
nand U6855 (N_6855,N_5466,N_5297);
xor U6856 (N_6856,N_5289,N_5113);
and U6857 (N_6857,N_5040,N_5190);
nand U6858 (N_6858,N_5531,N_5846);
nand U6859 (N_6859,N_5280,N_5083);
nand U6860 (N_6860,N_5924,N_5061);
or U6861 (N_6861,N_5755,N_5034);
nand U6862 (N_6862,N_5832,N_5382);
or U6863 (N_6863,N_5858,N_5521);
or U6864 (N_6864,N_5696,N_5189);
xnor U6865 (N_6865,N_5223,N_5878);
xnor U6866 (N_6866,N_5836,N_5614);
nor U6867 (N_6867,N_5702,N_5496);
or U6868 (N_6868,N_5781,N_5548);
and U6869 (N_6869,N_5976,N_5276);
xor U6870 (N_6870,N_5856,N_5872);
nor U6871 (N_6871,N_5873,N_5163);
nor U6872 (N_6872,N_5130,N_5931);
xor U6873 (N_6873,N_5480,N_5949);
nor U6874 (N_6874,N_5516,N_5854);
or U6875 (N_6875,N_5370,N_5382);
or U6876 (N_6876,N_5463,N_5714);
and U6877 (N_6877,N_5682,N_5298);
or U6878 (N_6878,N_5670,N_5029);
xnor U6879 (N_6879,N_5070,N_5527);
nand U6880 (N_6880,N_5929,N_5572);
nand U6881 (N_6881,N_5609,N_5389);
and U6882 (N_6882,N_5365,N_5716);
or U6883 (N_6883,N_5407,N_5236);
nand U6884 (N_6884,N_5500,N_5887);
or U6885 (N_6885,N_5743,N_5725);
or U6886 (N_6886,N_5154,N_5856);
xnor U6887 (N_6887,N_5355,N_5722);
nor U6888 (N_6888,N_5802,N_5578);
nor U6889 (N_6889,N_5201,N_5948);
and U6890 (N_6890,N_5565,N_5259);
and U6891 (N_6891,N_5805,N_5995);
and U6892 (N_6892,N_5665,N_5354);
or U6893 (N_6893,N_5270,N_5454);
nor U6894 (N_6894,N_5643,N_5674);
or U6895 (N_6895,N_5065,N_5783);
nand U6896 (N_6896,N_5382,N_5037);
nor U6897 (N_6897,N_5122,N_5721);
nor U6898 (N_6898,N_5478,N_5331);
or U6899 (N_6899,N_5089,N_5182);
nand U6900 (N_6900,N_5558,N_5272);
xnor U6901 (N_6901,N_5057,N_5169);
or U6902 (N_6902,N_5049,N_5552);
nor U6903 (N_6903,N_5967,N_5730);
or U6904 (N_6904,N_5735,N_5118);
nor U6905 (N_6905,N_5813,N_5601);
nor U6906 (N_6906,N_5304,N_5432);
nand U6907 (N_6907,N_5339,N_5527);
xor U6908 (N_6908,N_5494,N_5118);
or U6909 (N_6909,N_5129,N_5683);
nand U6910 (N_6910,N_5926,N_5016);
nor U6911 (N_6911,N_5461,N_5829);
xnor U6912 (N_6912,N_5096,N_5648);
nand U6913 (N_6913,N_5104,N_5798);
or U6914 (N_6914,N_5526,N_5676);
nor U6915 (N_6915,N_5860,N_5894);
and U6916 (N_6916,N_5659,N_5809);
xnor U6917 (N_6917,N_5132,N_5328);
nor U6918 (N_6918,N_5790,N_5090);
and U6919 (N_6919,N_5324,N_5014);
or U6920 (N_6920,N_5232,N_5569);
or U6921 (N_6921,N_5824,N_5148);
nand U6922 (N_6922,N_5914,N_5864);
nor U6923 (N_6923,N_5151,N_5019);
or U6924 (N_6924,N_5851,N_5714);
nand U6925 (N_6925,N_5294,N_5504);
nor U6926 (N_6926,N_5187,N_5103);
or U6927 (N_6927,N_5867,N_5416);
nor U6928 (N_6928,N_5662,N_5651);
or U6929 (N_6929,N_5692,N_5623);
or U6930 (N_6930,N_5165,N_5252);
or U6931 (N_6931,N_5625,N_5099);
or U6932 (N_6932,N_5409,N_5508);
and U6933 (N_6933,N_5363,N_5930);
and U6934 (N_6934,N_5375,N_5478);
nor U6935 (N_6935,N_5093,N_5974);
nor U6936 (N_6936,N_5368,N_5326);
xnor U6937 (N_6937,N_5775,N_5176);
nand U6938 (N_6938,N_5711,N_5971);
nor U6939 (N_6939,N_5926,N_5584);
and U6940 (N_6940,N_5971,N_5521);
nor U6941 (N_6941,N_5006,N_5140);
nor U6942 (N_6942,N_5549,N_5753);
or U6943 (N_6943,N_5281,N_5411);
or U6944 (N_6944,N_5164,N_5941);
xor U6945 (N_6945,N_5695,N_5375);
nand U6946 (N_6946,N_5140,N_5339);
nand U6947 (N_6947,N_5716,N_5465);
and U6948 (N_6948,N_5365,N_5350);
xnor U6949 (N_6949,N_5802,N_5072);
nand U6950 (N_6950,N_5739,N_5303);
and U6951 (N_6951,N_5553,N_5604);
xor U6952 (N_6952,N_5964,N_5545);
or U6953 (N_6953,N_5190,N_5206);
or U6954 (N_6954,N_5945,N_5066);
xnor U6955 (N_6955,N_5650,N_5936);
or U6956 (N_6956,N_5581,N_5666);
and U6957 (N_6957,N_5124,N_5643);
xnor U6958 (N_6958,N_5252,N_5730);
or U6959 (N_6959,N_5266,N_5537);
nor U6960 (N_6960,N_5116,N_5429);
nor U6961 (N_6961,N_5292,N_5931);
or U6962 (N_6962,N_5050,N_5956);
and U6963 (N_6963,N_5296,N_5616);
nand U6964 (N_6964,N_5446,N_5559);
and U6965 (N_6965,N_5222,N_5215);
nor U6966 (N_6966,N_5453,N_5349);
nor U6967 (N_6967,N_5873,N_5094);
nand U6968 (N_6968,N_5941,N_5260);
nand U6969 (N_6969,N_5569,N_5123);
nand U6970 (N_6970,N_5657,N_5416);
or U6971 (N_6971,N_5597,N_5271);
or U6972 (N_6972,N_5401,N_5737);
nor U6973 (N_6973,N_5811,N_5211);
xor U6974 (N_6974,N_5555,N_5331);
or U6975 (N_6975,N_5447,N_5308);
and U6976 (N_6976,N_5136,N_5446);
nor U6977 (N_6977,N_5225,N_5830);
nand U6978 (N_6978,N_5406,N_5586);
or U6979 (N_6979,N_5956,N_5409);
or U6980 (N_6980,N_5813,N_5737);
and U6981 (N_6981,N_5416,N_5553);
nor U6982 (N_6982,N_5045,N_5566);
xor U6983 (N_6983,N_5644,N_5518);
nor U6984 (N_6984,N_5052,N_5377);
or U6985 (N_6985,N_5500,N_5997);
xnor U6986 (N_6986,N_5284,N_5493);
and U6987 (N_6987,N_5323,N_5745);
nor U6988 (N_6988,N_5112,N_5208);
nand U6989 (N_6989,N_5799,N_5622);
and U6990 (N_6990,N_5529,N_5933);
nand U6991 (N_6991,N_5260,N_5424);
and U6992 (N_6992,N_5146,N_5999);
or U6993 (N_6993,N_5249,N_5976);
nor U6994 (N_6994,N_5817,N_5103);
and U6995 (N_6995,N_5031,N_5158);
and U6996 (N_6996,N_5309,N_5422);
and U6997 (N_6997,N_5012,N_5321);
and U6998 (N_6998,N_5533,N_5057);
nor U6999 (N_6999,N_5976,N_5271);
nand U7000 (N_7000,N_6326,N_6905);
nand U7001 (N_7001,N_6957,N_6968);
xor U7002 (N_7002,N_6658,N_6087);
or U7003 (N_7003,N_6132,N_6440);
nor U7004 (N_7004,N_6412,N_6312);
nor U7005 (N_7005,N_6064,N_6702);
xor U7006 (N_7006,N_6993,N_6677);
nor U7007 (N_7007,N_6519,N_6981);
xnor U7008 (N_7008,N_6305,N_6644);
nor U7009 (N_7009,N_6118,N_6296);
nor U7010 (N_7010,N_6217,N_6767);
nor U7011 (N_7011,N_6545,N_6816);
nand U7012 (N_7012,N_6778,N_6261);
nand U7013 (N_7013,N_6589,N_6593);
or U7014 (N_7014,N_6079,N_6980);
nor U7015 (N_7015,N_6600,N_6735);
and U7016 (N_7016,N_6060,N_6220);
and U7017 (N_7017,N_6512,N_6153);
xnor U7018 (N_7018,N_6035,N_6863);
and U7019 (N_7019,N_6002,N_6299);
nand U7020 (N_7020,N_6129,N_6345);
and U7021 (N_7021,N_6401,N_6994);
xnor U7022 (N_7022,N_6294,N_6173);
and U7023 (N_7023,N_6478,N_6361);
nand U7024 (N_7024,N_6694,N_6056);
or U7025 (N_7025,N_6280,N_6094);
nor U7026 (N_7026,N_6075,N_6281);
or U7027 (N_7027,N_6055,N_6530);
nand U7028 (N_7028,N_6329,N_6721);
nor U7029 (N_7029,N_6543,N_6167);
nor U7030 (N_7030,N_6308,N_6154);
or U7031 (N_7031,N_6469,N_6383);
nand U7032 (N_7032,N_6643,N_6573);
nor U7033 (N_7033,N_6441,N_6244);
nand U7034 (N_7034,N_6230,N_6316);
and U7035 (N_7035,N_6824,N_6013);
or U7036 (N_7036,N_6546,N_6366);
nand U7037 (N_7037,N_6459,N_6609);
or U7038 (N_7038,N_6920,N_6912);
nand U7039 (N_7039,N_6311,N_6632);
and U7040 (N_7040,N_6458,N_6391);
xnor U7041 (N_7041,N_6904,N_6768);
and U7042 (N_7042,N_6697,N_6488);
or U7043 (N_7043,N_6327,N_6286);
xor U7044 (N_7044,N_6836,N_6695);
nand U7045 (N_7045,N_6734,N_6936);
or U7046 (N_7046,N_6036,N_6707);
and U7047 (N_7047,N_6078,N_6477);
and U7048 (N_7048,N_6590,N_6524);
nand U7049 (N_7049,N_6647,N_6626);
or U7050 (N_7050,N_6787,N_6684);
nand U7051 (N_7051,N_6942,N_6017);
nand U7052 (N_7052,N_6319,N_6430);
nand U7053 (N_7053,N_6974,N_6499);
nor U7054 (N_7054,N_6948,N_6330);
or U7055 (N_7055,N_6359,N_6551);
nand U7056 (N_7056,N_6645,N_6601);
nor U7057 (N_7057,N_6983,N_6683);
and U7058 (N_7058,N_6933,N_6031);
and U7059 (N_7059,N_6322,N_6240);
nand U7060 (N_7060,N_6679,N_6771);
nand U7061 (N_7061,N_6856,N_6029);
nand U7062 (N_7062,N_6548,N_6318);
nand U7063 (N_7063,N_6045,N_6009);
and U7064 (N_7064,N_6197,N_6791);
or U7065 (N_7065,N_6368,N_6072);
xnor U7066 (N_7066,N_6229,N_6222);
and U7067 (N_7067,N_6585,N_6049);
nand U7068 (N_7068,N_6001,N_6067);
and U7069 (N_7069,N_6565,N_6352);
xor U7070 (N_7070,N_6044,N_6012);
nor U7071 (N_7071,N_6736,N_6803);
or U7072 (N_7072,N_6396,N_6509);
and U7073 (N_7073,N_6150,N_6579);
or U7074 (N_7074,N_6860,N_6878);
xnor U7075 (N_7075,N_6608,N_6131);
nor U7076 (N_7076,N_6429,N_6192);
nand U7077 (N_7077,N_6642,N_6757);
and U7078 (N_7078,N_6789,N_6179);
nor U7079 (N_7079,N_6358,N_6233);
nor U7080 (N_7080,N_6706,N_6283);
and U7081 (N_7081,N_6769,N_6404);
or U7082 (N_7082,N_6076,N_6620);
nor U7083 (N_7083,N_6680,N_6575);
and U7084 (N_7084,N_6894,N_6428);
or U7085 (N_7085,N_6723,N_6583);
and U7086 (N_7086,N_6651,N_6526);
nand U7087 (N_7087,N_6491,N_6451);
and U7088 (N_7088,N_6869,N_6264);
or U7089 (N_7089,N_6203,N_6796);
or U7090 (N_7090,N_6105,N_6051);
or U7091 (N_7091,N_6402,N_6985);
nand U7092 (N_7092,N_6117,N_6390);
nor U7093 (N_7093,N_6048,N_6270);
nor U7094 (N_7094,N_6300,N_6156);
or U7095 (N_7095,N_6603,N_6745);
nor U7096 (N_7096,N_6040,N_6959);
or U7097 (N_7097,N_6748,N_6168);
and U7098 (N_7098,N_6895,N_6475);
or U7099 (N_7099,N_6191,N_6272);
nor U7100 (N_7100,N_6618,N_6938);
xor U7101 (N_7101,N_6147,N_6092);
and U7102 (N_7102,N_6303,N_6490);
or U7103 (N_7103,N_6450,N_6982);
nand U7104 (N_7104,N_6825,N_6722);
or U7105 (N_7105,N_6393,N_6285);
or U7106 (N_7106,N_6761,N_6908);
nand U7107 (N_7107,N_6849,N_6143);
or U7108 (N_7108,N_6082,N_6937);
and U7109 (N_7109,N_6689,N_6950);
nand U7110 (N_7110,N_6766,N_6262);
or U7111 (N_7111,N_6328,N_6069);
nor U7112 (N_7112,N_6443,N_6570);
nand U7113 (N_7113,N_6587,N_6742);
xnor U7114 (N_7114,N_6198,N_6447);
and U7115 (N_7115,N_6978,N_6255);
nand U7116 (N_7116,N_6452,N_6639);
nor U7117 (N_7117,N_6989,N_6606);
or U7118 (N_7118,N_6988,N_6159);
and U7119 (N_7119,N_6425,N_6562);
nor U7120 (N_7120,N_6622,N_6185);
nand U7121 (N_7121,N_6884,N_6335);
nor U7122 (N_7122,N_6292,N_6817);
nand U7123 (N_7123,N_6657,N_6710);
xor U7124 (N_7124,N_6759,N_6896);
or U7125 (N_7125,N_6794,N_6193);
nand U7126 (N_7126,N_6612,N_6419);
xor U7127 (N_7127,N_6518,N_6627);
nor U7128 (N_7128,N_6151,N_6660);
nand U7129 (N_7129,N_6200,N_6254);
and U7130 (N_7130,N_6032,N_6614);
nor U7131 (N_7131,N_6915,N_6077);
nor U7132 (N_7132,N_6139,N_6389);
or U7133 (N_7133,N_6448,N_6288);
or U7134 (N_7134,N_6539,N_6212);
nor U7135 (N_7135,N_6411,N_6061);
or U7136 (N_7136,N_6636,N_6181);
nand U7137 (N_7137,N_6323,N_6779);
and U7138 (N_7138,N_6176,N_6542);
nor U7139 (N_7139,N_6619,N_6028);
nand U7140 (N_7140,N_6549,N_6165);
xnor U7141 (N_7141,N_6422,N_6089);
nand U7142 (N_7142,N_6175,N_6030);
or U7143 (N_7143,N_6487,N_6834);
nor U7144 (N_7144,N_6456,N_6416);
or U7145 (N_7145,N_6071,N_6865);
nand U7146 (N_7146,N_6113,N_6484);
and U7147 (N_7147,N_6298,N_6819);
nor U7148 (N_7148,N_6979,N_6841);
nand U7149 (N_7149,N_6837,N_6238);
and U7150 (N_7150,N_6195,N_6693);
and U7151 (N_7151,N_6126,N_6604);
and U7152 (N_7152,N_6502,N_6967);
or U7153 (N_7153,N_6672,N_6146);
nor U7154 (N_7154,N_6741,N_6558);
and U7155 (N_7155,N_6189,N_6027);
and U7156 (N_7156,N_6571,N_6753);
nand U7157 (N_7157,N_6828,N_6304);
and U7158 (N_7158,N_6461,N_6498);
nor U7159 (N_7159,N_6770,N_6387);
nor U7160 (N_7160,N_6553,N_6325);
and U7161 (N_7161,N_6861,N_6394);
or U7162 (N_7162,N_6569,N_6940);
nand U7163 (N_7163,N_6754,N_6395);
nor U7164 (N_7164,N_6893,N_6317);
or U7165 (N_7165,N_6501,N_6455);
nand U7166 (N_7166,N_6918,N_6821);
and U7167 (N_7167,N_6172,N_6804);
or U7168 (N_7168,N_6972,N_6005);
and U7169 (N_7169,N_6624,N_6144);
xnor U7170 (N_7170,N_6122,N_6662);
nor U7171 (N_7171,N_6091,N_6762);
nand U7172 (N_7172,N_6833,N_6862);
nor U7173 (N_7173,N_6084,N_6287);
nand U7174 (N_7174,N_6476,N_6987);
and U7175 (N_7175,N_6177,N_6696);
and U7176 (N_7176,N_6112,N_6617);
nand U7177 (N_7177,N_6164,N_6170);
nor U7178 (N_7178,N_6302,N_6634);
and U7179 (N_7179,N_6483,N_6535);
and U7180 (N_7180,N_6874,N_6661);
nand U7181 (N_7181,N_6086,N_6221);
nand U7182 (N_7182,N_6714,N_6307);
or U7183 (N_7183,N_6652,N_6656);
and U7184 (N_7184,N_6041,N_6909);
and U7185 (N_7185,N_6043,N_6764);
or U7186 (N_7186,N_6253,N_6554);
and U7187 (N_7187,N_6227,N_6251);
xor U7188 (N_7188,N_6310,N_6276);
nor U7189 (N_7189,N_6557,N_6047);
nand U7190 (N_7190,N_6591,N_6149);
nor U7191 (N_7191,N_6093,N_6206);
and U7192 (N_7192,N_6248,N_6665);
nand U7193 (N_7193,N_6566,N_6119);
or U7194 (N_7194,N_6355,N_6011);
nand U7195 (N_7195,N_6730,N_6977);
nor U7196 (N_7196,N_6740,N_6641);
or U7197 (N_7197,N_6482,N_6635);
or U7198 (N_7198,N_6353,N_6410);
nor U7199 (N_7199,N_6866,N_6289);
nand U7200 (N_7200,N_6962,N_6941);
nand U7201 (N_7201,N_6823,N_6555);
nor U7202 (N_7202,N_6463,N_6415);
xnor U7203 (N_7203,N_6236,N_6439);
xnor U7204 (N_7204,N_6529,N_6360);
and U7205 (N_7205,N_6128,N_6413);
nor U7206 (N_7206,N_6597,N_6595);
nor U7207 (N_7207,N_6399,N_6965);
or U7208 (N_7208,N_6515,N_6900);
and U7209 (N_7209,N_6324,N_6898);
and U7210 (N_7210,N_6855,N_6805);
or U7211 (N_7211,N_6659,N_6674);
and U7212 (N_7212,N_6525,N_6417);
nand U7213 (N_7213,N_6375,N_6125);
and U7214 (N_7214,N_6010,N_6961);
nand U7215 (N_7215,N_6725,N_6704);
or U7216 (N_7216,N_6370,N_6247);
nand U7217 (N_7217,N_6552,N_6685);
nor U7218 (N_7218,N_6398,N_6921);
and U7219 (N_7219,N_6582,N_6998);
nor U7220 (N_7220,N_6277,N_6629);
nand U7221 (N_7221,N_6882,N_6784);
nor U7222 (N_7222,N_6932,N_6135);
nor U7223 (N_7223,N_6931,N_6239);
or U7224 (N_7224,N_6640,N_6331);
nand U7225 (N_7225,N_6521,N_6424);
or U7226 (N_7226,N_6205,N_6169);
and U7227 (N_7227,N_6342,N_6357);
nand U7228 (N_7228,N_6480,N_6717);
or U7229 (N_7229,N_6103,N_6219);
nand U7230 (N_7230,N_6148,N_6949);
xnor U7231 (N_7231,N_6400,N_6916);
nand U7232 (N_7232,N_6100,N_6663);
nand U7233 (N_7233,N_6738,N_6199);
xor U7234 (N_7234,N_6607,N_6839);
nand U7235 (N_7235,N_6442,N_6210);
or U7236 (N_7236,N_6653,N_6688);
nand U7237 (N_7237,N_6881,N_6201);
nor U7238 (N_7238,N_6260,N_6503);
and U7239 (N_7239,N_6927,N_6615);
or U7240 (N_7240,N_6265,N_6892);
nand U7241 (N_7241,N_6226,N_6133);
xor U7242 (N_7242,N_6196,N_6510);
xnor U7243 (N_7243,N_6504,N_6719);
xnor U7244 (N_7244,N_6777,N_6848);
and U7245 (N_7245,N_6374,N_6901);
nor U7246 (N_7246,N_6602,N_6580);
and U7247 (N_7247,N_6667,N_6666);
nand U7248 (N_7248,N_6388,N_6726);
and U7249 (N_7249,N_6885,N_6246);
nor U7250 (N_7250,N_6405,N_6621);
nor U7251 (N_7251,N_6788,N_6765);
or U7252 (N_7252,N_6715,N_6356);
or U7253 (N_7253,N_6925,N_6373);
nor U7254 (N_7254,N_6145,N_6000);
or U7255 (N_7255,N_6245,N_6747);
nand U7256 (N_7256,N_6990,N_6868);
and U7257 (N_7257,N_6372,N_6397);
nand U7258 (N_7258,N_6806,N_6379);
nand U7259 (N_7259,N_6252,N_6369);
nand U7260 (N_7260,N_6107,N_6709);
nand U7261 (N_7261,N_6971,N_6537);
or U7262 (N_7262,N_6208,N_6190);
nand U7263 (N_7263,N_6268,N_6992);
nand U7264 (N_7264,N_6024,N_6584);
and U7265 (N_7265,N_6790,N_6489);
nor U7266 (N_7266,N_6025,N_6237);
xor U7267 (N_7267,N_6004,N_6454);
nor U7268 (N_7268,N_6003,N_6907);
nand U7269 (N_7269,N_6140,N_6313);
or U7270 (N_7270,N_6382,N_6158);
or U7271 (N_7271,N_6426,N_6633);
and U7272 (N_7272,N_6188,N_6339);
nor U7273 (N_7273,N_6801,N_6130);
nand U7274 (N_7274,N_6115,N_6121);
or U7275 (N_7275,N_6081,N_6864);
or U7276 (N_7276,N_6872,N_6728);
or U7277 (N_7277,N_6564,N_6586);
and U7278 (N_7278,N_6871,N_6610);
and U7279 (N_7279,N_6913,N_6963);
nand U7280 (N_7280,N_6711,N_6984);
nor U7281 (N_7281,N_6337,N_6724);
nand U7282 (N_7282,N_6059,N_6054);
nand U7283 (N_7283,N_6160,N_6997);
and U7284 (N_7284,N_6321,N_6531);
and U7285 (N_7285,N_6257,N_6567);
and U7286 (N_7286,N_6473,N_6223);
and U7287 (N_7287,N_6123,N_6336);
nor U7288 (N_7288,N_6433,N_6832);
or U7289 (N_7289,N_6334,N_6678);
and U7290 (N_7290,N_6471,N_6453);
or U7291 (N_7291,N_6939,N_6023);
and U7292 (N_7292,N_6496,N_6654);
nand U7293 (N_7293,N_6034,N_6814);
nand U7294 (N_7294,N_6810,N_6038);
and U7295 (N_7295,N_6014,N_6141);
or U7296 (N_7296,N_6842,N_6467);
xnor U7297 (N_7297,N_6780,N_6058);
nand U7298 (N_7298,N_6457,N_6544);
or U7299 (N_7299,N_6508,N_6827);
and U7300 (N_7300,N_6242,N_6377);
xor U7301 (N_7301,N_6134,N_6279);
nand U7302 (N_7302,N_6802,N_6042);
and U7303 (N_7303,N_6380,N_6187);
or U7304 (N_7304,N_6256,N_6267);
or U7305 (N_7305,N_6955,N_6446);
or U7306 (N_7306,N_6444,N_6018);
or U7307 (N_7307,N_6668,N_6171);
or U7308 (N_7308,N_6225,N_6138);
nand U7309 (N_7309,N_6516,N_6563);
nor U7310 (N_7310,N_6338,N_6533);
nor U7311 (N_7311,N_6935,N_6231);
or U7312 (N_7312,N_6408,N_6818);
or U7313 (N_7313,N_6623,N_6495);
or U7314 (N_7314,N_6110,N_6690);
nor U7315 (N_7315,N_6068,N_6578);
nand U7316 (N_7316,N_6792,N_6975);
nand U7317 (N_7317,N_6224,N_6592);
nand U7318 (N_7318,N_6161,N_6873);
and U7319 (N_7319,N_6681,N_6449);
or U7320 (N_7320,N_6846,N_6731);
and U7321 (N_7321,N_6120,N_6924);
and U7322 (N_7322,N_6781,N_6434);
and U7323 (N_7323,N_6877,N_6271);
xnor U7324 (N_7324,N_6859,N_6840);
and U7325 (N_7325,N_6407,N_6057);
or U7326 (N_7326,N_6556,N_6887);
nor U7327 (N_7327,N_6088,N_6070);
nand U7328 (N_7328,N_6956,N_6136);
nand U7329 (N_7329,N_6204,N_6384);
nand U7330 (N_7330,N_6637,N_6184);
and U7331 (N_7331,N_6782,N_6258);
or U7332 (N_7332,N_6889,N_6514);
xor U7333 (N_7333,N_6462,N_6275);
and U7334 (N_7334,N_6291,N_6934);
and U7335 (N_7335,N_6729,N_6216);
or U7336 (N_7336,N_6309,N_6232);
xnor U7337 (N_7337,N_6616,N_6347);
and U7338 (N_7338,N_6970,N_6507);
nand U7339 (N_7339,N_6050,N_6273);
nand U7340 (N_7340,N_6795,N_6333);
nand U7341 (N_7341,N_6180,N_6737);
and U7342 (N_7342,N_6891,N_6700);
nor U7343 (N_7343,N_6218,N_6016);
and U7344 (N_7344,N_6142,N_6576);
and U7345 (N_7345,N_6914,N_6080);
and U7346 (N_7346,N_6964,N_6421);
nand U7347 (N_7347,N_6182,N_6406);
xor U7348 (N_7348,N_6116,N_6207);
nand U7349 (N_7349,N_6815,N_6437);
and U7350 (N_7350,N_6705,N_6703);
nor U7351 (N_7351,N_6611,N_6235);
nand U7352 (N_7352,N_6763,N_6822);
nor U7353 (N_7353,N_6718,N_6344);
nand U7354 (N_7354,N_6854,N_6926);
nor U7355 (N_7355,N_6346,N_6249);
nor U7356 (N_7356,N_6708,N_6538);
nand U7357 (N_7357,N_6673,N_6157);
nor U7358 (N_7358,N_6492,N_6098);
nand U7359 (N_7359,N_6432,N_6186);
or U7360 (N_7360,N_6090,N_6183);
and U7361 (N_7361,N_6111,N_6445);
or U7362 (N_7362,N_6365,N_6494);
xor U7363 (N_7363,N_6493,N_6019);
or U7364 (N_7364,N_6341,N_6386);
and U7365 (N_7365,N_6743,N_6958);
and U7366 (N_7366,N_6420,N_6883);
or U7367 (N_7367,N_6851,N_6845);
nor U7368 (N_7368,N_6101,N_6460);
nor U7369 (N_7369,N_6945,N_6954);
nor U7370 (N_7370,N_6867,N_6888);
xnor U7371 (N_7371,N_6340,N_6550);
or U7372 (N_7372,N_6362,N_6811);
and U7373 (N_7373,N_6250,N_6650);
xor U7374 (N_7374,N_6969,N_6698);
or U7375 (N_7375,N_6099,N_6911);
nand U7376 (N_7376,N_6760,N_6381);
xnor U7377 (N_7377,N_6066,N_6108);
and U7378 (N_7378,N_6033,N_6943);
nor U7379 (N_7379,N_6194,N_6174);
nor U7380 (N_7380,N_6843,N_6798);
and U7381 (N_7381,N_6500,N_6732);
nand U7382 (N_7382,N_6613,N_6349);
or U7383 (N_7383,N_6751,N_6773);
nand U7384 (N_7384,N_6712,N_6414);
nand U7385 (N_7385,N_6039,N_6472);
nor U7386 (N_7386,N_6857,N_6713);
or U7387 (N_7387,N_6063,N_6692);
nand U7388 (N_7388,N_6351,N_6096);
nand U7389 (N_7389,N_6991,N_6435);
nand U7390 (N_7390,N_6953,N_6561);
and U7391 (N_7391,N_6572,N_6106);
or U7392 (N_7392,N_6202,N_6800);
nand U7393 (N_7393,N_6691,N_6973);
or U7394 (N_7394,N_6930,N_6137);
and U7395 (N_7395,N_6733,N_6015);
and U7396 (N_7396,N_6960,N_6053);
nand U7397 (N_7397,N_6903,N_6786);
and U7398 (N_7398,N_6910,N_6547);
nor U7399 (N_7399,N_6343,N_6392);
or U7400 (N_7400,N_6752,N_6234);
and U7401 (N_7401,N_6026,N_6104);
and U7402 (N_7402,N_6178,N_6065);
or U7403 (N_7403,N_6409,N_6073);
nor U7404 (N_7404,N_6638,N_6523);
or U7405 (N_7405,N_6675,N_6364);
nand U7406 (N_7406,N_6772,N_6946);
nor U7407 (N_7407,N_6716,N_6598);
nand U7408 (N_7408,N_6875,N_6812);
nand U7409 (N_7409,N_6809,N_6671);
xnor U7410 (N_7410,N_6727,N_6363);
or U7411 (N_7411,N_6295,N_6097);
and U7412 (N_7412,N_6922,N_6701);
nand U7413 (N_7413,N_6274,N_6259);
nand U7414 (N_7414,N_6906,N_6464);
nor U7415 (N_7415,N_6870,N_6020);
and U7416 (N_7416,N_6505,N_6720);
and U7417 (N_7417,N_6850,N_6807);
xor U7418 (N_7418,N_6750,N_6166);
or U7419 (N_7419,N_6215,N_6813);
nand U7420 (N_7420,N_6209,N_6669);
and U7421 (N_7421,N_6559,N_6481);
nor U7422 (N_7422,N_6858,N_6354);
or U7423 (N_7423,N_6799,N_6213);
nand U7424 (N_7424,N_6506,N_6581);
or U7425 (N_7425,N_6890,N_6520);
nor U7426 (N_7426,N_6944,N_6293);
and U7427 (N_7427,N_6403,N_6037);
or U7428 (N_7428,N_6022,N_6534);
nor U7429 (N_7429,N_6876,N_6540);
and U7430 (N_7430,N_6466,N_6631);
nor U7431 (N_7431,N_6835,N_6605);
nand U7432 (N_7432,N_6774,N_6052);
nor U7433 (N_7433,N_6418,N_6999);
and U7434 (N_7434,N_6046,N_6438);
nand U7435 (N_7435,N_6007,N_6479);
nand U7436 (N_7436,N_6532,N_6756);
nor U7437 (N_7437,N_6928,N_6655);
and U7438 (N_7438,N_6214,N_6062);
nand U7439 (N_7439,N_6006,N_6785);
nor U7440 (N_7440,N_6367,N_6830);
nand U7441 (N_7441,N_6127,N_6427);
nor U7442 (N_7442,N_6297,N_6880);
and U7443 (N_7443,N_6646,N_6560);
nor U7444 (N_7444,N_6332,N_6853);
or U7445 (N_7445,N_6599,N_6831);
and U7446 (N_7446,N_6522,N_6511);
and U7447 (N_7447,N_6838,N_6686);
or U7448 (N_7448,N_6630,N_6625);
nand U7449 (N_7449,N_6976,N_6162);
or U7450 (N_7450,N_6021,N_6568);
nor U7451 (N_7451,N_6102,N_6986);
or U7452 (N_7452,N_6241,N_6739);
or U7453 (N_7453,N_6074,N_6776);
or U7454 (N_7454,N_6474,N_6371);
or U7455 (N_7455,N_6749,N_6574);
xnor U7456 (N_7456,N_6793,N_6844);
xor U7457 (N_7457,N_6423,N_6376);
and U7458 (N_7458,N_6152,N_6290);
nand U7459 (N_7459,N_6588,N_6923);
and U7460 (N_7460,N_6385,N_6899);
nand U7461 (N_7461,N_6513,N_6755);
nor U7462 (N_7462,N_6902,N_6284);
xnor U7463 (N_7463,N_6670,N_6775);
nand U7464 (N_7464,N_6847,N_6436);
nand U7465 (N_7465,N_6952,N_6269);
or U7466 (N_7466,N_6852,N_6648);
nor U7467 (N_7467,N_6228,N_6114);
and U7468 (N_7468,N_6577,N_6485);
nor U7469 (N_7469,N_6947,N_6470);
and U7470 (N_7470,N_6431,N_6301);
nor U7471 (N_7471,N_6528,N_6917);
xor U7472 (N_7472,N_6744,N_6306);
nor U7473 (N_7473,N_6314,N_6829);
and U7474 (N_7474,N_6996,N_6919);
nand U7475 (N_7475,N_6995,N_6266);
nor U7476 (N_7476,N_6517,N_6682);
nand U7477 (N_7477,N_6008,N_6929);
nand U7478 (N_7478,N_6350,N_6124);
or U7479 (N_7479,N_6468,N_6211);
nand U7480 (N_7480,N_6596,N_6109);
xor U7481 (N_7481,N_6243,N_6649);
nor U7482 (N_7482,N_6687,N_6085);
nand U7483 (N_7483,N_6320,N_6664);
nand U7484 (N_7484,N_6808,N_6951);
or U7485 (N_7485,N_6348,N_6797);
nor U7486 (N_7486,N_6746,N_6378);
or U7487 (N_7487,N_6278,N_6263);
nor U7488 (N_7488,N_6465,N_6879);
xor U7489 (N_7489,N_6897,N_6676);
or U7490 (N_7490,N_6826,N_6095);
or U7491 (N_7491,N_6783,N_6758);
or U7492 (N_7492,N_6536,N_6527);
and U7493 (N_7493,N_6497,N_6594);
nand U7494 (N_7494,N_6966,N_6083);
and U7495 (N_7495,N_6699,N_6282);
nor U7496 (N_7496,N_6163,N_6628);
nand U7497 (N_7497,N_6155,N_6820);
and U7498 (N_7498,N_6541,N_6886);
nor U7499 (N_7499,N_6315,N_6486);
or U7500 (N_7500,N_6367,N_6520);
nand U7501 (N_7501,N_6733,N_6874);
xor U7502 (N_7502,N_6106,N_6692);
or U7503 (N_7503,N_6858,N_6824);
or U7504 (N_7504,N_6217,N_6990);
nand U7505 (N_7505,N_6996,N_6132);
xnor U7506 (N_7506,N_6766,N_6697);
nand U7507 (N_7507,N_6361,N_6449);
and U7508 (N_7508,N_6630,N_6726);
and U7509 (N_7509,N_6172,N_6624);
xor U7510 (N_7510,N_6491,N_6826);
or U7511 (N_7511,N_6308,N_6706);
nor U7512 (N_7512,N_6982,N_6136);
nand U7513 (N_7513,N_6370,N_6634);
or U7514 (N_7514,N_6710,N_6873);
or U7515 (N_7515,N_6086,N_6371);
nand U7516 (N_7516,N_6658,N_6600);
nor U7517 (N_7517,N_6292,N_6539);
or U7518 (N_7518,N_6650,N_6263);
xnor U7519 (N_7519,N_6783,N_6442);
and U7520 (N_7520,N_6549,N_6785);
or U7521 (N_7521,N_6563,N_6534);
nor U7522 (N_7522,N_6621,N_6403);
or U7523 (N_7523,N_6493,N_6550);
or U7524 (N_7524,N_6278,N_6252);
or U7525 (N_7525,N_6613,N_6662);
or U7526 (N_7526,N_6634,N_6970);
nand U7527 (N_7527,N_6602,N_6310);
nand U7528 (N_7528,N_6556,N_6200);
nand U7529 (N_7529,N_6367,N_6611);
or U7530 (N_7530,N_6582,N_6445);
nand U7531 (N_7531,N_6417,N_6407);
xnor U7532 (N_7532,N_6650,N_6712);
or U7533 (N_7533,N_6015,N_6658);
xor U7534 (N_7534,N_6599,N_6972);
nand U7535 (N_7535,N_6622,N_6731);
nor U7536 (N_7536,N_6826,N_6096);
and U7537 (N_7537,N_6645,N_6881);
or U7538 (N_7538,N_6113,N_6529);
xor U7539 (N_7539,N_6856,N_6828);
nor U7540 (N_7540,N_6293,N_6400);
and U7541 (N_7541,N_6816,N_6705);
nor U7542 (N_7542,N_6259,N_6998);
nand U7543 (N_7543,N_6800,N_6186);
nand U7544 (N_7544,N_6669,N_6850);
nand U7545 (N_7545,N_6055,N_6489);
nand U7546 (N_7546,N_6708,N_6020);
and U7547 (N_7547,N_6825,N_6010);
nand U7548 (N_7548,N_6744,N_6942);
and U7549 (N_7549,N_6551,N_6530);
nand U7550 (N_7550,N_6499,N_6689);
nand U7551 (N_7551,N_6028,N_6334);
or U7552 (N_7552,N_6765,N_6770);
nand U7553 (N_7553,N_6299,N_6169);
xor U7554 (N_7554,N_6294,N_6098);
and U7555 (N_7555,N_6757,N_6913);
nor U7556 (N_7556,N_6869,N_6560);
and U7557 (N_7557,N_6588,N_6934);
and U7558 (N_7558,N_6155,N_6324);
nand U7559 (N_7559,N_6753,N_6258);
and U7560 (N_7560,N_6242,N_6847);
nand U7561 (N_7561,N_6834,N_6737);
or U7562 (N_7562,N_6109,N_6025);
and U7563 (N_7563,N_6338,N_6416);
and U7564 (N_7564,N_6982,N_6240);
nor U7565 (N_7565,N_6502,N_6033);
and U7566 (N_7566,N_6051,N_6380);
nand U7567 (N_7567,N_6833,N_6912);
nor U7568 (N_7568,N_6620,N_6851);
and U7569 (N_7569,N_6910,N_6442);
or U7570 (N_7570,N_6075,N_6465);
nand U7571 (N_7571,N_6791,N_6921);
or U7572 (N_7572,N_6690,N_6062);
and U7573 (N_7573,N_6488,N_6555);
or U7574 (N_7574,N_6551,N_6474);
or U7575 (N_7575,N_6155,N_6024);
nor U7576 (N_7576,N_6197,N_6994);
nor U7577 (N_7577,N_6569,N_6789);
or U7578 (N_7578,N_6765,N_6196);
nor U7579 (N_7579,N_6108,N_6120);
nand U7580 (N_7580,N_6023,N_6972);
nand U7581 (N_7581,N_6776,N_6574);
and U7582 (N_7582,N_6383,N_6791);
or U7583 (N_7583,N_6629,N_6981);
nand U7584 (N_7584,N_6592,N_6002);
or U7585 (N_7585,N_6203,N_6512);
nor U7586 (N_7586,N_6142,N_6310);
nor U7587 (N_7587,N_6339,N_6153);
nand U7588 (N_7588,N_6473,N_6186);
and U7589 (N_7589,N_6486,N_6766);
nor U7590 (N_7590,N_6387,N_6290);
nand U7591 (N_7591,N_6627,N_6890);
xor U7592 (N_7592,N_6630,N_6452);
nor U7593 (N_7593,N_6805,N_6989);
nor U7594 (N_7594,N_6698,N_6359);
or U7595 (N_7595,N_6099,N_6510);
or U7596 (N_7596,N_6652,N_6968);
xor U7597 (N_7597,N_6931,N_6925);
and U7598 (N_7598,N_6715,N_6749);
and U7599 (N_7599,N_6460,N_6944);
and U7600 (N_7600,N_6537,N_6912);
nand U7601 (N_7601,N_6939,N_6178);
and U7602 (N_7602,N_6823,N_6369);
and U7603 (N_7603,N_6972,N_6821);
or U7604 (N_7604,N_6407,N_6126);
nand U7605 (N_7605,N_6526,N_6105);
or U7606 (N_7606,N_6214,N_6676);
and U7607 (N_7607,N_6369,N_6492);
and U7608 (N_7608,N_6832,N_6199);
nand U7609 (N_7609,N_6047,N_6672);
and U7610 (N_7610,N_6161,N_6260);
nor U7611 (N_7611,N_6298,N_6337);
and U7612 (N_7612,N_6310,N_6703);
nand U7613 (N_7613,N_6543,N_6362);
nor U7614 (N_7614,N_6988,N_6876);
nor U7615 (N_7615,N_6654,N_6383);
xor U7616 (N_7616,N_6575,N_6216);
and U7617 (N_7617,N_6596,N_6280);
xnor U7618 (N_7618,N_6516,N_6886);
or U7619 (N_7619,N_6937,N_6527);
nor U7620 (N_7620,N_6606,N_6745);
and U7621 (N_7621,N_6134,N_6021);
nand U7622 (N_7622,N_6362,N_6135);
nand U7623 (N_7623,N_6728,N_6490);
nor U7624 (N_7624,N_6473,N_6339);
and U7625 (N_7625,N_6342,N_6380);
nand U7626 (N_7626,N_6584,N_6511);
and U7627 (N_7627,N_6520,N_6108);
or U7628 (N_7628,N_6917,N_6321);
nor U7629 (N_7629,N_6628,N_6406);
and U7630 (N_7630,N_6462,N_6245);
nor U7631 (N_7631,N_6955,N_6634);
and U7632 (N_7632,N_6491,N_6293);
nor U7633 (N_7633,N_6089,N_6776);
or U7634 (N_7634,N_6446,N_6626);
nor U7635 (N_7635,N_6367,N_6915);
and U7636 (N_7636,N_6305,N_6926);
or U7637 (N_7637,N_6202,N_6219);
nor U7638 (N_7638,N_6126,N_6859);
and U7639 (N_7639,N_6192,N_6244);
nor U7640 (N_7640,N_6478,N_6672);
or U7641 (N_7641,N_6234,N_6145);
nor U7642 (N_7642,N_6468,N_6012);
nor U7643 (N_7643,N_6995,N_6288);
or U7644 (N_7644,N_6299,N_6211);
nor U7645 (N_7645,N_6208,N_6660);
nor U7646 (N_7646,N_6214,N_6194);
or U7647 (N_7647,N_6104,N_6474);
nor U7648 (N_7648,N_6304,N_6360);
nand U7649 (N_7649,N_6203,N_6355);
or U7650 (N_7650,N_6033,N_6024);
or U7651 (N_7651,N_6165,N_6404);
xnor U7652 (N_7652,N_6300,N_6184);
nand U7653 (N_7653,N_6551,N_6854);
or U7654 (N_7654,N_6602,N_6751);
nor U7655 (N_7655,N_6461,N_6799);
or U7656 (N_7656,N_6016,N_6997);
or U7657 (N_7657,N_6302,N_6735);
and U7658 (N_7658,N_6990,N_6310);
or U7659 (N_7659,N_6461,N_6277);
xor U7660 (N_7660,N_6447,N_6726);
or U7661 (N_7661,N_6536,N_6042);
nor U7662 (N_7662,N_6838,N_6542);
nand U7663 (N_7663,N_6406,N_6658);
and U7664 (N_7664,N_6006,N_6703);
nor U7665 (N_7665,N_6315,N_6328);
or U7666 (N_7666,N_6599,N_6477);
nand U7667 (N_7667,N_6162,N_6711);
nor U7668 (N_7668,N_6459,N_6436);
nor U7669 (N_7669,N_6512,N_6989);
xor U7670 (N_7670,N_6981,N_6125);
xnor U7671 (N_7671,N_6110,N_6716);
or U7672 (N_7672,N_6379,N_6939);
nor U7673 (N_7673,N_6039,N_6091);
or U7674 (N_7674,N_6194,N_6998);
or U7675 (N_7675,N_6273,N_6932);
and U7676 (N_7676,N_6125,N_6236);
xor U7677 (N_7677,N_6212,N_6041);
or U7678 (N_7678,N_6172,N_6061);
nand U7679 (N_7679,N_6746,N_6181);
or U7680 (N_7680,N_6493,N_6138);
xnor U7681 (N_7681,N_6095,N_6013);
nand U7682 (N_7682,N_6012,N_6531);
nor U7683 (N_7683,N_6168,N_6749);
or U7684 (N_7684,N_6893,N_6206);
or U7685 (N_7685,N_6847,N_6587);
or U7686 (N_7686,N_6517,N_6747);
nor U7687 (N_7687,N_6071,N_6779);
or U7688 (N_7688,N_6912,N_6960);
and U7689 (N_7689,N_6542,N_6855);
nand U7690 (N_7690,N_6438,N_6906);
xor U7691 (N_7691,N_6122,N_6124);
nand U7692 (N_7692,N_6899,N_6062);
xnor U7693 (N_7693,N_6687,N_6582);
nand U7694 (N_7694,N_6495,N_6747);
xnor U7695 (N_7695,N_6496,N_6685);
or U7696 (N_7696,N_6517,N_6446);
nand U7697 (N_7697,N_6483,N_6108);
nor U7698 (N_7698,N_6525,N_6156);
or U7699 (N_7699,N_6493,N_6992);
nor U7700 (N_7700,N_6239,N_6912);
nand U7701 (N_7701,N_6800,N_6668);
or U7702 (N_7702,N_6847,N_6682);
and U7703 (N_7703,N_6449,N_6965);
or U7704 (N_7704,N_6116,N_6911);
nor U7705 (N_7705,N_6384,N_6127);
and U7706 (N_7706,N_6604,N_6694);
nand U7707 (N_7707,N_6620,N_6455);
nand U7708 (N_7708,N_6564,N_6712);
or U7709 (N_7709,N_6418,N_6773);
or U7710 (N_7710,N_6006,N_6327);
nand U7711 (N_7711,N_6678,N_6570);
and U7712 (N_7712,N_6397,N_6101);
nand U7713 (N_7713,N_6251,N_6066);
nand U7714 (N_7714,N_6937,N_6203);
xor U7715 (N_7715,N_6074,N_6360);
nand U7716 (N_7716,N_6698,N_6782);
nor U7717 (N_7717,N_6956,N_6279);
nor U7718 (N_7718,N_6636,N_6260);
nand U7719 (N_7719,N_6573,N_6021);
or U7720 (N_7720,N_6270,N_6373);
nor U7721 (N_7721,N_6611,N_6854);
nor U7722 (N_7722,N_6387,N_6983);
nand U7723 (N_7723,N_6998,N_6240);
nor U7724 (N_7724,N_6560,N_6917);
or U7725 (N_7725,N_6478,N_6179);
nor U7726 (N_7726,N_6869,N_6377);
and U7727 (N_7727,N_6729,N_6756);
nand U7728 (N_7728,N_6452,N_6121);
and U7729 (N_7729,N_6911,N_6577);
and U7730 (N_7730,N_6320,N_6540);
xnor U7731 (N_7731,N_6699,N_6627);
or U7732 (N_7732,N_6307,N_6929);
and U7733 (N_7733,N_6111,N_6604);
nand U7734 (N_7734,N_6534,N_6256);
or U7735 (N_7735,N_6478,N_6316);
nor U7736 (N_7736,N_6875,N_6039);
nor U7737 (N_7737,N_6135,N_6091);
xor U7738 (N_7738,N_6996,N_6368);
and U7739 (N_7739,N_6580,N_6867);
xor U7740 (N_7740,N_6603,N_6531);
nand U7741 (N_7741,N_6104,N_6194);
nand U7742 (N_7742,N_6814,N_6461);
nand U7743 (N_7743,N_6896,N_6109);
nor U7744 (N_7744,N_6009,N_6079);
nand U7745 (N_7745,N_6831,N_6221);
nand U7746 (N_7746,N_6701,N_6395);
and U7747 (N_7747,N_6648,N_6204);
or U7748 (N_7748,N_6319,N_6420);
or U7749 (N_7749,N_6243,N_6346);
nor U7750 (N_7750,N_6399,N_6739);
nand U7751 (N_7751,N_6647,N_6780);
nand U7752 (N_7752,N_6130,N_6700);
nor U7753 (N_7753,N_6803,N_6111);
nor U7754 (N_7754,N_6473,N_6905);
xor U7755 (N_7755,N_6467,N_6594);
nand U7756 (N_7756,N_6388,N_6829);
xor U7757 (N_7757,N_6063,N_6310);
xor U7758 (N_7758,N_6938,N_6890);
nand U7759 (N_7759,N_6578,N_6648);
or U7760 (N_7760,N_6922,N_6336);
and U7761 (N_7761,N_6537,N_6250);
nor U7762 (N_7762,N_6482,N_6382);
nor U7763 (N_7763,N_6173,N_6222);
nor U7764 (N_7764,N_6690,N_6685);
nor U7765 (N_7765,N_6151,N_6209);
nor U7766 (N_7766,N_6263,N_6436);
or U7767 (N_7767,N_6446,N_6197);
nor U7768 (N_7768,N_6335,N_6216);
or U7769 (N_7769,N_6367,N_6182);
nand U7770 (N_7770,N_6540,N_6901);
or U7771 (N_7771,N_6222,N_6823);
nor U7772 (N_7772,N_6443,N_6338);
nand U7773 (N_7773,N_6213,N_6729);
or U7774 (N_7774,N_6692,N_6700);
and U7775 (N_7775,N_6979,N_6237);
or U7776 (N_7776,N_6285,N_6886);
or U7777 (N_7777,N_6746,N_6884);
or U7778 (N_7778,N_6573,N_6603);
nor U7779 (N_7779,N_6426,N_6650);
xnor U7780 (N_7780,N_6708,N_6824);
xnor U7781 (N_7781,N_6527,N_6070);
nand U7782 (N_7782,N_6867,N_6065);
nor U7783 (N_7783,N_6335,N_6270);
or U7784 (N_7784,N_6644,N_6446);
nand U7785 (N_7785,N_6685,N_6644);
and U7786 (N_7786,N_6144,N_6463);
nor U7787 (N_7787,N_6700,N_6190);
nor U7788 (N_7788,N_6042,N_6645);
and U7789 (N_7789,N_6272,N_6088);
nor U7790 (N_7790,N_6942,N_6200);
or U7791 (N_7791,N_6206,N_6823);
or U7792 (N_7792,N_6331,N_6359);
nand U7793 (N_7793,N_6479,N_6400);
nor U7794 (N_7794,N_6578,N_6206);
or U7795 (N_7795,N_6421,N_6083);
nand U7796 (N_7796,N_6209,N_6952);
and U7797 (N_7797,N_6167,N_6053);
and U7798 (N_7798,N_6750,N_6589);
xnor U7799 (N_7799,N_6140,N_6300);
nand U7800 (N_7800,N_6833,N_6463);
xnor U7801 (N_7801,N_6094,N_6421);
nand U7802 (N_7802,N_6724,N_6183);
nand U7803 (N_7803,N_6356,N_6551);
nand U7804 (N_7804,N_6261,N_6211);
xnor U7805 (N_7805,N_6445,N_6242);
nand U7806 (N_7806,N_6951,N_6385);
nand U7807 (N_7807,N_6988,N_6454);
nor U7808 (N_7808,N_6977,N_6648);
xnor U7809 (N_7809,N_6557,N_6488);
xnor U7810 (N_7810,N_6773,N_6892);
nand U7811 (N_7811,N_6932,N_6792);
and U7812 (N_7812,N_6669,N_6974);
and U7813 (N_7813,N_6799,N_6866);
xor U7814 (N_7814,N_6968,N_6345);
nor U7815 (N_7815,N_6667,N_6839);
and U7816 (N_7816,N_6481,N_6333);
and U7817 (N_7817,N_6440,N_6966);
xor U7818 (N_7818,N_6601,N_6610);
xnor U7819 (N_7819,N_6525,N_6776);
and U7820 (N_7820,N_6040,N_6240);
nor U7821 (N_7821,N_6703,N_6672);
xor U7822 (N_7822,N_6714,N_6194);
nor U7823 (N_7823,N_6416,N_6546);
nand U7824 (N_7824,N_6252,N_6349);
nand U7825 (N_7825,N_6723,N_6356);
nand U7826 (N_7826,N_6177,N_6955);
and U7827 (N_7827,N_6940,N_6089);
or U7828 (N_7828,N_6908,N_6295);
or U7829 (N_7829,N_6318,N_6460);
nor U7830 (N_7830,N_6137,N_6799);
and U7831 (N_7831,N_6906,N_6290);
or U7832 (N_7832,N_6177,N_6458);
xor U7833 (N_7833,N_6246,N_6757);
and U7834 (N_7834,N_6743,N_6377);
nor U7835 (N_7835,N_6148,N_6078);
and U7836 (N_7836,N_6814,N_6745);
nand U7837 (N_7837,N_6797,N_6202);
or U7838 (N_7838,N_6845,N_6201);
nand U7839 (N_7839,N_6763,N_6728);
and U7840 (N_7840,N_6473,N_6989);
nand U7841 (N_7841,N_6966,N_6786);
xor U7842 (N_7842,N_6387,N_6263);
and U7843 (N_7843,N_6723,N_6018);
and U7844 (N_7844,N_6108,N_6325);
nor U7845 (N_7845,N_6300,N_6703);
xnor U7846 (N_7846,N_6421,N_6090);
nand U7847 (N_7847,N_6676,N_6545);
or U7848 (N_7848,N_6597,N_6123);
nor U7849 (N_7849,N_6652,N_6553);
nor U7850 (N_7850,N_6926,N_6057);
nand U7851 (N_7851,N_6076,N_6760);
nand U7852 (N_7852,N_6010,N_6804);
nor U7853 (N_7853,N_6915,N_6238);
nor U7854 (N_7854,N_6433,N_6507);
or U7855 (N_7855,N_6502,N_6908);
nor U7856 (N_7856,N_6840,N_6619);
xnor U7857 (N_7857,N_6469,N_6290);
nand U7858 (N_7858,N_6677,N_6670);
or U7859 (N_7859,N_6039,N_6355);
nand U7860 (N_7860,N_6340,N_6994);
nand U7861 (N_7861,N_6537,N_6031);
xor U7862 (N_7862,N_6531,N_6091);
xnor U7863 (N_7863,N_6033,N_6371);
nand U7864 (N_7864,N_6710,N_6585);
or U7865 (N_7865,N_6070,N_6334);
nand U7866 (N_7866,N_6674,N_6002);
or U7867 (N_7867,N_6918,N_6303);
nand U7868 (N_7868,N_6828,N_6042);
and U7869 (N_7869,N_6499,N_6144);
or U7870 (N_7870,N_6956,N_6691);
nand U7871 (N_7871,N_6370,N_6702);
nand U7872 (N_7872,N_6294,N_6573);
and U7873 (N_7873,N_6857,N_6989);
nand U7874 (N_7874,N_6251,N_6498);
nand U7875 (N_7875,N_6212,N_6864);
nor U7876 (N_7876,N_6043,N_6794);
and U7877 (N_7877,N_6808,N_6831);
and U7878 (N_7878,N_6038,N_6248);
or U7879 (N_7879,N_6754,N_6358);
and U7880 (N_7880,N_6070,N_6386);
xor U7881 (N_7881,N_6939,N_6618);
or U7882 (N_7882,N_6173,N_6622);
or U7883 (N_7883,N_6406,N_6247);
and U7884 (N_7884,N_6229,N_6744);
nand U7885 (N_7885,N_6976,N_6870);
nor U7886 (N_7886,N_6314,N_6476);
xnor U7887 (N_7887,N_6742,N_6862);
or U7888 (N_7888,N_6733,N_6488);
or U7889 (N_7889,N_6306,N_6596);
and U7890 (N_7890,N_6549,N_6790);
nor U7891 (N_7891,N_6048,N_6676);
nand U7892 (N_7892,N_6688,N_6304);
and U7893 (N_7893,N_6509,N_6421);
nand U7894 (N_7894,N_6885,N_6606);
nand U7895 (N_7895,N_6935,N_6015);
and U7896 (N_7896,N_6615,N_6284);
nand U7897 (N_7897,N_6793,N_6649);
or U7898 (N_7898,N_6112,N_6810);
or U7899 (N_7899,N_6904,N_6421);
and U7900 (N_7900,N_6221,N_6223);
and U7901 (N_7901,N_6119,N_6891);
nor U7902 (N_7902,N_6618,N_6437);
nand U7903 (N_7903,N_6431,N_6185);
or U7904 (N_7904,N_6395,N_6941);
nor U7905 (N_7905,N_6617,N_6830);
or U7906 (N_7906,N_6550,N_6653);
nor U7907 (N_7907,N_6900,N_6119);
nand U7908 (N_7908,N_6853,N_6620);
xor U7909 (N_7909,N_6537,N_6578);
and U7910 (N_7910,N_6242,N_6383);
or U7911 (N_7911,N_6949,N_6200);
or U7912 (N_7912,N_6935,N_6335);
or U7913 (N_7913,N_6565,N_6184);
or U7914 (N_7914,N_6880,N_6783);
or U7915 (N_7915,N_6653,N_6964);
nor U7916 (N_7916,N_6762,N_6792);
or U7917 (N_7917,N_6918,N_6900);
xor U7918 (N_7918,N_6069,N_6616);
or U7919 (N_7919,N_6491,N_6746);
and U7920 (N_7920,N_6622,N_6427);
or U7921 (N_7921,N_6880,N_6748);
nand U7922 (N_7922,N_6208,N_6440);
xnor U7923 (N_7923,N_6203,N_6457);
nor U7924 (N_7924,N_6232,N_6670);
nand U7925 (N_7925,N_6288,N_6732);
nor U7926 (N_7926,N_6853,N_6298);
or U7927 (N_7927,N_6340,N_6285);
nand U7928 (N_7928,N_6495,N_6128);
nand U7929 (N_7929,N_6177,N_6751);
nor U7930 (N_7930,N_6743,N_6436);
and U7931 (N_7931,N_6290,N_6862);
and U7932 (N_7932,N_6364,N_6963);
nand U7933 (N_7933,N_6218,N_6919);
or U7934 (N_7934,N_6521,N_6011);
nand U7935 (N_7935,N_6085,N_6357);
and U7936 (N_7936,N_6424,N_6945);
or U7937 (N_7937,N_6368,N_6462);
and U7938 (N_7938,N_6421,N_6107);
nor U7939 (N_7939,N_6688,N_6841);
nor U7940 (N_7940,N_6747,N_6833);
and U7941 (N_7941,N_6680,N_6821);
nand U7942 (N_7942,N_6369,N_6799);
nand U7943 (N_7943,N_6911,N_6872);
xor U7944 (N_7944,N_6039,N_6642);
nand U7945 (N_7945,N_6608,N_6162);
or U7946 (N_7946,N_6398,N_6280);
and U7947 (N_7947,N_6315,N_6262);
nand U7948 (N_7948,N_6157,N_6530);
xor U7949 (N_7949,N_6613,N_6113);
nor U7950 (N_7950,N_6597,N_6413);
nor U7951 (N_7951,N_6422,N_6342);
nand U7952 (N_7952,N_6444,N_6913);
nor U7953 (N_7953,N_6612,N_6088);
nand U7954 (N_7954,N_6626,N_6833);
xor U7955 (N_7955,N_6895,N_6230);
nand U7956 (N_7956,N_6828,N_6461);
or U7957 (N_7957,N_6056,N_6785);
nor U7958 (N_7958,N_6666,N_6437);
nand U7959 (N_7959,N_6749,N_6385);
or U7960 (N_7960,N_6719,N_6332);
nor U7961 (N_7961,N_6490,N_6164);
nor U7962 (N_7962,N_6827,N_6769);
or U7963 (N_7963,N_6325,N_6027);
or U7964 (N_7964,N_6626,N_6592);
xnor U7965 (N_7965,N_6815,N_6231);
nand U7966 (N_7966,N_6615,N_6399);
nor U7967 (N_7967,N_6383,N_6238);
and U7968 (N_7968,N_6748,N_6030);
nand U7969 (N_7969,N_6263,N_6154);
nor U7970 (N_7970,N_6264,N_6796);
and U7971 (N_7971,N_6493,N_6228);
and U7972 (N_7972,N_6498,N_6468);
xor U7973 (N_7973,N_6277,N_6644);
nor U7974 (N_7974,N_6441,N_6057);
nor U7975 (N_7975,N_6483,N_6331);
or U7976 (N_7976,N_6131,N_6782);
nor U7977 (N_7977,N_6538,N_6856);
nand U7978 (N_7978,N_6897,N_6462);
xor U7979 (N_7979,N_6907,N_6295);
nor U7980 (N_7980,N_6070,N_6685);
or U7981 (N_7981,N_6923,N_6482);
nand U7982 (N_7982,N_6138,N_6268);
nand U7983 (N_7983,N_6554,N_6493);
nand U7984 (N_7984,N_6074,N_6698);
nand U7985 (N_7985,N_6708,N_6838);
xor U7986 (N_7986,N_6932,N_6779);
or U7987 (N_7987,N_6583,N_6020);
nand U7988 (N_7988,N_6705,N_6086);
nor U7989 (N_7989,N_6768,N_6973);
and U7990 (N_7990,N_6892,N_6089);
and U7991 (N_7991,N_6374,N_6179);
or U7992 (N_7992,N_6653,N_6955);
nand U7993 (N_7993,N_6274,N_6062);
or U7994 (N_7994,N_6673,N_6416);
or U7995 (N_7995,N_6317,N_6759);
or U7996 (N_7996,N_6277,N_6586);
xor U7997 (N_7997,N_6185,N_6944);
and U7998 (N_7998,N_6576,N_6063);
or U7999 (N_7999,N_6825,N_6680);
or U8000 (N_8000,N_7002,N_7430);
or U8001 (N_8001,N_7428,N_7336);
nand U8002 (N_8002,N_7383,N_7672);
nor U8003 (N_8003,N_7206,N_7947);
and U8004 (N_8004,N_7082,N_7326);
nor U8005 (N_8005,N_7315,N_7378);
and U8006 (N_8006,N_7354,N_7496);
and U8007 (N_8007,N_7524,N_7346);
nor U8008 (N_8008,N_7615,N_7787);
or U8009 (N_8009,N_7872,N_7299);
nand U8010 (N_8010,N_7003,N_7902);
and U8011 (N_8011,N_7553,N_7480);
or U8012 (N_8012,N_7358,N_7011);
nand U8013 (N_8013,N_7238,N_7666);
nor U8014 (N_8014,N_7382,N_7142);
xor U8015 (N_8015,N_7706,N_7085);
nand U8016 (N_8016,N_7412,N_7145);
nand U8017 (N_8017,N_7647,N_7867);
and U8018 (N_8018,N_7138,N_7931);
xnor U8019 (N_8019,N_7546,N_7053);
and U8020 (N_8020,N_7267,N_7555);
or U8021 (N_8021,N_7297,N_7864);
nor U8022 (N_8022,N_7376,N_7283);
nand U8023 (N_8023,N_7017,N_7848);
nor U8024 (N_8024,N_7102,N_7986);
nor U8025 (N_8025,N_7477,N_7934);
and U8026 (N_8026,N_7581,N_7605);
and U8027 (N_8027,N_7276,N_7628);
and U8028 (N_8028,N_7134,N_7410);
nand U8029 (N_8029,N_7368,N_7190);
nand U8030 (N_8030,N_7195,N_7865);
or U8031 (N_8031,N_7869,N_7791);
nand U8032 (N_8032,N_7655,N_7767);
nor U8033 (N_8033,N_7361,N_7303);
or U8034 (N_8034,N_7558,N_7693);
and U8035 (N_8035,N_7669,N_7226);
or U8036 (N_8036,N_7468,N_7527);
or U8037 (N_8037,N_7464,N_7112);
nor U8038 (N_8038,N_7419,N_7060);
nand U8039 (N_8039,N_7568,N_7294);
and U8040 (N_8040,N_7402,N_7813);
nor U8041 (N_8041,N_7632,N_7078);
or U8042 (N_8042,N_7900,N_7945);
nand U8043 (N_8043,N_7789,N_7652);
nor U8044 (N_8044,N_7933,N_7242);
or U8045 (N_8045,N_7857,N_7333);
or U8046 (N_8046,N_7440,N_7013);
and U8047 (N_8047,N_7456,N_7224);
nor U8048 (N_8048,N_7596,N_7510);
and U8049 (N_8049,N_7978,N_7021);
nand U8050 (N_8050,N_7778,N_7665);
nand U8051 (N_8051,N_7471,N_7979);
nor U8052 (N_8052,N_7274,N_7717);
and U8053 (N_8053,N_7390,N_7746);
xnor U8054 (N_8054,N_7006,N_7595);
and U8055 (N_8055,N_7451,N_7272);
nor U8056 (N_8056,N_7100,N_7816);
or U8057 (N_8057,N_7751,N_7146);
or U8058 (N_8058,N_7071,N_7159);
nand U8059 (N_8059,N_7579,N_7712);
or U8060 (N_8060,N_7830,N_7926);
or U8061 (N_8061,N_7629,N_7962);
nor U8062 (N_8062,N_7898,N_7690);
and U8063 (N_8063,N_7735,N_7413);
nor U8064 (N_8064,N_7443,N_7330);
nand U8065 (N_8065,N_7047,N_7876);
nand U8066 (N_8066,N_7044,N_7981);
nor U8067 (N_8067,N_7329,N_7453);
and U8068 (N_8068,N_7485,N_7526);
nor U8069 (N_8069,N_7936,N_7797);
and U8070 (N_8070,N_7842,N_7705);
nor U8071 (N_8071,N_7608,N_7269);
or U8072 (N_8072,N_7783,N_7509);
or U8073 (N_8073,N_7163,N_7247);
nand U8074 (N_8074,N_7135,N_7536);
nand U8075 (N_8075,N_7744,N_7481);
nand U8076 (N_8076,N_7221,N_7715);
and U8077 (N_8077,N_7548,N_7104);
nor U8078 (N_8078,N_7685,N_7811);
or U8079 (N_8079,N_7088,N_7364);
nor U8080 (N_8080,N_7461,N_7020);
nand U8081 (N_8081,N_7441,N_7356);
nor U8082 (N_8082,N_7278,N_7680);
nor U8083 (N_8083,N_7710,N_7923);
or U8084 (N_8084,N_7399,N_7331);
nand U8085 (N_8085,N_7182,N_7338);
nand U8086 (N_8086,N_7850,N_7856);
nor U8087 (N_8087,N_7774,N_7539);
and U8088 (N_8088,N_7362,N_7858);
or U8089 (N_8089,N_7367,N_7832);
or U8090 (N_8090,N_7503,N_7821);
or U8091 (N_8091,N_7156,N_7051);
nand U8092 (N_8092,N_7109,N_7826);
xor U8093 (N_8093,N_7279,N_7282);
nand U8094 (N_8094,N_7834,N_7016);
and U8095 (N_8095,N_7965,N_7952);
and U8096 (N_8096,N_7585,N_7349);
nor U8097 (N_8097,N_7042,N_7469);
nor U8098 (N_8098,N_7688,N_7630);
nor U8099 (N_8099,N_7252,N_7943);
nor U8100 (N_8100,N_7730,N_7955);
and U8101 (N_8101,N_7454,N_7411);
or U8102 (N_8102,N_7160,N_7270);
or U8103 (N_8103,N_7366,N_7466);
and U8104 (N_8104,N_7802,N_7048);
nand U8105 (N_8105,N_7124,N_7930);
and U8106 (N_8106,N_7779,N_7415);
and U8107 (N_8107,N_7301,N_7853);
or U8108 (N_8108,N_7452,N_7970);
xor U8109 (N_8109,N_7196,N_7552);
nor U8110 (N_8110,N_7960,N_7638);
and U8111 (N_8111,N_7186,N_7766);
nor U8112 (N_8112,N_7689,N_7198);
and U8113 (N_8113,N_7995,N_7959);
or U8114 (N_8114,N_7521,N_7069);
and U8115 (N_8115,N_7884,N_7506);
xnor U8116 (N_8116,N_7716,N_7760);
xnor U8117 (N_8117,N_7870,N_7839);
and U8118 (N_8118,N_7397,N_7677);
or U8119 (N_8119,N_7285,N_7447);
or U8120 (N_8120,N_7566,N_7380);
and U8121 (N_8121,N_7064,N_7009);
or U8122 (N_8122,N_7950,N_7866);
or U8123 (N_8123,N_7128,N_7609);
or U8124 (N_8124,N_7165,N_7067);
nor U8125 (N_8125,N_7562,N_7704);
nand U8126 (N_8126,N_7401,N_7005);
nor U8127 (N_8127,N_7572,N_7334);
and U8128 (N_8128,N_7360,N_7784);
xor U8129 (N_8129,N_7062,N_7000);
xor U8130 (N_8130,N_7851,N_7775);
or U8131 (N_8131,N_7050,N_7416);
or U8132 (N_8132,N_7115,N_7907);
and U8133 (N_8133,N_7248,N_7117);
and U8134 (N_8134,N_7939,N_7614);
or U8135 (N_8135,N_7586,N_7927);
and U8136 (N_8136,N_7417,N_7066);
and U8137 (N_8137,N_7687,N_7529);
nor U8138 (N_8138,N_7008,N_7482);
xnor U8139 (N_8139,N_7097,N_7332);
nor U8140 (N_8140,N_7559,N_7737);
or U8141 (N_8141,N_7321,N_7984);
or U8142 (N_8142,N_7734,N_7444);
or U8143 (N_8143,N_7395,N_7582);
or U8144 (N_8144,N_7880,N_7697);
and U8145 (N_8145,N_7547,N_7946);
or U8146 (N_8146,N_7545,N_7998);
nor U8147 (N_8147,N_7473,N_7941);
nor U8148 (N_8148,N_7486,N_7768);
or U8149 (N_8149,N_7091,N_7560);
nor U8150 (N_8150,N_7932,N_7845);
nand U8151 (N_8151,N_7694,N_7924);
nand U8152 (N_8152,N_7110,N_7670);
nand U8153 (N_8153,N_7445,N_7203);
nand U8154 (N_8154,N_7280,N_7184);
nand U8155 (N_8155,N_7126,N_7040);
xnor U8156 (N_8156,N_7286,N_7805);
nand U8157 (N_8157,N_7393,N_7339);
xor U8158 (N_8158,N_7713,N_7750);
nand U8159 (N_8159,N_7291,N_7218);
nand U8160 (N_8160,N_7571,N_7999);
xnor U8161 (N_8161,N_7041,N_7432);
and U8162 (N_8162,N_7249,N_7024);
nor U8163 (N_8163,N_7649,N_7076);
nor U8164 (N_8164,N_7389,N_7187);
nor U8165 (N_8165,N_7639,N_7894);
or U8166 (N_8166,N_7405,N_7036);
nand U8167 (N_8167,N_7534,N_7216);
and U8168 (N_8168,N_7426,N_7251);
and U8169 (N_8169,N_7167,N_7373);
nand U8170 (N_8170,N_7106,N_7273);
nor U8171 (N_8171,N_7037,N_7304);
nand U8172 (N_8172,N_7600,N_7137);
or U8173 (N_8173,N_7659,N_7788);
nor U8174 (N_8174,N_7904,N_7147);
or U8175 (N_8175,N_7173,N_7231);
nor U8176 (N_8176,N_7343,N_7501);
nand U8177 (N_8177,N_7818,N_7055);
xnor U8178 (N_8178,N_7194,N_7681);
nand U8179 (N_8179,N_7487,N_7084);
and U8180 (N_8180,N_7772,N_7829);
nand U8181 (N_8181,N_7578,N_7613);
nand U8182 (N_8182,N_7640,N_7513);
nor U8183 (N_8183,N_7022,N_7575);
xor U8184 (N_8184,N_7499,N_7027);
or U8185 (N_8185,N_7531,N_7045);
nor U8186 (N_8186,N_7949,N_7957);
xor U8187 (N_8187,N_7814,N_7136);
nand U8188 (N_8188,N_7287,N_7785);
nor U8189 (N_8189,N_7653,N_7488);
or U8190 (N_8190,N_7427,N_7989);
nand U8191 (N_8191,N_7754,N_7392);
and U8192 (N_8192,N_7831,N_7265);
nor U8193 (N_8193,N_7741,N_7234);
nand U8194 (N_8194,N_7458,N_7718);
xnor U8195 (N_8195,N_7337,N_7479);
or U8196 (N_8196,N_7262,N_7854);
and U8197 (N_8197,N_7861,N_7974);
xnor U8198 (N_8198,N_7782,N_7807);
or U8199 (N_8199,N_7958,N_7642);
or U8200 (N_8200,N_7835,N_7667);
or U8201 (N_8201,N_7701,N_7964);
and U8202 (N_8202,N_7985,N_7919);
nand U8203 (N_8203,N_7654,N_7598);
nor U8204 (N_8204,N_7912,N_7306);
nand U8205 (N_8205,N_7646,N_7460);
or U8206 (N_8206,N_7874,N_7824);
xnor U8207 (N_8207,N_7201,N_7075);
and U8208 (N_8208,N_7792,N_7462);
or U8209 (N_8209,N_7877,N_7664);
nor U8210 (N_8210,N_7859,N_7241);
xor U8211 (N_8211,N_7292,N_7293);
or U8212 (N_8212,N_7181,N_7624);
nand U8213 (N_8213,N_7275,N_7594);
xnor U8214 (N_8214,N_7174,N_7743);
nand U8215 (N_8215,N_7920,N_7183);
and U8216 (N_8216,N_7557,N_7729);
nor U8217 (N_8217,N_7388,N_7423);
and U8218 (N_8218,N_7179,N_7250);
nor U8219 (N_8219,N_7498,N_7891);
or U8220 (N_8220,N_7141,N_7374);
and U8221 (N_8221,N_7971,N_7796);
or U8222 (N_8222,N_7915,N_7726);
nand U8223 (N_8223,N_7656,N_7537);
or U8224 (N_8224,N_7246,N_7108);
nand U8225 (N_8225,N_7302,N_7465);
or U8226 (N_8226,N_7255,N_7863);
nor U8227 (N_8227,N_7208,N_7031);
nand U8228 (N_8228,N_7103,N_7722);
and U8229 (N_8229,N_7172,N_7387);
xnor U8230 (N_8230,N_7755,N_7626);
nand U8231 (N_8231,N_7612,N_7164);
or U8232 (N_8232,N_7966,N_7121);
nor U8233 (N_8233,N_7438,N_7313);
or U8234 (N_8234,N_7721,N_7414);
nor U8235 (N_8235,N_7833,N_7035);
and U8236 (N_8236,N_7090,N_7308);
xnor U8237 (N_8237,N_7494,N_7489);
and U8238 (N_8238,N_7209,N_7901);
nor U8239 (N_8239,N_7963,N_7341);
and U8240 (N_8240,N_7328,N_7455);
or U8241 (N_8241,N_7969,N_7938);
xor U8242 (N_8242,N_7404,N_7311);
nor U8243 (N_8243,N_7776,N_7113);
nand U8244 (N_8244,N_7061,N_7810);
nor U8245 (N_8245,N_7873,N_7025);
and U8246 (N_8246,N_7254,N_7673);
or U8247 (N_8247,N_7610,N_7457);
or U8248 (N_8248,N_7353,N_7243);
or U8249 (N_8249,N_7809,N_7663);
nand U8250 (N_8250,N_7335,N_7991);
nor U8251 (N_8251,N_7799,N_7497);
or U8252 (N_8252,N_7493,N_7806);
nor U8253 (N_8253,N_7258,N_7837);
nand U8254 (N_8254,N_7679,N_7063);
xor U8255 (N_8255,N_7227,N_7222);
xnor U8256 (N_8256,N_7709,N_7769);
and U8257 (N_8257,N_7570,N_7099);
xor U8258 (N_8258,N_7377,N_7152);
nor U8259 (N_8259,N_7972,N_7028);
and U8260 (N_8260,N_7565,N_7692);
nand U8261 (N_8261,N_7018,N_7519);
and U8262 (N_8262,N_7200,N_7153);
or U8263 (N_8263,N_7645,N_7483);
nand U8264 (N_8264,N_7073,N_7033);
nor U8265 (N_8265,N_7616,N_7199);
or U8266 (N_8266,N_7317,N_7120);
nand U8267 (N_8267,N_7010,N_7551);
xnor U8268 (N_8268,N_7259,N_7043);
nor U8269 (N_8269,N_7508,N_7937);
nor U8270 (N_8270,N_7727,N_7340);
and U8271 (N_8271,N_7838,N_7177);
and U8272 (N_8272,N_7815,N_7324);
nand U8273 (N_8273,N_7648,N_7214);
nand U8274 (N_8274,N_7323,N_7993);
nor U8275 (N_8275,N_7211,N_7910);
or U8276 (N_8276,N_7881,N_7220);
xnor U8277 (N_8277,N_7635,N_7736);
and U8278 (N_8278,N_7589,N_7463);
nor U8279 (N_8279,N_7144,N_7698);
and U8280 (N_8280,N_7849,N_7587);
and U8281 (N_8281,N_7636,N_7956);
or U8282 (N_8282,N_7997,N_7193);
nand U8283 (N_8283,N_7450,N_7913);
nor U8284 (N_8284,N_7723,N_7217);
or U8285 (N_8285,N_7948,N_7935);
or U8286 (N_8286,N_7072,N_7264);
nor U8287 (N_8287,N_7418,N_7525);
nand U8288 (N_8288,N_7188,N_7892);
nand U8289 (N_8289,N_7298,N_7054);
nand U8290 (N_8290,N_7475,N_7569);
or U8291 (N_8291,N_7987,N_7512);
xor U8292 (N_8292,N_7944,N_7786);
nor U8293 (N_8293,N_7800,N_7232);
and U8294 (N_8294,N_7749,N_7794);
or U8295 (N_8295,N_7549,N_7351);
nand U8296 (N_8296,N_7001,N_7140);
xnor U8297 (N_8297,N_7961,N_7550);
nor U8298 (N_8298,N_7803,N_7777);
nand U8299 (N_8299,N_7492,N_7355);
xnor U8300 (N_8300,N_7111,N_7149);
nand U8301 (N_8301,N_7756,N_7975);
xnor U8302 (N_8302,N_7307,N_7202);
and U8303 (N_8303,N_7762,N_7580);
or U8304 (N_8304,N_7192,N_7822);
or U8305 (N_8305,N_7682,N_7049);
nand U8306 (N_8306,N_7675,N_7977);
nor U8307 (N_8307,N_7256,N_7300);
nand U8308 (N_8308,N_7052,N_7089);
or U8309 (N_8309,N_7420,N_7281);
and U8310 (N_8310,N_7742,N_7660);
xnor U8311 (N_8311,N_7459,N_7083);
and U8312 (N_8312,N_7683,N_7883);
nor U8313 (N_8313,N_7719,N_7684);
nor U8314 (N_8314,N_7584,N_7678);
nor U8315 (N_8315,N_7094,N_7540);
nand U8316 (N_8316,N_7239,N_7442);
or U8317 (N_8317,N_7180,N_7812);
nand U8318 (N_8318,N_7421,N_7080);
and U8319 (N_8319,N_7846,N_7808);
nor U8320 (N_8320,N_7436,N_7268);
or U8321 (N_8321,N_7700,N_7823);
or U8322 (N_8322,N_7385,N_7210);
nand U8323 (N_8323,N_7070,N_7650);
nand U8324 (N_8324,N_7516,N_7906);
and U8325 (N_8325,N_7403,N_7068);
and U8326 (N_8326,N_7511,N_7236);
and U8327 (N_8327,N_7394,N_7437);
or U8328 (N_8328,N_7862,N_7905);
nand U8329 (N_8329,N_7176,N_7535);
or U8330 (N_8330,N_7474,N_7056);
or U8331 (N_8331,N_7745,N_7407);
or U8332 (N_8332,N_7542,N_7564);
nand U8333 (N_8333,N_7148,N_7058);
and U8334 (N_8334,N_7922,N_7714);
nor U8335 (N_8335,N_7765,N_7903);
and U8336 (N_8336,N_7739,N_7888);
nand U8337 (N_8337,N_7738,N_7490);
nand U8338 (N_8338,N_7899,N_7583);
and U8339 (N_8339,N_7561,N_7325);
and U8340 (N_8340,N_7625,N_7439);
xor U8341 (N_8341,N_7034,N_7429);
or U8342 (N_8342,N_7357,N_7606);
or U8343 (N_8343,N_7185,N_7651);
and U8344 (N_8344,N_7166,N_7836);
xnor U8345 (N_8345,N_7101,N_7914);
xor U8346 (N_8346,N_7607,N_7724);
xnor U8347 (N_8347,N_7538,N_7168);
and U8348 (N_8348,N_7593,N_7424);
and U8349 (N_8349,N_7092,N_7266);
nand U8350 (N_8350,N_7207,N_7391);
or U8351 (N_8351,N_7189,N_7590);
or U8352 (N_8352,N_7597,N_7178);
and U8353 (N_8353,N_7350,N_7522);
nand U8354 (N_8354,N_7171,N_7662);
or U8355 (N_8355,N_7476,N_7175);
nand U8356 (N_8356,N_7686,N_7691);
xor U8357 (N_8357,N_7817,N_7046);
or U8358 (N_8358,N_7918,N_7668);
nor U8359 (N_8359,N_7305,N_7940);
nand U8360 (N_8360,N_7795,N_7757);
nand U8361 (N_8361,N_7515,N_7344);
nand U8362 (N_8362,N_7720,N_7699);
and U8363 (N_8363,N_7643,N_7284);
xor U8364 (N_8364,N_7801,N_7711);
and U8365 (N_8365,N_7495,N_7014);
nor U8366 (N_8366,N_7409,N_7079);
or U8367 (N_8367,N_7644,N_7820);
or U8368 (N_8368,N_7911,N_7310);
xor U8369 (N_8369,N_7491,N_7191);
nor U8370 (N_8370,N_7620,N_7225);
nor U8371 (N_8371,N_7369,N_7573);
or U8372 (N_8372,N_7170,N_7348);
and U8373 (N_8373,N_7212,N_7763);
nand U8374 (N_8374,N_7633,N_7871);
or U8375 (N_8375,N_7223,N_7819);
xor U8376 (N_8376,N_7983,N_7219);
nand U8377 (N_8377,N_7517,N_7770);
nor U8378 (N_8378,N_7780,N_7370);
and U8379 (N_8379,N_7235,N_7885);
nor U8380 (N_8380,N_7502,N_7953);
nand U8381 (N_8381,N_7290,N_7520);
or U8382 (N_8382,N_7707,N_7747);
nor U8383 (N_8383,N_7532,N_7556);
or U8384 (N_8384,N_7038,N_7233);
nand U8385 (N_8385,N_7731,N_7518);
nor U8386 (N_8386,N_7728,N_7257);
nor U8387 (N_8387,N_7245,N_7618);
nand U8388 (N_8388,N_7197,N_7982);
or U8389 (N_8389,N_7887,N_7263);
or U8390 (N_8390,N_7352,N_7295);
and U8391 (N_8391,N_7237,N_7827);
nor U8392 (N_8392,N_7980,N_7996);
and U8393 (N_8393,N_7574,N_7130);
nor U8394 (N_8394,N_7764,N_7319);
nor U8395 (N_8395,N_7260,N_7314);
nand U8396 (N_8396,N_7081,N_7695);
nor U8397 (N_8397,N_7143,N_7320);
and U8398 (N_8398,N_7446,N_7123);
or U8399 (N_8399,N_7929,N_7781);
or U8400 (N_8400,N_7122,N_7541);
nand U8401 (N_8401,N_7386,N_7087);
nand U8402 (N_8402,N_7322,N_7004);
or U8403 (N_8403,N_7868,N_7886);
and U8404 (N_8404,N_7732,N_7967);
nand U8405 (N_8405,N_7793,N_7057);
or U8406 (N_8406,N_7213,N_7204);
or U8407 (N_8407,N_7576,N_7327);
or U8408 (N_8408,N_7703,N_7507);
or U8409 (N_8409,N_7215,N_7758);
and U8410 (N_8410,N_7676,N_7096);
nand U8411 (N_8411,N_7855,N_7592);
nand U8412 (N_8412,N_7434,N_7032);
or U8413 (N_8413,N_7470,N_7059);
nand U8414 (N_8414,N_7844,N_7131);
or U8415 (N_8415,N_7371,N_7702);
nor U8416 (N_8416,N_7895,N_7288);
nand U8417 (N_8417,N_7875,N_7925);
and U8418 (N_8418,N_7604,N_7406);
nand U8419 (N_8419,N_7928,N_7312);
xnor U8420 (N_8420,N_7882,N_7132);
or U8421 (N_8421,N_7748,N_7157);
nand U8422 (N_8422,N_7161,N_7840);
or U8423 (N_8423,N_7318,N_7954);
and U8424 (N_8424,N_7425,N_7105);
or U8425 (N_8425,N_7261,N_7631);
and U8426 (N_8426,N_7804,N_7271);
nor U8427 (N_8427,N_7841,N_7878);
nand U8428 (N_8428,N_7976,N_7316);
nor U8429 (N_8429,N_7740,N_7151);
nor U8430 (N_8430,N_7229,N_7449);
nand U8431 (N_8431,N_7623,N_7658);
nor U8432 (N_8432,N_7277,N_7500);
nor U8433 (N_8433,N_7637,N_7289);
nor U8434 (N_8434,N_7155,N_7375);
and U8435 (N_8435,N_7563,N_7591);
nand U8436 (N_8436,N_7077,N_7621);
nand U8437 (N_8437,N_7478,N_7909);
nor U8438 (N_8438,N_7893,N_7567);
or U8439 (N_8439,N_7847,N_7617);
nand U8440 (N_8440,N_7150,N_7448);
nand U8441 (N_8441,N_7012,N_7916);
or U8442 (N_8442,N_7896,N_7641);
or U8443 (N_8443,N_7828,N_7879);
or U8444 (N_8444,N_7661,N_7384);
and U8445 (N_8445,N_7696,N_7771);
nor U8446 (N_8446,N_7169,N_7852);
nor U8447 (N_8447,N_7244,N_7725);
or U8448 (N_8448,N_7602,N_7107);
nor U8449 (N_8449,N_7116,N_7381);
or U8450 (N_8450,N_7365,N_7359);
nor U8451 (N_8451,N_7504,N_7026);
and U8452 (N_8452,N_7733,N_7372);
or U8453 (N_8453,N_7530,N_7431);
nand U8454 (N_8454,N_7992,N_7523);
nand U8455 (N_8455,N_7619,N_7422);
xor U8456 (N_8456,N_7860,N_7065);
nand U8457 (N_8457,N_7118,N_7023);
nand U8458 (N_8458,N_7634,N_7467);
and U8459 (N_8459,N_7484,N_7345);
xnor U8460 (N_8460,N_7007,N_7086);
xor U8461 (N_8461,N_7753,N_7139);
and U8462 (N_8462,N_7889,N_7990);
xnor U8463 (N_8463,N_7029,N_7942);
nor U8464 (N_8464,N_7611,N_7129);
nor U8465 (N_8465,N_7752,N_7433);
nor U8466 (N_8466,N_7230,N_7622);
or U8467 (N_8467,N_7074,N_7396);
nand U8468 (N_8468,N_7921,N_7154);
nand U8469 (N_8469,N_7347,N_7988);
and U8470 (N_8470,N_7761,N_7627);
nand U8471 (N_8471,N_7554,N_7095);
or U8472 (N_8472,N_7588,N_7528);
nand U8473 (N_8473,N_7015,N_7162);
nor U8474 (N_8474,N_7127,N_7125);
nor U8475 (N_8475,N_7897,N_7408);
nand U8476 (N_8476,N_7514,N_7240);
nor U8477 (N_8477,N_7603,N_7657);
and U8478 (N_8478,N_7790,N_7533);
nand U8479 (N_8479,N_7544,N_7030);
or U8480 (N_8480,N_7601,N_7968);
nand U8481 (N_8481,N_7133,N_7098);
or U8482 (N_8482,N_7908,N_7674);
or U8483 (N_8483,N_7472,N_7773);
xor U8484 (N_8484,N_7119,N_7093);
and U8485 (N_8485,N_7253,N_7342);
nand U8486 (N_8486,N_7825,N_7039);
nand U8487 (N_8487,N_7363,N_7114);
xor U8488 (N_8488,N_7973,N_7843);
or U8489 (N_8489,N_7708,N_7398);
nor U8490 (N_8490,N_7759,N_7379);
and U8491 (N_8491,N_7309,N_7543);
or U8492 (N_8492,N_7890,N_7599);
nand U8493 (N_8493,N_7951,N_7228);
and U8494 (N_8494,N_7505,N_7400);
nand U8495 (N_8495,N_7435,N_7671);
or U8496 (N_8496,N_7577,N_7798);
or U8497 (N_8497,N_7296,N_7019);
and U8498 (N_8498,N_7994,N_7205);
xor U8499 (N_8499,N_7917,N_7158);
or U8500 (N_8500,N_7759,N_7597);
xnor U8501 (N_8501,N_7135,N_7511);
nor U8502 (N_8502,N_7597,N_7732);
and U8503 (N_8503,N_7188,N_7450);
or U8504 (N_8504,N_7594,N_7903);
nor U8505 (N_8505,N_7086,N_7990);
or U8506 (N_8506,N_7176,N_7891);
nand U8507 (N_8507,N_7147,N_7958);
and U8508 (N_8508,N_7266,N_7604);
nor U8509 (N_8509,N_7808,N_7791);
or U8510 (N_8510,N_7641,N_7449);
nand U8511 (N_8511,N_7080,N_7596);
nand U8512 (N_8512,N_7078,N_7841);
nor U8513 (N_8513,N_7116,N_7255);
and U8514 (N_8514,N_7799,N_7136);
nor U8515 (N_8515,N_7221,N_7430);
nand U8516 (N_8516,N_7411,N_7100);
nor U8517 (N_8517,N_7342,N_7002);
nand U8518 (N_8518,N_7066,N_7729);
nor U8519 (N_8519,N_7170,N_7793);
nand U8520 (N_8520,N_7144,N_7255);
nor U8521 (N_8521,N_7829,N_7095);
or U8522 (N_8522,N_7048,N_7069);
and U8523 (N_8523,N_7322,N_7635);
or U8524 (N_8524,N_7323,N_7678);
and U8525 (N_8525,N_7025,N_7222);
and U8526 (N_8526,N_7049,N_7578);
and U8527 (N_8527,N_7249,N_7848);
nor U8528 (N_8528,N_7006,N_7900);
or U8529 (N_8529,N_7249,N_7211);
and U8530 (N_8530,N_7303,N_7318);
or U8531 (N_8531,N_7519,N_7152);
or U8532 (N_8532,N_7931,N_7563);
and U8533 (N_8533,N_7685,N_7092);
or U8534 (N_8534,N_7403,N_7578);
or U8535 (N_8535,N_7108,N_7981);
nor U8536 (N_8536,N_7286,N_7997);
and U8537 (N_8537,N_7903,N_7784);
nand U8538 (N_8538,N_7477,N_7166);
and U8539 (N_8539,N_7677,N_7042);
nor U8540 (N_8540,N_7208,N_7601);
or U8541 (N_8541,N_7583,N_7754);
or U8542 (N_8542,N_7570,N_7659);
or U8543 (N_8543,N_7376,N_7752);
or U8544 (N_8544,N_7524,N_7981);
or U8545 (N_8545,N_7300,N_7780);
xor U8546 (N_8546,N_7592,N_7959);
nand U8547 (N_8547,N_7110,N_7153);
and U8548 (N_8548,N_7900,N_7277);
and U8549 (N_8549,N_7892,N_7363);
nor U8550 (N_8550,N_7874,N_7991);
nand U8551 (N_8551,N_7292,N_7239);
or U8552 (N_8552,N_7885,N_7895);
nor U8553 (N_8553,N_7959,N_7248);
and U8554 (N_8554,N_7897,N_7069);
and U8555 (N_8555,N_7749,N_7095);
nor U8556 (N_8556,N_7486,N_7520);
and U8557 (N_8557,N_7594,N_7480);
or U8558 (N_8558,N_7726,N_7821);
nor U8559 (N_8559,N_7971,N_7028);
and U8560 (N_8560,N_7767,N_7009);
nand U8561 (N_8561,N_7838,N_7720);
nor U8562 (N_8562,N_7201,N_7270);
nand U8563 (N_8563,N_7808,N_7289);
or U8564 (N_8564,N_7004,N_7921);
xnor U8565 (N_8565,N_7286,N_7792);
xor U8566 (N_8566,N_7814,N_7906);
or U8567 (N_8567,N_7893,N_7195);
nor U8568 (N_8568,N_7044,N_7560);
nor U8569 (N_8569,N_7877,N_7483);
nor U8570 (N_8570,N_7151,N_7867);
and U8571 (N_8571,N_7153,N_7598);
and U8572 (N_8572,N_7233,N_7565);
nand U8573 (N_8573,N_7076,N_7216);
nor U8574 (N_8574,N_7419,N_7059);
or U8575 (N_8575,N_7282,N_7641);
or U8576 (N_8576,N_7508,N_7619);
nand U8577 (N_8577,N_7453,N_7954);
or U8578 (N_8578,N_7868,N_7148);
or U8579 (N_8579,N_7890,N_7716);
or U8580 (N_8580,N_7522,N_7193);
or U8581 (N_8581,N_7421,N_7583);
nor U8582 (N_8582,N_7184,N_7253);
or U8583 (N_8583,N_7447,N_7103);
and U8584 (N_8584,N_7627,N_7881);
nor U8585 (N_8585,N_7084,N_7348);
and U8586 (N_8586,N_7584,N_7572);
nor U8587 (N_8587,N_7613,N_7310);
nand U8588 (N_8588,N_7463,N_7040);
nand U8589 (N_8589,N_7107,N_7007);
nor U8590 (N_8590,N_7853,N_7611);
or U8591 (N_8591,N_7835,N_7845);
nand U8592 (N_8592,N_7910,N_7283);
or U8593 (N_8593,N_7144,N_7005);
xor U8594 (N_8594,N_7709,N_7416);
or U8595 (N_8595,N_7192,N_7794);
xnor U8596 (N_8596,N_7348,N_7002);
and U8597 (N_8597,N_7588,N_7889);
xor U8598 (N_8598,N_7874,N_7008);
nand U8599 (N_8599,N_7185,N_7086);
or U8600 (N_8600,N_7266,N_7119);
or U8601 (N_8601,N_7989,N_7320);
and U8602 (N_8602,N_7645,N_7752);
nor U8603 (N_8603,N_7855,N_7341);
nand U8604 (N_8604,N_7999,N_7556);
nor U8605 (N_8605,N_7920,N_7887);
or U8606 (N_8606,N_7921,N_7007);
and U8607 (N_8607,N_7302,N_7047);
or U8608 (N_8608,N_7520,N_7922);
or U8609 (N_8609,N_7607,N_7447);
and U8610 (N_8610,N_7052,N_7210);
nor U8611 (N_8611,N_7527,N_7191);
nand U8612 (N_8612,N_7730,N_7501);
nand U8613 (N_8613,N_7522,N_7981);
and U8614 (N_8614,N_7463,N_7830);
or U8615 (N_8615,N_7846,N_7930);
or U8616 (N_8616,N_7114,N_7602);
nand U8617 (N_8617,N_7886,N_7022);
nand U8618 (N_8618,N_7756,N_7049);
nand U8619 (N_8619,N_7594,N_7444);
nor U8620 (N_8620,N_7677,N_7174);
nor U8621 (N_8621,N_7051,N_7254);
or U8622 (N_8622,N_7325,N_7064);
nand U8623 (N_8623,N_7479,N_7324);
nand U8624 (N_8624,N_7743,N_7399);
or U8625 (N_8625,N_7321,N_7358);
and U8626 (N_8626,N_7037,N_7118);
and U8627 (N_8627,N_7105,N_7991);
nor U8628 (N_8628,N_7899,N_7556);
nand U8629 (N_8629,N_7545,N_7702);
nor U8630 (N_8630,N_7180,N_7984);
nand U8631 (N_8631,N_7244,N_7475);
xor U8632 (N_8632,N_7390,N_7844);
or U8633 (N_8633,N_7965,N_7186);
nand U8634 (N_8634,N_7146,N_7463);
nand U8635 (N_8635,N_7796,N_7293);
nand U8636 (N_8636,N_7998,N_7159);
nor U8637 (N_8637,N_7285,N_7163);
and U8638 (N_8638,N_7972,N_7602);
nor U8639 (N_8639,N_7299,N_7979);
and U8640 (N_8640,N_7742,N_7871);
nand U8641 (N_8641,N_7485,N_7688);
nor U8642 (N_8642,N_7109,N_7686);
xor U8643 (N_8643,N_7820,N_7997);
or U8644 (N_8644,N_7186,N_7107);
nand U8645 (N_8645,N_7468,N_7552);
nand U8646 (N_8646,N_7101,N_7930);
nand U8647 (N_8647,N_7067,N_7212);
xnor U8648 (N_8648,N_7637,N_7738);
nand U8649 (N_8649,N_7840,N_7032);
nand U8650 (N_8650,N_7886,N_7689);
nand U8651 (N_8651,N_7387,N_7151);
or U8652 (N_8652,N_7645,N_7145);
xnor U8653 (N_8653,N_7343,N_7523);
or U8654 (N_8654,N_7777,N_7860);
nor U8655 (N_8655,N_7880,N_7750);
nor U8656 (N_8656,N_7094,N_7748);
nor U8657 (N_8657,N_7852,N_7238);
xnor U8658 (N_8658,N_7872,N_7986);
and U8659 (N_8659,N_7084,N_7514);
xnor U8660 (N_8660,N_7138,N_7203);
nand U8661 (N_8661,N_7586,N_7548);
or U8662 (N_8662,N_7896,N_7031);
or U8663 (N_8663,N_7962,N_7653);
nand U8664 (N_8664,N_7024,N_7727);
xnor U8665 (N_8665,N_7584,N_7330);
or U8666 (N_8666,N_7173,N_7284);
nand U8667 (N_8667,N_7906,N_7310);
or U8668 (N_8668,N_7266,N_7022);
nor U8669 (N_8669,N_7849,N_7202);
or U8670 (N_8670,N_7430,N_7397);
nor U8671 (N_8671,N_7803,N_7449);
nand U8672 (N_8672,N_7631,N_7698);
and U8673 (N_8673,N_7088,N_7125);
nand U8674 (N_8674,N_7624,N_7671);
or U8675 (N_8675,N_7592,N_7793);
nand U8676 (N_8676,N_7276,N_7066);
or U8677 (N_8677,N_7017,N_7456);
or U8678 (N_8678,N_7475,N_7721);
nor U8679 (N_8679,N_7136,N_7233);
nand U8680 (N_8680,N_7754,N_7460);
and U8681 (N_8681,N_7918,N_7879);
and U8682 (N_8682,N_7487,N_7222);
or U8683 (N_8683,N_7539,N_7713);
nor U8684 (N_8684,N_7232,N_7787);
and U8685 (N_8685,N_7581,N_7967);
or U8686 (N_8686,N_7282,N_7253);
and U8687 (N_8687,N_7671,N_7025);
xnor U8688 (N_8688,N_7907,N_7289);
or U8689 (N_8689,N_7224,N_7920);
nor U8690 (N_8690,N_7868,N_7675);
or U8691 (N_8691,N_7861,N_7693);
nor U8692 (N_8692,N_7000,N_7477);
nand U8693 (N_8693,N_7951,N_7096);
and U8694 (N_8694,N_7263,N_7071);
and U8695 (N_8695,N_7899,N_7139);
and U8696 (N_8696,N_7080,N_7654);
nand U8697 (N_8697,N_7221,N_7588);
nand U8698 (N_8698,N_7580,N_7333);
nand U8699 (N_8699,N_7977,N_7721);
and U8700 (N_8700,N_7732,N_7211);
nand U8701 (N_8701,N_7545,N_7035);
nor U8702 (N_8702,N_7493,N_7016);
or U8703 (N_8703,N_7655,N_7062);
nor U8704 (N_8704,N_7638,N_7741);
nor U8705 (N_8705,N_7991,N_7308);
or U8706 (N_8706,N_7443,N_7296);
nor U8707 (N_8707,N_7339,N_7251);
nor U8708 (N_8708,N_7695,N_7094);
nor U8709 (N_8709,N_7398,N_7353);
or U8710 (N_8710,N_7680,N_7577);
nand U8711 (N_8711,N_7661,N_7518);
nand U8712 (N_8712,N_7876,N_7717);
nand U8713 (N_8713,N_7151,N_7643);
nor U8714 (N_8714,N_7429,N_7119);
or U8715 (N_8715,N_7574,N_7459);
and U8716 (N_8716,N_7743,N_7301);
or U8717 (N_8717,N_7467,N_7085);
and U8718 (N_8718,N_7282,N_7059);
xor U8719 (N_8719,N_7305,N_7033);
or U8720 (N_8720,N_7941,N_7888);
or U8721 (N_8721,N_7528,N_7485);
or U8722 (N_8722,N_7710,N_7480);
xnor U8723 (N_8723,N_7052,N_7389);
nand U8724 (N_8724,N_7144,N_7380);
nand U8725 (N_8725,N_7907,N_7173);
nor U8726 (N_8726,N_7134,N_7443);
nand U8727 (N_8727,N_7370,N_7192);
or U8728 (N_8728,N_7985,N_7817);
xor U8729 (N_8729,N_7795,N_7690);
nand U8730 (N_8730,N_7817,N_7773);
nor U8731 (N_8731,N_7765,N_7812);
xnor U8732 (N_8732,N_7430,N_7135);
nand U8733 (N_8733,N_7685,N_7463);
xnor U8734 (N_8734,N_7745,N_7966);
nand U8735 (N_8735,N_7384,N_7548);
nor U8736 (N_8736,N_7566,N_7612);
nand U8737 (N_8737,N_7348,N_7214);
nand U8738 (N_8738,N_7874,N_7110);
or U8739 (N_8739,N_7766,N_7753);
xor U8740 (N_8740,N_7275,N_7601);
and U8741 (N_8741,N_7929,N_7144);
and U8742 (N_8742,N_7398,N_7764);
nand U8743 (N_8743,N_7925,N_7673);
nor U8744 (N_8744,N_7944,N_7714);
nor U8745 (N_8745,N_7527,N_7414);
nand U8746 (N_8746,N_7062,N_7257);
or U8747 (N_8747,N_7205,N_7743);
nand U8748 (N_8748,N_7643,N_7647);
nor U8749 (N_8749,N_7169,N_7935);
nand U8750 (N_8750,N_7813,N_7072);
xnor U8751 (N_8751,N_7086,N_7088);
xnor U8752 (N_8752,N_7377,N_7126);
nand U8753 (N_8753,N_7388,N_7804);
xnor U8754 (N_8754,N_7107,N_7031);
nor U8755 (N_8755,N_7234,N_7939);
or U8756 (N_8756,N_7099,N_7085);
or U8757 (N_8757,N_7237,N_7556);
nor U8758 (N_8758,N_7295,N_7442);
or U8759 (N_8759,N_7400,N_7959);
nor U8760 (N_8760,N_7656,N_7405);
and U8761 (N_8761,N_7605,N_7351);
or U8762 (N_8762,N_7527,N_7149);
nand U8763 (N_8763,N_7583,N_7003);
xnor U8764 (N_8764,N_7559,N_7020);
or U8765 (N_8765,N_7463,N_7476);
nor U8766 (N_8766,N_7404,N_7989);
xor U8767 (N_8767,N_7678,N_7534);
nor U8768 (N_8768,N_7501,N_7411);
or U8769 (N_8769,N_7878,N_7858);
xor U8770 (N_8770,N_7698,N_7903);
nand U8771 (N_8771,N_7853,N_7020);
nor U8772 (N_8772,N_7742,N_7783);
and U8773 (N_8773,N_7046,N_7767);
nand U8774 (N_8774,N_7097,N_7076);
nor U8775 (N_8775,N_7224,N_7565);
nand U8776 (N_8776,N_7789,N_7291);
nor U8777 (N_8777,N_7105,N_7171);
and U8778 (N_8778,N_7071,N_7829);
xor U8779 (N_8779,N_7501,N_7783);
nor U8780 (N_8780,N_7833,N_7270);
or U8781 (N_8781,N_7089,N_7497);
nor U8782 (N_8782,N_7872,N_7914);
nor U8783 (N_8783,N_7499,N_7548);
nand U8784 (N_8784,N_7382,N_7171);
nand U8785 (N_8785,N_7192,N_7116);
nand U8786 (N_8786,N_7466,N_7740);
nor U8787 (N_8787,N_7465,N_7129);
nor U8788 (N_8788,N_7269,N_7965);
xor U8789 (N_8789,N_7586,N_7958);
nor U8790 (N_8790,N_7008,N_7981);
or U8791 (N_8791,N_7233,N_7547);
nand U8792 (N_8792,N_7384,N_7396);
and U8793 (N_8793,N_7885,N_7522);
xor U8794 (N_8794,N_7248,N_7859);
nor U8795 (N_8795,N_7658,N_7300);
nand U8796 (N_8796,N_7412,N_7976);
nor U8797 (N_8797,N_7672,N_7156);
or U8798 (N_8798,N_7859,N_7681);
and U8799 (N_8799,N_7368,N_7170);
nand U8800 (N_8800,N_7330,N_7573);
and U8801 (N_8801,N_7381,N_7869);
xor U8802 (N_8802,N_7770,N_7554);
or U8803 (N_8803,N_7317,N_7340);
or U8804 (N_8804,N_7850,N_7601);
or U8805 (N_8805,N_7471,N_7367);
nor U8806 (N_8806,N_7117,N_7839);
xnor U8807 (N_8807,N_7575,N_7795);
nor U8808 (N_8808,N_7597,N_7319);
and U8809 (N_8809,N_7707,N_7824);
or U8810 (N_8810,N_7585,N_7869);
and U8811 (N_8811,N_7088,N_7780);
or U8812 (N_8812,N_7086,N_7625);
nor U8813 (N_8813,N_7993,N_7897);
nor U8814 (N_8814,N_7038,N_7883);
nor U8815 (N_8815,N_7676,N_7418);
nor U8816 (N_8816,N_7099,N_7826);
nand U8817 (N_8817,N_7132,N_7758);
nand U8818 (N_8818,N_7020,N_7181);
nor U8819 (N_8819,N_7140,N_7851);
or U8820 (N_8820,N_7783,N_7104);
or U8821 (N_8821,N_7351,N_7997);
nor U8822 (N_8822,N_7007,N_7911);
and U8823 (N_8823,N_7244,N_7247);
nor U8824 (N_8824,N_7995,N_7281);
or U8825 (N_8825,N_7616,N_7594);
nor U8826 (N_8826,N_7067,N_7991);
and U8827 (N_8827,N_7273,N_7566);
xor U8828 (N_8828,N_7512,N_7329);
and U8829 (N_8829,N_7706,N_7862);
nor U8830 (N_8830,N_7377,N_7755);
nor U8831 (N_8831,N_7237,N_7071);
xor U8832 (N_8832,N_7351,N_7251);
nor U8833 (N_8833,N_7516,N_7944);
nand U8834 (N_8834,N_7127,N_7906);
and U8835 (N_8835,N_7551,N_7237);
nand U8836 (N_8836,N_7513,N_7615);
and U8837 (N_8837,N_7704,N_7733);
nand U8838 (N_8838,N_7604,N_7353);
and U8839 (N_8839,N_7256,N_7880);
nor U8840 (N_8840,N_7795,N_7567);
or U8841 (N_8841,N_7791,N_7185);
nor U8842 (N_8842,N_7200,N_7384);
xor U8843 (N_8843,N_7178,N_7802);
or U8844 (N_8844,N_7554,N_7482);
nor U8845 (N_8845,N_7413,N_7436);
nand U8846 (N_8846,N_7046,N_7070);
nand U8847 (N_8847,N_7708,N_7764);
and U8848 (N_8848,N_7067,N_7160);
or U8849 (N_8849,N_7190,N_7672);
nand U8850 (N_8850,N_7718,N_7290);
nor U8851 (N_8851,N_7152,N_7329);
and U8852 (N_8852,N_7639,N_7546);
and U8853 (N_8853,N_7550,N_7769);
nor U8854 (N_8854,N_7984,N_7608);
or U8855 (N_8855,N_7546,N_7683);
and U8856 (N_8856,N_7918,N_7044);
or U8857 (N_8857,N_7955,N_7748);
and U8858 (N_8858,N_7083,N_7006);
xor U8859 (N_8859,N_7878,N_7322);
nor U8860 (N_8860,N_7291,N_7074);
nor U8861 (N_8861,N_7732,N_7780);
nor U8862 (N_8862,N_7867,N_7716);
nand U8863 (N_8863,N_7034,N_7405);
xnor U8864 (N_8864,N_7420,N_7237);
or U8865 (N_8865,N_7890,N_7589);
nand U8866 (N_8866,N_7613,N_7567);
nor U8867 (N_8867,N_7649,N_7662);
and U8868 (N_8868,N_7508,N_7827);
nand U8869 (N_8869,N_7258,N_7872);
nor U8870 (N_8870,N_7113,N_7356);
nor U8871 (N_8871,N_7219,N_7462);
nor U8872 (N_8872,N_7461,N_7139);
nand U8873 (N_8873,N_7552,N_7601);
nor U8874 (N_8874,N_7219,N_7818);
nor U8875 (N_8875,N_7548,N_7664);
and U8876 (N_8876,N_7727,N_7725);
and U8877 (N_8877,N_7869,N_7645);
and U8878 (N_8878,N_7823,N_7799);
nand U8879 (N_8879,N_7258,N_7353);
nor U8880 (N_8880,N_7545,N_7920);
nor U8881 (N_8881,N_7490,N_7547);
and U8882 (N_8882,N_7033,N_7961);
xnor U8883 (N_8883,N_7327,N_7629);
nor U8884 (N_8884,N_7961,N_7060);
nor U8885 (N_8885,N_7963,N_7625);
or U8886 (N_8886,N_7826,N_7822);
or U8887 (N_8887,N_7659,N_7792);
nor U8888 (N_8888,N_7104,N_7100);
and U8889 (N_8889,N_7470,N_7323);
xnor U8890 (N_8890,N_7745,N_7972);
or U8891 (N_8891,N_7320,N_7669);
nand U8892 (N_8892,N_7080,N_7822);
or U8893 (N_8893,N_7731,N_7901);
nor U8894 (N_8894,N_7904,N_7057);
nor U8895 (N_8895,N_7843,N_7590);
nand U8896 (N_8896,N_7241,N_7887);
nor U8897 (N_8897,N_7251,N_7478);
or U8898 (N_8898,N_7062,N_7839);
or U8899 (N_8899,N_7577,N_7785);
or U8900 (N_8900,N_7969,N_7691);
and U8901 (N_8901,N_7522,N_7306);
nor U8902 (N_8902,N_7669,N_7279);
nand U8903 (N_8903,N_7914,N_7220);
or U8904 (N_8904,N_7920,N_7962);
nand U8905 (N_8905,N_7681,N_7401);
xnor U8906 (N_8906,N_7266,N_7409);
or U8907 (N_8907,N_7906,N_7576);
or U8908 (N_8908,N_7960,N_7723);
or U8909 (N_8909,N_7296,N_7185);
xor U8910 (N_8910,N_7189,N_7271);
nand U8911 (N_8911,N_7802,N_7269);
and U8912 (N_8912,N_7271,N_7068);
xor U8913 (N_8913,N_7138,N_7328);
or U8914 (N_8914,N_7689,N_7421);
nand U8915 (N_8915,N_7003,N_7839);
or U8916 (N_8916,N_7035,N_7022);
or U8917 (N_8917,N_7455,N_7348);
or U8918 (N_8918,N_7330,N_7341);
nor U8919 (N_8919,N_7884,N_7504);
nand U8920 (N_8920,N_7439,N_7817);
nor U8921 (N_8921,N_7447,N_7667);
nor U8922 (N_8922,N_7092,N_7988);
and U8923 (N_8923,N_7707,N_7533);
nand U8924 (N_8924,N_7919,N_7071);
and U8925 (N_8925,N_7288,N_7557);
or U8926 (N_8926,N_7847,N_7312);
and U8927 (N_8927,N_7120,N_7620);
xor U8928 (N_8928,N_7684,N_7634);
and U8929 (N_8929,N_7778,N_7948);
nand U8930 (N_8930,N_7196,N_7144);
nor U8931 (N_8931,N_7900,N_7511);
nand U8932 (N_8932,N_7131,N_7376);
and U8933 (N_8933,N_7339,N_7602);
nand U8934 (N_8934,N_7537,N_7286);
or U8935 (N_8935,N_7015,N_7201);
or U8936 (N_8936,N_7437,N_7592);
nand U8937 (N_8937,N_7703,N_7511);
xnor U8938 (N_8938,N_7157,N_7489);
nand U8939 (N_8939,N_7444,N_7474);
and U8940 (N_8940,N_7864,N_7329);
nor U8941 (N_8941,N_7917,N_7728);
and U8942 (N_8942,N_7301,N_7877);
nand U8943 (N_8943,N_7922,N_7048);
nor U8944 (N_8944,N_7085,N_7932);
nand U8945 (N_8945,N_7116,N_7807);
and U8946 (N_8946,N_7879,N_7309);
nand U8947 (N_8947,N_7915,N_7064);
and U8948 (N_8948,N_7875,N_7142);
nand U8949 (N_8949,N_7561,N_7302);
and U8950 (N_8950,N_7655,N_7821);
nand U8951 (N_8951,N_7126,N_7586);
nor U8952 (N_8952,N_7370,N_7843);
nand U8953 (N_8953,N_7648,N_7288);
nand U8954 (N_8954,N_7232,N_7259);
nand U8955 (N_8955,N_7656,N_7576);
and U8956 (N_8956,N_7716,N_7756);
or U8957 (N_8957,N_7603,N_7665);
and U8958 (N_8958,N_7808,N_7647);
nand U8959 (N_8959,N_7606,N_7865);
nand U8960 (N_8960,N_7656,N_7174);
nand U8961 (N_8961,N_7134,N_7197);
and U8962 (N_8962,N_7312,N_7791);
nor U8963 (N_8963,N_7791,N_7800);
or U8964 (N_8964,N_7577,N_7320);
nor U8965 (N_8965,N_7547,N_7692);
or U8966 (N_8966,N_7328,N_7348);
nand U8967 (N_8967,N_7191,N_7360);
nor U8968 (N_8968,N_7101,N_7962);
nor U8969 (N_8969,N_7473,N_7396);
and U8970 (N_8970,N_7462,N_7412);
nor U8971 (N_8971,N_7837,N_7079);
nand U8972 (N_8972,N_7918,N_7014);
and U8973 (N_8973,N_7223,N_7370);
and U8974 (N_8974,N_7401,N_7690);
nor U8975 (N_8975,N_7073,N_7895);
and U8976 (N_8976,N_7508,N_7551);
and U8977 (N_8977,N_7478,N_7645);
or U8978 (N_8978,N_7696,N_7240);
nand U8979 (N_8979,N_7058,N_7045);
or U8980 (N_8980,N_7612,N_7173);
or U8981 (N_8981,N_7320,N_7144);
or U8982 (N_8982,N_7373,N_7514);
and U8983 (N_8983,N_7500,N_7023);
and U8984 (N_8984,N_7662,N_7386);
or U8985 (N_8985,N_7515,N_7595);
and U8986 (N_8986,N_7893,N_7911);
xor U8987 (N_8987,N_7312,N_7563);
xnor U8988 (N_8988,N_7097,N_7048);
or U8989 (N_8989,N_7365,N_7625);
nand U8990 (N_8990,N_7101,N_7008);
and U8991 (N_8991,N_7278,N_7069);
and U8992 (N_8992,N_7023,N_7966);
or U8993 (N_8993,N_7697,N_7202);
and U8994 (N_8994,N_7807,N_7781);
nand U8995 (N_8995,N_7907,N_7600);
or U8996 (N_8996,N_7127,N_7280);
and U8997 (N_8997,N_7613,N_7645);
xnor U8998 (N_8998,N_7701,N_7634);
nor U8999 (N_8999,N_7057,N_7977);
and U9000 (N_9000,N_8907,N_8996);
xnor U9001 (N_9001,N_8259,N_8779);
nor U9002 (N_9002,N_8335,N_8309);
and U9003 (N_9003,N_8227,N_8545);
xnor U9004 (N_9004,N_8810,N_8372);
and U9005 (N_9005,N_8363,N_8154);
nor U9006 (N_9006,N_8846,N_8013);
nand U9007 (N_9007,N_8539,N_8870);
nor U9008 (N_9008,N_8394,N_8754);
and U9009 (N_9009,N_8404,N_8410);
and U9010 (N_9010,N_8225,N_8074);
xor U9011 (N_9011,N_8934,N_8274);
or U9012 (N_9012,N_8703,N_8078);
nor U9013 (N_9013,N_8106,N_8733);
nand U9014 (N_9014,N_8064,N_8627);
or U9015 (N_9015,N_8306,N_8911);
nand U9016 (N_9016,N_8378,N_8576);
or U9017 (N_9017,N_8774,N_8347);
nor U9018 (N_9018,N_8128,N_8617);
nor U9019 (N_9019,N_8801,N_8088);
or U9020 (N_9020,N_8023,N_8280);
nand U9021 (N_9021,N_8654,N_8805);
xnor U9022 (N_9022,N_8294,N_8340);
nand U9023 (N_9023,N_8398,N_8928);
nand U9024 (N_9024,N_8022,N_8011);
or U9025 (N_9025,N_8897,N_8483);
nor U9026 (N_9026,N_8960,N_8898);
nand U9027 (N_9027,N_8766,N_8058);
or U9028 (N_9028,N_8656,N_8828);
or U9029 (N_9029,N_8256,N_8217);
nor U9030 (N_9030,N_8111,N_8487);
and U9031 (N_9031,N_8970,N_8508);
nor U9032 (N_9032,N_8091,N_8524);
nor U9033 (N_9033,N_8126,N_8231);
nor U9034 (N_9034,N_8051,N_8437);
or U9035 (N_9035,N_8269,N_8476);
and U9036 (N_9036,N_8124,N_8788);
and U9037 (N_9037,N_8729,N_8165);
nand U9038 (N_9038,N_8370,N_8209);
nor U9039 (N_9039,N_8017,N_8270);
nor U9040 (N_9040,N_8691,N_8208);
nor U9041 (N_9041,N_8332,N_8602);
or U9042 (N_9042,N_8246,N_8042);
nor U9043 (N_9043,N_8122,N_8169);
and U9044 (N_9044,N_8344,N_8419);
xnor U9045 (N_9045,N_8250,N_8546);
nand U9046 (N_9046,N_8678,N_8661);
nand U9047 (N_9047,N_8860,N_8040);
nor U9048 (N_9048,N_8355,N_8232);
xnor U9049 (N_9049,N_8257,N_8178);
or U9050 (N_9050,N_8299,N_8686);
or U9051 (N_9051,N_8515,N_8995);
nor U9052 (N_9052,N_8093,N_8226);
or U9053 (N_9053,N_8955,N_8374);
and U9054 (N_9054,N_8830,N_8184);
xor U9055 (N_9055,N_8035,N_8041);
and U9056 (N_9056,N_8454,N_8004);
nand U9057 (N_9057,N_8929,N_8979);
and U9058 (N_9058,N_8429,N_8424);
nor U9059 (N_9059,N_8940,N_8599);
or U9060 (N_9060,N_8525,N_8851);
and U9061 (N_9061,N_8720,N_8358);
and U9062 (N_9062,N_8314,N_8997);
and U9063 (N_9063,N_8393,N_8481);
nand U9064 (N_9064,N_8382,N_8685);
and U9065 (N_9065,N_8914,N_8859);
or U9066 (N_9066,N_8189,N_8477);
nand U9067 (N_9067,N_8186,N_8384);
nor U9068 (N_9068,N_8200,N_8185);
and U9069 (N_9069,N_8281,N_8988);
nand U9070 (N_9070,N_8760,N_8461);
nor U9071 (N_9071,N_8562,N_8839);
nor U9072 (N_9072,N_8066,N_8591);
nand U9073 (N_9073,N_8919,N_8367);
nand U9074 (N_9074,N_8923,N_8390);
and U9075 (N_9075,N_8359,N_8116);
and U9076 (N_9076,N_8303,N_8962);
nand U9077 (N_9077,N_8565,N_8119);
and U9078 (N_9078,N_8808,N_8882);
and U9079 (N_9079,N_8557,N_8386);
nor U9080 (N_9080,N_8307,N_8762);
or U9081 (N_9081,N_8141,N_8236);
nand U9082 (N_9082,N_8071,N_8594);
or U9083 (N_9083,N_8373,N_8784);
nand U9084 (N_9084,N_8908,N_8123);
and U9085 (N_9085,N_8473,N_8060);
nand U9086 (N_9086,N_8688,N_8974);
nand U9087 (N_9087,N_8936,N_8958);
or U9088 (N_9088,N_8098,N_8913);
nor U9089 (N_9089,N_8567,N_8712);
nor U9090 (N_9090,N_8369,N_8021);
nor U9091 (N_9091,N_8036,N_8138);
nor U9092 (N_9092,N_8149,N_8694);
or U9093 (N_9093,N_8749,N_8713);
or U9094 (N_9094,N_8511,N_8059);
nor U9095 (N_9095,N_8350,N_8318);
xor U9096 (N_9096,N_8939,N_8527);
or U9097 (N_9097,N_8738,N_8921);
nor U9098 (N_9098,N_8623,N_8849);
nand U9099 (N_9099,N_8304,N_8379);
nand U9100 (N_9100,N_8388,N_8652);
nand U9101 (N_9101,N_8696,N_8285);
or U9102 (N_9102,N_8467,N_8218);
or U9103 (N_9103,N_8994,N_8628);
nor U9104 (N_9104,N_8811,N_8560);
or U9105 (N_9105,N_8224,N_8864);
and U9106 (N_9106,N_8737,N_8789);
nor U9107 (N_9107,N_8173,N_8311);
nand U9108 (N_9108,N_8118,N_8957);
or U9109 (N_9109,N_8422,N_8426);
nor U9110 (N_9110,N_8619,N_8799);
or U9111 (N_9111,N_8360,N_8778);
nor U9112 (N_9112,N_8951,N_8079);
nand U9113 (N_9113,N_8679,N_8544);
and U9114 (N_9114,N_8814,N_8276);
or U9115 (N_9115,N_8287,N_8411);
nand U9116 (N_9116,N_8201,N_8781);
nor U9117 (N_9117,N_8109,N_8170);
or U9118 (N_9118,N_8620,N_8491);
xor U9119 (N_9119,N_8931,N_8573);
or U9120 (N_9120,N_8765,N_8353);
and U9121 (N_9121,N_8077,N_8438);
nand U9122 (N_9122,N_8146,N_8847);
or U9123 (N_9123,N_8858,N_8721);
xor U9124 (N_9124,N_8107,N_8183);
or U9125 (N_9125,N_8547,N_8967);
nand U9126 (N_9126,N_8181,N_8191);
nand U9127 (N_9127,N_8197,N_8439);
and U9128 (N_9128,N_8717,N_8484);
nor U9129 (N_9129,N_8991,N_8513);
or U9130 (N_9130,N_8272,N_8728);
or U9131 (N_9131,N_8552,N_8884);
nor U9132 (N_9132,N_8159,N_8924);
or U9133 (N_9133,N_8930,N_8655);
nor U9134 (N_9134,N_8470,N_8650);
and U9135 (N_9135,N_8094,N_8603);
nor U9136 (N_9136,N_8220,N_8012);
xor U9137 (N_9137,N_8877,N_8657);
and U9138 (N_9138,N_8130,N_8081);
xor U9139 (N_9139,N_8708,N_8229);
nor U9140 (N_9140,N_8516,N_8521);
nand U9141 (N_9141,N_8916,N_8982);
or U9142 (N_9142,N_8561,N_8407);
xor U9143 (N_9143,N_8613,N_8634);
and U9144 (N_9144,N_8406,N_8937);
nand U9145 (N_9145,N_8647,N_8326);
nand U9146 (N_9146,N_8512,N_8635);
and U9147 (N_9147,N_8669,N_8554);
nor U9148 (N_9148,N_8179,N_8769);
or U9149 (N_9149,N_8767,N_8443);
nand U9150 (N_9150,N_8726,N_8313);
nand U9151 (N_9151,N_8659,N_8056);
or U9152 (N_9152,N_8342,N_8168);
or U9153 (N_9153,N_8329,N_8984);
xor U9154 (N_9154,N_8216,N_8945);
nand U9155 (N_9155,N_8289,N_8638);
nor U9156 (N_9156,N_8277,N_8596);
and U9157 (N_9157,N_8442,N_8947);
nand U9158 (N_9158,N_8015,N_8356);
nor U9159 (N_9159,N_8549,N_8933);
nand U9160 (N_9160,N_8687,N_8609);
and U9161 (N_9161,N_8469,N_8776);
and U9162 (N_9162,N_8574,N_8338);
or U9163 (N_9163,N_8075,N_8938);
nor U9164 (N_9164,N_8155,N_8380);
or U9165 (N_9165,N_8027,N_8291);
and U9166 (N_9166,N_8867,N_8998);
nand U9167 (N_9167,N_8537,N_8676);
nor U9168 (N_9168,N_8785,N_8876);
and U9169 (N_9169,N_8813,N_8375);
or U9170 (N_9170,N_8742,N_8089);
nor U9171 (N_9171,N_8435,N_8850);
or U9172 (N_9172,N_8436,N_8063);
xnor U9173 (N_9173,N_8145,N_8462);
or U9174 (N_9174,N_8275,N_8920);
nor U9175 (N_9175,N_8608,N_8297);
or U9176 (N_9176,N_8211,N_8626);
nand U9177 (N_9177,N_8698,N_8744);
and U9178 (N_9178,N_8631,N_8577);
or U9179 (N_9179,N_8134,N_8301);
nor U9180 (N_9180,N_8362,N_8731);
nand U9181 (N_9181,N_8503,N_8381);
nor U9182 (N_9182,N_8653,N_8743);
or U9183 (N_9183,N_8018,N_8963);
or U9184 (N_9184,N_8777,N_8457);
xnor U9185 (N_9185,N_8556,N_8910);
nor U9186 (N_9186,N_8589,N_8330);
xor U9187 (N_9187,N_8065,N_8964);
nor U9188 (N_9188,N_8684,N_8976);
nand U9189 (N_9189,N_8621,N_8357);
and U9190 (N_9190,N_8214,N_8113);
and U9191 (N_9191,N_8352,N_8010);
and U9192 (N_9192,N_8090,N_8474);
or U9193 (N_9193,N_8495,N_8346);
and U9194 (N_9194,N_8579,N_8566);
xnor U9195 (N_9195,N_8153,N_8792);
or U9196 (N_9196,N_8247,N_8981);
xnor U9197 (N_9197,N_8701,N_8000);
or U9198 (N_9198,N_8049,N_8416);
or U9199 (N_9199,N_8383,N_8003);
xnor U9200 (N_9200,N_8499,N_8115);
xnor U9201 (N_9201,N_8399,N_8400);
nand U9202 (N_9202,N_8233,N_8842);
and U9203 (N_9203,N_8016,N_8334);
nor U9204 (N_9204,N_8674,N_8459);
and U9205 (N_9205,N_8798,N_8192);
nand U9206 (N_9206,N_8905,N_8990);
or U9207 (N_9207,N_8328,N_8782);
nand U9208 (N_9208,N_8033,N_8219);
nor U9209 (N_9209,N_8651,N_8447);
and U9210 (N_9210,N_8592,N_8230);
nor U9211 (N_9211,N_8711,N_8543);
nand U9212 (N_9212,N_8127,N_8317);
and U9213 (N_9213,N_8992,N_8880);
nand U9214 (N_9214,N_8194,N_8868);
nand U9215 (N_9215,N_8188,N_8019);
nor U9216 (N_9216,N_8826,N_8148);
xnor U9217 (N_9217,N_8031,N_8395);
nor U9218 (N_9218,N_8665,N_8520);
and U9219 (N_9219,N_8180,N_8497);
or U9220 (N_9220,N_8879,N_8458);
nand U9221 (N_9221,N_8752,N_8986);
and U9222 (N_9222,N_8862,N_8260);
nor U9223 (N_9223,N_8709,N_8008);
nand U9224 (N_9224,N_8377,N_8486);
nor U9225 (N_9225,N_8136,N_8172);
and U9226 (N_9226,N_8104,N_8946);
nand U9227 (N_9227,N_8812,N_8434);
xor U9228 (N_9228,N_8187,N_8349);
nor U9229 (N_9229,N_8604,N_8327);
or U9230 (N_9230,N_8135,N_8643);
nor U9231 (N_9231,N_8848,N_8542);
or U9232 (N_9232,N_8034,N_8455);
nor U9233 (N_9233,N_8875,N_8150);
or U9234 (N_9234,N_8530,N_8922);
nor U9235 (N_9235,N_8787,N_8954);
xor U9236 (N_9236,N_8465,N_8872);
nand U9237 (N_9237,N_8649,N_8783);
nor U9238 (N_9238,N_8587,N_8593);
and U9239 (N_9239,N_8615,N_8772);
and U9240 (N_9240,N_8892,N_8658);
nor U9241 (N_9241,N_8255,N_8293);
and U9242 (N_9242,N_8244,N_8509);
xnor U9243 (N_9243,N_8901,N_8087);
nand U9244 (N_9244,N_8949,N_8501);
and U9245 (N_9245,N_8702,N_8730);
nand U9246 (N_9246,N_8271,N_8747);
and U9247 (N_9247,N_8973,N_8639);
or U9248 (N_9248,N_8129,N_8715);
nand U9249 (N_9249,N_8748,N_8727);
or U9250 (N_9250,N_8054,N_8909);
or U9251 (N_9251,N_8773,N_8614);
or U9252 (N_9252,N_8529,N_8835);
and U9253 (N_9253,N_8719,N_8563);
or U9254 (N_9254,N_8953,N_8820);
and U9255 (N_9255,N_8637,N_8047);
nor U9256 (N_9256,N_8866,N_8354);
nand U9257 (N_9257,N_8993,N_8348);
nor U9258 (N_9258,N_8223,N_8475);
nand U9259 (N_9259,N_8020,N_8261);
nor U9260 (N_9260,N_8445,N_8863);
nor U9261 (N_9261,N_8132,N_8433);
nand U9262 (N_9262,N_8452,N_8736);
nor U9263 (N_9263,N_8072,N_8391);
nand U9264 (N_9264,N_8489,N_8836);
nand U9265 (N_9265,N_8239,N_8213);
nor U9266 (N_9266,N_8468,N_8724);
nor U9267 (N_9267,N_8874,N_8944);
and U9268 (N_9268,N_8630,N_8258);
xor U9269 (N_9269,N_8112,N_8807);
xnor U9270 (N_9270,N_8403,N_8550);
or U9271 (N_9271,N_8800,N_8158);
nor U9272 (N_9272,N_8286,N_8199);
or U9273 (N_9273,N_8775,N_8283);
and U9274 (N_9274,N_8043,N_8941);
nand U9275 (N_9275,N_8084,N_8324);
nand U9276 (N_9276,N_8926,N_8662);
and U9277 (N_9277,N_8666,N_8840);
or U9278 (N_9278,N_8590,N_8315);
and U9279 (N_9279,N_8558,N_8401);
nor U9280 (N_9280,N_8045,N_8298);
nor U9281 (N_9281,N_8222,N_8413);
and U9282 (N_9282,N_8819,N_8405);
and U9283 (N_9283,N_8450,N_8718);
xor U9284 (N_9284,N_8584,N_8086);
nand U9285 (N_9285,N_8507,N_8918);
nor U9286 (N_9286,N_8430,N_8580);
and U9287 (N_9287,N_8305,N_8073);
and U9288 (N_9288,N_8163,N_8843);
xor U9289 (N_9289,N_8266,N_8460);
or U9290 (N_9290,N_8221,N_8999);
nand U9291 (N_9291,N_8758,N_8680);
and U9292 (N_9292,N_8444,N_8364);
nand U9293 (N_9293,N_8166,N_8714);
nor U9294 (N_9294,N_8095,N_8841);
nor U9295 (N_9295,N_8682,N_8583);
or U9296 (N_9296,N_8253,N_8818);
and U9297 (N_9297,N_8716,N_8345);
nand U9298 (N_9298,N_8001,N_8618);
and U9299 (N_9299,N_8570,N_8177);
nor U9300 (N_9300,N_8479,N_8959);
and U9301 (N_9301,N_8108,N_8797);
nand U9302 (N_9302,N_8493,N_8616);
nand U9303 (N_9303,N_8241,N_8983);
nand U9304 (N_9304,N_8190,N_8735);
nand U9305 (N_9305,N_8564,N_8541);
or U9306 (N_9306,N_8157,N_8480);
nand U9307 (N_9307,N_8642,N_8553);
or U9308 (N_9308,N_8500,N_8829);
nand U9309 (N_9309,N_8068,N_8548);
and U9310 (N_9310,N_8531,N_8598);
nand U9311 (N_9311,N_8279,N_8014);
nand U9312 (N_9312,N_8409,N_8965);
nor U9313 (N_9313,N_8741,N_8196);
and U9314 (N_9314,N_8645,N_8816);
and U9315 (N_9315,N_8425,N_8795);
xnor U9316 (N_9316,N_8977,N_8446);
nand U9317 (N_9317,N_8228,N_8510);
nor U9318 (N_9318,N_8024,N_8532);
nor U9319 (N_9319,N_8252,N_8092);
xnor U9320 (N_9320,N_8641,N_8295);
or U9321 (N_9321,N_8873,N_8025);
and U9322 (N_9322,N_8677,N_8895);
or U9323 (N_9323,N_8496,N_8292);
or U9324 (N_9324,N_8451,N_8822);
nand U9325 (N_9325,N_8249,N_8823);
and U9326 (N_9326,N_8707,N_8915);
nor U9327 (N_9327,N_8526,N_8368);
nor U9328 (N_9328,N_8756,N_8421);
nand U9329 (N_9329,N_8710,N_8026);
nor U9330 (N_9330,N_8827,N_8648);
or U9331 (N_9331,N_8174,N_8336);
xnor U9332 (N_9332,N_8853,N_8505);
nor U9333 (N_9333,N_8817,N_8575);
xnor U9334 (N_9334,N_8935,N_8578);
and U9335 (N_9335,N_8597,N_8248);
and U9336 (N_9336,N_8193,N_8551);
nor U9337 (N_9337,N_8831,N_8453);
nand U9338 (N_9338,N_8069,N_8402);
nand U9339 (N_9339,N_8053,N_8449);
nand U9340 (N_9340,N_8278,N_8855);
nand U9341 (N_9341,N_8725,N_8878);
and U9342 (N_9342,N_8706,N_8240);
nand U9343 (N_9343,N_8825,N_8952);
and U9344 (N_9344,N_8343,N_8062);
or U9345 (N_9345,N_8588,N_8005);
and U9346 (N_9346,N_8610,N_8761);
or U9347 (N_9347,N_8950,N_8282);
xor U9348 (N_9348,N_8131,N_8699);
or U9349 (N_9349,N_8205,N_8385);
nand U9350 (N_9350,N_8085,N_8692);
nor U9351 (N_9351,N_8753,N_8423);
or U9352 (N_9352,N_8366,N_8917);
and U9353 (N_9353,N_8504,N_8441);
nor U9354 (N_9354,N_8176,N_8943);
nor U9355 (N_9355,N_8412,N_8485);
nor U9356 (N_9356,N_8103,N_8755);
nor U9357 (N_9357,N_8865,N_8308);
nor U9358 (N_9358,N_8414,N_8606);
or U9359 (N_9359,N_8883,N_8514);
and U9360 (N_9360,N_8243,N_8055);
nor U9361 (N_9361,N_8365,N_8534);
xor U9362 (N_9362,N_8151,N_8478);
or U9363 (N_9363,N_8881,N_8492);
nand U9364 (N_9364,N_8331,N_8582);
xnor U9365 (N_9365,N_8607,N_8082);
and U9366 (N_9366,N_8771,N_8147);
nand U9367 (N_9367,N_8900,N_8764);
nor U9368 (N_9368,N_8806,N_8745);
and U9369 (N_9369,N_8175,N_8763);
and U9370 (N_9370,N_8076,N_8300);
nand U9371 (N_9371,N_8632,N_8912);
and U9372 (N_9372,N_8972,N_8804);
and U9373 (N_9373,N_8927,N_8740);
nand U9374 (N_9374,N_8466,N_8268);
nor U9375 (N_9375,N_8683,N_8768);
nand U9376 (N_9376,N_8083,N_8844);
nand U9377 (N_9377,N_8202,N_8312);
nand U9378 (N_9378,N_8237,N_8009);
nand U9379 (N_9379,N_8044,N_8284);
or U9380 (N_9380,N_8431,N_8490);
or U9381 (N_9381,N_8262,N_8971);
and U9382 (N_9382,N_8793,N_8052);
or U9383 (N_9383,N_8581,N_8668);
and U9384 (N_9384,N_8096,N_8100);
and U9385 (N_9385,N_8519,N_8207);
and U9386 (N_9386,N_8671,N_8705);
nor U9387 (N_9387,N_8288,N_8322);
and U9388 (N_9388,N_8114,N_8102);
nor U9389 (N_9389,N_8050,N_8101);
nor U9390 (N_9390,N_8408,N_8057);
and U9391 (N_9391,N_8029,N_8522);
or U9392 (N_9392,N_8675,N_8803);
and U9393 (N_9393,N_8889,N_8361);
and U9394 (N_9394,N_8472,N_8039);
nand U9395 (N_9395,N_8061,N_8622);
xor U9396 (N_9396,N_8689,N_8321);
and U9397 (N_9397,N_8857,N_8975);
nand U9398 (N_9398,N_8387,N_8488);
xnor U9399 (N_9399,N_8376,N_8833);
nor U9400 (N_9400,N_8746,N_8969);
and U9401 (N_9401,N_8624,N_8471);
or U9402 (N_9402,N_8734,N_8320);
nand U9403 (N_9403,N_8886,N_8245);
and U9404 (N_9404,N_8234,N_8167);
nor U9405 (N_9405,N_8203,N_8533);
nand U9406 (N_9406,N_8903,N_8586);
and U9407 (N_9407,N_8099,N_8722);
and U9408 (N_9408,N_8144,N_8948);
and U9409 (N_9409,N_8750,N_8251);
nand U9410 (N_9410,N_8852,N_8601);
nor U9411 (N_9411,N_8681,N_8821);
xor U9412 (N_9412,N_8834,N_8371);
and U9413 (N_9413,N_8837,N_8296);
nor U9414 (N_9414,N_8757,N_8891);
and U9415 (N_9415,N_8006,N_8673);
nor U9416 (N_9416,N_8448,N_8535);
and U9417 (N_9417,N_8418,N_8142);
nor U9418 (N_9418,N_8629,N_8323);
or U9419 (N_9419,N_8732,N_8351);
nor U9420 (N_9420,N_8885,N_8464);
and U9421 (N_9421,N_8871,N_8536);
or U9422 (N_9422,N_8572,N_8143);
and U9423 (N_9423,N_8397,N_8007);
or U9424 (N_9424,N_8980,N_8456);
nor U9425 (N_9425,N_8796,N_8759);
or U9426 (N_9426,N_8117,N_8636);
and U9427 (N_9427,N_8290,N_8046);
or U9428 (N_9428,N_8463,N_8595);
and U9429 (N_9429,N_8032,N_8125);
or U9430 (N_9430,N_8585,N_8518);
nand U9431 (N_9431,N_8978,N_8600);
nor U9432 (N_9432,N_8815,N_8161);
nor U9433 (N_9433,N_8791,N_8786);
and U9434 (N_9434,N_8802,N_8670);
and U9435 (N_9435,N_8838,N_8700);
nand U9436 (N_9436,N_8182,N_8506);
nor U9437 (N_9437,N_8568,N_8212);
or U9438 (N_9438,N_8198,N_8273);
nand U9439 (N_9439,N_8646,N_8832);
nor U9440 (N_9440,N_8896,N_8152);
and U9441 (N_9441,N_8887,N_8693);
or U9442 (N_9442,N_8569,N_8316);
or U9443 (N_9443,N_8028,N_8325);
or U9444 (N_9444,N_8644,N_8097);
xor U9445 (N_9445,N_8845,N_8235);
nand U9446 (N_9446,N_8440,N_8389);
nand U9447 (N_9447,N_8048,N_8140);
nand U9448 (N_9448,N_8660,N_8195);
nor U9449 (N_9449,N_8968,N_8133);
nor U9450 (N_9450,N_8392,N_8110);
xor U9451 (N_9451,N_8672,N_8899);
nand U9452 (N_9452,N_8210,N_8987);
nor U9453 (N_9453,N_8961,N_8482);
nor U9454 (N_9454,N_8664,N_8861);
and U9455 (N_9455,N_8751,N_8697);
and U9456 (N_9456,N_8121,N_8517);
nor U9457 (N_9457,N_8164,N_8932);
and U9458 (N_9458,N_8310,N_8498);
nor U9459 (N_9459,N_8555,N_8906);
or U9460 (N_9460,N_8341,N_8396);
and U9461 (N_9461,N_8605,N_8942);
nor U9462 (N_9462,N_8612,N_8319);
or U9463 (N_9463,N_8494,N_8571);
nor U9464 (N_9464,N_8427,N_8030);
xnor U9465 (N_9465,N_8540,N_8162);
nand U9466 (N_9466,N_8264,N_8856);
or U9467 (N_9467,N_8204,N_8267);
and U9468 (N_9468,N_8302,N_8502);
and U9469 (N_9469,N_8037,N_8238);
or U9470 (N_9470,N_8611,N_8254);
nand U9471 (N_9471,N_8902,N_8067);
nand U9472 (N_9472,N_8888,N_8432);
and U9473 (N_9473,N_8215,N_8770);
and U9474 (N_9474,N_8869,N_8739);
and U9475 (N_9475,N_8704,N_8854);
and U9476 (N_9476,N_8428,N_8080);
nor U9477 (N_9477,N_8415,N_8780);
nand U9478 (N_9478,N_8038,N_8824);
and U9479 (N_9479,N_8120,N_8723);
nor U9480 (N_9480,N_8538,N_8890);
nor U9481 (N_9481,N_8690,N_8985);
nor U9482 (N_9482,N_8956,N_8790);
nand U9483 (N_9483,N_8242,N_8633);
and U9484 (N_9484,N_8139,N_8989);
nor U9485 (N_9485,N_8523,N_8265);
or U9486 (N_9486,N_8625,N_8966);
nand U9487 (N_9487,N_8339,N_8663);
nor U9488 (N_9488,N_8904,N_8667);
xor U9489 (N_9489,N_8263,N_8925);
or U9490 (N_9490,N_8137,N_8171);
or U9491 (N_9491,N_8206,N_8559);
nor U9492 (N_9492,N_8105,N_8070);
nor U9493 (N_9493,N_8156,N_8893);
nand U9494 (N_9494,N_8809,N_8002);
nand U9495 (N_9495,N_8640,N_8695);
or U9496 (N_9496,N_8894,N_8417);
or U9497 (N_9497,N_8420,N_8333);
nor U9498 (N_9498,N_8528,N_8160);
or U9499 (N_9499,N_8794,N_8337);
nand U9500 (N_9500,N_8485,N_8898);
nor U9501 (N_9501,N_8210,N_8342);
nand U9502 (N_9502,N_8311,N_8337);
or U9503 (N_9503,N_8242,N_8497);
nand U9504 (N_9504,N_8639,N_8908);
nor U9505 (N_9505,N_8206,N_8657);
and U9506 (N_9506,N_8844,N_8926);
or U9507 (N_9507,N_8069,N_8950);
xor U9508 (N_9508,N_8421,N_8996);
and U9509 (N_9509,N_8150,N_8323);
nand U9510 (N_9510,N_8439,N_8778);
xor U9511 (N_9511,N_8122,N_8092);
or U9512 (N_9512,N_8923,N_8818);
or U9513 (N_9513,N_8266,N_8911);
nand U9514 (N_9514,N_8133,N_8837);
and U9515 (N_9515,N_8256,N_8727);
or U9516 (N_9516,N_8058,N_8312);
nor U9517 (N_9517,N_8425,N_8682);
nand U9518 (N_9518,N_8309,N_8799);
and U9519 (N_9519,N_8791,N_8728);
nor U9520 (N_9520,N_8318,N_8938);
xor U9521 (N_9521,N_8968,N_8934);
or U9522 (N_9522,N_8034,N_8520);
xnor U9523 (N_9523,N_8136,N_8970);
or U9524 (N_9524,N_8267,N_8104);
nand U9525 (N_9525,N_8431,N_8435);
xor U9526 (N_9526,N_8897,N_8279);
nor U9527 (N_9527,N_8059,N_8456);
nor U9528 (N_9528,N_8465,N_8952);
nand U9529 (N_9529,N_8620,N_8916);
nor U9530 (N_9530,N_8281,N_8292);
nand U9531 (N_9531,N_8212,N_8810);
nand U9532 (N_9532,N_8132,N_8763);
nand U9533 (N_9533,N_8596,N_8679);
nand U9534 (N_9534,N_8129,N_8704);
xor U9535 (N_9535,N_8866,N_8811);
nor U9536 (N_9536,N_8815,N_8222);
nand U9537 (N_9537,N_8749,N_8576);
nor U9538 (N_9538,N_8857,N_8054);
nand U9539 (N_9539,N_8262,N_8487);
nor U9540 (N_9540,N_8523,N_8468);
or U9541 (N_9541,N_8928,N_8170);
nand U9542 (N_9542,N_8842,N_8756);
xnor U9543 (N_9543,N_8793,N_8226);
or U9544 (N_9544,N_8011,N_8519);
nand U9545 (N_9545,N_8802,N_8933);
nand U9546 (N_9546,N_8921,N_8878);
nand U9547 (N_9547,N_8447,N_8645);
nand U9548 (N_9548,N_8386,N_8100);
or U9549 (N_9549,N_8495,N_8130);
nand U9550 (N_9550,N_8478,N_8722);
and U9551 (N_9551,N_8700,N_8366);
nand U9552 (N_9552,N_8642,N_8991);
or U9553 (N_9553,N_8528,N_8984);
nand U9554 (N_9554,N_8158,N_8642);
nor U9555 (N_9555,N_8265,N_8967);
or U9556 (N_9556,N_8786,N_8283);
nand U9557 (N_9557,N_8680,N_8622);
nor U9558 (N_9558,N_8506,N_8082);
nor U9559 (N_9559,N_8164,N_8257);
and U9560 (N_9560,N_8267,N_8913);
or U9561 (N_9561,N_8082,N_8028);
nor U9562 (N_9562,N_8092,N_8460);
xnor U9563 (N_9563,N_8605,N_8270);
or U9564 (N_9564,N_8679,N_8051);
nand U9565 (N_9565,N_8424,N_8799);
xnor U9566 (N_9566,N_8339,N_8842);
or U9567 (N_9567,N_8116,N_8385);
and U9568 (N_9568,N_8578,N_8483);
or U9569 (N_9569,N_8406,N_8132);
nand U9570 (N_9570,N_8635,N_8320);
nand U9571 (N_9571,N_8551,N_8874);
xor U9572 (N_9572,N_8388,N_8868);
nand U9573 (N_9573,N_8399,N_8354);
and U9574 (N_9574,N_8235,N_8639);
nand U9575 (N_9575,N_8925,N_8569);
nor U9576 (N_9576,N_8242,N_8608);
and U9577 (N_9577,N_8985,N_8693);
and U9578 (N_9578,N_8913,N_8995);
nand U9579 (N_9579,N_8500,N_8147);
nor U9580 (N_9580,N_8990,N_8292);
nand U9581 (N_9581,N_8006,N_8084);
nand U9582 (N_9582,N_8245,N_8686);
nand U9583 (N_9583,N_8161,N_8576);
or U9584 (N_9584,N_8839,N_8240);
nor U9585 (N_9585,N_8671,N_8412);
nand U9586 (N_9586,N_8649,N_8734);
xnor U9587 (N_9587,N_8179,N_8658);
or U9588 (N_9588,N_8548,N_8405);
nand U9589 (N_9589,N_8987,N_8710);
xnor U9590 (N_9590,N_8520,N_8821);
or U9591 (N_9591,N_8205,N_8806);
xnor U9592 (N_9592,N_8120,N_8012);
nand U9593 (N_9593,N_8312,N_8024);
nand U9594 (N_9594,N_8814,N_8785);
nand U9595 (N_9595,N_8395,N_8616);
and U9596 (N_9596,N_8163,N_8591);
nand U9597 (N_9597,N_8370,N_8219);
nand U9598 (N_9598,N_8857,N_8198);
nand U9599 (N_9599,N_8269,N_8556);
and U9600 (N_9600,N_8949,N_8492);
or U9601 (N_9601,N_8952,N_8064);
or U9602 (N_9602,N_8330,N_8851);
or U9603 (N_9603,N_8126,N_8117);
or U9604 (N_9604,N_8575,N_8795);
or U9605 (N_9605,N_8990,N_8861);
nand U9606 (N_9606,N_8306,N_8468);
nor U9607 (N_9607,N_8256,N_8252);
or U9608 (N_9608,N_8337,N_8701);
nand U9609 (N_9609,N_8351,N_8581);
and U9610 (N_9610,N_8114,N_8549);
nand U9611 (N_9611,N_8011,N_8554);
nor U9612 (N_9612,N_8489,N_8364);
or U9613 (N_9613,N_8062,N_8180);
xnor U9614 (N_9614,N_8020,N_8574);
and U9615 (N_9615,N_8259,N_8899);
or U9616 (N_9616,N_8253,N_8924);
nor U9617 (N_9617,N_8838,N_8321);
and U9618 (N_9618,N_8872,N_8414);
xnor U9619 (N_9619,N_8092,N_8330);
or U9620 (N_9620,N_8964,N_8048);
nor U9621 (N_9621,N_8298,N_8624);
nor U9622 (N_9622,N_8245,N_8534);
and U9623 (N_9623,N_8833,N_8116);
or U9624 (N_9624,N_8679,N_8334);
nand U9625 (N_9625,N_8896,N_8380);
and U9626 (N_9626,N_8799,N_8743);
nand U9627 (N_9627,N_8633,N_8863);
or U9628 (N_9628,N_8064,N_8370);
nor U9629 (N_9629,N_8473,N_8538);
nor U9630 (N_9630,N_8704,N_8724);
and U9631 (N_9631,N_8072,N_8286);
nor U9632 (N_9632,N_8198,N_8687);
and U9633 (N_9633,N_8450,N_8956);
or U9634 (N_9634,N_8723,N_8787);
nor U9635 (N_9635,N_8279,N_8125);
nor U9636 (N_9636,N_8552,N_8907);
or U9637 (N_9637,N_8154,N_8149);
nand U9638 (N_9638,N_8208,N_8894);
nand U9639 (N_9639,N_8624,N_8808);
and U9640 (N_9640,N_8774,N_8307);
xor U9641 (N_9641,N_8530,N_8349);
and U9642 (N_9642,N_8261,N_8877);
or U9643 (N_9643,N_8775,N_8795);
xor U9644 (N_9644,N_8394,N_8496);
nor U9645 (N_9645,N_8616,N_8835);
and U9646 (N_9646,N_8715,N_8773);
nor U9647 (N_9647,N_8605,N_8227);
or U9648 (N_9648,N_8463,N_8780);
or U9649 (N_9649,N_8454,N_8808);
nand U9650 (N_9650,N_8987,N_8314);
xnor U9651 (N_9651,N_8852,N_8759);
or U9652 (N_9652,N_8339,N_8371);
or U9653 (N_9653,N_8330,N_8577);
and U9654 (N_9654,N_8055,N_8722);
nor U9655 (N_9655,N_8717,N_8149);
nand U9656 (N_9656,N_8798,N_8061);
and U9657 (N_9657,N_8446,N_8676);
nand U9658 (N_9658,N_8534,N_8858);
nand U9659 (N_9659,N_8487,N_8414);
and U9660 (N_9660,N_8999,N_8003);
or U9661 (N_9661,N_8525,N_8596);
or U9662 (N_9662,N_8901,N_8813);
nor U9663 (N_9663,N_8252,N_8005);
or U9664 (N_9664,N_8725,N_8302);
xnor U9665 (N_9665,N_8093,N_8289);
nor U9666 (N_9666,N_8402,N_8360);
and U9667 (N_9667,N_8834,N_8916);
or U9668 (N_9668,N_8561,N_8751);
nand U9669 (N_9669,N_8645,N_8178);
nor U9670 (N_9670,N_8653,N_8012);
and U9671 (N_9671,N_8698,N_8972);
and U9672 (N_9672,N_8873,N_8887);
nor U9673 (N_9673,N_8355,N_8825);
nand U9674 (N_9674,N_8793,N_8027);
xnor U9675 (N_9675,N_8422,N_8110);
and U9676 (N_9676,N_8091,N_8299);
nor U9677 (N_9677,N_8936,N_8115);
nor U9678 (N_9678,N_8676,N_8896);
nand U9679 (N_9679,N_8134,N_8928);
and U9680 (N_9680,N_8202,N_8536);
or U9681 (N_9681,N_8658,N_8080);
xor U9682 (N_9682,N_8825,N_8654);
nand U9683 (N_9683,N_8551,N_8649);
nor U9684 (N_9684,N_8781,N_8534);
xor U9685 (N_9685,N_8580,N_8253);
xor U9686 (N_9686,N_8393,N_8304);
or U9687 (N_9687,N_8637,N_8342);
nor U9688 (N_9688,N_8893,N_8915);
nor U9689 (N_9689,N_8176,N_8512);
and U9690 (N_9690,N_8557,N_8372);
and U9691 (N_9691,N_8269,N_8710);
nand U9692 (N_9692,N_8473,N_8596);
nor U9693 (N_9693,N_8971,N_8910);
nand U9694 (N_9694,N_8189,N_8550);
nand U9695 (N_9695,N_8658,N_8940);
nor U9696 (N_9696,N_8659,N_8369);
nor U9697 (N_9697,N_8535,N_8342);
xor U9698 (N_9698,N_8652,N_8556);
nor U9699 (N_9699,N_8326,N_8645);
nor U9700 (N_9700,N_8948,N_8923);
or U9701 (N_9701,N_8758,N_8983);
nor U9702 (N_9702,N_8929,N_8640);
and U9703 (N_9703,N_8501,N_8718);
and U9704 (N_9704,N_8522,N_8125);
xor U9705 (N_9705,N_8732,N_8550);
or U9706 (N_9706,N_8483,N_8402);
and U9707 (N_9707,N_8151,N_8808);
xnor U9708 (N_9708,N_8451,N_8958);
nand U9709 (N_9709,N_8656,N_8584);
nand U9710 (N_9710,N_8808,N_8337);
or U9711 (N_9711,N_8054,N_8563);
and U9712 (N_9712,N_8171,N_8222);
or U9713 (N_9713,N_8055,N_8986);
xnor U9714 (N_9714,N_8289,N_8330);
and U9715 (N_9715,N_8424,N_8081);
nand U9716 (N_9716,N_8406,N_8860);
and U9717 (N_9717,N_8181,N_8286);
nand U9718 (N_9718,N_8279,N_8957);
xnor U9719 (N_9719,N_8878,N_8104);
nand U9720 (N_9720,N_8828,N_8038);
nand U9721 (N_9721,N_8034,N_8789);
and U9722 (N_9722,N_8839,N_8946);
and U9723 (N_9723,N_8118,N_8163);
nor U9724 (N_9724,N_8379,N_8637);
nand U9725 (N_9725,N_8643,N_8319);
xor U9726 (N_9726,N_8866,N_8463);
nand U9727 (N_9727,N_8036,N_8446);
nand U9728 (N_9728,N_8178,N_8029);
xnor U9729 (N_9729,N_8757,N_8869);
nand U9730 (N_9730,N_8235,N_8262);
xor U9731 (N_9731,N_8910,N_8249);
or U9732 (N_9732,N_8736,N_8345);
nand U9733 (N_9733,N_8158,N_8862);
nor U9734 (N_9734,N_8000,N_8201);
and U9735 (N_9735,N_8897,N_8110);
and U9736 (N_9736,N_8102,N_8714);
nor U9737 (N_9737,N_8141,N_8882);
and U9738 (N_9738,N_8504,N_8875);
or U9739 (N_9739,N_8462,N_8082);
and U9740 (N_9740,N_8840,N_8871);
nor U9741 (N_9741,N_8720,N_8007);
and U9742 (N_9742,N_8187,N_8516);
or U9743 (N_9743,N_8544,N_8624);
nand U9744 (N_9744,N_8631,N_8522);
and U9745 (N_9745,N_8498,N_8909);
and U9746 (N_9746,N_8344,N_8617);
nor U9747 (N_9747,N_8908,N_8294);
and U9748 (N_9748,N_8770,N_8302);
nor U9749 (N_9749,N_8764,N_8142);
nand U9750 (N_9750,N_8407,N_8773);
nand U9751 (N_9751,N_8451,N_8739);
or U9752 (N_9752,N_8138,N_8730);
and U9753 (N_9753,N_8107,N_8287);
or U9754 (N_9754,N_8388,N_8114);
nor U9755 (N_9755,N_8467,N_8281);
nor U9756 (N_9756,N_8627,N_8605);
xor U9757 (N_9757,N_8519,N_8575);
and U9758 (N_9758,N_8501,N_8395);
nand U9759 (N_9759,N_8619,N_8741);
nand U9760 (N_9760,N_8517,N_8049);
nor U9761 (N_9761,N_8276,N_8365);
or U9762 (N_9762,N_8797,N_8602);
or U9763 (N_9763,N_8030,N_8135);
or U9764 (N_9764,N_8945,N_8416);
and U9765 (N_9765,N_8356,N_8074);
nor U9766 (N_9766,N_8562,N_8941);
nor U9767 (N_9767,N_8341,N_8668);
xor U9768 (N_9768,N_8450,N_8015);
and U9769 (N_9769,N_8005,N_8319);
nor U9770 (N_9770,N_8559,N_8368);
nor U9771 (N_9771,N_8327,N_8858);
or U9772 (N_9772,N_8653,N_8714);
nand U9773 (N_9773,N_8377,N_8346);
or U9774 (N_9774,N_8035,N_8218);
or U9775 (N_9775,N_8515,N_8699);
nor U9776 (N_9776,N_8888,N_8030);
and U9777 (N_9777,N_8256,N_8182);
or U9778 (N_9778,N_8546,N_8566);
or U9779 (N_9779,N_8448,N_8882);
and U9780 (N_9780,N_8350,N_8717);
and U9781 (N_9781,N_8337,N_8235);
nand U9782 (N_9782,N_8161,N_8011);
or U9783 (N_9783,N_8589,N_8869);
nand U9784 (N_9784,N_8371,N_8148);
or U9785 (N_9785,N_8482,N_8908);
or U9786 (N_9786,N_8702,N_8860);
nor U9787 (N_9787,N_8651,N_8587);
and U9788 (N_9788,N_8825,N_8643);
nand U9789 (N_9789,N_8279,N_8782);
and U9790 (N_9790,N_8865,N_8473);
or U9791 (N_9791,N_8974,N_8007);
and U9792 (N_9792,N_8642,N_8734);
xor U9793 (N_9793,N_8523,N_8357);
and U9794 (N_9794,N_8930,N_8926);
nor U9795 (N_9795,N_8829,N_8588);
and U9796 (N_9796,N_8354,N_8225);
nand U9797 (N_9797,N_8613,N_8143);
nand U9798 (N_9798,N_8175,N_8793);
or U9799 (N_9799,N_8281,N_8692);
and U9800 (N_9800,N_8633,N_8768);
or U9801 (N_9801,N_8828,N_8278);
xor U9802 (N_9802,N_8101,N_8838);
or U9803 (N_9803,N_8513,N_8844);
and U9804 (N_9804,N_8524,N_8250);
nand U9805 (N_9805,N_8021,N_8060);
nor U9806 (N_9806,N_8034,N_8768);
or U9807 (N_9807,N_8479,N_8717);
xor U9808 (N_9808,N_8658,N_8009);
nand U9809 (N_9809,N_8712,N_8520);
nor U9810 (N_9810,N_8339,N_8529);
nand U9811 (N_9811,N_8145,N_8899);
nor U9812 (N_9812,N_8845,N_8583);
or U9813 (N_9813,N_8633,N_8430);
nor U9814 (N_9814,N_8459,N_8324);
xnor U9815 (N_9815,N_8691,N_8554);
nor U9816 (N_9816,N_8722,N_8543);
nand U9817 (N_9817,N_8357,N_8864);
or U9818 (N_9818,N_8382,N_8792);
nand U9819 (N_9819,N_8307,N_8562);
xor U9820 (N_9820,N_8982,N_8740);
nor U9821 (N_9821,N_8574,N_8647);
nand U9822 (N_9822,N_8232,N_8260);
and U9823 (N_9823,N_8712,N_8528);
nand U9824 (N_9824,N_8414,N_8643);
or U9825 (N_9825,N_8165,N_8368);
nand U9826 (N_9826,N_8680,N_8337);
nor U9827 (N_9827,N_8517,N_8877);
and U9828 (N_9828,N_8636,N_8737);
nor U9829 (N_9829,N_8625,N_8795);
nor U9830 (N_9830,N_8133,N_8913);
nor U9831 (N_9831,N_8537,N_8990);
nand U9832 (N_9832,N_8157,N_8594);
or U9833 (N_9833,N_8391,N_8780);
or U9834 (N_9834,N_8072,N_8635);
nor U9835 (N_9835,N_8246,N_8969);
and U9836 (N_9836,N_8959,N_8302);
and U9837 (N_9837,N_8045,N_8704);
nand U9838 (N_9838,N_8037,N_8283);
nor U9839 (N_9839,N_8373,N_8994);
nand U9840 (N_9840,N_8071,N_8724);
and U9841 (N_9841,N_8349,N_8402);
nor U9842 (N_9842,N_8642,N_8429);
or U9843 (N_9843,N_8416,N_8054);
or U9844 (N_9844,N_8320,N_8341);
or U9845 (N_9845,N_8754,N_8784);
nor U9846 (N_9846,N_8123,N_8965);
or U9847 (N_9847,N_8617,N_8485);
or U9848 (N_9848,N_8531,N_8928);
and U9849 (N_9849,N_8182,N_8964);
xor U9850 (N_9850,N_8219,N_8603);
xnor U9851 (N_9851,N_8826,N_8899);
xnor U9852 (N_9852,N_8246,N_8571);
or U9853 (N_9853,N_8121,N_8928);
nor U9854 (N_9854,N_8761,N_8984);
or U9855 (N_9855,N_8596,N_8673);
nand U9856 (N_9856,N_8438,N_8143);
nand U9857 (N_9857,N_8357,N_8059);
and U9858 (N_9858,N_8971,N_8040);
or U9859 (N_9859,N_8022,N_8583);
nor U9860 (N_9860,N_8153,N_8428);
xor U9861 (N_9861,N_8698,N_8218);
nand U9862 (N_9862,N_8353,N_8559);
or U9863 (N_9863,N_8121,N_8161);
nor U9864 (N_9864,N_8738,N_8182);
or U9865 (N_9865,N_8881,N_8518);
nor U9866 (N_9866,N_8587,N_8406);
nand U9867 (N_9867,N_8802,N_8070);
and U9868 (N_9868,N_8846,N_8806);
and U9869 (N_9869,N_8074,N_8809);
nand U9870 (N_9870,N_8167,N_8282);
or U9871 (N_9871,N_8464,N_8243);
or U9872 (N_9872,N_8586,N_8243);
and U9873 (N_9873,N_8851,N_8942);
nand U9874 (N_9874,N_8329,N_8419);
nand U9875 (N_9875,N_8568,N_8174);
nor U9876 (N_9876,N_8013,N_8110);
nor U9877 (N_9877,N_8527,N_8730);
or U9878 (N_9878,N_8533,N_8388);
or U9879 (N_9879,N_8404,N_8180);
and U9880 (N_9880,N_8985,N_8176);
nand U9881 (N_9881,N_8242,N_8278);
nand U9882 (N_9882,N_8646,N_8893);
xnor U9883 (N_9883,N_8792,N_8905);
nand U9884 (N_9884,N_8600,N_8959);
and U9885 (N_9885,N_8283,N_8967);
xnor U9886 (N_9886,N_8854,N_8368);
nand U9887 (N_9887,N_8068,N_8443);
nor U9888 (N_9888,N_8322,N_8300);
xnor U9889 (N_9889,N_8189,N_8391);
or U9890 (N_9890,N_8887,N_8058);
or U9891 (N_9891,N_8951,N_8471);
or U9892 (N_9892,N_8587,N_8682);
and U9893 (N_9893,N_8798,N_8769);
and U9894 (N_9894,N_8530,N_8842);
and U9895 (N_9895,N_8832,N_8395);
nor U9896 (N_9896,N_8885,N_8156);
nand U9897 (N_9897,N_8166,N_8665);
and U9898 (N_9898,N_8524,N_8601);
nor U9899 (N_9899,N_8971,N_8444);
or U9900 (N_9900,N_8048,N_8786);
nand U9901 (N_9901,N_8828,N_8111);
or U9902 (N_9902,N_8534,N_8035);
xor U9903 (N_9903,N_8219,N_8488);
nor U9904 (N_9904,N_8393,N_8792);
or U9905 (N_9905,N_8502,N_8224);
and U9906 (N_9906,N_8462,N_8582);
and U9907 (N_9907,N_8335,N_8850);
xnor U9908 (N_9908,N_8364,N_8225);
nand U9909 (N_9909,N_8068,N_8511);
or U9910 (N_9910,N_8037,N_8156);
and U9911 (N_9911,N_8127,N_8500);
or U9912 (N_9912,N_8081,N_8986);
and U9913 (N_9913,N_8138,N_8934);
and U9914 (N_9914,N_8983,N_8539);
xnor U9915 (N_9915,N_8760,N_8604);
and U9916 (N_9916,N_8593,N_8501);
nor U9917 (N_9917,N_8655,N_8517);
or U9918 (N_9918,N_8814,N_8343);
and U9919 (N_9919,N_8690,N_8062);
nand U9920 (N_9920,N_8174,N_8272);
or U9921 (N_9921,N_8156,N_8696);
or U9922 (N_9922,N_8871,N_8006);
or U9923 (N_9923,N_8764,N_8055);
nor U9924 (N_9924,N_8790,N_8213);
and U9925 (N_9925,N_8093,N_8551);
or U9926 (N_9926,N_8728,N_8221);
or U9927 (N_9927,N_8246,N_8323);
and U9928 (N_9928,N_8923,N_8293);
nand U9929 (N_9929,N_8135,N_8725);
and U9930 (N_9930,N_8069,N_8312);
and U9931 (N_9931,N_8574,N_8306);
xnor U9932 (N_9932,N_8541,N_8468);
or U9933 (N_9933,N_8273,N_8789);
and U9934 (N_9934,N_8247,N_8263);
nand U9935 (N_9935,N_8326,N_8425);
xnor U9936 (N_9936,N_8102,N_8310);
or U9937 (N_9937,N_8311,N_8683);
nand U9938 (N_9938,N_8508,N_8393);
nor U9939 (N_9939,N_8828,N_8733);
xnor U9940 (N_9940,N_8058,N_8031);
and U9941 (N_9941,N_8908,N_8069);
nand U9942 (N_9942,N_8525,N_8799);
xnor U9943 (N_9943,N_8294,N_8654);
xnor U9944 (N_9944,N_8694,N_8000);
xor U9945 (N_9945,N_8874,N_8013);
nor U9946 (N_9946,N_8268,N_8733);
nand U9947 (N_9947,N_8275,N_8553);
nand U9948 (N_9948,N_8908,N_8558);
nor U9949 (N_9949,N_8973,N_8396);
nand U9950 (N_9950,N_8181,N_8014);
or U9951 (N_9951,N_8160,N_8600);
or U9952 (N_9952,N_8692,N_8691);
or U9953 (N_9953,N_8798,N_8681);
or U9954 (N_9954,N_8793,N_8836);
xnor U9955 (N_9955,N_8259,N_8611);
nor U9956 (N_9956,N_8170,N_8245);
or U9957 (N_9957,N_8084,N_8616);
nor U9958 (N_9958,N_8098,N_8512);
and U9959 (N_9959,N_8083,N_8650);
or U9960 (N_9960,N_8506,N_8444);
and U9961 (N_9961,N_8634,N_8978);
nand U9962 (N_9962,N_8689,N_8906);
nand U9963 (N_9963,N_8433,N_8607);
nand U9964 (N_9964,N_8521,N_8988);
nand U9965 (N_9965,N_8165,N_8561);
nand U9966 (N_9966,N_8066,N_8795);
and U9967 (N_9967,N_8115,N_8040);
and U9968 (N_9968,N_8013,N_8014);
and U9969 (N_9969,N_8314,N_8282);
nor U9970 (N_9970,N_8852,N_8128);
nor U9971 (N_9971,N_8878,N_8206);
nand U9972 (N_9972,N_8959,N_8494);
or U9973 (N_9973,N_8473,N_8075);
nand U9974 (N_9974,N_8845,N_8313);
nand U9975 (N_9975,N_8708,N_8889);
or U9976 (N_9976,N_8525,N_8705);
and U9977 (N_9977,N_8228,N_8775);
nor U9978 (N_9978,N_8687,N_8162);
nor U9979 (N_9979,N_8436,N_8302);
or U9980 (N_9980,N_8336,N_8410);
nand U9981 (N_9981,N_8671,N_8498);
and U9982 (N_9982,N_8236,N_8204);
nor U9983 (N_9983,N_8720,N_8817);
nand U9984 (N_9984,N_8348,N_8035);
and U9985 (N_9985,N_8323,N_8646);
and U9986 (N_9986,N_8393,N_8617);
and U9987 (N_9987,N_8382,N_8627);
or U9988 (N_9988,N_8340,N_8782);
nor U9989 (N_9989,N_8705,N_8489);
xnor U9990 (N_9990,N_8600,N_8084);
nor U9991 (N_9991,N_8498,N_8739);
xor U9992 (N_9992,N_8444,N_8571);
nor U9993 (N_9993,N_8269,N_8910);
nor U9994 (N_9994,N_8175,N_8792);
and U9995 (N_9995,N_8070,N_8348);
nand U9996 (N_9996,N_8413,N_8104);
and U9997 (N_9997,N_8356,N_8062);
nor U9998 (N_9998,N_8635,N_8763);
and U9999 (N_9999,N_8002,N_8305);
nand UO_0 (O_0,N_9624,N_9908);
and UO_1 (O_1,N_9094,N_9698);
and UO_2 (O_2,N_9933,N_9174);
or UO_3 (O_3,N_9727,N_9447);
nor UO_4 (O_4,N_9921,N_9873);
or UO_5 (O_5,N_9822,N_9243);
xor UO_6 (O_6,N_9187,N_9758);
nor UO_7 (O_7,N_9423,N_9355);
xor UO_8 (O_8,N_9363,N_9362);
and UO_9 (O_9,N_9018,N_9345);
or UO_10 (O_10,N_9219,N_9204);
and UO_11 (O_11,N_9651,N_9022);
or UO_12 (O_12,N_9033,N_9769);
or UO_13 (O_13,N_9158,N_9878);
and UO_14 (O_14,N_9353,N_9124);
nor UO_15 (O_15,N_9713,N_9602);
nand UO_16 (O_16,N_9257,N_9482);
or UO_17 (O_17,N_9675,N_9852);
and UO_18 (O_18,N_9929,N_9129);
nor UO_19 (O_19,N_9863,N_9173);
xor UO_20 (O_20,N_9808,N_9207);
and UO_21 (O_21,N_9632,N_9048);
nand UO_22 (O_22,N_9284,N_9154);
or UO_23 (O_23,N_9339,N_9752);
nand UO_24 (O_24,N_9945,N_9637);
nand UO_25 (O_25,N_9568,N_9517);
nand UO_26 (O_26,N_9014,N_9025);
and UO_27 (O_27,N_9116,N_9749);
and UO_28 (O_28,N_9575,N_9202);
and UO_29 (O_29,N_9135,N_9098);
or UO_30 (O_30,N_9712,N_9398);
nand UO_31 (O_31,N_9413,N_9589);
nand UO_32 (O_32,N_9709,N_9601);
and UO_33 (O_33,N_9010,N_9816);
nand UO_34 (O_34,N_9036,N_9962);
nor UO_35 (O_35,N_9733,N_9839);
nor UO_36 (O_36,N_9114,N_9145);
and UO_37 (O_37,N_9854,N_9007);
xor UO_38 (O_38,N_9799,N_9058);
nor UO_39 (O_39,N_9842,N_9941);
xor UO_40 (O_40,N_9337,N_9740);
and UO_41 (O_41,N_9720,N_9288);
xor UO_42 (O_42,N_9907,N_9453);
or UO_43 (O_43,N_9293,N_9429);
or UO_44 (O_44,N_9618,N_9800);
and UO_45 (O_45,N_9461,N_9325);
nor UO_46 (O_46,N_9558,N_9235);
and UO_47 (O_47,N_9569,N_9894);
nand UO_48 (O_48,N_9579,N_9877);
or UO_49 (O_49,N_9732,N_9090);
or UO_50 (O_50,N_9326,N_9495);
nand UO_51 (O_51,N_9970,N_9797);
nand UO_52 (O_52,N_9920,N_9590);
nand UO_53 (O_53,N_9975,N_9350);
nor UO_54 (O_54,N_9346,N_9947);
or UO_55 (O_55,N_9383,N_9582);
nor UO_56 (O_56,N_9296,N_9703);
and UO_57 (O_57,N_9216,N_9109);
or UO_58 (O_58,N_9278,N_9315);
nor UO_59 (O_59,N_9859,N_9672);
or UO_60 (O_60,N_9684,N_9940);
xnor UO_61 (O_61,N_9678,N_9107);
nor UO_62 (O_62,N_9912,N_9340);
nand UO_63 (O_63,N_9327,N_9591);
and UO_64 (O_64,N_9400,N_9457);
and UO_65 (O_65,N_9131,N_9001);
nand UO_66 (O_66,N_9421,N_9371);
nor UO_67 (O_67,N_9404,N_9813);
and UO_68 (O_68,N_9702,N_9472);
nand UO_69 (O_69,N_9511,N_9742);
and UO_70 (O_70,N_9445,N_9016);
xnor UO_71 (O_71,N_9239,N_9984);
nand UO_72 (O_72,N_9711,N_9074);
nor UO_73 (O_73,N_9600,N_9963);
nor UO_74 (O_74,N_9256,N_9264);
and UO_75 (O_75,N_9654,N_9083);
nand UO_76 (O_76,N_9251,N_9226);
nor UO_77 (O_77,N_9375,N_9831);
xor UO_78 (O_78,N_9829,N_9305);
nor UO_79 (O_79,N_9052,N_9244);
and UO_80 (O_80,N_9367,N_9440);
and UO_81 (O_81,N_9465,N_9368);
and UO_82 (O_82,N_9960,N_9099);
nor UO_83 (O_83,N_9882,N_9452);
nand UO_84 (O_84,N_9778,N_9292);
or UO_85 (O_85,N_9723,N_9258);
nor UO_86 (O_86,N_9186,N_9825);
nor UO_87 (O_87,N_9053,N_9369);
or UO_88 (O_88,N_9227,N_9232);
and UO_89 (O_89,N_9697,N_9608);
or UO_90 (O_90,N_9837,N_9250);
and UO_91 (O_91,N_9365,N_9621);
nor UO_92 (O_92,N_9312,N_9140);
nand UO_93 (O_93,N_9596,N_9895);
and UO_94 (O_94,N_9085,N_9520);
and UO_95 (O_95,N_9660,N_9834);
or UO_96 (O_96,N_9230,N_9387);
nand UO_97 (O_97,N_9903,N_9537);
or UO_98 (O_98,N_9639,N_9436);
and UO_99 (O_99,N_9714,N_9300);
and UO_100 (O_100,N_9838,N_9277);
nor UO_101 (O_101,N_9701,N_9281);
nor UO_102 (O_102,N_9081,N_9731);
xor UO_103 (O_103,N_9027,N_9306);
nor UO_104 (O_104,N_9468,N_9299);
or UO_105 (O_105,N_9845,N_9223);
nand UO_106 (O_106,N_9943,N_9160);
and UO_107 (O_107,N_9208,N_9587);
nand UO_108 (O_108,N_9781,N_9125);
or UO_109 (O_109,N_9844,N_9307);
nand UO_110 (O_110,N_9390,N_9994);
nor UO_111 (O_111,N_9646,N_9162);
or UO_112 (O_112,N_9717,N_9008);
nor UO_113 (O_113,N_9329,N_9944);
and UO_114 (O_114,N_9273,N_9377);
nor UO_115 (O_115,N_9650,N_9567);
nor UO_116 (O_116,N_9950,N_9320);
and UO_117 (O_117,N_9879,N_9221);
or UO_118 (O_118,N_9199,N_9764);
and UO_119 (O_119,N_9780,N_9864);
or UO_120 (O_120,N_9662,N_9466);
nor UO_121 (O_121,N_9557,N_9737);
nand UO_122 (O_122,N_9862,N_9510);
nor UO_123 (O_123,N_9088,N_9519);
and UO_124 (O_124,N_9473,N_9127);
and UO_125 (O_125,N_9610,N_9946);
or UO_126 (O_126,N_9455,N_9351);
nor UO_127 (O_127,N_9751,N_9642);
nor UO_128 (O_128,N_9795,N_9655);
or UO_129 (O_129,N_9640,N_9184);
xor UO_130 (O_130,N_9006,N_9763);
or UO_131 (O_131,N_9747,N_9285);
nand UO_132 (O_132,N_9932,N_9700);
nor UO_133 (O_133,N_9754,N_9420);
and UO_134 (O_134,N_9501,N_9527);
nor UO_135 (O_135,N_9123,N_9528);
nor UO_136 (O_136,N_9938,N_9869);
nor UO_137 (O_137,N_9021,N_9885);
or UO_138 (O_138,N_9989,N_9024);
nand UO_139 (O_139,N_9068,N_9934);
and UO_140 (O_140,N_9571,N_9964);
nand UO_141 (O_141,N_9134,N_9741);
or UO_142 (O_142,N_9046,N_9229);
and UO_143 (O_143,N_9463,N_9324);
nand UO_144 (O_144,N_9987,N_9530);
or UO_145 (O_145,N_9166,N_9043);
or UO_146 (O_146,N_9647,N_9454);
nor UO_147 (O_147,N_9756,N_9674);
nand UO_148 (O_148,N_9372,N_9347);
or UO_149 (O_149,N_9005,N_9034);
xnor UO_150 (O_150,N_9225,N_9937);
nor UO_151 (O_151,N_9693,N_9980);
or UO_152 (O_152,N_9595,N_9020);
nor UO_153 (O_153,N_9040,N_9710);
nand UO_154 (O_154,N_9426,N_9668);
and UO_155 (O_155,N_9597,N_9695);
and UO_156 (O_156,N_9531,N_9084);
and UO_157 (O_157,N_9237,N_9641);
or UO_158 (O_158,N_9614,N_9103);
nand UO_159 (O_159,N_9648,N_9067);
and UO_160 (O_160,N_9978,N_9178);
nor UO_161 (O_161,N_9378,N_9556);
nand UO_162 (O_162,N_9917,N_9211);
and UO_163 (O_163,N_9181,N_9164);
and UO_164 (O_164,N_9746,N_9512);
or UO_165 (O_165,N_9889,N_9354);
nor UO_166 (O_166,N_9490,N_9849);
nor UO_167 (O_167,N_9197,N_9884);
nor UO_168 (O_168,N_9026,N_9586);
nor UO_169 (O_169,N_9146,N_9991);
and UO_170 (O_170,N_9965,N_9986);
xor UO_171 (O_171,N_9999,N_9868);
and UO_172 (O_172,N_9827,N_9193);
and UO_173 (O_173,N_9985,N_9604);
or UO_174 (O_174,N_9011,N_9359);
and UO_175 (O_175,N_9673,N_9979);
nand UO_176 (O_176,N_9079,N_9035);
or UO_177 (O_177,N_9196,N_9657);
nand UO_178 (O_178,N_9524,N_9357);
or UO_179 (O_179,N_9771,N_9928);
or UO_180 (O_180,N_9638,N_9102);
nor UO_181 (O_181,N_9607,N_9952);
and UO_182 (O_182,N_9425,N_9464);
or UO_183 (O_183,N_9798,N_9002);
nor UO_184 (O_184,N_9228,N_9248);
and UO_185 (O_185,N_9543,N_9832);
and UO_186 (O_186,N_9593,N_9899);
and UO_187 (O_187,N_9442,N_9126);
nand UO_188 (O_188,N_9704,N_9896);
and UO_189 (O_189,N_9522,N_9730);
nand UO_190 (O_190,N_9031,N_9508);
and UO_191 (O_191,N_9765,N_9157);
and UO_192 (O_192,N_9113,N_9396);
and UO_193 (O_193,N_9456,N_9328);
or UO_194 (O_194,N_9955,N_9149);
nor UO_195 (O_195,N_9176,N_9222);
xnor UO_196 (O_196,N_9152,N_9677);
nor UO_197 (O_197,N_9552,N_9267);
xor UO_198 (O_198,N_9201,N_9833);
xnor UO_199 (O_199,N_9439,N_9653);
xnor UO_200 (O_200,N_9424,N_9785);
nor UO_201 (O_201,N_9828,N_9860);
nand UO_202 (O_202,N_9290,N_9268);
or UO_203 (O_203,N_9971,N_9988);
nand UO_204 (O_204,N_9993,N_9616);
nand UO_205 (O_205,N_9951,N_9432);
or UO_206 (O_206,N_9494,N_9821);
nor UO_207 (O_207,N_9169,N_9269);
nor UO_208 (O_208,N_9259,N_9066);
or UO_209 (O_209,N_9167,N_9956);
nand UO_210 (O_210,N_9385,N_9625);
and UO_211 (O_211,N_9075,N_9574);
nand UO_212 (O_212,N_9939,N_9138);
nor UO_213 (O_213,N_9664,N_9634);
and UO_214 (O_214,N_9009,N_9190);
nor UO_215 (O_215,N_9548,N_9460);
and UO_216 (O_216,N_9620,N_9478);
nand UO_217 (O_217,N_9973,N_9911);
nand UO_218 (O_218,N_9119,N_9914);
nor UO_219 (O_219,N_9846,N_9509);
or UO_220 (O_220,N_9893,N_9722);
nand UO_221 (O_221,N_9841,N_9289);
or UO_222 (O_222,N_9724,N_9395);
and UO_223 (O_223,N_9403,N_9386);
or UO_224 (O_224,N_9245,N_9263);
and UO_225 (O_225,N_9297,N_9533);
and UO_226 (O_226,N_9093,N_9743);
and UO_227 (O_227,N_9851,N_9716);
nor UO_228 (O_228,N_9037,N_9505);
nor UO_229 (O_229,N_9738,N_9405);
nor UO_230 (O_230,N_9438,N_9957);
nand UO_231 (O_231,N_9847,N_9483);
and UO_232 (O_232,N_9203,N_9753);
nand UO_233 (O_233,N_9360,N_9394);
nor UO_234 (O_234,N_9000,N_9810);
nand UO_235 (O_235,N_9298,N_9142);
nand UO_236 (O_236,N_9959,N_9603);
nand UO_237 (O_237,N_9130,N_9694);
xnor UO_238 (O_238,N_9811,N_9388);
and UO_239 (O_239,N_9481,N_9699);
nor UO_240 (O_240,N_9760,N_9352);
nand UO_241 (O_241,N_9295,N_9333);
nor UO_242 (O_242,N_9412,N_9807);
nor UO_243 (O_243,N_9995,N_9949);
and UO_244 (O_244,N_9309,N_9872);
or UO_245 (O_245,N_9282,N_9393);
nand UO_246 (O_246,N_9252,N_9974);
or UO_247 (O_247,N_9692,N_9990);
and UO_248 (O_248,N_9559,N_9023);
and UO_249 (O_249,N_9739,N_9815);
and UO_250 (O_250,N_9861,N_9380);
nor UO_251 (O_251,N_9376,N_9332);
and UO_252 (O_252,N_9476,N_9437);
nand UO_253 (O_253,N_9496,N_9317);
or UO_254 (O_254,N_9391,N_9361);
and UO_255 (O_255,N_9547,N_9110);
or UO_256 (O_256,N_9217,N_9562);
nand UO_257 (O_257,N_9057,N_9658);
or UO_258 (O_258,N_9766,N_9526);
nor UO_259 (O_259,N_9215,N_9534);
and UO_260 (O_260,N_9392,N_9015);
nand UO_261 (O_261,N_9843,N_9630);
nand UO_262 (O_262,N_9240,N_9086);
nand UO_263 (O_263,N_9247,N_9507);
nor UO_264 (O_264,N_9584,N_9576);
xor UO_265 (O_265,N_9294,N_9205);
nor UO_266 (O_266,N_9623,N_9968);
xnor UO_267 (O_267,N_9892,N_9171);
and UO_268 (O_268,N_9656,N_9062);
and UO_269 (O_269,N_9012,N_9283);
nor UO_270 (O_270,N_9865,N_9177);
nand UO_271 (O_271,N_9789,N_9491);
xor UO_272 (O_272,N_9794,N_9613);
or UO_273 (O_273,N_9824,N_9118);
and UO_274 (O_274,N_9803,N_9279);
nand UO_275 (O_275,N_9898,N_9477);
nand UO_276 (O_276,N_9812,N_9049);
or UO_277 (O_277,N_9314,N_9560);
nand UO_278 (O_278,N_9930,N_9063);
nand UO_279 (O_279,N_9792,N_9583);
or UO_280 (O_280,N_9523,N_9136);
and UO_281 (O_281,N_9449,N_9271);
or UO_282 (O_282,N_9967,N_9143);
nor UO_283 (O_283,N_9629,N_9611);
nand UO_284 (O_284,N_9356,N_9626);
nand UO_285 (O_285,N_9089,N_9475);
and UO_286 (O_286,N_9728,N_9935);
and UO_287 (O_287,N_9092,N_9200);
nand UO_288 (O_288,N_9686,N_9408);
nor UO_289 (O_289,N_9249,N_9925);
or UO_290 (O_290,N_9786,N_9101);
nor UO_291 (O_291,N_9304,N_9669);
nand UO_292 (O_292,N_9667,N_9242);
nor UO_293 (O_293,N_9253,N_9707);
nor UO_294 (O_294,N_9170,N_9735);
nand UO_295 (O_295,N_9095,N_9411);
and UO_296 (O_296,N_9071,N_9514);
nand UO_297 (O_297,N_9788,N_9106);
nor UO_298 (O_298,N_9876,N_9998);
and UO_299 (O_299,N_9518,N_9546);
or UO_300 (O_300,N_9047,N_9622);
and UO_301 (O_301,N_9310,N_9906);
nor UO_302 (O_302,N_9549,N_9787);
and UO_303 (O_303,N_9718,N_9880);
nand UO_304 (O_304,N_9080,N_9382);
nor UO_305 (O_305,N_9705,N_9690);
nand UO_306 (O_306,N_9888,N_9826);
nand UO_307 (O_307,N_9588,N_9185);
and UO_308 (O_308,N_9050,N_9891);
nor UO_309 (O_309,N_9539,N_9308);
or UO_310 (O_310,N_9680,N_9450);
and UO_311 (O_311,N_9924,N_9545);
nand UO_312 (O_312,N_9335,N_9688);
or UO_313 (O_313,N_9238,N_9983);
nand UO_314 (O_314,N_9804,N_9497);
xnor UO_315 (O_315,N_9814,N_9783);
or UO_316 (O_316,N_9105,N_9076);
or UO_317 (O_317,N_9159,N_9682);
nand UO_318 (O_318,N_9137,N_9330);
nand UO_319 (O_319,N_9725,N_9209);
and UO_320 (O_320,N_9077,N_9691);
xor UO_321 (O_321,N_9516,N_9996);
nor UO_322 (O_322,N_9819,N_9782);
nand UO_323 (O_323,N_9897,N_9358);
or UO_324 (O_324,N_9768,N_9260);
and UO_325 (O_325,N_9192,N_9078);
or UO_326 (O_326,N_9774,N_9044);
nor UO_327 (O_327,N_9577,N_9434);
or UO_328 (O_328,N_9082,N_9401);
nand UO_329 (O_329,N_9767,N_9636);
xnor UO_330 (O_330,N_9721,N_9820);
nand UO_331 (O_331,N_9471,N_9744);
or UO_332 (O_332,N_9028,N_9073);
and UO_333 (O_333,N_9536,N_9503);
nor UO_334 (O_334,N_9762,N_9958);
or UO_335 (O_335,N_9492,N_9441);
nor UO_336 (O_336,N_9661,N_9652);
and UO_337 (O_337,N_9316,N_9823);
nor UO_338 (O_338,N_9858,N_9370);
nor UO_339 (O_339,N_9343,N_9580);
xnor UO_340 (O_340,N_9644,N_9506);
nor UO_341 (O_341,N_9670,N_9064);
nor UO_342 (O_342,N_9342,N_9649);
nor UO_343 (O_343,N_9554,N_9561);
or UO_344 (O_344,N_9659,N_9121);
or UO_345 (O_345,N_9916,N_9555);
and UO_346 (O_346,N_9541,N_9270);
or UO_347 (O_347,N_9665,N_9748);
nand UO_348 (O_348,N_9904,N_9915);
nor UO_349 (O_349,N_9276,N_9696);
xnor UO_350 (O_350,N_9341,N_9498);
nand UO_351 (O_351,N_9141,N_9224);
nor UO_352 (O_352,N_9840,N_9961);
nor UO_353 (O_353,N_9019,N_9755);
and UO_354 (O_354,N_9881,N_9901);
xor UO_355 (O_355,N_9430,N_9213);
nor UO_356 (O_356,N_9091,N_9427);
or UO_357 (O_357,N_9633,N_9419);
and UO_358 (O_358,N_9761,N_9902);
nor UO_359 (O_359,N_9480,N_9029);
or UO_360 (O_360,N_9627,N_9488);
or UO_361 (O_361,N_9416,N_9060);
nand UO_362 (O_362,N_9502,N_9384);
or UO_363 (O_363,N_9349,N_9133);
or UO_364 (O_364,N_9318,N_9262);
nor UO_365 (O_365,N_9214,N_9275);
or UO_366 (O_366,N_9525,N_9397);
and UO_367 (O_367,N_9218,N_9606);
nand UO_368 (O_368,N_9338,N_9521);
nand UO_369 (O_369,N_9806,N_9041);
nand UO_370 (O_370,N_9163,N_9234);
or UO_371 (O_371,N_9617,N_9890);
and UO_372 (O_372,N_9389,N_9926);
nand UO_373 (O_373,N_9096,N_9719);
and UO_374 (O_374,N_9605,N_9982);
and UO_375 (O_375,N_9830,N_9817);
nor UO_376 (O_376,N_9151,N_9115);
nor UO_377 (O_377,N_9479,N_9848);
and UO_378 (O_378,N_9147,N_9274);
nand UO_379 (O_379,N_9188,N_9261);
xor UO_380 (O_380,N_9045,N_9619);
or UO_381 (O_381,N_9493,N_9153);
and UO_382 (O_382,N_9791,N_9286);
nand UO_383 (O_383,N_9905,N_9189);
nand UO_384 (O_384,N_9687,N_9883);
and UO_385 (O_385,N_9553,N_9435);
and UO_386 (O_386,N_9323,N_9069);
and UO_387 (O_387,N_9474,N_9966);
or UO_388 (O_388,N_9676,N_9236);
or UO_389 (O_389,N_9120,N_9504);
nand UO_390 (O_390,N_9550,N_9409);
nand UO_391 (O_391,N_9104,N_9265);
nor UO_392 (O_392,N_9931,N_9535);
nor UO_393 (O_393,N_9663,N_9540);
and UO_394 (O_394,N_9948,N_9364);
nand UO_395 (O_395,N_9210,N_9570);
xnor UO_396 (O_396,N_9489,N_9017);
or UO_397 (O_397,N_9855,N_9128);
nor UO_398 (O_398,N_9168,N_9809);
nand UO_399 (O_399,N_9220,N_9870);
nand UO_400 (O_400,N_9231,N_9195);
and UO_401 (O_401,N_9004,N_9111);
and UO_402 (O_402,N_9287,N_9255);
nor UO_403 (O_403,N_9433,N_9183);
nor UO_404 (O_404,N_9487,N_9628);
nor UO_405 (O_405,N_9566,N_9331);
nand UO_406 (O_406,N_9805,N_9565);
nor UO_407 (O_407,N_9032,N_9451);
or UO_408 (O_408,N_9233,N_9759);
and UO_409 (O_409,N_9871,N_9757);
or UO_410 (O_410,N_9165,N_9191);
nor UO_411 (O_411,N_9072,N_9467);
and UO_412 (O_412,N_9706,N_9402);
nand UO_413 (O_413,N_9581,N_9303);
nor UO_414 (O_414,N_9212,N_9857);
or UO_415 (O_415,N_9344,N_9156);
and UO_416 (O_416,N_9484,N_9500);
and UO_417 (O_417,N_9462,N_9180);
nand UO_418 (O_418,N_9708,N_9366);
xor UO_419 (O_419,N_9038,N_9643);
nand UO_420 (O_420,N_9866,N_9486);
or UO_421 (O_421,N_9594,N_9802);
xnor UO_422 (O_422,N_9198,N_9779);
nor UO_423 (O_423,N_9499,N_9977);
xor UO_424 (O_424,N_9321,N_9726);
or UO_425 (O_425,N_9381,N_9407);
and UO_426 (O_426,N_9969,N_9246);
and UO_427 (O_427,N_9039,N_9139);
nor UO_428 (O_428,N_9334,N_9112);
nor UO_429 (O_429,N_9513,N_9175);
or UO_430 (O_430,N_9059,N_9150);
nand UO_431 (O_431,N_9194,N_9301);
nor UO_432 (O_432,N_9322,N_9936);
nor UO_433 (O_433,N_9172,N_9348);
nand UO_434 (O_434,N_9910,N_9336);
and UO_435 (O_435,N_9291,N_9850);
or UO_436 (O_436,N_9671,N_9777);
nand UO_437 (O_437,N_9161,N_9458);
and UO_438 (O_438,N_9054,N_9042);
nand UO_439 (O_439,N_9529,N_9919);
or UO_440 (O_440,N_9874,N_9772);
and UO_441 (O_441,N_9087,N_9206);
xor UO_442 (O_442,N_9790,N_9972);
and UO_443 (O_443,N_9563,N_9241);
or UO_444 (O_444,N_9148,N_9051);
nand UO_445 (O_445,N_9736,N_9373);
or UO_446 (O_446,N_9313,N_9544);
and UO_447 (O_447,N_9784,N_9485);
nand UO_448 (O_448,N_9750,N_9900);
and UO_449 (O_449,N_9302,N_9446);
nor UO_450 (O_450,N_9578,N_9003);
or UO_451 (O_451,N_9532,N_9431);
nand UO_452 (O_452,N_9254,N_9070);
nor UO_453 (O_453,N_9681,N_9635);
or UO_454 (O_454,N_9418,N_9417);
and UO_455 (O_455,N_9448,N_9272);
nand UO_456 (O_456,N_9927,N_9399);
xnor UO_457 (O_457,N_9679,N_9796);
or UO_458 (O_458,N_9573,N_9918);
nand UO_459 (O_459,N_9428,N_9108);
or UO_460 (O_460,N_9923,N_9122);
and UO_461 (O_461,N_9773,N_9867);
and UO_462 (O_462,N_9572,N_9801);
or UO_463 (O_463,N_9144,N_9818);
and UO_464 (O_464,N_9470,N_9976);
nand UO_465 (O_465,N_9793,N_9887);
nand UO_466 (O_466,N_9836,N_9551);
nand UO_467 (O_467,N_9055,N_9415);
nand UO_468 (O_468,N_9745,N_9909);
nor UO_469 (O_469,N_9997,N_9954);
or UO_470 (O_470,N_9609,N_9683);
or UO_471 (O_471,N_9319,N_9666);
nor UO_472 (O_472,N_9922,N_9266);
nand UO_473 (O_473,N_9689,N_9875);
xnor UO_474 (O_474,N_9645,N_9715);
or UO_475 (O_475,N_9117,N_9459);
and UO_476 (O_476,N_9444,N_9942);
nor UO_477 (O_477,N_9056,N_9913);
or UO_478 (O_478,N_9097,N_9013);
nand UO_479 (O_479,N_9953,N_9564);
or UO_480 (O_480,N_9061,N_9631);
nand UO_481 (O_481,N_9585,N_9065);
nand UO_482 (O_482,N_9443,N_9100);
nor UO_483 (O_483,N_9685,N_9311);
nor UO_484 (O_484,N_9612,N_9132);
nor UO_485 (O_485,N_9182,N_9835);
nand UO_486 (O_486,N_9179,N_9422);
nand UO_487 (O_487,N_9775,N_9379);
nor UO_488 (O_488,N_9406,N_9729);
nand UO_489 (O_489,N_9981,N_9615);
nand UO_490 (O_490,N_9992,N_9469);
nor UO_491 (O_491,N_9280,N_9030);
or UO_492 (O_492,N_9886,N_9414);
and UO_493 (O_493,N_9592,N_9776);
and UO_494 (O_494,N_9542,N_9374);
nand UO_495 (O_495,N_9410,N_9770);
nor UO_496 (O_496,N_9734,N_9598);
and UO_497 (O_497,N_9856,N_9515);
nor UO_498 (O_498,N_9155,N_9853);
nor UO_499 (O_499,N_9599,N_9538);
and UO_500 (O_500,N_9006,N_9514);
and UO_501 (O_501,N_9144,N_9329);
or UO_502 (O_502,N_9150,N_9577);
and UO_503 (O_503,N_9894,N_9748);
nand UO_504 (O_504,N_9508,N_9493);
and UO_505 (O_505,N_9966,N_9494);
or UO_506 (O_506,N_9706,N_9507);
nand UO_507 (O_507,N_9847,N_9871);
nor UO_508 (O_508,N_9536,N_9824);
or UO_509 (O_509,N_9737,N_9179);
or UO_510 (O_510,N_9446,N_9905);
and UO_511 (O_511,N_9795,N_9108);
and UO_512 (O_512,N_9059,N_9840);
xnor UO_513 (O_513,N_9201,N_9223);
nand UO_514 (O_514,N_9867,N_9078);
xor UO_515 (O_515,N_9859,N_9647);
nor UO_516 (O_516,N_9447,N_9214);
nor UO_517 (O_517,N_9700,N_9676);
nor UO_518 (O_518,N_9156,N_9905);
nor UO_519 (O_519,N_9935,N_9943);
and UO_520 (O_520,N_9329,N_9504);
and UO_521 (O_521,N_9456,N_9109);
or UO_522 (O_522,N_9645,N_9983);
nand UO_523 (O_523,N_9377,N_9740);
nand UO_524 (O_524,N_9111,N_9622);
nand UO_525 (O_525,N_9500,N_9726);
and UO_526 (O_526,N_9474,N_9375);
and UO_527 (O_527,N_9536,N_9890);
xor UO_528 (O_528,N_9459,N_9986);
and UO_529 (O_529,N_9915,N_9107);
nand UO_530 (O_530,N_9475,N_9639);
nor UO_531 (O_531,N_9206,N_9068);
xnor UO_532 (O_532,N_9374,N_9040);
nor UO_533 (O_533,N_9086,N_9991);
nor UO_534 (O_534,N_9593,N_9349);
nor UO_535 (O_535,N_9082,N_9098);
nor UO_536 (O_536,N_9775,N_9599);
nand UO_537 (O_537,N_9828,N_9835);
xor UO_538 (O_538,N_9500,N_9793);
and UO_539 (O_539,N_9366,N_9672);
nor UO_540 (O_540,N_9909,N_9974);
nor UO_541 (O_541,N_9412,N_9257);
or UO_542 (O_542,N_9498,N_9565);
xor UO_543 (O_543,N_9328,N_9976);
nand UO_544 (O_544,N_9029,N_9114);
xor UO_545 (O_545,N_9568,N_9108);
nand UO_546 (O_546,N_9349,N_9898);
and UO_547 (O_547,N_9718,N_9365);
or UO_548 (O_548,N_9680,N_9479);
and UO_549 (O_549,N_9939,N_9701);
xor UO_550 (O_550,N_9827,N_9680);
nor UO_551 (O_551,N_9370,N_9685);
nand UO_552 (O_552,N_9287,N_9852);
and UO_553 (O_553,N_9024,N_9542);
nand UO_554 (O_554,N_9857,N_9529);
or UO_555 (O_555,N_9770,N_9209);
or UO_556 (O_556,N_9565,N_9643);
or UO_557 (O_557,N_9341,N_9032);
nor UO_558 (O_558,N_9015,N_9776);
or UO_559 (O_559,N_9155,N_9612);
or UO_560 (O_560,N_9105,N_9092);
nand UO_561 (O_561,N_9531,N_9384);
nor UO_562 (O_562,N_9431,N_9023);
and UO_563 (O_563,N_9457,N_9594);
or UO_564 (O_564,N_9575,N_9104);
or UO_565 (O_565,N_9390,N_9801);
and UO_566 (O_566,N_9437,N_9222);
and UO_567 (O_567,N_9341,N_9810);
nor UO_568 (O_568,N_9693,N_9566);
nand UO_569 (O_569,N_9621,N_9591);
or UO_570 (O_570,N_9753,N_9233);
nor UO_571 (O_571,N_9915,N_9594);
and UO_572 (O_572,N_9923,N_9207);
nand UO_573 (O_573,N_9120,N_9203);
nand UO_574 (O_574,N_9231,N_9379);
xor UO_575 (O_575,N_9559,N_9259);
nor UO_576 (O_576,N_9290,N_9800);
nand UO_577 (O_577,N_9199,N_9169);
or UO_578 (O_578,N_9695,N_9191);
xnor UO_579 (O_579,N_9633,N_9854);
nand UO_580 (O_580,N_9099,N_9893);
nand UO_581 (O_581,N_9946,N_9042);
nand UO_582 (O_582,N_9768,N_9393);
or UO_583 (O_583,N_9680,N_9743);
xnor UO_584 (O_584,N_9926,N_9746);
or UO_585 (O_585,N_9754,N_9102);
nor UO_586 (O_586,N_9244,N_9845);
or UO_587 (O_587,N_9413,N_9788);
nor UO_588 (O_588,N_9786,N_9459);
and UO_589 (O_589,N_9098,N_9185);
nand UO_590 (O_590,N_9983,N_9689);
and UO_591 (O_591,N_9109,N_9669);
xor UO_592 (O_592,N_9358,N_9266);
and UO_593 (O_593,N_9012,N_9179);
nor UO_594 (O_594,N_9002,N_9851);
nor UO_595 (O_595,N_9402,N_9453);
nand UO_596 (O_596,N_9498,N_9406);
xnor UO_597 (O_597,N_9396,N_9760);
nand UO_598 (O_598,N_9552,N_9981);
and UO_599 (O_599,N_9347,N_9856);
nand UO_600 (O_600,N_9047,N_9452);
xor UO_601 (O_601,N_9706,N_9958);
nand UO_602 (O_602,N_9515,N_9028);
and UO_603 (O_603,N_9832,N_9890);
nand UO_604 (O_604,N_9840,N_9063);
and UO_605 (O_605,N_9563,N_9858);
and UO_606 (O_606,N_9306,N_9443);
nor UO_607 (O_607,N_9217,N_9693);
or UO_608 (O_608,N_9185,N_9900);
or UO_609 (O_609,N_9670,N_9079);
or UO_610 (O_610,N_9504,N_9436);
or UO_611 (O_611,N_9286,N_9016);
nor UO_612 (O_612,N_9951,N_9777);
and UO_613 (O_613,N_9674,N_9115);
or UO_614 (O_614,N_9761,N_9917);
and UO_615 (O_615,N_9311,N_9244);
nand UO_616 (O_616,N_9311,N_9133);
nand UO_617 (O_617,N_9028,N_9117);
nand UO_618 (O_618,N_9642,N_9082);
xnor UO_619 (O_619,N_9851,N_9807);
nand UO_620 (O_620,N_9445,N_9348);
and UO_621 (O_621,N_9332,N_9414);
nand UO_622 (O_622,N_9135,N_9346);
nor UO_623 (O_623,N_9037,N_9619);
and UO_624 (O_624,N_9285,N_9339);
nor UO_625 (O_625,N_9946,N_9435);
nand UO_626 (O_626,N_9305,N_9964);
nor UO_627 (O_627,N_9752,N_9536);
nor UO_628 (O_628,N_9993,N_9842);
nor UO_629 (O_629,N_9446,N_9554);
nor UO_630 (O_630,N_9198,N_9919);
xor UO_631 (O_631,N_9587,N_9064);
or UO_632 (O_632,N_9308,N_9576);
and UO_633 (O_633,N_9591,N_9764);
nor UO_634 (O_634,N_9381,N_9852);
or UO_635 (O_635,N_9379,N_9346);
or UO_636 (O_636,N_9169,N_9790);
or UO_637 (O_637,N_9263,N_9469);
or UO_638 (O_638,N_9670,N_9236);
or UO_639 (O_639,N_9797,N_9319);
and UO_640 (O_640,N_9578,N_9690);
and UO_641 (O_641,N_9187,N_9542);
nor UO_642 (O_642,N_9012,N_9466);
or UO_643 (O_643,N_9156,N_9533);
nand UO_644 (O_644,N_9032,N_9749);
and UO_645 (O_645,N_9662,N_9058);
nor UO_646 (O_646,N_9523,N_9498);
nor UO_647 (O_647,N_9759,N_9338);
nand UO_648 (O_648,N_9397,N_9752);
nor UO_649 (O_649,N_9989,N_9975);
nand UO_650 (O_650,N_9605,N_9518);
nor UO_651 (O_651,N_9814,N_9465);
nand UO_652 (O_652,N_9399,N_9482);
or UO_653 (O_653,N_9994,N_9929);
nor UO_654 (O_654,N_9603,N_9619);
and UO_655 (O_655,N_9449,N_9915);
nand UO_656 (O_656,N_9592,N_9841);
or UO_657 (O_657,N_9850,N_9023);
nor UO_658 (O_658,N_9588,N_9825);
nor UO_659 (O_659,N_9432,N_9912);
nor UO_660 (O_660,N_9046,N_9324);
and UO_661 (O_661,N_9326,N_9562);
nand UO_662 (O_662,N_9552,N_9471);
or UO_663 (O_663,N_9920,N_9560);
nor UO_664 (O_664,N_9292,N_9386);
or UO_665 (O_665,N_9415,N_9459);
and UO_666 (O_666,N_9794,N_9623);
or UO_667 (O_667,N_9181,N_9160);
xor UO_668 (O_668,N_9896,N_9594);
and UO_669 (O_669,N_9401,N_9739);
or UO_670 (O_670,N_9322,N_9604);
nor UO_671 (O_671,N_9179,N_9380);
nor UO_672 (O_672,N_9730,N_9221);
nor UO_673 (O_673,N_9128,N_9705);
nor UO_674 (O_674,N_9291,N_9191);
nor UO_675 (O_675,N_9701,N_9097);
and UO_676 (O_676,N_9278,N_9909);
nand UO_677 (O_677,N_9733,N_9244);
nor UO_678 (O_678,N_9791,N_9098);
nor UO_679 (O_679,N_9858,N_9416);
or UO_680 (O_680,N_9876,N_9292);
or UO_681 (O_681,N_9658,N_9562);
and UO_682 (O_682,N_9203,N_9767);
nor UO_683 (O_683,N_9119,N_9630);
xor UO_684 (O_684,N_9837,N_9818);
xor UO_685 (O_685,N_9127,N_9074);
or UO_686 (O_686,N_9773,N_9156);
nor UO_687 (O_687,N_9122,N_9511);
nand UO_688 (O_688,N_9735,N_9838);
and UO_689 (O_689,N_9732,N_9665);
and UO_690 (O_690,N_9236,N_9313);
nand UO_691 (O_691,N_9148,N_9890);
nand UO_692 (O_692,N_9975,N_9885);
xnor UO_693 (O_693,N_9191,N_9985);
nor UO_694 (O_694,N_9353,N_9491);
and UO_695 (O_695,N_9203,N_9555);
or UO_696 (O_696,N_9581,N_9918);
and UO_697 (O_697,N_9508,N_9339);
nor UO_698 (O_698,N_9181,N_9021);
nor UO_699 (O_699,N_9472,N_9103);
or UO_700 (O_700,N_9105,N_9999);
nor UO_701 (O_701,N_9639,N_9066);
or UO_702 (O_702,N_9856,N_9404);
nand UO_703 (O_703,N_9227,N_9824);
nand UO_704 (O_704,N_9493,N_9813);
and UO_705 (O_705,N_9494,N_9552);
and UO_706 (O_706,N_9124,N_9354);
and UO_707 (O_707,N_9768,N_9595);
nor UO_708 (O_708,N_9154,N_9366);
nor UO_709 (O_709,N_9681,N_9690);
nand UO_710 (O_710,N_9918,N_9360);
nand UO_711 (O_711,N_9954,N_9828);
nor UO_712 (O_712,N_9902,N_9922);
and UO_713 (O_713,N_9656,N_9699);
nand UO_714 (O_714,N_9607,N_9782);
and UO_715 (O_715,N_9672,N_9843);
or UO_716 (O_716,N_9178,N_9880);
nor UO_717 (O_717,N_9069,N_9096);
or UO_718 (O_718,N_9695,N_9864);
nor UO_719 (O_719,N_9218,N_9280);
and UO_720 (O_720,N_9800,N_9622);
nor UO_721 (O_721,N_9056,N_9409);
nand UO_722 (O_722,N_9692,N_9396);
or UO_723 (O_723,N_9447,N_9585);
and UO_724 (O_724,N_9865,N_9634);
or UO_725 (O_725,N_9478,N_9552);
or UO_726 (O_726,N_9876,N_9651);
xor UO_727 (O_727,N_9010,N_9522);
nand UO_728 (O_728,N_9123,N_9207);
nor UO_729 (O_729,N_9247,N_9552);
nor UO_730 (O_730,N_9222,N_9866);
nand UO_731 (O_731,N_9642,N_9793);
or UO_732 (O_732,N_9244,N_9044);
nor UO_733 (O_733,N_9376,N_9237);
and UO_734 (O_734,N_9521,N_9093);
nor UO_735 (O_735,N_9956,N_9323);
nand UO_736 (O_736,N_9276,N_9653);
nand UO_737 (O_737,N_9014,N_9371);
nor UO_738 (O_738,N_9903,N_9327);
and UO_739 (O_739,N_9278,N_9950);
nand UO_740 (O_740,N_9266,N_9708);
and UO_741 (O_741,N_9228,N_9731);
nor UO_742 (O_742,N_9082,N_9281);
and UO_743 (O_743,N_9913,N_9052);
nand UO_744 (O_744,N_9793,N_9874);
nand UO_745 (O_745,N_9904,N_9890);
or UO_746 (O_746,N_9505,N_9412);
or UO_747 (O_747,N_9201,N_9876);
nand UO_748 (O_748,N_9695,N_9520);
nor UO_749 (O_749,N_9714,N_9978);
nand UO_750 (O_750,N_9111,N_9600);
and UO_751 (O_751,N_9287,N_9384);
nand UO_752 (O_752,N_9811,N_9422);
or UO_753 (O_753,N_9575,N_9882);
and UO_754 (O_754,N_9480,N_9673);
nand UO_755 (O_755,N_9239,N_9336);
nand UO_756 (O_756,N_9157,N_9821);
nor UO_757 (O_757,N_9993,N_9662);
or UO_758 (O_758,N_9159,N_9703);
nand UO_759 (O_759,N_9420,N_9646);
and UO_760 (O_760,N_9358,N_9189);
and UO_761 (O_761,N_9790,N_9281);
xor UO_762 (O_762,N_9671,N_9603);
nor UO_763 (O_763,N_9298,N_9107);
nand UO_764 (O_764,N_9163,N_9275);
nand UO_765 (O_765,N_9841,N_9565);
nand UO_766 (O_766,N_9958,N_9622);
nand UO_767 (O_767,N_9212,N_9795);
nand UO_768 (O_768,N_9618,N_9844);
nand UO_769 (O_769,N_9866,N_9376);
xnor UO_770 (O_770,N_9711,N_9124);
nor UO_771 (O_771,N_9084,N_9719);
or UO_772 (O_772,N_9553,N_9213);
or UO_773 (O_773,N_9717,N_9522);
and UO_774 (O_774,N_9275,N_9489);
or UO_775 (O_775,N_9438,N_9465);
or UO_776 (O_776,N_9735,N_9808);
nand UO_777 (O_777,N_9601,N_9730);
nand UO_778 (O_778,N_9194,N_9086);
and UO_779 (O_779,N_9360,N_9939);
nand UO_780 (O_780,N_9707,N_9609);
nor UO_781 (O_781,N_9055,N_9539);
or UO_782 (O_782,N_9896,N_9549);
nand UO_783 (O_783,N_9999,N_9349);
nand UO_784 (O_784,N_9043,N_9873);
or UO_785 (O_785,N_9876,N_9497);
and UO_786 (O_786,N_9912,N_9672);
nand UO_787 (O_787,N_9208,N_9138);
or UO_788 (O_788,N_9155,N_9778);
nand UO_789 (O_789,N_9847,N_9711);
and UO_790 (O_790,N_9559,N_9650);
or UO_791 (O_791,N_9573,N_9376);
xnor UO_792 (O_792,N_9829,N_9941);
and UO_793 (O_793,N_9193,N_9911);
nor UO_794 (O_794,N_9197,N_9653);
and UO_795 (O_795,N_9196,N_9251);
or UO_796 (O_796,N_9669,N_9931);
nand UO_797 (O_797,N_9645,N_9532);
nor UO_798 (O_798,N_9322,N_9392);
and UO_799 (O_799,N_9503,N_9098);
nor UO_800 (O_800,N_9450,N_9527);
nor UO_801 (O_801,N_9497,N_9811);
and UO_802 (O_802,N_9742,N_9864);
nor UO_803 (O_803,N_9292,N_9660);
nor UO_804 (O_804,N_9027,N_9217);
and UO_805 (O_805,N_9020,N_9699);
nand UO_806 (O_806,N_9777,N_9040);
nand UO_807 (O_807,N_9378,N_9520);
nand UO_808 (O_808,N_9087,N_9668);
and UO_809 (O_809,N_9771,N_9378);
xnor UO_810 (O_810,N_9691,N_9150);
or UO_811 (O_811,N_9333,N_9484);
nand UO_812 (O_812,N_9963,N_9572);
nor UO_813 (O_813,N_9414,N_9031);
or UO_814 (O_814,N_9639,N_9373);
nand UO_815 (O_815,N_9768,N_9163);
and UO_816 (O_816,N_9904,N_9491);
and UO_817 (O_817,N_9563,N_9952);
nor UO_818 (O_818,N_9265,N_9963);
nor UO_819 (O_819,N_9821,N_9984);
xor UO_820 (O_820,N_9280,N_9356);
and UO_821 (O_821,N_9393,N_9104);
nand UO_822 (O_822,N_9161,N_9499);
nor UO_823 (O_823,N_9686,N_9532);
and UO_824 (O_824,N_9745,N_9375);
and UO_825 (O_825,N_9841,N_9149);
or UO_826 (O_826,N_9119,N_9790);
nor UO_827 (O_827,N_9173,N_9529);
and UO_828 (O_828,N_9994,N_9818);
xor UO_829 (O_829,N_9141,N_9872);
nor UO_830 (O_830,N_9022,N_9554);
nor UO_831 (O_831,N_9048,N_9942);
nand UO_832 (O_832,N_9352,N_9412);
or UO_833 (O_833,N_9934,N_9238);
or UO_834 (O_834,N_9517,N_9171);
or UO_835 (O_835,N_9909,N_9503);
or UO_836 (O_836,N_9562,N_9285);
or UO_837 (O_837,N_9256,N_9580);
and UO_838 (O_838,N_9538,N_9805);
and UO_839 (O_839,N_9134,N_9350);
nand UO_840 (O_840,N_9162,N_9464);
and UO_841 (O_841,N_9736,N_9124);
nor UO_842 (O_842,N_9568,N_9921);
and UO_843 (O_843,N_9778,N_9816);
or UO_844 (O_844,N_9404,N_9883);
nand UO_845 (O_845,N_9299,N_9977);
or UO_846 (O_846,N_9060,N_9511);
and UO_847 (O_847,N_9821,N_9760);
and UO_848 (O_848,N_9348,N_9995);
and UO_849 (O_849,N_9971,N_9788);
or UO_850 (O_850,N_9883,N_9616);
and UO_851 (O_851,N_9783,N_9107);
nand UO_852 (O_852,N_9727,N_9826);
nor UO_853 (O_853,N_9563,N_9628);
or UO_854 (O_854,N_9101,N_9402);
nand UO_855 (O_855,N_9768,N_9589);
nand UO_856 (O_856,N_9718,N_9389);
nor UO_857 (O_857,N_9204,N_9467);
or UO_858 (O_858,N_9219,N_9891);
nor UO_859 (O_859,N_9252,N_9511);
or UO_860 (O_860,N_9777,N_9908);
or UO_861 (O_861,N_9371,N_9468);
nor UO_862 (O_862,N_9798,N_9776);
or UO_863 (O_863,N_9181,N_9009);
nand UO_864 (O_864,N_9541,N_9794);
nand UO_865 (O_865,N_9356,N_9769);
nand UO_866 (O_866,N_9005,N_9941);
xnor UO_867 (O_867,N_9814,N_9935);
nand UO_868 (O_868,N_9206,N_9147);
nand UO_869 (O_869,N_9526,N_9239);
nor UO_870 (O_870,N_9660,N_9397);
and UO_871 (O_871,N_9501,N_9342);
or UO_872 (O_872,N_9705,N_9781);
nand UO_873 (O_873,N_9013,N_9528);
nor UO_874 (O_874,N_9410,N_9981);
nand UO_875 (O_875,N_9941,N_9967);
or UO_876 (O_876,N_9650,N_9414);
and UO_877 (O_877,N_9866,N_9933);
or UO_878 (O_878,N_9076,N_9182);
or UO_879 (O_879,N_9486,N_9327);
nand UO_880 (O_880,N_9051,N_9653);
nand UO_881 (O_881,N_9524,N_9144);
nand UO_882 (O_882,N_9438,N_9272);
and UO_883 (O_883,N_9906,N_9849);
nand UO_884 (O_884,N_9825,N_9865);
xnor UO_885 (O_885,N_9284,N_9781);
nor UO_886 (O_886,N_9838,N_9080);
nand UO_887 (O_887,N_9817,N_9321);
nand UO_888 (O_888,N_9736,N_9049);
and UO_889 (O_889,N_9515,N_9651);
nor UO_890 (O_890,N_9247,N_9123);
and UO_891 (O_891,N_9461,N_9108);
xor UO_892 (O_892,N_9526,N_9527);
nor UO_893 (O_893,N_9209,N_9037);
nor UO_894 (O_894,N_9991,N_9700);
and UO_895 (O_895,N_9734,N_9069);
or UO_896 (O_896,N_9916,N_9864);
xor UO_897 (O_897,N_9304,N_9985);
and UO_898 (O_898,N_9459,N_9355);
nand UO_899 (O_899,N_9642,N_9580);
or UO_900 (O_900,N_9468,N_9232);
or UO_901 (O_901,N_9362,N_9250);
xnor UO_902 (O_902,N_9456,N_9295);
or UO_903 (O_903,N_9546,N_9435);
nor UO_904 (O_904,N_9952,N_9608);
or UO_905 (O_905,N_9712,N_9832);
and UO_906 (O_906,N_9938,N_9410);
or UO_907 (O_907,N_9605,N_9409);
and UO_908 (O_908,N_9973,N_9512);
or UO_909 (O_909,N_9973,N_9754);
xor UO_910 (O_910,N_9169,N_9230);
nand UO_911 (O_911,N_9224,N_9104);
nor UO_912 (O_912,N_9576,N_9246);
and UO_913 (O_913,N_9055,N_9839);
and UO_914 (O_914,N_9683,N_9681);
nor UO_915 (O_915,N_9269,N_9540);
nand UO_916 (O_916,N_9100,N_9562);
xor UO_917 (O_917,N_9195,N_9130);
nand UO_918 (O_918,N_9701,N_9871);
nor UO_919 (O_919,N_9941,N_9550);
or UO_920 (O_920,N_9327,N_9113);
or UO_921 (O_921,N_9597,N_9036);
or UO_922 (O_922,N_9125,N_9829);
xnor UO_923 (O_923,N_9816,N_9110);
nor UO_924 (O_924,N_9855,N_9517);
nor UO_925 (O_925,N_9602,N_9818);
nor UO_926 (O_926,N_9651,N_9678);
xnor UO_927 (O_927,N_9783,N_9480);
nor UO_928 (O_928,N_9309,N_9359);
nand UO_929 (O_929,N_9425,N_9937);
xnor UO_930 (O_930,N_9086,N_9792);
or UO_931 (O_931,N_9701,N_9083);
and UO_932 (O_932,N_9457,N_9576);
nor UO_933 (O_933,N_9578,N_9903);
nand UO_934 (O_934,N_9859,N_9781);
nand UO_935 (O_935,N_9993,N_9259);
or UO_936 (O_936,N_9810,N_9945);
nor UO_937 (O_937,N_9782,N_9268);
nand UO_938 (O_938,N_9714,N_9998);
nand UO_939 (O_939,N_9671,N_9977);
and UO_940 (O_940,N_9852,N_9186);
nand UO_941 (O_941,N_9726,N_9064);
and UO_942 (O_942,N_9064,N_9951);
or UO_943 (O_943,N_9980,N_9138);
and UO_944 (O_944,N_9986,N_9319);
and UO_945 (O_945,N_9096,N_9651);
or UO_946 (O_946,N_9854,N_9737);
or UO_947 (O_947,N_9821,N_9435);
nand UO_948 (O_948,N_9988,N_9328);
and UO_949 (O_949,N_9564,N_9660);
or UO_950 (O_950,N_9429,N_9425);
nand UO_951 (O_951,N_9850,N_9880);
nor UO_952 (O_952,N_9061,N_9907);
or UO_953 (O_953,N_9802,N_9615);
nand UO_954 (O_954,N_9154,N_9615);
or UO_955 (O_955,N_9972,N_9919);
nand UO_956 (O_956,N_9107,N_9374);
nand UO_957 (O_957,N_9230,N_9398);
xor UO_958 (O_958,N_9105,N_9154);
or UO_959 (O_959,N_9009,N_9788);
nor UO_960 (O_960,N_9211,N_9289);
nor UO_961 (O_961,N_9873,N_9717);
and UO_962 (O_962,N_9455,N_9221);
nand UO_963 (O_963,N_9577,N_9423);
nor UO_964 (O_964,N_9768,N_9217);
and UO_965 (O_965,N_9315,N_9989);
xor UO_966 (O_966,N_9174,N_9122);
or UO_967 (O_967,N_9313,N_9655);
or UO_968 (O_968,N_9699,N_9175);
xor UO_969 (O_969,N_9215,N_9538);
nand UO_970 (O_970,N_9283,N_9629);
or UO_971 (O_971,N_9526,N_9929);
or UO_972 (O_972,N_9689,N_9249);
nor UO_973 (O_973,N_9021,N_9899);
nor UO_974 (O_974,N_9476,N_9351);
and UO_975 (O_975,N_9363,N_9234);
nor UO_976 (O_976,N_9212,N_9809);
or UO_977 (O_977,N_9663,N_9231);
and UO_978 (O_978,N_9180,N_9554);
or UO_979 (O_979,N_9679,N_9998);
and UO_980 (O_980,N_9289,N_9194);
or UO_981 (O_981,N_9071,N_9896);
and UO_982 (O_982,N_9278,N_9056);
nor UO_983 (O_983,N_9785,N_9463);
xor UO_984 (O_984,N_9861,N_9975);
nand UO_985 (O_985,N_9738,N_9205);
nor UO_986 (O_986,N_9947,N_9115);
and UO_987 (O_987,N_9889,N_9777);
and UO_988 (O_988,N_9722,N_9918);
nor UO_989 (O_989,N_9924,N_9630);
and UO_990 (O_990,N_9213,N_9046);
or UO_991 (O_991,N_9228,N_9178);
nand UO_992 (O_992,N_9522,N_9718);
nand UO_993 (O_993,N_9561,N_9132);
and UO_994 (O_994,N_9919,N_9024);
and UO_995 (O_995,N_9947,N_9413);
and UO_996 (O_996,N_9625,N_9443);
or UO_997 (O_997,N_9465,N_9304);
nand UO_998 (O_998,N_9874,N_9039);
and UO_999 (O_999,N_9470,N_9531);
or UO_1000 (O_1000,N_9690,N_9630);
xor UO_1001 (O_1001,N_9193,N_9498);
or UO_1002 (O_1002,N_9329,N_9773);
nor UO_1003 (O_1003,N_9624,N_9041);
nand UO_1004 (O_1004,N_9102,N_9923);
xor UO_1005 (O_1005,N_9558,N_9693);
nor UO_1006 (O_1006,N_9984,N_9721);
or UO_1007 (O_1007,N_9036,N_9505);
nor UO_1008 (O_1008,N_9305,N_9564);
nor UO_1009 (O_1009,N_9813,N_9009);
or UO_1010 (O_1010,N_9613,N_9110);
and UO_1011 (O_1011,N_9561,N_9743);
nand UO_1012 (O_1012,N_9107,N_9066);
nand UO_1013 (O_1013,N_9089,N_9808);
nand UO_1014 (O_1014,N_9360,N_9203);
nor UO_1015 (O_1015,N_9759,N_9358);
xnor UO_1016 (O_1016,N_9916,N_9638);
or UO_1017 (O_1017,N_9157,N_9225);
nand UO_1018 (O_1018,N_9816,N_9200);
and UO_1019 (O_1019,N_9898,N_9087);
or UO_1020 (O_1020,N_9805,N_9083);
or UO_1021 (O_1021,N_9346,N_9643);
nand UO_1022 (O_1022,N_9406,N_9262);
or UO_1023 (O_1023,N_9276,N_9735);
nor UO_1024 (O_1024,N_9551,N_9872);
xor UO_1025 (O_1025,N_9077,N_9748);
xor UO_1026 (O_1026,N_9217,N_9474);
or UO_1027 (O_1027,N_9111,N_9983);
and UO_1028 (O_1028,N_9646,N_9332);
nand UO_1029 (O_1029,N_9662,N_9289);
nand UO_1030 (O_1030,N_9695,N_9222);
nand UO_1031 (O_1031,N_9420,N_9461);
nor UO_1032 (O_1032,N_9740,N_9884);
nand UO_1033 (O_1033,N_9853,N_9368);
nand UO_1034 (O_1034,N_9875,N_9787);
nor UO_1035 (O_1035,N_9813,N_9348);
xnor UO_1036 (O_1036,N_9517,N_9781);
or UO_1037 (O_1037,N_9899,N_9519);
and UO_1038 (O_1038,N_9203,N_9367);
and UO_1039 (O_1039,N_9221,N_9125);
xor UO_1040 (O_1040,N_9993,N_9529);
nor UO_1041 (O_1041,N_9463,N_9911);
or UO_1042 (O_1042,N_9862,N_9203);
xnor UO_1043 (O_1043,N_9229,N_9767);
nor UO_1044 (O_1044,N_9947,N_9423);
and UO_1045 (O_1045,N_9929,N_9145);
nand UO_1046 (O_1046,N_9424,N_9102);
nor UO_1047 (O_1047,N_9714,N_9207);
nand UO_1048 (O_1048,N_9132,N_9707);
nor UO_1049 (O_1049,N_9916,N_9387);
nand UO_1050 (O_1050,N_9347,N_9212);
nor UO_1051 (O_1051,N_9435,N_9746);
nor UO_1052 (O_1052,N_9012,N_9444);
and UO_1053 (O_1053,N_9189,N_9117);
nand UO_1054 (O_1054,N_9722,N_9025);
xor UO_1055 (O_1055,N_9095,N_9318);
and UO_1056 (O_1056,N_9210,N_9555);
and UO_1057 (O_1057,N_9343,N_9615);
or UO_1058 (O_1058,N_9537,N_9727);
nand UO_1059 (O_1059,N_9614,N_9672);
nor UO_1060 (O_1060,N_9237,N_9619);
nand UO_1061 (O_1061,N_9604,N_9678);
nor UO_1062 (O_1062,N_9995,N_9805);
nor UO_1063 (O_1063,N_9365,N_9059);
or UO_1064 (O_1064,N_9865,N_9542);
nand UO_1065 (O_1065,N_9537,N_9639);
and UO_1066 (O_1066,N_9593,N_9452);
nand UO_1067 (O_1067,N_9091,N_9311);
nand UO_1068 (O_1068,N_9951,N_9399);
nor UO_1069 (O_1069,N_9129,N_9298);
and UO_1070 (O_1070,N_9564,N_9518);
nand UO_1071 (O_1071,N_9075,N_9867);
nand UO_1072 (O_1072,N_9372,N_9476);
nand UO_1073 (O_1073,N_9393,N_9182);
or UO_1074 (O_1074,N_9152,N_9774);
nand UO_1075 (O_1075,N_9922,N_9699);
nand UO_1076 (O_1076,N_9885,N_9395);
xor UO_1077 (O_1077,N_9048,N_9352);
nand UO_1078 (O_1078,N_9906,N_9418);
xnor UO_1079 (O_1079,N_9375,N_9617);
nand UO_1080 (O_1080,N_9869,N_9441);
or UO_1081 (O_1081,N_9589,N_9563);
or UO_1082 (O_1082,N_9419,N_9126);
and UO_1083 (O_1083,N_9569,N_9148);
or UO_1084 (O_1084,N_9583,N_9710);
nand UO_1085 (O_1085,N_9024,N_9820);
or UO_1086 (O_1086,N_9758,N_9813);
and UO_1087 (O_1087,N_9717,N_9275);
and UO_1088 (O_1088,N_9124,N_9882);
and UO_1089 (O_1089,N_9091,N_9758);
nand UO_1090 (O_1090,N_9873,N_9483);
and UO_1091 (O_1091,N_9448,N_9599);
nand UO_1092 (O_1092,N_9480,N_9489);
nand UO_1093 (O_1093,N_9866,N_9554);
nor UO_1094 (O_1094,N_9468,N_9745);
or UO_1095 (O_1095,N_9333,N_9253);
nand UO_1096 (O_1096,N_9396,N_9507);
nand UO_1097 (O_1097,N_9966,N_9585);
or UO_1098 (O_1098,N_9405,N_9797);
and UO_1099 (O_1099,N_9838,N_9545);
or UO_1100 (O_1100,N_9902,N_9103);
and UO_1101 (O_1101,N_9210,N_9069);
nor UO_1102 (O_1102,N_9962,N_9089);
xnor UO_1103 (O_1103,N_9594,N_9720);
nor UO_1104 (O_1104,N_9559,N_9149);
and UO_1105 (O_1105,N_9032,N_9368);
xnor UO_1106 (O_1106,N_9748,N_9531);
and UO_1107 (O_1107,N_9895,N_9611);
xor UO_1108 (O_1108,N_9705,N_9908);
nand UO_1109 (O_1109,N_9734,N_9313);
or UO_1110 (O_1110,N_9770,N_9257);
and UO_1111 (O_1111,N_9392,N_9351);
nand UO_1112 (O_1112,N_9473,N_9826);
and UO_1113 (O_1113,N_9514,N_9902);
and UO_1114 (O_1114,N_9577,N_9746);
and UO_1115 (O_1115,N_9860,N_9485);
nand UO_1116 (O_1116,N_9428,N_9339);
or UO_1117 (O_1117,N_9435,N_9978);
and UO_1118 (O_1118,N_9592,N_9803);
nand UO_1119 (O_1119,N_9345,N_9550);
nand UO_1120 (O_1120,N_9782,N_9527);
or UO_1121 (O_1121,N_9768,N_9925);
nor UO_1122 (O_1122,N_9082,N_9784);
and UO_1123 (O_1123,N_9132,N_9360);
nor UO_1124 (O_1124,N_9871,N_9109);
or UO_1125 (O_1125,N_9679,N_9460);
nand UO_1126 (O_1126,N_9997,N_9776);
xnor UO_1127 (O_1127,N_9786,N_9444);
or UO_1128 (O_1128,N_9094,N_9701);
or UO_1129 (O_1129,N_9093,N_9598);
or UO_1130 (O_1130,N_9546,N_9696);
and UO_1131 (O_1131,N_9342,N_9960);
and UO_1132 (O_1132,N_9872,N_9443);
xnor UO_1133 (O_1133,N_9425,N_9308);
and UO_1134 (O_1134,N_9370,N_9589);
nor UO_1135 (O_1135,N_9098,N_9894);
nor UO_1136 (O_1136,N_9711,N_9515);
and UO_1137 (O_1137,N_9234,N_9598);
or UO_1138 (O_1138,N_9498,N_9374);
xor UO_1139 (O_1139,N_9995,N_9089);
and UO_1140 (O_1140,N_9889,N_9113);
nor UO_1141 (O_1141,N_9186,N_9120);
and UO_1142 (O_1142,N_9426,N_9410);
and UO_1143 (O_1143,N_9590,N_9362);
and UO_1144 (O_1144,N_9222,N_9943);
nand UO_1145 (O_1145,N_9753,N_9054);
and UO_1146 (O_1146,N_9997,N_9511);
nor UO_1147 (O_1147,N_9570,N_9693);
nand UO_1148 (O_1148,N_9027,N_9509);
nor UO_1149 (O_1149,N_9659,N_9352);
nor UO_1150 (O_1150,N_9351,N_9767);
or UO_1151 (O_1151,N_9473,N_9012);
or UO_1152 (O_1152,N_9523,N_9027);
xnor UO_1153 (O_1153,N_9072,N_9567);
xor UO_1154 (O_1154,N_9150,N_9078);
nor UO_1155 (O_1155,N_9314,N_9619);
and UO_1156 (O_1156,N_9517,N_9997);
nand UO_1157 (O_1157,N_9752,N_9612);
or UO_1158 (O_1158,N_9417,N_9774);
nand UO_1159 (O_1159,N_9917,N_9939);
and UO_1160 (O_1160,N_9015,N_9991);
and UO_1161 (O_1161,N_9014,N_9599);
nor UO_1162 (O_1162,N_9033,N_9120);
nor UO_1163 (O_1163,N_9267,N_9123);
nor UO_1164 (O_1164,N_9295,N_9610);
nand UO_1165 (O_1165,N_9168,N_9310);
and UO_1166 (O_1166,N_9121,N_9315);
and UO_1167 (O_1167,N_9481,N_9137);
or UO_1168 (O_1168,N_9582,N_9134);
nand UO_1169 (O_1169,N_9627,N_9508);
xor UO_1170 (O_1170,N_9435,N_9726);
nor UO_1171 (O_1171,N_9115,N_9203);
nand UO_1172 (O_1172,N_9647,N_9819);
and UO_1173 (O_1173,N_9593,N_9887);
nand UO_1174 (O_1174,N_9459,N_9958);
and UO_1175 (O_1175,N_9594,N_9522);
or UO_1176 (O_1176,N_9418,N_9021);
and UO_1177 (O_1177,N_9764,N_9638);
xnor UO_1178 (O_1178,N_9968,N_9979);
xnor UO_1179 (O_1179,N_9135,N_9283);
and UO_1180 (O_1180,N_9717,N_9660);
nor UO_1181 (O_1181,N_9817,N_9469);
and UO_1182 (O_1182,N_9385,N_9437);
and UO_1183 (O_1183,N_9898,N_9922);
and UO_1184 (O_1184,N_9713,N_9679);
or UO_1185 (O_1185,N_9515,N_9862);
or UO_1186 (O_1186,N_9185,N_9108);
nand UO_1187 (O_1187,N_9317,N_9547);
and UO_1188 (O_1188,N_9007,N_9376);
and UO_1189 (O_1189,N_9059,N_9506);
xor UO_1190 (O_1190,N_9239,N_9710);
and UO_1191 (O_1191,N_9076,N_9207);
nand UO_1192 (O_1192,N_9874,N_9371);
nand UO_1193 (O_1193,N_9646,N_9008);
xnor UO_1194 (O_1194,N_9366,N_9348);
or UO_1195 (O_1195,N_9606,N_9873);
and UO_1196 (O_1196,N_9701,N_9207);
nand UO_1197 (O_1197,N_9645,N_9618);
nor UO_1198 (O_1198,N_9699,N_9727);
xor UO_1199 (O_1199,N_9393,N_9158);
or UO_1200 (O_1200,N_9463,N_9803);
nor UO_1201 (O_1201,N_9215,N_9996);
xnor UO_1202 (O_1202,N_9604,N_9007);
or UO_1203 (O_1203,N_9603,N_9414);
nand UO_1204 (O_1204,N_9757,N_9685);
and UO_1205 (O_1205,N_9216,N_9324);
or UO_1206 (O_1206,N_9568,N_9849);
nor UO_1207 (O_1207,N_9188,N_9329);
and UO_1208 (O_1208,N_9872,N_9624);
xnor UO_1209 (O_1209,N_9025,N_9143);
and UO_1210 (O_1210,N_9886,N_9380);
nor UO_1211 (O_1211,N_9107,N_9713);
xnor UO_1212 (O_1212,N_9343,N_9649);
nand UO_1213 (O_1213,N_9856,N_9086);
nand UO_1214 (O_1214,N_9600,N_9264);
or UO_1215 (O_1215,N_9214,N_9267);
or UO_1216 (O_1216,N_9633,N_9652);
nand UO_1217 (O_1217,N_9089,N_9489);
and UO_1218 (O_1218,N_9589,N_9890);
xnor UO_1219 (O_1219,N_9525,N_9605);
or UO_1220 (O_1220,N_9440,N_9492);
nand UO_1221 (O_1221,N_9732,N_9591);
and UO_1222 (O_1222,N_9943,N_9187);
or UO_1223 (O_1223,N_9547,N_9842);
nor UO_1224 (O_1224,N_9013,N_9050);
nor UO_1225 (O_1225,N_9455,N_9005);
nand UO_1226 (O_1226,N_9683,N_9870);
or UO_1227 (O_1227,N_9505,N_9824);
nor UO_1228 (O_1228,N_9663,N_9484);
nor UO_1229 (O_1229,N_9700,N_9727);
and UO_1230 (O_1230,N_9461,N_9540);
nor UO_1231 (O_1231,N_9696,N_9192);
and UO_1232 (O_1232,N_9270,N_9479);
nand UO_1233 (O_1233,N_9378,N_9335);
and UO_1234 (O_1234,N_9094,N_9442);
nor UO_1235 (O_1235,N_9282,N_9481);
xnor UO_1236 (O_1236,N_9271,N_9283);
and UO_1237 (O_1237,N_9644,N_9612);
xor UO_1238 (O_1238,N_9368,N_9743);
or UO_1239 (O_1239,N_9709,N_9489);
and UO_1240 (O_1240,N_9380,N_9025);
nor UO_1241 (O_1241,N_9432,N_9787);
nor UO_1242 (O_1242,N_9723,N_9339);
nand UO_1243 (O_1243,N_9108,N_9433);
or UO_1244 (O_1244,N_9462,N_9718);
nand UO_1245 (O_1245,N_9610,N_9720);
nor UO_1246 (O_1246,N_9192,N_9933);
or UO_1247 (O_1247,N_9386,N_9470);
or UO_1248 (O_1248,N_9753,N_9166);
nand UO_1249 (O_1249,N_9049,N_9507);
or UO_1250 (O_1250,N_9480,N_9664);
nand UO_1251 (O_1251,N_9144,N_9165);
nor UO_1252 (O_1252,N_9866,N_9415);
nand UO_1253 (O_1253,N_9316,N_9875);
nor UO_1254 (O_1254,N_9259,N_9793);
nand UO_1255 (O_1255,N_9969,N_9886);
and UO_1256 (O_1256,N_9799,N_9395);
and UO_1257 (O_1257,N_9519,N_9939);
or UO_1258 (O_1258,N_9295,N_9872);
or UO_1259 (O_1259,N_9148,N_9355);
nor UO_1260 (O_1260,N_9993,N_9720);
or UO_1261 (O_1261,N_9077,N_9641);
nand UO_1262 (O_1262,N_9784,N_9101);
or UO_1263 (O_1263,N_9199,N_9812);
xor UO_1264 (O_1264,N_9052,N_9896);
nand UO_1265 (O_1265,N_9371,N_9422);
nand UO_1266 (O_1266,N_9857,N_9376);
nor UO_1267 (O_1267,N_9117,N_9164);
xor UO_1268 (O_1268,N_9225,N_9750);
or UO_1269 (O_1269,N_9316,N_9464);
nand UO_1270 (O_1270,N_9720,N_9984);
or UO_1271 (O_1271,N_9674,N_9585);
nand UO_1272 (O_1272,N_9605,N_9347);
xor UO_1273 (O_1273,N_9664,N_9032);
nor UO_1274 (O_1274,N_9296,N_9290);
xnor UO_1275 (O_1275,N_9756,N_9899);
and UO_1276 (O_1276,N_9705,N_9151);
and UO_1277 (O_1277,N_9486,N_9031);
nand UO_1278 (O_1278,N_9251,N_9009);
xor UO_1279 (O_1279,N_9875,N_9361);
nand UO_1280 (O_1280,N_9221,N_9608);
nor UO_1281 (O_1281,N_9451,N_9758);
xnor UO_1282 (O_1282,N_9119,N_9024);
nor UO_1283 (O_1283,N_9888,N_9908);
and UO_1284 (O_1284,N_9166,N_9973);
or UO_1285 (O_1285,N_9750,N_9993);
or UO_1286 (O_1286,N_9977,N_9184);
nand UO_1287 (O_1287,N_9898,N_9825);
and UO_1288 (O_1288,N_9289,N_9459);
or UO_1289 (O_1289,N_9846,N_9028);
nand UO_1290 (O_1290,N_9825,N_9990);
or UO_1291 (O_1291,N_9239,N_9390);
or UO_1292 (O_1292,N_9150,N_9117);
nor UO_1293 (O_1293,N_9877,N_9156);
xor UO_1294 (O_1294,N_9862,N_9474);
nand UO_1295 (O_1295,N_9654,N_9663);
and UO_1296 (O_1296,N_9734,N_9384);
or UO_1297 (O_1297,N_9616,N_9041);
nand UO_1298 (O_1298,N_9298,N_9942);
or UO_1299 (O_1299,N_9786,N_9100);
nand UO_1300 (O_1300,N_9163,N_9962);
nand UO_1301 (O_1301,N_9894,N_9369);
and UO_1302 (O_1302,N_9848,N_9174);
xnor UO_1303 (O_1303,N_9447,N_9280);
or UO_1304 (O_1304,N_9933,N_9744);
xnor UO_1305 (O_1305,N_9736,N_9625);
and UO_1306 (O_1306,N_9570,N_9002);
or UO_1307 (O_1307,N_9921,N_9376);
or UO_1308 (O_1308,N_9469,N_9423);
xor UO_1309 (O_1309,N_9602,N_9527);
and UO_1310 (O_1310,N_9146,N_9902);
nand UO_1311 (O_1311,N_9308,N_9968);
and UO_1312 (O_1312,N_9041,N_9710);
nor UO_1313 (O_1313,N_9776,N_9237);
xnor UO_1314 (O_1314,N_9652,N_9862);
nand UO_1315 (O_1315,N_9059,N_9340);
or UO_1316 (O_1316,N_9410,N_9175);
nor UO_1317 (O_1317,N_9542,N_9115);
or UO_1318 (O_1318,N_9932,N_9790);
or UO_1319 (O_1319,N_9367,N_9015);
and UO_1320 (O_1320,N_9698,N_9779);
nor UO_1321 (O_1321,N_9479,N_9256);
nand UO_1322 (O_1322,N_9811,N_9515);
nand UO_1323 (O_1323,N_9340,N_9982);
xor UO_1324 (O_1324,N_9848,N_9120);
nor UO_1325 (O_1325,N_9316,N_9003);
nand UO_1326 (O_1326,N_9781,N_9522);
or UO_1327 (O_1327,N_9702,N_9670);
nor UO_1328 (O_1328,N_9219,N_9860);
nor UO_1329 (O_1329,N_9773,N_9134);
nor UO_1330 (O_1330,N_9775,N_9178);
nand UO_1331 (O_1331,N_9384,N_9895);
or UO_1332 (O_1332,N_9432,N_9336);
and UO_1333 (O_1333,N_9569,N_9548);
or UO_1334 (O_1334,N_9021,N_9264);
nor UO_1335 (O_1335,N_9023,N_9312);
or UO_1336 (O_1336,N_9622,N_9794);
nor UO_1337 (O_1337,N_9859,N_9502);
xnor UO_1338 (O_1338,N_9718,N_9656);
and UO_1339 (O_1339,N_9115,N_9073);
nand UO_1340 (O_1340,N_9459,N_9418);
and UO_1341 (O_1341,N_9054,N_9108);
and UO_1342 (O_1342,N_9729,N_9683);
nor UO_1343 (O_1343,N_9702,N_9776);
xor UO_1344 (O_1344,N_9409,N_9421);
and UO_1345 (O_1345,N_9055,N_9093);
nand UO_1346 (O_1346,N_9451,N_9766);
nor UO_1347 (O_1347,N_9520,N_9930);
nor UO_1348 (O_1348,N_9735,N_9410);
xnor UO_1349 (O_1349,N_9302,N_9343);
and UO_1350 (O_1350,N_9043,N_9437);
or UO_1351 (O_1351,N_9596,N_9285);
xor UO_1352 (O_1352,N_9362,N_9496);
and UO_1353 (O_1353,N_9784,N_9284);
nand UO_1354 (O_1354,N_9766,N_9283);
nand UO_1355 (O_1355,N_9112,N_9272);
or UO_1356 (O_1356,N_9785,N_9158);
or UO_1357 (O_1357,N_9443,N_9264);
and UO_1358 (O_1358,N_9413,N_9944);
and UO_1359 (O_1359,N_9134,N_9284);
and UO_1360 (O_1360,N_9093,N_9054);
nand UO_1361 (O_1361,N_9864,N_9421);
and UO_1362 (O_1362,N_9443,N_9440);
or UO_1363 (O_1363,N_9269,N_9279);
or UO_1364 (O_1364,N_9043,N_9732);
nand UO_1365 (O_1365,N_9831,N_9474);
nand UO_1366 (O_1366,N_9554,N_9809);
nor UO_1367 (O_1367,N_9530,N_9944);
or UO_1368 (O_1368,N_9730,N_9710);
or UO_1369 (O_1369,N_9140,N_9587);
or UO_1370 (O_1370,N_9657,N_9636);
or UO_1371 (O_1371,N_9112,N_9761);
nor UO_1372 (O_1372,N_9479,N_9412);
or UO_1373 (O_1373,N_9271,N_9277);
nor UO_1374 (O_1374,N_9538,N_9627);
nand UO_1375 (O_1375,N_9980,N_9945);
nor UO_1376 (O_1376,N_9292,N_9625);
and UO_1377 (O_1377,N_9520,N_9179);
and UO_1378 (O_1378,N_9178,N_9992);
nand UO_1379 (O_1379,N_9505,N_9105);
xnor UO_1380 (O_1380,N_9921,N_9703);
and UO_1381 (O_1381,N_9102,N_9165);
nor UO_1382 (O_1382,N_9466,N_9272);
and UO_1383 (O_1383,N_9407,N_9352);
nand UO_1384 (O_1384,N_9729,N_9830);
or UO_1385 (O_1385,N_9223,N_9064);
nor UO_1386 (O_1386,N_9429,N_9173);
and UO_1387 (O_1387,N_9370,N_9584);
or UO_1388 (O_1388,N_9536,N_9903);
or UO_1389 (O_1389,N_9482,N_9481);
and UO_1390 (O_1390,N_9653,N_9041);
nand UO_1391 (O_1391,N_9326,N_9315);
xnor UO_1392 (O_1392,N_9949,N_9346);
nand UO_1393 (O_1393,N_9173,N_9721);
xor UO_1394 (O_1394,N_9646,N_9777);
and UO_1395 (O_1395,N_9174,N_9659);
and UO_1396 (O_1396,N_9887,N_9723);
nand UO_1397 (O_1397,N_9003,N_9213);
or UO_1398 (O_1398,N_9644,N_9423);
nor UO_1399 (O_1399,N_9936,N_9150);
or UO_1400 (O_1400,N_9371,N_9690);
and UO_1401 (O_1401,N_9099,N_9436);
and UO_1402 (O_1402,N_9341,N_9993);
and UO_1403 (O_1403,N_9074,N_9309);
nand UO_1404 (O_1404,N_9393,N_9942);
and UO_1405 (O_1405,N_9767,N_9014);
or UO_1406 (O_1406,N_9446,N_9312);
nand UO_1407 (O_1407,N_9195,N_9067);
or UO_1408 (O_1408,N_9435,N_9944);
or UO_1409 (O_1409,N_9770,N_9107);
nor UO_1410 (O_1410,N_9072,N_9689);
nand UO_1411 (O_1411,N_9368,N_9058);
or UO_1412 (O_1412,N_9893,N_9373);
or UO_1413 (O_1413,N_9091,N_9359);
xnor UO_1414 (O_1414,N_9126,N_9372);
nand UO_1415 (O_1415,N_9025,N_9930);
and UO_1416 (O_1416,N_9017,N_9358);
or UO_1417 (O_1417,N_9470,N_9606);
nor UO_1418 (O_1418,N_9786,N_9876);
nor UO_1419 (O_1419,N_9507,N_9501);
nor UO_1420 (O_1420,N_9598,N_9350);
nand UO_1421 (O_1421,N_9316,N_9046);
or UO_1422 (O_1422,N_9113,N_9247);
nor UO_1423 (O_1423,N_9318,N_9327);
nand UO_1424 (O_1424,N_9662,N_9004);
and UO_1425 (O_1425,N_9410,N_9500);
nor UO_1426 (O_1426,N_9621,N_9955);
nor UO_1427 (O_1427,N_9554,N_9102);
and UO_1428 (O_1428,N_9993,N_9464);
nor UO_1429 (O_1429,N_9890,N_9594);
or UO_1430 (O_1430,N_9238,N_9024);
nor UO_1431 (O_1431,N_9600,N_9629);
or UO_1432 (O_1432,N_9281,N_9788);
nand UO_1433 (O_1433,N_9577,N_9318);
or UO_1434 (O_1434,N_9817,N_9020);
nand UO_1435 (O_1435,N_9610,N_9281);
nand UO_1436 (O_1436,N_9356,N_9784);
nand UO_1437 (O_1437,N_9278,N_9280);
and UO_1438 (O_1438,N_9837,N_9407);
or UO_1439 (O_1439,N_9117,N_9234);
xnor UO_1440 (O_1440,N_9316,N_9253);
and UO_1441 (O_1441,N_9220,N_9720);
or UO_1442 (O_1442,N_9240,N_9283);
xor UO_1443 (O_1443,N_9643,N_9405);
nand UO_1444 (O_1444,N_9895,N_9667);
or UO_1445 (O_1445,N_9799,N_9487);
or UO_1446 (O_1446,N_9798,N_9807);
xnor UO_1447 (O_1447,N_9801,N_9985);
or UO_1448 (O_1448,N_9035,N_9998);
nand UO_1449 (O_1449,N_9972,N_9498);
xor UO_1450 (O_1450,N_9744,N_9946);
nor UO_1451 (O_1451,N_9675,N_9088);
or UO_1452 (O_1452,N_9850,N_9824);
or UO_1453 (O_1453,N_9018,N_9674);
or UO_1454 (O_1454,N_9195,N_9650);
or UO_1455 (O_1455,N_9146,N_9646);
and UO_1456 (O_1456,N_9100,N_9619);
and UO_1457 (O_1457,N_9381,N_9348);
or UO_1458 (O_1458,N_9022,N_9761);
xor UO_1459 (O_1459,N_9893,N_9905);
nand UO_1460 (O_1460,N_9617,N_9940);
or UO_1461 (O_1461,N_9084,N_9080);
nor UO_1462 (O_1462,N_9681,N_9928);
nand UO_1463 (O_1463,N_9535,N_9419);
nor UO_1464 (O_1464,N_9730,N_9961);
and UO_1465 (O_1465,N_9651,N_9531);
and UO_1466 (O_1466,N_9044,N_9029);
nand UO_1467 (O_1467,N_9028,N_9014);
or UO_1468 (O_1468,N_9331,N_9825);
or UO_1469 (O_1469,N_9710,N_9747);
and UO_1470 (O_1470,N_9255,N_9799);
nor UO_1471 (O_1471,N_9047,N_9831);
nor UO_1472 (O_1472,N_9701,N_9706);
or UO_1473 (O_1473,N_9985,N_9599);
nand UO_1474 (O_1474,N_9687,N_9606);
or UO_1475 (O_1475,N_9028,N_9425);
and UO_1476 (O_1476,N_9193,N_9495);
nor UO_1477 (O_1477,N_9293,N_9478);
or UO_1478 (O_1478,N_9102,N_9163);
or UO_1479 (O_1479,N_9688,N_9906);
nor UO_1480 (O_1480,N_9249,N_9814);
nor UO_1481 (O_1481,N_9806,N_9215);
or UO_1482 (O_1482,N_9063,N_9459);
and UO_1483 (O_1483,N_9096,N_9759);
nand UO_1484 (O_1484,N_9066,N_9920);
and UO_1485 (O_1485,N_9746,N_9519);
nor UO_1486 (O_1486,N_9289,N_9622);
nor UO_1487 (O_1487,N_9943,N_9462);
or UO_1488 (O_1488,N_9059,N_9417);
or UO_1489 (O_1489,N_9330,N_9052);
nor UO_1490 (O_1490,N_9233,N_9718);
and UO_1491 (O_1491,N_9412,N_9308);
nor UO_1492 (O_1492,N_9338,N_9015);
xor UO_1493 (O_1493,N_9757,N_9485);
or UO_1494 (O_1494,N_9477,N_9347);
and UO_1495 (O_1495,N_9064,N_9275);
nand UO_1496 (O_1496,N_9376,N_9728);
nand UO_1497 (O_1497,N_9221,N_9841);
and UO_1498 (O_1498,N_9394,N_9668);
and UO_1499 (O_1499,N_9039,N_9106);
endmodule