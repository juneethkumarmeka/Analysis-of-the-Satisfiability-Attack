module basic_1000_10000_1500_100_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_247,In_585);
nor U1 (N_1,In_806,In_305);
or U2 (N_2,In_377,In_203);
or U3 (N_3,In_626,In_907);
nand U4 (N_4,In_942,In_749);
and U5 (N_5,In_498,In_571);
nor U6 (N_6,In_224,In_861);
and U7 (N_7,In_429,In_135);
or U8 (N_8,In_627,In_278);
nor U9 (N_9,In_120,In_478);
nor U10 (N_10,In_386,In_988);
nor U11 (N_11,In_49,In_857);
nand U12 (N_12,In_887,In_670);
nor U13 (N_13,In_338,In_950);
nor U14 (N_14,In_650,In_816);
nand U15 (N_15,In_449,In_606);
and U16 (N_16,In_383,In_916);
or U17 (N_17,In_629,In_704);
nand U18 (N_18,In_503,In_763);
or U19 (N_19,In_355,In_698);
nor U20 (N_20,In_924,In_727);
nand U21 (N_21,In_785,In_294);
nand U22 (N_22,In_753,In_163);
xnor U23 (N_23,In_274,In_989);
or U24 (N_24,In_209,In_463);
and U25 (N_25,In_853,In_660);
nand U26 (N_26,In_783,In_738);
nor U27 (N_27,In_175,In_152);
nor U28 (N_28,In_779,In_872);
and U29 (N_29,In_584,In_51);
and U30 (N_30,In_953,In_179);
or U31 (N_31,In_373,In_101);
or U32 (N_32,In_288,In_107);
and U33 (N_33,In_244,In_636);
nand U34 (N_34,In_888,In_919);
or U35 (N_35,In_524,In_41);
nand U36 (N_36,In_233,In_128);
or U37 (N_37,In_882,In_119);
nor U38 (N_38,In_781,In_60);
or U39 (N_39,In_893,In_889);
or U40 (N_40,In_746,In_789);
or U41 (N_41,In_948,In_743);
or U42 (N_42,In_969,In_741);
nand U43 (N_43,In_612,In_379);
nand U44 (N_44,In_675,In_923);
nor U45 (N_45,In_3,In_103);
nor U46 (N_46,In_326,In_920);
nor U47 (N_47,In_681,In_546);
nor U48 (N_48,In_602,In_508);
and U49 (N_49,In_534,In_501);
and U50 (N_50,In_93,In_553);
nand U51 (N_51,In_620,In_390);
and U52 (N_52,In_207,In_122);
or U53 (N_53,In_809,In_499);
nand U54 (N_54,In_801,In_666);
and U55 (N_55,In_800,In_531);
nand U56 (N_56,In_526,In_655);
or U57 (N_57,In_360,In_631);
nand U58 (N_58,In_72,In_621);
nor U59 (N_59,In_487,In_562);
and U60 (N_60,In_228,In_19);
nand U61 (N_61,In_777,In_140);
and U62 (N_62,In_164,In_593);
or U63 (N_63,In_549,In_538);
and U64 (N_64,In_381,In_929);
nand U65 (N_65,In_730,In_460);
nand U66 (N_66,In_454,In_554);
and U67 (N_67,In_284,In_563);
nand U68 (N_68,In_395,In_413);
and U69 (N_69,In_344,In_346);
or U70 (N_70,In_837,In_664);
nor U71 (N_71,In_514,In_723);
and U72 (N_72,In_48,In_2);
nor U73 (N_73,In_804,In_814);
nand U74 (N_74,In_669,In_637);
nand U75 (N_75,In_291,In_428);
nor U76 (N_76,In_160,In_95);
nand U77 (N_77,In_913,In_261);
and U78 (N_78,In_223,In_699);
or U79 (N_79,In_649,In_695);
nor U80 (N_80,In_201,In_740);
and U81 (N_81,In_263,In_335);
and U82 (N_82,In_40,In_162);
nor U83 (N_83,In_84,In_711);
nor U84 (N_84,In_188,In_46);
nand U85 (N_85,In_974,In_597);
or U86 (N_86,In_232,In_959);
and U87 (N_87,In_547,In_32);
nor U88 (N_88,In_251,In_925);
nand U89 (N_89,In_324,In_735);
or U90 (N_90,In_736,In_427);
and U91 (N_91,In_522,In_677);
nor U92 (N_92,In_174,In_641);
nand U93 (N_93,In_301,In_142);
nand U94 (N_94,In_88,In_517);
or U95 (N_95,In_751,In_716);
nor U96 (N_96,In_805,In_459);
nand U97 (N_97,In_213,In_533);
or U98 (N_98,In_258,In_906);
nand U99 (N_99,In_397,In_333);
and U100 (N_100,In_880,N_88);
nand U101 (N_101,In_292,In_170);
nand U102 (N_102,N_53,In_748);
nand U103 (N_103,In_940,In_29);
nor U104 (N_104,In_802,In_860);
nand U105 (N_105,In_280,In_985);
and U106 (N_106,In_56,In_180);
nor U107 (N_107,In_532,In_234);
nand U108 (N_108,In_218,In_774);
or U109 (N_109,In_370,In_194);
and U110 (N_110,N_33,In_550);
nand U111 (N_111,In_854,N_84);
nand U112 (N_112,In_790,In_874);
nor U113 (N_113,In_693,In_187);
and U114 (N_114,In_718,In_63);
nor U115 (N_115,In_132,In_791);
and U116 (N_116,In_281,In_254);
and U117 (N_117,In_582,N_58);
nand U118 (N_118,N_86,In_473);
or U119 (N_119,In_195,In_976);
nor U120 (N_120,In_839,In_823);
xnor U121 (N_121,In_412,In_944);
or U122 (N_122,In_506,In_239);
and U123 (N_123,In_240,In_462);
nor U124 (N_124,In_375,In_516);
or U125 (N_125,In_332,In_440);
nand U126 (N_126,In_193,In_567);
and U127 (N_127,In_613,In_105);
and U128 (N_128,In_886,In_368);
nor U129 (N_129,In_17,In_795);
nor U130 (N_130,N_97,In_75);
nand U131 (N_131,In_578,In_775);
nor U132 (N_132,In_451,In_0);
and U133 (N_133,In_481,In_868);
or U134 (N_134,In_883,In_200);
and U135 (N_135,In_496,In_938);
nand U136 (N_136,In_756,In_987);
nor U137 (N_137,In_894,N_47);
and U138 (N_138,In_576,In_512);
and U139 (N_139,In_876,In_965);
nand U140 (N_140,In_309,In_958);
or U141 (N_141,N_66,In_124);
nand U142 (N_142,In_519,In_384);
or U143 (N_143,In_125,In_928);
nor U144 (N_144,In_903,In_337);
or U145 (N_145,In_488,In_81);
nand U146 (N_146,In_687,In_729);
nand U147 (N_147,N_15,In_780);
nand U148 (N_148,In_573,N_64);
or U149 (N_149,In_520,In_471);
nor U150 (N_150,N_52,In_22);
or U151 (N_151,In_838,In_416);
nand U152 (N_152,In_156,N_91);
and U153 (N_153,In_461,In_154);
and U154 (N_154,In_173,In_910);
nor U155 (N_155,In_502,In_892);
and U156 (N_156,In_216,In_979);
and U157 (N_157,In_273,In_879);
or U158 (N_158,In_319,In_268);
nor U159 (N_159,In_935,In_235);
or U160 (N_160,In_798,In_21);
or U161 (N_161,In_282,N_79);
or U162 (N_162,In_143,N_34);
nor U163 (N_163,N_51,In_114);
and U164 (N_164,In_214,In_285);
and U165 (N_165,In_971,In_731);
and U166 (N_166,In_432,In_766);
nor U167 (N_167,In_102,In_453);
and U168 (N_168,In_587,In_447);
and U169 (N_169,In_477,In_155);
or U170 (N_170,In_653,In_825);
nand U171 (N_171,In_245,N_70);
nor U172 (N_172,In_89,In_657);
and U173 (N_173,In_212,In_275);
nor U174 (N_174,In_492,In_414);
xnor U175 (N_175,In_850,In_820);
or U176 (N_176,In_867,N_4);
or U177 (N_177,N_10,In_78);
or U178 (N_178,In_583,In_722);
nand U179 (N_179,In_830,In_821);
xor U180 (N_180,In_607,In_991);
or U181 (N_181,N_48,In_912);
nor U182 (N_182,In_742,In_560);
nand U183 (N_183,In_662,In_656);
nor U184 (N_184,In_35,In_425);
and U185 (N_185,In_37,In_541);
nor U186 (N_186,In_8,In_100);
nand U187 (N_187,In_276,In_786);
and U188 (N_188,N_69,In_359);
nor U189 (N_189,In_286,In_69);
nor U190 (N_190,In_392,In_984);
or U191 (N_191,N_85,In_467);
nand U192 (N_192,In_28,In_199);
xor U193 (N_193,In_34,N_43);
or U194 (N_194,In_497,In_856);
and U195 (N_195,In_895,In_761);
or U196 (N_196,N_9,In_181);
nand U197 (N_197,In_642,In_446);
and U198 (N_198,In_443,In_537);
and U199 (N_199,In_436,In_66);
or U200 (N_200,In_972,In_376);
nor U201 (N_201,In_401,N_105);
nor U202 (N_202,In_864,In_166);
nor U203 (N_203,In_954,N_135);
or U204 (N_204,In_82,In_702);
nor U205 (N_205,In_57,N_149);
nor U206 (N_206,In_189,In_115);
and U207 (N_207,N_36,In_847);
or U208 (N_208,N_130,In_130);
or U209 (N_209,In_126,In_172);
nand U210 (N_210,In_283,In_431);
nor U211 (N_211,In_904,N_41);
or U212 (N_212,N_198,In_248);
and U213 (N_213,N_113,In_202);
and U214 (N_214,In_339,N_154);
and U215 (N_215,In_515,In_683);
nor U216 (N_216,In_588,N_155);
and U217 (N_217,In_772,In_523);
and U218 (N_218,In_243,In_437);
nor U219 (N_219,In_387,N_195);
nor U220 (N_220,N_147,N_168);
and U221 (N_221,N_29,In_225);
nor U222 (N_222,In_577,In_411);
nor U223 (N_223,In_262,In_53);
and U224 (N_224,In_430,In_851);
xnor U225 (N_225,In_109,In_267);
nor U226 (N_226,N_136,In_651);
nor U227 (N_227,In_625,In_967);
and U228 (N_228,N_127,In_362);
nand U229 (N_229,In_726,In_192);
nor U230 (N_230,In_956,In_369);
and U231 (N_231,In_827,In_198);
and U232 (N_232,In_6,In_391);
and U233 (N_233,In_638,N_106);
nand U234 (N_234,In_231,In_83);
nor U235 (N_235,In_983,N_131);
nand U236 (N_236,In_659,N_199);
nand U237 (N_237,In_870,In_771);
nor U238 (N_238,In_226,In_685);
nand U239 (N_239,In_765,In_978);
nand U240 (N_240,N_189,In_450);
or U241 (N_241,In_494,N_7);
nand U242 (N_242,In_371,In_529);
nand U243 (N_243,In_993,N_151);
nor U244 (N_244,In_306,In_848);
or U245 (N_245,In_921,In_891);
and U246 (N_246,N_188,In_684);
and U247 (N_247,In_632,In_485);
or U248 (N_248,In_551,N_143);
nand U249 (N_249,N_187,In_253);
nor U250 (N_250,In_590,N_122);
or U251 (N_251,In_14,In_323);
nor U252 (N_252,In_438,In_776);
or U253 (N_253,In_465,N_44);
nor U254 (N_254,In_559,In_828);
nand U255 (N_255,In_250,In_961);
or U256 (N_256,In_493,N_111);
nor U257 (N_257,In_707,In_222);
and U258 (N_258,In_968,In_768);
nor U259 (N_259,N_139,In_778);
xor U260 (N_260,N_197,In_30);
nand U261 (N_261,In_113,In_25);
nor U262 (N_262,In_121,In_604);
nand U263 (N_263,In_490,In_7);
and U264 (N_264,In_236,In_62);
nor U265 (N_265,In_530,In_106);
or U266 (N_266,In_605,In_215);
and U267 (N_267,In_564,In_665);
or U268 (N_268,In_676,In_782);
nand U269 (N_269,In_873,In_327);
nand U270 (N_270,In_720,N_186);
or U271 (N_271,In_74,In_586);
or U272 (N_272,N_27,In_445);
and U273 (N_273,In_65,In_405);
or U274 (N_274,In_183,In_382);
and U275 (N_275,In_843,In_316);
nand U276 (N_276,In_943,In_992);
or U277 (N_277,In_813,N_180);
and U278 (N_278,N_123,In_509);
nand U279 (N_279,In_673,In_350);
or U280 (N_280,In_518,In_762);
or U281 (N_281,In_456,In_812);
nor U282 (N_282,In_271,N_171);
and U283 (N_283,In_16,In_378);
nor U284 (N_284,In_527,In_308);
nand U285 (N_285,In_73,In_952);
nand U286 (N_286,In_97,In_340);
or U287 (N_287,N_173,In_982);
nand U288 (N_288,In_939,In_930);
nand U289 (N_289,In_246,In_832);
or U290 (N_290,In_737,In_354);
nor U291 (N_291,In_668,In_468);
or U292 (N_292,In_70,In_334);
nand U293 (N_293,In_259,In_616);
and U294 (N_294,In_544,In_936);
nand U295 (N_295,N_83,In_739);
nand U296 (N_296,N_163,In_858);
xor U297 (N_297,In_455,N_183);
nor U298 (N_298,In_433,N_71);
nor U299 (N_299,N_121,In_208);
and U300 (N_300,In_205,In_141);
nor U301 (N_301,N_264,N_277);
nand U302 (N_302,In_315,In_165);
or U303 (N_303,N_169,In_400);
nor U304 (N_304,In_557,In_866);
nand U305 (N_305,N_179,N_279);
nand U306 (N_306,In_824,In_941);
nor U307 (N_307,N_112,N_270);
nand U308 (N_308,In_725,In_347);
nand U309 (N_309,In_365,N_0);
and U310 (N_310,In_622,In_482);
or U311 (N_311,In_300,In_901);
and U312 (N_312,In_787,In_513);
nand U313 (N_313,In_877,N_45);
and U314 (N_314,N_203,In_915);
and U315 (N_315,N_204,N_231);
and U316 (N_316,N_172,In_238);
or U317 (N_317,In_568,In_998);
and U318 (N_318,In_389,In_962);
nor U319 (N_319,In_363,N_22);
nand U320 (N_320,In_426,In_321);
nor U321 (N_321,N_108,In_525);
nor U322 (N_322,In_331,N_35);
and U323 (N_323,N_117,In_634);
and U324 (N_324,N_274,N_242);
and U325 (N_325,In_840,In_191);
and U326 (N_326,In_628,In_717);
and U327 (N_327,In_313,In_618);
nand U328 (N_328,In_47,N_75);
nand U329 (N_329,In_701,In_980);
and U330 (N_330,In_922,In_819);
nor U331 (N_331,N_298,N_82);
nand U332 (N_332,In_815,In_808);
nand U333 (N_333,In_311,In_754);
xnor U334 (N_334,In_548,In_177);
nand U335 (N_335,In_591,In_317);
nand U336 (N_336,N_252,In_706);
nand U337 (N_337,In_85,N_296);
and U338 (N_338,In_20,N_220);
nand U339 (N_339,In_862,N_262);
nand U340 (N_340,In_667,In_277);
nor U341 (N_341,N_156,In_398);
nor U342 (N_342,In_844,In_932);
and U343 (N_343,N_80,In_713);
nand U344 (N_344,In_421,In_734);
and U345 (N_345,In_5,In_750);
and U346 (N_346,In_303,In_169);
or U347 (N_347,In_764,In_957);
nand U348 (N_348,In_836,In_36);
or U349 (N_349,N_176,N_282);
nor U350 (N_350,In_26,In_594);
or U351 (N_351,In_186,In_144);
or U352 (N_352,In_279,In_320);
nor U353 (N_353,In_715,N_213);
and U354 (N_354,In_402,N_124);
nand U355 (N_355,N_193,In_648);
nand U356 (N_356,In_674,In_964);
or U357 (N_357,N_225,In_690);
nand U358 (N_358,In_33,N_3);
and U359 (N_359,N_288,In_803);
and U360 (N_360,N_60,In_325);
or U361 (N_361,N_177,In_349);
or U362 (N_362,In_403,In_946);
nor U363 (N_363,In_543,In_671);
or U364 (N_364,In_732,In_176);
nor U365 (N_365,In_849,In_457);
and U366 (N_366,In_875,In_977);
nor U367 (N_367,In_127,N_20);
or U368 (N_368,In_408,N_251);
or U369 (N_369,In_792,In_747);
or U370 (N_370,N_54,In_452);
nor U371 (N_371,In_329,In_694);
or U372 (N_372,N_164,N_243);
and U373 (N_373,In_10,In_710);
and U374 (N_374,In_146,N_216);
nand U375 (N_375,N_275,In_111);
nor U376 (N_376,In_491,In_788);
nand U377 (N_377,In_52,N_87);
and U378 (N_378,In_855,In_799);
and U379 (N_379,N_217,In_973);
nand U380 (N_380,In_96,N_258);
nor U381 (N_381,In_769,In_380);
and U382 (N_382,In_500,In_15);
nor U383 (N_383,In_934,In_117);
nor U384 (N_384,N_161,N_272);
or U385 (N_385,In_296,In_709);
nor U386 (N_386,N_240,In_909);
and U387 (N_387,N_56,In_302);
nand U388 (N_388,In_150,N_283);
nor U389 (N_389,In_592,N_207);
nand U390 (N_390,In_635,In_572);
and U391 (N_391,In_947,In_406);
or U392 (N_392,N_294,N_93);
or U393 (N_393,N_61,N_30);
or U394 (N_394,N_185,N_192);
nor U395 (N_395,N_98,N_221);
nand U396 (N_396,In_996,In_77);
nor U397 (N_397,N_158,N_201);
and U398 (N_398,In_185,N_18);
and U399 (N_399,In_797,N_153);
nand U400 (N_400,N_101,N_342);
xnor U401 (N_401,N_336,In_841);
nand U402 (N_402,In_345,In_831);
and U403 (N_403,N_137,In_184);
or U404 (N_404,In_61,In_417);
nand U405 (N_405,In_700,N_394);
nand U406 (N_406,N_381,N_134);
or U407 (N_407,In_86,N_109);
and U408 (N_408,In_385,In_71);
nand U409 (N_409,In_511,In_639);
or U410 (N_410,N_212,In_611);
nand U411 (N_411,N_307,N_306);
nor U412 (N_412,N_19,N_194);
or U413 (N_413,In_811,N_219);
or U414 (N_414,N_73,N_318);
or U415 (N_415,In_24,In_342);
nand U416 (N_416,In_104,In_39);
and U417 (N_417,In_558,N_59);
and U418 (N_418,N_377,N_326);
nand U419 (N_419,N_315,In_31);
nand U420 (N_420,In_569,N_133);
nand U421 (N_421,N_14,N_364);
nand U422 (N_422,In_647,In_679);
and U423 (N_423,N_317,In_990);
nand U424 (N_424,In_341,In_640);
and U425 (N_425,In_817,In_474);
nand U426 (N_426,N_202,In_298);
or U427 (N_427,In_691,In_242);
nor U428 (N_428,In_328,N_360);
nor U429 (N_429,In_835,In_744);
or U430 (N_430,In_322,N_375);
and U431 (N_431,In_505,N_150);
nand U432 (N_432,In_859,In_834);
nand U433 (N_433,In_682,In_241);
nor U434 (N_434,N_370,In_353);
and U435 (N_435,N_6,In_937);
nor U436 (N_436,N_140,In_469);
and U437 (N_437,N_353,In_507);
or U438 (N_438,In_266,N_266);
nand U439 (N_439,N_392,In_926);
or U440 (N_440,N_387,In_139);
or U441 (N_441,N_119,N_365);
and U442 (N_442,In_536,In_396);
nor U443 (N_443,N_68,In_908);
nand U444 (N_444,In_483,In_999);
nand U445 (N_445,N_398,N_23);
xor U446 (N_446,N_99,N_196);
nand U447 (N_447,N_8,N_289);
nor U448 (N_448,N_238,N_182);
nand U449 (N_449,In_419,In_479);
nand U450 (N_450,In_129,In_609);
nor U451 (N_451,In_168,In_884);
and U452 (N_452,N_312,In_80);
or U453 (N_453,N_178,N_241);
nor U454 (N_454,In_272,N_284);
and U455 (N_455,In_68,In_4);
nand U456 (N_456,In_480,N_391);
or U457 (N_457,In_237,In_204);
nand U458 (N_458,In_917,N_40);
and U459 (N_459,In_364,N_148);
nor U460 (N_460,In_914,N_354);
nor U461 (N_461,N_367,In_435);
or U462 (N_462,In_661,In_151);
nand U463 (N_463,N_371,In_295);
nand U464 (N_464,In_595,In_409);
and U465 (N_465,In_423,In_58);
and U466 (N_466,N_335,In_133);
or U467 (N_467,N_361,In_94);
nor U468 (N_468,In_489,In_18);
and U469 (N_469,N_222,N_349);
or U470 (N_470,N_286,N_292);
nand U471 (N_471,N_362,N_1);
nand U472 (N_472,In_178,N_350);
and U473 (N_473,N_146,In_970);
and U474 (N_474,In_846,N_248);
nor U475 (N_475,In_312,In_424);
and U476 (N_476,N_311,N_107);
nor U477 (N_477,In_986,In_336);
nor U478 (N_478,N_190,In_829);
and U479 (N_479,In_818,N_114);
nor U480 (N_480,N_17,In_442);
xnor U481 (N_481,In_878,N_285);
nand U482 (N_482,In_255,N_141);
nand U483 (N_483,N_366,N_309);
nor U484 (N_484,In_955,N_230);
and U485 (N_485,N_94,In_42);
and U486 (N_486,N_323,N_55);
nor U487 (N_487,N_74,N_281);
nand U488 (N_488,In_918,In_692);
xnor U489 (N_489,In_608,In_310);
or U490 (N_490,In_356,N_343);
or U491 (N_491,In_615,In_902);
or U492 (N_492,In_314,In_504);
or U493 (N_493,N_256,In_897);
and U494 (N_494,N_390,In_374);
or U495 (N_495,N_234,N_351);
nor U496 (N_496,In_589,N_162);
nor U497 (N_497,N_316,N_12);
nor U498 (N_498,In_475,In_148);
nor U499 (N_499,N_16,In_367);
nand U500 (N_500,N_499,In_357);
nor U501 (N_501,N_62,N_409);
nor U502 (N_502,N_175,N_303);
nand U503 (N_503,N_125,N_466);
nand U504 (N_504,N_77,In_997);
or U505 (N_505,N_407,In_610);
and U506 (N_506,In_784,In_542);
nand U507 (N_507,In_171,In_911);
nor U508 (N_508,In_869,N_340);
nor U509 (N_509,In_257,In_249);
and U510 (N_510,N_310,In_833);
and U511 (N_511,N_430,N_115);
or U512 (N_512,N_411,In_287);
nand U513 (N_513,N_450,In_822);
or U514 (N_514,In_528,N_498);
or U515 (N_515,N_302,N_299);
nand U516 (N_516,In_458,N_226);
and U517 (N_517,In_535,In_394);
and U518 (N_518,N_301,N_287);
and U519 (N_519,N_260,N_254);
nand U520 (N_520,In_905,N_305);
and U521 (N_521,N_257,In_566);
and U522 (N_522,In_221,In_646);
nand U523 (N_523,In_949,N_293);
or U524 (N_524,N_482,N_273);
nand U525 (N_525,In_76,In_299);
nand U526 (N_526,In_210,N_261);
nor U527 (N_527,N_157,N_434);
nand U528 (N_528,In_933,N_21);
nor U529 (N_529,In_420,N_104);
nor U530 (N_530,In_770,In_404);
or U531 (N_531,N_400,In_318);
nor U532 (N_532,In_697,In_190);
nand U533 (N_533,In_11,N_470);
nand U534 (N_534,N_457,N_278);
nor U535 (N_535,In_719,In_79);
or U536 (N_536,N_31,In_900);
nor U537 (N_537,N_170,N_223);
nand U538 (N_538,In_182,In_466);
or U539 (N_539,N_489,N_441);
and U540 (N_540,In_12,In_898);
nor U541 (N_541,In_598,In_863);
nand U542 (N_542,N_465,N_235);
and U543 (N_543,In_624,N_237);
nand U544 (N_544,In_773,N_355);
or U545 (N_545,N_428,In_845);
nor U546 (N_546,In_108,N_356);
nor U547 (N_547,N_330,N_13);
or U548 (N_548,N_280,In_724);
nor U549 (N_549,In_663,N_167);
and U550 (N_550,N_333,N_493);
and U551 (N_551,N_89,In_149);
nor U552 (N_552,N_295,In_206);
and U553 (N_553,In_269,N_92);
nor U554 (N_554,N_422,N_291);
or U555 (N_555,N_246,N_11);
xor U556 (N_556,N_420,In_721);
nand U557 (N_557,N_232,N_473);
nor U558 (N_558,In_219,In_539);
and U559 (N_559,In_112,In_118);
nand U560 (N_560,In_220,In_90);
and U561 (N_561,N_346,N_247);
nand U562 (N_562,N_477,N_385);
and U563 (N_563,N_455,N_81);
nor U564 (N_564,N_494,In_654);
or U565 (N_565,N_447,N_384);
and U566 (N_566,In_44,N_379);
or U567 (N_567,In_495,N_78);
nor U568 (N_568,In_393,N_142);
nand U569 (N_569,N_308,In_601);
and U570 (N_570,N_438,In_960);
nand U571 (N_571,N_200,In_145);
nor U572 (N_572,N_174,N_191);
nand U573 (N_573,In_230,N_250);
or U574 (N_574,N_96,N_476);
nor U575 (N_575,In_561,N_345);
or U576 (N_576,In_439,In_197);
and U577 (N_577,In_13,In_758);
nor U578 (N_578,In_658,In_50);
nor U579 (N_579,N_358,In_91);
or U580 (N_580,In_510,N_244);
nor U581 (N_581,N_459,In_330);
or U582 (N_582,In_352,In_167);
or U583 (N_583,N_205,In_422);
nor U584 (N_584,N_485,N_57);
nor U585 (N_585,N_253,In_600);
nor U586 (N_586,In_289,In_927);
nand U587 (N_587,In_521,N_472);
and U588 (N_588,In_565,N_374);
and U589 (N_589,In_159,In_229);
nand U590 (N_590,In_434,In_871);
nor U591 (N_591,N_263,N_159);
nor U592 (N_592,In_472,N_116);
nand U593 (N_593,N_456,In_38);
nor U594 (N_594,In_767,In_484);
or U595 (N_595,N_396,N_389);
or U596 (N_596,In_297,In_304);
or U597 (N_597,In_64,In_540);
or U598 (N_598,N_432,In_161);
or U599 (N_599,In_116,N_458);
and U600 (N_600,N_368,N_118);
nand U601 (N_601,In_556,In_796);
nand U602 (N_602,N_581,N_423);
and U603 (N_603,N_512,N_442);
nand U604 (N_604,In_358,N_344);
or U605 (N_605,In_705,N_320);
and U606 (N_606,In_623,N_388);
or U607 (N_607,In_633,N_506);
nand U608 (N_608,N_592,N_297);
and U609 (N_609,In_388,N_545);
or U610 (N_610,N_559,N_443);
nor U611 (N_611,In_696,N_495);
nor U612 (N_612,In_966,In_826);
or U613 (N_613,N_478,N_215);
nand U614 (N_614,N_380,N_401);
nor U615 (N_615,In_27,In_464);
nor U616 (N_616,N_427,N_322);
and U617 (N_617,N_525,N_555);
nand U618 (N_618,In_852,N_313);
nand U619 (N_619,N_469,N_576);
and U620 (N_620,N_414,N_540);
nor U621 (N_621,In_652,In_963);
and U622 (N_622,In_153,N_503);
nor U623 (N_623,N_321,In_410);
nor U624 (N_624,In_614,N_547);
nand U625 (N_625,N_590,N_586);
and U626 (N_626,In_415,N_339);
nor U627 (N_627,N_446,N_208);
nor U628 (N_628,N_424,In_366);
nand U629 (N_629,N_558,N_399);
nor U630 (N_630,In_55,N_550);
and U631 (N_631,N_425,In_945);
nor U632 (N_632,N_564,N_429);
or U633 (N_633,N_519,In_728);
nor U634 (N_634,N_276,N_544);
and U635 (N_635,In_994,In_137);
or U636 (N_636,N_413,N_583);
nor U637 (N_637,In_759,N_239);
or U638 (N_638,In_348,N_166);
nor U639 (N_639,N_37,N_484);
or U640 (N_640,In_545,In_689);
or U641 (N_641,N_445,N_483);
nor U642 (N_642,N_419,N_341);
nand U643 (N_643,N_562,N_67);
nor U644 (N_644,N_488,N_566);
nor U645 (N_645,In_678,N_210);
or U646 (N_646,N_541,N_319);
nand U647 (N_647,N_408,In_43);
or U648 (N_648,N_265,N_329);
nand U649 (N_649,N_145,N_211);
nand U650 (N_650,N_426,N_572);
or U651 (N_651,In_448,N_599);
xor U652 (N_652,N_505,N_460);
and U653 (N_653,N_501,N_249);
nor U654 (N_654,N_363,N_132);
and U655 (N_655,N_152,N_593);
nand U656 (N_656,In_899,N_421);
and U657 (N_657,In_147,N_463);
and U658 (N_658,N_492,N_334);
and U659 (N_659,In_110,N_65);
and U660 (N_660,N_481,N_383);
or U661 (N_661,N_435,N_449);
or U662 (N_662,In_157,N_556);
or U663 (N_663,In_476,N_487);
and U664 (N_664,N_72,In_307);
or U665 (N_665,N_528,N_209);
nand U666 (N_666,In_59,In_619);
nor U667 (N_667,N_454,N_395);
nor U668 (N_668,In_418,In_580);
or U669 (N_669,N_259,N_522);
or U670 (N_670,N_557,In_931);
and U671 (N_671,In_570,N_575);
and U672 (N_672,N_596,N_582);
nor U673 (N_673,N_28,N_521);
or U674 (N_674,N_453,N_526);
or U675 (N_675,N_475,N_589);
nor U676 (N_676,N_497,N_144);
nor U677 (N_677,In_865,N_38);
and U678 (N_678,N_338,In_842);
nand U679 (N_679,N_448,N_537);
or U680 (N_680,N_32,In_441);
or U681 (N_681,N_378,N_439);
nor U682 (N_682,In_270,N_382);
or U683 (N_683,N_26,N_569);
nand U684 (N_684,N_510,In_293);
nand U685 (N_685,N_165,N_103);
nand U686 (N_686,In_995,N_507);
and U687 (N_687,N_224,In_67);
nor U688 (N_688,N_328,In_703);
nor U689 (N_689,N_417,N_160);
or U690 (N_690,N_227,N_406);
and U691 (N_691,N_267,N_245);
and U692 (N_692,N_546,In_351);
nand U693 (N_693,In_686,In_290);
nand U694 (N_694,N_444,In_712);
and U695 (N_695,N_534,In_158);
and U696 (N_696,N_184,N_515);
or U697 (N_697,N_517,N_128);
or U698 (N_698,In_951,In_575);
nand U699 (N_699,In_981,N_595);
nor U700 (N_700,In_555,N_467);
and U701 (N_701,N_615,N_620);
or U702 (N_702,N_669,N_337);
nor U703 (N_703,N_46,N_348);
nand U704 (N_704,N_551,N_479);
or U705 (N_705,In_680,N_491);
nand U706 (N_706,N_588,N_416);
or U707 (N_707,N_233,In_211);
nand U708 (N_708,In_596,N_535);
nand U709 (N_709,N_674,N_580);
nand U710 (N_710,N_325,N_471);
or U711 (N_711,N_613,N_561);
nand U712 (N_712,In_881,N_508);
and U713 (N_713,In_644,N_689);
and U714 (N_714,N_542,In_794);
nand U715 (N_715,N_630,In_54);
nor U716 (N_716,N_636,N_431);
or U717 (N_717,N_633,In_733);
xor U718 (N_718,N_181,N_656);
nor U719 (N_719,N_665,N_655);
or U720 (N_720,N_587,In_885);
and U721 (N_721,In_45,N_598);
or U722 (N_722,N_486,N_623);
and U723 (N_723,N_269,In_810);
or U724 (N_724,N_24,N_5);
nand U725 (N_725,In_227,N_357);
nor U726 (N_726,N_677,In_708);
nand U727 (N_727,N_39,N_645);
nand U728 (N_728,N_662,N_440);
nand U729 (N_729,N_638,N_553);
nand U730 (N_730,N_462,In_9);
nand U731 (N_731,N_402,In_87);
nor U732 (N_732,N_410,In_552);
nor U733 (N_733,N_681,N_678);
and U734 (N_734,N_110,N_602);
nor U735 (N_735,N_290,In_131);
nor U736 (N_736,N_625,N_412);
and U737 (N_737,N_403,N_527);
nand U738 (N_738,In_23,N_516);
or U739 (N_739,N_352,N_324);
or U740 (N_740,N_331,N_639);
nor U741 (N_741,N_650,N_304);
or U742 (N_742,N_415,In_196);
nor U743 (N_743,In_630,N_671);
nor U744 (N_744,N_138,N_609);
or U745 (N_745,N_579,N_691);
and U746 (N_746,N_666,In_599);
or U747 (N_747,N_663,In_361);
and U748 (N_748,In_890,N_622);
nor U749 (N_749,N_628,In_757);
and U750 (N_750,N_271,N_653);
or U751 (N_751,N_659,In_688);
nand U752 (N_752,N_605,N_654);
nor U753 (N_753,In_645,N_675);
and U754 (N_754,N_397,N_42);
or U755 (N_755,N_464,N_643);
or U756 (N_756,In_217,N_372);
nand U757 (N_757,N_687,N_529);
and U758 (N_758,N_601,In_444);
and U759 (N_759,N_696,N_533);
nand U760 (N_760,N_206,N_651);
and U761 (N_761,N_120,In_264);
nor U762 (N_762,N_695,N_634);
and U763 (N_763,In_260,N_359);
nor U764 (N_764,In_975,N_574);
and U765 (N_765,N_619,N_536);
nand U766 (N_766,N_490,N_560);
nor U767 (N_767,N_693,N_538);
nor U768 (N_768,In_752,N_218);
nor U769 (N_769,In_793,N_514);
nand U770 (N_770,N_692,N_608);
nor U771 (N_771,N_660,In_617);
or U772 (N_772,N_618,N_658);
nor U773 (N_773,N_376,N_688);
nor U774 (N_774,N_631,In_486);
and U775 (N_775,N_474,In_399);
and U776 (N_776,N_554,N_698);
or U777 (N_777,N_641,N_25);
or U778 (N_778,In_123,N_679);
nand U779 (N_779,N_690,In_134);
or U780 (N_780,N_578,N_667);
or U781 (N_781,N_255,N_567);
nand U782 (N_782,N_332,N_228);
or U783 (N_783,N_452,N_617);
or U784 (N_784,N_451,N_480);
nor U785 (N_785,N_606,N_511);
nand U786 (N_786,N_577,N_664);
and U787 (N_787,N_612,In_603);
and U788 (N_788,In_760,N_642);
and U789 (N_789,N_63,N_552);
nor U790 (N_790,N_647,In_745);
nor U791 (N_791,In_714,N_386);
nand U792 (N_792,N_649,N_548);
or U793 (N_793,N_699,In_252);
and U794 (N_794,N_697,N_102);
nor U795 (N_795,N_657,N_661);
and U796 (N_796,N_673,N_585);
and U797 (N_797,N_90,N_314);
and U798 (N_798,N_646,In_470);
nand U799 (N_799,N_129,N_597);
nor U800 (N_800,N_229,N_716);
and U801 (N_801,N_758,N_502);
and U802 (N_802,N_749,N_773);
and U803 (N_803,N_733,N_707);
nor U804 (N_804,N_761,N_781);
nand U805 (N_805,N_685,N_539);
nor U806 (N_806,N_794,N_702);
nor U807 (N_807,N_727,N_746);
and U808 (N_808,In_136,N_327);
nor U809 (N_809,N_76,N_621);
nand U810 (N_810,N_635,N_571);
xor U811 (N_811,N_783,N_709);
nor U812 (N_812,In_643,N_752);
or U813 (N_813,N_762,N_787);
nor U814 (N_814,In_574,N_763);
or U815 (N_815,N_437,N_607);
or U816 (N_816,N_748,N_710);
and U817 (N_817,N_404,N_772);
and U818 (N_818,N_790,N_543);
nor U819 (N_819,N_686,In_672);
and U820 (N_820,N_683,N_523);
and U821 (N_821,N_680,N_524);
and U822 (N_822,N_672,N_405);
nor U823 (N_823,N_676,N_518);
or U824 (N_824,N_573,N_779);
nor U825 (N_825,N_670,N_744);
nor U826 (N_826,N_776,N_706);
and U827 (N_827,N_730,N_624);
and U828 (N_828,N_268,N_629);
nor U829 (N_829,N_784,N_775);
or U830 (N_830,In_807,N_714);
and U831 (N_831,N_728,N_718);
or U832 (N_832,N_789,N_725);
and U833 (N_833,N_369,N_49);
and U834 (N_834,N_782,In_407);
or U835 (N_835,N_610,N_513);
or U836 (N_836,In_92,N_726);
and U837 (N_837,N_770,N_591);
and U838 (N_838,N_721,N_739);
or U839 (N_839,N_682,N_766);
and U840 (N_840,N_715,N_594);
nand U841 (N_841,N_461,N_720);
nor U842 (N_842,N_694,N_793);
and U843 (N_843,In_343,N_756);
nor U844 (N_844,N_757,N_703);
nor U845 (N_845,In_896,N_504);
nor U846 (N_846,N_765,N_743);
nand U847 (N_847,N_614,N_640);
nand U848 (N_848,N_436,N_236);
nor U849 (N_849,N_767,N_719);
nor U850 (N_850,N_759,N_214);
or U851 (N_851,N_668,N_632);
nor U852 (N_852,N_126,N_785);
nand U853 (N_853,N_788,N_393);
nand U854 (N_854,N_532,N_717);
and U855 (N_855,N_791,N_611);
nor U856 (N_856,N_565,In_1);
and U857 (N_857,N_627,N_700);
or U858 (N_858,N_745,N_786);
nor U859 (N_859,N_778,N_652);
nor U860 (N_860,N_373,N_780);
and U861 (N_861,N_734,N_755);
nand U862 (N_862,N_704,N_637);
and U863 (N_863,N_732,N_712);
or U864 (N_864,In_581,N_729);
or U865 (N_865,N_549,N_722);
nand U866 (N_866,N_747,N_735);
nor U867 (N_867,In_99,In_579);
nor U868 (N_868,N_626,N_563);
or U869 (N_869,N_496,N_764);
nor U870 (N_870,N_468,In_98);
and U871 (N_871,N_705,N_568);
and U872 (N_872,N_797,In_138);
nor U873 (N_873,N_713,N_95);
and U874 (N_874,N_711,N_520);
or U875 (N_875,N_570,In_265);
or U876 (N_876,N_648,N_530);
nor U877 (N_877,N_708,N_500);
and U878 (N_878,N_799,N_531);
or U879 (N_879,N_300,N_701);
nor U880 (N_880,N_600,N_731);
and U881 (N_881,N_796,N_603);
and U882 (N_882,N_741,N_753);
nand U883 (N_883,In_256,N_724);
and U884 (N_884,N_777,N_737);
nand U885 (N_885,N_792,In_755);
nand U886 (N_886,N_509,N_751);
and U887 (N_887,N_768,N_644);
and U888 (N_888,N_740,N_750);
nor U889 (N_889,N_798,In_372);
or U890 (N_890,N_736,N_771);
nand U891 (N_891,N_2,N_769);
nand U892 (N_892,N_604,N_616);
nor U893 (N_893,N_684,N_347);
and U894 (N_894,N_742,N_738);
xnor U895 (N_895,N_584,N_433);
nor U896 (N_896,N_100,N_754);
and U897 (N_897,N_723,N_760);
and U898 (N_898,N_774,N_795);
or U899 (N_899,N_418,N_50);
and U900 (N_900,N_849,N_824);
nand U901 (N_901,N_836,N_886);
nand U902 (N_902,N_855,N_827);
nor U903 (N_903,N_882,N_876);
nor U904 (N_904,N_837,N_877);
or U905 (N_905,N_852,N_872);
and U906 (N_906,N_897,N_833);
or U907 (N_907,N_864,N_845);
nor U908 (N_908,N_854,N_846);
xor U909 (N_909,N_853,N_899);
or U910 (N_910,N_868,N_856);
nand U911 (N_911,N_875,N_890);
nor U912 (N_912,N_832,N_884);
or U913 (N_913,N_857,N_835);
nor U914 (N_914,N_848,N_851);
or U915 (N_915,N_870,N_802);
nor U916 (N_916,N_804,N_831);
or U917 (N_917,N_883,N_895);
or U918 (N_918,N_841,N_859);
nor U919 (N_919,N_823,N_842);
nor U920 (N_920,N_879,N_892);
nor U921 (N_921,N_838,N_821);
or U922 (N_922,N_801,N_828);
nor U923 (N_923,N_881,N_820);
nand U924 (N_924,N_812,N_826);
or U925 (N_925,N_850,N_865);
nand U926 (N_926,N_816,N_805);
and U927 (N_927,N_810,N_803);
and U928 (N_928,N_874,N_834);
nand U929 (N_929,N_861,N_825);
nor U930 (N_930,N_893,N_887);
nor U931 (N_931,N_817,N_822);
xor U932 (N_932,N_871,N_896);
nor U933 (N_933,N_869,N_847);
or U934 (N_934,N_800,N_830);
or U935 (N_935,N_843,N_819);
nand U936 (N_936,N_840,N_889);
nand U937 (N_937,N_862,N_813);
and U938 (N_938,N_807,N_814);
or U939 (N_939,N_860,N_809);
or U940 (N_940,N_878,N_808);
or U941 (N_941,N_811,N_818);
or U942 (N_942,N_894,N_863);
nor U943 (N_943,N_858,N_880);
or U944 (N_944,N_888,N_885);
and U945 (N_945,N_866,N_829);
or U946 (N_946,N_844,N_839);
and U947 (N_947,N_806,N_891);
or U948 (N_948,N_898,N_873);
nor U949 (N_949,N_867,N_815);
nor U950 (N_950,N_843,N_844);
or U951 (N_951,N_871,N_877);
or U952 (N_952,N_859,N_842);
or U953 (N_953,N_837,N_823);
nand U954 (N_954,N_880,N_897);
nor U955 (N_955,N_888,N_891);
nor U956 (N_956,N_897,N_852);
or U957 (N_957,N_805,N_803);
and U958 (N_958,N_893,N_812);
nand U959 (N_959,N_895,N_882);
nor U960 (N_960,N_845,N_833);
nand U961 (N_961,N_874,N_888);
or U962 (N_962,N_811,N_890);
nor U963 (N_963,N_844,N_818);
nor U964 (N_964,N_834,N_805);
and U965 (N_965,N_846,N_820);
nand U966 (N_966,N_880,N_830);
nor U967 (N_967,N_829,N_816);
nor U968 (N_968,N_827,N_814);
nor U969 (N_969,N_827,N_864);
nand U970 (N_970,N_835,N_812);
or U971 (N_971,N_898,N_889);
and U972 (N_972,N_888,N_823);
nor U973 (N_973,N_898,N_835);
and U974 (N_974,N_806,N_872);
or U975 (N_975,N_842,N_896);
and U976 (N_976,N_816,N_874);
nor U977 (N_977,N_890,N_830);
nor U978 (N_978,N_862,N_860);
or U979 (N_979,N_861,N_889);
or U980 (N_980,N_888,N_886);
nor U981 (N_981,N_889,N_877);
nor U982 (N_982,N_820,N_818);
or U983 (N_983,N_882,N_834);
nor U984 (N_984,N_859,N_892);
nor U985 (N_985,N_859,N_855);
nand U986 (N_986,N_807,N_834);
or U987 (N_987,N_859,N_860);
nand U988 (N_988,N_892,N_880);
nand U989 (N_989,N_858,N_865);
nand U990 (N_990,N_822,N_838);
nor U991 (N_991,N_863,N_812);
and U992 (N_992,N_816,N_864);
nand U993 (N_993,N_878,N_807);
or U994 (N_994,N_898,N_803);
or U995 (N_995,N_819,N_876);
and U996 (N_996,N_870,N_801);
and U997 (N_997,N_808,N_861);
and U998 (N_998,N_820,N_869);
or U999 (N_999,N_805,N_883);
nor U1000 (N_1000,N_945,N_961);
nor U1001 (N_1001,N_902,N_968);
nor U1002 (N_1002,N_924,N_977);
nand U1003 (N_1003,N_931,N_900);
and U1004 (N_1004,N_957,N_989);
nor U1005 (N_1005,N_998,N_903);
or U1006 (N_1006,N_986,N_951);
and U1007 (N_1007,N_978,N_935);
or U1008 (N_1008,N_904,N_948);
and U1009 (N_1009,N_907,N_939);
nor U1010 (N_1010,N_991,N_925);
nor U1011 (N_1011,N_912,N_954);
and U1012 (N_1012,N_938,N_901);
nand U1013 (N_1013,N_930,N_949);
nor U1014 (N_1014,N_990,N_956);
and U1015 (N_1015,N_987,N_959);
and U1016 (N_1016,N_965,N_985);
nor U1017 (N_1017,N_974,N_932);
and U1018 (N_1018,N_972,N_967);
or U1019 (N_1019,N_958,N_993);
nand U1020 (N_1020,N_955,N_909);
xnor U1021 (N_1021,N_992,N_919);
nor U1022 (N_1022,N_914,N_941);
or U1023 (N_1023,N_973,N_952);
nand U1024 (N_1024,N_934,N_969);
and U1025 (N_1025,N_996,N_975);
nand U1026 (N_1026,N_908,N_927);
or U1027 (N_1027,N_971,N_984);
and U1028 (N_1028,N_918,N_950);
or U1029 (N_1029,N_940,N_979);
nand U1030 (N_1030,N_983,N_933);
and U1031 (N_1031,N_923,N_929);
and U1032 (N_1032,N_966,N_916);
or U1033 (N_1033,N_910,N_982);
or U1034 (N_1034,N_917,N_981);
and U1035 (N_1035,N_905,N_988);
nand U1036 (N_1036,N_928,N_937);
nand U1037 (N_1037,N_994,N_920);
or U1038 (N_1038,N_922,N_964);
or U1039 (N_1039,N_936,N_976);
or U1040 (N_1040,N_980,N_947);
nand U1041 (N_1041,N_943,N_963);
xnor U1042 (N_1042,N_960,N_921);
or U1043 (N_1043,N_942,N_999);
or U1044 (N_1044,N_911,N_995);
or U1045 (N_1045,N_997,N_962);
nand U1046 (N_1046,N_913,N_946);
nor U1047 (N_1047,N_970,N_944);
and U1048 (N_1048,N_926,N_915);
nand U1049 (N_1049,N_953,N_906);
and U1050 (N_1050,N_995,N_966);
or U1051 (N_1051,N_930,N_993);
nand U1052 (N_1052,N_944,N_903);
nor U1053 (N_1053,N_975,N_977);
or U1054 (N_1054,N_988,N_968);
nand U1055 (N_1055,N_905,N_971);
nor U1056 (N_1056,N_946,N_916);
nor U1057 (N_1057,N_958,N_964);
and U1058 (N_1058,N_999,N_956);
nor U1059 (N_1059,N_916,N_967);
or U1060 (N_1060,N_936,N_908);
or U1061 (N_1061,N_934,N_922);
and U1062 (N_1062,N_994,N_956);
nand U1063 (N_1063,N_943,N_926);
and U1064 (N_1064,N_950,N_965);
nor U1065 (N_1065,N_987,N_967);
or U1066 (N_1066,N_993,N_943);
or U1067 (N_1067,N_941,N_952);
or U1068 (N_1068,N_907,N_925);
or U1069 (N_1069,N_954,N_969);
nor U1070 (N_1070,N_971,N_989);
or U1071 (N_1071,N_906,N_905);
and U1072 (N_1072,N_979,N_994);
nor U1073 (N_1073,N_981,N_907);
and U1074 (N_1074,N_946,N_945);
nor U1075 (N_1075,N_988,N_996);
and U1076 (N_1076,N_988,N_961);
or U1077 (N_1077,N_951,N_999);
or U1078 (N_1078,N_905,N_941);
and U1079 (N_1079,N_987,N_912);
nor U1080 (N_1080,N_947,N_953);
nor U1081 (N_1081,N_999,N_914);
nand U1082 (N_1082,N_996,N_971);
nor U1083 (N_1083,N_960,N_989);
nand U1084 (N_1084,N_954,N_956);
nand U1085 (N_1085,N_970,N_912);
nand U1086 (N_1086,N_989,N_962);
nand U1087 (N_1087,N_918,N_949);
and U1088 (N_1088,N_919,N_991);
or U1089 (N_1089,N_944,N_908);
nor U1090 (N_1090,N_910,N_930);
nand U1091 (N_1091,N_924,N_965);
and U1092 (N_1092,N_986,N_988);
nand U1093 (N_1093,N_962,N_906);
and U1094 (N_1094,N_938,N_998);
nor U1095 (N_1095,N_925,N_922);
nor U1096 (N_1096,N_931,N_961);
nand U1097 (N_1097,N_980,N_956);
nor U1098 (N_1098,N_912,N_917);
nor U1099 (N_1099,N_962,N_978);
and U1100 (N_1100,N_1045,N_1014);
nor U1101 (N_1101,N_1054,N_1028);
and U1102 (N_1102,N_1005,N_1034);
or U1103 (N_1103,N_1077,N_1060);
nand U1104 (N_1104,N_1010,N_1013);
and U1105 (N_1105,N_1074,N_1071);
xnor U1106 (N_1106,N_1050,N_1059);
or U1107 (N_1107,N_1058,N_1092);
nand U1108 (N_1108,N_1020,N_1062);
nor U1109 (N_1109,N_1035,N_1007);
and U1110 (N_1110,N_1085,N_1066);
nor U1111 (N_1111,N_1022,N_1097);
nor U1112 (N_1112,N_1027,N_1069);
and U1113 (N_1113,N_1011,N_1082);
or U1114 (N_1114,N_1078,N_1099);
nand U1115 (N_1115,N_1033,N_1038);
nor U1116 (N_1116,N_1008,N_1090);
nor U1117 (N_1117,N_1006,N_1023);
and U1118 (N_1118,N_1041,N_1031);
nand U1119 (N_1119,N_1009,N_1075);
and U1120 (N_1120,N_1000,N_1021);
and U1121 (N_1121,N_1056,N_1043);
or U1122 (N_1122,N_1055,N_1076);
and U1123 (N_1123,N_1080,N_1088);
nand U1124 (N_1124,N_1002,N_1095);
and U1125 (N_1125,N_1040,N_1089);
nand U1126 (N_1126,N_1086,N_1019);
and U1127 (N_1127,N_1037,N_1098);
and U1128 (N_1128,N_1091,N_1003);
and U1129 (N_1129,N_1015,N_1083);
or U1130 (N_1130,N_1029,N_1026);
or U1131 (N_1131,N_1096,N_1064);
and U1132 (N_1132,N_1017,N_1044);
nand U1133 (N_1133,N_1052,N_1065);
nor U1134 (N_1134,N_1063,N_1061);
nor U1135 (N_1135,N_1084,N_1081);
or U1136 (N_1136,N_1024,N_1036);
nand U1137 (N_1137,N_1072,N_1042);
nand U1138 (N_1138,N_1032,N_1068);
or U1139 (N_1139,N_1004,N_1001);
nand U1140 (N_1140,N_1025,N_1047);
and U1141 (N_1141,N_1070,N_1053);
nor U1142 (N_1142,N_1051,N_1046);
or U1143 (N_1143,N_1094,N_1073);
nor U1144 (N_1144,N_1057,N_1039);
nor U1145 (N_1145,N_1067,N_1030);
nand U1146 (N_1146,N_1079,N_1093);
nand U1147 (N_1147,N_1012,N_1016);
nor U1148 (N_1148,N_1049,N_1048);
or U1149 (N_1149,N_1018,N_1087);
nor U1150 (N_1150,N_1060,N_1086);
nand U1151 (N_1151,N_1028,N_1091);
or U1152 (N_1152,N_1012,N_1075);
nor U1153 (N_1153,N_1035,N_1032);
nor U1154 (N_1154,N_1008,N_1065);
nor U1155 (N_1155,N_1016,N_1096);
and U1156 (N_1156,N_1056,N_1079);
nor U1157 (N_1157,N_1074,N_1093);
nor U1158 (N_1158,N_1014,N_1010);
or U1159 (N_1159,N_1092,N_1008);
or U1160 (N_1160,N_1024,N_1069);
and U1161 (N_1161,N_1096,N_1085);
or U1162 (N_1162,N_1020,N_1071);
nor U1163 (N_1163,N_1073,N_1028);
nand U1164 (N_1164,N_1095,N_1086);
and U1165 (N_1165,N_1078,N_1034);
and U1166 (N_1166,N_1082,N_1030);
and U1167 (N_1167,N_1027,N_1033);
or U1168 (N_1168,N_1048,N_1081);
xor U1169 (N_1169,N_1056,N_1069);
and U1170 (N_1170,N_1089,N_1085);
nor U1171 (N_1171,N_1007,N_1068);
nor U1172 (N_1172,N_1028,N_1050);
nand U1173 (N_1173,N_1050,N_1045);
or U1174 (N_1174,N_1041,N_1069);
nand U1175 (N_1175,N_1067,N_1021);
and U1176 (N_1176,N_1074,N_1063);
or U1177 (N_1177,N_1098,N_1083);
or U1178 (N_1178,N_1084,N_1020);
and U1179 (N_1179,N_1021,N_1088);
or U1180 (N_1180,N_1049,N_1065);
or U1181 (N_1181,N_1010,N_1091);
nand U1182 (N_1182,N_1039,N_1023);
xor U1183 (N_1183,N_1033,N_1076);
or U1184 (N_1184,N_1042,N_1068);
and U1185 (N_1185,N_1046,N_1003);
or U1186 (N_1186,N_1097,N_1021);
nand U1187 (N_1187,N_1061,N_1045);
or U1188 (N_1188,N_1019,N_1031);
or U1189 (N_1189,N_1078,N_1028);
nand U1190 (N_1190,N_1010,N_1031);
nand U1191 (N_1191,N_1096,N_1030);
nor U1192 (N_1192,N_1003,N_1063);
and U1193 (N_1193,N_1015,N_1086);
or U1194 (N_1194,N_1052,N_1068);
nand U1195 (N_1195,N_1064,N_1013);
or U1196 (N_1196,N_1008,N_1075);
or U1197 (N_1197,N_1011,N_1034);
nor U1198 (N_1198,N_1010,N_1093);
nor U1199 (N_1199,N_1058,N_1088);
or U1200 (N_1200,N_1198,N_1194);
nor U1201 (N_1201,N_1112,N_1152);
or U1202 (N_1202,N_1115,N_1185);
nor U1203 (N_1203,N_1147,N_1168);
nand U1204 (N_1204,N_1195,N_1182);
nand U1205 (N_1205,N_1102,N_1101);
and U1206 (N_1206,N_1190,N_1163);
nand U1207 (N_1207,N_1193,N_1135);
nor U1208 (N_1208,N_1129,N_1188);
or U1209 (N_1209,N_1142,N_1110);
xnor U1210 (N_1210,N_1122,N_1113);
nor U1211 (N_1211,N_1145,N_1196);
or U1212 (N_1212,N_1128,N_1106);
nor U1213 (N_1213,N_1159,N_1133);
nand U1214 (N_1214,N_1107,N_1109);
nand U1215 (N_1215,N_1164,N_1170);
and U1216 (N_1216,N_1178,N_1160);
nor U1217 (N_1217,N_1121,N_1184);
or U1218 (N_1218,N_1166,N_1123);
or U1219 (N_1219,N_1179,N_1161);
nor U1220 (N_1220,N_1119,N_1100);
and U1221 (N_1221,N_1156,N_1181);
or U1222 (N_1222,N_1180,N_1169);
nand U1223 (N_1223,N_1162,N_1132);
or U1224 (N_1224,N_1105,N_1199);
or U1225 (N_1225,N_1146,N_1117);
nor U1226 (N_1226,N_1144,N_1171);
or U1227 (N_1227,N_1165,N_1150);
nand U1228 (N_1228,N_1143,N_1148);
nor U1229 (N_1229,N_1176,N_1191);
nand U1230 (N_1230,N_1155,N_1139);
nand U1231 (N_1231,N_1154,N_1158);
and U1232 (N_1232,N_1103,N_1136);
nand U1233 (N_1233,N_1104,N_1149);
nand U1234 (N_1234,N_1174,N_1189);
nand U1235 (N_1235,N_1172,N_1134);
nand U1236 (N_1236,N_1131,N_1124);
nand U1237 (N_1237,N_1108,N_1186);
and U1238 (N_1238,N_1167,N_1137);
and U1239 (N_1239,N_1111,N_1126);
nand U1240 (N_1240,N_1157,N_1116);
and U1241 (N_1241,N_1153,N_1120);
nand U1242 (N_1242,N_1183,N_1175);
nor U1243 (N_1243,N_1118,N_1192);
nor U1244 (N_1244,N_1125,N_1177);
nand U1245 (N_1245,N_1138,N_1151);
nand U1246 (N_1246,N_1114,N_1140);
or U1247 (N_1247,N_1130,N_1127);
and U1248 (N_1248,N_1173,N_1187);
nand U1249 (N_1249,N_1197,N_1141);
nand U1250 (N_1250,N_1120,N_1186);
nand U1251 (N_1251,N_1137,N_1132);
nand U1252 (N_1252,N_1108,N_1139);
nand U1253 (N_1253,N_1171,N_1164);
nor U1254 (N_1254,N_1153,N_1162);
nand U1255 (N_1255,N_1148,N_1186);
nand U1256 (N_1256,N_1166,N_1142);
or U1257 (N_1257,N_1133,N_1148);
and U1258 (N_1258,N_1133,N_1196);
xnor U1259 (N_1259,N_1176,N_1151);
nand U1260 (N_1260,N_1116,N_1169);
or U1261 (N_1261,N_1130,N_1157);
and U1262 (N_1262,N_1116,N_1195);
or U1263 (N_1263,N_1120,N_1142);
nand U1264 (N_1264,N_1151,N_1188);
nor U1265 (N_1265,N_1113,N_1152);
and U1266 (N_1266,N_1137,N_1134);
xnor U1267 (N_1267,N_1156,N_1123);
nor U1268 (N_1268,N_1140,N_1135);
nor U1269 (N_1269,N_1140,N_1155);
nand U1270 (N_1270,N_1173,N_1160);
or U1271 (N_1271,N_1138,N_1118);
nand U1272 (N_1272,N_1193,N_1188);
and U1273 (N_1273,N_1193,N_1164);
nor U1274 (N_1274,N_1132,N_1187);
nor U1275 (N_1275,N_1118,N_1191);
or U1276 (N_1276,N_1135,N_1134);
nand U1277 (N_1277,N_1123,N_1196);
and U1278 (N_1278,N_1169,N_1143);
nor U1279 (N_1279,N_1161,N_1125);
nand U1280 (N_1280,N_1161,N_1166);
or U1281 (N_1281,N_1115,N_1146);
or U1282 (N_1282,N_1115,N_1151);
nand U1283 (N_1283,N_1102,N_1142);
nor U1284 (N_1284,N_1116,N_1192);
nor U1285 (N_1285,N_1168,N_1153);
and U1286 (N_1286,N_1140,N_1180);
nand U1287 (N_1287,N_1153,N_1188);
nor U1288 (N_1288,N_1173,N_1105);
nor U1289 (N_1289,N_1191,N_1127);
nand U1290 (N_1290,N_1170,N_1106);
nor U1291 (N_1291,N_1135,N_1123);
or U1292 (N_1292,N_1136,N_1167);
nand U1293 (N_1293,N_1139,N_1128);
nor U1294 (N_1294,N_1141,N_1104);
nand U1295 (N_1295,N_1139,N_1158);
nand U1296 (N_1296,N_1147,N_1169);
nor U1297 (N_1297,N_1183,N_1166);
and U1298 (N_1298,N_1141,N_1109);
or U1299 (N_1299,N_1193,N_1132);
nor U1300 (N_1300,N_1221,N_1239);
nor U1301 (N_1301,N_1251,N_1207);
and U1302 (N_1302,N_1258,N_1272);
nand U1303 (N_1303,N_1255,N_1231);
nor U1304 (N_1304,N_1241,N_1277);
or U1305 (N_1305,N_1252,N_1278);
nor U1306 (N_1306,N_1284,N_1237);
or U1307 (N_1307,N_1286,N_1238);
nand U1308 (N_1308,N_1204,N_1254);
and U1309 (N_1309,N_1240,N_1280);
nand U1310 (N_1310,N_1244,N_1215);
nand U1311 (N_1311,N_1216,N_1271);
or U1312 (N_1312,N_1213,N_1225);
nor U1313 (N_1313,N_1297,N_1208);
and U1314 (N_1314,N_1218,N_1253);
and U1315 (N_1315,N_1201,N_1222);
and U1316 (N_1316,N_1220,N_1275);
nand U1317 (N_1317,N_1269,N_1230);
or U1318 (N_1318,N_1203,N_1268);
and U1319 (N_1319,N_1288,N_1282);
nor U1320 (N_1320,N_1212,N_1266);
and U1321 (N_1321,N_1287,N_1246);
nor U1322 (N_1322,N_1223,N_1293);
or U1323 (N_1323,N_1205,N_1295);
or U1324 (N_1324,N_1298,N_1233);
nand U1325 (N_1325,N_1226,N_1290);
nor U1326 (N_1326,N_1292,N_1267);
or U1327 (N_1327,N_1200,N_1262);
nand U1328 (N_1328,N_1210,N_1211);
nand U1329 (N_1329,N_1265,N_1285);
nand U1330 (N_1330,N_1264,N_1256);
nand U1331 (N_1331,N_1219,N_1234);
or U1332 (N_1332,N_1281,N_1279);
or U1333 (N_1333,N_1242,N_1243);
or U1334 (N_1334,N_1235,N_1236);
or U1335 (N_1335,N_1299,N_1248);
nand U1336 (N_1336,N_1206,N_1232);
and U1337 (N_1337,N_1289,N_1250);
nand U1338 (N_1338,N_1217,N_1247);
nand U1339 (N_1339,N_1283,N_1270);
nand U1340 (N_1340,N_1273,N_1227);
nor U1341 (N_1341,N_1229,N_1224);
nand U1342 (N_1342,N_1276,N_1214);
nand U1343 (N_1343,N_1209,N_1249);
and U1344 (N_1344,N_1260,N_1228);
nand U1345 (N_1345,N_1202,N_1296);
nor U1346 (N_1346,N_1294,N_1263);
nand U1347 (N_1347,N_1291,N_1274);
and U1348 (N_1348,N_1245,N_1257);
and U1349 (N_1349,N_1259,N_1261);
nand U1350 (N_1350,N_1273,N_1225);
and U1351 (N_1351,N_1207,N_1289);
nor U1352 (N_1352,N_1275,N_1290);
and U1353 (N_1353,N_1218,N_1245);
nand U1354 (N_1354,N_1221,N_1291);
or U1355 (N_1355,N_1248,N_1200);
and U1356 (N_1356,N_1246,N_1249);
nor U1357 (N_1357,N_1280,N_1208);
nor U1358 (N_1358,N_1248,N_1219);
nor U1359 (N_1359,N_1211,N_1274);
or U1360 (N_1360,N_1292,N_1209);
nor U1361 (N_1361,N_1296,N_1207);
nand U1362 (N_1362,N_1260,N_1211);
nor U1363 (N_1363,N_1290,N_1230);
nor U1364 (N_1364,N_1234,N_1249);
and U1365 (N_1365,N_1263,N_1237);
nand U1366 (N_1366,N_1228,N_1241);
nand U1367 (N_1367,N_1205,N_1280);
and U1368 (N_1368,N_1283,N_1244);
nand U1369 (N_1369,N_1263,N_1256);
nand U1370 (N_1370,N_1281,N_1291);
or U1371 (N_1371,N_1201,N_1280);
or U1372 (N_1372,N_1209,N_1248);
and U1373 (N_1373,N_1200,N_1284);
and U1374 (N_1374,N_1247,N_1205);
nor U1375 (N_1375,N_1276,N_1205);
nand U1376 (N_1376,N_1203,N_1265);
nor U1377 (N_1377,N_1284,N_1278);
and U1378 (N_1378,N_1263,N_1261);
nand U1379 (N_1379,N_1224,N_1299);
or U1380 (N_1380,N_1235,N_1225);
and U1381 (N_1381,N_1208,N_1296);
and U1382 (N_1382,N_1252,N_1286);
and U1383 (N_1383,N_1267,N_1261);
nor U1384 (N_1384,N_1230,N_1256);
or U1385 (N_1385,N_1295,N_1209);
or U1386 (N_1386,N_1213,N_1269);
nand U1387 (N_1387,N_1287,N_1258);
nor U1388 (N_1388,N_1263,N_1234);
nand U1389 (N_1389,N_1296,N_1227);
nand U1390 (N_1390,N_1210,N_1247);
or U1391 (N_1391,N_1228,N_1280);
and U1392 (N_1392,N_1202,N_1282);
nand U1393 (N_1393,N_1208,N_1268);
and U1394 (N_1394,N_1215,N_1241);
xnor U1395 (N_1395,N_1267,N_1211);
nand U1396 (N_1396,N_1294,N_1200);
and U1397 (N_1397,N_1252,N_1276);
xnor U1398 (N_1398,N_1205,N_1231);
nand U1399 (N_1399,N_1201,N_1200);
and U1400 (N_1400,N_1361,N_1396);
xnor U1401 (N_1401,N_1359,N_1328);
nand U1402 (N_1402,N_1362,N_1302);
and U1403 (N_1403,N_1356,N_1379);
nor U1404 (N_1404,N_1397,N_1332);
nand U1405 (N_1405,N_1307,N_1347);
nor U1406 (N_1406,N_1335,N_1330);
and U1407 (N_1407,N_1375,N_1370);
nand U1408 (N_1408,N_1314,N_1366);
nand U1409 (N_1409,N_1349,N_1331);
or U1410 (N_1410,N_1334,N_1371);
or U1411 (N_1411,N_1309,N_1390);
nand U1412 (N_1412,N_1344,N_1369);
nand U1413 (N_1413,N_1348,N_1394);
and U1414 (N_1414,N_1385,N_1322);
or U1415 (N_1415,N_1360,N_1311);
nor U1416 (N_1416,N_1382,N_1377);
and U1417 (N_1417,N_1373,N_1319);
or U1418 (N_1418,N_1387,N_1372);
xnor U1419 (N_1419,N_1383,N_1345);
nor U1420 (N_1420,N_1323,N_1381);
and U1421 (N_1421,N_1395,N_1368);
nor U1422 (N_1422,N_1399,N_1312);
and U1423 (N_1423,N_1324,N_1315);
nor U1424 (N_1424,N_1310,N_1300);
nand U1425 (N_1425,N_1355,N_1318);
nor U1426 (N_1426,N_1343,N_1374);
and U1427 (N_1427,N_1380,N_1376);
or U1428 (N_1428,N_1350,N_1325);
nand U1429 (N_1429,N_1389,N_1320);
or U1430 (N_1430,N_1316,N_1303);
and U1431 (N_1431,N_1354,N_1308);
nand U1432 (N_1432,N_1327,N_1329);
nor U1433 (N_1433,N_1386,N_1306);
nand U1434 (N_1434,N_1358,N_1367);
nand U1435 (N_1435,N_1321,N_1336);
or U1436 (N_1436,N_1353,N_1338);
and U1437 (N_1437,N_1313,N_1365);
or U1438 (N_1438,N_1305,N_1342);
or U1439 (N_1439,N_1384,N_1364);
and U1440 (N_1440,N_1341,N_1363);
or U1441 (N_1441,N_1391,N_1301);
nand U1442 (N_1442,N_1398,N_1339);
and U1443 (N_1443,N_1333,N_1351);
nor U1444 (N_1444,N_1346,N_1317);
nor U1445 (N_1445,N_1352,N_1378);
or U1446 (N_1446,N_1340,N_1392);
or U1447 (N_1447,N_1388,N_1393);
and U1448 (N_1448,N_1337,N_1357);
or U1449 (N_1449,N_1304,N_1326);
and U1450 (N_1450,N_1343,N_1314);
nand U1451 (N_1451,N_1303,N_1370);
and U1452 (N_1452,N_1334,N_1390);
or U1453 (N_1453,N_1303,N_1336);
nand U1454 (N_1454,N_1381,N_1371);
or U1455 (N_1455,N_1399,N_1324);
or U1456 (N_1456,N_1330,N_1355);
or U1457 (N_1457,N_1355,N_1356);
or U1458 (N_1458,N_1331,N_1321);
nor U1459 (N_1459,N_1355,N_1373);
and U1460 (N_1460,N_1319,N_1311);
nand U1461 (N_1461,N_1316,N_1344);
and U1462 (N_1462,N_1300,N_1324);
or U1463 (N_1463,N_1365,N_1366);
or U1464 (N_1464,N_1380,N_1379);
nand U1465 (N_1465,N_1357,N_1327);
nand U1466 (N_1466,N_1330,N_1332);
nor U1467 (N_1467,N_1375,N_1369);
and U1468 (N_1468,N_1391,N_1312);
nor U1469 (N_1469,N_1376,N_1300);
or U1470 (N_1470,N_1379,N_1307);
or U1471 (N_1471,N_1333,N_1397);
nand U1472 (N_1472,N_1398,N_1389);
nand U1473 (N_1473,N_1343,N_1369);
nor U1474 (N_1474,N_1314,N_1342);
and U1475 (N_1475,N_1374,N_1346);
nand U1476 (N_1476,N_1309,N_1301);
and U1477 (N_1477,N_1341,N_1370);
or U1478 (N_1478,N_1356,N_1361);
or U1479 (N_1479,N_1337,N_1334);
nand U1480 (N_1480,N_1345,N_1366);
or U1481 (N_1481,N_1376,N_1342);
nand U1482 (N_1482,N_1326,N_1309);
nor U1483 (N_1483,N_1341,N_1343);
nor U1484 (N_1484,N_1326,N_1394);
or U1485 (N_1485,N_1313,N_1361);
xnor U1486 (N_1486,N_1383,N_1354);
xnor U1487 (N_1487,N_1345,N_1378);
and U1488 (N_1488,N_1332,N_1305);
nor U1489 (N_1489,N_1324,N_1398);
and U1490 (N_1490,N_1301,N_1371);
nor U1491 (N_1491,N_1395,N_1330);
or U1492 (N_1492,N_1393,N_1350);
or U1493 (N_1493,N_1327,N_1318);
and U1494 (N_1494,N_1343,N_1388);
nand U1495 (N_1495,N_1365,N_1314);
nand U1496 (N_1496,N_1341,N_1394);
nand U1497 (N_1497,N_1372,N_1373);
nor U1498 (N_1498,N_1353,N_1397);
nor U1499 (N_1499,N_1342,N_1322);
nand U1500 (N_1500,N_1487,N_1413);
and U1501 (N_1501,N_1495,N_1483);
or U1502 (N_1502,N_1451,N_1467);
nor U1503 (N_1503,N_1411,N_1440);
nand U1504 (N_1504,N_1432,N_1447);
nand U1505 (N_1505,N_1499,N_1464);
and U1506 (N_1506,N_1473,N_1416);
nand U1507 (N_1507,N_1409,N_1421);
or U1508 (N_1508,N_1491,N_1446);
and U1509 (N_1509,N_1482,N_1492);
and U1510 (N_1510,N_1434,N_1458);
or U1511 (N_1511,N_1450,N_1488);
nand U1512 (N_1512,N_1459,N_1405);
nand U1513 (N_1513,N_1497,N_1470);
or U1514 (N_1514,N_1493,N_1402);
or U1515 (N_1515,N_1478,N_1449);
and U1516 (N_1516,N_1417,N_1455);
and U1517 (N_1517,N_1429,N_1474);
nor U1518 (N_1518,N_1476,N_1453);
or U1519 (N_1519,N_1438,N_1481);
or U1520 (N_1520,N_1433,N_1424);
and U1521 (N_1521,N_1456,N_1466);
or U1522 (N_1522,N_1400,N_1454);
nand U1523 (N_1523,N_1475,N_1498);
nor U1524 (N_1524,N_1419,N_1472);
and U1525 (N_1525,N_1463,N_1457);
nand U1526 (N_1526,N_1496,N_1418);
nor U1527 (N_1527,N_1445,N_1403);
nor U1528 (N_1528,N_1414,N_1431);
or U1529 (N_1529,N_1435,N_1443);
and U1530 (N_1530,N_1422,N_1460);
or U1531 (N_1531,N_1426,N_1439);
nor U1532 (N_1532,N_1479,N_1462);
and U1533 (N_1533,N_1410,N_1437);
nand U1534 (N_1534,N_1404,N_1477);
nor U1535 (N_1535,N_1494,N_1427);
or U1536 (N_1536,N_1452,N_1412);
nor U1537 (N_1537,N_1425,N_1468);
or U1538 (N_1538,N_1480,N_1415);
or U1539 (N_1539,N_1465,N_1489);
or U1540 (N_1540,N_1461,N_1436);
or U1541 (N_1541,N_1420,N_1406);
nor U1542 (N_1542,N_1408,N_1471);
nor U1543 (N_1543,N_1423,N_1430);
nand U1544 (N_1544,N_1448,N_1490);
or U1545 (N_1545,N_1407,N_1484);
nand U1546 (N_1546,N_1428,N_1441);
nor U1547 (N_1547,N_1485,N_1486);
nor U1548 (N_1548,N_1401,N_1444);
nor U1549 (N_1549,N_1442,N_1469);
or U1550 (N_1550,N_1477,N_1461);
nor U1551 (N_1551,N_1452,N_1489);
nor U1552 (N_1552,N_1454,N_1422);
or U1553 (N_1553,N_1498,N_1473);
or U1554 (N_1554,N_1484,N_1434);
nand U1555 (N_1555,N_1437,N_1482);
and U1556 (N_1556,N_1447,N_1413);
or U1557 (N_1557,N_1471,N_1475);
nor U1558 (N_1558,N_1407,N_1471);
or U1559 (N_1559,N_1437,N_1402);
nor U1560 (N_1560,N_1474,N_1496);
and U1561 (N_1561,N_1472,N_1408);
and U1562 (N_1562,N_1490,N_1489);
or U1563 (N_1563,N_1448,N_1443);
or U1564 (N_1564,N_1431,N_1439);
nor U1565 (N_1565,N_1472,N_1442);
nand U1566 (N_1566,N_1447,N_1451);
or U1567 (N_1567,N_1478,N_1404);
and U1568 (N_1568,N_1495,N_1423);
or U1569 (N_1569,N_1416,N_1463);
nor U1570 (N_1570,N_1443,N_1446);
nand U1571 (N_1571,N_1470,N_1427);
nor U1572 (N_1572,N_1463,N_1473);
or U1573 (N_1573,N_1441,N_1477);
and U1574 (N_1574,N_1496,N_1412);
and U1575 (N_1575,N_1423,N_1461);
nand U1576 (N_1576,N_1404,N_1430);
nand U1577 (N_1577,N_1493,N_1451);
or U1578 (N_1578,N_1416,N_1436);
nand U1579 (N_1579,N_1463,N_1407);
and U1580 (N_1580,N_1401,N_1441);
nor U1581 (N_1581,N_1421,N_1437);
nor U1582 (N_1582,N_1416,N_1467);
and U1583 (N_1583,N_1405,N_1429);
nand U1584 (N_1584,N_1480,N_1445);
nor U1585 (N_1585,N_1418,N_1457);
and U1586 (N_1586,N_1408,N_1494);
nand U1587 (N_1587,N_1418,N_1405);
nor U1588 (N_1588,N_1443,N_1419);
or U1589 (N_1589,N_1479,N_1421);
nor U1590 (N_1590,N_1478,N_1470);
or U1591 (N_1591,N_1459,N_1485);
nor U1592 (N_1592,N_1414,N_1450);
and U1593 (N_1593,N_1436,N_1422);
nand U1594 (N_1594,N_1480,N_1490);
and U1595 (N_1595,N_1444,N_1480);
and U1596 (N_1596,N_1470,N_1484);
nand U1597 (N_1597,N_1483,N_1463);
nor U1598 (N_1598,N_1485,N_1458);
nand U1599 (N_1599,N_1451,N_1477);
or U1600 (N_1600,N_1580,N_1586);
or U1601 (N_1601,N_1588,N_1564);
or U1602 (N_1602,N_1510,N_1542);
nor U1603 (N_1603,N_1515,N_1535);
nor U1604 (N_1604,N_1512,N_1598);
and U1605 (N_1605,N_1562,N_1554);
nor U1606 (N_1606,N_1579,N_1563);
or U1607 (N_1607,N_1590,N_1573);
and U1608 (N_1608,N_1571,N_1560);
and U1609 (N_1609,N_1575,N_1544);
nor U1610 (N_1610,N_1524,N_1525);
and U1611 (N_1611,N_1578,N_1561);
and U1612 (N_1612,N_1589,N_1584);
nand U1613 (N_1613,N_1540,N_1595);
nand U1614 (N_1614,N_1568,N_1550);
or U1615 (N_1615,N_1519,N_1514);
and U1616 (N_1616,N_1551,N_1527);
and U1617 (N_1617,N_1532,N_1511);
or U1618 (N_1618,N_1577,N_1518);
and U1619 (N_1619,N_1558,N_1592);
nor U1620 (N_1620,N_1506,N_1509);
or U1621 (N_1621,N_1530,N_1537);
or U1622 (N_1622,N_1557,N_1520);
nor U1623 (N_1623,N_1502,N_1545);
and U1624 (N_1624,N_1576,N_1565);
or U1625 (N_1625,N_1599,N_1533);
and U1626 (N_1626,N_1596,N_1553);
or U1627 (N_1627,N_1529,N_1543);
nand U1628 (N_1628,N_1591,N_1523);
or U1629 (N_1629,N_1521,N_1594);
or U1630 (N_1630,N_1556,N_1526);
or U1631 (N_1631,N_1513,N_1503);
nand U1632 (N_1632,N_1559,N_1539);
and U1633 (N_1633,N_1581,N_1534);
and U1634 (N_1634,N_1574,N_1507);
nand U1635 (N_1635,N_1528,N_1508);
nor U1636 (N_1636,N_1567,N_1522);
or U1637 (N_1637,N_1546,N_1504);
and U1638 (N_1638,N_1531,N_1548);
or U1639 (N_1639,N_1597,N_1547);
or U1640 (N_1640,N_1500,N_1569);
nor U1641 (N_1641,N_1570,N_1582);
nand U1642 (N_1642,N_1517,N_1587);
xnor U1643 (N_1643,N_1555,N_1585);
nand U1644 (N_1644,N_1583,N_1572);
nor U1645 (N_1645,N_1549,N_1541);
or U1646 (N_1646,N_1538,N_1593);
or U1647 (N_1647,N_1501,N_1505);
nor U1648 (N_1648,N_1552,N_1566);
or U1649 (N_1649,N_1516,N_1536);
nand U1650 (N_1650,N_1539,N_1540);
xor U1651 (N_1651,N_1546,N_1560);
nand U1652 (N_1652,N_1529,N_1533);
and U1653 (N_1653,N_1590,N_1578);
or U1654 (N_1654,N_1557,N_1594);
nor U1655 (N_1655,N_1530,N_1557);
and U1656 (N_1656,N_1506,N_1561);
nor U1657 (N_1657,N_1528,N_1536);
nand U1658 (N_1658,N_1504,N_1575);
nor U1659 (N_1659,N_1535,N_1505);
xor U1660 (N_1660,N_1523,N_1567);
nand U1661 (N_1661,N_1588,N_1500);
and U1662 (N_1662,N_1548,N_1580);
nor U1663 (N_1663,N_1596,N_1539);
and U1664 (N_1664,N_1527,N_1504);
nor U1665 (N_1665,N_1511,N_1571);
or U1666 (N_1666,N_1588,N_1586);
or U1667 (N_1667,N_1597,N_1509);
and U1668 (N_1668,N_1551,N_1510);
or U1669 (N_1669,N_1552,N_1567);
and U1670 (N_1670,N_1575,N_1582);
nand U1671 (N_1671,N_1546,N_1567);
nor U1672 (N_1672,N_1590,N_1562);
and U1673 (N_1673,N_1552,N_1575);
and U1674 (N_1674,N_1534,N_1597);
or U1675 (N_1675,N_1533,N_1587);
or U1676 (N_1676,N_1587,N_1535);
or U1677 (N_1677,N_1552,N_1539);
and U1678 (N_1678,N_1519,N_1543);
nand U1679 (N_1679,N_1582,N_1549);
and U1680 (N_1680,N_1562,N_1571);
nor U1681 (N_1681,N_1569,N_1542);
nor U1682 (N_1682,N_1556,N_1552);
nand U1683 (N_1683,N_1516,N_1511);
or U1684 (N_1684,N_1595,N_1510);
and U1685 (N_1685,N_1583,N_1567);
or U1686 (N_1686,N_1553,N_1509);
and U1687 (N_1687,N_1585,N_1528);
or U1688 (N_1688,N_1531,N_1572);
nand U1689 (N_1689,N_1522,N_1538);
nor U1690 (N_1690,N_1579,N_1547);
or U1691 (N_1691,N_1505,N_1595);
nor U1692 (N_1692,N_1551,N_1547);
and U1693 (N_1693,N_1588,N_1515);
or U1694 (N_1694,N_1517,N_1573);
nor U1695 (N_1695,N_1507,N_1575);
nor U1696 (N_1696,N_1538,N_1511);
and U1697 (N_1697,N_1500,N_1521);
and U1698 (N_1698,N_1588,N_1558);
nand U1699 (N_1699,N_1590,N_1530);
and U1700 (N_1700,N_1634,N_1665);
and U1701 (N_1701,N_1627,N_1682);
nand U1702 (N_1702,N_1604,N_1631);
nand U1703 (N_1703,N_1690,N_1698);
nor U1704 (N_1704,N_1629,N_1656);
or U1705 (N_1705,N_1681,N_1676);
or U1706 (N_1706,N_1619,N_1680);
or U1707 (N_1707,N_1638,N_1697);
or U1708 (N_1708,N_1671,N_1670);
nor U1709 (N_1709,N_1688,N_1605);
xnor U1710 (N_1710,N_1679,N_1639);
and U1711 (N_1711,N_1614,N_1612);
and U1712 (N_1712,N_1641,N_1600);
and U1713 (N_1713,N_1657,N_1613);
or U1714 (N_1714,N_1695,N_1643);
nor U1715 (N_1715,N_1636,N_1608);
nor U1716 (N_1716,N_1622,N_1646);
nand U1717 (N_1717,N_1696,N_1632);
or U1718 (N_1718,N_1610,N_1694);
nor U1719 (N_1719,N_1642,N_1699);
and U1720 (N_1720,N_1675,N_1677);
or U1721 (N_1721,N_1635,N_1616);
nand U1722 (N_1722,N_1658,N_1652);
nand U1723 (N_1723,N_1689,N_1691);
nand U1724 (N_1724,N_1630,N_1687);
nor U1725 (N_1725,N_1692,N_1645);
nand U1726 (N_1726,N_1668,N_1623);
nand U1727 (N_1727,N_1662,N_1603);
nand U1728 (N_1728,N_1674,N_1659);
nor U1729 (N_1729,N_1649,N_1661);
nor U1730 (N_1730,N_1683,N_1669);
or U1731 (N_1731,N_1611,N_1609);
nand U1732 (N_1732,N_1655,N_1625);
nand U1733 (N_1733,N_1628,N_1606);
or U1734 (N_1734,N_1648,N_1647);
and U1735 (N_1735,N_1644,N_1640);
and U1736 (N_1736,N_1693,N_1621);
and U1737 (N_1737,N_1654,N_1653);
nand U1738 (N_1738,N_1664,N_1602);
nand U1739 (N_1739,N_1620,N_1660);
nand U1740 (N_1740,N_1651,N_1673);
or U1741 (N_1741,N_1663,N_1684);
or U1742 (N_1742,N_1667,N_1601);
nor U1743 (N_1743,N_1617,N_1618);
or U1744 (N_1744,N_1672,N_1615);
nand U1745 (N_1745,N_1633,N_1666);
or U1746 (N_1746,N_1686,N_1607);
or U1747 (N_1747,N_1637,N_1624);
nor U1748 (N_1748,N_1678,N_1685);
nand U1749 (N_1749,N_1626,N_1650);
xor U1750 (N_1750,N_1639,N_1615);
and U1751 (N_1751,N_1638,N_1627);
nor U1752 (N_1752,N_1640,N_1696);
or U1753 (N_1753,N_1633,N_1600);
or U1754 (N_1754,N_1660,N_1679);
nor U1755 (N_1755,N_1686,N_1629);
and U1756 (N_1756,N_1658,N_1604);
nor U1757 (N_1757,N_1679,N_1671);
and U1758 (N_1758,N_1691,N_1652);
and U1759 (N_1759,N_1626,N_1619);
or U1760 (N_1760,N_1600,N_1670);
nor U1761 (N_1761,N_1699,N_1679);
or U1762 (N_1762,N_1664,N_1657);
or U1763 (N_1763,N_1601,N_1612);
nand U1764 (N_1764,N_1620,N_1616);
nor U1765 (N_1765,N_1623,N_1657);
or U1766 (N_1766,N_1656,N_1663);
nand U1767 (N_1767,N_1685,N_1669);
or U1768 (N_1768,N_1642,N_1661);
nand U1769 (N_1769,N_1684,N_1672);
nor U1770 (N_1770,N_1686,N_1685);
or U1771 (N_1771,N_1620,N_1692);
nor U1772 (N_1772,N_1610,N_1638);
nand U1773 (N_1773,N_1649,N_1636);
or U1774 (N_1774,N_1614,N_1609);
nor U1775 (N_1775,N_1679,N_1625);
nand U1776 (N_1776,N_1638,N_1674);
nand U1777 (N_1777,N_1602,N_1617);
nor U1778 (N_1778,N_1624,N_1678);
nor U1779 (N_1779,N_1660,N_1623);
or U1780 (N_1780,N_1611,N_1625);
nand U1781 (N_1781,N_1645,N_1690);
and U1782 (N_1782,N_1617,N_1623);
nor U1783 (N_1783,N_1672,N_1642);
and U1784 (N_1784,N_1684,N_1611);
xnor U1785 (N_1785,N_1643,N_1688);
nor U1786 (N_1786,N_1608,N_1675);
nand U1787 (N_1787,N_1600,N_1645);
nand U1788 (N_1788,N_1647,N_1620);
and U1789 (N_1789,N_1605,N_1658);
nor U1790 (N_1790,N_1669,N_1607);
nor U1791 (N_1791,N_1694,N_1660);
nand U1792 (N_1792,N_1691,N_1623);
nand U1793 (N_1793,N_1650,N_1668);
and U1794 (N_1794,N_1636,N_1630);
nand U1795 (N_1795,N_1642,N_1669);
or U1796 (N_1796,N_1699,N_1696);
nor U1797 (N_1797,N_1651,N_1601);
or U1798 (N_1798,N_1671,N_1632);
or U1799 (N_1799,N_1657,N_1637);
or U1800 (N_1800,N_1780,N_1758);
xor U1801 (N_1801,N_1790,N_1742);
and U1802 (N_1802,N_1760,N_1772);
and U1803 (N_1803,N_1717,N_1770);
nand U1804 (N_1804,N_1749,N_1778);
nor U1805 (N_1805,N_1748,N_1730);
or U1806 (N_1806,N_1714,N_1737);
and U1807 (N_1807,N_1769,N_1765);
nand U1808 (N_1808,N_1719,N_1729);
and U1809 (N_1809,N_1783,N_1756);
or U1810 (N_1810,N_1745,N_1740);
nor U1811 (N_1811,N_1736,N_1784);
and U1812 (N_1812,N_1789,N_1757);
and U1813 (N_1813,N_1726,N_1715);
or U1814 (N_1814,N_1732,N_1773);
nor U1815 (N_1815,N_1766,N_1799);
nand U1816 (N_1816,N_1753,N_1791);
nor U1817 (N_1817,N_1703,N_1702);
nor U1818 (N_1818,N_1767,N_1762);
or U1819 (N_1819,N_1711,N_1704);
nor U1820 (N_1820,N_1768,N_1779);
or U1821 (N_1821,N_1793,N_1727);
nor U1822 (N_1822,N_1716,N_1755);
or U1823 (N_1823,N_1733,N_1752);
nor U1824 (N_1824,N_1731,N_1771);
nand U1825 (N_1825,N_1792,N_1777);
and U1826 (N_1826,N_1735,N_1787);
and U1827 (N_1827,N_1746,N_1759);
nor U1828 (N_1828,N_1738,N_1744);
nand U1829 (N_1829,N_1734,N_1797);
and U1830 (N_1830,N_1705,N_1710);
or U1831 (N_1831,N_1796,N_1798);
nand U1832 (N_1832,N_1713,N_1782);
xor U1833 (N_1833,N_1712,N_1786);
and U1834 (N_1834,N_1718,N_1725);
nand U1835 (N_1835,N_1728,N_1761);
and U1836 (N_1836,N_1764,N_1774);
nand U1837 (N_1837,N_1776,N_1739);
and U1838 (N_1838,N_1721,N_1788);
and U1839 (N_1839,N_1750,N_1708);
nand U1840 (N_1840,N_1795,N_1775);
nor U1841 (N_1841,N_1722,N_1707);
or U1842 (N_1842,N_1751,N_1743);
and U1843 (N_1843,N_1754,N_1724);
nor U1844 (N_1844,N_1720,N_1785);
and U1845 (N_1845,N_1763,N_1701);
nand U1846 (N_1846,N_1794,N_1741);
and U1847 (N_1847,N_1781,N_1709);
or U1848 (N_1848,N_1700,N_1706);
nor U1849 (N_1849,N_1723,N_1747);
and U1850 (N_1850,N_1705,N_1723);
nor U1851 (N_1851,N_1748,N_1783);
nand U1852 (N_1852,N_1766,N_1764);
or U1853 (N_1853,N_1708,N_1779);
or U1854 (N_1854,N_1724,N_1744);
or U1855 (N_1855,N_1783,N_1774);
nand U1856 (N_1856,N_1750,N_1714);
or U1857 (N_1857,N_1783,N_1708);
or U1858 (N_1858,N_1765,N_1784);
and U1859 (N_1859,N_1735,N_1729);
or U1860 (N_1860,N_1704,N_1762);
and U1861 (N_1861,N_1748,N_1777);
nand U1862 (N_1862,N_1774,N_1706);
and U1863 (N_1863,N_1758,N_1719);
xor U1864 (N_1864,N_1764,N_1751);
nand U1865 (N_1865,N_1761,N_1700);
and U1866 (N_1866,N_1705,N_1728);
or U1867 (N_1867,N_1726,N_1750);
or U1868 (N_1868,N_1743,N_1790);
nor U1869 (N_1869,N_1756,N_1705);
nor U1870 (N_1870,N_1749,N_1741);
and U1871 (N_1871,N_1789,N_1704);
nor U1872 (N_1872,N_1747,N_1791);
nor U1873 (N_1873,N_1710,N_1722);
and U1874 (N_1874,N_1726,N_1751);
and U1875 (N_1875,N_1706,N_1776);
or U1876 (N_1876,N_1735,N_1737);
nand U1877 (N_1877,N_1762,N_1742);
or U1878 (N_1878,N_1786,N_1777);
or U1879 (N_1879,N_1742,N_1771);
nor U1880 (N_1880,N_1702,N_1785);
or U1881 (N_1881,N_1758,N_1755);
nand U1882 (N_1882,N_1771,N_1788);
or U1883 (N_1883,N_1734,N_1714);
and U1884 (N_1884,N_1706,N_1770);
nor U1885 (N_1885,N_1729,N_1772);
nand U1886 (N_1886,N_1754,N_1730);
or U1887 (N_1887,N_1718,N_1757);
nor U1888 (N_1888,N_1739,N_1760);
and U1889 (N_1889,N_1744,N_1705);
nand U1890 (N_1890,N_1749,N_1768);
nor U1891 (N_1891,N_1757,N_1717);
nand U1892 (N_1892,N_1779,N_1772);
and U1893 (N_1893,N_1746,N_1770);
or U1894 (N_1894,N_1717,N_1753);
nor U1895 (N_1895,N_1754,N_1787);
or U1896 (N_1896,N_1723,N_1776);
nor U1897 (N_1897,N_1771,N_1758);
nor U1898 (N_1898,N_1773,N_1791);
nor U1899 (N_1899,N_1704,N_1792);
nor U1900 (N_1900,N_1871,N_1835);
and U1901 (N_1901,N_1837,N_1815);
and U1902 (N_1902,N_1842,N_1824);
or U1903 (N_1903,N_1847,N_1849);
nand U1904 (N_1904,N_1879,N_1851);
nand U1905 (N_1905,N_1858,N_1861);
nand U1906 (N_1906,N_1800,N_1892);
nor U1907 (N_1907,N_1897,N_1888);
and U1908 (N_1908,N_1802,N_1896);
nor U1909 (N_1909,N_1881,N_1829);
or U1910 (N_1910,N_1838,N_1865);
or U1911 (N_1911,N_1852,N_1878);
or U1912 (N_1912,N_1821,N_1809);
nor U1913 (N_1913,N_1883,N_1820);
nand U1914 (N_1914,N_1876,N_1813);
nand U1915 (N_1915,N_1827,N_1845);
nor U1916 (N_1916,N_1836,N_1886);
and U1917 (N_1917,N_1895,N_1808);
nor U1918 (N_1918,N_1859,N_1863);
nor U1919 (N_1919,N_1898,N_1823);
or U1920 (N_1920,N_1862,N_1833);
nand U1921 (N_1921,N_1812,N_1857);
and U1922 (N_1922,N_1814,N_1854);
nand U1923 (N_1923,N_1848,N_1828);
nor U1924 (N_1924,N_1855,N_1872);
or U1925 (N_1925,N_1834,N_1831);
and U1926 (N_1926,N_1846,N_1880);
or U1927 (N_1927,N_1843,N_1840);
nand U1928 (N_1928,N_1864,N_1841);
nand U1929 (N_1929,N_1819,N_1811);
nor U1930 (N_1930,N_1894,N_1850);
and U1931 (N_1931,N_1891,N_1869);
nand U1932 (N_1932,N_1885,N_1866);
nand U1933 (N_1933,N_1822,N_1804);
and U1934 (N_1934,N_1887,N_1817);
nor U1935 (N_1935,N_1884,N_1826);
and U1936 (N_1936,N_1873,N_1839);
or U1937 (N_1937,N_1818,N_1856);
or U1938 (N_1938,N_1807,N_1801);
nor U1939 (N_1939,N_1806,N_1874);
or U1940 (N_1940,N_1844,N_1810);
or U1941 (N_1941,N_1882,N_1893);
nor U1942 (N_1942,N_1853,N_1889);
and U1943 (N_1943,N_1867,N_1860);
nand U1944 (N_1944,N_1868,N_1816);
and U1945 (N_1945,N_1899,N_1832);
nand U1946 (N_1946,N_1875,N_1805);
nor U1947 (N_1947,N_1890,N_1830);
and U1948 (N_1948,N_1803,N_1870);
or U1949 (N_1949,N_1825,N_1877);
and U1950 (N_1950,N_1899,N_1827);
nor U1951 (N_1951,N_1847,N_1897);
and U1952 (N_1952,N_1893,N_1825);
nand U1953 (N_1953,N_1896,N_1820);
nor U1954 (N_1954,N_1822,N_1854);
and U1955 (N_1955,N_1803,N_1862);
nor U1956 (N_1956,N_1823,N_1838);
or U1957 (N_1957,N_1883,N_1868);
and U1958 (N_1958,N_1846,N_1838);
and U1959 (N_1959,N_1838,N_1857);
nand U1960 (N_1960,N_1839,N_1841);
nor U1961 (N_1961,N_1850,N_1821);
and U1962 (N_1962,N_1827,N_1877);
and U1963 (N_1963,N_1861,N_1851);
nand U1964 (N_1964,N_1875,N_1839);
or U1965 (N_1965,N_1804,N_1802);
and U1966 (N_1966,N_1812,N_1878);
nand U1967 (N_1967,N_1815,N_1851);
nand U1968 (N_1968,N_1870,N_1837);
or U1969 (N_1969,N_1867,N_1872);
nand U1970 (N_1970,N_1842,N_1819);
and U1971 (N_1971,N_1870,N_1898);
or U1972 (N_1972,N_1887,N_1897);
or U1973 (N_1973,N_1814,N_1879);
nor U1974 (N_1974,N_1809,N_1818);
nor U1975 (N_1975,N_1836,N_1843);
and U1976 (N_1976,N_1870,N_1832);
or U1977 (N_1977,N_1817,N_1828);
and U1978 (N_1978,N_1890,N_1847);
and U1979 (N_1979,N_1824,N_1807);
nor U1980 (N_1980,N_1842,N_1840);
and U1981 (N_1981,N_1879,N_1880);
nor U1982 (N_1982,N_1887,N_1827);
nor U1983 (N_1983,N_1890,N_1807);
nor U1984 (N_1984,N_1863,N_1893);
or U1985 (N_1985,N_1804,N_1820);
and U1986 (N_1986,N_1802,N_1881);
nor U1987 (N_1987,N_1847,N_1879);
and U1988 (N_1988,N_1883,N_1889);
and U1989 (N_1989,N_1859,N_1882);
nor U1990 (N_1990,N_1891,N_1872);
xnor U1991 (N_1991,N_1843,N_1857);
and U1992 (N_1992,N_1890,N_1832);
nor U1993 (N_1993,N_1897,N_1832);
nand U1994 (N_1994,N_1864,N_1843);
nor U1995 (N_1995,N_1816,N_1886);
xor U1996 (N_1996,N_1808,N_1888);
and U1997 (N_1997,N_1863,N_1818);
and U1998 (N_1998,N_1840,N_1816);
nor U1999 (N_1999,N_1870,N_1894);
and U2000 (N_2000,N_1983,N_1964);
nor U2001 (N_2001,N_1940,N_1925);
and U2002 (N_2002,N_1961,N_1921);
and U2003 (N_2003,N_1965,N_1957);
or U2004 (N_2004,N_1912,N_1933);
nand U2005 (N_2005,N_1974,N_1929);
nand U2006 (N_2006,N_1942,N_1910);
and U2007 (N_2007,N_1950,N_1979);
and U2008 (N_2008,N_1996,N_1915);
nor U2009 (N_2009,N_1937,N_1911);
nand U2010 (N_2010,N_1984,N_1934);
or U2011 (N_2011,N_1938,N_1977);
nor U2012 (N_2012,N_1926,N_1995);
nor U2013 (N_2013,N_1902,N_1955);
nor U2014 (N_2014,N_1953,N_1907);
or U2015 (N_2015,N_1993,N_1956);
nand U2016 (N_2016,N_1903,N_1987);
nand U2017 (N_2017,N_1997,N_1927);
or U2018 (N_2018,N_1999,N_1905);
nor U2019 (N_2019,N_1988,N_1919);
nand U2020 (N_2020,N_1962,N_1917);
nand U2021 (N_2021,N_1949,N_1931);
nor U2022 (N_2022,N_1967,N_1948);
or U2023 (N_2023,N_1994,N_1951);
and U2024 (N_2024,N_1930,N_1980);
nor U2025 (N_2025,N_1991,N_1981);
nor U2026 (N_2026,N_1990,N_1900);
and U2027 (N_2027,N_1963,N_1992);
nand U2028 (N_2028,N_1906,N_1928);
nand U2029 (N_2029,N_1909,N_1944);
nand U2030 (N_2030,N_1901,N_1914);
nand U2031 (N_2031,N_1932,N_1976);
nor U2032 (N_2032,N_1972,N_1978);
and U2033 (N_2033,N_1998,N_1952);
nor U2034 (N_2034,N_1924,N_1986);
nand U2035 (N_2035,N_1941,N_1947);
and U2036 (N_2036,N_1973,N_1935);
nand U2037 (N_2037,N_1939,N_1982);
nor U2038 (N_2038,N_1985,N_1975);
and U2039 (N_2039,N_1954,N_1918);
nand U2040 (N_2040,N_1904,N_1971);
nand U2041 (N_2041,N_1968,N_1946);
xnor U2042 (N_2042,N_1960,N_1922);
nor U2043 (N_2043,N_1936,N_1966);
or U2044 (N_2044,N_1970,N_1959);
and U2045 (N_2045,N_1945,N_1958);
nor U2046 (N_2046,N_1908,N_1943);
or U2047 (N_2047,N_1989,N_1916);
nand U2048 (N_2048,N_1913,N_1920);
nand U2049 (N_2049,N_1969,N_1923);
and U2050 (N_2050,N_1902,N_1910);
and U2051 (N_2051,N_1918,N_1958);
or U2052 (N_2052,N_1991,N_1941);
or U2053 (N_2053,N_1941,N_1970);
or U2054 (N_2054,N_1926,N_1990);
nand U2055 (N_2055,N_1916,N_1990);
nand U2056 (N_2056,N_1937,N_1993);
and U2057 (N_2057,N_1935,N_1944);
and U2058 (N_2058,N_1902,N_1913);
or U2059 (N_2059,N_1904,N_1945);
nor U2060 (N_2060,N_1942,N_1906);
and U2061 (N_2061,N_1953,N_1966);
and U2062 (N_2062,N_1931,N_1919);
nand U2063 (N_2063,N_1989,N_1975);
and U2064 (N_2064,N_1906,N_1959);
nand U2065 (N_2065,N_1903,N_1958);
nor U2066 (N_2066,N_1979,N_1953);
and U2067 (N_2067,N_1983,N_1922);
nand U2068 (N_2068,N_1913,N_1915);
or U2069 (N_2069,N_1990,N_1907);
and U2070 (N_2070,N_1960,N_1929);
and U2071 (N_2071,N_1994,N_1903);
nand U2072 (N_2072,N_1979,N_1997);
or U2073 (N_2073,N_1941,N_1939);
or U2074 (N_2074,N_1953,N_1959);
or U2075 (N_2075,N_1915,N_1906);
and U2076 (N_2076,N_1916,N_1904);
nand U2077 (N_2077,N_1988,N_1936);
nor U2078 (N_2078,N_1927,N_1920);
and U2079 (N_2079,N_1937,N_1995);
or U2080 (N_2080,N_1945,N_1932);
nor U2081 (N_2081,N_1962,N_1969);
nor U2082 (N_2082,N_1931,N_1956);
and U2083 (N_2083,N_1918,N_1936);
and U2084 (N_2084,N_1988,N_1984);
nand U2085 (N_2085,N_1953,N_1976);
nand U2086 (N_2086,N_1975,N_1910);
or U2087 (N_2087,N_1947,N_1902);
nand U2088 (N_2088,N_1999,N_1904);
nand U2089 (N_2089,N_1911,N_1934);
and U2090 (N_2090,N_1972,N_1987);
nand U2091 (N_2091,N_1953,N_1949);
nand U2092 (N_2092,N_1951,N_1911);
nand U2093 (N_2093,N_1983,N_1906);
nand U2094 (N_2094,N_1980,N_1918);
nor U2095 (N_2095,N_1996,N_1929);
nor U2096 (N_2096,N_1955,N_1986);
xor U2097 (N_2097,N_1908,N_1903);
nor U2098 (N_2098,N_1961,N_1903);
or U2099 (N_2099,N_1980,N_1965);
or U2100 (N_2100,N_2046,N_2018);
and U2101 (N_2101,N_2082,N_2033);
nand U2102 (N_2102,N_2050,N_2080);
and U2103 (N_2103,N_2006,N_2067);
nor U2104 (N_2104,N_2026,N_2072);
nor U2105 (N_2105,N_2055,N_2058);
nand U2106 (N_2106,N_2030,N_2049);
and U2107 (N_2107,N_2066,N_2071);
or U2108 (N_2108,N_2073,N_2008);
and U2109 (N_2109,N_2028,N_2098);
nor U2110 (N_2110,N_2007,N_2031);
nor U2111 (N_2111,N_2012,N_2069);
nor U2112 (N_2112,N_2086,N_2019);
or U2113 (N_2113,N_2083,N_2005);
and U2114 (N_2114,N_2078,N_2063);
and U2115 (N_2115,N_2087,N_2035);
nand U2116 (N_2116,N_2088,N_2037);
nand U2117 (N_2117,N_2045,N_2014);
nand U2118 (N_2118,N_2084,N_2032);
xor U2119 (N_2119,N_2016,N_2054);
and U2120 (N_2120,N_2023,N_2094);
and U2121 (N_2121,N_2074,N_2051);
and U2122 (N_2122,N_2043,N_2089);
nor U2123 (N_2123,N_2060,N_2097);
nand U2124 (N_2124,N_2081,N_2021);
or U2125 (N_2125,N_2011,N_2062);
xnor U2126 (N_2126,N_2053,N_2009);
or U2127 (N_2127,N_2002,N_2027);
or U2128 (N_2128,N_2047,N_2039);
and U2129 (N_2129,N_2024,N_2076);
nor U2130 (N_2130,N_2079,N_2052);
nand U2131 (N_2131,N_2059,N_2095);
or U2132 (N_2132,N_2034,N_2000);
nand U2133 (N_2133,N_2003,N_2096);
or U2134 (N_2134,N_2022,N_2093);
and U2135 (N_2135,N_2036,N_2038);
nor U2136 (N_2136,N_2077,N_2013);
nand U2137 (N_2137,N_2099,N_2068);
and U2138 (N_2138,N_2001,N_2004);
nor U2139 (N_2139,N_2091,N_2041);
nand U2140 (N_2140,N_2065,N_2044);
or U2141 (N_2141,N_2085,N_2029);
nor U2142 (N_2142,N_2040,N_2092);
or U2143 (N_2143,N_2010,N_2090);
and U2144 (N_2144,N_2064,N_2017);
or U2145 (N_2145,N_2061,N_2025);
nand U2146 (N_2146,N_2042,N_2015);
nand U2147 (N_2147,N_2075,N_2070);
xnor U2148 (N_2148,N_2048,N_2057);
nand U2149 (N_2149,N_2056,N_2020);
nor U2150 (N_2150,N_2047,N_2060);
nand U2151 (N_2151,N_2041,N_2060);
nor U2152 (N_2152,N_2039,N_2012);
nand U2153 (N_2153,N_2073,N_2042);
or U2154 (N_2154,N_2067,N_2097);
nor U2155 (N_2155,N_2085,N_2075);
and U2156 (N_2156,N_2005,N_2073);
or U2157 (N_2157,N_2026,N_2053);
and U2158 (N_2158,N_2039,N_2051);
or U2159 (N_2159,N_2005,N_2011);
nor U2160 (N_2160,N_2050,N_2054);
or U2161 (N_2161,N_2016,N_2070);
or U2162 (N_2162,N_2021,N_2093);
or U2163 (N_2163,N_2090,N_2022);
or U2164 (N_2164,N_2079,N_2075);
and U2165 (N_2165,N_2061,N_2071);
nand U2166 (N_2166,N_2006,N_2076);
nand U2167 (N_2167,N_2051,N_2023);
nor U2168 (N_2168,N_2052,N_2065);
and U2169 (N_2169,N_2040,N_2039);
or U2170 (N_2170,N_2046,N_2083);
and U2171 (N_2171,N_2067,N_2017);
and U2172 (N_2172,N_2066,N_2074);
nand U2173 (N_2173,N_2098,N_2054);
xor U2174 (N_2174,N_2048,N_2086);
nor U2175 (N_2175,N_2001,N_2070);
nand U2176 (N_2176,N_2054,N_2066);
nor U2177 (N_2177,N_2010,N_2085);
and U2178 (N_2178,N_2022,N_2079);
nand U2179 (N_2179,N_2041,N_2067);
nand U2180 (N_2180,N_2029,N_2019);
nand U2181 (N_2181,N_2081,N_2075);
nor U2182 (N_2182,N_2040,N_2099);
or U2183 (N_2183,N_2075,N_2033);
nor U2184 (N_2184,N_2010,N_2059);
nand U2185 (N_2185,N_2040,N_2047);
or U2186 (N_2186,N_2027,N_2073);
and U2187 (N_2187,N_2015,N_2049);
or U2188 (N_2188,N_2043,N_2051);
nand U2189 (N_2189,N_2006,N_2099);
or U2190 (N_2190,N_2055,N_2065);
and U2191 (N_2191,N_2032,N_2090);
or U2192 (N_2192,N_2086,N_2097);
nor U2193 (N_2193,N_2035,N_2050);
and U2194 (N_2194,N_2063,N_2020);
nand U2195 (N_2195,N_2054,N_2056);
and U2196 (N_2196,N_2096,N_2034);
and U2197 (N_2197,N_2034,N_2061);
or U2198 (N_2198,N_2041,N_2055);
and U2199 (N_2199,N_2088,N_2071);
or U2200 (N_2200,N_2115,N_2188);
and U2201 (N_2201,N_2177,N_2175);
or U2202 (N_2202,N_2113,N_2185);
nand U2203 (N_2203,N_2184,N_2157);
nor U2204 (N_2204,N_2171,N_2196);
nor U2205 (N_2205,N_2139,N_2160);
or U2206 (N_2206,N_2126,N_2194);
nor U2207 (N_2207,N_2152,N_2192);
nand U2208 (N_2208,N_2125,N_2140);
nand U2209 (N_2209,N_2101,N_2150);
nor U2210 (N_2210,N_2151,N_2114);
nand U2211 (N_2211,N_2165,N_2195);
or U2212 (N_2212,N_2121,N_2166);
nand U2213 (N_2213,N_2102,N_2111);
nand U2214 (N_2214,N_2147,N_2168);
and U2215 (N_2215,N_2190,N_2162);
nor U2216 (N_2216,N_2135,N_2183);
nand U2217 (N_2217,N_2136,N_2138);
nor U2218 (N_2218,N_2134,N_2180);
nor U2219 (N_2219,N_2143,N_2104);
nor U2220 (N_2220,N_2187,N_2119);
nand U2221 (N_2221,N_2129,N_2176);
nor U2222 (N_2222,N_2169,N_2178);
nor U2223 (N_2223,N_2182,N_2193);
or U2224 (N_2224,N_2112,N_2120);
and U2225 (N_2225,N_2145,N_2132);
nor U2226 (N_2226,N_2164,N_2161);
nand U2227 (N_2227,N_2133,N_2103);
and U2228 (N_2228,N_2197,N_2153);
nand U2229 (N_2229,N_2156,N_2148);
nand U2230 (N_2230,N_2141,N_2186);
or U2231 (N_2231,N_2149,N_2172);
or U2232 (N_2232,N_2117,N_2105);
nand U2233 (N_2233,N_2154,N_2198);
and U2234 (N_2234,N_2118,N_2124);
and U2235 (N_2235,N_2181,N_2106);
nand U2236 (N_2236,N_2110,N_2130);
nor U2237 (N_2237,N_2100,N_2142);
nor U2238 (N_2238,N_2199,N_2128);
nor U2239 (N_2239,N_2173,N_2144);
or U2240 (N_2240,N_2158,N_2107);
nand U2241 (N_2241,N_2179,N_2137);
nor U2242 (N_2242,N_2163,N_2191);
nor U2243 (N_2243,N_2109,N_2167);
and U2244 (N_2244,N_2174,N_2122);
nor U2245 (N_2245,N_2146,N_2189);
nand U2246 (N_2246,N_2127,N_2108);
nor U2247 (N_2247,N_2155,N_2159);
nor U2248 (N_2248,N_2170,N_2131);
and U2249 (N_2249,N_2116,N_2123);
nor U2250 (N_2250,N_2123,N_2176);
and U2251 (N_2251,N_2142,N_2193);
or U2252 (N_2252,N_2194,N_2129);
nor U2253 (N_2253,N_2152,N_2189);
nor U2254 (N_2254,N_2166,N_2156);
and U2255 (N_2255,N_2182,N_2197);
and U2256 (N_2256,N_2165,N_2190);
nor U2257 (N_2257,N_2148,N_2149);
nand U2258 (N_2258,N_2107,N_2111);
or U2259 (N_2259,N_2159,N_2133);
nand U2260 (N_2260,N_2107,N_2149);
nand U2261 (N_2261,N_2196,N_2161);
nand U2262 (N_2262,N_2135,N_2127);
and U2263 (N_2263,N_2186,N_2190);
or U2264 (N_2264,N_2109,N_2156);
and U2265 (N_2265,N_2189,N_2149);
nand U2266 (N_2266,N_2164,N_2132);
and U2267 (N_2267,N_2132,N_2156);
nand U2268 (N_2268,N_2199,N_2193);
and U2269 (N_2269,N_2115,N_2135);
or U2270 (N_2270,N_2183,N_2115);
nand U2271 (N_2271,N_2130,N_2122);
nand U2272 (N_2272,N_2123,N_2186);
nor U2273 (N_2273,N_2111,N_2135);
or U2274 (N_2274,N_2139,N_2178);
or U2275 (N_2275,N_2103,N_2140);
nand U2276 (N_2276,N_2131,N_2145);
nor U2277 (N_2277,N_2194,N_2111);
or U2278 (N_2278,N_2130,N_2106);
or U2279 (N_2279,N_2174,N_2193);
or U2280 (N_2280,N_2195,N_2182);
nand U2281 (N_2281,N_2140,N_2143);
nor U2282 (N_2282,N_2181,N_2101);
nand U2283 (N_2283,N_2108,N_2147);
or U2284 (N_2284,N_2172,N_2168);
and U2285 (N_2285,N_2189,N_2103);
nor U2286 (N_2286,N_2171,N_2197);
or U2287 (N_2287,N_2100,N_2195);
and U2288 (N_2288,N_2188,N_2181);
nand U2289 (N_2289,N_2136,N_2102);
nor U2290 (N_2290,N_2135,N_2116);
and U2291 (N_2291,N_2105,N_2190);
nor U2292 (N_2292,N_2131,N_2189);
nand U2293 (N_2293,N_2167,N_2134);
nand U2294 (N_2294,N_2178,N_2122);
or U2295 (N_2295,N_2124,N_2155);
or U2296 (N_2296,N_2183,N_2104);
and U2297 (N_2297,N_2192,N_2120);
or U2298 (N_2298,N_2116,N_2160);
or U2299 (N_2299,N_2107,N_2164);
or U2300 (N_2300,N_2283,N_2258);
and U2301 (N_2301,N_2231,N_2282);
nand U2302 (N_2302,N_2277,N_2223);
nor U2303 (N_2303,N_2217,N_2244);
and U2304 (N_2304,N_2238,N_2284);
or U2305 (N_2305,N_2232,N_2260);
and U2306 (N_2306,N_2220,N_2264);
or U2307 (N_2307,N_2221,N_2270);
and U2308 (N_2308,N_2285,N_2255);
and U2309 (N_2309,N_2237,N_2214);
or U2310 (N_2310,N_2202,N_2215);
xnor U2311 (N_2311,N_2204,N_2261);
or U2312 (N_2312,N_2286,N_2248);
nand U2313 (N_2313,N_2265,N_2250);
or U2314 (N_2314,N_2245,N_2252);
nand U2315 (N_2315,N_2299,N_2256);
or U2316 (N_2316,N_2266,N_2227);
nand U2317 (N_2317,N_2254,N_2276);
nor U2318 (N_2318,N_2210,N_2251);
nand U2319 (N_2319,N_2236,N_2280);
or U2320 (N_2320,N_2262,N_2200);
or U2321 (N_2321,N_2208,N_2212);
nor U2322 (N_2322,N_2239,N_2281);
nand U2323 (N_2323,N_2267,N_2201);
or U2324 (N_2324,N_2293,N_2297);
nor U2325 (N_2325,N_2218,N_2230);
nor U2326 (N_2326,N_2290,N_2288);
or U2327 (N_2327,N_2203,N_2213);
nand U2328 (N_2328,N_2224,N_2211);
nor U2329 (N_2329,N_2219,N_2226);
nand U2330 (N_2330,N_2234,N_2249);
and U2331 (N_2331,N_2205,N_2207);
nand U2332 (N_2332,N_2206,N_2259);
nand U2333 (N_2333,N_2287,N_2272);
and U2334 (N_2334,N_2243,N_2228);
or U2335 (N_2335,N_2296,N_2257);
or U2336 (N_2336,N_2298,N_2225);
nand U2337 (N_2337,N_2246,N_2229);
nor U2338 (N_2338,N_2273,N_2235);
nand U2339 (N_2339,N_2271,N_2269);
nor U2340 (N_2340,N_2253,N_2268);
nand U2341 (N_2341,N_2247,N_2291);
and U2342 (N_2342,N_2275,N_2292);
and U2343 (N_2343,N_2278,N_2295);
xnor U2344 (N_2344,N_2289,N_2222);
nand U2345 (N_2345,N_2279,N_2241);
xor U2346 (N_2346,N_2294,N_2240);
nor U2347 (N_2347,N_2216,N_2233);
or U2348 (N_2348,N_2242,N_2263);
nor U2349 (N_2349,N_2209,N_2274);
nor U2350 (N_2350,N_2242,N_2218);
nand U2351 (N_2351,N_2215,N_2276);
nand U2352 (N_2352,N_2288,N_2275);
nand U2353 (N_2353,N_2284,N_2206);
nand U2354 (N_2354,N_2211,N_2271);
or U2355 (N_2355,N_2229,N_2275);
and U2356 (N_2356,N_2226,N_2253);
nand U2357 (N_2357,N_2256,N_2252);
nand U2358 (N_2358,N_2229,N_2293);
nand U2359 (N_2359,N_2212,N_2205);
nand U2360 (N_2360,N_2261,N_2256);
or U2361 (N_2361,N_2209,N_2255);
or U2362 (N_2362,N_2205,N_2244);
nand U2363 (N_2363,N_2275,N_2298);
or U2364 (N_2364,N_2248,N_2283);
and U2365 (N_2365,N_2267,N_2243);
nor U2366 (N_2366,N_2298,N_2260);
nor U2367 (N_2367,N_2251,N_2288);
or U2368 (N_2368,N_2228,N_2292);
or U2369 (N_2369,N_2222,N_2234);
and U2370 (N_2370,N_2267,N_2265);
or U2371 (N_2371,N_2244,N_2294);
or U2372 (N_2372,N_2232,N_2268);
nand U2373 (N_2373,N_2237,N_2211);
and U2374 (N_2374,N_2282,N_2226);
nand U2375 (N_2375,N_2280,N_2230);
or U2376 (N_2376,N_2241,N_2265);
nand U2377 (N_2377,N_2288,N_2269);
nand U2378 (N_2378,N_2297,N_2288);
and U2379 (N_2379,N_2289,N_2248);
xor U2380 (N_2380,N_2260,N_2274);
and U2381 (N_2381,N_2202,N_2276);
nor U2382 (N_2382,N_2277,N_2219);
nand U2383 (N_2383,N_2282,N_2287);
or U2384 (N_2384,N_2270,N_2236);
or U2385 (N_2385,N_2215,N_2286);
and U2386 (N_2386,N_2291,N_2264);
or U2387 (N_2387,N_2221,N_2203);
nand U2388 (N_2388,N_2220,N_2200);
and U2389 (N_2389,N_2242,N_2291);
nand U2390 (N_2390,N_2237,N_2278);
and U2391 (N_2391,N_2205,N_2230);
nand U2392 (N_2392,N_2244,N_2254);
or U2393 (N_2393,N_2212,N_2297);
or U2394 (N_2394,N_2286,N_2268);
nand U2395 (N_2395,N_2293,N_2211);
nand U2396 (N_2396,N_2289,N_2247);
nor U2397 (N_2397,N_2225,N_2223);
nor U2398 (N_2398,N_2245,N_2255);
and U2399 (N_2399,N_2288,N_2202);
nand U2400 (N_2400,N_2320,N_2373);
or U2401 (N_2401,N_2348,N_2381);
or U2402 (N_2402,N_2333,N_2384);
nand U2403 (N_2403,N_2365,N_2380);
and U2404 (N_2404,N_2356,N_2395);
nor U2405 (N_2405,N_2353,N_2379);
and U2406 (N_2406,N_2351,N_2307);
xor U2407 (N_2407,N_2350,N_2327);
nor U2408 (N_2408,N_2300,N_2382);
nor U2409 (N_2409,N_2397,N_2367);
nor U2410 (N_2410,N_2352,N_2389);
and U2411 (N_2411,N_2363,N_2328);
or U2412 (N_2412,N_2383,N_2368);
nand U2413 (N_2413,N_2372,N_2360);
nand U2414 (N_2414,N_2309,N_2336);
nand U2415 (N_2415,N_2387,N_2334);
or U2416 (N_2416,N_2347,N_2325);
nand U2417 (N_2417,N_2326,N_2362);
nor U2418 (N_2418,N_2303,N_2331);
nand U2419 (N_2419,N_2302,N_2354);
nor U2420 (N_2420,N_2371,N_2345);
nand U2421 (N_2421,N_2310,N_2393);
and U2422 (N_2422,N_2340,N_2337);
or U2423 (N_2423,N_2330,N_2305);
or U2424 (N_2424,N_2304,N_2378);
and U2425 (N_2425,N_2306,N_2313);
nand U2426 (N_2426,N_2388,N_2358);
or U2427 (N_2427,N_2343,N_2359);
nand U2428 (N_2428,N_2369,N_2376);
nor U2429 (N_2429,N_2315,N_2385);
and U2430 (N_2430,N_2392,N_2366);
or U2431 (N_2431,N_2349,N_2391);
nand U2432 (N_2432,N_2386,N_2318);
nor U2433 (N_2433,N_2374,N_2312);
or U2434 (N_2434,N_2342,N_2341);
nand U2435 (N_2435,N_2332,N_2317);
or U2436 (N_2436,N_2399,N_2339);
nor U2437 (N_2437,N_2324,N_2390);
and U2438 (N_2438,N_2323,N_2329);
nand U2439 (N_2439,N_2346,N_2322);
nand U2440 (N_2440,N_2321,N_2355);
and U2441 (N_2441,N_2357,N_2370);
nand U2442 (N_2442,N_2311,N_2338);
nor U2443 (N_2443,N_2394,N_2377);
nor U2444 (N_2444,N_2319,N_2398);
and U2445 (N_2445,N_2335,N_2301);
xnor U2446 (N_2446,N_2316,N_2361);
and U2447 (N_2447,N_2344,N_2375);
nand U2448 (N_2448,N_2364,N_2308);
or U2449 (N_2449,N_2396,N_2314);
nor U2450 (N_2450,N_2380,N_2307);
or U2451 (N_2451,N_2372,N_2342);
or U2452 (N_2452,N_2320,N_2377);
or U2453 (N_2453,N_2363,N_2382);
or U2454 (N_2454,N_2325,N_2336);
or U2455 (N_2455,N_2391,N_2335);
and U2456 (N_2456,N_2379,N_2303);
or U2457 (N_2457,N_2368,N_2385);
and U2458 (N_2458,N_2368,N_2358);
nand U2459 (N_2459,N_2334,N_2322);
and U2460 (N_2460,N_2379,N_2307);
nor U2461 (N_2461,N_2351,N_2361);
nand U2462 (N_2462,N_2383,N_2336);
nand U2463 (N_2463,N_2334,N_2359);
xor U2464 (N_2464,N_2365,N_2301);
nor U2465 (N_2465,N_2318,N_2349);
nor U2466 (N_2466,N_2307,N_2399);
and U2467 (N_2467,N_2331,N_2333);
or U2468 (N_2468,N_2306,N_2346);
and U2469 (N_2469,N_2385,N_2389);
nor U2470 (N_2470,N_2367,N_2357);
nor U2471 (N_2471,N_2313,N_2359);
or U2472 (N_2472,N_2385,N_2388);
nor U2473 (N_2473,N_2341,N_2306);
nor U2474 (N_2474,N_2329,N_2332);
and U2475 (N_2475,N_2388,N_2312);
or U2476 (N_2476,N_2360,N_2387);
and U2477 (N_2477,N_2325,N_2303);
nor U2478 (N_2478,N_2370,N_2365);
nor U2479 (N_2479,N_2346,N_2335);
or U2480 (N_2480,N_2393,N_2390);
and U2481 (N_2481,N_2374,N_2340);
nor U2482 (N_2482,N_2309,N_2365);
nor U2483 (N_2483,N_2383,N_2366);
and U2484 (N_2484,N_2313,N_2341);
nand U2485 (N_2485,N_2343,N_2374);
and U2486 (N_2486,N_2339,N_2318);
or U2487 (N_2487,N_2305,N_2388);
nor U2488 (N_2488,N_2371,N_2362);
nor U2489 (N_2489,N_2301,N_2352);
or U2490 (N_2490,N_2302,N_2325);
nand U2491 (N_2491,N_2365,N_2310);
or U2492 (N_2492,N_2310,N_2348);
nand U2493 (N_2493,N_2315,N_2301);
nand U2494 (N_2494,N_2399,N_2337);
or U2495 (N_2495,N_2374,N_2359);
and U2496 (N_2496,N_2303,N_2382);
and U2497 (N_2497,N_2387,N_2369);
nand U2498 (N_2498,N_2387,N_2305);
or U2499 (N_2499,N_2397,N_2336);
and U2500 (N_2500,N_2490,N_2455);
nand U2501 (N_2501,N_2466,N_2419);
nand U2502 (N_2502,N_2489,N_2407);
nand U2503 (N_2503,N_2423,N_2408);
nor U2504 (N_2504,N_2422,N_2417);
nand U2505 (N_2505,N_2406,N_2413);
or U2506 (N_2506,N_2452,N_2410);
nand U2507 (N_2507,N_2404,N_2454);
or U2508 (N_2508,N_2480,N_2465);
nand U2509 (N_2509,N_2471,N_2497);
nor U2510 (N_2510,N_2459,N_2478);
and U2511 (N_2511,N_2446,N_2482);
nand U2512 (N_2512,N_2400,N_2424);
or U2513 (N_2513,N_2470,N_2418);
nand U2514 (N_2514,N_2428,N_2405);
nor U2515 (N_2515,N_2475,N_2439);
nand U2516 (N_2516,N_2484,N_2457);
and U2517 (N_2517,N_2412,N_2491);
nand U2518 (N_2518,N_2434,N_2421);
nand U2519 (N_2519,N_2473,N_2458);
nand U2520 (N_2520,N_2462,N_2479);
nor U2521 (N_2521,N_2453,N_2444);
and U2522 (N_2522,N_2450,N_2432);
and U2523 (N_2523,N_2415,N_2425);
or U2524 (N_2524,N_2441,N_2477);
nor U2525 (N_2525,N_2416,N_2445);
or U2526 (N_2526,N_2456,N_2488);
or U2527 (N_2527,N_2436,N_2483);
and U2528 (N_2528,N_2437,N_2487);
and U2529 (N_2529,N_2496,N_2427);
nor U2530 (N_2530,N_2440,N_2467);
or U2531 (N_2531,N_2414,N_2420);
nor U2532 (N_2532,N_2449,N_2433);
nor U2533 (N_2533,N_2468,N_2442);
and U2534 (N_2534,N_2429,N_2451);
nand U2535 (N_2535,N_2460,N_2426);
nor U2536 (N_2536,N_2499,N_2463);
nand U2537 (N_2537,N_2493,N_2435);
and U2538 (N_2538,N_2461,N_2492);
and U2539 (N_2539,N_2402,N_2495);
or U2540 (N_2540,N_2438,N_2430);
or U2541 (N_2541,N_2498,N_2474);
nor U2542 (N_2542,N_2472,N_2401);
and U2543 (N_2543,N_2485,N_2411);
nand U2544 (N_2544,N_2447,N_2476);
nor U2545 (N_2545,N_2486,N_2481);
or U2546 (N_2546,N_2494,N_2431);
or U2547 (N_2547,N_2469,N_2403);
or U2548 (N_2548,N_2448,N_2464);
nand U2549 (N_2549,N_2409,N_2443);
nor U2550 (N_2550,N_2479,N_2468);
nor U2551 (N_2551,N_2439,N_2412);
or U2552 (N_2552,N_2424,N_2440);
or U2553 (N_2553,N_2411,N_2469);
or U2554 (N_2554,N_2459,N_2407);
or U2555 (N_2555,N_2466,N_2468);
nor U2556 (N_2556,N_2418,N_2484);
nand U2557 (N_2557,N_2429,N_2420);
nor U2558 (N_2558,N_2406,N_2467);
or U2559 (N_2559,N_2489,N_2415);
and U2560 (N_2560,N_2415,N_2495);
nand U2561 (N_2561,N_2424,N_2466);
or U2562 (N_2562,N_2469,N_2483);
and U2563 (N_2563,N_2454,N_2406);
and U2564 (N_2564,N_2431,N_2463);
and U2565 (N_2565,N_2482,N_2477);
nor U2566 (N_2566,N_2483,N_2424);
nor U2567 (N_2567,N_2457,N_2416);
and U2568 (N_2568,N_2483,N_2403);
and U2569 (N_2569,N_2407,N_2430);
or U2570 (N_2570,N_2426,N_2479);
nor U2571 (N_2571,N_2423,N_2484);
nor U2572 (N_2572,N_2404,N_2471);
or U2573 (N_2573,N_2451,N_2434);
and U2574 (N_2574,N_2429,N_2441);
and U2575 (N_2575,N_2491,N_2498);
and U2576 (N_2576,N_2406,N_2430);
nor U2577 (N_2577,N_2477,N_2438);
or U2578 (N_2578,N_2487,N_2469);
or U2579 (N_2579,N_2412,N_2474);
or U2580 (N_2580,N_2411,N_2477);
nand U2581 (N_2581,N_2497,N_2467);
nand U2582 (N_2582,N_2458,N_2419);
and U2583 (N_2583,N_2477,N_2474);
or U2584 (N_2584,N_2401,N_2415);
and U2585 (N_2585,N_2473,N_2499);
or U2586 (N_2586,N_2481,N_2453);
nand U2587 (N_2587,N_2447,N_2410);
and U2588 (N_2588,N_2473,N_2437);
nor U2589 (N_2589,N_2496,N_2455);
and U2590 (N_2590,N_2433,N_2457);
nor U2591 (N_2591,N_2412,N_2488);
nand U2592 (N_2592,N_2429,N_2434);
and U2593 (N_2593,N_2458,N_2484);
and U2594 (N_2594,N_2453,N_2438);
or U2595 (N_2595,N_2494,N_2423);
nand U2596 (N_2596,N_2493,N_2438);
nor U2597 (N_2597,N_2411,N_2429);
nor U2598 (N_2598,N_2421,N_2481);
nor U2599 (N_2599,N_2475,N_2446);
nor U2600 (N_2600,N_2522,N_2559);
and U2601 (N_2601,N_2558,N_2526);
or U2602 (N_2602,N_2560,N_2553);
nand U2603 (N_2603,N_2568,N_2516);
nor U2604 (N_2604,N_2571,N_2535);
nand U2605 (N_2605,N_2500,N_2514);
and U2606 (N_2606,N_2504,N_2542);
and U2607 (N_2607,N_2590,N_2557);
nand U2608 (N_2608,N_2588,N_2589);
or U2609 (N_2609,N_2567,N_2544);
and U2610 (N_2610,N_2524,N_2531);
nor U2611 (N_2611,N_2538,N_2505);
xor U2612 (N_2612,N_2562,N_2579);
and U2613 (N_2613,N_2599,N_2595);
or U2614 (N_2614,N_2545,N_2597);
nand U2615 (N_2615,N_2541,N_2549);
or U2616 (N_2616,N_2528,N_2577);
nor U2617 (N_2617,N_2540,N_2585);
and U2618 (N_2618,N_2527,N_2591);
nor U2619 (N_2619,N_2561,N_2520);
nand U2620 (N_2620,N_2564,N_2525);
and U2621 (N_2621,N_2547,N_2569);
and U2622 (N_2622,N_2552,N_2530);
nor U2623 (N_2623,N_2573,N_2537);
or U2624 (N_2624,N_2501,N_2555);
nor U2625 (N_2625,N_2575,N_2512);
or U2626 (N_2626,N_2529,N_2521);
nand U2627 (N_2627,N_2532,N_2566);
or U2628 (N_2628,N_2515,N_2570);
nor U2629 (N_2629,N_2518,N_2513);
xnor U2630 (N_2630,N_2572,N_2596);
or U2631 (N_2631,N_2507,N_2533);
or U2632 (N_2632,N_2581,N_2509);
nand U2633 (N_2633,N_2594,N_2578);
or U2634 (N_2634,N_2565,N_2554);
and U2635 (N_2635,N_2517,N_2587);
or U2636 (N_2636,N_2586,N_2506);
and U2637 (N_2637,N_2502,N_2510);
or U2638 (N_2638,N_2576,N_2551);
or U2639 (N_2639,N_2539,N_2592);
and U2640 (N_2640,N_2563,N_2580);
and U2641 (N_2641,N_2534,N_2543);
nand U2642 (N_2642,N_2523,N_2550);
nor U2643 (N_2643,N_2511,N_2593);
or U2644 (N_2644,N_2519,N_2556);
nand U2645 (N_2645,N_2584,N_2503);
nand U2646 (N_2646,N_2598,N_2536);
or U2647 (N_2647,N_2574,N_2546);
and U2648 (N_2648,N_2582,N_2583);
and U2649 (N_2649,N_2508,N_2548);
nand U2650 (N_2650,N_2557,N_2592);
and U2651 (N_2651,N_2552,N_2562);
or U2652 (N_2652,N_2570,N_2530);
and U2653 (N_2653,N_2579,N_2539);
nand U2654 (N_2654,N_2536,N_2550);
or U2655 (N_2655,N_2513,N_2540);
and U2656 (N_2656,N_2530,N_2592);
nor U2657 (N_2657,N_2581,N_2540);
nand U2658 (N_2658,N_2513,N_2585);
or U2659 (N_2659,N_2527,N_2509);
or U2660 (N_2660,N_2522,N_2582);
nor U2661 (N_2661,N_2557,N_2569);
or U2662 (N_2662,N_2500,N_2507);
and U2663 (N_2663,N_2543,N_2505);
nor U2664 (N_2664,N_2575,N_2566);
nor U2665 (N_2665,N_2585,N_2552);
nand U2666 (N_2666,N_2577,N_2524);
and U2667 (N_2667,N_2544,N_2504);
nor U2668 (N_2668,N_2568,N_2586);
or U2669 (N_2669,N_2565,N_2564);
nand U2670 (N_2670,N_2532,N_2595);
nor U2671 (N_2671,N_2549,N_2568);
nand U2672 (N_2672,N_2513,N_2575);
and U2673 (N_2673,N_2583,N_2510);
and U2674 (N_2674,N_2512,N_2578);
nand U2675 (N_2675,N_2592,N_2553);
nor U2676 (N_2676,N_2501,N_2512);
nor U2677 (N_2677,N_2508,N_2584);
and U2678 (N_2678,N_2588,N_2501);
and U2679 (N_2679,N_2538,N_2531);
nor U2680 (N_2680,N_2573,N_2539);
nor U2681 (N_2681,N_2516,N_2512);
and U2682 (N_2682,N_2520,N_2548);
nand U2683 (N_2683,N_2531,N_2511);
and U2684 (N_2684,N_2595,N_2510);
and U2685 (N_2685,N_2588,N_2578);
and U2686 (N_2686,N_2586,N_2523);
or U2687 (N_2687,N_2534,N_2597);
nand U2688 (N_2688,N_2509,N_2598);
nor U2689 (N_2689,N_2520,N_2509);
or U2690 (N_2690,N_2511,N_2509);
nand U2691 (N_2691,N_2590,N_2536);
nor U2692 (N_2692,N_2540,N_2516);
nor U2693 (N_2693,N_2535,N_2583);
nor U2694 (N_2694,N_2535,N_2555);
nand U2695 (N_2695,N_2560,N_2552);
and U2696 (N_2696,N_2566,N_2523);
nand U2697 (N_2697,N_2551,N_2565);
and U2698 (N_2698,N_2555,N_2557);
and U2699 (N_2699,N_2519,N_2555);
nor U2700 (N_2700,N_2673,N_2633);
nor U2701 (N_2701,N_2662,N_2696);
and U2702 (N_2702,N_2691,N_2601);
nand U2703 (N_2703,N_2652,N_2609);
and U2704 (N_2704,N_2643,N_2617);
nor U2705 (N_2705,N_2659,N_2669);
nand U2706 (N_2706,N_2663,N_2654);
nor U2707 (N_2707,N_2641,N_2648);
nor U2708 (N_2708,N_2699,N_2618);
nor U2709 (N_2709,N_2676,N_2620);
or U2710 (N_2710,N_2610,N_2622);
or U2711 (N_2711,N_2637,N_2685);
nor U2712 (N_2712,N_2636,N_2645);
nand U2713 (N_2713,N_2665,N_2640);
nor U2714 (N_2714,N_2613,N_2615);
or U2715 (N_2715,N_2688,N_2630);
and U2716 (N_2716,N_2625,N_2693);
nand U2717 (N_2717,N_2672,N_2683);
nor U2718 (N_2718,N_2612,N_2655);
nor U2719 (N_2719,N_2670,N_2689);
or U2720 (N_2720,N_2661,N_2681);
nor U2721 (N_2721,N_2639,N_2664);
nand U2722 (N_2722,N_2646,N_2651);
or U2723 (N_2723,N_2627,N_2623);
and U2724 (N_2724,N_2629,N_2628);
nor U2725 (N_2725,N_2671,N_2649);
nor U2726 (N_2726,N_2631,N_2607);
or U2727 (N_2727,N_2658,N_2667);
nand U2728 (N_2728,N_2695,N_2621);
nand U2729 (N_2729,N_2614,N_2638);
or U2730 (N_2730,N_2602,N_2647);
nand U2731 (N_2731,N_2666,N_2656);
or U2732 (N_2732,N_2660,N_2626);
nand U2733 (N_2733,N_2686,N_2611);
nor U2734 (N_2734,N_2674,N_2679);
and U2735 (N_2735,N_2608,N_2635);
and U2736 (N_2736,N_2657,N_2604);
or U2737 (N_2737,N_2687,N_2678);
or U2738 (N_2738,N_2644,N_2697);
nand U2739 (N_2739,N_2653,N_2650);
or U2740 (N_2740,N_2642,N_2690);
and U2741 (N_2741,N_2677,N_2634);
or U2742 (N_2742,N_2624,N_2680);
and U2743 (N_2743,N_2600,N_2682);
nand U2744 (N_2744,N_2692,N_2698);
nand U2745 (N_2745,N_2684,N_2606);
nor U2746 (N_2746,N_2619,N_2675);
nand U2747 (N_2747,N_2603,N_2616);
or U2748 (N_2748,N_2632,N_2694);
or U2749 (N_2749,N_2605,N_2668);
and U2750 (N_2750,N_2659,N_2630);
nand U2751 (N_2751,N_2621,N_2673);
nand U2752 (N_2752,N_2615,N_2693);
nand U2753 (N_2753,N_2604,N_2600);
nor U2754 (N_2754,N_2631,N_2672);
and U2755 (N_2755,N_2626,N_2688);
nor U2756 (N_2756,N_2691,N_2662);
and U2757 (N_2757,N_2639,N_2653);
or U2758 (N_2758,N_2654,N_2653);
nor U2759 (N_2759,N_2662,N_2656);
nand U2760 (N_2760,N_2661,N_2653);
nand U2761 (N_2761,N_2672,N_2695);
or U2762 (N_2762,N_2666,N_2623);
or U2763 (N_2763,N_2633,N_2676);
nand U2764 (N_2764,N_2619,N_2667);
nor U2765 (N_2765,N_2654,N_2615);
nand U2766 (N_2766,N_2643,N_2622);
and U2767 (N_2767,N_2684,N_2682);
or U2768 (N_2768,N_2631,N_2627);
nor U2769 (N_2769,N_2662,N_2694);
nand U2770 (N_2770,N_2699,N_2667);
or U2771 (N_2771,N_2665,N_2621);
and U2772 (N_2772,N_2621,N_2683);
or U2773 (N_2773,N_2683,N_2664);
or U2774 (N_2774,N_2636,N_2607);
or U2775 (N_2775,N_2659,N_2671);
nand U2776 (N_2776,N_2619,N_2620);
nand U2777 (N_2777,N_2647,N_2652);
and U2778 (N_2778,N_2651,N_2645);
and U2779 (N_2779,N_2681,N_2673);
and U2780 (N_2780,N_2671,N_2654);
and U2781 (N_2781,N_2676,N_2648);
nor U2782 (N_2782,N_2690,N_2636);
nor U2783 (N_2783,N_2642,N_2640);
and U2784 (N_2784,N_2660,N_2667);
nor U2785 (N_2785,N_2647,N_2609);
nor U2786 (N_2786,N_2685,N_2620);
and U2787 (N_2787,N_2623,N_2604);
or U2788 (N_2788,N_2651,N_2678);
or U2789 (N_2789,N_2621,N_2622);
nor U2790 (N_2790,N_2672,N_2678);
or U2791 (N_2791,N_2637,N_2611);
and U2792 (N_2792,N_2616,N_2602);
nor U2793 (N_2793,N_2649,N_2672);
and U2794 (N_2794,N_2647,N_2674);
or U2795 (N_2795,N_2656,N_2693);
or U2796 (N_2796,N_2698,N_2691);
and U2797 (N_2797,N_2607,N_2680);
and U2798 (N_2798,N_2674,N_2684);
or U2799 (N_2799,N_2681,N_2685);
or U2800 (N_2800,N_2785,N_2724);
nand U2801 (N_2801,N_2784,N_2778);
nor U2802 (N_2802,N_2715,N_2753);
nand U2803 (N_2803,N_2775,N_2717);
or U2804 (N_2804,N_2712,N_2777);
or U2805 (N_2805,N_2770,N_2706);
and U2806 (N_2806,N_2704,N_2702);
nand U2807 (N_2807,N_2740,N_2786);
and U2808 (N_2808,N_2767,N_2795);
nor U2809 (N_2809,N_2743,N_2781);
nor U2810 (N_2810,N_2727,N_2719);
nand U2811 (N_2811,N_2783,N_2738);
nor U2812 (N_2812,N_2730,N_2747);
nor U2813 (N_2813,N_2737,N_2762);
nand U2814 (N_2814,N_2739,N_2725);
or U2815 (N_2815,N_2797,N_2799);
and U2816 (N_2816,N_2703,N_2755);
or U2817 (N_2817,N_2701,N_2736);
nor U2818 (N_2818,N_2741,N_2776);
or U2819 (N_2819,N_2731,N_2732);
nor U2820 (N_2820,N_2752,N_2750);
or U2821 (N_2821,N_2794,N_2721);
nand U2822 (N_2822,N_2726,N_2707);
nand U2823 (N_2823,N_2742,N_2733);
nand U2824 (N_2824,N_2735,N_2760);
or U2825 (N_2825,N_2711,N_2718);
or U2826 (N_2826,N_2798,N_2757);
and U2827 (N_2827,N_2708,N_2723);
or U2828 (N_2828,N_2714,N_2769);
nand U2829 (N_2829,N_2746,N_2754);
nand U2830 (N_2830,N_2796,N_2745);
and U2831 (N_2831,N_2788,N_2748);
or U2832 (N_2832,N_2779,N_2751);
nor U2833 (N_2833,N_2792,N_2728);
or U2834 (N_2834,N_2780,N_2766);
and U2835 (N_2835,N_2709,N_2710);
or U2836 (N_2836,N_2763,N_2722);
and U2837 (N_2837,N_2756,N_2758);
nand U2838 (N_2838,N_2782,N_2765);
and U2839 (N_2839,N_2761,N_2749);
nand U2840 (N_2840,N_2700,N_2759);
nor U2841 (N_2841,N_2744,N_2713);
or U2842 (N_2842,N_2771,N_2790);
nand U2843 (N_2843,N_2764,N_2791);
nor U2844 (N_2844,N_2705,N_2729);
or U2845 (N_2845,N_2773,N_2774);
and U2846 (N_2846,N_2716,N_2787);
nor U2847 (N_2847,N_2720,N_2768);
nor U2848 (N_2848,N_2734,N_2772);
nor U2849 (N_2849,N_2793,N_2789);
and U2850 (N_2850,N_2780,N_2763);
nor U2851 (N_2851,N_2786,N_2755);
nor U2852 (N_2852,N_2712,N_2783);
and U2853 (N_2853,N_2754,N_2727);
nor U2854 (N_2854,N_2709,N_2740);
and U2855 (N_2855,N_2794,N_2781);
nand U2856 (N_2856,N_2770,N_2781);
or U2857 (N_2857,N_2749,N_2783);
nand U2858 (N_2858,N_2743,N_2724);
nor U2859 (N_2859,N_2781,N_2728);
nand U2860 (N_2860,N_2761,N_2792);
nand U2861 (N_2861,N_2717,N_2772);
xor U2862 (N_2862,N_2774,N_2786);
and U2863 (N_2863,N_2741,N_2755);
nand U2864 (N_2864,N_2748,N_2761);
nor U2865 (N_2865,N_2731,N_2724);
nor U2866 (N_2866,N_2723,N_2715);
nor U2867 (N_2867,N_2753,N_2702);
or U2868 (N_2868,N_2750,N_2727);
nor U2869 (N_2869,N_2792,N_2741);
nor U2870 (N_2870,N_2744,N_2785);
or U2871 (N_2871,N_2775,N_2744);
and U2872 (N_2872,N_2779,N_2730);
nor U2873 (N_2873,N_2754,N_2700);
or U2874 (N_2874,N_2734,N_2735);
and U2875 (N_2875,N_2710,N_2743);
nand U2876 (N_2876,N_2728,N_2747);
and U2877 (N_2877,N_2720,N_2725);
nor U2878 (N_2878,N_2728,N_2754);
and U2879 (N_2879,N_2768,N_2725);
nand U2880 (N_2880,N_2742,N_2780);
nor U2881 (N_2881,N_2790,N_2741);
nand U2882 (N_2882,N_2799,N_2705);
or U2883 (N_2883,N_2777,N_2738);
nand U2884 (N_2884,N_2779,N_2775);
and U2885 (N_2885,N_2700,N_2736);
nand U2886 (N_2886,N_2747,N_2726);
nor U2887 (N_2887,N_2752,N_2766);
nor U2888 (N_2888,N_2754,N_2759);
and U2889 (N_2889,N_2771,N_2760);
nor U2890 (N_2890,N_2783,N_2728);
nor U2891 (N_2891,N_2767,N_2734);
nand U2892 (N_2892,N_2791,N_2785);
nor U2893 (N_2893,N_2735,N_2717);
nand U2894 (N_2894,N_2785,N_2755);
nand U2895 (N_2895,N_2706,N_2766);
nand U2896 (N_2896,N_2776,N_2705);
nor U2897 (N_2897,N_2733,N_2723);
nand U2898 (N_2898,N_2706,N_2798);
and U2899 (N_2899,N_2749,N_2701);
or U2900 (N_2900,N_2865,N_2859);
or U2901 (N_2901,N_2847,N_2809);
or U2902 (N_2902,N_2843,N_2826);
or U2903 (N_2903,N_2889,N_2842);
nand U2904 (N_2904,N_2858,N_2891);
nand U2905 (N_2905,N_2844,N_2830);
or U2906 (N_2906,N_2881,N_2806);
and U2907 (N_2907,N_2839,N_2890);
nor U2908 (N_2908,N_2835,N_2895);
and U2909 (N_2909,N_2805,N_2833);
or U2910 (N_2910,N_2845,N_2894);
nor U2911 (N_2911,N_2896,N_2818);
nor U2912 (N_2912,N_2803,N_2866);
and U2913 (N_2913,N_2888,N_2823);
nand U2914 (N_2914,N_2837,N_2814);
and U2915 (N_2915,N_2852,N_2838);
or U2916 (N_2916,N_2868,N_2807);
and U2917 (N_2917,N_2878,N_2829);
or U2918 (N_2918,N_2808,N_2886);
and U2919 (N_2919,N_2819,N_2812);
and U2920 (N_2920,N_2867,N_2892);
nor U2921 (N_2921,N_2853,N_2804);
or U2922 (N_2922,N_2813,N_2815);
nand U2923 (N_2923,N_2848,N_2817);
nor U2924 (N_2924,N_2834,N_2884);
and U2925 (N_2925,N_2810,N_2821);
and U2926 (N_2926,N_2824,N_2864);
and U2927 (N_2927,N_2828,N_2877);
nor U2928 (N_2928,N_2822,N_2872);
or U2929 (N_2929,N_2863,N_2855);
nor U2930 (N_2930,N_2825,N_2841);
nand U2931 (N_2931,N_2876,N_2871);
nor U2932 (N_2932,N_2801,N_2870);
nand U2933 (N_2933,N_2869,N_2882);
nand U2934 (N_2934,N_2827,N_2893);
and U2935 (N_2935,N_2800,N_2851);
nand U2936 (N_2936,N_2880,N_2873);
or U2937 (N_2937,N_2856,N_2850);
nor U2938 (N_2938,N_2899,N_2846);
or U2939 (N_2939,N_2861,N_2849);
nor U2940 (N_2940,N_2862,N_2887);
nand U2941 (N_2941,N_2874,N_2816);
nor U2942 (N_2942,N_2883,N_2857);
nand U2943 (N_2943,N_2836,N_2811);
or U2944 (N_2944,N_2875,N_2832);
nor U2945 (N_2945,N_2879,N_2897);
nor U2946 (N_2946,N_2831,N_2854);
nor U2947 (N_2947,N_2885,N_2860);
or U2948 (N_2948,N_2840,N_2820);
nand U2949 (N_2949,N_2802,N_2898);
and U2950 (N_2950,N_2851,N_2881);
nand U2951 (N_2951,N_2887,N_2884);
nand U2952 (N_2952,N_2848,N_2834);
and U2953 (N_2953,N_2892,N_2850);
nand U2954 (N_2954,N_2840,N_2893);
or U2955 (N_2955,N_2863,N_2815);
and U2956 (N_2956,N_2804,N_2864);
nand U2957 (N_2957,N_2827,N_2843);
nor U2958 (N_2958,N_2827,N_2811);
nor U2959 (N_2959,N_2874,N_2835);
or U2960 (N_2960,N_2858,N_2803);
or U2961 (N_2961,N_2868,N_2800);
and U2962 (N_2962,N_2845,N_2827);
nand U2963 (N_2963,N_2810,N_2885);
or U2964 (N_2964,N_2814,N_2888);
nand U2965 (N_2965,N_2823,N_2849);
or U2966 (N_2966,N_2881,N_2877);
and U2967 (N_2967,N_2856,N_2849);
nand U2968 (N_2968,N_2893,N_2881);
and U2969 (N_2969,N_2832,N_2884);
nand U2970 (N_2970,N_2818,N_2893);
and U2971 (N_2971,N_2849,N_2818);
nor U2972 (N_2972,N_2888,N_2838);
or U2973 (N_2973,N_2848,N_2872);
nor U2974 (N_2974,N_2838,N_2802);
nor U2975 (N_2975,N_2869,N_2864);
or U2976 (N_2976,N_2884,N_2816);
nor U2977 (N_2977,N_2817,N_2841);
nor U2978 (N_2978,N_2839,N_2884);
nor U2979 (N_2979,N_2837,N_2874);
or U2980 (N_2980,N_2807,N_2865);
and U2981 (N_2981,N_2842,N_2869);
or U2982 (N_2982,N_2841,N_2882);
nor U2983 (N_2983,N_2833,N_2836);
and U2984 (N_2984,N_2877,N_2872);
and U2985 (N_2985,N_2802,N_2865);
nand U2986 (N_2986,N_2837,N_2884);
nor U2987 (N_2987,N_2854,N_2840);
nor U2988 (N_2988,N_2838,N_2847);
or U2989 (N_2989,N_2830,N_2877);
or U2990 (N_2990,N_2811,N_2847);
and U2991 (N_2991,N_2875,N_2819);
nand U2992 (N_2992,N_2821,N_2860);
or U2993 (N_2993,N_2838,N_2880);
nor U2994 (N_2994,N_2857,N_2894);
or U2995 (N_2995,N_2898,N_2862);
nor U2996 (N_2996,N_2849,N_2883);
nor U2997 (N_2997,N_2858,N_2814);
nand U2998 (N_2998,N_2854,N_2860);
nand U2999 (N_2999,N_2817,N_2893);
nand U3000 (N_3000,N_2946,N_2982);
nor U3001 (N_3001,N_2983,N_2994);
nand U3002 (N_3002,N_2930,N_2923);
nand U3003 (N_3003,N_2965,N_2928);
xnor U3004 (N_3004,N_2948,N_2926);
or U3005 (N_3005,N_2997,N_2999);
xor U3006 (N_3006,N_2958,N_2966);
nor U3007 (N_3007,N_2914,N_2955);
or U3008 (N_3008,N_2905,N_2990);
nand U3009 (N_3009,N_2913,N_2929);
and U3010 (N_3010,N_2974,N_2962);
nor U3011 (N_3011,N_2900,N_2978);
nor U3012 (N_3012,N_2992,N_2985);
and U3013 (N_3013,N_2935,N_2980);
nor U3014 (N_3014,N_2931,N_2957);
or U3015 (N_3015,N_2961,N_2991);
nand U3016 (N_3016,N_2995,N_2959);
nand U3017 (N_3017,N_2939,N_2981);
or U3018 (N_3018,N_2952,N_2996);
and U3019 (N_3019,N_2979,N_2944);
or U3020 (N_3020,N_2902,N_2989);
and U3021 (N_3021,N_2916,N_2922);
nand U3022 (N_3022,N_2921,N_2951);
or U3023 (N_3023,N_2911,N_2940);
and U3024 (N_3024,N_2917,N_2986);
nor U3025 (N_3025,N_2925,N_2901);
nor U3026 (N_3026,N_2950,N_2936);
nand U3027 (N_3027,N_2919,N_2938);
nand U3028 (N_3028,N_2903,N_2988);
and U3029 (N_3029,N_2956,N_2967);
nor U3030 (N_3030,N_2918,N_2932);
nand U3031 (N_3031,N_2972,N_2907);
nand U3032 (N_3032,N_2910,N_2976);
nand U3033 (N_3033,N_2953,N_2984);
nor U3034 (N_3034,N_2947,N_2924);
or U3035 (N_3035,N_2941,N_2934);
nand U3036 (N_3036,N_2964,N_2970);
nand U3037 (N_3037,N_2993,N_2977);
nand U3038 (N_3038,N_2942,N_2975);
nand U3039 (N_3039,N_2904,N_2943);
and U3040 (N_3040,N_2933,N_2960);
nand U3041 (N_3041,N_2949,N_2968);
nand U3042 (N_3042,N_2971,N_2987);
nand U3043 (N_3043,N_2915,N_2945);
or U3044 (N_3044,N_2920,N_2954);
nor U3045 (N_3045,N_2998,N_2906);
or U3046 (N_3046,N_2912,N_2969);
or U3047 (N_3047,N_2909,N_2937);
and U3048 (N_3048,N_2927,N_2963);
nor U3049 (N_3049,N_2973,N_2908);
or U3050 (N_3050,N_2910,N_2965);
nor U3051 (N_3051,N_2928,N_2924);
and U3052 (N_3052,N_2981,N_2912);
nand U3053 (N_3053,N_2947,N_2987);
and U3054 (N_3054,N_2900,N_2984);
nor U3055 (N_3055,N_2902,N_2980);
nand U3056 (N_3056,N_2991,N_2917);
and U3057 (N_3057,N_2969,N_2924);
nand U3058 (N_3058,N_2963,N_2907);
or U3059 (N_3059,N_2944,N_2933);
nor U3060 (N_3060,N_2996,N_2977);
nand U3061 (N_3061,N_2919,N_2914);
and U3062 (N_3062,N_2947,N_2932);
or U3063 (N_3063,N_2973,N_2957);
nor U3064 (N_3064,N_2953,N_2910);
nand U3065 (N_3065,N_2933,N_2936);
nand U3066 (N_3066,N_2915,N_2992);
nand U3067 (N_3067,N_2945,N_2981);
nor U3068 (N_3068,N_2911,N_2974);
nand U3069 (N_3069,N_2954,N_2925);
nand U3070 (N_3070,N_2928,N_2988);
nor U3071 (N_3071,N_2940,N_2991);
or U3072 (N_3072,N_2991,N_2972);
nor U3073 (N_3073,N_2972,N_2943);
nand U3074 (N_3074,N_2966,N_2921);
nand U3075 (N_3075,N_2953,N_2905);
nor U3076 (N_3076,N_2962,N_2956);
and U3077 (N_3077,N_2954,N_2953);
and U3078 (N_3078,N_2907,N_2980);
nor U3079 (N_3079,N_2938,N_2980);
or U3080 (N_3080,N_2903,N_2967);
and U3081 (N_3081,N_2992,N_2925);
nand U3082 (N_3082,N_2916,N_2990);
or U3083 (N_3083,N_2988,N_2934);
and U3084 (N_3084,N_2940,N_2957);
or U3085 (N_3085,N_2993,N_2999);
or U3086 (N_3086,N_2929,N_2983);
or U3087 (N_3087,N_2917,N_2938);
nand U3088 (N_3088,N_2944,N_2943);
nand U3089 (N_3089,N_2937,N_2977);
or U3090 (N_3090,N_2977,N_2905);
or U3091 (N_3091,N_2983,N_2911);
nor U3092 (N_3092,N_2918,N_2941);
nor U3093 (N_3093,N_2926,N_2902);
and U3094 (N_3094,N_2903,N_2949);
nor U3095 (N_3095,N_2902,N_2962);
and U3096 (N_3096,N_2900,N_2939);
and U3097 (N_3097,N_2905,N_2902);
or U3098 (N_3098,N_2961,N_2939);
nor U3099 (N_3099,N_2936,N_2984);
nand U3100 (N_3100,N_3081,N_3031);
nand U3101 (N_3101,N_3041,N_3093);
and U3102 (N_3102,N_3011,N_3032);
and U3103 (N_3103,N_3068,N_3072);
nand U3104 (N_3104,N_3026,N_3019);
nor U3105 (N_3105,N_3087,N_3062);
and U3106 (N_3106,N_3048,N_3013);
and U3107 (N_3107,N_3022,N_3029);
nand U3108 (N_3108,N_3015,N_3001);
nand U3109 (N_3109,N_3063,N_3005);
nor U3110 (N_3110,N_3092,N_3037);
nand U3111 (N_3111,N_3060,N_3052);
and U3112 (N_3112,N_3058,N_3077);
nor U3113 (N_3113,N_3085,N_3044);
nand U3114 (N_3114,N_3054,N_3059);
nand U3115 (N_3115,N_3099,N_3027);
or U3116 (N_3116,N_3073,N_3034);
or U3117 (N_3117,N_3089,N_3050);
nand U3118 (N_3118,N_3074,N_3096);
nor U3119 (N_3119,N_3075,N_3083);
nor U3120 (N_3120,N_3000,N_3040);
or U3121 (N_3121,N_3051,N_3009);
or U3122 (N_3122,N_3008,N_3091);
nor U3123 (N_3123,N_3082,N_3086);
or U3124 (N_3124,N_3038,N_3080);
or U3125 (N_3125,N_3036,N_3056);
nand U3126 (N_3126,N_3084,N_3018);
and U3127 (N_3127,N_3098,N_3014);
nor U3128 (N_3128,N_3066,N_3053);
and U3129 (N_3129,N_3003,N_3006);
nor U3130 (N_3130,N_3007,N_3065);
and U3131 (N_3131,N_3021,N_3049);
or U3132 (N_3132,N_3078,N_3070);
or U3133 (N_3133,N_3002,N_3088);
nand U3134 (N_3134,N_3076,N_3020);
or U3135 (N_3135,N_3017,N_3024);
or U3136 (N_3136,N_3064,N_3039);
and U3137 (N_3137,N_3094,N_3035);
nor U3138 (N_3138,N_3016,N_3079);
nand U3139 (N_3139,N_3042,N_3043);
nand U3140 (N_3140,N_3045,N_3046);
nand U3141 (N_3141,N_3023,N_3055);
nor U3142 (N_3142,N_3033,N_3010);
and U3143 (N_3143,N_3069,N_3090);
and U3144 (N_3144,N_3047,N_3097);
nor U3145 (N_3145,N_3067,N_3028);
nor U3146 (N_3146,N_3061,N_3004);
or U3147 (N_3147,N_3025,N_3071);
and U3148 (N_3148,N_3057,N_3030);
and U3149 (N_3149,N_3095,N_3012);
and U3150 (N_3150,N_3057,N_3027);
nor U3151 (N_3151,N_3096,N_3088);
nor U3152 (N_3152,N_3093,N_3045);
or U3153 (N_3153,N_3014,N_3060);
nor U3154 (N_3154,N_3024,N_3097);
and U3155 (N_3155,N_3029,N_3076);
or U3156 (N_3156,N_3029,N_3048);
and U3157 (N_3157,N_3057,N_3069);
and U3158 (N_3158,N_3002,N_3075);
or U3159 (N_3159,N_3033,N_3055);
or U3160 (N_3160,N_3086,N_3003);
and U3161 (N_3161,N_3048,N_3049);
nand U3162 (N_3162,N_3019,N_3079);
or U3163 (N_3163,N_3069,N_3048);
nand U3164 (N_3164,N_3016,N_3073);
nor U3165 (N_3165,N_3040,N_3045);
and U3166 (N_3166,N_3013,N_3087);
nor U3167 (N_3167,N_3040,N_3019);
nor U3168 (N_3168,N_3063,N_3020);
or U3169 (N_3169,N_3007,N_3017);
nand U3170 (N_3170,N_3079,N_3063);
nor U3171 (N_3171,N_3086,N_3029);
nor U3172 (N_3172,N_3034,N_3089);
nand U3173 (N_3173,N_3004,N_3019);
and U3174 (N_3174,N_3081,N_3054);
or U3175 (N_3175,N_3024,N_3057);
nand U3176 (N_3176,N_3013,N_3071);
or U3177 (N_3177,N_3085,N_3031);
or U3178 (N_3178,N_3037,N_3058);
nand U3179 (N_3179,N_3035,N_3091);
and U3180 (N_3180,N_3094,N_3073);
and U3181 (N_3181,N_3097,N_3006);
and U3182 (N_3182,N_3040,N_3090);
xor U3183 (N_3183,N_3029,N_3089);
nand U3184 (N_3184,N_3041,N_3005);
nand U3185 (N_3185,N_3049,N_3011);
and U3186 (N_3186,N_3075,N_3088);
nand U3187 (N_3187,N_3073,N_3054);
nand U3188 (N_3188,N_3019,N_3091);
or U3189 (N_3189,N_3089,N_3071);
nand U3190 (N_3190,N_3074,N_3011);
nor U3191 (N_3191,N_3075,N_3099);
and U3192 (N_3192,N_3058,N_3026);
nand U3193 (N_3193,N_3004,N_3052);
or U3194 (N_3194,N_3084,N_3027);
or U3195 (N_3195,N_3066,N_3065);
and U3196 (N_3196,N_3043,N_3005);
xnor U3197 (N_3197,N_3032,N_3090);
or U3198 (N_3198,N_3099,N_3070);
nand U3199 (N_3199,N_3041,N_3029);
nor U3200 (N_3200,N_3155,N_3147);
nor U3201 (N_3201,N_3128,N_3110);
or U3202 (N_3202,N_3143,N_3125);
nor U3203 (N_3203,N_3184,N_3108);
and U3204 (N_3204,N_3153,N_3131);
or U3205 (N_3205,N_3197,N_3148);
nand U3206 (N_3206,N_3168,N_3192);
or U3207 (N_3207,N_3100,N_3119);
xnor U3208 (N_3208,N_3144,N_3134);
nor U3209 (N_3209,N_3123,N_3109);
nor U3210 (N_3210,N_3111,N_3198);
and U3211 (N_3211,N_3179,N_3118);
or U3212 (N_3212,N_3142,N_3178);
and U3213 (N_3213,N_3103,N_3190);
or U3214 (N_3214,N_3139,N_3107);
and U3215 (N_3215,N_3149,N_3194);
nor U3216 (N_3216,N_3124,N_3158);
and U3217 (N_3217,N_3195,N_3120);
or U3218 (N_3218,N_3191,N_3122);
nor U3219 (N_3219,N_3173,N_3170);
and U3220 (N_3220,N_3127,N_3150);
and U3221 (N_3221,N_3183,N_3193);
nand U3222 (N_3222,N_3164,N_3105);
nor U3223 (N_3223,N_3176,N_3136);
or U3224 (N_3224,N_3199,N_3181);
and U3225 (N_3225,N_3115,N_3146);
and U3226 (N_3226,N_3104,N_3174);
nand U3227 (N_3227,N_3160,N_3186);
or U3228 (N_3228,N_3152,N_3172);
nor U3229 (N_3229,N_3135,N_3171);
nand U3230 (N_3230,N_3163,N_3133);
nand U3231 (N_3231,N_3156,N_3113);
nor U3232 (N_3232,N_3185,N_3101);
nand U3233 (N_3233,N_3151,N_3138);
nand U3234 (N_3234,N_3169,N_3188);
nor U3235 (N_3235,N_3157,N_3166);
nand U3236 (N_3236,N_3159,N_3196);
and U3237 (N_3237,N_3126,N_3106);
nand U3238 (N_3238,N_3154,N_3140);
or U3239 (N_3239,N_3116,N_3141);
or U3240 (N_3240,N_3132,N_3137);
or U3241 (N_3241,N_3165,N_3130);
nand U3242 (N_3242,N_3162,N_3102);
nor U3243 (N_3243,N_3121,N_3112);
nand U3244 (N_3244,N_3182,N_3175);
and U3245 (N_3245,N_3187,N_3177);
or U3246 (N_3246,N_3189,N_3114);
or U3247 (N_3247,N_3180,N_3167);
nand U3248 (N_3248,N_3161,N_3117);
or U3249 (N_3249,N_3145,N_3129);
nor U3250 (N_3250,N_3195,N_3153);
and U3251 (N_3251,N_3133,N_3190);
and U3252 (N_3252,N_3179,N_3137);
and U3253 (N_3253,N_3185,N_3193);
or U3254 (N_3254,N_3147,N_3166);
nand U3255 (N_3255,N_3108,N_3168);
nand U3256 (N_3256,N_3100,N_3150);
nand U3257 (N_3257,N_3174,N_3170);
or U3258 (N_3258,N_3118,N_3124);
nor U3259 (N_3259,N_3170,N_3190);
or U3260 (N_3260,N_3189,N_3182);
and U3261 (N_3261,N_3138,N_3116);
nor U3262 (N_3262,N_3179,N_3117);
xor U3263 (N_3263,N_3139,N_3129);
and U3264 (N_3264,N_3119,N_3194);
or U3265 (N_3265,N_3167,N_3193);
and U3266 (N_3266,N_3192,N_3198);
and U3267 (N_3267,N_3133,N_3141);
nor U3268 (N_3268,N_3196,N_3128);
or U3269 (N_3269,N_3123,N_3193);
nor U3270 (N_3270,N_3109,N_3199);
nor U3271 (N_3271,N_3172,N_3168);
nand U3272 (N_3272,N_3131,N_3172);
and U3273 (N_3273,N_3100,N_3177);
or U3274 (N_3274,N_3128,N_3179);
nor U3275 (N_3275,N_3156,N_3131);
and U3276 (N_3276,N_3153,N_3188);
nand U3277 (N_3277,N_3115,N_3125);
nand U3278 (N_3278,N_3138,N_3180);
nor U3279 (N_3279,N_3170,N_3189);
nor U3280 (N_3280,N_3104,N_3189);
and U3281 (N_3281,N_3101,N_3189);
nand U3282 (N_3282,N_3156,N_3136);
and U3283 (N_3283,N_3117,N_3154);
or U3284 (N_3284,N_3113,N_3110);
or U3285 (N_3285,N_3175,N_3135);
and U3286 (N_3286,N_3172,N_3130);
nor U3287 (N_3287,N_3137,N_3174);
and U3288 (N_3288,N_3126,N_3191);
nand U3289 (N_3289,N_3118,N_3163);
nand U3290 (N_3290,N_3147,N_3102);
nor U3291 (N_3291,N_3110,N_3148);
or U3292 (N_3292,N_3151,N_3103);
nand U3293 (N_3293,N_3116,N_3144);
and U3294 (N_3294,N_3135,N_3149);
nor U3295 (N_3295,N_3173,N_3136);
or U3296 (N_3296,N_3185,N_3171);
or U3297 (N_3297,N_3165,N_3118);
nand U3298 (N_3298,N_3104,N_3127);
nand U3299 (N_3299,N_3150,N_3117);
and U3300 (N_3300,N_3256,N_3277);
nor U3301 (N_3301,N_3204,N_3246);
nor U3302 (N_3302,N_3251,N_3274);
nand U3303 (N_3303,N_3235,N_3258);
nor U3304 (N_3304,N_3212,N_3252);
or U3305 (N_3305,N_3264,N_3210);
and U3306 (N_3306,N_3208,N_3278);
and U3307 (N_3307,N_3205,N_3203);
nor U3308 (N_3308,N_3298,N_3218);
nor U3309 (N_3309,N_3269,N_3202);
and U3310 (N_3310,N_3261,N_3248);
and U3311 (N_3311,N_3223,N_3280);
or U3312 (N_3312,N_3228,N_3247);
or U3313 (N_3313,N_3272,N_3282);
nor U3314 (N_3314,N_3214,N_3236);
or U3315 (N_3315,N_3279,N_3233);
or U3316 (N_3316,N_3283,N_3263);
and U3317 (N_3317,N_3267,N_3265);
or U3318 (N_3318,N_3294,N_3255);
nand U3319 (N_3319,N_3234,N_3297);
nand U3320 (N_3320,N_3201,N_3220);
and U3321 (N_3321,N_3270,N_3206);
and U3322 (N_3322,N_3275,N_3242);
nor U3323 (N_3323,N_3253,N_3215);
or U3324 (N_3324,N_3250,N_3211);
nor U3325 (N_3325,N_3260,N_3229);
or U3326 (N_3326,N_3225,N_3217);
nand U3327 (N_3327,N_3266,N_3259);
xor U3328 (N_3328,N_3240,N_3292);
nor U3329 (N_3329,N_3271,N_3213);
nand U3330 (N_3330,N_3296,N_3243);
and U3331 (N_3331,N_3232,N_3239);
nand U3332 (N_3332,N_3245,N_3221);
nor U3333 (N_3333,N_3281,N_3257);
and U3334 (N_3334,N_3268,N_3226);
or U3335 (N_3335,N_3295,N_3286);
nor U3336 (N_3336,N_3237,N_3230);
or U3337 (N_3337,N_3284,N_3273);
and U3338 (N_3338,N_3238,N_3289);
and U3339 (N_3339,N_3288,N_3293);
and U3340 (N_3340,N_3285,N_3254);
or U3341 (N_3341,N_3249,N_3227);
nor U3342 (N_3342,N_3200,N_3290);
and U3343 (N_3343,N_3287,N_3276);
nor U3344 (N_3344,N_3222,N_3216);
and U3345 (N_3345,N_3241,N_3207);
and U3346 (N_3346,N_3209,N_3244);
or U3347 (N_3347,N_3262,N_3231);
nor U3348 (N_3348,N_3219,N_3224);
nor U3349 (N_3349,N_3291,N_3299);
or U3350 (N_3350,N_3237,N_3249);
and U3351 (N_3351,N_3208,N_3274);
or U3352 (N_3352,N_3243,N_3211);
nor U3353 (N_3353,N_3218,N_3212);
nor U3354 (N_3354,N_3241,N_3201);
and U3355 (N_3355,N_3234,N_3268);
and U3356 (N_3356,N_3231,N_3257);
nand U3357 (N_3357,N_3276,N_3257);
and U3358 (N_3358,N_3244,N_3297);
xnor U3359 (N_3359,N_3227,N_3293);
nor U3360 (N_3360,N_3285,N_3206);
nor U3361 (N_3361,N_3262,N_3294);
and U3362 (N_3362,N_3202,N_3236);
or U3363 (N_3363,N_3205,N_3281);
or U3364 (N_3364,N_3267,N_3269);
nand U3365 (N_3365,N_3243,N_3286);
nand U3366 (N_3366,N_3202,N_3283);
nand U3367 (N_3367,N_3225,N_3272);
nor U3368 (N_3368,N_3287,N_3210);
nor U3369 (N_3369,N_3225,N_3263);
nor U3370 (N_3370,N_3219,N_3239);
nor U3371 (N_3371,N_3231,N_3260);
and U3372 (N_3372,N_3298,N_3248);
nor U3373 (N_3373,N_3262,N_3271);
or U3374 (N_3374,N_3252,N_3289);
and U3375 (N_3375,N_3282,N_3225);
nand U3376 (N_3376,N_3264,N_3232);
nand U3377 (N_3377,N_3238,N_3222);
or U3378 (N_3378,N_3291,N_3285);
nor U3379 (N_3379,N_3233,N_3295);
and U3380 (N_3380,N_3257,N_3220);
nand U3381 (N_3381,N_3263,N_3210);
or U3382 (N_3382,N_3291,N_3202);
and U3383 (N_3383,N_3243,N_3245);
nor U3384 (N_3384,N_3292,N_3268);
and U3385 (N_3385,N_3293,N_3263);
nor U3386 (N_3386,N_3285,N_3240);
or U3387 (N_3387,N_3277,N_3282);
nor U3388 (N_3388,N_3228,N_3295);
nor U3389 (N_3389,N_3200,N_3262);
or U3390 (N_3390,N_3207,N_3270);
nand U3391 (N_3391,N_3214,N_3298);
nor U3392 (N_3392,N_3244,N_3255);
or U3393 (N_3393,N_3243,N_3224);
nand U3394 (N_3394,N_3280,N_3254);
or U3395 (N_3395,N_3284,N_3234);
nand U3396 (N_3396,N_3218,N_3205);
nor U3397 (N_3397,N_3284,N_3265);
or U3398 (N_3398,N_3222,N_3299);
or U3399 (N_3399,N_3272,N_3204);
nor U3400 (N_3400,N_3348,N_3375);
and U3401 (N_3401,N_3305,N_3387);
nand U3402 (N_3402,N_3377,N_3302);
or U3403 (N_3403,N_3351,N_3315);
nor U3404 (N_3404,N_3382,N_3341);
or U3405 (N_3405,N_3309,N_3331);
nor U3406 (N_3406,N_3352,N_3364);
nand U3407 (N_3407,N_3399,N_3333);
nor U3408 (N_3408,N_3329,N_3355);
nor U3409 (N_3409,N_3363,N_3304);
nand U3410 (N_3410,N_3332,N_3318);
or U3411 (N_3411,N_3335,N_3350);
and U3412 (N_3412,N_3383,N_3396);
nand U3413 (N_3413,N_3349,N_3371);
nand U3414 (N_3414,N_3374,N_3321);
nand U3415 (N_3415,N_3312,N_3311);
or U3416 (N_3416,N_3313,N_3395);
nand U3417 (N_3417,N_3365,N_3353);
nand U3418 (N_3418,N_3389,N_3356);
or U3419 (N_3419,N_3336,N_3325);
nand U3420 (N_3420,N_3337,N_3393);
or U3421 (N_3421,N_3378,N_3347);
nand U3422 (N_3422,N_3345,N_3324);
nand U3423 (N_3423,N_3301,N_3323);
or U3424 (N_3424,N_3328,N_3361);
and U3425 (N_3425,N_3385,N_3386);
or U3426 (N_3426,N_3392,N_3362);
nand U3427 (N_3427,N_3340,N_3381);
nand U3428 (N_3428,N_3370,N_3376);
nand U3429 (N_3429,N_3391,N_3369);
nand U3430 (N_3430,N_3317,N_3358);
nor U3431 (N_3431,N_3339,N_3368);
or U3432 (N_3432,N_3344,N_3379);
or U3433 (N_3433,N_3366,N_3354);
or U3434 (N_3434,N_3394,N_3346);
or U3435 (N_3435,N_3320,N_3380);
and U3436 (N_3436,N_3319,N_3300);
and U3437 (N_3437,N_3307,N_3327);
nor U3438 (N_3438,N_3306,N_3397);
and U3439 (N_3439,N_3342,N_3384);
nor U3440 (N_3440,N_3373,N_3314);
and U3441 (N_3441,N_3330,N_3308);
and U3442 (N_3442,N_3360,N_3359);
or U3443 (N_3443,N_3343,N_3398);
nor U3444 (N_3444,N_3334,N_3388);
or U3445 (N_3445,N_3390,N_3367);
nor U3446 (N_3446,N_3372,N_3338);
or U3447 (N_3447,N_3322,N_3316);
and U3448 (N_3448,N_3310,N_3357);
and U3449 (N_3449,N_3326,N_3303);
nor U3450 (N_3450,N_3307,N_3325);
and U3451 (N_3451,N_3367,N_3337);
nor U3452 (N_3452,N_3392,N_3365);
or U3453 (N_3453,N_3380,N_3346);
or U3454 (N_3454,N_3324,N_3374);
xor U3455 (N_3455,N_3367,N_3338);
or U3456 (N_3456,N_3327,N_3316);
and U3457 (N_3457,N_3316,N_3330);
nor U3458 (N_3458,N_3303,N_3387);
nor U3459 (N_3459,N_3327,N_3306);
and U3460 (N_3460,N_3387,N_3330);
nor U3461 (N_3461,N_3326,N_3389);
nand U3462 (N_3462,N_3378,N_3364);
nor U3463 (N_3463,N_3349,N_3397);
or U3464 (N_3464,N_3393,N_3318);
and U3465 (N_3465,N_3341,N_3365);
xnor U3466 (N_3466,N_3356,N_3361);
and U3467 (N_3467,N_3362,N_3394);
or U3468 (N_3468,N_3362,N_3390);
nor U3469 (N_3469,N_3348,N_3314);
nand U3470 (N_3470,N_3388,N_3355);
or U3471 (N_3471,N_3354,N_3344);
or U3472 (N_3472,N_3310,N_3398);
or U3473 (N_3473,N_3338,N_3319);
or U3474 (N_3474,N_3380,N_3383);
and U3475 (N_3475,N_3313,N_3376);
and U3476 (N_3476,N_3385,N_3363);
nand U3477 (N_3477,N_3386,N_3398);
nor U3478 (N_3478,N_3350,N_3345);
nand U3479 (N_3479,N_3315,N_3378);
xor U3480 (N_3480,N_3318,N_3329);
and U3481 (N_3481,N_3309,N_3398);
nand U3482 (N_3482,N_3335,N_3399);
nand U3483 (N_3483,N_3334,N_3311);
nor U3484 (N_3484,N_3361,N_3357);
or U3485 (N_3485,N_3339,N_3352);
and U3486 (N_3486,N_3327,N_3380);
nand U3487 (N_3487,N_3396,N_3314);
xor U3488 (N_3488,N_3394,N_3355);
nor U3489 (N_3489,N_3359,N_3369);
nor U3490 (N_3490,N_3302,N_3352);
nand U3491 (N_3491,N_3367,N_3361);
and U3492 (N_3492,N_3370,N_3329);
nand U3493 (N_3493,N_3311,N_3381);
or U3494 (N_3494,N_3339,N_3335);
nor U3495 (N_3495,N_3331,N_3385);
nor U3496 (N_3496,N_3328,N_3355);
nor U3497 (N_3497,N_3342,N_3337);
and U3498 (N_3498,N_3346,N_3313);
nand U3499 (N_3499,N_3314,N_3311);
nand U3500 (N_3500,N_3491,N_3477);
nand U3501 (N_3501,N_3404,N_3459);
and U3502 (N_3502,N_3428,N_3436);
nand U3503 (N_3503,N_3425,N_3418);
or U3504 (N_3504,N_3458,N_3471);
and U3505 (N_3505,N_3416,N_3445);
and U3506 (N_3506,N_3492,N_3464);
and U3507 (N_3507,N_3497,N_3450);
and U3508 (N_3508,N_3410,N_3430);
nor U3509 (N_3509,N_3481,N_3472);
or U3510 (N_3510,N_3442,N_3400);
nand U3511 (N_3511,N_3493,N_3438);
or U3512 (N_3512,N_3454,N_3403);
or U3513 (N_3513,N_3435,N_3417);
xor U3514 (N_3514,N_3432,N_3476);
nand U3515 (N_3515,N_3440,N_3478);
nand U3516 (N_3516,N_3426,N_3489);
and U3517 (N_3517,N_3499,N_3486);
nand U3518 (N_3518,N_3439,N_3437);
nand U3519 (N_3519,N_3451,N_3427);
nor U3520 (N_3520,N_3452,N_3414);
nand U3521 (N_3521,N_3480,N_3470);
nor U3522 (N_3522,N_3468,N_3469);
and U3523 (N_3523,N_3495,N_3429);
or U3524 (N_3524,N_3401,N_3457);
nor U3525 (N_3525,N_3463,N_3409);
and U3526 (N_3526,N_3446,N_3494);
and U3527 (N_3527,N_3433,N_3484);
and U3528 (N_3528,N_3465,N_3473);
nor U3529 (N_3529,N_3462,N_3431);
or U3530 (N_3530,N_3482,N_3461);
and U3531 (N_3531,N_3420,N_3443);
or U3532 (N_3532,N_3474,N_3402);
and U3533 (N_3533,N_3422,N_3467);
nand U3534 (N_3534,N_3415,N_3413);
nor U3535 (N_3535,N_3424,N_3448);
or U3536 (N_3536,N_3460,N_3408);
or U3537 (N_3537,N_3498,N_3485);
or U3538 (N_3538,N_3444,N_3447);
nor U3539 (N_3539,N_3488,N_3479);
nand U3540 (N_3540,N_3449,N_3496);
or U3541 (N_3541,N_3405,N_3407);
and U3542 (N_3542,N_3441,N_3455);
or U3543 (N_3543,N_3406,N_3419);
nand U3544 (N_3544,N_3421,N_3412);
and U3545 (N_3545,N_3483,N_3490);
or U3546 (N_3546,N_3475,N_3456);
nand U3547 (N_3547,N_3487,N_3466);
or U3548 (N_3548,N_3434,N_3423);
nand U3549 (N_3549,N_3411,N_3453);
and U3550 (N_3550,N_3425,N_3401);
or U3551 (N_3551,N_3420,N_3429);
or U3552 (N_3552,N_3424,N_3489);
or U3553 (N_3553,N_3464,N_3475);
nand U3554 (N_3554,N_3486,N_3441);
and U3555 (N_3555,N_3491,N_3456);
and U3556 (N_3556,N_3484,N_3498);
nand U3557 (N_3557,N_3440,N_3416);
and U3558 (N_3558,N_3419,N_3498);
nor U3559 (N_3559,N_3449,N_3431);
nand U3560 (N_3560,N_3444,N_3423);
and U3561 (N_3561,N_3417,N_3402);
or U3562 (N_3562,N_3459,N_3495);
nand U3563 (N_3563,N_3444,N_3412);
and U3564 (N_3564,N_3409,N_3408);
nor U3565 (N_3565,N_3422,N_3414);
and U3566 (N_3566,N_3456,N_3493);
nor U3567 (N_3567,N_3481,N_3446);
nor U3568 (N_3568,N_3470,N_3484);
nor U3569 (N_3569,N_3409,N_3461);
nor U3570 (N_3570,N_3453,N_3483);
nor U3571 (N_3571,N_3486,N_3452);
nand U3572 (N_3572,N_3432,N_3487);
and U3573 (N_3573,N_3402,N_3425);
or U3574 (N_3574,N_3485,N_3460);
nand U3575 (N_3575,N_3416,N_3420);
nand U3576 (N_3576,N_3401,N_3469);
nor U3577 (N_3577,N_3485,N_3402);
nor U3578 (N_3578,N_3448,N_3405);
nand U3579 (N_3579,N_3416,N_3435);
or U3580 (N_3580,N_3410,N_3429);
or U3581 (N_3581,N_3452,N_3413);
or U3582 (N_3582,N_3421,N_3446);
nand U3583 (N_3583,N_3407,N_3454);
nand U3584 (N_3584,N_3412,N_3431);
and U3585 (N_3585,N_3486,N_3480);
and U3586 (N_3586,N_3497,N_3453);
and U3587 (N_3587,N_3402,N_3473);
or U3588 (N_3588,N_3430,N_3428);
or U3589 (N_3589,N_3473,N_3460);
and U3590 (N_3590,N_3488,N_3423);
nand U3591 (N_3591,N_3423,N_3469);
and U3592 (N_3592,N_3472,N_3400);
nand U3593 (N_3593,N_3451,N_3454);
nand U3594 (N_3594,N_3441,N_3468);
or U3595 (N_3595,N_3428,N_3407);
xor U3596 (N_3596,N_3413,N_3403);
or U3597 (N_3597,N_3411,N_3498);
nand U3598 (N_3598,N_3401,N_3498);
and U3599 (N_3599,N_3436,N_3407);
nand U3600 (N_3600,N_3527,N_3541);
nor U3601 (N_3601,N_3564,N_3523);
and U3602 (N_3602,N_3501,N_3553);
nor U3603 (N_3603,N_3515,N_3558);
nor U3604 (N_3604,N_3570,N_3508);
or U3605 (N_3605,N_3519,N_3506);
and U3606 (N_3606,N_3547,N_3557);
nand U3607 (N_3607,N_3571,N_3516);
nand U3608 (N_3608,N_3584,N_3545);
xor U3609 (N_3609,N_3534,N_3577);
nor U3610 (N_3610,N_3537,N_3532);
or U3611 (N_3611,N_3544,N_3569);
nand U3612 (N_3612,N_3580,N_3525);
or U3613 (N_3613,N_3517,N_3511);
and U3614 (N_3614,N_3591,N_3575);
and U3615 (N_3615,N_3589,N_3529);
nand U3616 (N_3616,N_3581,N_3554);
nand U3617 (N_3617,N_3596,N_3518);
and U3618 (N_3618,N_3574,N_3546);
nand U3619 (N_3619,N_3524,N_3543);
nor U3620 (N_3620,N_3526,N_3559);
nand U3621 (N_3621,N_3521,N_3504);
nand U3622 (N_3622,N_3520,N_3552);
and U3623 (N_3623,N_3563,N_3513);
nor U3624 (N_3624,N_3565,N_3592);
and U3625 (N_3625,N_3510,N_3549);
nand U3626 (N_3626,N_3502,N_3560);
nand U3627 (N_3627,N_3530,N_3599);
nor U3628 (N_3628,N_3590,N_3548);
or U3629 (N_3629,N_3503,N_3556);
or U3630 (N_3630,N_3588,N_3568);
and U3631 (N_3631,N_3507,N_3587);
nand U3632 (N_3632,N_3539,N_3540);
and U3633 (N_3633,N_3598,N_3582);
nand U3634 (N_3634,N_3595,N_3594);
nor U3635 (N_3635,N_3538,N_3509);
nor U3636 (N_3636,N_3578,N_3573);
and U3637 (N_3637,N_3555,N_3535);
nand U3638 (N_3638,N_3542,N_3550);
or U3639 (N_3639,N_3567,N_3522);
nor U3640 (N_3640,N_3579,N_3583);
nor U3641 (N_3641,N_3533,N_3566);
nor U3642 (N_3642,N_3514,N_3572);
and U3643 (N_3643,N_3505,N_3536);
or U3644 (N_3644,N_3500,N_3576);
nor U3645 (N_3645,N_3593,N_3562);
and U3646 (N_3646,N_3585,N_3597);
and U3647 (N_3647,N_3512,N_3531);
and U3648 (N_3648,N_3561,N_3551);
nand U3649 (N_3649,N_3586,N_3528);
and U3650 (N_3650,N_3533,N_3541);
and U3651 (N_3651,N_3567,N_3556);
and U3652 (N_3652,N_3538,N_3541);
or U3653 (N_3653,N_3501,N_3530);
and U3654 (N_3654,N_3591,N_3543);
nor U3655 (N_3655,N_3590,N_3520);
nor U3656 (N_3656,N_3516,N_3512);
or U3657 (N_3657,N_3566,N_3549);
nor U3658 (N_3658,N_3556,N_3510);
or U3659 (N_3659,N_3597,N_3537);
or U3660 (N_3660,N_3517,N_3586);
and U3661 (N_3661,N_3541,N_3505);
nor U3662 (N_3662,N_3590,N_3580);
or U3663 (N_3663,N_3592,N_3571);
nand U3664 (N_3664,N_3568,N_3533);
nor U3665 (N_3665,N_3522,N_3570);
and U3666 (N_3666,N_3538,N_3581);
or U3667 (N_3667,N_3590,N_3577);
or U3668 (N_3668,N_3537,N_3577);
and U3669 (N_3669,N_3569,N_3545);
nand U3670 (N_3670,N_3594,N_3515);
nor U3671 (N_3671,N_3595,N_3518);
and U3672 (N_3672,N_3596,N_3507);
or U3673 (N_3673,N_3520,N_3506);
nor U3674 (N_3674,N_3510,N_3584);
and U3675 (N_3675,N_3593,N_3525);
and U3676 (N_3676,N_3587,N_3570);
nor U3677 (N_3677,N_3575,N_3530);
and U3678 (N_3678,N_3534,N_3547);
nand U3679 (N_3679,N_3517,N_3519);
nand U3680 (N_3680,N_3559,N_3540);
nand U3681 (N_3681,N_3591,N_3526);
nand U3682 (N_3682,N_3565,N_3503);
or U3683 (N_3683,N_3524,N_3521);
nand U3684 (N_3684,N_3546,N_3594);
or U3685 (N_3685,N_3563,N_3532);
or U3686 (N_3686,N_3527,N_3555);
or U3687 (N_3687,N_3582,N_3505);
or U3688 (N_3688,N_3547,N_3570);
nor U3689 (N_3689,N_3581,N_3589);
or U3690 (N_3690,N_3586,N_3534);
or U3691 (N_3691,N_3502,N_3588);
and U3692 (N_3692,N_3575,N_3576);
nand U3693 (N_3693,N_3598,N_3544);
or U3694 (N_3694,N_3520,N_3527);
nand U3695 (N_3695,N_3509,N_3573);
or U3696 (N_3696,N_3578,N_3530);
or U3697 (N_3697,N_3530,N_3536);
nor U3698 (N_3698,N_3525,N_3567);
or U3699 (N_3699,N_3502,N_3583);
and U3700 (N_3700,N_3671,N_3604);
nand U3701 (N_3701,N_3676,N_3665);
nor U3702 (N_3702,N_3607,N_3695);
and U3703 (N_3703,N_3615,N_3696);
nand U3704 (N_3704,N_3687,N_3699);
nand U3705 (N_3705,N_3634,N_3682);
or U3706 (N_3706,N_3673,N_3606);
nand U3707 (N_3707,N_3628,N_3670);
nand U3708 (N_3708,N_3638,N_3609);
nand U3709 (N_3709,N_3698,N_3602);
or U3710 (N_3710,N_3605,N_3667);
or U3711 (N_3711,N_3645,N_3689);
and U3712 (N_3712,N_3601,N_3622);
or U3713 (N_3713,N_3653,N_3681);
nand U3714 (N_3714,N_3657,N_3618);
nor U3715 (N_3715,N_3621,N_3686);
nor U3716 (N_3716,N_3678,N_3651);
nand U3717 (N_3717,N_3635,N_3692);
and U3718 (N_3718,N_3614,N_3631);
nor U3719 (N_3719,N_3603,N_3637);
nor U3720 (N_3720,N_3663,N_3672);
nand U3721 (N_3721,N_3639,N_3674);
and U3722 (N_3722,N_3697,N_3694);
nor U3723 (N_3723,N_3640,N_3680);
nand U3724 (N_3724,N_3612,N_3652);
and U3725 (N_3725,N_3688,N_3629);
nor U3726 (N_3726,N_3660,N_3644);
and U3727 (N_3727,N_3611,N_3600);
and U3728 (N_3728,N_3669,N_3642);
nor U3729 (N_3729,N_3630,N_3675);
or U3730 (N_3730,N_3679,N_3647);
and U3731 (N_3731,N_3643,N_3662);
nand U3732 (N_3732,N_3650,N_3668);
nor U3733 (N_3733,N_3626,N_3613);
and U3734 (N_3734,N_3656,N_3661);
or U3735 (N_3735,N_3632,N_3636);
nor U3736 (N_3736,N_3655,N_3693);
nor U3737 (N_3737,N_3685,N_3619);
and U3738 (N_3738,N_3608,N_3654);
or U3739 (N_3739,N_3624,N_3690);
and U3740 (N_3740,N_3641,N_3633);
nand U3741 (N_3741,N_3684,N_3646);
nand U3742 (N_3742,N_3666,N_3610);
or U3743 (N_3743,N_3627,N_3620);
nor U3744 (N_3744,N_3691,N_3648);
and U3745 (N_3745,N_3658,N_3659);
xnor U3746 (N_3746,N_3683,N_3617);
nand U3747 (N_3747,N_3677,N_3649);
and U3748 (N_3748,N_3616,N_3625);
nor U3749 (N_3749,N_3623,N_3664);
and U3750 (N_3750,N_3676,N_3612);
nand U3751 (N_3751,N_3675,N_3638);
nor U3752 (N_3752,N_3625,N_3685);
and U3753 (N_3753,N_3667,N_3698);
nand U3754 (N_3754,N_3683,N_3649);
nand U3755 (N_3755,N_3658,N_3618);
nor U3756 (N_3756,N_3656,N_3647);
and U3757 (N_3757,N_3631,N_3634);
or U3758 (N_3758,N_3611,N_3660);
or U3759 (N_3759,N_3648,N_3692);
and U3760 (N_3760,N_3612,N_3660);
nor U3761 (N_3761,N_3642,N_3621);
nand U3762 (N_3762,N_3600,N_3613);
and U3763 (N_3763,N_3625,N_3661);
nand U3764 (N_3764,N_3610,N_3623);
or U3765 (N_3765,N_3679,N_3649);
nor U3766 (N_3766,N_3663,N_3647);
nor U3767 (N_3767,N_3633,N_3653);
nor U3768 (N_3768,N_3648,N_3602);
nor U3769 (N_3769,N_3632,N_3618);
nand U3770 (N_3770,N_3668,N_3639);
and U3771 (N_3771,N_3681,N_3649);
and U3772 (N_3772,N_3676,N_3680);
or U3773 (N_3773,N_3676,N_3609);
and U3774 (N_3774,N_3611,N_3602);
or U3775 (N_3775,N_3631,N_3635);
and U3776 (N_3776,N_3631,N_3662);
nand U3777 (N_3777,N_3672,N_3639);
nand U3778 (N_3778,N_3613,N_3615);
or U3779 (N_3779,N_3685,N_3603);
and U3780 (N_3780,N_3699,N_3604);
nand U3781 (N_3781,N_3694,N_3635);
and U3782 (N_3782,N_3655,N_3607);
nor U3783 (N_3783,N_3698,N_3675);
and U3784 (N_3784,N_3681,N_3606);
nor U3785 (N_3785,N_3667,N_3602);
or U3786 (N_3786,N_3693,N_3669);
nand U3787 (N_3787,N_3613,N_3638);
and U3788 (N_3788,N_3687,N_3605);
nand U3789 (N_3789,N_3619,N_3615);
nand U3790 (N_3790,N_3618,N_3636);
and U3791 (N_3791,N_3643,N_3650);
nor U3792 (N_3792,N_3613,N_3609);
nor U3793 (N_3793,N_3662,N_3644);
nand U3794 (N_3794,N_3654,N_3693);
or U3795 (N_3795,N_3696,N_3621);
or U3796 (N_3796,N_3668,N_3653);
nor U3797 (N_3797,N_3672,N_3667);
or U3798 (N_3798,N_3639,N_3643);
or U3799 (N_3799,N_3689,N_3655);
nand U3800 (N_3800,N_3726,N_3771);
or U3801 (N_3801,N_3796,N_3709);
nand U3802 (N_3802,N_3795,N_3743);
nand U3803 (N_3803,N_3770,N_3721);
and U3804 (N_3804,N_3786,N_3780);
nand U3805 (N_3805,N_3753,N_3792);
nor U3806 (N_3806,N_3711,N_3798);
nor U3807 (N_3807,N_3791,N_3778);
and U3808 (N_3808,N_3751,N_3730);
and U3809 (N_3809,N_3738,N_3745);
nand U3810 (N_3810,N_3723,N_3799);
or U3811 (N_3811,N_3732,N_3757);
or U3812 (N_3812,N_3740,N_3765);
nor U3813 (N_3813,N_3719,N_3772);
or U3814 (N_3814,N_3735,N_3737);
nor U3815 (N_3815,N_3766,N_3702);
and U3816 (N_3816,N_3731,N_3742);
nand U3817 (N_3817,N_3750,N_3705);
nor U3818 (N_3818,N_3774,N_3769);
nor U3819 (N_3819,N_3787,N_3734);
nor U3820 (N_3820,N_3728,N_3718);
or U3821 (N_3821,N_3785,N_3748);
and U3822 (N_3822,N_3788,N_3746);
and U3823 (N_3823,N_3704,N_3777);
or U3824 (N_3824,N_3763,N_3717);
and U3825 (N_3825,N_3720,N_3700);
nor U3826 (N_3826,N_3794,N_3790);
and U3827 (N_3827,N_3782,N_3755);
or U3828 (N_3828,N_3760,N_3716);
and U3829 (N_3829,N_3736,N_3758);
and U3830 (N_3830,N_3725,N_3775);
and U3831 (N_3831,N_3789,N_3797);
and U3832 (N_3832,N_3701,N_3722);
nand U3833 (N_3833,N_3714,N_3713);
and U3834 (N_3834,N_3761,N_3781);
or U3835 (N_3835,N_3773,N_3741);
nor U3836 (N_3836,N_3724,N_3707);
nand U3837 (N_3837,N_3747,N_3779);
xnor U3838 (N_3838,N_3703,N_3784);
and U3839 (N_3839,N_3729,N_3708);
nand U3840 (N_3840,N_3754,N_3752);
or U3841 (N_3841,N_3793,N_3727);
or U3842 (N_3842,N_3733,N_3756);
nor U3843 (N_3843,N_3749,N_3744);
or U3844 (N_3844,N_3783,N_3762);
or U3845 (N_3845,N_3764,N_3712);
nor U3846 (N_3846,N_3739,N_3776);
nand U3847 (N_3847,N_3710,N_3767);
or U3848 (N_3848,N_3715,N_3768);
nor U3849 (N_3849,N_3759,N_3706);
or U3850 (N_3850,N_3756,N_3730);
and U3851 (N_3851,N_3778,N_3770);
nand U3852 (N_3852,N_3761,N_3786);
or U3853 (N_3853,N_3716,N_3783);
and U3854 (N_3854,N_3752,N_3721);
nor U3855 (N_3855,N_3787,N_3713);
nand U3856 (N_3856,N_3776,N_3729);
and U3857 (N_3857,N_3706,N_3729);
and U3858 (N_3858,N_3722,N_3715);
nand U3859 (N_3859,N_3783,N_3722);
nand U3860 (N_3860,N_3743,N_3777);
nand U3861 (N_3861,N_3745,N_3755);
nand U3862 (N_3862,N_3726,N_3738);
nor U3863 (N_3863,N_3793,N_3788);
and U3864 (N_3864,N_3723,N_3767);
nor U3865 (N_3865,N_3793,N_3715);
or U3866 (N_3866,N_3701,N_3794);
nor U3867 (N_3867,N_3745,N_3767);
and U3868 (N_3868,N_3768,N_3707);
nor U3869 (N_3869,N_3715,N_3781);
nor U3870 (N_3870,N_3714,N_3717);
nor U3871 (N_3871,N_3716,N_3720);
nor U3872 (N_3872,N_3723,N_3741);
nand U3873 (N_3873,N_3728,N_3778);
nor U3874 (N_3874,N_3754,N_3758);
and U3875 (N_3875,N_3705,N_3760);
or U3876 (N_3876,N_3784,N_3750);
and U3877 (N_3877,N_3784,N_3765);
nor U3878 (N_3878,N_3786,N_3721);
and U3879 (N_3879,N_3789,N_3783);
xor U3880 (N_3880,N_3744,N_3705);
or U3881 (N_3881,N_3737,N_3739);
nor U3882 (N_3882,N_3708,N_3789);
xnor U3883 (N_3883,N_3758,N_3738);
nor U3884 (N_3884,N_3737,N_3755);
nand U3885 (N_3885,N_3782,N_3767);
and U3886 (N_3886,N_3775,N_3771);
or U3887 (N_3887,N_3731,N_3774);
or U3888 (N_3888,N_3792,N_3762);
or U3889 (N_3889,N_3702,N_3771);
or U3890 (N_3890,N_3780,N_3747);
and U3891 (N_3891,N_3795,N_3746);
nand U3892 (N_3892,N_3759,N_3709);
or U3893 (N_3893,N_3730,N_3721);
and U3894 (N_3894,N_3770,N_3756);
nor U3895 (N_3895,N_3789,N_3750);
nand U3896 (N_3896,N_3728,N_3738);
nor U3897 (N_3897,N_3796,N_3790);
nand U3898 (N_3898,N_3784,N_3799);
nand U3899 (N_3899,N_3732,N_3725);
nand U3900 (N_3900,N_3876,N_3814);
and U3901 (N_3901,N_3888,N_3816);
nor U3902 (N_3902,N_3813,N_3829);
nor U3903 (N_3903,N_3810,N_3800);
or U3904 (N_3904,N_3834,N_3818);
nand U3905 (N_3905,N_3866,N_3828);
and U3906 (N_3906,N_3808,N_3820);
or U3907 (N_3907,N_3862,N_3805);
nor U3908 (N_3908,N_3826,N_3833);
or U3909 (N_3909,N_3847,N_3863);
or U3910 (N_3910,N_3822,N_3899);
and U3911 (N_3911,N_3883,N_3864);
nand U3912 (N_3912,N_3880,N_3853);
or U3913 (N_3913,N_3801,N_3850);
nand U3914 (N_3914,N_3804,N_3841);
nor U3915 (N_3915,N_3849,N_3815);
or U3916 (N_3916,N_3823,N_3858);
nor U3917 (N_3917,N_3869,N_3836);
and U3918 (N_3918,N_3885,N_3806);
nor U3919 (N_3919,N_3868,N_3803);
nor U3920 (N_3920,N_3879,N_3898);
or U3921 (N_3921,N_3838,N_3846);
or U3922 (N_3922,N_3819,N_3835);
and U3923 (N_3923,N_3892,N_3854);
and U3924 (N_3924,N_3875,N_3860);
and U3925 (N_3925,N_3889,N_3881);
and U3926 (N_3926,N_3891,N_3857);
nor U3927 (N_3927,N_3845,N_3837);
and U3928 (N_3928,N_3855,N_3830);
and U3929 (N_3929,N_3832,N_3852);
or U3930 (N_3930,N_3895,N_3861);
and U3931 (N_3931,N_3843,N_3894);
and U3932 (N_3932,N_3831,N_3886);
nand U3933 (N_3933,N_3807,N_3827);
nand U3934 (N_3934,N_3839,N_3817);
nand U3935 (N_3935,N_3851,N_3856);
and U3936 (N_3936,N_3865,N_3884);
nor U3937 (N_3937,N_3872,N_3844);
nand U3938 (N_3938,N_3887,N_3874);
xor U3939 (N_3939,N_3859,N_3871);
nor U3940 (N_3940,N_3848,N_3897);
nand U3941 (N_3941,N_3890,N_3842);
nand U3942 (N_3942,N_3824,N_3802);
and U3943 (N_3943,N_3877,N_3825);
or U3944 (N_3944,N_3812,N_3811);
nand U3945 (N_3945,N_3867,N_3870);
or U3946 (N_3946,N_3878,N_3882);
nor U3947 (N_3947,N_3821,N_3873);
or U3948 (N_3948,N_3809,N_3896);
and U3949 (N_3949,N_3893,N_3840);
and U3950 (N_3950,N_3837,N_3824);
and U3951 (N_3951,N_3850,N_3865);
nor U3952 (N_3952,N_3873,N_3884);
nor U3953 (N_3953,N_3838,N_3835);
and U3954 (N_3954,N_3876,N_3811);
nand U3955 (N_3955,N_3837,N_3885);
nand U3956 (N_3956,N_3871,N_3854);
nand U3957 (N_3957,N_3829,N_3840);
and U3958 (N_3958,N_3834,N_3823);
nand U3959 (N_3959,N_3845,N_3831);
or U3960 (N_3960,N_3843,N_3886);
and U3961 (N_3961,N_3881,N_3856);
nor U3962 (N_3962,N_3883,N_3823);
nor U3963 (N_3963,N_3879,N_3868);
and U3964 (N_3964,N_3877,N_3807);
and U3965 (N_3965,N_3867,N_3895);
or U3966 (N_3966,N_3858,N_3891);
or U3967 (N_3967,N_3861,N_3825);
and U3968 (N_3968,N_3894,N_3820);
or U3969 (N_3969,N_3882,N_3822);
nand U3970 (N_3970,N_3865,N_3828);
nor U3971 (N_3971,N_3872,N_3833);
nand U3972 (N_3972,N_3822,N_3832);
xnor U3973 (N_3973,N_3873,N_3828);
and U3974 (N_3974,N_3830,N_3874);
and U3975 (N_3975,N_3884,N_3864);
nor U3976 (N_3976,N_3812,N_3876);
nor U3977 (N_3977,N_3853,N_3898);
or U3978 (N_3978,N_3856,N_3891);
and U3979 (N_3979,N_3802,N_3833);
nor U3980 (N_3980,N_3821,N_3841);
or U3981 (N_3981,N_3844,N_3839);
or U3982 (N_3982,N_3883,N_3824);
and U3983 (N_3983,N_3855,N_3814);
nor U3984 (N_3984,N_3805,N_3893);
and U3985 (N_3985,N_3837,N_3847);
nor U3986 (N_3986,N_3868,N_3827);
or U3987 (N_3987,N_3853,N_3804);
nor U3988 (N_3988,N_3803,N_3865);
nor U3989 (N_3989,N_3837,N_3844);
or U3990 (N_3990,N_3880,N_3898);
nor U3991 (N_3991,N_3828,N_3877);
nor U3992 (N_3992,N_3815,N_3805);
and U3993 (N_3993,N_3821,N_3899);
and U3994 (N_3994,N_3884,N_3899);
or U3995 (N_3995,N_3838,N_3866);
and U3996 (N_3996,N_3853,N_3824);
nor U3997 (N_3997,N_3819,N_3828);
and U3998 (N_3998,N_3866,N_3827);
nand U3999 (N_3999,N_3832,N_3866);
nor U4000 (N_4000,N_3906,N_3905);
or U4001 (N_4001,N_3935,N_3968);
nand U4002 (N_4002,N_3930,N_3931);
nor U4003 (N_4003,N_3948,N_3945);
nand U4004 (N_4004,N_3916,N_3972);
and U4005 (N_4005,N_3953,N_3942);
or U4006 (N_4006,N_3951,N_3977);
or U4007 (N_4007,N_3970,N_3964);
nor U4008 (N_4008,N_3940,N_3903);
nor U4009 (N_4009,N_3941,N_3901);
or U4010 (N_4010,N_3909,N_3947);
and U4011 (N_4011,N_3933,N_3936);
and U4012 (N_4012,N_3912,N_3969);
and U4013 (N_4013,N_3934,N_3959);
or U4014 (N_4014,N_3961,N_3928);
or U4015 (N_4015,N_3975,N_3985);
nand U4016 (N_4016,N_3925,N_3954);
nor U4017 (N_4017,N_3996,N_3918);
nand U4018 (N_4018,N_3990,N_3913);
nand U4019 (N_4019,N_3956,N_3910);
and U4020 (N_4020,N_3908,N_3929);
or U4021 (N_4021,N_3900,N_3960);
and U4022 (N_4022,N_3920,N_3965);
and U4023 (N_4023,N_3938,N_3962);
nor U4024 (N_4024,N_3997,N_3995);
or U4025 (N_4025,N_3988,N_3994);
nand U4026 (N_4026,N_3999,N_3957);
and U4027 (N_4027,N_3949,N_3915);
xnor U4028 (N_4028,N_3958,N_3989);
nor U4029 (N_4029,N_3981,N_3932);
nor U4030 (N_4030,N_3982,N_3907);
nor U4031 (N_4031,N_3998,N_3939);
nor U4032 (N_4032,N_3986,N_3921);
or U4033 (N_4033,N_3919,N_3978);
and U4034 (N_4034,N_3902,N_3944);
or U4035 (N_4035,N_3966,N_3923);
and U4036 (N_4036,N_3926,N_3984);
nand U4037 (N_4037,N_3987,N_3971);
nor U4038 (N_4038,N_3937,N_3927);
nand U4039 (N_4039,N_3973,N_3924);
xor U4040 (N_4040,N_3922,N_3983);
nand U4041 (N_4041,N_3946,N_3911);
nand U4042 (N_4042,N_3976,N_3950);
nor U4043 (N_4043,N_3917,N_3993);
nor U4044 (N_4044,N_3963,N_3914);
and U4045 (N_4045,N_3974,N_3991);
or U4046 (N_4046,N_3967,N_3904);
and U4047 (N_4047,N_3955,N_3979);
nor U4048 (N_4048,N_3943,N_3952);
nand U4049 (N_4049,N_3992,N_3980);
nor U4050 (N_4050,N_3941,N_3993);
and U4051 (N_4051,N_3912,N_3932);
nand U4052 (N_4052,N_3969,N_3953);
or U4053 (N_4053,N_3918,N_3904);
or U4054 (N_4054,N_3939,N_3920);
nand U4055 (N_4055,N_3973,N_3911);
nor U4056 (N_4056,N_3938,N_3908);
nor U4057 (N_4057,N_3980,N_3977);
nand U4058 (N_4058,N_3947,N_3979);
nor U4059 (N_4059,N_3939,N_3966);
nand U4060 (N_4060,N_3928,N_3904);
and U4061 (N_4061,N_3926,N_3908);
and U4062 (N_4062,N_3932,N_3909);
or U4063 (N_4063,N_3936,N_3920);
nand U4064 (N_4064,N_3990,N_3932);
or U4065 (N_4065,N_3944,N_3962);
and U4066 (N_4066,N_3921,N_3990);
and U4067 (N_4067,N_3940,N_3901);
or U4068 (N_4068,N_3951,N_3947);
nor U4069 (N_4069,N_3955,N_3957);
or U4070 (N_4070,N_3982,N_3942);
or U4071 (N_4071,N_3930,N_3915);
and U4072 (N_4072,N_3946,N_3976);
or U4073 (N_4073,N_3976,N_3909);
or U4074 (N_4074,N_3951,N_3948);
nand U4075 (N_4075,N_3995,N_3973);
and U4076 (N_4076,N_3962,N_3910);
nor U4077 (N_4077,N_3947,N_3945);
and U4078 (N_4078,N_3945,N_3910);
nor U4079 (N_4079,N_3928,N_3908);
and U4080 (N_4080,N_3938,N_3924);
nor U4081 (N_4081,N_3931,N_3964);
nor U4082 (N_4082,N_3920,N_3962);
and U4083 (N_4083,N_3984,N_3906);
or U4084 (N_4084,N_3951,N_3991);
and U4085 (N_4085,N_3936,N_3956);
nor U4086 (N_4086,N_3985,N_3935);
and U4087 (N_4087,N_3991,N_3935);
and U4088 (N_4088,N_3944,N_3937);
nand U4089 (N_4089,N_3972,N_3987);
and U4090 (N_4090,N_3970,N_3960);
or U4091 (N_4091,N_3971,N_3903);
nor U4092 (N_4092,N_3968,N_3932);
nand U4093 (N_4093,N_3982,N_3941);
and U4094 (N_4094,N_3925,N_3951);
and U4095 (N_4095,N_3964,N_3980);
nand U4096 (N_4096,N_3914,N_3934);
nor U4097 (N_4097,N_3930,N_3939);
nor U4098 (N_4098,N_3927,N_3976);
or U4099 (N_4099,N_3933,N_3992);
and U4100 (N_4100,N_4027,N_4095);
or U4101 (N_4101,N_4010,N_4087);
or U4102 (N_4102,N_4053,N_4046);
and U4103 (N_4103,N_4011,N_4018);
nand U4104 (N_4104,N_4093,N_4050);
and U4105 (N_4105,N_4075,N_4073);
nor U4106 (N_4106,N_4031,N_4012);
and U4107 (N_4107,N_4054,N_4005);
and U4108 (N_4108,N_4070,N_4091);
and U4109 (N_4109,N_4056,N_4035);
or U4110 (N_4110,N_4017,N_4066);
and U4111 (N_4111,N_4055,N_4041);
and U4112 (N_4112,N_4030,N_4077);
nand U4113 (N_4113,N_4076,N_4088);
or U4114 (N_4114,N_4081,N_4084);
or U4115 (N_4115,N_4045,N_4057);
or U4116 (N_4116,N_4047,N_4092);
nor U4117 (N_4117,N_4067,N_4021);
and U4118 (N_4118,N_4000,N_4072);
nand U4119 (N_4119,N_4090,N_4007);
nand U4120 (N_4120,N_4025,N_4097);
nand U4121 (N_4121,N_4079,N_4006);
or U4122 (N_4122,N_4028,N_4032);
xor U4123 (N_4123,N_4002,N_4082);
or U4124 (N_4124,N_4065,N_4034);
and U4125 (N_4125,N_4022,N_4023);
or U4126 (N_4126,N_4004,N_4029);
and U4127 (N_4127,N_4051,N_4060);
or U4128 (N_4128,N_4009,N_4015);
nor U4129 (N_4129,N_4042,N_4052);
nand U4130 (N_4130,N_4094,N_4098);
nand U4131 (N_4131,N_4099,N_4024);
nand U4132 (N_4132,N_4074,N_4020);
or U4133 (N_4133,N_4083,N_4068);
or U4134 (N_4134,N_4078,N_4064);
nor U4135 (N_4135,N_4036,N_4016);
nand U4136 (N_4136,N_4049,N_4003);
nor U4137 (N_4137,N_4019,N_4040);
nand U4138 (N_4138,N_4039,N_4013);
or U4139 (N_4139,N_4048,N_4026);
and U4140 (N_4140,N_4089,N_4043);
nor U4141 (N_4141,N_4062,N_4071);
nor U4142 (N_4142,N_4008,N_4038);
nand U4143 (N_4143,N_4044,N_4033);
nor U4144 (N_4144,N_4085,N_4014);
nor U4145 (N_4145,N_4037,N_4059);
and U4146 (N_4146,N_4061,N_4096);
nor U4147 (N_4147,N_4058,N_4086);
nand U4148 (N_4148,N_4069,N_4001);
and U4149 (N_4149,N_4080,N_4063);
and U4150 (N_4150,N_4053,N_4036);
nor U4151 (N_4151,N_4016,N_4092);
nor U4152 (N_4152,N_4068,N_4019);
nand U4153 (N_4153,N_4032,N_4009);
and U4154 (N_4154,N_4038,N_4080);
nand U4155 (N_4155,N_4039,N_4021);
nand U4156 (N_4156,N_4050,N_4021);
or U4157 (N_4157,N_4082,N_4084);
or U4158 (N_4158,N_4051,N_4098);
nand U4159 (N_4159,N_4058,N_4089);
nor U4160 (N_4160,N_4052,N_4027);
and U4161 (N_4161,N_4075,N_4068);
or U4162 (N_4162,N_4013,N_4047);
and U4163 (N_4163,N_4036,N_4063);
or U4164 (N_4164,N_4035,N_4073);
nand U4165 (N_4165,N_4085,N_4031);
nor U4166 (N_4166,N_4084,N_4027);
nor U4167 (N_4167,N_4020,N_4069);
nor U4168 (N_4168,N_4000,N_4011);
or U4169 (N_4169,N_4009,N_4092);
nand U4170 (N_4170,N_4044,N_4079);
nor U4171 (N_4171,N_4049,N_4036);
nor U4172 (N_4172,N_4046,N_4056);
and U4173 (N_4173,N_4044,N_4011);
or U4174 (N_4174,N_4020,N_4019);
nor U4175 (N_4175,N_4007,N_4020);
nand U4176 (N_4176,N_4071,N_4051);
nand U4177 (N_4177,N_4007,N_4014);
nand U4178 (N_4178,N_4017,N_4039);
or U4179 (N_4179,N_4003,N_4039);
and U4180 (N_4180,N_4030,N_4083);
nand U4181 (N_4181,N_4070,N_4060);
nand U4182 (N_4182,N_4044,N_4030);
nor U4183 (N_4183,N_4072,N_4039);
nor U4184 (N_4184,N_4019,N_4038);
or U4185 (N_4185,N_4078,N_4072);
and U4186 (N_4186,N_4097,N_4053);
or U4187 (N_4187,N_4080,N_4046);
nand U4188 (N_4188,N_4076,N_4008);
or U4189 (N_4189,N_4074,N_4084);
and U4190 (N_4190,N_4047,N_4039);
and U4191 (N_4191,N_4043,N_4051);
nand U4192 (N_4192,N_4018,N_4041);
or U4193 (N_4193,N_4088,N_4011);
or U4194 (N_4194,N_4055,N_4027);
nor U4195 (N_4195,N_4080,N_4068);
nor U4196 (N_4196,N_4067,N_4025);
or U4197 (N_4197,N_4094,N_4036);
or U4198 (N_4198,N_4005,N_4048);
nand U4199 (N_4199,N_4032,N_4076);
and U4200 (N_4200,N_4148,N_4174);
and U4201 (N_4201,N_4155,N_4121);
nor U4202 (N_4202,N_4194,N_4100);
or U4203 (N_4203,N_4182,N_4188);
or U4204 (N_4204,N_4109,N_4179);
or U4205 (N_4205,N_4125,N_4161);
nor U4206 (N_4206,N_4167,N_4163);
nor U4207 (N_4207,N_4172,N_4169);
and U4208 (N_4208,N_4127,N_4110);
nand U4209 (N_4209,N_4142,N_4158);
nor U4210 (N_4210,N_4160,N_4187);
or U4211 (N_4211,N_4137,N_4101);
nand U4212 (N_4212,N_4126,N_4146);
and U4213 (N_4213,N_4135,N_4189);
or U4214 (N_4214,N_4143,N_4139);
nand U4215 (N_4215,N_4173,N_4128);
nand U4216 (N_4216,N_4131,N_4168);
or U4217 (N_4217,N_4176,N_4104);
or U4218 (N_4218,N_4198,N_4145);
nor U4219 (N_4219,N_4113,N_4193);
or U4220 (N_4220,N_4154,N_4156);
nand U4221 (N_4221,N_4181,N_4153);
and U4222 (N_4222,N_4196,N_4134);
nand U4223 (N_4223,N_4195,N_4190);
or U4224 (N_4224,N_4183,N_4149);
or U4225 (N_4225,N_4197,N_4150);
nand U4226 (N_4226,N_4122,N_4152);
nand U4227 (N_4227,N_4118,N_4114);
and U4228 (N_4228,N_4120,N_4186);
or U4229 (N_4229,N_4103,N_4138);
and U4230 (N_4230,N_4166,N_4151);
or U4231 (N_4231,N_4105,N_4171);
nand U4232 (N_4232,N_4165,N_4164);
nor U4233 (N_4233,N_4116,N_4129);
and U4234 (N_4234,N_4123,N_4136);
or U4235 (N_4235,N_4185,N_4147);
nand U4236 (N_4236,N_4117,N_4111);
or U4237 (N_4237,N_4124,N_4170);
and U4238 (N_4238,N_4107,N_4112);
or U4239 (N_4239,N_4140,N_4157);
and U4240 (N_4240,N_4108,N_4119);
and U4241 (N_4241,N_4133,N_4184);
nand U4242 (N_4242,N_4144,N_4177);
nor U4243 (N_4243,N_4106,N_4199);
nor U4244 (N_4244,N_4162,N_4115);
or U4245 (N_4245,N_4180,N_4141);
nand U4246 (N_4246,N_4191,N_4102);
or U4247 (N_4247,N_4175,N_4192);
or U4248 (N_4248,N_4178,N_4159);
and U4249 (N_4249,N_4130,N_4132);
or U4250 (N_4250,N_4133,N_4189);
and U4251 (N_4251,N_4179,N_4101);
nor U4252 (N_4252,N_4139,N_4179);
or U4253 (N_4253,N_4156,N_4153);
or U4254 (N_4254,N_4162,N_4176);
nor U4255 (N_4255,N_4130,N_4139);
xor U4256 (N_4256,N_4107,N_4137);
xnor U4257 (N_4257,N_4116,N_4115);
and U4258 (N_4258,N_4135,N_4119);
or U4259 (N_4259,N_4159,N_4128);
and U4260 (N_4260,N_4128,N_4162);
nor U4261 (N_4261,N_4141,N_4139);
and U4262 (N_4262,N_4182,N_4155);
nor U4263 (N_4263,N_4124,N_4103);
nand U4264 (N_4264,N_4109,N_4163);
and U4265 (N_4265,N_4156,N_4112);
nand U4266 (N_4266,N_4125,N_4173);
or U4267 (N_4267,N_4135,N_4145);
and U4268 (N_4268,N_4110,N_4180);
or U4269 (N_4269,N_4168,N_4116);
nand U4270 (N_4270,N_4159,N_4168);
and U4271 (N_4271,N_4147,N_4170);
nand U4272 (N_4272,N_4175,N_4117);
nor U4273 (N_4273,N_4178,N_4163);
and U4274 (N_4274,N_4135,N_4157);
nor U4275 (N_4275,N_4161,N_4170);
or U4276 (N_4276,N_4137,N_4142);
and U4277 (N_4277,N_4195,N_4146);
nor U4278 (N_4278,N_4188,N_4150);
nor U4279 (N_4279,N_4109,N_4124);
nand U4280 (N_4280,N_4133,N_4110);
and U4281 (N_4281,N_4114,N_4133);
or U4282 (N_4282,N_4149,N_4166);
and U4283 (N_4283,N_4171,N_4199);
nor U4284 (N_4284,N_4106,N_4193);
or U4285 (N_4285,N_4184,N_4143);
nand U4286 (N_4286,N_4146,N_4192);
and U4287 (N_4287,N_4168,N_4169);
or U4288 (N_4288,N_4110,N_4164);
nor U4289 (N_4289,N_4186,N_4157);
and U4290 (N_4290,N_4112,N_4118);
or U4291 (N_4291,N_4134,N_4102);
and U4292 (N_4292,N_4132,N_4169);
or U4293 (N_4293,N_4108,N_4167);
and U4294 (N_4294,N_4189,N_4115);
nand U4295 (N_4295,N_4149,N_4117);
or U4296 (N_4296,N_4189,N_4100);
nor U4297 (N_4297,N_4116,N_4120);
and U4298 (N_4298,N_4140,N_4103);
or U4299 (N_4299,N_4163,N_4104);
xnor U4300 (N_4300,N_4215,N_4262);
and U4301 (N_4301,N_4264,N_4288);
and U4302 (N_4302,N_4290,N_4242);
nor U4303 (N_4303,N_4225,N_4258);
xnor U4304 (N_4304,N_4236,N_4287);
or U4305 (N_4305,N_4220,N_4248);
nand U4306 (N_4306,N_4255,N_4200);
and U4307 (N_4307,N_4274,N_4231);
nand U4308 (N_4308,N_4284,N_4240);
xnor U4309 (N_4309,N_4203,N_4279);
nor U4310 (N_4310,N_4273,N_4235);
or U4311 (N_4311,N_4283,N_4252);
nand U4312 (N_4312,N_4210,N_4232);
or U4313 (N_4313,N_4239,N_4263);
nor U4314 (N_4314,N_4265,N_4269);
nor U4315 (N_4315,N_4238,N_4268);
or U4316 (N_4316,N_4295,N_4272);
nand U4317 (N_4317,N_4243,N_4297);
nor U4318 (N_4318,N_4233,N_4204);
or U4319 (N_4319,N_4219,N_4271);
nand U4320 (N_4320,N_4213,N_4275);
nand U4321 (N_4321,N_4223,N_4276);
nand U4322 (N_4322,N_4205,N_4254);
nand U4323 (N_4323,N_4292,N_4230);
or U4324 (N_4324,N_4299,N_4244);
and U4325 (N_4325,N_4209,N_4208);
and U4326 (N_4326,N_4266,N_4257);
and U4327 (N_4327,N_4237,N_4222);
and U4328 (N_4328,N_4251,N_4250);
and U4329 (N_4329,N_4286,N_4277);
and U4330 (N_4330,N_4216,N_4256);
and U4331 (N_4331,N_4278,N_4247);
or U4332 (N_4332,N_4259,N_4212);
nor U4333 (N_4333,N_4298,N_4280);
and U4334 (N_4334,N_4228,N_4217);
nor U4335 (N_4335,N_4294,N_4221);
nor U4336 (N_4336,N_4282,N_4207);
or U4337 (N_4337,N_4234,N_4291);
or U4338 (N_4338,N_4293,N_4214);
nor U4339 (N_4339,N_4227,N_4246);
nor U4340 (N_4340,N_4206,N_4201);
nor U4341 (N_4341,N_4267,N_4218);
and U4342 (N_4342,N_4289,N_4281);
or U4343 (N_4343,N_4253,N_4285);
nor U4344 (N_4344,N_4226,N_4224);
nand U4345 (N_4345,N_4296,N_4241);
nand U4346 (N_4346,N_4270,N_4229);
or U4347 (N_4347,N_4260,N_4202);
and U4348 (N_4348,N_4245,N_4249);
or U4349 (N_4349,N_4261,N_4211);
or U4350 (N_4350,N_4263,N_4207);
and U4351 (N_4351,N_4289,N_4245);
and U4352 (N_4352,N_4211,N_4224);
nand U4353 (N_4353,N_4220,N_4263);
or U4354 (N_4354,N_4263,N_4287);
and U4355 (N_4355,N_4284,N_4279);
and U4356 (N_4356,N_4243,N_4281);
nand U4357 (N_4357,N_4231,N_4203);
or U4358 (N_4358,N_4223,N_4208);
nand U4359 (N_4359,N_4247,N_4222);
nand U4360 (N_4360,N_4215,N_4212);
nor U4361 (N_4361,N_4292,N_4236);
and U4362 (N_4362,N_4201,N_4296);
nor U4363 (N_4363,N_4237,N_4280);
or U4364 (N_4364,N_4255,N_4219);
nand U4365 (N_4365,N_4236,N_4215);
or U4366 (N_4366,N_4293,N_4278);
and U4367 (N_4367,N_4283,N_4269);
or U4368 (N_4368,N_4285,N_4271);
nor U4369 (N_4369,N_4222,N_4280);
or U4370 (N_4370,N_4230,N_4235);
and U4371 (N_4371,N_4208,N_4213);
or U4372 (N_4372,N_4206,N_4243);
and U4373 (N_4373,N_4297,N_4231);
nand U4374 (N_4374,N_4270,N_4213);
nand U4375 (N_4375,N_4213,N_4274);
and U4376 (N_4376,N_4235,N_4221);
and U4377 (N_4377,N_4289,N_4214);
nand U4378 (N_4378,N_4282,N_4213);
nor U4379 (N_4379,N_4228,N_4211);
nor U4380 (N_4380,N_4232,N_4265);
nand U4381 (N_4381,N_4253,N_4205);
or U4382 (N_4382,N_4243,N_4220);
or U4383 (N_4383,N_4262,N_4257);
nand U4384 (N_4384,N_4282,N_4263);
nand U4385 (N_4385,N_4279,N_4229);
nor U4386 (N_4386,N_4262,N_4284);
nor U4387 (N_4387,N_4270,N_4261);
nor U4388 (N_4388,N_4262,N_4233);
and U4389 (N_4389,N_4221,N_4213);
nand U4390 (N_4390,N_4223,N_4291);
nor U4391 (N_4391,N_4212,N_4245);
nor U4392 (N_4392,N_4256,N_4226);
nand U4393 (N_4393,N_4276,N_4218);
nor U4394 (N_4394,N_4269,N_4241);
or U4395 (N_4395,N_4290,N_4245);
and U4396 (N_4396,N_4216,N_4236);
nor U4397 (N_4397,N_4251,N_4229);
nor U4398 (N_4398,N_4254,N_4248);
and U4399 (N_4399,N_4246,N_4287);
or U4400 (N_4400,N_4389,N_4390);
or U4401 (N_4401,N_4355,N_4314);
or U4402 (N_4402,N_4338,N_4317);
and U4403 (N_4403,N_4304,N_4363);
and U4404 (N_4404,N_4313,N_4375);
and U4405 (N_4405,N_4386,N_4398);
and U4406 (N_4406,N_4336,N_4309);
nand U4407 (N_4407,N_4394,N_4372);
or U4408 (N_4408,N_4347,N_4315);
nor U4409 (N_4409,N_4345,N_4301);
or U4410 (N_4410,N_4340,N_4388);
nor U4411 (N_4411,N_4332,N_4391);
and U4412 (N_4412,N_4361,N_4341);
nand U4413 (N_4413,N_4342,N_4376);
or U4414 (N_4414,N_4353,N_4343);
and U4415 (N_4415,N_4371,N_4331);
or U4416 (N_4416,N_4365,N_4378);
or U4417 (N_4417,N_4377,N_4333);
or U4418 (N_4418,N_4381,N_4323);
or U4419 (N_4419,N_4370,N_4351);
nor U4420 (N_4420,N_4369,N_4397);
nand U4421 (N_4421,N_4360,N_4362);
nor U4422 (N_4422,N_4325,N_4348);
nand U4423 (N_4423,N_4344,N_4352);
nand U4424 (N_4424,N_4319,N_4380);
or U4425 (N_4425,N_4316,N_4357);
or U4426 (N_4426,N_4393,N_4327);
nor U4427 (N_4427,N_4373,N_4382);
and U4428 (N_4428,N_4328,N_4311);
nand U4429 (N_4429,N_4359,N_4392);
and U4430 (N_4430,N_4334,N_4395);
and U4431 (N_4431,N_4366,N_4308);
and U4432 (N_4432,N_4396,N_4337);
nor U4433 (N_4433,N_4330,N_4368);
nand U4434 (N_4434,N_4318,N_4322);
or U4435 (N_4435,N_4320,N_4374);
and U4436 (N_4436,N_4302,N_4310);
nor U4437 (N_4437,N_4329,N_4358);
nor U4438 (N_4438,N_4324,N_4356);
nand U4439 (N_4439,N_4321,N_4307);
or U4440 (N_4440,N_4350,N_4367);
or U4441 (N_4441,N_4305,N_4349);
nand U4442 (N_4442,N_4312,N_4384);
nand U4443 (N_4443,N_4346,N_4387);
nand U4444 (N_4444,N_4306,N_4335);
and U4445 (N_4445,N_4339,N_4364);
nand U4446 (N_4446,N_4383,N_4354);
nand U4447 (N_4447,N_4326,N_4385);
or U4448 (N_4448,N_4303,N_4399);
and U4449 (N_4449,N_4300,N_4379);
and U4450 (N_4450,N_4345,N_4379);
and U4451 (N_4451,N_4303,N_4383);
or U4452 (N_4452,N_4384,N_4345);
or U4453 (N_4453,N_4321,N_4311);
or U4454 (N_4454,N_4371,N_4361);
or U4455 (N_4455,N_4385,N_4376);
and U4456 (N_4456,N_4351,N_4396);
or U4457 (N_4457,N_4324,N_4345);
and U4458 (N_4458,N_4397,N_4364);
nand U4459 (N_4459,N_4306,N_4321);
and U4460 (N_4460,N_4388,N_4356);
nor U4461 (N_4461,N_4392,N_4303);
nor U4462 (N_4462,N_4345,N_4387);
and U4463 (N_4463,N_4342,N_4389);
nor U4464 (N_4464,N_4385,N_4350);
nor U4465 (N_4465,N_4303,N_4309);
and U4466 (N_4466,N_4390,N_4342);
or U4467 (N_4467,N_4325,N_4363);
and U4468 (N_4468,N_4311,N_4347);
and U4469 (N_4469,N_4381,N_4380);
and U4470 (N_4470,N_4371,N_4315);
or U4471 (N_4471,N_4302,N_4304);
nand U4472 (N_4472,N_4353,N_4326);
nor U4473 (N_4473,N_4311,N_4366);
or U4474 (N_4474,N_4378,N_4361);
and U4475 (N_4475,N_4395,N_4303);
or U4476 (N_4476,N_4355,N_4312);
nor U4477 (N_4477,N_4319,N_4303);
nor U4478 (N_4478,N_4324,N_4301);
or U4479 (N_4479,N_4380,N_4357);
nor U4480 (N_4480,N_4348,N_4384);
and U4481 (N_4481,N_4340,N_4327);
nand U4482 (N_4482,N_4373,N_4312);
or U4483 (N_4483,N_4399,N_4338);
or U4484 (N_4484,N_4388,N_4396);
and U4485 (N_4485,N_4314,N_4388);
or U4486 (N_4486,N_4302,N_4368);
nand U4487 (N_4487,N_4311,N_4308);
and U4488 (N_4488,N_4398,N_4357);
or U4489 (N_4489,N_4364,N_4306);
nor U4490 (N_4490,N_4316,N_4342);
and U4491 (N_4491,N_4333,N_4312);
nor U4492 (N_4492,N_4327,N_4361);
nor U4493 (N_4493,N_4355,N_4389);
nand U4494 (N_4494,N_4365,N_4356);
nand U4495 (N_4495,N_4347,N_4303);
or U4496 (N_4496,N_4321,N_4394);
nand U4497 (N_4497,N_4306,N_4369);
or U4498 (N_4498,N_4320,N_4382);
or U4499 (N_4499,N_4341,N_4306);
nand U4500 (N_4500,N_4470,N_4434);
nor U4501 (N_4501,N_4452,N_4489);
nor U4502 (N_4502,N_4408,N_4497);
nor U4503 (N_4503,N_4411,N_4436);
nand U4504 (N_4504,N_4413,N_4400);
nor U4505 (N_4505,N_4499,N_4402);
nor U4506 (N_4506,N_4473,N_4433);
and U4507 (N_4507,N_4430,N_4485);
nor U4508 (N_4508,N_4403,N_4409);
or U4509 (N_4509,N_4492,N_4468);
nand U4510 (N_4510,N_4460,N_4426);
and U4511 (N_4511,N_4466,N_4440);
and U4512 (N_4512,N_4478,N_4459);
or U4513 (N_4513,N_4476,N_4447);
nor U4514 (N_4514,N_4417,N_4421);
and U4515 (N_4515,N_4483,N_4463);
and U4516 (N_4516,N_4423,N_4446);
nand U4517 (N_4517,N_4450,N_4406);
or U4518 (N_4518,N_4401,N_4456);
nand U4519 (N_4519,N_4441,N_4458);
or U4520 (N_4520,N_4484,N_4453);
nand U4521 (N_4521,N_4474,N_4491);
nor U4522 (N_4522,N_4418,N_4419);
and U4523 (N_4523,N_4486,N_4455);
nand U4524 (N_4524,N_4429,N_4444);
and U4525 (N_4525,N_4449,N_4439);
nand U4526 (N_4526,N_4465,N_4487);
nor U4527 (N_4527,N_4425,N_4480);
or U4528 (N_4528,N_4495,N_4442);
nor U4529 (N_4529,N_4431,N_4404);
and U4530 (N_4530,N_4490,N_4405);
or U4531 (N_4531,N_4414,N_4472);
nand U4532 (N_4532,N_4479,N_4475);
and U4533 (N_4533,N_4428,N_4469);
nor U4534 (N_4534,N_4443,N_4420);
nor U4535 (N_4535,N_4438,N_4427);
nor U4536 (N_4536,N_4445,N_4407);
or U4537 (N_4537,N_4424,N_4432);
and U4538 (N_4538,N_4494,N_4464);
or U4539 (N_4539,N_4454,N_4496);
nand U4540 (N_4540,N_4477,N_4488);
nor U4541 (N_4541,N_4435,N_4493);
and U4542 (N_4542,N_4481,N_4467);
and U4543 (N_4543,N_4471,N_4410);
nor U4544 (N_4544,N_4448,N_4422);
or U4545 (N_4545,N_4457,N_4462);
and U4546 (N_4546,N_4461,N_4416);
and U4547 (N_4547,N_4482,N_4498);
nand U4548 (N_4548,N_4415,N_4451);
or U4549 (N_4549,N_4412,N_4437);
nand U4550 (N_4550,N_4465,N_4428);
nand U4551 (N_4551,N_4465,N_4490);
or U4552 (N_4552,N_4412,N_4401);
or U4553 (N_4553,N_4443,N_4461);
nor U4554 (N_4554,N_4473,N_4458);
nor U4555 (N_4555,N_4416,N_4411);
or U4556 (N_4556,N_4400,N_4448);
or U4557 (N_4557,N_4449,N_4400);
or U4558 (N_4558,N_4405,N_4429);
nor U4559 (N_4559,N_4447,N_4419);
nand U4560 (N_4560,N_4427,N_4422);
nand U4561 (N_4561,N_4410,N_4418);
and U4562 (N_4562,N_4438,N_4458);
nor U4563 (N_4563,N_4426,N_4450);
nand U4564 (N_4564,N_4458,N_4426);
nor U4565 (N_4565,N_4451,N_4432);
and U4566 (N_4566,N_4410,N_4486);
nand U4567 (N_4567,N_4437,N_4440);
nor U4568 (N_4568,N_4415,N_4426);
nand U4569 (N_4569,N_4405,N_4433);
nand U4570 (N_4570,N_4469,N_4476);
nor U4571 (N_4571,N_4440,N_4406);
or U4572 (N_4572,N_4418,N_4422);
nor U4573 (N_4573,N_4413,N_4429);
and U4574 (N_4574,N_4467,N_4474);
xnor U4575 (N_4575,N_4484,N_4424);
nor U4576 (N_4576,N_4410,N_4484);
nand U4577 (N_4577,N_4499,N_4487);
xnor U4578 (N_4578,N_4415,N_4468);
and U4579 (N_4579,N_4452,N_4445);
nand U4580 (N_4580,N_4453,N_4427);
and U4581 (N_4581,N_4409,N_4479);
and U4582 (N_4582,N_4482,N_4423);
and U4583 (N_4583,N_4488,N_4438);
and U4584 (N_4584,N_4461,N_4424);
nand U4585 (N_4585,N_4421,N_4404);
or U4586 (N_4586,N_4401,N_4422);
nor U4587 (N_4587,N_4460,N_4452);
nor U4588 (N_4588,N_4403,N_4472);
nor U4589 (N_4589,N_4476,N_4481);
or U4590 (N_4590,N_4438,N_4407);
nor U4591 (N_4591,N_4410,N_4402);
and U4592 (N_4592,N_4488,N_4417);
and U4593 (N_4593,N_4437,N_4484);
nand U4594 (N_4594,N_4402,N_4490);
or U4595 (N_4595,N_4410,N_4462);
nand U4596 (N_4596,N_4443,N_4472);
nor U4597 (N_4597,N_4432,N_4439);
nor U4598 (N_4598,N_4480,N_4471);
nor U4599 (N_4599,N_4465,N_4414);
or U4600 (N_4600,N_4524,N_4578);
and U4601 (N_4601,N_4555,N_4503);
or U4602 (N_4602,N_4595,N_4550);
or U4603 (N_4603,N_4553,N_4552);
or U4604 (N_4604,N_4585,N_4587);
and U4605 (N_4605,N_4518,N_4547);
nand U4606 (N_4606,N_4565,N_4525);
nor U4607 (N_4607,N_4516,N_4544);
nand U4608 (N_4608,N_4599,N_4536);
nor U4609 (N_4609,N_4582,N_4515);
nor U4610 (N_4610,N_4566,N_4590);
nor U4611 (N_4611,N_4513,N_4532);
nor U4612 (N_4612,N_4558,N_4569);
xnor U4613 (N_4613,N_4589,N_4546);
and U4614 (N_4614,N_4548,N_4531);
nor U4615 (N_4615,N_4593,N_4564);
or U4616 (N_4616,N_4511,N_4586);
or U4617 (N_4617,N_4522,N_4562);
or U4618 (N_4618,N_4554,N_4551);
and U4619 (N_4619,N_4567,N_4584);
and U4620 (N_4620,N_4523,N_4514);
or U4621 (N_4621,N_4530,N_4542);
or U4622 (N_4622,N_4537,N_4538);
nor U4623 (N_4623,N_4570,N_4594);
nand U4624 (N_4624,N_4543,N_4533);
nor U4625 (N_4625,N_4520,N_4568);
or U4626 (N_4626,N_4541,N_4576);
and U4627 (N_4627,N_4574,N_4592);
and U4628 (N_4628,N_4539,N_4598);
nor U4629 (N_4629,N_4540,N_4529);
nor U4630 (N_4630,N_4577,N_4561);
nand U4631 (N_4631,N_4507,N_4559);
or U4632 (N_4632,N_4583,N_4591);
nor U4633 (N_4633,N_4596,N_4512);
and U4634 (N_4634,N_4560,N_4517);
nand U4635 (N_4635,N_4573,N_4509);
and U4636 (N_4636,N_4501,N_4579);
nand U4637 (N_4637,N_4528,N_4556);
nand U4638 (N_4638,N_4575,N_4597);
nor U4639 (N_4639,N_4500,N_4534);
nand U4640 (N_4640,N_4505,N_4504);
and U4641 (N_4641,N_4549,N_4526);
nand U4642 (N_4642,N_4535,N_4510);
or U4643 (N_4643,N_4527,N_4521);
nor U4644 (N_4644,N_4588,N_4572);
or U4645 (N_4645,N_4506,N_4580);
and U4646 (N_4646,N_4545,N_4563);
and U4647 (N_4647,N_4508,N_4557);
nor U4648 (N_4648,N_4519,N_4571);
or U4649 (N_4649,N_4502,N_4581);
and U4650 (N_4650,N_4554,N_4525);
and U4651 (N_4651,N_4507,N_4593);
nor U4652 (N_4652,N_4549,N_4564);
nand U4653 (N_4653,N_4549,N_4586);
nor U4654 (N_4654,N_4546,N_4500);
and U4655 (N_4655,N_4599,N_4592);
and U4656 (N_4656,N_4564,N_4514);
nand U4657 (N_4657,N_4558,N_4500);
and U4658 (N_4658,N_4546,N_4592);
nor U4659 (N_4659,N_4593,N_4545);
or U4660 (N_4660,N_4581,N_4591);
and U4661 (N_4661,N_4588,N_4510);
nor U4662 (N_4662,N_4542,N_4534);
nand U4663 (N_4663,N_4578,N_4504);
or U4664 (N_4664,N_4590,N_4571);
or U4665 (N_4665,N_4575,N_4594);
nand U4666 (N_4666,N_4517,N_4543);
nor U4667 (N_4667,N_4580,N_4594);
and U4668 (N_4668,N_4561,N_4520);
and U4669 (N_4669,N_4504,N_4569);
nand U4670 (N_4670,N_4599,N_4556);
or U4671 (N_4671,N_4568,N_4543);
and U4672 (N_4672,N_4516,N_4581);
xnor U4673 (N_4673,N_4595,N_4572);
nor U4674 (N_4674,N_4588,N_4543);
nor U4675 (N_4675,N_4513,N_4510);
and U4676 (N_4676,N_4529,N_4536);
and U4677 (N_4677,N_4590,N_4514);
or U4678 (N_4678,N_4517,N_4525);
or U4679 (N_4679,N_4539,N_4538);
nor U4680 (N_4680,N_4548,N_4592);
nand U4681 (N_4681,N_4564,N_4577);
nand U4682 (N_4682,N_4548,N_4527);
nand U4683 (N_4683,N_4567,N_4539);
nor U4684 (N_4684,N_4568,N_4521);
nand U4685 (N_4685,N_4555,N_4540);
and U4686 (N_4686,N_4535,N_4565);
nand U4687 (N_4687,N_4589,N_4576);
nor U4688 (N_4688,N_4582,N_4547);
or U4689 (N_4689,N_4589,N_4540);
nand U4690 (N_4690,N_4550,N_4588);
nor U4691 (N_4691,N_4520,N_4572);
nor U4692 (N_4692,N_4531,N_4573);
nand U4693 (N_4693,N_4595,N_4537);
or U4694 (N_4694,N_4557,N_4518);
nand U4695 (N_4695,N_4519,N_4559);
nand U4696 (N_4696,N_4547,N_4599);
xor U4697 (N_4697,N_4571,N_4540);
nor U4698 (N_4698,N_4593,N_4542);
nor U4699 (N_4699,N_4536,N_4520);
nor U4700 (N_4700,N_4620,N_4692);
nand U4701 (N_4701,N_4630,N_4629);
nor U4702 (N_4702,N_4635,N_4636);
nand U4703 (N_4703,N_4662,N_4698);
and U4704 (N_4704,N_4677,N_4697);
and U4705 (N_4705,N_4661,N_4628);
or U4706 (N_4706,N_4648,N_4615);
and U4707 (N_4707,N_4601,N_4600);
or U4708 (N_4708,N_4666,N_4606);
nor U4709 (N_4709,N_4689,N_4667);
nand U4710 (N_4710,N_4610,N_4619);
nand U4711 (N_4711,N_4611,N_4690);
nand U4712 (N_4712,N_4694,N_4656);
and U4713 (N_4713,N_4634,N_4678);
or U4714 (N_4714,N_4608,N_4602);
and U4715 (N_4715,N_4655,N_4642);
and U4716 (N_4716,N_4604,N_4699);
nor U4717 (N_4717,N_4652,N_4663);
nor U4718 (N_4718,N_4673,N_4668);
nand U4719 (N_4719,N_4681,N_4609);
or U4720 (N_4720,N_4633,N_4646);
nor U4721 (N_4721,N_4679,N_4624);
nand U4722 (N_4722,N_4685,N_4641);
and U4723 (N_4723,N_4644,N_4674);
nand U4724 (N_4724,N_4675,N_4603);
and U4725 (N_4725,N_4613,N_4664);
or U4726 (N_4726,N_4639,N_4682);
or U4727 (N_4727,N_4658,N_4625);
and U4728 (N_4728,N_4627,N_4612);
or U4729 (N_4729,N_4680,N_4622);
nand U4730 (N_4730,N_4614,N_4695);
nand U4731 (N_4731,N_4657,N_4649);
nor U4732 (N_4732,N_4638,N_4686);
or U4733 (N_4733,N_4653,N_4691);
nor U4734 (N_4734,N_4659,N_4616);
or U4735 (N_4735,N_4672,N_4637);
nor U4736 (N_4736,N_4626,N_4670);
and U4737 (N_4737,N_4650,N_4643);
or U4738 (N_4738,N_4671,N_4618);
nand U4739 (N_4739,N_4617,N_4631);
nand U4740 (N_4740,N_4669,N_4696);
and U4741 (N_4741,N_4688,N_4621);
nor U4742 (N_4742,N_4645,N_4683);
nor U4743 (N_4743,N_4693,N_4654);
nand U4744 (N_4744,N_4684,N_4647);
nand U4745 (N_4745,N_4623,N_4660);
or U4746 (N_4746,N_4607,N_4665);
nand U4747 (N_4747,N_4651,N_4605);
nand U4748 (N_4748,N_4640,N_4687);
nor U4749 (N_4749,N_4676,N_4632);
or U4750 (N_4750,N_4613,N_4608);
nor U4751 (N_4751,N_4644,N_4677);
nor U4752 (N_4752,N_4613,N_4615);
or U4753 (N_4753,N_4633,N_4617);
nor U4754 (N_4754,N_4672,N_4628);
or U4755 (N_4755,N_4626,N_4651);
nand U4756 (N_4756,N_4631,N_4604);
nand U4757 (N_4757,N_4636,N_4662);
or U4758 (N_4758,N_4644,N_4645);
or U4759 (N_4759,N_4679,N_4622);
or U4760 (N_4760,N_4663,N_4619);
or U4761 (N_4761,N_4656,N_4664);
nor U4762 (N_4762,N_4641,N_4625);
or U4763 (N_4763,N_4622,N_4687);
and U4764 (N_4764,N_4694,N_4624);
or U4765 (N_4765,N_4684,N_4672);
nand U4766 (N_4766,N_4686,N_4641);
and U4767 (N_4767,N_4696,N_4676);
and U4768 (N_4768,N_4610,N_4683);
nand U4769 (N_4769,N_4652,N_4675);
nand U4770 (N_4770,N_4655,N_4665);
nand U4771 (N_4771,N_4612,N_4673);
and U4772 (N_4772,N_4651,N_4638);
nand U4773 (N_4773,N_4696,N_4663);
nand U4774 (N_4774,N_4622,N_4672);
or U4775 (N_4775,N_4613,N_4649);
nand U4776 (N_4776,N_4649,N_4698);
or U4777 (N_4777,N_4677,N_4626);
nand U4778 (N_4778,N_4638,N_4645);
or U4779 (N_4779,N_4610,N_4681);
and U4780 (N_4780,N_4643,N_4630);
and U4781 (N_4781,N_4646,N_4642);
and U4782 (N_4782,N_4616,N_4600);
nand U4783 (N_4783,N_4603,N_4638);
or U4784 (N_4784,N_4613,N_4684);
nand U4785 (N_4785,N_4669,N_4613);
nand U4786 (N_4786,N_4682,N_4608);
nor U4787 (N_4787,N_4691,N_4679);
and U4788 (N_4788,N_4681,N_4615);
nor U4789 (N_4789,N_4644,N_4648);
and U4790 (N_4790,N_4662,N_4601);
and U4791 (N_4791,N_4628,N_4655);
nor U4792 (N_4792,N_4671,N_4673);
nand U4793 (N_4793,N_4690,N_4693);
nand U4794 (N_4794,N_4616,N_4612);
xnor U4795 (N_4795,N_4636,N_4677);
and U4796 (N_4796,N_4689,N_4668);
or U4797 (N_4797,N_4642,N_4622);
or U4798 (N_4798,N_4625,N_4673);
or U4799 (N_4799,N_4682,N_4643);
and U4800 (N_4800,N_4742,N_4722);
xor U4801 (N_4801,N_4733,N_4710);
or U4802 (N_4802,N_4796,N_4781);
nor U4803 (N_4803,N_4758,N_4789);
nor U4804 (N_4804,N_4790,N_4754);
or U4805 (N_4805,N_4721,N_4746);
or U4806 (N_4806,N_4798,N_4731);
or U4807 (N_4807,N_4704,N_4776);
or U4808 (N_4808,N_4719,N_4730);
and U4809 (N_4809,N_4755,N_4744);
or U4810 (N_4810,N_4727,N_4720);
nor U4811 (N_4811,N_4784,N_4786);
nand U4812 (N_4812,N_4708,N_4797);
nor U4813 (N_4813,N_4734,N_4769);
nor U4814 (N_4814,N_4768,N_4773);
and U4815 (N_4815,N_4702,N_4703);
nor U4816 (N_4816,N_4756,N_4737);
or U4817 (N_4817,N_4766,N_4767);
nor U4818 (N_4818,N_4739,N_4771);
and U4819 (N_4819,N_4774,N_4757);
nor U4820 (N_4820,N_4750,N_4788);
and U4821 (N_4821,N_4794,N_4782);
and U4822 (N_4822,N_4752,N_4792);
or U4823 (N_4823,N_4785,N_4772);
and U4824 (N_4824,N_4743,N_4759);
or U4825 (N_4825,N_4749,N_4783);
or U4826 (N_4826,N_4723,N_4748);
and U4827 (N_4827,N_4740,N_4716);
nand U4828 (N_4828,N_4700,N_4793);
and U4829 (N_4829,N_4717,N_4764);
nor U4830 (N_4830,N_4777,N_4711);
nor U4831 (N_4831,N_4795,N_4726);
nand U4832 (N_4832,N_4718,N_4762);
or U4833 (N_4833,N_4770,N_4706);
nand U4834 (N_4834,N_4741,N_4715);
and U4835 (N_4835,N_4763,N_4724);
or U4836 (N_4836,N_4736,N_4761);
nand U4837 (N_4837,N_4751,N_4765);
and U4838 (N_4838,N_4701,N_4787);
or U4839 (N_4839,N_4729,N_4799);
nand U4840 (N_4840,N_4745,N_4728);
nor U4841 (N_4841,N_4779,N_4778);
or U4842 (N_4842,N_4713,N_4753);
nor U4843 (N_4843,N_4760,N_4747);
or U4844 (N_4844,N_4775,N_4709);
and U4845 (N_4845,N_4714,N_4780);
nand U4846 (N_4846,N_4738,N_4705);
nand U4847 (N_4847,N_4725,N_4791);
nor U4848 (N_4848,N_4712,N_4732);
and U4849 (N_4849,N_4735,N_4707);
nor U4850 (N_4850,N_4704,N_4714);
nand U4851 (N_4851,N_4780,N_4724);
nor U4852 (N_4852,N_4712,N_4797);
or U4853 (N_4853,N_4719,N_4749);
nor U4854 (N_4854,N_4796,N_4754);
and U4855 (N_4855,N_4792,N_4722);
nor U4856 (N_4856,N_4772,N_4782);
or U4857 (N_4857,N_4722,N_4712);
or U4858 (N_4858,N_4797,N_4737);
nand U4859 (N_4859,N_4725,N_4702);
and U4860 (N_4860,N_4790,N_4788);
nand U4861 (N_4861,N_4743,N_4739);
and U4862 (N_4862,N_4734,N_4794);
or U4863 (N_4863,N_4760,N_4766);
nand U4864 (N_4864,N_4758,N_4774);
or U4865 (N_4865,N_4745,N_4782);
nand U4866 (N_4866,N_4774,N_4779);
and U4867 (N_4867,N_4705,N_4785);
or U4868 (N_4868,N_4787,N_4717);
nor U4869 (N_4869,N_4799,N_4756);
and U4870 (N_4870,N_4769,N_4708);
or U4871 (N_4871,N_4744,N_4775);
and U4872 (N_4872,N_4748,N_4710);
and U4873 (N_4873,N_4703,N_4777);
nand U4874 (N_4874,N_4702,N_4755);
nand U4875 (N_4875,N_4741,N_4796);
nand U4876 (N_4876,N_4740,N_4794);
or U4877 (N_4877,N_4761,N_4784);
or U4878 (N_4878,N_4702,N_4784);
nand U4879 (N_4879,N_4783,N_4734);
nor U4880 (N_4880,N_4703,N_4752);
and U4881 (N_4881,N_4789,N_4724);
and U4882 (N_4882,N_4774,N_4700);
nor U4883 (N_4883,N_4770,N_4793);
and U4884 (N_4884,N_4738,N_4789);
and U4885 (N_4885,N_4765,N_4752);
nor U4886 (N_4886,N_4733,N_4782);
nor U4887 (N_4887,N_4711,N_4745);
or U4888 (N_4888,N_4737,N_4759);
nor U4889 (N_4889,N_4711,N_4707);
nor U4890 (N_4890,N_4721,N_4773);
and U4891 (N_4891,N_4760,N_4786);
nand U4892 (N_4892,N_4791,N_4775);
or U4893 (N_4893,N_4706,N_4702);
and U4894 (N_4894,N_4793,N_4767);
nor U4895 (N_4895,N_4708,N_4721);
nor U4896 (N_4896,N_4752,N_4788);
nand U4897 (N_4897,N_4718,N_4736);
or U4898 (N_4898,N_4777,N_4728);
and U4899 (N_4899,N_4775,N_4733);
and U4900 (N_4900,N_4806,N_4873);
or U4901 (N_4901,N_4889,N_4897);
or U4902 (N_4902,N_4899,N_4832);
nand U4903 (N_4903,N_4828,N_4801);
nand U4904 (N_4904,N_4893,N_4850);
nor U4905 (N_4905,N_4840,N_4898);
and U4906 (N_4906,N_4821,N_4862);
nor U4907 (N_4907,N_4831,N_4812);
and U4908 (N_4908,N_4884,N_4849);
or U4909 (N_4909,N_4867,N_4854);
nand U4910 (N_4910,N_4891,N_4800);
nor U4911 (N_4911,N_4835,N_4841);
and U4912 (N_4912,N_4846,N_4857);
nor U4913 (N_4913,N_4853,N_4880);
nand U4914 (N_4914,N_4834,N_4804);
and U4915 (N_4915,N_4874,N_4878);
and U4916 (N_4916,N_4805,N_4895);
nor U4917 (N_4917,N_4845,N_4870);
nor U4918 (N_4918,N_4839,N_4843);
nand U4919 (N_4919,N_4819,N_4861);
and U4920 (N_4920,N_4872,N_4852);
and U4921 (N_4921,N_4875,N_4815);
or U4922 (N_4922,N_4816,N_4881);
nor U4923 (N_4923,N_4856,N_4825);
nor U4924 (N_4924,N_4887,N_4820);
or U4925 (N_4925,N_4838,N_4892);
nand U4926 (N_4926,N_4822,N_4866);
or U4927 (N_4927,N_4869,N_4871);
nor U4928 (N_4928,N_4859,N_4829);
nor U4929 (N_4929,N_4847,N_4817);
or U4930 (N_4930,N_4809,N_4811);
and U4931 (N_4931,N_4876,N_4848);
nor U4932 (N_4932,N_4810,N_4863);
nand U4933 (N_4933,N_4814,N_4836);
nor U4934 (N_4934,N_4833,N_4883);
or U4935 (N_4935,N_4827,N_4807);
or U4936 (N_4936,N_4858,N_4888);
or U4937 (N_4937,N_4885,N_4890);
and U4938 (N_4938,N_4879,N_4864);
or U4939 (N_4939,N_4802,N_4824);
or U4940 (N_4940,N_4860,N_4855);
and U4941 (N_4941,N_4830,N_4886);
and U4942 (N_4942,N_4868,N_4882);
nor U4943 (N_4943,N_4818,N_4844);
nand U4944 (N_4944,N_4851,N_4865);
or U4945 (N_4945,N_4877,N_4842);
and U4946 (N_4946,N_4823,N_4826);
nor U4947 (N_4947,N_4813,N_4808);
nor U4948 (N_4948,N_4896,N_4894);
and U4949 (N_4949,N_4837,N_4803);
and U4950 (N_4950,N_4816,N_4849);
or U4951 (N_4951,N_4892,N_4822);
nand U4952 (N_4952,N_4876,N_4852);
nor U4953 (N_4953,N_4851,N_4807);
xor U4954 (N_4954,N_4895,N_4817);
or U4955 (N_4955,N_4878,N_4828);
or U4956 (N_4956,N_4882,N_4835);
nor U4957 (N_4957,N_4872,N_4803);
nand U4958 (N_4958,N_4810,N_4867);
or U4959 (N_4959,N_4854,N_4819);
or U4960 (N_4960,N_4898,N_4836);
and U4961 (N_4961,N_4850,N_4848);
nand U4962 (N_4962,N_4876,N_4896);
nand U4963 (N_4963,N_4875,N_4806);
or U4964 (N_4964,N_4880,N_4845);
or U4965 (N_4965,N_4899,N_4824);
nor U4966 (N_4966,N_4848,N_4812);
nor U4967 (N_4967,N_4812,N_4804);
nand U4968 (N_4968,N_4818,N_4857);
or U4969 (N_4969,N_4854,N_4862);
nand U4970 (N_4970,N_4811,N_4854);
nor U4971 (N_4971,N_4813,N_4823);
or U4972 (N_4972,N_4899,N_4800);
and U4973 (N_4973,N_4841,N_4802);
nor U4974 (N_4974,N_4844,N_4802);
nor U4975 (N_4975,N_4806,N_4866);
or U4976 (N_4976,N_4849,N_4818);
nand U4977 (N_4977,N_4811,N_4838);
and U4978 (N_4978,N_4822,N_4893);
nor U4979 (N_4979,N_4878,N_4863);
nand U4980 (N_4980,N_4802,N_4800);
nand U4981 (N_4981,N_4883,N_4809);
nand U4982 (N_4982,N_4832,N_4848);
and U4983 (N_4983,N_4806,N_4893);
nand U4984 (N_4984,N_4880,N_4823);
nand U4985 (N_4985,N_4890,N_4862);
nand U4986 (N_4986,N_4803,N_4806);
or U4987 (N_4987,N_4870,N_4820);
nand U4988 (N_4988,N_4817,N_4858);
nor U4989 (N_4989,N_4834,N_4838);
nand U4990 (N_4990,N_4802,N_4850);
nand U4991 (N_4991,N_4835,N_4865);
or U4992 (N_4992,N_4826,N_4852);
nand U4993 (N_4993,N_4815,N_4809);
or U4994 (N_4994,N_4896,N_4844);
nand U4995 (N_4995,N_4803,N_4825);
nand U4996 (N_4996,N_4884,N_4840);
nor U4997 (N_4997,N_4804,N_4847);
and U4998 (N_4998,N_4825,N_4849);
nor U4999 (N_4999,N_4873,N_4842);
nand U5000 (N_5000,N_4990,N_4972);
nand U5001 (N_5001,N_4902,N_4935);
nor U5002 (N_5002,N_4939,N_4904);
and U5003 (N_5003,N_4978,N_4970);
and U5004 (N_5004,N_4998,N_4958);
nor U5005 (N_5005,N_4937,N_4924);
nor U5006 (N_5006,N_4999,N_4919);
nor U5007 (N_5007,N_4986,N_4992);
and U5008 (N_5008,N_4965,N_4964);
or U5009 (N_5009,N_4930,N_4967);
nor U5010 (N_5010,N_4980,N_4903);
nor U5011 (N_5011,N_4966,N_4934);
nor U5012 (N_5012,N_4963,N_4932);
or U5013 (N_5013,N_4982,N_4920);
nand U5014 (N_5014,N_4910,N_4951);
or U5015 (N_5015,N_4988,N_4907);
nor U5016 (N_5016,N_4914,N_4969);
and U5017 (N_5017,N_4906,N_4971);
nor U5018 (N_5018,N_4941,N_4947);
nand U5019 (N_5019,N_4901,N_4912);
nor U5020 (N_5020,N_4926,N_4929);
or U5021 (N_5021,N_4962,N_4940);
or U5022 (N_5022,N_4949,N_4995);
and U5023 (N_5023,N_4994,N_4985);
or U5024 (N_5024,N_4960,N_4900);
and U5025 (N_5025,N_4957,N_4989);
and U5026 (N_5026,N_4931,N_4956);
nor U5027 (N_5027,N_4977,N_4959);
and U5028 (N_5028,N_4983,N_4950);
and U5029 (N_5029,N_4942,N_4954);
nor U5030 (N_5030,N_4984,N_4952);
nor U5031 (N_5031,N_4955,N_4943);
and U5032 (N_5032,N_4909,N_4973);
xnor U5033 (N_5033,N_4925,N_4968);
nand U5034 (N_5034,N_4915,N_4936);
nor U5035 (N_5035,N_4921,N_4991);
and U5036 (N_5036,N_4918,N_4928);
nor U5037 (N_5037,N_4938,N_4923);
nor U5038 (N_5038,N_4933,N_4913);
nand U5039 (N_5039,N_4961,N_4948);
nor U5040 (N_5040,N_4993,N_4996);
nor U5041 (N_5041,N_4927,N_4911);
nor U5042 (N_5042,N_4945,N_4922);
and U5043 (N_5043,N_4917,N_4987);
and U5044 (N_5044,N_4979,N_4916);
and U5045 (N_5045,N_4953,N_4975);
and U5046 (N_5046,N_4908,N_4905);
or U5047 (N_5047,N_4976,N_4997);
nor U5048 (N_5048,N_4974,N_4981);
nand U5049 (N_5049,N_4944,N_4946);
or U5050 (N_5050,N_4913,N_4981);
or U5051 (N_5051,N_4971,N_4944);
nor U5052 (N_5052,N_4960,N_4912);
nor U5053 (N_5053,N_4974,N_4982);
or U5054 (N_5054,N_4918,N_4965);
nand U5055 (N_5055,N_4978,N_4943);
nand U5056 (N_5056,N_4902,N_4958);
and U5057 (N_5057,N_4962,N_4992);
nor U5058 (N_5058,N_4943,N_4983);
or U5059 (N_5059,N_4901,N_4915);
and U5060 (N_5060,N_4943,N_4914);
or U5061 (N_5061,N_4984,N_4990);
and U5062 (N_5062,N_4973,N_4974);
nand U5063 (N_5063,N_4901,N_4951);
nor U5064 (N_5064,N_4990,N_4943);
and U5065 (N_5065,N_4987,N_4998);
nand U5066 (N_5066,N_4911,N_4975);
or U5067 (N_5067,N_4973,N_4944);
or U5068 (N_5068,N_4978,N_4919);
nand U5069 (N_5069,N_4926,N_4902);
or U5070 (N_5070,N_4908,N_4900);
nor U5071 (N_5071,N_4913,N_4977);
nor U5072 (N_5072,N_4901,N_4999);
nand U5073 (N_5073,N_4983,N_4916);
or U5074 (N_5074,N_4984,N_4944);
or U5075 (N_5075,N_4997,N_4915);
or U5076 (N_5076,N_4922,N_4946);
nor U5077 (N_5077,N_4974,N_4904);
or U5078 (N_5078,N_4911,N_4932);
nor U5079 (N_5079,N_4910,N_4919);
nor U5080 (N_5080,N_4904,N_4994);
nor U5081 (N_5081,N_4989,N_4988);
nand U5082 (N_5082,N_4949,N_4933);
or U5083 (N_5083,N_4951,N_4990);
and U5084 (N_5084,N_4958,N_4943);
nor U5085 (N_5085,N_4952,N_4920);
and U5086 (N_5086,N_4974,N_4993);
or U5087 (N_5087,N_4902,N_4979);
nand U5088 (N_5088,N_4954,N_4970);
and U5089 (N_5089,N_4972,N_4947);
and U5090 (N_5090,N_4970,N_4967);
nand U5091 (N_5091,N_4968,N_4999);
and U5092 (N_5092,N_4926,N_4964);
xnor U5093 (N_5093,N_4984,N_4938);
and U5094 (N_5094,N_4988,N_4965);
nor U5095 (N_5095,N_4915,N_4959);
or U5096 (N_5096,N_4996,N_4986);
or U5097 (N_5097,N_4958,N_4999);
and U5098 (N_5098,N_4950,N_4959);
and U5099 (N_5099,N_4955,N_4909);
nand U5100 (N_5100,N_5093,N_5096);
nand U5101 (N_5101,N_5049,N_5073);
or U5102 (N_5102,N_5026,N_5004);
nand U5103 (N_5103,N_5042,N_5092);
or U5104 (N_5104,N_5037,N_5031);
or U5105 (N_5105,N_5005,N_5057);
nand U5106 (N_5106,N_5063,N_5035);
and U5107 (N_5107,N_5008,N_5002);
or U5108 (N_5108,N_5065,N_5019);
nand U5109 (N_5109,N_5023,N_5082);
nand U5110 (N_5110,N_5059,N_5090);
nor U5111 (N_5111,N_5016,N_5034);
and U5112 (N_5112,N_5069,N_5064);
nor U5113 (N_5113,N_5044,N_5033);
nand U5114 (N_5114,N_5097,N_5085);
nand U5115 (N_5115,N_5055,N_5078);
nand U5116 (N_5116,N_5083,N_5017);
nand U5117 (N_5117,N_5025,N_5009);
nor U5118 (N_5118,N_5070,N_5077);
and U5119 (N_5119,N_5054,N_5013);
and U5120 (N_5120,N_5050,N_5071);
nand U5121 (N_5121,N_5036,N_5081);
or U5122 (N_5122,N_5053,N_5000);
and U5123 (N_5123,N_5074,N_5084);
and U5124 (N_5124,N_5014,N_5039);
nand U5125 (N_5125,N_5045,N_5068);
or U5126 (N_5126,N_5028,N_5091);
and U5127 (N_5127,N_5032,N_5046);
nand U5128 (N_5128,N_5024,N_5040);
nand U5129 (N_5129,N_5048,N_5021);
xnor U5130 (N_5130,N_5007,N_5003);
nand U5131 (N_5131,N_5094,N_5020);
and U5132 (N_5132,N_5011,N_5061);
and U5133 (N_5133,N_5047,N_5088);
nand U5134 (N_5134,N_5099,N_5038);
nor U5135 (N_5135,N_5027,N_5079);
or U5136 (N_5136,N_5066,N_5006);
and U5137 (N_5137,N_5072,N_5067);
nand U5138 (N_5138,N_5052,N_5058);
nand U5139 (N_5139,N_5087,N_5051);
nor U5140 (N_5140,N_5001,N_5043);
and U5141 (N_5141,N_5015,N_5029);
and U5142 (N_5142,N_5098,N_5095);
nand U5143 (N_5143,N_5075,N_5010);
or U5144 (N_5144,N_5056,N_5076);
nand U5145 (N_5145,N_5062,N_5041);
and U5146 (N_5146,N_5030,N_5060);
nor U5147 (N_5147,N_5089,N_5022);
or U5148 (N_5148,N_5018,N_5012);
nand U5149 (N_5149,N_5086,N_5080);
or U5150 (N_5150,N_5012,N_5072);
and U5151 (N_5151,N_5094,N_5084);
or U5152 (N_5152,N_5081,N_5051);
or U5153 (N_5153,N_5065,N_5040);
nand U5154 (N_5154,N_5030,N_5083);
and U5155 (N_5155,N_5076,N_5075);
nor U5156 (N_5156,N_5022,N_5059);
nor U5157 (N_5157,N_5038,N_5003);
and U5158 (N_5158,N_5040,N_5022);
and U5159 (N_5159,N_5004,N_5056);
nand U5160 (N_5160,N_5044,N_5087);
nor U5161 (N_5161,N_5093,N_5003);
nor U5162 (N_5162,N_5093,N_5009);
nor U5163 (N_5163,N_5090,N_5027);
nand U5164 (N_5164,N_5083,N_5070);
nand U5165 (N_5165,N_5022,N_5075);
and U5166 (N_5166,N_5046,N_5023);
nand U5167 (N_5167,N_5063,N_5097);
nand U5168 (N_5168,N_5038,N_5070);
nor U5169 (N_5169,N_5099,N_5089);
nor U5170 (N_5170,N_5035,N_5018);
or U5171 (N_5171,N_5087,N_5010);
nor U5172 (N_5172,N_5097,N_5066);
nor U5173 (N_5173,N_5040,N_5020);
nor U5174 (N_5174,N_5000,N_5046);
nand U5175 (N_5175,N_5095,N_5066);
nor U5176 (N_5176,N_5050,N_5034);
and U5177 (N_5177,N_5036,N_5018);
nor U5178 (N_5178,N_5059,N_5014);
and U5179 (N_5179,N_5052,N_5010);
and U5180 (N_5180,N_5022,N_5056);
nor U5181 (N_5181,N_5042,N_5009);
nand U5182 (N_5182,N_5083,N_5081);
nor U5183 (N_5183,N_5098,N_5037);
nand U5184 (N_5184,N_5030,N_5015);
and U5185 (N_5185,N_5072,N_5060);
or U5186 (N_5186,N_5060,N_5039);
and U5187 (N_5187,N_5079,N_5004);
and U5188 (N_5188,N_5027,N_5065);
nand U5189 (N_5189,N_5045,N_5083);
nand U5190 (N_5190,N_5029,N_5037);
and U5191 (N_5191,N_5017,N_5003);
or U5192 (N_5192,N_5060,N_5045);
or U5193 (N_5193,N_5092,N_5035);
nor U5194 (N_5194,N_5088,N_5083);
nand U5195 (N_5195,N_5082,N_5094);
and U5196 (N_5196,N_5019,N_5075);
or U5197 (N_5197,N_5084,N_5038);
or U5198 (N_5198,N_5081,N_5048);
nor U5199 (N_5199,N_5099,N_5016);
or U5200 (N_5200,N_5114,N_5193);
nand U5201 (N_5201,N_5189,N_5195);
or U5202 (N_5202,N_5153,N_5178);
and U5203 (N_5203,N_5108,N_5161);
nand U5204 (N_5204,N_5110,N_5147);
nor U5205 (N_5205,N_5182,N_5134);
or U5206 (N_5206,N_5177,N_5160);
nand U5207 (N_5207,N_5126,N_5164);
or U5208 (N_5208,N_5140,N_5112);
nor U5209 (N_5209,N_5124,N_5152);
or U5210 (N_5210,N_5101,N_5192);
nor U5211 (N_5211,N_5163,N_5165);
nor U5212 (N_5212,N_5106,N_5169);
nor U5213 (N_5213,N_5174,N_5118);
nand U5214 (N_5214,N_5107,N_5128);
nand U5215 (N_5215,N_5141,N_5132);
nor U5216 (N_5216,N_5183,N_5103);
nand U5217 (N_5217,N_5117,N_5127);
nor U5218 (N_5218,N_5149,N_5133);
nand U5219 (N_5219,N_5173,N_5186);
or U5220 (N_5220,N_5190,N_5199);
and U5221 (N_5221,N_5162,N_5129);
nor U5222 (N_5222,N_5187,N_5191);
nand U5223 (N_5223,N_5113,N_5179);
nor U5224 (N_5224,N_5185,N_5125);
nand U5225 (N_5225,N_5121,N_5100);
or U5226 (N_5226,N_5197,N_5138);
and U5227 (N_5227,N_5156,N_5154);
nor U5228 (N_5228,N_5181,N_5139);
and U5229 (N_5229,N_5196,N_5159);
nand U5230 (N_5230,N_5176,N_5198);
nor U5231 (N_5231,N_5170,N_5109);
nor U5232 (N_5232,N_5102,N_5172);
or U5233 (N_5233,N_5122,N_5180);
and U5234 (N_5234,N_5111,N_5168);
nand U5235 (N_5235,N_5135,N_5145);
or U5236 (N_5236,N_5155,N_5151);
nor U5237 (N_5237,N_5116,N_5157);
or U5238 (N_5238,N_5148,N_5105);
xnor U5239 (N_5239,N_5130,N_5123);
nor U5240 (N_5240,N_5150,N_5175);
nand U5241 (N_5241,N_5171,N_5144);
nor U5242 (N_5242,N_5142,N_5136);
or U5243 (N_5243,N_5167,N_5166);
or U5244 (N_5244,N_5146,N_5188);
xnor U5245 (N_5245,N_5131,N_5104);
nand U5246 (N_5246,N_5120,N_5143);
nand U5247 (N_5247,N_5184,N_5115);
and U5248 (N_5248,N_5119,N_5137);
and U5249 (N_5249,N_5194,N_5158);
nand U5250 (N_5250,N_5105,N_5165);
nor U5251 (N_5251,N_5163,N_5128);
nor U5252 (N_5252,N_5103,N_5190);
and U5253 (N_5253,N_5195,N_5178);
nand U5254 (N_5254,N_5173,N_5138);
or U5255 (N_5255,N_5102,N_5105);
and U5256 (N_5256,N_5182,N_5119);
or U5257 (N_5257,N_5152,N_5155);
and U5258 (N_5258,N_5164,N_5142);
and U5259 (N_5259,N_5145,N_5127);
nor U5260 (N_5260,N_5105,N_5167);
nor U5261 (N_5261,N_5149,N_5155);
and U5262 (N_5262,N_5105,N_5120);
or U5263 (N_5263,N_5199,N_5188);
nor U5264 (N_5264,N_5100,N_5165);
nand U5265 (N_5265,N_5111,N_5147);
and U5266 (N_5266,N_5122,N_5148);
nor U5267 (N_5267,N_5180,N_5133);
and U5268 (N_5268,N_5199,N_5173);
nor U5269 (N_5269,N_5140,N_5132);
nor U5270 (N_5270,N_5168,N_5148);
nand U5271 (N_5271,N_5162,N_5125);
and U5272 (N_5272,N_5138,N_5199);
or U5273 (N_5273,N_5156,N_5124);
or U5274 (N_5274,N_5170,N_5117);
or U5275 (N_5275,N_5141,N_5179);
nand U5276 (N_5276,N_5141,N_5192);
or U5277 (N_5277,N_5193,N_5146);
xor U5278 (N_5278,N_5104,N_5177);
nand U5279 (N_5279,N_5185,N_5141);
and U5280 (N_5280,N_5189,N_5187);
nor U5281 (N_5281,N_5183,N_5165);
or U5282 (N_5282,N_5166,N_5150);
or U5283 (N_5283,N_5195,N_5192);
or U5284 (N_5284,N_5164,N_5136);
nand U5285 (N_5285,N_5123,N_5149);
or U5286 (N_5286,N_5108,N_5153);
and U5287 (N_5287,N_5145,N_5174);
nand U5288 (N_5288,N_5119,N_5109);
nor U5289 (N_5289,N_5182,N_5133);
or U5290 (N_5290,N_5133,N_5115);
nor U5291 (N_5291,N_5186,N_5181);
or U5292 (N_5292,N_5180,N_5117);
and U5293 (N_5293,N_5104,N_5109);
or U5294 (N_5294,N_5103,N_5122);
and U5295 (N_5295,N_5194,N_5180);
or U5296 (N_5296,N_5106,N_5190);
and U5297 (N_5297,N_5178,N_5194);
or U5298 (N_5298,N_5154,N_5178);
nand U5299 (N_5299,N_5108,N_5198);
nor U5300 (N_5300,N_5216,N_5290);
and U5301 (N_5301,N_5268,N_5276);
or U5302 (N_5302,N_5248,N_5225);
nand U5303 (N_5303,N_5264,N_5230);
nand U5304 (N_5304,N_5223,N_5274);
and U5305 (N_5305,N_5210,N_5288);
nor U5306 (N_5306,N_5251,N_5218);
nor U5307 (N_5307,N_5203,N_5289);
or U5308 (N_5308,N_5281,N_5241);
nand U5309 (N_5309,N_5212,N_5227);
and U5310 (N_5310,N_5253,N_5220);
or U5311 (N_5311,N_5217,N_5242);
and U5312 (N_5312,N_5247,N_5243);
or U5313 (N_5313,N_5266,N_5226);
or U5314 (N_5314,N_5228,N_5263);
or U5315 (N_5315,N_5267,N_5273);
xor U5316 (N_5316,N_5272,N_5209);
nand U5317 (N_5317,N_5233,N_5238);
nor U5318 (N_5318,N_5255,N_5229);
xnor U5319 (N_5319,N_5222,N_5283);
nand U5320 (N_5320,N_5246,N_5256);
and U5321 (N_5321,N_5285,N_5239);
nor U5322 (N_5322,N_5284,N_5292);
and U5323 (N_5323,N_5234,N_5249);
or U5324 (N_5324,N_5250,N_5277);
or U5325 (N_5325,N_5282,N_5213);
nand U5326 (N_5326,N_5207,N_5236);
or U5327 (N_5327,N_5291,N_5245);
and U5328 (N_5328,N_5280,N_5299);
nor U5329 (N_5329,N_5270,N_5219);
and U5330 (N_5330,N_5293,N_5279);
and U5331 (N_5331,N_5224,N_5206);
nand U5332 (N_5332,N_5244,N_5278);
or U5333 (N_5333,N_5232,N_5231);
nand U5334 (N_5334,N_5262,N_5296);
or U5335 (N_5335,N_5254,N_5211);
nor U5336 (N_5336,N_5265,N_5235);
xnor U5337 (N_5337,N_5258,N_5205);
nand U5338 (N_5338,N_5237,N_5200);
nand U5339 (N_5339,N_5261,N_5202);
nor U5340 (N_5340,N_5252,N_5208);
nor U5341 (N_5341,N_5214,N_5221);
nand U5342 (N_5342,N_5287,N_5294);
or U5343 (N_5343,N_5240,N_5259);
or U5344 (N_5344,N_5201,N_5297);
and U5345 (N_5345,N_5257,N_5271);
and U5346 (N_5346,N_5286,N_5260);
nor U5347 (N_5347,N_5298,N_5204);
nor U5348 (N_5348,N_5295,N_5275);
nor U5349 (N_5349,N_5269,N_5215);
nand U5350 (N_5350,N_5257,N_5252);
or U5351 (N_5351,N_5275,N_5226);
nor U5352 (N_5352,N_5280,N_5290);
nor U5353 (N_5353,N_5237,N_5222);
and U5354 (N_5354,N_5273,N_5284);
nor U5355 (N_5355,N_5261,N_5240);
nor U5356 (N_5356,N_5238,N_5266);
and U5357 (N_5357,N_5293,N_5284);
nand U5358 (N_5358,N_5268,N_5287);
nand U5359 (N_5359,N_5201,N_5225);
and U5360 (N_5360,N_5265,N_5222);
and U5361 (N_5361,N_5206,N_5244);
nor U5362 (N_5362,N_5210,N_5229);
nor U5363 (N_5363,N_5255,N_5222);
or U5364 (N_5364,N_5266,N_5274);
or U5365 (N_5365,N_5290,N_5283);
nor U5366 (N_5366,N_5279,N_5204);
or U5367 (N_5367,N_5227,N_5263);
and U5368 (N_5368,N_5230,N_5294);
nor U5369 (N_5369,N_5236,N_5299);
and U5370 (N_5370,N_5202,N_5221);
nor U5371 (N_5371,N_5260,N_5296);
and U5372 (N_5372,N_5204,N_5216);
nor U5373 (N_5373,N_5203,N_5211);
nor U5374 (N_5374,N_5249,N_5236);
and U5375 (N_5375,N_5222,N_5285);
nor U5376 (N_5376,N_5284,N_5249);
nor U5377 (N_5377,N_5232,N_5281);
nand U5378 (N_5378,N_5276,N_5220);
nand U5379 (N_5379,N_5290,N_5254);
and U5380 (N_5380,N_5243,N_5294);
and U5381 (N_5381,N_5273,N_5240);
nand U5382 (N_5382,N_5277,N_5233);
and U5383 (N_5383,N_5243,N_5223);
and U5384 (N_5384,N_5287,N_5201);
and U5385 (N_5385,N_5242,N_5207);
or U5386 (N_5386,N_5220,N_5234);
or U5387 (N_5387,N_5236,N_5255);
nand U5388 (N_5388,N_5267,N_5269);
and U5389 (N_5389,N_5283,N_5200);
nand U5390 (N_5390,N_5241,N_5217);
nor U5391 (N_5391,N_5291,N_5202);
nor U5392 (N_5392,N_5218,N_5267);
nor U5393 (N_5393,N_5299,N_5275);
nor U5394 (N_5394,N_5214,N_5245);
nand U5395 (N_5395,N_5289,N_5261);
nand U5396 (N_5396,N_5253,N_5208);
nor U5397 (N_5397,N_5261,N_5247);
and U5398 (N_5398,N_5270,N_5283);
nor U5399 (N_5399,N_5297,N_5237);
nand U5400 (N_5400,N_5360,N_5378);
nand U5401 (N_5401,N_5388,N_5312);
and U5402 (N_5402,N_5343,N_5375);
or U5403 (N_5403,N_5361,N_5385);
and U5404 (N_5404,N_5397,N_5308);
and U5405 (N_5405,N_5354,N_5314);
or U5406 (N_5406,N_5326,N_5331);
nand U5407 (N_5407,N_5353,N_5323);
nor U5408 (N_5408,N_5368,N_5338);
nand U5409 (N_5409,N_5327,N_5339);
nand U5410 (N_5410,N_5356,N_5391);
nand U5411 (N_5411,N_5352,N_5381);
nand U5412 (N_5412,N_5351,N_5396);
or U5413 (N_5413,N_5382,N_5325);
or U5414 (N_5414,N_5377,N_5362);
nand U5415 (N_5415,N_5347,N_5334);
nand U5416 (N_5416,N_5380,N_5333);
or U5417 (N_5417,N_5317,N_5349);
or U5418 (N_5418,N_5320,N_5307);
nand U5419 (N_5419,N_5329,N_5379);
nand U5420 (N_5420,N_5364,N_5309);
nand U5421 (N_5421,N_5328,N_5336);
or U5422 (N_5422,N_5315,N_5366);
nand U5423 (N_5423,N_5393,N_5346);
nor U5424 (N_5424,N_5358,N_5370);
or U5425 (N_5425,N_5332,N_5373);
nand U5426 (N_5426,N_5340,N_5363);
or U5427 (N_5427,N_5344,N_5399);
and U5428 (N_5428,N_5310,N_5394);
nor U5429 (N_5429,N_5300,N_5355);
nand U5430 (N_5430,N_5335,N_5371);
and U5431 (N_5431,N_5383,N_5392);
and U5432 (N_5432,N_5345,N_5322);
and U5433 (N_5433,N_5348,N_5330);
and U5434 (N_5434,N_5390,N_5342);
or U5435 (N_5435,N_5374,N_5357);
or U5436 (N_5436,N_5367,N_5387);
nand U5437 (N_5437,N_5313,N_5319);
and U5438 (N_5438,N_5386,N_5318);
nand U5439 (N_5439,N_5376,N_5341);
nor U5440 (N_5440,N_5395,N_5337);
and U5441 (N_5441,N_5311,N_5359);
and U5442 (N_5442,N_5306,N_5305);
nand U5443 (N_5443,N_5384,N_5365);
or U5444 (N_5444,N_5389,N_5369);
or U5445 (N_5445,N_5316,N_5324);
nor U5446 (N_5446,N_5321,N_5303);
and U5447 (N_5447,N_5350,N_5304);
and U5448 (N_5448,N_5301,N_5398);
nand U5449 (N_5449,N_5302,N_5372);
nand U5450 (N_5450,N_5334,N_5370);
xnor U5451 (N_5451,N_5334,N_5338);
nand U5452 (N_5452,N_5328,N_5313);
nor U5453 (N_5453,N_5316,N_5377);
and U5454 (N_5454,N_5354,N_5399);
or U5455 (N_5455,N_5354,N_5374);
nand U5456 (N_5456,N_5358,N_5365);
nor U5457 (N_5457,N_5397,N_5362);
and U5458 (N_5458,N_5312,N_5387);
and U5459 (N_5459,N_5329,N_5361);
or U5460 (N_5460,N_5362,N_5379);
nor U5461 (N_5461,N_5394,N_5374);
nor U5462 (N_5462,N_5339,N_5383);
or U5463 (N_5463,N_5399,N_5372);
or U5464 (N_5464,N_5313,N_5340);
and U5465 (N_5465,N_5359,N_5361);
and U5466 (N_5466,N_5339,N_5311);
nand U5467 (N_5467,N_5380,N_5361);
nand U5468 (N_5468,N_5312,N_5347);
nand U5469 (N_5469,N_5318,N_5353);
or U5470 (N_5470,N_5308,N_5339);
or U5471 (N_5471,N_5318,N_5389);
nand U5472 (N_5472,N_5335,N_5394);
nand U5473 (N_5473,N_5357,N_5308);
nand U5474 (N_5474,N_5366,N_5332);
nand U5475 (N_5475,N_5364,N_5343);
nand U5476 (N_5476,N_5321,N_5335);
or U5477 (N_5477,N_5335,N_5386);
or U5478 (N_5478,N_5311,N_5309);
and U5479 (N_5479,N_5397,N_5392);
nor U5480 (N_5480,N_5334,N_5398);
or U5481 (N_5481,N_5306,N_5313);
nor U5482 (N_5482,N_5311,N_5330);
nand U5483 (N_5483,N_5386,N_5375);
or U5484 (N_5484,N_5383,N_5388);
and U5485 (N_5485,N_5348,N_5301);
nor U5486 (N_5486,N_5379,N_5397);
or U5487 (N_5487,N_5306,N_5377);
and U5488 (N_5488,N_5304,N_5348);
or U5489 (N_5489,N_5310,N_5398);
and U5490 (N_5490,N_5378,N_5366);
nor U5491 (N_5491,N_5348,N_5349);
or U5492 (N_5492,N_5308,N_5310);
nand U5493 (N_5493,N_5347,N_5309);
xor U5494 (N_5494,N_5314,N_5318);
nand U5495 (N_5495,N_5370,N_5397);
nor U5496 (N_5496,N_5305,N_5368);
and U5497 (N_5497,N_5384,N_5332);
and U5498 (N_5498,N_5326,N_5322);
or U5499 (N_5499,N_5350,N_5375);
nor U5500 (N_5500,N_5443,N_5497);
nor U5501 (N_5501,N_5428,N_5486);
nor U5502 (N_5502,N_5483,N_5467);
nand U5503 (N_5503,N_5456,N_5491);
or U5504 (N_5504,N_5406,N_5429);
nand U5505 (N_5505,N_5457,N_5444);
nor U5506 (N_5506,N_5415,N_5401);
and U5507 (N_5507,N_5427,N_5446);
or U5508 (N_5508,N_5464,N_5481);
nand U5509 (N_5509,N_5437,N_5466);
nand U5510 (N_5510,N_5421,N_5441);
and U5511 (N_5511,N_5422,N_5450);
nor U5512 (N_5512,N_5408,N_5434);
nand U5513 (N_5513,N_5479,N_5471);
nand U5514 (N_5514,N_5420,N_5414);
or U5515 (N_5515,N_5413,N_5468);
nand U5516 (N_5516,N_5431,N_5487);
and U5517 (N_5517,N_5494,N_5485);
nor U5518 (N_5518,N_5489,N_5436);
nor U5519 (N_5519,N_5448,N_5425);
and U5520 (N_5520,N_5475,N_5453);
nand U5521 (N_5521,N_5488,N_5493);
nand U5522 (N_5522,N_5407,N_5411);
or U5523 (N_5523,N_5442,N_5459);
nand U5524 (N_5524,N_5476,N_5465);
and U5525 (N_5525,N_5423,N_5424);
or U5526 (N_5526,N_5462,N_5439);
nor U5527 (N_5527,N_5419,N_5452);
nand U5528 (N_5528,N_5482,N_5430);
or U5529 (N_5529,N_5499,N_5418);
and U5530 (N_5530,N_5417,N_5498);
nor U5531 (N_5531,N_5405,N_5463);
nor U5532 (N_5532,N_5412,N_5404);
nor U5533 (N_5533,N_5496,N_5472);
and U5534 (N_5534,N_5403,N_5473);
or U5535 (N_5535,N_5474,N_5440);
nand U5536 (N_5536,N_5410,N_5402);
nor U5537 (N_5537,N_5460,N_5470);
and U5538 (N_5538,N_5447,N_5469);
and U5539 (N_5539,N_5492,N_5455);
and U5540 (N_5540,N_5458,N_5484);
nor U5541 (N_5541,N_5480,N_5435);
nor U5542 (N_5542,N_5432,N_5454);
nand U5543 (N_5543,N_5433,N_5478);
nor U5544 (N_5544,N_5461,N_5416);
nor U5545 (N_5545,N_5490,N_5449);
and U5546 (N_5546,N_5400,N_5477);
nor U5547 (N_5547,N_5445,N_5495);
or U5548 (N_5548,N_5438,N_5426);
or U5549 (N_5549,N_5451,N_5409);
and U5550 (N_5550,N_5416,N_5409);
and U5551 (N_5551,N_5463,N_5420);
and U5552 (N_5552,N_5491,N_5461);
and U5553 (N_5553,N_5479,N_5493);
nand U5554 (N_5554,N_5497,N_5475);
nand U5555 (N_5555,N_5489,N_5493);
nor U5556 (N_5556,N_5401,N_5471);
or U5557 (N_5557,N_5479,N_5484);
nor U5558 (N_5558,N_5407,N_5455);
nor U5559 (N_5559,N_5439,N_5490);
and U5560 (N_5560,N_5491,N_5499);
or U5561 (N_5561,N_5401,N_5439);
nand U5562 (N_5562,N_5456,N_5477);
and U5563 (N_5563,N_5411,N_5441);
or U5564 (N_5564,N_5454,N_5459);
nor U5565 (N_5565,N_5492,N_5434);
nand U5566 (N_5566,N_5405,N_5478);
and U5567 (N_5567,N_5462,N_5416);
nand U5568 (N_5568,N_5408,N_5482);
and U5569 (N_5569,N_5498,N_5440);
and U5570 (N_5570,N_5400,N_5483);
or U5571 (N_5571,N_5440,N_5450);
nand U5572 (N_5572,N_5435,N_5485);
nand U5573 (N_5573,N_5459,N_5432);
nand U5574 (N_5574,N_5466,N_5496);
nand U5575 (N_5575,N_5470,N_5436);
or U5576 (N_5576,N_5441,N_5468);
or U5577 (N_5577,N_5488,N_5490);
nor U5578 (N_5578,N_5425,N_5473);
and U5579 (N_5579,N_5498,N_5419);
nand U5580 (N_5580,N_5454,N_5423);
nand U5581 (N_5581,N_5403,N_5472);
and U5582 (N_5582,N_5418,N_5484);
and U5583 (N_5583,N_5486,N_5400);
and U5584 (N_5584,N_5461,N_5458);
nand U5585 (N_5585,N_5457,N_5498);
nand U5586 (N_5586,N_5474,N_5475);
and U5587 (N_5587,N_5420,N_5456);
and U5588 (N_5588,N_5414,N_5431);
nor U5589 (N_5589,N_5417,N_5458);
nand U5590 (N_5590,N_5481,N_5475);
nand U5591 (N_5591,N_5470,N_5475);
xnor U5592 (N_5592,N_5421,N_5475);
nor U5593 (N_5593,N_5470,N_5440);
and U5594 (N_5594,N_5494,N_5496);
nand U5595 (N_5595,N_5486,N_5499);
or U5596 (N_5596,N_5447,N_5450);
or U5597 (N_5597,N_5491,N_5486);
or U5598 (N_5598,N_5484,N_5495);
nand U5599 (N_5599,N_5445,N_5417);
nand U5600 (N_5600,N_5563,N_5560);
or U5601 (N_5601,N_5586,N_5549);
nor U5602 (N_5602,N_5515,N_5535);
nor U5603 (N_5603,N_5512,N_5522);
and U5604 (N_5604,N_5546,N_5584);
or U5605 (N_5605,N_5565,N_5556);
nand U5606 (N_5606,N_5521,N_5553);
or U5607 (N_5607,N_5578,N_5593);
nand U5608 (N_5608,N_5577,N_5507);
nand U5609 (N_5609,N_5504,N_5513);
nand U5610 (N_5610,N_5597,N_5518);
nand U5611 (N_5611,N_5508,N_5533);
nor U5612 (N_5612,N_5548,N_5530);
and U5613 (N_5613,N_5592,N_5501);
or U5614 (N_5614,N_5509,N_5526);
nor U5615 (N_5615,N_5527,N_5542);
nand U5616 (N_5616,N_5557,N_5514);
nor U5617 (N_5617,N_5591,N_5540);
nor U5618 (N_5618,N_5579,N_5599);
nor U5619 (N_5619,N_5519,N_5590);
nand U5620 (N_5620,N_5581,N_5529);
and U5621 (N_5621,N_5523,N_5571);
nand U5622 (N_5622,N_5567,N_5511);
or U5623 (N_5623,N_5531,N_5541);
and U5624 (N_5624,N_5532,N_5595);
nand U5625 (N_5625,N_5550,N_5547);
and U5626 (N_5626,N_5502,N_5543);
nand U5627 (N_5627,N_5517,N_5552);
nand U5628 (N_5628,N_5561,N_5524);
and U5629 (N_5629,N_5570,N_5596);
or U5630 (N_5630,N_5516,N_5594);
nor U5631 (N_5631,N_5539,N_5505);
nand U5632 (N_5632,N_5580,N_5525);
nand U5633 (N_5633,N_5534,N_5572);
nand U5634 (N_5634,N_5583,N_5558);
nand U5635 (N_5635,N_5588,N_5503);
and U5636 (N_5636,N_5585,N_5574);
nor U5637 (N_5637,N_5538,N_5564);
or U5638 (N_5638,N_5500,N_5545);
nand U5639 (N_5639,N_5582,N_5569);
nor U5640 (N_5640,N_5559,N_5554);
nand U5641 (N_5641,N_5589,N_5587);
and U5642 (N_5642,N_5536,N_5562);
nor U5643 (N_5643,N_5544,N_5506);
xnor U5644 (N_5644,N_5510,N_5551);
and U5645 (N_5645,N_5537,N_5576);
and U5646 (N_5646,N_5568,N_5575);
or U5647 (N_5647,N_5528,N_5520);
and U5648 (N_5648,N_5555,N_5598);
nand U5649 (N_5649,N_5573,N_5566);
or U5650 (N_5650,N_5554,N_5530);
or U5651 (N_5651,N_5573,N_5506);
and U5652 (N_5652,N_5584,N_5533);
and U5653 (N_5653,N_5519,N_5512);
nor U5654 (N_5654,N_5586,N_5527);
nor U5655 (N_5655,N_5530,N_5531);
and U5656 (N_5656,N_5583,N_5596);
nand U5657 (N_5657,N_5570,N_5516);
nor U5658 (N_5658,N_5581,N_5504);
and U5659 (N_5659,N_5544,N_5504);
or U5660 (N_5660,N_5523,N_5567);
nor U5661 (N_5661,N_5593,N_5566);
or U5662 (N_5662,N_5532,N_5594);
and U5663 (N_5663,N_5500,N_5503);
xor U5664 (N_5664,N_5548,N_5555);
nand U5665 (N_5665,N_5577,N_5501);
nor U5666 (N_5666,N_5549,N_5568);
nand U5667 (N_5667,N_5543,N_5571);
and U5668 (N_5668,N_5584,N_5543);
or U5669 (N_5669,N_5540,N_5576);
or U5670 (N_5670,N_5553,N_5529);
nand U5671 (N_5671,N_5526,N_5598);
or U5672 (N_5672,N_5574,N_5531);
nand U5673 (N_5673,N_5549,N_5585);
and U5674 (N_5674,N_5548,N_5506);
nor U5675 (N_5675,N_5585,N_5586);
and U5676 (N_5676,N_5517,N_5574);
or U5677 (N_5677,N_5563,N_5582);
nor U5678 (N_5678,N_5549,N_5507);
nor U5679 (N_5679,N_5541,N_5540);
and U5680 (N_5680,N_5558,N_5527);
nand U5681 (N_5681,N_5579,N_5562);
nor U5682 (N_5682,N_5541,N_5571);
nand U5683 (N_5683,N_5519,N_5544);
or U5684 (N_5684,N_5575,N_5513);
or U5685 (N_5685,N_5573,N_5561);
nand U5686 (N_5686,N_5567,N_5578);
nand U5687 (N_5687,N_5559,N_5595);
or U5688 (N_5688,N_5571,N_5516);
and U5689 (N_5689,N_5541,N_5567);
or U5690 (N_5690,N_5594,N_5564);
nand U5691 (N_5691,N_5556,N_5525);
nor U5692 (N_5692,N_5593,N_5567);
nand U5693 (N_5693,N_5544,N_5574);
nand U5694 (N_5694,N_5515,N_5559);
and U5695 (N_5695,N_5585,N_5556);
nand U5696 (N_5696,N_5552,N_5511);
nand U5697 (N_5697,N_5568,N_5505);
and U5698 (N_5698,N_5527,N_5534);
and U5699 (N_5699,N_5596,N_5565);
nand U5700 (N_5700,N_5694,N_5679);
nor U5701 (N_5701,N_5650,N_5698);
and U5702 (N_5702,N_5699,N_5622);
or U5703 (N_5703,N_5633,N_5677);
nand U5704 (N_5704,N_5670,N_5682);
nor U5705 (N_5705,N_5610,N_5647);
and U5706 (N_5706,N_5672,N_5632);
and U5707 (N_5707,N_5608,N_5630);
nand U5708 (N_5708,N_5619,N_5638);
or U5709 (N_5709,N_5675,N_5642);
or U5710 (N_5710,N_5613,N_5648);
and U5711 (N_5711,N_5640,N_5602);
or U5712 (N_5712,N_5649,N_5697);
or U5713 (N_5713,N_5646,N_5686);
nand U5714 (N_5714,N_5629,N_5687);
and U5715 (N_5715,N_5681,N_5688);
nand U5716 (N_5716,N_5685,N_5668);
or U5717 (N_5717,N_5643,N_5606);
nand U5718 (N_5718,N_5660,N_5628);
or U5719 (N_5719,N_5653,N_5673);
and U5720 (N_5720,N_5678,N_5695);
nor U5721 (N_5721,N_5639,N_5645);
or U5722 (N_5722,N_5644,N_5626);
nand U5723 (N_5723,N_5661,N_5654);
nor U5724 (N_5724,N_5696,N_5680);
nor U5725 (N_5725,N_5690,N_5669);
nand U5726 (N_5726,N_5612,N_5616);
and U5727 (N_5727,N_5665,N_5667);
or U5728 (N_5728,N_5691,N_5674);
nand U5729 (N_5729,N_5692,N_5621);
and U5730 (N_5730,N_5601,N_5618);
or U5731 (N_5731,N_5655,N_5617);
or U5732 (N_5732,N_5605,N_5614);
or U5733 (N_5733,N_5651,N_5607);
or U5734 (N_5734,N_5689,N_5666);
and U5735 (N_5735,N_5662,N_5664);
and U5736 (N_5736,N_5631,N_5658);
nor U5737 (N_5737,N_5659,N_5637);
or U5738 (N_5738,N_5634,N_5636);
or U5739 (N_5739,N_5641,N_5683);
and U5740 (N_5740,N_5609,N_5671);
and U5741 (N_5741,N_5600,N_5657);
or U5742 (N_5742,N_5615,N_5625);
nor U5743 (N_5743,N_5623,N_5676);
and U5744 (N_5744,N_5635,N_5684);
or U5745 (N_5745,N_5603,N_5624);
and U5746 (N_5746,N_5627,N_5604);
and U5747 (N_5747,N_5693,N_5663);
nor U5748 (N_5748,N_5611,N_5620);
or U5749 (N_5749,N_5652,N_5656);
nand U5750 (N_5750,N_5666,N_5677);
and U5751 (N_5751,N_5677,N_5637);
or U5752 (N_5752,N_5614,N_5663);
and U5753 (N_5753,N_5615,N_5673);
or U5754 (N_5754,N_5655,N_5682);
nor U5755 (N_5755,N_5605,N_5688);
or U5756 (N_5756,N_5610,N_5613);
nor U5757 (N_5757,N_5690,N_5667);
nor U5758 (N_5758,N_5680,N_5645);
nor U5759 (N_5759,N_5627,N_5623);
nor U5760 (N_5760,N_5604,N_5601);
or U5761 (N_5761,N_5672,N_5622);
nand U5762 (N_5762,N_5645,N_5624);
nand U5763 (N_5763,N_5609,N_5618);
or U5764 (N_5764,N_5680,N_5606);
and U5765 (N_5765,N_5663,N_5687);
or U5766 (N_5766,N_5671,N_5626);
and U5767 (N_5767,N_5678,N_5655);
or U5768 (N_5768,N_5635,N_5672);
and U5769 (N_5769,N_5692,N_5636);
or U5770 (N_5770,N_5686,N_5606);
and U5771 (N_5771,N_5656,N_5675);
and U5772 (N_5772,N_5620,N_5679);
nand U5773 (N_5773,N_5648,N_5654);
nor U5774 (N_5774,N_5619,N_5636);
and U5775 (N_5775,N_5685,N_5659);
nor U5776 (N_5776,N_5615,N_5644);
and U5777 (N_5777,N_5686,N_5650);
nor U5778 (N_5778,N_5627,N_5676);
nand U5779 (N_5779,N_5682,N_5626);
nor U5780 (N_5780,N_5640,N_5620);
and U5781 (N_5781,N_5670,N_5620);
or U5782 (N_5782,N_5664,N_5615);
nor U5783 (N_5783,N_5687,N_5640);
or U5784 (N_5784,N_5606,N_5602);
nor U5785 (N_5785,N_5676,N_5610);
and U5786 (N_5786,N_5684,N_5651);
and U5787 (N_5787,N_5694,N_5667);
and U5788 (N_5788,N_5660,N_5634);
or U5789 (N_5789,N_5648,N_5610);
nand U5790 (N_5790,N_5692,N_5677);
nand U5791 (N_5791,N_5641,N_5689);
nor U5792 (N_5792,N_5697,N_5666);
or U5793 (N_5793,N_5624,N_5614);
and U5794 (N_5794,N_5695,N_5617);
nand U5795 (N_5795,N_5632,N_5620);
or U5796 (N_5796,N_5628,N_5636);
or U5797 (N_5797,N_5692,N_5699);
nor U5798 (N_5798,N_5606,N_5610);
and U5799 (N_5799,N_5671,N_5665);
nor U5800 (N_5800,N_5787,N_5778);
or U5801 (N_5801,N_5750,N_5716);
nor U5802 (N_5802,N_5761,N_5772);
and U5803 (N_5803,N_5799,N_5707);
and U5804 (N_5804,N_5700,N_5704);
nand U5805 (N_5805,N_5710,N_5759);
and U5806 (N_5806,N_5781,N_5724);
nand U5807 (N_5807,N_5791,N_5786);
or U5808 (N_5808,N_5784,N_5727);
and U5809 (N_5809,N_5764,N_5729);
nor U5810 (N_5810,N_5755,N_5776);
nand U5811 (N_5811,N_5735,N_5734);
and U5812 (N_5812,N_5726,N_5733);
or U5813 (N_5813,N_5771,N_5797);
nor U5814 (N_5814,N_5752,N_5708);
nor U5815 (N_5815,N_5779,N_5768);
and U5816 (N_5816,N_5722,N_5789);
nand U5817 (N_5817,N_5715,N_5739);
or U5818 (N_5818,N_5774,N_5712);
and U5819 (N_5819,N_5703,N_5717);
nand U5820 (N_5820,N_5743,N_5706);
nand U5821 (N_5821,N_5762,N_5782);
nor U5822 (N_5822,N_5795,N_5731);
or U5823 (N_5823,N_5758,N_5780);
and U5824 (N_5824,N_5792,N_5713);
and U5825 (N_5825,N_5738,N_5736);
or U5826 (N_5826,N_5741,N_5767);
nand U5827 (N_5827,N_5760,N_5766);
or U5828 (N_5828,N_5796,N_5777);
or U5829 (N_5829,N_5785,N_5740);
nand U5830 (N_5830,N_5751,N_5709);
and U5831 (N_5831,N_5745,N_5702);
and U5832 (N_5832,N_5746,N_5793);
or U5833 (N_5833,N_5794,N_5773);
or U5834 (N_5834,N_5747,N_5757);
nor U5835 (N_5835,N_5719,N_5749);
nor U5836 (N_5836,N_5775,N_5705);
nand U5837 (N_5837,N_5720,N_5756);
or U5838 (N_5838,N_5737,N_5783);
nand U5839 (N_5839,N_5732,N_5754);
or U5840 (N_5840,N_5765,N_5711);
or U5841 (N_5841,N_5728,N_5714);
or U5842 (N_5842,N_5742,N_5769);
or U5843 (N_5843,N_5730,N_5718);
or U5844 (N_5844,N_5763,N_5798);
nor U5845 (N_5845,N_5721,N_5788);
nand U5846 (N_5846,N_5748,N_5770);
or U5847 (N_5847,N_5790,N_5723);
nor U5848 (N_5848,N_5725,N_5744);
nand U5849 (N_5849,N_5753,N_5701);
nand U5850 (N_5850,N_5788,N_5715);
nand U5851 (N_5851,N_5761,N_5742);
nor U5852 (N_5852,N_5759,N_5751);
nor U5853 (N_5853,N_5719,N_5722);
nor U5854 (N_5854,N_5724,N_5789);
and U5855 (N_5855,N_5700,N_5748);
nand U5856 (N_5856,N_5709,N_5758);
nor U5857 (N_5857,N_5762,N_5774);
nor U5858 (N_5858,N_5751,N_5788);
or U5859 (N_5859,N_5733,N_5760);
and U5860 (N_5860,N_5791,N_5729);
and U5861 (N_5861,N_5772,N_5754);
nor U5862 (N_5862,N_5709,N_5738);
nand U5863 (N_5863,N_5721,N_5716);
and U5864 (N_5864,N_5716,N_5724);
and U5865 (N_5865,N_5776,N_5726);
or U5866 (N_5866,N_5761,N_5717);
nor U5867 (N_5867,N_5723,N_5711);
nand U5868 (N_5868,N_5703,N_5797);
or U5869 (N_5869,N_5745,N_5741);
or U5870 (N_5870,N_5798,N_5702);
and U5871 (N_5871,N_5780,N_5716);
or U5872 (N_5872,N_5773,N_5754);
or U5873 (N_5873,N_5736,N_5710);
nor U5874 (N_5874,N_5762,N_5768);
nor U5875 (N_5875,N_5789,N_5726);
nor U5876 (N_5876,N_5748,N_5783);
and U5877 (N_5877,N_5700,N_5756);
or U5878 (N_5878,N_5752,N_5770);
nor U5879 (N_5879,N_5710,N_5781);
nand U5880 (N_5880,N_5780,N_5776);
or U5881 (N_5881,N_5763,N_5764);
nand U5882 (N_5882,N_5726,N_5734);
and U5883 (N_5883,N_5764,N_5756);
nand U5884 (N_5884,N_5709,N_5774);
nor U5885 (N_5885,N_5725,N_5739);
and U5886 (N_5886,N_5758,N_5701);
or U5887 (N_5887,N_5752,N_5767);
or U5888 (N_5888,N_5718,N_5793);
or U5889 (N_5889,N_5747,N_5731);
nand U5890 (N_5890,N_5798,N_5716);
and U5891 (N_5891,N_5772,N_5703);
and U5892 (N_5892,N_5780,N_5767);
nor U5893 (N_5893,N_5777,N_5709);
nand U5894 (N_5894,N_5727,N_5746);
or U5895 (N_5895,N_5791,N_5751);
nand U5896 (N_5896,N_5754,N_5705);
nor U5897 (N_5897,N_5765,N_5705);
nand U5898 (N_5898,N_5719,N_5795);
or U5899 (N_5899,N_5784,N_5785);
and U5900 (N_5900,N_5879,N_5841);
nor U5901 (N_5901,N_5877,N_5881);
or U5902 (N_5902,N_5855,N_5829);
and U5903 (N_5903,N_5826,N_5810);
nand U5904 (N_5904,N_5883,N_5822);
nor U5905 (N_5905,N_5885,N_5825);
or U5906 (N_5906,N_5876,N_5840);
nor U5907 (N_5907,N_5849,N_5846);
nor U5908 (N_5908,N_5897,N_5802);
nor U5909 (N_5909,N_5856,N_5867);
nor U5910 (N_5910,N_5860,N_5821);
or U5911 (N_5911,N_5870,N_5820);
and U5912 (N_5912,N_5853,N_5854);
and U5913 (N_5913,N_5865,N_5816);
or U5914 (N_5914,N_5812,N_5839);
nor U5915 (N_5915,N_5868,N_5845);
nand U5916 (N_5916,N_5836,N_5838);
nor U5917 (N_5917,N_5880,N_5857);
nand U5918 (N_5918,N_5890,N_5891);
or U5919 (N_5919,N_5837,N_5887);
and U5920 (N_5920,N_5817,N_5896);
nand U5921 (N_5921,N_5842,N_5863);
nor U5922 (N_5922,N_5894,N_5882);
nand U5923 (N_5923,N_5828,N_5801);
nand U5924 (N_5924,N_5831,N_5844);
nand U5925 (N_5925,N_5811,N_5818);
or U5926 (N_5926,N_5851,N_5804);
or U5927 (N_5927,N_5886,N_5835);
nor U5928 (N_5928,N_5871,N_5852);
nor U5929 (N_5929,N_5808,N_5830);
or U5930 (N_5930,N_5819,N_5843);
nand U5931 (N_5931,N_5872,N_5809);
nand U5932 (N_5932,N_5814,N_5895);
and U5933 (N_5933,N_5833,N_5834);
or U5934 (N_5934,N_5866,N_5858);
and U5935 (N_5935,N_5878,N_5888);
and U5936 (N_5936,N_5893,N_5800);
nor U5937 (N_5937,N_5862,N_5806);
nor U5938 (N_5938,N_5864,N_5873);
nor U5939 (N_5939,N_5832,N_5892);
nor U5940 (N_5940,N_5847,N_5859);
nor U5941 (N_5941,N_5827,N_5898);
nor U5942 (N_5942,N_5884,N_5869);
nand U5943 (N_5943,N_5813,N_5823);
nor U5944 (N_5944,N_5805,N_5874);
and U5945 (N_5945,N_5803,N_5899);
or U5946 (N_5946,N_5848,N_5824);
nand U5947 (N_5947,N_5807,N_5815);
nand U5948 (N_5948,N_5889,N_5861);
or U5949 (N_5949,N_5850,N_5875);
nor U5950 (N_5950,N_5888,N_5858);
or U5951 (N_5951,N_5838,N_5831);
nand U5952 (N_5952,N_5869,N_5806);
nor U5953 (N_5953,N_5891,N_5819);
and U5954 (N_5954,N_5893,N_5805);
and U5955 (N_5955,N_5824,N_5853);
nand U5956 (N_5956,N_5826,N_5862);
nor U5957 (N_5957,N_5835,N_5852);
or U5958 (N_5958,N_5832,N_5836);
nor U5959 (N_5959,N_5860,N_5831);
nor U5960 (N_5960,N_5834,N_5885);
or U5961 (N_5961,N_5889,N_5875);
or U5962 (N_5962,N_5876,N_5886);
nor U5963 (N_5963,N_5816,N_5843);
xor U5964 (N_5964,N_5843,N_5858);
and U5965 (N_5965,N_5845,N_5872);
nand U5966 (N_5966,N_5812,N_5886);
and U5967 (N_5967,N_5866,N_5800);
and U5968 (N_5968,N_5858,N_5839);
nor U5969 (N_5969,N_5838,N_5808);
or U5970 (N_5970,N_5845,N_5867);
nor U5971 (N_5971,N_5849,N_5853);
nand U5972 (N_5972,N_5878,N_5885);
nand U5973 (N_5973,N_5854,N_5892);
and U5974 (N_5974,N_5870,N_5875);
nor U5975 (N_5975,N_5854,N_5890);
nor U5976 (N_5976,N_5810,N_5832);
nor U5977 (N_5977,N_5837,N_5882);
nand U5978 (N_5978,N_5888,N_5874);
or U5979 (N_5979,N_5887,N_5883);
or U5980 (N_5980,N_5860,N_5805);
nor U5981 (N_5981,N_5812,N_5803);
and U5982 (N_5982,N_5894,N_5876);
nor U5983 (N_5983,N_5860,N_5812);
and U5984 (N_5984,N_5853,N_5828);
nand U5985 (N_5985,N_5885,N_5827);
or U5986 (N_5986,N_5827,N_5871);
nor U5987 (N_5987,N_5825,N_5844);
nor U5988 (N_5988,N_5801,N_5816);
or U5989 (N_5989,N_5853,N_5818);
or U5990 (N_5990,N_5875,N_5891);
and U5991 (N_5991,N_5898,N_5835);
or U5992 (N_5992,N_5858,N_5832);
nand U5993 (N_5993,N_5867,N_5826);
nor U5994 (N_5994,N_5886,N_5881);
and U5995 (N_5995,N_5803,N_5881);
nor U5996 (N_5996,N_5869,N_5834);
and U5997 (N_5997,N_5827,N_5819);
nor U5998 (N_5998,N_5844,N_5864);
or U5999 (N_5999,N_5857,N_5827);
and U6000 (N_6000,N_5965,N_5998);
or U6001 (N_6001,N_5984,N_5944);
or U6002 (N_6002,N_5981,N_5949);
nor U6003 (N_6003,N_5992,N_5921);
and U6004 (N_6004,N_5990,N_5976);
nand U6005 (N_6005,N_5956,N_5963);
nor U6006 (N_6006,N_5945,N_5940);
nand U6007 (N_6007,N_5957,N_5985);
or U6008 (N_6008,N_5910,N_5915);
and U6009 (N_6009,N_5930,N_5916);
and U6010 (N_6010,N_5982,N_5914);
and U6011 (N_6011,N_5959,N_5901);
nor U6012 (N_6012,N_5929,N_5954);
nand U6013 (N_6013,N_5922,N_5967);
and U6014 (N_6014,N_5909,N_5947);
nand U6015 (N_6015,N_5932,N_5958);
nor U6016 (N_6016,N_5993,N_5908);
and U6017 (N_6017,N_5988,N_5994);
nor U6018 (N_6018,N_5934,N_5964);
and U6019 (N_6019,N_5996,N_5975);
or U6020 (N_6020,N_5923,N_5971);
and U6021 (N_6021,N_5997,N_5969);
nor U6022 (N_6022,N_5973,N_5902);
or U6023 (N_6023,N_5977,N_5920);
and U6024 (N_6024,N_5938,N_5995);
nand U6025 (N_6025,N_5952,N_5962);
or U6026 (N_6026,N_5904,N_5970);
nand U6027 (N_6027,N_5999,N_5935);
nor U6028 (N_6028,N_5926,N_5925);
nor U6029 (N_6029,N_5978,N_5939);
and U6030 (N_6030,N_5905,N_5961);
or U6031 (N_6031,N_5943,N_5900);
nor U6032 (N_6032,N_5960,N_5991);
and U6033 (N_6033,N_5924,N_5968);
nand U6034 (N_6034,N_5917,N_5912);
or U6035 (N_6035,N_5937,N_5931);
and U6036 (N_6036,N_5955,N_5946);
nor U6037 (N_6037,N_5918,N_5986);
or U6038 (N_6038,N_5987,N_5941);
nand U6039 (N_6039,N_5974,N_5948);
or U6040 (N_6040,N_5919,N_5979);
and U6041 (N_6041,N_5972,N_5911);
or U6042 (N_6042,N_5953,N_5983);
and U6043 (N_6043,N_5951,N_5933);
or U6044 (N_6044,N_5942,N_5936);
nand U6045 (N_6045,N_5980,N_5927);
and U6046 (N_6046,N_5989,N_5950);
or U6047 (N_6047,N_5903,N_5906);
nand U6048 (N_6048,N_5966,N_5907);
nand U6049 (N_6049,N_5913,N_5928);
or U6050 (N_6050,N_5963,N_5998);
and U6051 (N_6051,N_5987,N_5919);
and U6052 (N_6052,N_5982,N_5984);
and U6053 (N_6053,N_5929,N_5902);
and U6054 (N_6054,N_5936,N_5958);
or U6055 (N_6055,N_5914,N_5962);
and U6056 (N_6056,N_5966,N_5939);
and U6057 (N_6057,N_5971,N_5970);
and U6058 (N_6058,N_5963,N_5993);
and U6059 (N_6059,N_5909,N_5908);
or U6060 (N_6060,N_5919,N_5928);
nor U6061 (N_6061,N_5914,N_5946);
nand U6062 (N_6062,N_5901,N_5951);
nor U6063 (N_6063,N_5976,N_5930);
or U6064 (N_6064,N_5931,N_5964);
and U6065 (N_6065,N_5990,N_5927);
or U6066 (N_6066,N_5973,N_5943);
nor U6067 (N_6067,N_5923,N_5901);
or U6068 (N_6068,N_5922,N_5963);
nand U6069 (N_6069,N_5942,N_5900);
or U6070 (N_6070,N_5998,N_5918);
nand U6071 (N_6071,N_5933,N_5932);
nor U6072 (N_6072,N_5903,N_5919);
nor U6073 (N_6073,N_5917,N_5927);
or U6074 (N_6074,N_5934,N_5902);
xnor U6075 (N_6075,N_5975,N_5970);
nand U6076 (N_6076,N_5916,N_5962);
and U6077 (N_6077,N_5996,N_5998);
nor U6078 (N_6078,N_5936,N_5929);
or U6079 (N_6079,N_5968,N_5997);
and U6080 (N_6080,N_5946,N_5947);
and U6081 (N_6081,N_5993,N_5943);
or U6082 (N_6082,N_5950,N_5924);
or U6083 (N_6083,N_5989,N_5973);
nor U6084 (N_6084,N_5980,N_5992);
nor U6085 (N_6085,N_5925,N_5975);
and U6086 (N_6086,N_5954,N_5976);
nor U6087 (N_6087,N_5933,N_5948);
nand U6088 (N_6088,N_5984,N_5923);
nand U6089 (N_6089,N_5931,N_5922);
or U6090 (N_6090,N_5998,N_5942);
nor U6091 (N_6091,N_5946,N_5939);
nor U6092 (N_6092,N_5918,N_5980);
and U6093 (N_6093,N_5959,N_5986);
and U6094 (N_6094,N_5904,N_5901);
nand U6095 (N_6095,N_5985,N_5992);
or U6096 (N_6096,N_5957,N_5916);
or U6097 (N_6097,N_5987,N_5985);
and U6098 (N_6098,N_5901,N_5999);
nand U6099 (N_6099,N_5922,N_5995);
and U6100 (N_6100,N_6043,N_6090);
nand U6101 (N_6101,N_6033,N_6096);
nand U6102 (N_6102,N_6029,N_6038);
nand U6103 (N_6103,N_6070,N_6042);
nor U6104 (N_6104,N_6046,N_6075);
nor U6105 (N_6105,N_6079,N_6063);
nor U6106 (N_6106,N_6002,N_6094);
and U6107 (N_6107,N_6084,N_6028);
nand U6108 (N_6108,N_6056,N_6013);
nor U6109 (N_6109,N_6053,N_6019);
nand U6110 (N_6110,N_6060,N_6024);
and U6111 (N_6111,N_6091,N_6098);
and U6112 (N_6112,N_6011,N_6010);
nor U6113 (N_6113,N_6040,N_6045);
or U6114 (N_6114,N_6021,N_6064);
and U6115 (N_6115,N_6080,N_6081);
and U6116 (N_6116,N_6037,N_6059);
and U6117 (N_6117,N_6077,N_6027);
nor U6118 (N_6118,N_6018,N_6052);
or U6119 (N_6119,N_6032,N_6001);
nand U6120 (N_6120,N_6066,N_6082);
and U6121 (N_6121,N_6044,N_6007);
and U6122 (N_6122,N_6099,N_6062);
nor U6123 (N_6123,N_6097,N_6031);
or U6124 (N_6124,N_6008,N_6069);
nand U6125 (N_6125,N_6078,N_6017);
or U6126 (N_6126,N_6023,N_6073);
xor U6127 (N_6127,N_6014,N_6047);
or U6128 (N_6128,N_6039,N_6005);
nand U6129 (N_6129,N_6095,N_6036);
and U6130 (N_6130,N_6026,N_6050);
or U6131 (N_6131,N_6076,N_6074);
and U6132 (N_6132,N_6089,N_6068);
nand U6133 (N_6133,N_6049,N_6016);
nand U6134 (N_6134,N_6025,N_6012);
and U6135 (N_6135,N_6088,N_6003);
xor U6136 (N_6136,N_6004,N_6015);
nor U6137 (N_6137,N_6054,N_6065);
or U6138 (N_6138,N_6055,N_6034);
nand U6139 (N_6139,N_6020,N_6057);
or U6140 (N_6140,N_6006,N_6072);
and U6141 (N_6141,N_6071,N_6087);
and U6142 (N_6142,N_6000,N_6061);
nand U6143 (N_6143,N_6048,N_6041);
or U6144 (N_6144,N_6093,N_6092);
nor U6145 (N_6145,N_6030,N_6035);
and U6146 (N_6146,N_6051,N_6067);
nand U6147 (N_6147,N_6022,N_6086);
nand U6148 (N_6148,N_6085,N_6083);
nor U6149 (N_6149,N_6009,N_6058);
nand U6150 (N_6150,N_6079,N_6028);
or U6151 (N_6151,N_6015,N_6065);
nor U6152 (N_6152,N_6070,N_6044);
nor U6153 (N_6153,N_6089,N_6014);
and U6154 (N_6154,N_6047,N_6097);
nand U6155 (N_6155,N_6085,N_6000);
nand U6156 (N_6156,N_6090,N_6095);
or U6157 (N_6157,N_6041,N_6071);
or U6158 (N_6158,N_6014,N_6077);
nor U6159 (N_6159,N_6011,N_6018);
nor U6160 (N_6160,N_6014,N_6023);
and U6161 (N_6161,N_6062,N_6011);
and U6162 (N_6162,N_6022,N_6054);
nor U6163 (N_6163,N_6017,N_6073);
and U6164 (N_6164,N_6041,N_6035);
nand U6165 (N_6165,N_6067,N_6004);
and U6166 (N_6166,N_6001,N_6096);
or U6167 (N_6167,N_6003,N_6043);
or U6168 (N_6168,N_6085,N_6033);
nor U6169 (N_6169,N_6096,N_6018);
nor U6170 (N_6170,N_6065,N_6013);
or U6171 (N_6171,N_6092,N_6008);
nand U6172 (N_6172,N_6013,N_6068);
nand U6173 (N_6173,N_6003,N_6059);
and U6174 (N_6174,N_6076,N_6042);
nor U6175 (N_6175,N_6072,N_6065);
and U6176 (N_6176,N_6021,N_6074);
or U6177 (N_6177,N_6029,N_6033);
nor U6178 (N_6178,N_6027,N_6024);
nor U6179 (N_6179,N_6045,N_6037);
nand U6180 (N_6180,N_6075,N_6074);
and U6181 (N_6181,N_6071,N_6092);
nand U6182 (N_6182,N_6030,N_6023);
or U6183 (N_6183,N_6010,N_6001);
and U6184 (N_6184,N_6055,N_6048);
and U6185 (N_6185,N_6094,N_6052);
nor U6186 (N_6186,N_6045,N_6036);
nor U6187 (N_6187,N_6074,N_6001);
or U6188 (N_6188,N_6023,N_6097);
xor U6189 (N_6189,N_6035,N_6071);
or U6190 (N_6190,N_6067,N_6056);
nand U6191 (N_6191,N_6065,N_6060);
or U6192 (N_6192,N_6005,N_6078);
nor U6193 (N_6193,N_6076,N_6070);
and U6194 (N_6194,N_6018,N_6066);
nand U6195 (N_6195,N_6095,N_6021);
or U6196 (N_6196,N_6021,N_6056);
or U6197 (N_6197,N_6013,N_6095);
nand U6198 (N_6198,N_6093,N_6018);
nand U6199 (N_6199,N_6011,N_6063);
nand U6200 (N_6200,N_6191,N_6177);
nor U6201 (N_6201,N_6132,N_6138);
nand U6202 (N_6202,N_6110,N_6149);
and U6203 (N_6203,N_6183,N_6126);
or U6204 (N_6204,N_6100,N_6170);
or U6205 (N_6205,N_6134,N_6130);
nand U6206 (N_6206,N_6199,N_6162);
xor U6207 (N_6207,N_6153,N_6168);
nand U6208 (N_6208,N_6197,N_6135);
or U6209 (N_6209,N_6169,N_6158);
nand U6210 (N_6210,N_6127,N_6163);
or U6211 (N_6211,N_6125,N_6151);
or U6212 (N_6212,N_6154,N_6184);
nor U6213 (N_6213,N_6144,N_6150);
nor U6214 (N_6214,N_6147,N_6120);
nor U6215 (N_6215,N_6196,N_6121);
and U6216 (N_6216,N_6142,N_6175);
and U6217 (N_6217,N_6189,N_6145);
nand U6218 (N_6218,N_6166,N_6123);
and U6219 (N_6219,N_6114,N_6124);
or U6220 (N_6220,N_6140,N_6108);
and U6221 (N_6221,N_6185,N_6139);
and U6222 (N_6222,N_6186,N_6180);
nand U6223 (N_6223,N_6137,N_6146);
nand U6224 (N_6224,N_6174,N_6172);
nand U6225 (N_6225,N_6133,N_6187);
nand U6226 (N_6226,N_6103,N_6102);
or U6227 (N_6227,N_6198,N_6176);
and U6228 (N_6228,N_6107,N_6141);
and U6229 (N_6229,N_6115,N_6122);
and U6230 (N_6230,N_6109,N_6160);
and U6231 (N_6231,N_6171,N_6101);
or U6232 (N_6232,N_6112,N_6113);
or U6233 (N_6233,N_6159,N_6136);
nand U6234 (N_6234,N_6190,N_6111);
or U6235 (N_6235,N_6116,N_6119);
nor U6236 (N_6236,N_6192,N_6156);
nor U6237 (N_6237,N_6161,N_6104);
or U6238 (N_6238,N_6167,N_6182);
nor U6239 (N_6239,N_6157,N_6155);
nand U6240 (N_6240,N_6188,N_6164);
nor U6241 (N_6241,N_6194,N_6105);
nor U6242 (N_6242,N_6117,N_6193);
and U6243 (N_6243,N_6143,N_6181);
and U6244 (N_6244,N_6129,N_6195);
nor U6245 (N_6245,N_6152,N_6118);
and U6246 (N_6246,N_6173,N_6179);
or U6247 (N_6247,N_6106,N_6128);
or U6248 (N_6248,N_6131,N_6165);
or U6249 (N_6249,N_6148,N_6178);
nand U6250 (N_6250,N_6150,N_6142);
and U6251 (N_6251,N_6181,N_6133);
nand U6252 (N_6252,N_6126,N_6184);
and U6253 (N_6253,N_6198,N_6139);
xor U6254 (N_6254,N_6161,N_6162);
nor U6255 (N_6255,N_6187,N_6154);
or U6256 (N_6256,N_6112,N_6137);
and U6257 (N_6257,N_6100,N_6124);
nor U6258 (N_6258,N_6152,N_6135);
nand U6259 (N_6259,N_6183,N_6110);
nand U6260 (N_6260,N_6114,N_6111);
nor U6261 (N_6261,N_6123,N_6185);
or U6262 (N_6262,N_6170,N_6138);
or U6263 (N_6263,N_6116,N_6167);
nor U6264 (N_6264,N_6195,N_6161);
and U6265 (N_6265,N_6182,N_6144);
nor U6266 (N_6266,N_6172,N_6154);
nand U6267 (N_6267,N_6124,N_6183);
nand U6268 (N_6268,N_6160,N_6135);
and U6269 (N_6269,N_6189,N_6177);
nor U6270 (N_6270,N_6158,N_6168);
nor U6271 (N_6271,N_6107,N_6134);
or U6272 (N_6272,N_6143,N_6138);
or U6273 (N_6273,N_6125,N_6133);
and U6274 (N_6274,N_6132,N_6104);
nand U6275 (N_6275,N_6103,N_6144);
nor U6276 (N_6276,N_6172,N_6101);
nand U6277 (N_6277,N_6122,N_6183);
or U6278 (N_6278,N_6117,N_6144);
nand U6279 (N_6279,N_6107,N_6174);
or U6280 (N_6280,N_6170,N_6169);
or U6281 (N_6281,N_6186,N_6136);
and U6282 (N_6282,N_6121,N_6138);
or U6283 (N_6283,N_6164,N_6167);
and U6284 (N_6284,N_6150,N_6133);
nor U6285 (N_6285,N_6131,N_6105);
nor U6286 (N_6286,N_6174,N_6133);
or U6287 (N_6287,N_6107,N_6166);
or U6288 (N_6288,N_6138,N_6169);
and U6289 (N_6289,N_6183,N_6114);
nor U6290 (N_6290,N_6134,N_6194);
or U6291 (N_6291,N_6131,N_6185);
and U6292 (N_6292,N_6161,N_6194);
nor U6293 (N_6293,N_6178,N_6132);
and U6294 (N_6294,N_6170,N_6120);
nand U6295 (N_6295,N_6139,N_6173);
nor U6296 (N_6296,N_6111,N_6112);
nor U6297 (N_6297,N_6166,N_6121);
and U6298 (N_6298,N_6109,N_6142);
and U6299 (N_6299,N_6165,N_6129);
nand U6300 (N_6300,N_6243,N_6215);
nand U6301 (N_6301,N_6294,N_6207);
and U6302 (N_6302,N_6240,N_6217);
or U6303 (N_6303,N_6253,N_6283);
and U6304 (N_6304,N_6291,N_6261);
nor U6305 (N_6305,N_6264,N_6234);
or U6306 (N_6306,N_6259,N_6216);
and U6307 (N_6307,N_6200,N_6286);
nand U6308 (N_6308,N_6206,N_6227);
nand U6309 (N_6309,N_6296,N_6235);
or U6310 (N_6310,N_6201,N_6208);
xnor U6311 (N_6311,N_6226,N_6238);
and U6312 (N_6312,N_6298,N_6265);
nor U6313 (N_6313,N_6248,N_6275);
and U6314 (N_6314,N_6221,N_6269);
and U6315 (N_6315,N_6239,N_6287);
nand U6316 (N_6316,N_6297,N_6276);
nor U6317 (N_6317,N_6255,N_6203);
and U6318 (N_6318,N_6236,N_6233);
nand U6319 (N_6319,N_6272,N_6256);
or U6320 (N_6320,N_6252,N_6254);
nor U6321 (N_6321,N_6222,N_6277);
nor U6322 (N_6322,N_6263,N_6281);
and U6323 (N_6323,N_6258,N_6224);
and U6324 (N_6324,N_6246,N_6229);
nor U6325 (N_6325,N_6266,N_6295);
and U6326 (N_6326,N_6232,N_6242);
nand U6327 (N_6327,N_6225,N_6213);
nor U6328 (N_6328,N_6202,N_6218);
nor U6329 (N_6329,N_6204,N_6279);
and U6330 (N_6330,N_6267,N_6249);
nor U6331 (N_6331,N_6274,N_6260);
nand U6332 (N_6332,N_6299,N_6223);
or U6333 (N_6333,N_6257,N_6205);
and U6334 (N_6334,N_6211,N_6241);
or U6335 (N_6335,N_6270,N_6220);
nor U6336 (N_6336,N_6214,N_6282);
nand U6337 (N_6337,N_6244,N_6273);
or U6338 (N_6338,N_6228,N_6292);
nand U6339 (N_6339,N_6247,N_6288);
or U6340 (N_6340,N_6230,N_6268);
nor U6341 (N_6341,N_6293,N_6209);
and U6342 (N_6342,N_6262,N_6285);
or U6343 (N_6343,N_6245,N_6290);
and U6344 (N_6344,N_6210,N_6284);
nand U6345 (N_6345,N_6231,N_6278);
or U6346 (N_6346,N_6280,N_6212);
nor U6347 (N_6347,N_6251,N_6289);
and U6348 (N_6348,N_6250,N_6219);
nand U6349 (N_6349,N_6237,N_6271);
or U6350 (N_6350,N_6277,N_6233);
or U6351 (N_6351,N_6211,N_6295);
nand U6352 (N_6352,N_6206,N_6280);
nor U6353 (N_6353,N_6263,N_6283);
nor U6354 (N_6354,N_6296,N_6217);
nor U6355 (N_6355,N_6211,N_6279);
nor U6356 (N_6356,N_6229,N_6230);
nor U6357 (N_6357,N_6250,N_6287);
and U6358 (N_6358,N_6296,N_6268);
nand U6359 (N_6359,N_6254,N_6210);
nor U6360 (N_6360,N_6229,N_6254);
or U6361 (N_6361,N_6255,N_6220);
nor U6362 (N_6362,N_6262,N_6219);
or U6363 (N_6363,N_6239,N_6260);
nand U6364 (N_6364,N_6214,N_6287);
and U6365 (N_6365,N_6299,N_6206);
and U6366 (N_6366,N_6263,N_6276);
nor U6367 (N_6367,N_6231,N_6261);
and U6368 (N_6368,N_6253,N_6297);
nor U6369 (N_6369,N_6271,N_6207);
nor U6370 (N_6370,N_6265,N_6208);
nand U6371 (N_6371,N_6262,N_6283);
nand U6372 (N_6372,N_6290,N_6221);
nor U6373 (N_6373,N_6265,N_6296);
nand U6374 (N_6374,N_6281,N_6292);
and U6375 (N_6375,N_6224,N_6252);
and U6376 (N_6376,N_6202,N_6280);
nand U6377 (N_6377,N_6246,N_6270);
and U6378 (N_6378,N_6276,N_6288);
or U6379 (N_6379,N_6279,N_6288);
nand U6380 (N_6380,N_6271,N_6201);
or U6381 (N_6381,N_6282,N_6266);
nor U6382 (N_6382,N_6243,N_6209);
nor U6383 (N_6383,N_6205,N_6221);
and U6384 (N_6384,N_6237,N_6286);
and U6385 (N_6385,N_6236,N_6221);
or U6386 (N_6386,N_6287,N_6252);
nor U6387 (N_6387,N_6256,N_6289);
nor U6388 (N_6388,N_6253,N_6243);
or U6389 (N_6389,N_6289,N_6238);
nand U6390 (N_6390,N_6221,N_6242);
nor U6391 (N_6391,N_6277,N_6265);
or U6392 (N_6392,N_6291,N_6221);
and U6393 (N_6393,N_6274,N_6216);
nor U6394 (N_6394,N_6284,N_6285);
or U6395 (N_6395,N_6279,N_6242);
nor U6396 (N_6396,N_6252,N_6283);
nand U6397 (N_6397,N_6200,N_6232);
nor U6398 (N_6398,N_6209,N_6236);
nand U6399 (N_6399,N_6290,N_6223);
and U6400 (N_6400,N_6354,N_6315);
nor U6401 (N_6401,N_6399,N_6327);
nand U6402 (N_6402,N_6322,N_6324);
nand U6403 (N_6403,N_6300,N_6370);
and U6404 (N_6404,N_6387,N_6371);
nor U6405 (N_6405,N_6325,N_6314);
and U6406 (N_6406,N_6332,N_6383);
or U6407 (N_6407,N_6356,N_6363);
or U6408 (N_6408,N_6360,N_6318);
nand U6409 (N_6409,N_6373,N_6397);
and U6410 (N_6410,N_6312,N_6331);
and U6411 (N_6411,N_6358,N_6301);
and U6412 (N_6412,N_6342,N_6391);
nor U6413 (N_6413,N_6348,N_6398);
nand U6414 (N_6414,N_6393,N_6390);
nand U6415 (N_6415,N_6323,N_6344);
nor U6416 (N_6416,N_6345,N_6346);
nor U6417 (N_6417,N_6352,N_6364);
nand U6418 (N_6418,N_6376,N_6326);
nand U6419 (N_6419,N_6377,N_6336);
nor U6420 (N_6420,N_6389,N_6333);
nor U6421 (N_6421,N_6350,N_6334);
nor U6422 (N_6422,N_6355,N_6379);
nor U6423 (N_6423,N_6362,N_6310);
or U6424 (N_6424,N_6367,N_6349);
and U6425 (N_6425,N_6319,N_6388);
or U6426 (N_6426,N_6321,N_6316);
or U6427 (N_6427,N_6307,N_6382);
nand U6428 (N_6428,N_6384,N_6396);
or U6429 (N_6429,N_6392,N_6353);
or U6430 (N_6430,N_6385,N_6306);
and U6431 (N_6431,N_6308,N_6340);
and U6432 (N_6432,N_6304,N_6338);
and U6433 (N_6433,N_6328,N_6378);
nor U6434 (N_6434,N_6351,N_6317);
nor U6435 (N_6435,N_6330,N_6372);
or U6436 (N_6436,N_6386,N_6369);
and U6437 (N_6437,N_6357,N_6361);
nor U6438 (N_6438,N_6311,N_6305);
and U6439 (N_6439,N_6380,N_6337);
nand U6440 (N_6440,N_6302,N_6375);
nand U6441 (N_6441,N_6343,N_6339);
nand U6442 (N_6442,N_6359,N_6347);
or U6443 (N_6443,N_6303,N_6320);
xnor U6444 (N_6444,N_6395,N_6309);
nand U6445 (N_6445,N_6368,N_6335);
and U6446 (N_6446,N_6365,N_6394);
nor U6447 (N_6447,N_6313,N_6381);
nand U6448 (N_6448,N_6366,N_6374);
and U6449 (N_6449,N_6329,N_6341);
and U6450 (N_6450,N_6365,N_6388);
nand U6451 (N_6451,N_6349,N_6306);
nand U6452 (N_6452,N_6373,N_6356);
nor U6453 (N_6453,N_6318,N_6327);
or U6454 (N_6454,N_6373,N_6323);
or U6455 (N_6455,N_6312,N_6303);
nand U6456 (N_6456,N_6384,N_6379);
or U6457 (N_6457,N_6309,N_6386);
nand U6458 (N_6458,N_6355,N_6398);
nor U6459 (N_6459,N_6316,N_6397);
nor U6460 (N_6460,N_6387,N_6388);
or U6461 (N_6461,N_6337,N_6333);
or U6462 (N_6462,N_6325,N_6365);
nor U6463 (N_6463,N_6306,N_6393);
nor U6464 (N_6464,N_6311,N_6398);
nand U6465 (N_6465,N_6337,N_6326);
and U6466 (N_6466,N_6345,N_6325);
or U6467 (N_6467,N_6306,N_6344);
nor U6468 (N_6468,N_6339,N_6395);
nand U6469 (N_6469,N_6320,N_6313);
and U6470 (N_6470,N_6394,N_6306);
nand U6471 (N_6471,N_6377,N_6341);
nor U6472 (N_6472,N_6320,N_6329);
and U6473 (N_6473,N_6319,N_6365);
or U6474 (N_6474,N_6392,N_6329);
or U6475 (N_6475,N_6362,N_6383);
and U6476 (N_6476,N_6378,N_6324);
nand U6477 (N_6477,N_6354,N_6355);
and U6478 (N_6478,N_6350,N_6338);
xor U6479 (N_6479,N_6317,N_6330);
and U6480 (N_6480,N_6383,N_6343);
nor U6481 (N_6481,N_6335,N_6315);
nand U6482 (N_6482,N_6331,N_6340);
nand U6483 (N_6483,N_6390,N_6363);
and U6484 (N_6484,N_6327,N_6378);
or U6485 (N_6485,N_6312,N_6327);
nor U6486 (N_6486,N_6301,N_6346);
or U6487 (N_6487,N_6348,N_6378);
or U6488 (N_6488,N_6370,N_6327);
nor U6489 (N_6489,N_6375,N_6379);
or U6490 (N_6490,N_6393,N_6398);
nor U6491 (N_6491,N_6308,N_6335);
nor U6492 (N_6492,N_6328,N_6399);
nor U6493 (N_6493,N_6352,N_6326);
or U6494 (N_6494,N_6365,N_6367);
and U6495 (N_6495,N_6387,N_6314);
and U6496 (N_6496,N_6327,N_6337);
nand U6497 (N_6497,N_6382,N_6392);
nand U6498 (N_6498,N_6331,N_6354);
nor U6499 (N_6499,N_6393,N_6375);
nand U6500 (N_6500,N_6453,N_6475);
nor U6501 (N_6501,N_6480,N_6420);
nor U6502 (N_6502,N_6403,N_6405);
nor U6503 (N_6503,N_6465,N_6459);
or U6504 (N_6504,N_6424,N_6434);
and U6505 (N_6505,N_6442,N_6401);
or U6506 (N_6506,N_6439,N_6478);
or U6507 (N_6507,N_6444,N_6423);
nor U6508 (N_6508,N_6489,N_6414);
and U6509 (N_6509,N_6448,N_6441);
or U6510 (N_6510,N_6422,N_6494);
nand U6511 (N_6511,N_6493,N_6470);
and U6512 (N_6512,N_6450,N_6429);
or U6513 (N_6513,N_6486,N_6435);
nor U6514 (N_6514,N_6445,N_6467);
or U6515 (N_6515,N_6419,N_6432);
and U6516 (N_6516,N_6454,N_6458);
nand U6517 (N_6517,N_6498,N_6411);
nand U6518 (N_6518,N_6404,N_6447);
nand U6519 (N_6519,N_6416,N_6438);
nand U6520 (N_6520,N_6468,N_6460);
and U6521 (N_6521,N_6483,N_6449);
nor U6522 (N_6522,N_6499,N_6437);
or U6523 (N_6523,N_6410,N_6407);
and U6524 (N_6524,N_6400,N_6473);
nand U6525 (N_6525,N_6463,N_6451);
nor U6526 (N_6526,N_6466,N_6491);
and U6527 (N_6527,N_6477,N_6488);
nor U6528 (N_6528,N_6485,N_6440);
nand U6529 (N_6529,N_6443,N_6479);
nor U6530 (N_6530,N_6430,N_6436);
xor U6531 (N_6531,N_6496,N_6462);
nand U6532 (N_6532,N_6452,N_6408);
and U6533 (N_6533,N_6412,N_6428);
nor U6534 (N_6534,N_6472,N_6476);
and U6535 (N_6535,N_6481,N_6464);
nor U6536 (N_6536,N_6433,N_6409);
and U6537 (N_6537,N_6469,N_6457);
or U6538 (N_6538,N_6431,N_6492);
nand U6539 (N_6539,N_6495,N_6482);
and U6540 (N_6540,N_6455,N_6418);
nand U6541 (N_6541,N_6402,N_6406);
and U6542 (N_6542,N_6484,N_6456);
and U6543 (N_6543,N_6446,N_6421);
nor U6544 (N_6544,N_6487,N_6417);
nor U6545 (N_6545,N_6426,N_6474);
or U6546 (N_6546,N_6415,N_6413);
and U6547 (N_6547,N_6427,N_6471);
or U6548 (N_6548,N_6497,N_6425);
nand U6549 (N_6549,N_6490,N_6461);
nor U6550 (N_6550,N_6402,N_6411);
or U6551 (N_6551,N_6467,N_6491);
nand U6552 (N_6552,N_6409,N_6432);
or U6553 (N_6553,N_6452,N_6422);
or U6554 (N_6554,N_6459,N_6469);
and U6555 (N_6555,N_6439,N_6415);
and U6556 (N_6556,N_6478,N_6423);
or U6557 (N_6557,N_6449,N_6487);
nand U6558 (N_6558,N_6415,N_6483);
or U6559 (N_6559,N_6416,N_6404);
and U6560 (N_6560,N_6409,N_6492);
or U6561 (N_6561,N_6447,N_6488);
or U6562 (N_6562,N_6444,N_6408);
nand U6563 (N_6563,N_6432,N_6415);
nand U6564 (N_6564,N_6478,N_6428);
nand U6565 (N_6565,N_6491,N_6453);
or U6566 (N_6566,N_6426,N_6422);
nor U6567 (N_6567,N_6495,N_6476);
nand U6568 (N_6568,N_6491,N_6454);
nor U6569 (N_6569,N_6496,N_6428);
nand U6570 (N_6570,N_6493,N_6477);
or U6571 (N_6571,N_6451,N_6487);
and U6572 (N_6572,N_6473,N_6476);
nor U6573 (N_6573,N_6447,N_6405);
or U6574 (N_6574,N_6465,N_6485);
nor U6575 (N_6575,N_6470,N_6433);
and U6576 (N_6576,N_6445,N_6452);
nand U6577 (N_6577,N_6429,N_6404);
or U6578 (N_6578,N_6422,N_6400);
nor U6579 (N_6579,N_6453,N_6443);
or U6580 (N_6580,N_6406,N_6454);
and U6581 (N_6581,N_6410,N_6455);
and U6582 (N_6582,N_6416,N_6458);
or U6583 (N_6583,N_6441,N_6432);
nand U6584 (N_6584,N_6465,N_6409);
nand U6585 (N_6585,N_6435,N_6475);
nor U6586 (N_6586,N_6488,N_6438);
nand U6587 (N_6587,N_6464,N_6477);
nand U6588 (N_6588,N_6428,N_6456);
nor U6589 (N_6589,N_6457,N_6463);
nor U6590 (N_6590,N_6455,N_6486);
and U6591 (N_6591,N_6423,N_6469);
nor U6592 (N_6592,N_6425,N_6448);
or U6593 (N_6593,N_6405,N_6445);
nand U6594 (N_6594,N_6416,N_6400);
and U6595 (N_6595,N_6419,N_6454);
or U6596 (N_6596,N_6413,N_6402);
and U6597 (N_6597,N_6478,N_6472);
nand U6598 (N_6598,N_6404,N_6412);
xnor U6599 (N_6599,N_6417,N_6410);
nand U6600 (N_6600,N_6554,N_6511);
or U6601 (N_6601,N_6584,N_6540);
nor U6602 (N_6602,N_6567,N_6575);
nand U6603 (N_6603,N_6520,N_6512);
and U6604 (N_6604,N_6542,N_6592);
or U6605 (N_6605,N_6589,N_6558);
nor U6606 (N_6606,N_6515,N_6591);
and U6607 (N_6607,N_6545,N_6559);
nor U6608 (N_6608,N_6578,N_6583);
and U6609 (N_6609,N_6562,N_6510);
and U6610 (N_6610,N_6555,N_6570);
nand U6611 (N_6611,N_6568,N_6533);
nor U6612 (N_6612,N_6585,N_6576);
nor U6613 (N_6613,N_6560,N_6595);
nand U6614 (N_6614,N_6596,N_6549);
nand U6615 (N_6615,N_6566,N_6507);
nor U6616 (N_6616,N_6594,N_6535);
and U6617 (N_6617,N_6593,N_6504);
nand U6618 (N_6618,N_6538,N_6571);
nor U6619 (N_6619,N_6505,N_6530);
nor U6620 (N_6620,N_6531,N_6574);
nor U6621 (N_6621,N_6541,N_6546);
and U6622 (N_6622,N_6519,N_6527);
nor U6623 (N_6623,N_6547,N_6597);
nand U6624 (N_6624,N_6524,N_6518);
nand U6625 (N_6625,N_6551,N_6572);
or U6626 (N_6626,N_6506,N_6521);
nand U6627 (N_6627,N_6564,N_6561);
and U6628 (N_6628,N_6598,N_6523);
nand U6629 (N_6629,N_6522,N_6586);
nand U6630 (N_6630,N_6563,N_6579);
nand U6631 (N_6631,N_6552,N_6532);
or U6632 (N_6632,N_6543,N_6509);
or U6633 (N_6633,N_6548,N_6588);
nor U6634 (N_6634,N_6526,N_6556);
nor U6635 (N_6635,N_6550,N_6513);
or U6636 (N_6636,N_6581,N_6565);
nor U6637 (N_6637,N_6503,N_6516);
nand U6638 (N_6638,N_6544,N_6577);
nor U6639 (N_6639,N_6514,N_6590);
and U6640 (N_6640,N_6508,N_6539);
nor U6641 (N_6641,N_6582,N_6536);
and U6642 (N_6642,N_6573,N_6557);
nand U6643 (N_6643,N_6537,N_6501);
or U6644 (N_6644,N_6569,N_6553);
or U6645 (N_6645,N_6599,N_6529);
and U6646 (N_6646,N_6500,N_6587);
nor U6647 (N_6647,N_6525,N_6580);
nand U6648 (N_6648,N_6502,N_6517);
nor U6649 (N_6649,N_6534,N_6528);
nor U6650 (N_6650,N_6508,N_6550);
or U6651 (N_6651,N_6595,N_6578);
or U6652 (N_6652,N_6593,N_6579);
nand U6653 (N_6653,N_6539,N_6561);
and U6654 (N_6654,N_6569,N_6547);
nor U6655 (N_6655,N_6536,N_6501);
nor U6656 (N_6656,N_6532,N_6523);
and U6657 (N_6657,N_6584,N_6530);
nand U6658 (N_6658,N_6571,N_6566);
nor U6659 (N_6659,N_6536,N_6506);
or U6660 (N_6660,N_6502,N_6539);
nor U6661 (N_6661,N_6559,N_6509);
and U6662 (N_6662,N_6504,N_6539);
nand U6663 (N_6663,N_6577,N_6536);
and U6664 (N_6664,N_6569,N_6520);
or U6665 (N_6665,N_6500,N_6583);
and U6666 (N_6666,N_6534,N_6550);
nand U6667 (N_6667,N_6534,N_6532);
or U6668 (N_6668,N_6519,N_6591);
or U6669 (N_6669,N_6508,N_6520);
or U6670 (N_6670,N_6590,N_6560);
or U6671 (N_6671,N_6572,N_6524);
or U6672 (N_6672,N_6543,N_6563);
or U6673 (N_6673,N_6569,N_6587);
and U6674 (N_6674,N_6514,N_6535);
and U6675 (N_6675,N_6529,N_6573);
nor U6676 (N_6676,N_6535,N_6516);
nor U6677 (N_6677,N_6555,N_6510);
and U6678 (N_6678,N_6512,N_6507);
nor U6679 (N_6679,N_6569,N_6519);
nand U6680 (N_6680,N_6550,N_6526);
and U6681 (N_6681,N_6532,N_6511);
nor U6682 (N_6682,N_6500,N_6594);
nand U6683 (N_6683,N_6583,N_6590);
nor U6684 (N_6684,N_6543,N_6534);
or U6685 (N_6685,N_6584,N_6559);
or U6686 (N_6686,N_6567,N_6554);
nor U6687 (N_6687,N_6569,N_6552);
nand U6688 (N_6688,N_6523,N_6557);
nand U6689 (N_6689,N_6549,N_6542);
nor U6690 (N_6690,N_6595,N_6516);
or U6691 (N_6691,N_6575,N_6565);
or U6692 (N_6692,N_6597,N_6568);
nand U6693 (N_6693,N_6536,N_6592);
nand U6694 (N_6694,N_6568,N_6535);
nand U6695 (N_6695,N_6574,N_6587);
nand U6696 (N_6696,N_6585,N_6586);
and U6697 (N_6697,N_6516,N_6598);
or U6698 (N_6698,N_6574,N_6538);
nand U6699 (N_6699,N_6567,N_6514);
or U6700 (N_6700,N_6617,N_6650);
or U6701 (N_6701,N_6682,N_6676);
nor U6702 (N_6702,N_6618,N_6606);
nand U6703 (N_6703,N_6655,N_6622);
or U6704 (N_6704,N_6607,N_6610);
nor U6705 (N_6705,N_6604,N_6647);
nand U6706 (N_6706,N_6609,N_6693);
or U6707 (N_6707,N_6602,N_6670);
and U6708 (N_6708,N_6681,N_6654);
nand U6709 (N_6709,N_6687,N_6678);
and U6710 (N_6710,N_6611,N_6661);
nor U6711 (N_6711,N_6630,N_6635);
and U6712 (N_6712,N_6658,N_6633);
or U6713 (N_6713,N_6652,N_6694);
nand U6714 (N_6714,N_6667,N_6668);
nand U6715 (N_6715,N_6675,N_6615);
nand U6716 (N_6716,N_6686,N_6638);
nand U6717 (N_6717,N_6651,N_6653);
nand U6718 (N_6718,N_6628,N_6621);
or U6719 (N_6719,N_6688,N_6665);
and U6720 (N_6720,N_6649,N_6613);
nand U6721 (N_6721,N_6616,N_6679);
and U6722 (N_6722,N_6680,N_6608);
nand U6723 (N_6723,N_6677,N_6674);
nor U6724 (N_6724,N_6657,N_6620);
or U6725 (N_6725,N_6690,N_6669);
and U6726 (N_6726,N_6600,N_6699);
or U6727 (N_6727,N_6637,N_6624);
nand U6728 (N_6728,N_6683,N_6656);
and U6729 (N_6729,N_6629,N_6612);
nor U6730 (N_6730,N_6631,N_6684);
or U6731 (N_6731,N_6696,N_6697);
nor U6732 (N_6732,N_6627,N_6641);
nand U6733 (N_6733,N_6695,N_6634);
and U6734 (N_6734,N_6698,N_6644);
or U6735 (N_6735,N_6645,N_6689);
nor U6736 (N_6736,N_6643,N_6663);
nand U6737 (N_6737,N_6625,N_6660);
and U6738 (N_6738,N_6659,N_6685);
and U6739 (N_6739,N_6691,N_6601);
nand U6740 (N_6740,N_6673,N_6639);
or U6741 (N_6741,N_6664,N_6692);
or U6742 (N_6742,N_6603,N_6626);
nor U6743 (N_6743,N_6605,N_6648);
nand U6744 (N_6744,N_6671,N_6614);
nand U6745 (N_6745,N_6666,N_6636);
nand U6746 (N_6746,N_6619,N_6632);
and U6747 (N_6747,N_6623,N_6662);
nand U6748 (N_6748,N_6646,N_6642);
nor U6749 (N_6749,N_6672,N_6640);
or U6750 (N_6750,N_6651,N_6695);
nand U6751 (N_6751,N_6687,N_6660);
nor U6752 (N_6752,N_6672,N_6658);
or U6753 (N_6753,N_6614,N_6627);
nor U6754 (N_6754,N_6635,N_6610);
and U6755 (N_6755,N_6666,N_6679);
nor U6756 (N_6756,N_6692,N_6630);
or U6757 (N_6757,N_6603,N_6675);
or U6758 (N_6758,N_6630,N_6625);
and U6759 (N_6759,N_6674,N_6632);
or U6760 (N_6760,N_6638,N_6692);
nor U6761 (N_6761,N_6682,N_6688);
and U6762 (N_6762,N_6632,N_6641);
nand U6763 (N_6763,N_6651,N_6661);
nor U6764 (N_6764,N_6683,N_6661);
nor U6765 (N_6765,N_6617,N_6629);
nor U6766 (N_6766,N_6605,N_6626);
nand U6767 (N_6767,N_6614,N_6655);
nor U6768 (N_6768,N_6665,N_6661);
or U6769 (N_6769,N_6666,N_6695);
nand U6770 (N_6770,N_6696,N_6670);
nor U6771 (N_6771,N_6600,N_6631);
nor U6772 (N_6772,N_6650,N_6638);
nor U6773 (N_6773,N_6654,N_6698);
and U6774 (N_6774,N_6602,N_6682);
or U6775 (N_6775,N_6631,N_6642);
nand U6776 (N_6776,N_6647,N_6677);
and U6777 (N_6777,N_6690,N_6623);
or U6778 (N_6778,N_6604,N_6653);
or U6779 (N_6779,N_6656,N_6650);
nand U6780 (N_6780,N_6695,N_6608);
xnor U6781 (N_6781,N_6679,N_6614);
nor U6782 (N_6782,N_6664,N_6601);
and U6783 (N_6783,N_6692,N_6637);
nand U6784 (N_6784,N_6673,N_6602);
nor U6785 (N_6785,N_6646,N_6628);
and U6786 (N_6786,N_6650,N_6647);
nand U6787 (N_6787,N_6647,N_6667);
and U6788 (N_6788,N_6604,N_6641);
nor U6789 (N_6789,N_6677,N_6635);
or U6790 (N_6790,N_6649,N_6636);
nand U6791 (N_6791,N_6657,N_6681);
or U6792 (N_6792,N_6689,N_6669);
nor U6793 (N_6793,N_6662,N_6602);
and U6794 (N_6794,N_6616,N_6655);
nand U6795 (N_6795,N_6622,N_6618);
or U6796 (N_6796,N_6601,N_6661);
nand U6797 (N_6797,N_6662,N_6686);
nand U6798 (N_6798,N_6669,N_6625);
nand U6799 (N_6799,N_6614,N_6693);
nor U6800 (N_6800,N_6774,N_6767);
nor U6801 (N_6801,N_6732,N_6714);
or U6802 (N_6802,N_6758,N_6706);
nor U6803 (N_6803,N_6721,N_6704);
nor U6804 (N_6804,N_6763,N_6727);
and U6805 (N_6805,N_6777,N_6784);
nand U6806 (N_6806,N_6792,N_6779);
or U6807 (N_6807,N_6772,N_6701);
or U6808 (N_6808,N_6768,N_6731);
or U6809 (N_6809,N_6796,N_6776);
nor U6810 (N_6810,N_6755,N_6761);
or U6811 (N_6811,N_6765,N_6798);
and U6812 (N_6812,N_6750,N_6766);
nor U6813 (N_6813,N_6756,N_6795);
or U6814 (N_6814,N_6744,N_6791);
and U6815 (N_6815,N_6726,N_6786);
xnor U6816 (N_6816,N_6753,N_6762);
nand U6817 (N_6817,N_6705,N_6769);
or U6818 (N_6818,N_6720,N_6743);
nand U6819 (N_6819,N_6735,N_6760);
nand U6820 (N_6820,N_6710,N_6700);
or U6821 (N_6821,N_6722,N_6778);
nor U6822 (N_6822,N_6783,N_6738);
nand U6823 (N_6823,N_6707,N_6730);
and U6824 (N_6824,N_6729,N_6747);
nand U6825 (N_6825,N_6703,N_6781);
nand U6826 (N_6826,N_6715,N_6745);
and U6827 (N_6827,N_6718,N_6764);
or U6828 (N_6828,N_6719,N_6742);
and U6829 (N_6829,N_6736,N_6752);
and U6830 (N_6830,N_6788,N_6793);
nand U6831 (N_6831,N_6739,N_6741);
nor U6832 (N_6832,N_6771,N_6787);
and U6833 (N_6833,N_6790,N_6751);
and U6834 (N_6834,N_6757,N_6716);
nand U6835 (N_6835,N_6754,N_6737);
or U6836 (N_6836,N_6717,N_6746);
or U6837 (N_6837,N_6748,N_6711);
and U6838 (N_6838,N_6734,N_6728);
nor U6839 (N_6839,N_6797,N_6780);
nor U6840 (N_6840,N_6799,N_6709);
nor U6841 (N_6841,N_6702,N_6794);
nor U6842 (N_6842,N_6733,N_6785);
nor U6843 (N_6843,N_6740,N_6713);
nor U6844 (N_6844,N_6770,N_6773);
and U6845 (N_6845,N_6789,N_6723);
or U6846 (N_6846,N_6775,N_6708);
or U6847 (N_6847,N_6724,N_6725);
and U6848 (N_6848,N_6759,N_6749);
nor U6849 (N_6849,N_6712,N_6782);
xor U6850 (N_6850,N_6705,N_6794);
and U6851 (N_6851,N_6786,N_6770);
nor U6852 (N_6852,N_6753,N_6795);
nor U6853 (N_6853,N_6774,N_6702);
or U6854 (N_6854,N_6778,N_6710);
nand U6855 (N_6855,N_6721,N_6754);
or U6856 (N_6856,N_6709,N_6756);
nand U6857 (N_6857,N_6712,N_6727);
nor U6858 (N_6858,N_6771,N_6714);
or U6859 (N_6859,N_6736,N_6728);
nor U6860 (N_6860,N_6753,N_6718);
nand U6861 (N_6861,N_6762,N_6749);
nand U6862 (N_6862,N_6769,N_6772);
nor U6863 (N_6863,N_6799,N_6772);
and U6864 (N_6864,N_6716,N_6727);
and U6865 (N_6865,N_6726,N_6788);
or U6866 (N_6866,N_6732,N_6766);
or U6867 (N_6867,N_6763,N_6703);
and U6868 (N_6868,N_6789,N_6704);
and U6869 (N_6869,N_6784,N_6733);
and U6870 (N_6870,N_6769,N_6714);
nand U6871 (N_6871,N_6749,N_6787);
and U6872 (N_6872,N_6783,N_6780);
nand U6873 (N_6873,N_6799,N_6703);
and U6874 (N_6874,N_6733,N_6758);
and U6875 (N_6875,N_6731,N_6788);
or U6876 (N_6876,N_6708,N_6784);
or U6877 (N_6877,N_6744,N_6784);
nand U6878 (N_6878,N_6778,N_6705);
and U6879 (N_6879,N_6768,N_6786);
nand U6880 (N_6880,N_6712,N_6764);
nor U6881 (N_6881,N_6759,N_6765);
and U6882 (N_6882,N_6744,N_6775);
or U6883 (N_6883,N_6786,N_6795);
nor U6884 (N_6884,N_6737,N_6789);
and U6885 (N_6885,N_6739,N_6743);
and U6886 (N_6886,N_6793,N_6723);
or U6887 (N_6887,N_6729,N_6743);
nor U6888 (N_6888,N_6787,N_6729);
nor U6889 (N_6889,N_6710,N_6773);
nand U6890 (N_6890,N_6775,N_6776);
nand U6891 (N_6891,N_6732,N_6749);
xor U6892 (N_6892,N_6707,N_6784);
or U6893 (N_6893,N_6706,N_6734);
nand U6894 (N_6894,N_6752,N_6779);
nand U6895 (N_6895,N_6700,N_6718);
nand U6896 (N_6896,N_6761,N_6723);
nor U6897 (N_6897,N_6794,N_6755);
or U6898 (N_6898,N_6757,N_6712);
nand U6899 (N_6899,N_6747,N_6777);
nand U6900 (N_6900,N_6888,N_6828);
and U6901 (N_6901,N_6887,N_6801);
nand U6902 (N_6902,N_6841,N_6890);
nor U6903 (N_6903,N_6820,N_6860);
and U6904 (N_6904,N_6842,N_6897);
nand U6905 (N_6905,N_6822,N_6800);
or U6906 (N_6906,N_6829,N_6813);
or U6907 (N_6907,N_6864,N_6831);
or U6908 (N_6908,N_6825,N_6858);
nand U6909 (N_6909,N_6830,N_6861);
nor U6910 (N_6910,N_6877,N_6810);
and U6911 (N_6911,N_6847,N_6856);
and U6912 (N_6912,N_6863,N_6803);
nand U6913 (N_6913,N_6804,N_6815);
nor U6914 (N_6914,N_6846,N_6859);
or U6915 (N_6915,N_6816,N_6896);
and U6916 (N_6916,N_6806,N_6850);
and U6917 (N_6917,N_6873,N_6870);
nor U6918 (N_6918,N_6805,N_6811);
nand U6919 (N_6919,N_6840,N_6832);
or U6920 (N_6920,N_6817,N_6876);
nand U6921 (N_6921,N_6882,N_6869);
nor U6922 (N_6922,N_6821,N_6866);
and U6923 (N_6923,N_6892,N_6855);
nor U6924 (N_6924,N_6885,N_6871);
or U6925 (N_6925,N_6898,N_6853);
nor U6926 (N_6926,N_6894,N_6835);
nand U6927 (N_6927,N_6891,N_6844);
nor U6928 (N_6928,N_6867,N_6893);
or U6929 (N_6929,N_6838,N_6807);
and U6930 (N_6930,N_6833,N_6818);
nor U6931 (N_6931,N_6884,N_6843);
nor U6932 (N_6932,N_6880,N_6845);
nand U6933 (N_6933,N_6854,N_6883);
or U6934 (N_6934,N_6879,N_6851);
nor U6935 (N_6935,N_6862,N_6819);
and U6936 (N_6936,N_6872,N_6834);
and U6937 (N_6937,N_6823,N_6899);
nor U6938 (N_6938,N_6802,N_6881);
or U6939 (N_6939,N_6865,N_6848);
or U6940 (N_6940,N_6827,N_6812);
and U6941 (N_6941,N_6889,N_6874);
nor U6942 (N_6942,N_6878,N_6849);
nor U6943 (N_6943,N_6857,N_6852);
and U6944 (N_6944,N_6886,N_6824);
and U6945 (N_6945,N_6814,N_6839);
and U6946 (N_6946,N_6895,N_6826);
nor U6947 (N_6947,N_6875,N_6836);
and U6948 (N_6948,N_6809,N_6837);
or U6949 (N_6949,N_6808,N_6868);
or U6950 (N_6950,N_6835,N_6843);
nor U6951 (N_6951,N_6833,N_6847);
or U6952 (N_6952,N_6873,N_6825);
nor U6953 (N_6953,N_6852,N_6856);
and U6954 (N_6954,N_6862,N_6842);
or U6955 (N_6955,N_6840,N_6830);
nand U6956 (N_6956,N_6800,N_6834);
and U6957 (N_6957,N_6832,N_6873);
or U6958 (N_6958,N_6868,N_6819);
and U6959 (N_6959,N_6800,N_6864);
and U6960 (N_6960,N_6875,N_6838);
and U6961 (N_6961,N_6836,N_6833);
or U6962 (N_6962,N_6867,N_6817);
and U6963 (N_6963,N_6878,N_6888);
nand U6964 (N_6964,N_6806,N_6868);
nand U6965 (N_6965,N_6857,N_6836);
or U6966 (N_6966,N_6844,N_6848);
nand U6967 (N_6967,N_6804,N_6845);
or U6968 (N_6968,N_6836,N_6865);
nand U6969 (N_6969,N_6877,N_6862);
or U6970 (N_6970,N_6835,N_6818);
nand U6971 (N_6971,N_6849,N_6860);
and U6972 (N_6972,N_6834,N_6863);
and U6973 (N_6973,N_6852,N_6827);
xor U6974 (N_6974,N_6865,N_6810);
nand U6975 (N_6975,N_6847,N_6864);
nand U6976 (N_6976,N_6871,N_6808);
and U6977 (N_6977,N_6866,N_6809);
and U6978 (N_6978,N_6843,N_6877);
or U6979 (N_6979,N_6826,N_6879);
nand U6980 (N_6980,N_6885,N_6876);
or U6981 (N_6981,N_6847,N_6898);
or U6982 (N_6982,N_6899,N_6861);
and U6983 (N_6983,N_6817,N_6863);
or U6984 (N_6984,N_6837,N_6831);
nor U6985 (N_6985,N_6857,N_6896);
and U6986 (N_6986,N_6883,N_6868);
nor U6987 (N_6987,N_6861,N_6843);
nand U6988 (N_6988,N_6813,N_6815);
or U6989 (N_6989,N_6805,N_6842);
and U6990 (N_6990,N_6831,N_6886);
nand U6991 (N_6991,N_6893,N_6865);
and U6992 (N_6992,N_6890,N_6842);
nand U6993 (N_6993,N_6899,N_6820);
nand U6994 (N_6994,N_6892,N_6899);
or U6995 (N_6995,N_6893,N_6837);
nor U6996 (N_6996,N_6872,N_6894);
and U6997 (N_6997,N_6882,N_6802);
xor U6998 (N_6998,N_6806,N_6829);
xnor U6999 (N_6999,N_6850,N_6883);
or U7000 (N_7000,N_6977,N_6986);
nand U7001 (N_7001,N_6962,N_6918);
nand U7002 (N_7002,N_6942,N_6923);
nand U7003 (N_7003,N_6961,N_6906);
nor U7004 (N_7004,N_6936,N_6985);
and U7005 (N_7005,N_6904,N_6957);
and U7006 (N_7006,N_6975,N_6968);
or U7007 (N_7007,N_6970,N_6994);
nand U7008 (N_7008,N_6967,N_6955);
or U7009 (N_7009,N_6914,N_6941);
nor U7010 (N_7010,N_6979,N_6954);
nand U7011 (N_7011,N_6921,N_6989);
nand U7012 (N_7012,N_6964,N_6971);
nand U7013 (N_7013,N_6931,N_6963);
and U7014 (N_7014,N_6910,N_6908);
or U7015 (N_7015,N_6902,N_6912);
nor U7016 (N_7016,N_6987,N_6973);
and U7017 (N_7017,N_6956,N_6980);
nand U7018 (N_7018,N_6969,N_6903);
nand U7019 (N_7019,N_6959,N_6927);
nand U7020 (N_7020,N_6983,N_6911);
nor U7021 (N_7021,N_6992,N_6938);
nor U7022 (N_7022,N_6990,N_6966);
or U7023 (N_7023,N_6976,N_6993);
nor U7024 (N_7024,N_6939,N_6972);
nand U7025 (N_7025,N_6949,N_6948);
nor U7026 (N_7026,N_6947,N_6926);
or U7027 (N_7027,N_6943,N_6929);
and U7028 (N_7028,N_6999,N_6919);
nor U7029 (N_7029,N_6981,N_6960);
and U7030 (N_7030,N_6982,N_6998);
or U7031 (N_7031,N_6924,N_6900);
or U7032 (N_7032,N_6984,N_6917);
nand U7033 (N_7033,N_6934,N_6952);
and U7034 (N_7034,N_6925,N_6913);
or U7035 (N_7035,N_6928,N_6920);
or U7036 (N_7036,N_6953,N_6915);
or U7037 (N_7037,N_6901,N_6940);
nand U7038 (N_7038,N_6944,N_6951);
or U7039 (N_7039,N_6974,N_6988);
or U7040 (N_7040,N_6996,N_6933);
nor U7041 (N_7041,N_6909,N_6995);
or U7042 (N_7042,N_6932,N_6907);
nor U7043 (N_7043,N_6997,N_6978);
nand U7044 (N_7044,N_6946,N_6950);
and U7045 (N_7045,N_6922,N_6916);
nor U7046 (N_7046,N_6937,N_6958);
xnor U7047 (N_7047,N_6991,N_6945);
nand U7048 (N_7048,N_6965,N_6935);
nand U7049 (N_7049,N_6930,N_6905);
nor U7050 (N_7050,N_6909,N_6968);
and U7051 (N_7051,N_6949,N_6964);
nor U7052 (N_7052,N_6955,N_6996);
nor U7053 (N_7053,N_6975,N_6938);
and U7054 (N_7054,N_6947,N_6973);
and U7055 (N_7055,N_6993,N_6945);
nor U7056 (N_7056,N_6972,N_6989);
or U7057 (N_7057,N_6947,N_6982);
and U7058 (N_7058,N_6992,N_6936);
nor U7059 (N_7059,N_6920,N_6927);
nand U7060 (N_7060,N_6970,N_6981);
nor U7061 (N_7061,N_6909,N_6925);
and U7062 (N_7062,N_6962,N_6953);
nor U7063 (N_7063,N_6958,N_6924);
nor U7064 (N_7064,N_6944,N_6980);
or U7065 (N_7065,N_6977,N_6972);
or U7066 (N_7066,N_6941,N_6958);
or U7067 (N_7067,N_6963,N_6949);
nand U7068 (N_7068,N_6903,N_6992);
nand U7069 (N_7069,N_6995,N_6987);
nor U7070 (N_7070,N_6961,N_6992);
or U7071 (N_7071,N_6924,N_6934);
or U7072 (N_7072,N_6996,N_6989);
and U7073 (N_7073,N_6980,N_6996);
nand U7074 (N_7074,N_6926,N_6986);
and U7075 (N_7075,N_6900,N_6940);
or U7076 (N_7076,N_6999,N_6958);
or U7077 (N_7077,N_6983,N_6976);
and U7078 (N_7078,N_6918,N_6933);
and U7079 (N_7079,N_6963,N_6962);
nor U7080 (N_7080,N_6968,N_6956);
nand U7081 (N_7081,N_6984,N_6926);
nand U7082 (N_7082,N_6924,N_6921);
nand U7083 (N_7083,N_6954,N_6984);
nor U7084 (N_7084,N_6916,N_6915);
and U7085 (N_7085,N_6951,N_6990);
or U7086 (N_7086,N_6994,N_6943);
and U7087 (N_7087,N_6923,N_6953);
nand U7088 (N_7088,N_6926,N_6901);
and U7089 (N_7089,N_6949,N_6936);
and U7090 (N_7090,N_6930,N_6944);
nor U7091 (N_7091,N_6959,N_6905);
nand U7092 (N_7092,N_6993,N_6989);
nor U7093 (N_7093,N_6980,N_6925);
nand U7094 (N_7094,N_6933,N_6964);
and U7095 (N_7095,N_6926,N_6982);
or U7096 (N_7096,N_6954,N_6987);
nand U7097 (N_7097,N_6908,N_6920);
and U7098 (N_7098,N_6901,N_6914);
or U7099 (N_7099,N_6916,N_6988);
and U7100 (N_7100,N_7030,N_7016);
and U7101 (N_7101,N_7058,N_7036);
nand U7102 (N_7102,N_7096,N_7064);
or U7103 (N_7103,N_7060,N_7006);
nor U7104 (N_7104,N_7057,N_7054);
and U7105 (N_7105,N_7012,N_7069);
and U7106 (N_7106,N_7004,N_7075);
and U7107 (N_7107,N_7090,N_7098);
nor U7108 (N_7108,N_7003,N_7034);
nor U7109 (N_7109,N_7013,N_7040);
and U7110 (N_7110,N_7084,N_7053);
and U7111 (N_7111,N_7005,N_7026);
nor U7112 (N_7112,N_7021,N_7094);
and U7113 (N_7113,N_7091,N_7068);
nor U7114 (N_7114,N_7048,N_7043);
or U7115 (N_7115,N_7056,N_7024);
and U7116 (N_7116,N_7038,N_7039);
nor U7117 (N_7117,N_7059,N_7099);
nand U7118 (N_7118,N_7033,N_7015);
nand U7119 (N_7119,N_7007,N_7028);
and U7120 (N_7120,N_7000,N_7001);
and U7121 (N_7121,N_7083,N_7041);
nand U7122 (N_7122,N_7020,N_7002);
nand U7123 (N_7123,N_7049,N_7022);
or U7124 (N_7124,N_7087,N_7050);
or U7125 (N_7125,N_7080,N_7037);
nor U7126 (N_7126,N_7070,N_7067);
nand U7127 (N_7127,N_7044,N_7093);
and U7128 (N_7128,N_7063,N_7011);
or U7129 (N_7129,N_7092,N_7079);
nor U7130 (N_7130,N_7074,N_7061);
and U7131 (N_7131,N_7081,N_7095);
or U7132 (N_7132,N_7086,N_7023);
and U7133 (N_7133,N_7029,N_7066);
and U7134 (N_7134,N_7010,N_7042);
xor U7135 (N_7135,N_7027,N_7089);
and U7136 (N_7136,N_7065,N_7035);
and U7137 (N_7137,N_7045,N_7097);
and U7138 (N_7138,N_7076,N_7078);
or U7139 (N_7139,N_7077,N_7052);
and U7140 (N_7140,N_7062,N_7009);
nand U7141 (N_7141,N_7072,N_7071);
nor U7142 (N_7142,N_7082,N_7019);
and U7143 (N_7143,N_7073,N_7031);
or U7144 (N_7144,N_7008,N_7085);
nand U7145 (N_7145,N_7046,N_7018);
nor U7146 (N_7146,N_7088,N_7017);
and U7147 (N_7147,N_7032,N_7025);
or U7148 (N_7148,N_7055,N_7047);
nor U7149 (N_7149,N_7051,N_7014);
or U7150 (N_7150,N_7040,N_7017);
and U7151 (N_7151,N_7071,N_7064);
and U7152 (N_7152,N_7001,N_7057);
and U7153 (N_7153,N_7055,N_7028);
nand U7154 (N_7154,N_7035,N_7008);
nand U7155 (N_7155,N_7093,N_7014);
nand U7156 (N_7156,N_7010,N_7076);
nand U7157 (N_7157,N_7077,N_7066);
and U7158 (N_7158,N_7058,N_7020);
and U7159 (N_7159,N_7042,N_7001);
and U7160 (N_7160,N_7070,N_7029);
nor U7161 (N_7161,N_7071,N_7030);
and U7162 (N_7162,N_7079,N_7016);
and U7163 (N_7163,N_7085,N_7014);
and U7164 (N_7164,N_7015,N_7068);
nor U7165 (N_7165,N_7064,N_7091);
nand U7166 (N_7166,N_7081,N_7096);
nand U7167 (N_7167,N_7078,N_7001);
nand U7168 (N_7168,N_7014,N_7087);
nor U7169 (N_7169,N_7054,N_7097);
nand U7170 (N_7170,N_7024,N_7009);
nor U7171 (N_7171,N_7062,N_7029);
nand U7172 (N_7172,N_7056,N_7079);
nand U7173 (N_7173,N_7086,N_7093);
or U7174 (N_7174,N_7086,N_7053);
nand U7175 (N_7175,N_7002,N_7059);
and U7176 (N_7176,N_7065,N_7097);
nor U7177 (N_7177,N_7000,N_7073);
and U7178 (N_7178,N_7091,N_7076);
nor U7179 (N_7179,N_7020,N_7029);
nor U7180 (N_7180,N_7008,N_7081);
nor U7181 (N_7181,N_7055,N_7061);
nor U7182 (N_7182,N_7099,N_7046);
and U7183 (N_7183,N_7037,N_7031);
nand U7184 (N_7184,N_7086,N_7015);
nand U7185 (N_7185,N_7022,N_7038);
nor U7186 (N_7186,N_7092,N_7055);
nor U7187 (N_7187,N_7002,N_7019);
nor U7188 (N_7188,N_7033,N_7077);
or U7189 (N_7189,N_7010,N_7064);
nand U7190 (N_7190,N_7018,N_7050);
and U7191 (N_7191,N_7026,N_7041);
nand U7192 (N_7192,N_7040,N_7084);
and U7193 (N_7193,N_7087,N_7034);
nand U7194 (N_7194,N_7092,N_7030);
or U7195 (N_7195,N_7079,N_7002);
nor U7196 (N_7196,N_7020,N_7038);
nor U7197 (N_7197,N_7051,N_7076);
nand U7198 (N_7198,N_7052,N_7027);
nand U7199 (N_7199,N_7031,N_7066);
or U7200 (N_7200,N_7188,N_7197);
and U7201 (N_7201,N_7160,N_7155);
and U7202 (N_7202,N_7169,N_7178);
or U7203 (N_7203,N_7193,N_7116);
and U7204 (N_7204,N_7183,N_7107);
nor U7205 (N_7205,N_7121,N_7196);
nand U7206 (N_7206,N_7198,N_7148);
nand U7207 (N_7207,N_7125,N_7119);
nand U7208 (N_7208,N_7152,N_7165);
or U7209 (N_7209,N_7129,N_7156);
and U7210 (N_7210,N_7130,N_7115);
nor U7211 (N_7211,N_7185,N_7147);
nand U7212 (N_7212,N_7184,N_7162);
nand U7213 (N_7213,N_7138,N_7164);
or U7214 (N_7214,N_7131,N_7114);
and U7215 (N_7215,N_7167,N_7109);
nor U7216 (N_7216,N_7182,N_7199);
nand U7217 (N_7217,N_7179,N_7166);
and U7218 (N_7218,N_7157,N_7192);
nand U7219 (N_7219,N_7117,N_7126);
and U7220 (N_7220,N_7105,N_7144);
nand U7221 (N_7221,N_7139,N_7189);
or U7222 (N_7222,N_7175,N_7103);
or U7223 (N_7223,N_7151,N_7123);
nor U7224 (N_7224,N_7141,N_7191);
nor U7225 (N_7225,N_7195,N_7140);
nand U7226 (N_7226,N_7146,N_7186);
or U7227 (N_7227,N_7137,N_7190);
nor U7228 (N_7228,N_7106,N_7118);
nand U7229 (N_7229,N_7120,N_7172);
or U7230 (N_7230,N_7154,N_7110);
nor U7231 (N_7231,N_7142,N_7122);
nor U7232 (N_7232,N_7127,N_7145);
nand U7233 (N_7233,N_7168,N_7149);
and U7234 (N_7234,N_7171,N_7143);
and U7235 (N_7235,N_7134,N_7111);
or U7236 (N_7236,N_7101,N_7163);
or U7237 (N_7237,N_7187,N_7108);
nor U7238 (N_7238,N_7124,N_7159);
or U7239 (N_7239,N_7100,N_7136);
and U7240 (N_7240,N_7181,N_7112);
or U7241 (N_7241,N_7102,N_7150);
nand U7242 (N_7242,N_7128,N_7174);
nor U7243 (N_7243,N_7135,N_7161);
nor U7244 (N_7244,N_7158,N_7170);
nand U7245 (N_7245,N_7104,N_7194);
or U7246 (N_7246,N_7177,N_7176);
or U7247 (N_7247,N_7133,N_7180);
nand U7248 (N_7248,N_7173,N_7132);
or U7249 (N_7249,N_7113,N_7153);
nand U7250 (N_7250,N_7159,N_7137);
nand U7251 (N_7251,N_7195,N_7121);
and U7252 (N_7252,N_7172,N_7162);
or U7253 (N_7253,N_7104,N_7114);
nand U7254 (N_7254,N_7123,N_7165);
nor U7255 (N_7255,N_7182,N_7124);
and U7256 (N_7256,N_7145,N_7111);
nor U7257 (N_7257,N_7162,N_7165);
nand U7258 (N_7258,N_7140,N_7141);
nor U7259 (N_7259,N_7198,N_7121);
and U7260 (N_7260,N_7115,N_7132);
or U7261 (N_7261,N_7114,N_7137);
nor U7262 (N_7262,N_7172,N_7152);
nand U7263 (N_7263,N_7135,N_7126);
nand U7264 (N_7264,N_7100,N_7110);
or U7265 (N_7265,N_7196,N_7151);
nand U7266 (N_7266,N_7124,N_7101);
nand U7267 (N_7267,N_7158,N_7141);
nor U7268 (N_7268,N_7160,N_7131);
and U7269 (N_7269,N_7158,N_7125);
or U7270 (N_7270,N_7101,N_7195);
nor U7271 (N_7271,N_7149,N_7161);
or U7272 (N_7272,N_7114,N_7153);
nor U7273 (N_7273,N_7116,N_7173);
and U7274 (N_7274,N_7130,N_7122);
and U7275 (N_7275,N_7141,N_7165);
nand U7276 (N_7276,N_7148,N_7115);
and U7277 (N_7277,N_7190,N_7121);
and U7278 (N_7278,N_7176,N_7187);
nor U7279 (N_7279,N_7197,N_7104);
and U7280 (N_7280,N_7166,N_7156);
nand U7281 (N_7281,N_7173,N_7155);
and U7282 (N_7282,N_7177,N_7191);
and U7283 (N_7283,N_7153,N_7198);
or U7284 (N_7284,N_7106,N_7193);
and U7285 (N_7285,N_7127,N_7164);
and U7286 (N_7286,N_7194,N_7181);
nand U7287 (N_7287,N_7140,N_7148);
and U7288 (N_7288,N_7112,N_7190);
nor U7289 (N_7289,N_7178,N_7163);
and U7290 (N_7290,N_7195,N_7134);
nand U7291 (N_7291,N_7127,N_7105);
and U7292 (N_7292,N_7131,N_7135);
nor U7293 (N_7293,N_7103,N_7181);
nand U7294 (N_7294,N_7145,N_7112);
or U7295 (N_7295,N_7141,N_7187);
or U7296 (N_7296,N_7112,N_7108);
nor U7297 (N_7297,N_7182,N_7144);
or U7298 (N_7298,N_7118,N_7145);
nand U7299 (N_7299,N_7189,N_7149);
nor U7300 (N_7300,N_7221,N_7232);
and U7301 (N_7301,N_7200,N_7275);
nor U7302 (N_7302,N_7210,N_7294);
or U7303 (N_7303,N_7278,N_7204);
or U7304 (N_7304,N_7226,N_7218);
and U7305 (N_7305,N_7240,N_7276);
nor U7306 (N_7306,N_7252,N_7260);
nor U7307 (N_7307,N_7238,N_7215);
nand U7308 (N_7308,N_7250,N_7243);
nor U7309 (N_7309,N_7203,N_7245);
or U7310 (N_7310,N_7220,N_7213);
nor U7311 (N_7311,N_7290,N_7239);
nor U7312 (N_7312,N_7255,N_7228);
nand U7313 (N_7313,N_7280,N_7265);
nor U7314 (N_7314,N_7281,N_7216);
and U7315 (N_7315,N_7282,N_7211);
nand U7316 (N_7316,N_7296,N_7268);
and U7317 (N_7317,N_7297,N_7225);
or U7318 (N_7318,N_7230,N_7235);
xnor U7319 (N_7319,N_7234,N_7244);
and U7320 (N_7320,N_7246,N_7273);
or U7321 (N_7321,N_7269,N_7242);
or U7322 (N_7322,N_7262,N_7208);
or U7323 (N_7323,N_7298,N_7258);
nand U7324 (N_7324,N_7251,N_7287);
and U7325 (N_7325,N_7267,N_7272);
and U7326 (N_7326,N_7224,N_7249);
or U7327 (N_7327,N_7241,N_7285);
nand U7328 (N_7328,N_7299,N_7219);
and U7329 (N_7329,N_7233,N_7217);
or U7330 (N_7330,N_7236,N_7266);
nand U7331 (N_7331,N_7205,N_7231);
and U7332 (N_7332,N_7214,N_7286);
nand U7333 (N_7333,N_7229,N_7289);
and U7334 (N_7334,N_7209,N_7253);
nor U7335 (N_7335,N_7259,N_7206);
xor U7336 (N_7336,N_7207,N_7254);
and U7337 (N_7337,N_7222,N_7270);
or U7338 (N_7338,N_7248,N_7293);
nand U7339 (N_7339,N_7295,N_7201);
and U7340 (N_7340,N_7263,N_7256);
or U7341 (N_7341,N_7212,N_7202);
nand U7342 (N_7342,N_7257,N_7247);
and U7343 (N_7343,N_7227,N_7274);
or U7344 (N_7344,N_7261,N_7292);
nor U7345 (N_7345,N_7277,N_7264);
or U7346 (N_7346,N_7237,N_7284);
and U7347 (N_7347,N_7279,N_7271);
or U7348 (N_7348,N_7291,N_7288);
and U7349 (N_7349,N_7223,N_7283);
or U7350 (N_7350,N_7269,N_7239);
or U7351 (N_7351,N_7231,N_7282);
or U7352 (N_7352,N_7203,N_7246);
nand U7353 (N_7353,N_7206,N_7264);
and U7354 (N_7354,N_7268,N_7248);
nand U7355 (N_7355,N_7259,N_7201);
nand U7356 (N_7356,N_7267,N_7283);
nor U7357 (N_7357,N_7236,N_7240);
nor U7358 (N_7358,N_7203,N_7205);
nand U7359 (N_7359,N_7212,N_7205);
xnor U7360 (N_7360,N_7200,N_7204);
or U7361 (N_7361,N_7246,N_7223);
or U7362 (N_7362,N_7236,N_7285);
nand U7363 (N_7363,N_7271,N_7241);
nand U7364 (N_7364,N_7236,N_7256);
or U7365 (N_7365,N_7222,N_7248);
or U7366 (N_7366,N_7245,N_7248);
nand U7367 (N_7367,N_7206,N_7201);
nand U7368 (N_7368,N_7254,N_7242);
and U7369 (N_7369,N_7287,N_7228);
nor U7370 (N_7370,N_7246,N_7209);
and U7371 (N_7371,N_7247,N_7276);
and U7372 (N_7372,N_7203,N_7278);
nand U7373 (N_7373,N_7267,N_7206);
and U7374 (N_7374,N_7280,N_7248);
and U7375 (N_7375,N_7217,N_7222);
and U7376 (N_7376,N_7217,N_7223);
nand U7377 (N_7377,N_7274,N_7281);
or U7378 (N_7378,N_7290,N_7255);
or U7379 (N_7379,N_7278,N_7234);
and U7380 (N_7380,N_7266,N_7247);
or U7381 (N_7381,N_7227,N_7263);
and U7382 (N_7382,N_7284,N_7293);
or U7383 (N_7383,N_7213,N_7247);
and U7384 (N_7384,N_7273,N_7235);
nand U7385 (N_7385,N_7262,N_7201);
nand U7386 (N_7386,N_7221,N_7207);
nor U7387 (N_7387,N_7296,N_7244);
and U7388 (N_7388,N_7270,N_7230);
and U7389 (N_7389,N_7237,N_7236);
and U7390 (N_7390,N_7246,N_7241);
nand U7391 (N_7391,N_7252,N_7208);
and U7392 (N_7392,N_7285,N_7244);
nor U7393 (N_7393,N_7245,N_7223);
and U7394 (N_7394,N_7257,N_7209);
nand U7395 (N_7395,N_7293,N_7230);
or U7396 (N_7396,N_7216,N_7285);
or U7397 (N_7397,N_7284,N_7297);
nor U7398 (N_7398,N_7204,N_7270);
nand U7399 (N_7399,N_7214,N_7257);
nor U7400 (N_7400,N_7329,N_7326);
and U7401 (N_7401,N_7324,N_7355);
nand U7402 (N_7402,N_7320,N_7399);
nor U7403 (N_7403,N_7304,N_7305);
and U7404 (N_7404,N_7354,N_7358);
nor U7405 (N_7405,N_7362,N_7378);
nor U7406 (N_7406,N_7350,N_7356);
nor U7407 (N_7407,N_7353,N_7366);
nor U7408 (N_7408,N_7322,N_7334);
and U7409 (N_7409,N_7365,N_7376);
and U7410 (N_7410,N_7339,N_7300);
nor U7411 (N_7411,N_7340,N_7374);
nand U7412 (N_7412,N_7335,N_7333);
nor U7413 (N_7413,N_7342,N_7313);
nand U7414 (N_7414,N_7372,N_7325);
nand U7415 (N_7415,N_7397,N_7386);
or U7416 (N_7416,N_7381,N_7363);
or U7417 (N_7417,N_7343,N_7392);
nor U7418 (N_7418,N_7337,N_7341);
and U7419 (N_7419,N_7328,N_7383);
nor U7420 (N_7420,N_7314,N_7375);
nand U7421 (N_7421,N_7323,N_7351);
and U7422 (N_7422,N_7308,N_7389);
or U7423 (N_7423,N_7338,N_7385);
and U7424 (N_7424,N_7331,N_7315);
nand U7425 (N_7425,N_7371,N_7349);
nand U7426 (N_7426,N_7307,N_7398);
or U7427 (N_7427,N_7318,N_7346);
or U7428 (N_7428,N_7306,N_7391);
and U7429 (N_7429,N_7317,N_7367);
nand U7430 (N_7430,N_7312,N_7319);
nand U7431 (N_7431,N_7384,N_7332);
and U7432 (N_7432,N_7388,N_7345);
nor U7433 (N_7433,N_7327,N_7368);
nand U7434 (N_7434,N_7379,N_7382);
or U7435 (N_7435,N_7393,N_7321);
nand U7436 (N_7436,N_7380,N_7373);
nand U7437 (N_7437,N_7396,N_7336);
nand U7438 (N_7438,N_7344,N_7361);
or U7439 (N_7439,N_7301,N_7348);
and U7440 (N_7440,N_7360,N_7359);
or U7441 (N_7441,N_7387,N_7302);
and U7442 (N_7442,N_7311,N_7309);
nor U7443 (N_7443,N_7316,N_7394);
or U7444 (N_7444,N_7330,N_7395);
and U7445 (N_7445,N_7370,N_7310);
nand U7446 (N_7446,N_7369,N_7364);
or U7447 (N_7447,N_7352,N_7357);
and U7448 (N_7448,N_7377,N_7390);
and U7449 (N_7449,N_7303,N_7347);
nand U7450 (N_7450,N_7342,N_7390);
nand U7451 (N_7451,N_7397,N_7326);
nor U7452 (N_7452,N_7395,N_7327);
or U7453 (N_7453,N_7379,N_7344);
and U7454 (N_7454,N_7350,N_7392);
or U7455 (N_7455,N_7307,N_7325);
nand U7456 (N_7456,N_7315,N_7384);
or U7457 (N_7457,N_7340,N_7391);
nand U7458 (N_7458,N_7381,N_7334);
nand U7459 (N_7459,N_7368,N_7381);
nor U7460 (N_7460,N_7370,N_7320);
and U7461 (N_7461,N_7320,N_7338);
or U7462 (N_7462,N_7332,N_7351);
nand U7463 (N_7463,N_7375,N_7341);
or U7464 (N_7464,N_7321,N_7351);
and U7465 (N_7465,N_7362,N_7381);
nand U7466 (N_7466,N_7346,N_7366);
or U7467 (N_7467,N_7310,N_7362);
nor U7468 (N_7468,N_7358,N_7311);
nor U7469 (N_7469,N_7390,N_7364);
and U7470 (N_7470,N_7306,N_7302);
nand U7471 (N_7471,N_7317,N_7387);
nor U7472 (N_7472,N_7341,N_7352);
nand U7473 (N_7473,N_7388,N_7327);
or U7474 (N_7474,N_7302,N_7394);
or U7475 (N_7475,N_7338,N_7394);
nand U7476 (N_7476,N_7349,N_7302);
nand U7477 (N_7477,N_7336,N_7393);
nor U7478 (N_7478,N_7394,N_7354);
and U7479 (N_7479,N_7385,N_7378);
and U7480 (N_7480,N_7316,N_7355);
nand U7481 (N_7481,N_7394,N_7374);
nor U7482 (N_7482,N_7368,N_7385);
or U7483 (N_7483,N_7366,N_7345);
and U7484 (N_7484,N_7394,N_7339);
nand U7485 (N_7485,N_7396,N_7303);
nand U7486 (N_7486,N_7371,N_7311);
nor U7487 (N_7487,N_7319,N_7302);
or U7488 (N_7488,N_7304,N_7331);
nor U7489 (N_7489,N_7388,N_7343);
and U7490 (N_7490,N_7386,N_7365);
nor U7491 (N_7491,N_7361,N_7387);
nor U7492 (N_7492,N_7334,N_7336);
or U7493 (N_7493,N_7377,N_7360);
nand U7494 (N_7494,N_7373,N_7318);
nor U7495 (N_7495,N_7337,N_7375);
or U7496 (N_7496,N_7393,N_7318);
nand U7497 (N_7497,N_7310,N_7390);
or U7498 (N_7498,N_7388,N_7318);
or U7499 (N_7499,N_7397,N_7366);
nand U7500 (N_7500,N_7495,N_7434);
and U7501 (N_7501,N_7449,N_7462);
nand U7502 (N_7502,N_7498,N_7458);
nor U7503 (N_7503,N_7418,N_7461);
or U7504 (N_7504,N_7435,N_7417);
nand U7505 (N_7505,N_7481,N_7452);
and U7506 (N_7506,N_7478,N_7402);
and U7507 (N_7507,N_7406,N_7493);
and U7508 (N_7508,N_7499,N_7484);
or U7509 (N_7509,N_7487,N_7473);
or U7510 (N_7510,N_7467,N_7422);
nand U7511 (N_7511,N_7455,N_7491);
nand U7512 (N_7512,N_7486,N_7414);
nand U7513 (N_7513,N_7446,N_7415);
or U7514 (N_7514,N_7450,N_7469);
and U7515 (N_7515,N_7483,N_7423);
or U7516 (N_7516,N_7447,N_7464);
and U7517 (N_7517,N_7477,N_7416);
and U7518 (N_7518,N_7408,N_7465);
and U7519 (N_7519,N_7492,N_7440);
or U7520 (N_7520,N_7488,N_7419);
nor U7521 (N_7521,N_7456,N_7468);
nor U7522 (N_7522,N_7438,N_7411);
nand U7523 (N_7523,N_7427,N_7454);
and U7524 (N_7524,N_7403,N_7496);
nor U7525 (N_7525,N_7448,N_7489);
or U7526 (N_7526,N_7437,N_7407);
and U7527 (N_7527,N_7404,N_7401);
nor U7528 (N_7528,N_7453,N_7480);
and U7529 (N_7529,N_7466,N_7428);
nand U7530 (N_7530,N_7460,N_7429);
or U7531 (N_7531,N_7443,N_7420);
or U7532 (N_7532,N_7441,N_7436);
and U7533 (N_7533,N_7444,N_7459);
and U7534 (N_7534,N_7490,N_7439);
or U7535 (N_7535,N_7421,N_7471);
or U7536 (N_7536,N_7463,N_7425);
nor U7537 (N_7537,N_7426,N_7472);
and U7538 (N_7538,N_7445,N_7424);
nand U7539 (N_7539,N_7409,N_7412);
nor U7540 (N_7540,N_7470,N_7433);
nand U7541 (N_7541,N_7474,N_7482);
nor U7542 (N_7542,N_7405,N_7442);
nor U7543 (N_7543,N_7475,N_7410);
nand U7544 (N_7544,N_7494,N_7497);
nand U7545 (N_7545,N_7432,N_7457);
nor U7546 (N_7546,N_7485,N_7400);
nand U7547 (N_7547,N_7431,N_7430);
and U7548 (N_7548,N_7451,N_7476);
or U7549 (N_7549,N_7413,N_7479);
nor U7550 (N_7550,N_7471,N_7404);
nor U7551 (N_7551,N_7425,N_7448);
and U7552 (N_7552,N_7419,N_7401);
nor U7553 (N_7553,N_7431,N_7475);
and U7554 (N_7554,N_7437,N_7478);
nor U7555 (N_7555,N_7460,N_7428);
or U7556 (N_7556,N_7465,N_7439);
nor U7557 (N_7557,N_7484,N_7400);
nand U7558 (N_7558,N_7460,N_7445);
or U7559 (N_7559,N_7493,N_7453);
nor U7560 (N_7560,N_7404,N_7403);
and U7561 (N_7561,N_7463,N_7412);
nor U7562 (N_7562,N_7442,N_7486);
and U7563 (N_7563,N_7410,N_7418);
and U7564 (N_7564,N_7421,N_7425);
or U7565 (N_7565,N_7426,N_7497);
and U7566 (N_7566,N_7448,N_7463);
or U7567 (N_7567,N_7482,N_7498);
nor U7568 (N_7568,N_7432,N_7428);
nor U7569 (N_7569,N_7487,N_7427);
nand U7570 (N_7570,N_7435,N_7425);
or U7571 (N_7571,N_7405,N_7466);
and U7572 (N_7572,N_7413,N_7483);
nor U7573 (N_7573,N_7488,N_7460);
or U7574 (N_7574,N_7442,N_7448);
and U7575 (N_7575,N_7459,N_7407);
nand U7576 (N_7576,N_7434,N_7479);
nor U7577 (N_7577,N_7479,N_7446);
nand U7578 (N_7578,N_7421,N_7495);
or U7579 (N_7579,N_7460,N_7478);
xnor U7580 (N_7580,N_7453,N_7470);
nor U7581 (N_7581,N_7499,N_7408);
nand U7582 (N_7582,N_7413,N_7404);
nor U7583 (N_7583,N_7459,N_7464);
nand U7584 (N_7584,N_7481,N_7459);
nand U7585 (N_7585,N_7445,N_7450);
and U7586 (N_7586,N_7496,N_7400);
nand U7587 (N_7587,N_7414,N_7481);
nand U7588 (N_7588,N_7426,N_7489);
or U7589 (N_7589,N_7404,N_7408);
nor U7590 (N_7590,N_7443,N_7495);
nand U7591 (N_7591,N_7436,N_7489);
nand U7592 (N_7592,N_7470,N_7437);
nand U7593 (N_7593,N_7419,N_7405);
or U7594 (N_7594,N_7475,N_7423);
nand U7595 (N_7595,N_7412,N_7426);
nand U7596 (N_7596,N_7435,N_7493);
nand U7597 (N_7597,N_7447,N_7429);
nand U7598 (N_7598,N_7497,N_7408);
and U7599 (N_7599,N_7446,N_7495);
and U7600 (N_7600,N_7594,N_7508);
and U7601 (N_7601,N_7579,N_7539);
nor U7602 (N_7602,N_7564,N_7575);
or U7603 (N_7603,N_7515,N_7514);
nand U7604 (N_7604,N_7561,N_7519);
nor U7605 (N_7605,N_7590,N_7517);
or U7606 (N_7606,N_7563,N_7562);
nor U7607 (N_7607,N_7500,N_7531);
or U7608 (N_7608,N_7584,N_7526);
nor U7609 (N_7609,N_7552,N_7581);
nand U7610 (N_7610,N_7521,N_7559);
nor U7611 (N_7611,N_7553,N_7572);
and U7612 (N_7612,N_7598,N_7542);
and U7613 (N_7613,N_7556,N_7545);
nand U7614 (N_7614,N_7554,N_7568);
nand U7615 (N_7615,N_7523,N_7593);
or U7616 (N_7616,N_7533,N_7548);
nand U7617 (N_7617,N_7520,N_7546);
and U7618 (N_7618,N_7527,N_7507);
nand U7619 (N_7619,N_7510,N_7576);
and U7620 (N_7620,N_7511,N_7516);
or U7621 (N_7621,N_7530,N_7528);
nand U7622 (N_7622,N_7583,N_7540);
or U7623 (N_7623,N_7504,N_7578);
or U7624 (N_7624,N_7587,N_7558);
and U7625 (N_7625,N_7509,N_7595);
nor U7626 (N_7626,N_7565,N_7524);
nor U7627 (N_7627,N_7535,N_7522);
or U7628 (N_7628,N_7544,N_7574);
nand U7629 (N_7629,N_7543,N_7569);
and U7630 (N_7630,N_7577,N_7525);
nand U7631 (N_7631,N_7597,N_7555);
and U7632 (N_7632,N_7585,N_7529);
nor U7633 (N_7633,N_7518,N_7502);
nor U7634 (N_7634,N_7534,N_7506);
or U7635 (N_7635,N_7541,N_7582);
nor U7636 (N_7636,N_7580,N_7503);
or U7637 (N_7637,N_7513,N_7596);
nor U7638 (N_7638,N_7588,N_7550);
and U7639 (N_7639,N_7566,N_7573);
or U7640 (N_7640,N_7589,N_7549);
nand U7641 (N_7641,N_7512,N_7557);
nor U7642 (N_7642,N_7586,N_7571);
and U7643 (N_7643,N_7532,N_7560);
nand U7644 (N_7644,N_7592,N_7547);
and U7645 (N_7645,N_7505,N_7536);
nand U7646 (N_7646,N_7570,N_7537);
nand U7647 (N_7647,N_7551,N_7591);
and U7648 (N_7648,N_7538,N_7567);
nand U7649 (N_7649,N_7501,N_7599);
nor U7650 (N_7650,N_7563,N_7504);
or U7651 (N_7651,N_7582,N_7513);
and U7652 (N_7652,N_7551,N_7581);
or U7653 (N_7653,N_7568,N_7500);
and U7654 (N_7654,N_7581,N_7516);
or U7655 (N_7655,N_7571,N_7526);
and U7656 (N_7656,N_7594,N_7501);
or U7657 (N_7657,N_7524,N_7525);
or U7658 (N_7658,N_7513,N_7573);
nand U7659 (N_7659,N_7599,N_7575);
and U7660 (N_7660,N_7548,N_7507);
nor U7661 (N_7661,N_7587,N_7507);
nand U7662 (N_7662,N_7580,N_7519);
nor U7663 (N_7663,N_7568,N_7587);
or U7664 (N_7664,N_7547,N_7570);
nor U7665 (N_7665,N_7594,N_7587);
and U7666 (N_7666,N_7595,N_7573);
nor U7667 (N_7667,N_7546,N_7593);
nand U7668 (N_7668,N_7503,N_7502);
nor U7669 (N_7669,N_7515,N_7580);
nor U7670 (N_7670,N_7588,N_7571);
nand U7671 (N_7671,N_7504,N_7555);
and U7672 (N_7672,N_7539,N_7507);
or U7673 (N_7673,N_7518,N_7596);
and U7674 (N_7674,N_7576,N_7599);
and U7675 (N_7675,N_7501,N_7534);
and U7676 (N_7676,N_7502,N_7572);
or U7677 (N_7677,N_7511,N_7539);
nand U7678 (N_7678,N_7518,N_7555);
nand U7679 (N_7679,N_7517,N_7500);
nor U7680 (N_7680,N_7571,N_7590);
nor U7681 (N_7681,N_7505,N_7506);
or U7682 (N_7682,N_7567,N_7507);
or U7683 (N_7683,N_7531,N_7529);
or U7684 (N_7684,N_7519,N_7593);
nor U7685 (N_7685,N_7558,N_7506);
nand U7686 (N_7686,N_7519,N_7540);
and U7687 (N_7687,N_7527,N_7509);
or U7688 (N_7688,N_7519,N_7528);
or U7689 (N_7689,N_7556,N_7566);
and U7690 (N_7690,N_7521,N_7590);
nor U7691 (N_7691,N_7540,N_7553);
and U7692 (N_7692,N_7520,N_7581);
nor U7693 (N_7693,N_7501,N_7518);
nand U7694 (N_7694,N_7510,N_7526);
and U7695 (N_7695,N_7504,N_7582);
and U7696 (N_7696,N_7505,N_7568);
and U7697 (N_7697,N_7540,N_7597);
and U7698 (N_7698,N_7546,N_7584);
nor U7699 (N_7699,N_7531,N_7563);
nor U7700 (N_7700,N_7610,N_7695);
or U7701 (N_7701,N_7602,N_7697);
and U7702 (N_7702,N_7687,N_7689);
or U7703 (N_7703,N_7617,N_7693);
nand U7704 (N_7704,N_7682,N_7678);
and U7705 (N_7705,N_7686,N_7612);
nand U7706 (N_7706,N_7603,N_7611);
nand U7707 (N_7707,N_7609,N_7677);
nand U7708 (N_7708,N_7636,N_7663);
nand U7709 (N_7709,N_7614,N_7645);
or U7710 (N_7710,N_7681,N_7608);
or U7711 (N_7711,N_7616,N_7641);
or U7712 (N_7712,N_7692,N_7667);
or U7713 (N_7713,N_7623,N_7696);
nor U7714 (N_7714,N_7655,N_7634);
or U7715 (N_7715,N_7675,N_7654);
or U7716 (N_7716,N_7633,N_7604);
or U7717 (N_7717,N_7606,N_7652);
and U7718 (N_7718,N_7651,N_7683);
nand U7719 (N_7719,N_7621,N_7618);
or U7720 (N_7720,N_7662,N_7622);
and U7721 (N_7721,N_7660,N_7601);
and U7722 (N_7722,N_7679,N_7605);
xor U7723 (N_7723,N_7628,N_7632);
nor U7724 (N_7724,N_7640,N_7672);
nand U7725 (N_7725,N_7698,N_7669);
nor U7726 (N_7726,N_7690,N_7657);
xnor U7727 (N_7727,N_7627,N_7664);
and U7728 (N_7728,N_7650,N_7649);
and U7729 (N_7729,N_7648,N_7613);
nor U7730 (N_7730,N_7688,N_7631);
nand U7731 (N_7731,N_7624,N_7626);
nand U7732 (N_7732,N_7638,N_7625);
nor U7733 (N_7733,N_7684,N_7630);
nand U7734 (N_7734,N_7685,N_7680);
and U7735 (N_7735,N_7629,N_7619);
and U7736 (N_7736,N_7661,N_7668);
nor U7737 (N_7737,N_7670,N_7620);
and U7738 (N_7738,N_7666,N_7658);
or U7739 (N_7739,N_7646,N_7607);
or U7740 (N_7740,N_7656,N_7659);
or U7741 (N_7741,N_7637,N_7644);
and U7742 (N_7742,N_7674,N_7600);
nor U7743 (N_7743,N_7653,N_7615);
and U7744 (N_7744,N_7673,N_7691);
nor U7745 (N_7745,N_7671,N_7665);
nand U7746 (N_7746,N_7676,N_7694);
or U7747 (N_7747,N_7635,N_7639);
or U7748 (N_7748,N_7699,N_7643);
nand U7749 (N_7749,N_7647,N_7642);
or U7750 (N_7750,N_7697,N_7672);
nand U7751 (N_7751,N_7664,N_7657);
and U7752 (N_7752,N_7611,N_7608);
or U7753 (N_7753,N_7673,N_7694);
nand U7754 (N_7754,N_7695,N_7612);
or U7755 (N_7755,N_7624,N_7687);
nand U7756 (N_7756,N_7641,N_7696);
nor U7757 (N_7757,N_7679,N_7671);
and U7758 (N_7758,N_7654,N_7656);
and U7759 (N_7759,N_7627,N_7613);
or U7760 (N_7760,N_7644,N_7674);
nand U7761 (N_7761,N_7687,N_7695);
or U7762 (N_7762,N_7625,N_7679);
nor U7763 (N_7763,N_7631,N_7641);
nor U7764 (N_7764,N_7669,N_7687);
xor U7765 (N_7765,N_7628,N_7671);
nor U7766 (N_7766,N_7644,N_7602);
or U7767 (N_7767,N_7649,N_7661);
and U7768 (N_7768,N_7648,N_7629);
nand U7769 (N_7769,N_7645,N_7654);
nand U7770 (N_7770,N_7694,N_7695);
nand U7771 (N_7771,N_7624,N_7676);
and U7772 (N_7772,N_7699,N_7637);
and U7773 (N_7773,N_7644,N_7617);
or U7774 (N_7774,N_7684,N_7600);
nand U7775 (N_7775,N_7661,N_7697);
and U7776 (N_7776,N_7646,N_7625);
nor U7777 (N_7777,N_7683,N_7629);
nor U7778 (N_7778,N_7625,N_7630);
and U7779 (N_7779,N_7654,N_7613);
and U7780 (N_7780,N_7602,N_7607);
nor U7781 (N_7781,N_7617,N_7670);
nor U7782 (N_7782,N_7607,N_7637);
or U7783 (N_7783,N_7638,N_7664);
nor U7784 (N_7784,N_7683,N_7678);
and U7785 (N_7785,N_7615,N_7648);
and U7786 (N_7786,N_7647,N_7686);
and U7787 (N_7787,N_7601,N_7650);
or U7788 (N_7788,N_7629,N_7600);
nor U7789 (N_7789,N_7669,N_7674);
nand U7790 (N_7790,N_7676,N_7699);
or U7791 (N_7791,N_7608,N_7615);
and U7792 (N_7792,N_7649,N_7691);
nand U7793 (N_7793,N_7653,N_7674);
nand U7794 (N_7794,N_7683,N_7620);
nand U7795 (N_7795,N_7620,N_7692);
nand U7796 (N_7796,N_7646,N_7638);
nor U7797 (N_7797,N_7642,N_7620);
and U7798 (N_7798,N_7653,N_7652);
nor U7799 (N_7799,N_7684,N_7699);
nand U7800 (N_7800,N_7716,N_7763);
xor U7801 (N_7801,N_7758,N_7742);
nor U7802 (N_7802,N_7796,N_7726);
or U7803 (N_7803,N_7732,N_7770);
and U7804 (N_7804,N_7745,N_7705);
and U7805 (N_7805,N_7783,N_7768);
and U7806 (N_7806,N_7712,N_7746);
nand U7807 (N_7807,N_7749,N_7722);
nand U7808 (N_7808,N_7702,N_7755);
or U7809 (N_7809,N_7789,N_7795);
and U7810 (N_7810,N_7747,N_7711);
nor U7811 (N_7811,N_7757,N_7773);
nand U7812 (N_7812,N_7764,N_7703);
xor U7813 (N_7813,N_7734,N_7786);
or U7814 (N_7814,N_7774,N_7767);
and U7815 (N_7815,N_7794,N_7718);
and U7816 (N_7816,N_7790,N_7724);
and U7817 (N_7817,N_7765,N_7762);
and U7818 (N_7818,N_7710,N_7756);
nand U7819 (N_7819,N_7776,N_7717);
and U7820 (N_7820,N_7743,N_7738);
nor U7821 (N_7821,N_7727,N_7701);
and U7822 (N_7822,N_7769,N_7736);
nor U7823 (N_7823,N_7708,N_7787);
or U7824 (N_7824,N_7772,N_7784);
and U7825 (N_7825,N_7761,N_7771);
and U7826 (N_7826,N_7704,N_7791);
xnor U7827 (N_7827,N_7754,N_7728);
or U7828 (N_7828,N_7700,N_7797);
nor U7829 (N_7829,N_7719,N_7750);
nor U7830 (N_7830,N_7729,N_7782);
or U7831 (N_7831,N_7741,N_7735);
or U7832 (N_7832,N_7744,N_7709);
nor U7833 (N_7833,N_7779,N_7793);
nor U7834 (N_7834,N_7751,N_7778);
nand U7835 (N_7835,N_7766,N_7731);
nand U7836 (N_7836,N_7781,N_7799);
nor U7837 (N_7837,N_7733,N_7739);
or U7838 (N_7838,N_7753,N_7785);
nand U7839 (N_7839,N_7798,N_7713);
and U7840 (N_7840,N_7707,N_7760);
and U7841 (N_7841,N_7721,N_7788);
xor U7842 (N_7842,N_7720,N_7706);
or U7843 (N_7843,N_7715,N_7723);
nor U7844 (N_7844,N_7792,N_7748);
and U7845 (N_7845,N_7775,N_7759);
or U7846 (N_7846,N_7740,N_7752);
nor U7847 (N_7847,N_7714,N_7780);
nor U7848 (N_7848,N_7730,N_7777);
nor U7849 (N_7849,N_7725,N_7737);
nor U7850 (N_7850,N_7769,N_7797);
or U7851 (N_7851,N_7722,N_7755);
or U7852 (N_7852,N_7721,N_7727);
nor U7853 (N_7853,N_7774,N_7788);
xor U7854 (N_7854,N_7737,N_7715);
nand U7855 (N_7855,N_7775,N_7779);
or U7856 (N_7856,N_7784,N_7753);
and U7857 (N_7857,N_7726,N_7731);
or U7858 (N_7858,N_7753,N_7714);
nor U7859 (N_7859,N_7736,N_7743);
or U7860 (N_7860,N_7777,N_7766);
and U7861 (N_7861,N_7739,N_7750);
nand U7862 (N_7862,N_7717,N_7747);
nand U7863 (N_7863,N_7722,N_7770);
nor U7864 (N_7864,N_7709,N_7767);
nor U7865 (N_7865,N_7744,N_7797);
and U7866 (N_7866,N_7750,N_7778);
and U7867 (N_7867,N_7704,N_7731);
nor U7868 (N_7868,N_7768,N_7729);
and U7869 (N_7869,N_7730,N_7745);
or U7870 (N_7870,N_7773,N_7717);
nor U7871 (N_7871,N_7705,N_7746);
and U7872 (N_7872,N_7785,N_7762);
nor U7873 (N_7873,N_7789,N_7753);
nand U7874 (N_7874,N_7705,N_7708);
or U7875 (N_7875,N_7715,N_7714);
and U7876 (N_7876,N_7773,N_7783);
nor U7877 (N_7877,N_7788,N_7771);
nor U7878 (N_7878,N_7787,N_7715);
and U7879 (N_7879,N_7754,N_7770);
nor U7880 (N_7880,N_7715,N_7790);
nand U7881 (N_7881,N_7770,N_7775);
or U7882 (N_7882,N_7731,N_7756);
nor U7883 (N_7883,N_7774,N_7796);
nand U7884 (N_7884,N_7750,N_7751);
and U7885 (N_7885,N_7764,N_7774);
or U7886 (N_7886,N_7701,N_7779);
or U7887 (N_7887,N_7777,N_7718);
nor U7888 (N_7888,N_7717,N_7771);
nand U7889 (N_7889,N_7712,N_7766);
nor U7890 (N_7890,N_7759,N_7778);
nand U7891 (N_7891,N_7750,N_7715);
or U7892 (N_7892,N_7727,N_7790);
nor U7893 (N_7893,N_7754,N_7718);
nand U7894 (N_7894,N_7751,N_7743);
or U7895 (N_7895,N_7757,N_7703);
or U7896 (N_7896,N_7729,N_7764);
or U7897 (N_7897,N_7729,N_7777);
nand U7898 (N_7898,N_7735,N_7732);
and U7899 (N_7899,N_7777,N_7721);
or U7900 (N_7900,N_7859,N_7805);
and U7901 (N_7901,N_7876,N_7880);
nor U7902 (N_7902,N_7841,N_7827);
or U7903 (N_7903,N_7896,N_7844);
or U7904 (N_7904,N_7855,N_7838);
and U7905 (N_7905,N_7810,N_7825);
or U7906 (N_7906,N_7868,N_7821);
and U7907 (N_7907,N_7804,N_7817);
and U7908 (N_7908,N_7815,N_7871);
nand U7909 (N_7909,N_7801,N_7853);
or U7910 (N_7910,N_7864,N_7829);
or U7911 (N_7911,N_7856,N_7802);
nand U7912 (N_7912,N_7832,N_7834);
and U7913 (N_7913,N_7851,N_7800);
or U7914 (N_7914,N_7807,N_7837);
nor U7915 (N_7915,N_7893,N_7885);
nand U7916 (N_7916,N_7803,N_7886);
and U7917 (N_7917,N_7877,N_7823);
nand U7918 (N_7918,N_7883,N_7862);
nor U7919 (N_7919,N_7884,N_7852);
nor U7920 (N_7920,N_7891,N_7846);
and U7921 (N_7921,N_7820,N_7809);
and U7922 (N_7922,N_7869,N_7808);
and U7923 (N_7923,N_7889,N_7857);
or U7924 (N_7924,N_7835,N_7861);
nor U7925 (N_7925,N_7858,N_7887);
or U7926 (N_7926,N_7845,N_7870);
nor U7927 (N_7927,N_7847,N_7867);
and U7928 (N_7928,N_7872,N_7874);
or U7929 (N_7929,N_7848,N_7850);
nor U7930 (N_7930,N_7866,N_7881);
or U7931 (N_7931,N_7890,N_7819);
nand U7932 (N_7932,N_7894,N_7863);
and U7933 (N_7933,N_7882,N_7826);
nand U7934 (N_7934,N_7836,N_7831);
nor U7935 (N_7935,N_7833,N_7895);
or U7936 (N_7936,N_7878,N_7811);
nand U7937 (N_7937,N_7843,N_7818);
or U7938 (N_7938,N_7824,N_7860);
and U7939 (N_7939,N_7813,N_7830);
nor U7940 (N_7940,N_7875,N_7840);
nor U7941 (N_7941,N_7849,N_7828);
nand U7942 (N_7942,N_7839,N_7816);
or U7943 (N_7943,N_7897,N_7806);
and U7944 (N_7944,N_7892,N_7812);
or U7945 (N_7945,N_7814,N_7865);
and U7946 (N_7946,N_7873,N_7842);
nor U7947 (N_7947,N_7879,N_7888);
nor U7948 (N_7948,N_7898,N_7899);
and U7949 (N_7949,N_7822,N_7854);
or U7950 (N_7950,N_7816,N_7807);
xor U7951 (N_7951,N_7800,N_7876);
nand U7952 (N_7952,N_7825,N_7814);
and U7953 (N_7953,N_7838,N_7885);
or U7954 (N_7954,N_7855,N_7875);
or U7955 (N_7955,N_7873,N_7894);
and U7956 (N_7956,N_7861,N_7866);
or U7957 (N_7957,N_7892,N_7863);
nand U7958 (N_7958,N_7864,N_7812);
nor U7959 (N_7959,N_7881,N_7836);
nor U7960 (N_7960,N_7847,N_7834);
and U7961 (N_7961,N_7875,N_7878);
or U7962 (N_7962,N_7876,N_7867);
and U7963 (N_7963,N_7847,N_7895);
nand U7964 (N_7964,N_7829,N_7866);
and U7965 (N_7965,N_7821,N_7871);
or U7966 (N_7966,N_7848,N_7871);
nand U7967 (N_7967,N_7819,N_7824);
nand U7968 (N_7968,N_7881,N_7826);
nor U7969 (N_7969,N_7829,N_7811);
or U7970 (N_7970,N_7859,N_7887);
nor U7971 (N_7971,N_7881,N_7890);
nor U7972 (N_7972,N_7869,N_7894);
nand U7973 (N_7973,N_7839,N_7896);
or U7974 (N_7974,N_7819,N_7860);
or U7975 (N_7975,N_7809,N_7835);
and U7976 (N_7976,N_7825,N_7841);
nor U7977 (N_7977,N_7835,N_7810);
or U7978 (N_7978,N_7865,N_7831);
and U7979 (N_7979,N_7868,N_7846);
or U7980 (N_7980,N_7855,N_7879);
and U7981 (N_7981,N_7848,N_7804);
nor U7982 (N_7982,N_7867,N_7836);
and U7983 (N_7983,N_7806,N_7888);
nand U7984 (N_7984,N_7803,N_7883);
nor U7985 (N_7985,N_7832,N_7804);
nand U7986 (N_7986,N_7880,N_7842);
and U7987 (N_7987,N_7839,N_7892);
nor U7988 (N_7988,N_7802,N_7850);
nor U7989 (N_7989,N_7807,N_7888);
and U7990 (N_7990,N_7859,N_7893);
and U7991 (N_7991,N_7883,N_7841);
nor U7992 (N_7992,N_7869,N_7835);
nor U7993 (N_7993,N_7861,N_7893);
nand U7994 (N_7994,N_7873,N_7828);
nor U7995 (N_7995,N_7892,N_7811);
or U7996 (N_7996,N_7851,N_7812);
and U7997 (N_7997,N_7839,N_7864);
xor U7998 (N_7998,N_7821,N_7893);
and U7999 (N_7999,N_7813,N_7866);
nand U8000 (N_8000,N_7972,N_7978);
nor U8001 (N_8001,N_7953,N_7979);
nor U8002 (N_8002,N_7930,N_7989);
nand U8003 (N_8003,N_7915,N_7961);
or U8004 (N_8004,N_7909,N_7906);
or U8005 (N_8005,N_7981,N_7903);
nor U8006 (N_8006,N_7913,N_7947);
nand U8007 (N_8007,N_7971,N_7982);
and U8008 (N_8008,N_7988,N_7960);
and U8009 (N_8009,N_7998,N_7991);
or U8010 (N_8010,N_7924,N_7937);
nor U8011 (N_8011,N_7922,N_7984);
nand U8012 (N_8012,N_7928,N_7992);
nor U8013 (N_8013,N_7911,N_7945);
nand U8014 (N_8014,N_7902,N_7963);
nor U8015 (N_8015,N_7934,N_7997);
xor U8016 (N_8016,N_7976,N_7951);
or U8017 (N_8017,N_7942,N_7949);
nor U8018 (N_8018,N_7970,N_7983);
nand U8019 (N_8019,N_7962,N_7940);
and U8020 (N_8020,N_7996,N_7939);
nor U8021 (N_8021,N_7926,N_7904);
or U8022 (N_8022,N_7966,N_7944);
nor U8023 (N_8023,N_7935,N_7946);
nor U8024 (N_8024,N_7936,N_7994);
nor U8025 (N_8025,N_7927,N_7931);
or U8026 (N_8026,N_7932,N_7973);
and U8027 (N_8027,N_7938,N_7987);
nor U8028 (N_8028,N_7923,N_7977);
or U8029 (N_8029,N_7954,N_7965);
or U8030 (N_8030,N_7918,N_7990);
nor U8031 (N_8031,N_7920,N_7993);
or U8032 (N_8032,N_7916,N_7986);
nand U8033 (N_8033,N_7907,N_7955);
nand U8034 (N_8034,N_7925,N_7958);
nor U8035 (N_8035,N_7999,N_7967);
nor U8036 (N_8036,N_7912,N_7952);
nand U8037 (N_8037,N_7948,N_7969);
or U8038 (N_8038,N_7964,N_7943);
and U8039 (N_8039,N_7933,N_7985);
nand U8040 (N_8040,N_7950,N_7908);
nand U8041 (N_8041,N_7975,N_7910);
or U8042 (N_8042,N_7905,N_7917);
and U8043 (N_8043,N_7929,N_7900);
nor U8044 (N_8044,N_7921,N_7995);
and U8045 (N_8045,N_7941,N_7914);
nor U8046 (N_8046,N_7974,N_7919);
and U8047 (N_8047,N_7980,N_7959);
and U8048 (N_8048,N_7901,N_7968);
nand U8049 (N_8049,N_7957,N_7956);
nand U8050 (N_8050,N_7949,N_7914);
and U8051 (N_8051,N_7901,N_7954);
nor U8052 (N_8052,N_7979,N_7901);
nor U8053 (N_8053,N_7964,N_7925);
or U8054 (N_8054,N_7994,N_7915);
nand U8055 (N_8055,N_7984,N_7928);
or U8056 (N_8056,N_7903,N_7936);
nor U8057 (N_8057,N_7924,N_7915);
nor U8058 (N_8058,N_7958,N_7972);
and U8059 (N_8059,N_7969,N_7992);
nand U8060 (N_8060,N_7979,N_7909);
nand U8061 (N_8061,N_7989,N_7927);
or U8062 (N_8062,N_7926,N_7900);
or U8063 (N_8063,N_7925,N_7977);
or U8064 (N_8064,N_7945,N_7971);
and U8065 (N_8065,N_7963,N_7997);
and U8066 (N_8066,N_7984,N_7906);
nor U8067 (N_8067,N_7902,N_7933);
nand U8068 (N_8068,N_7945,N_7922);
nand U8069 (N_8069,N_7962,N_7924);
nand U8070 (N_8070,N_7934,N_7963);
and U8071 (N_8071,N_7926,N_7912);
and U8072 (N_8072,N_7939,N_7927);
and U8073 (N_8073,N_7977,N_7965);
and U8074 (N_8074,N_7903,N_7919);
or U8075 (N_8075,N_7919,N_7965);
nand U8076 (N_8076,N_7927,N_7901);
and U8077 (N_8077,N_7910,N_7962);
nor U8078 (N_8078,N_7901,N_7931);
nand U8079 (N_8079,N_7974,N_7921);
nor U8080 (N_8080,N_7991,N_7934);
nand U8081 (N_8081,N_7917,N_7910);
and U8082 (N_8082,N_7941,N_7917);
nand U8083 (N_8083,N_7953,N_7903);
nand U8084 (N_8084,N_7980,N_7965);
or U8085 (N_8085,N_7973,N_7924);
xnor U8086 (N_8086,N_7931,N_7999);
and U8087 (N_8087,N_7943,N_7945);
nand U8088 (N_8088,N_7949,N_7993);
nor U8089 (N_8089,N_7970,N_7984);
nand U8090 (N_8090,N_7996,N_7983);
or U8091 (N_8091,N_7951,N_7905);
nand U8092 (N_8092,N_7948,N_7953);
or U8093 (N_8093,N_7933,N_7963);
nand U8094 (N_8094,N_7975,N_7972);
and U8095 (N_8095,N_7900,N_7976);
nand U8096 (N_8096,N_7906,N_7952);
and U8097 (N_8097,N_7930,N_7994);
and U8098 (N_8098,N_7995,N_7981);
and U8099 (N_8099,N_7905,N_7960);
nor U8100 (N_8100,N_8049,N_8031);
nor U8101 (N_8101,N_8024,N_8006);
or U8102 (N_8102,N_8016,N_8088);
and U8103 (N_8103,N_8052,N_8033);
nor U8104 (N_8104,N_8067,N_8023);
or U8105 (N_8105,N_8096,N_8090);
or U8106 (N_8106,N_8004,N_8097);
nand U8107 (N_8107,N_8072,N_8061);
nor U8108 (N_8108,N_8065,N_8009);
nand U8109 (N_8109,N_8038,N_8080);
nor U8110 (N_8110,N_8000,N_8058);
or U8111 (N_8111,N_8047,N_8078);
and U8112 (N_8112,N_8050,N_8099);
nand U8113 (N_8113,N_8055,N_8010);
nor U8114 (N_8114,N_8071,N_8045);
and U8115 (N_8115,N_8054,N_8070);
or U8116 (N_8116,N_8076,N_8056);
nor U8117 (N_8117,N_8069,N_8001);
nand U8118 (N_8118,N_8011,N_8034);
nand U8119 (N_8119,N_8064,N_8003);
or U8120 (N_8120,N_8017,N_8085);
or U8121 (N_8121,N_8093,N_8020);
nor U8122 (N_8122,N_8028,N_8087);
and U8123 (N_8123,N_8013,N_8012);
nor U8124 (N_8124,N_8027,N_8044);
nand U8125 (N_8125,N_8007,N_8059);
or U8126 (N_8126,N_8095,N_8066);
nand U8127 (N_8127,N_8025,N_8068);
or U8128 (N_8128,N_8086,N_8029);
nor U8129 (N_8129,N_8039,N_8015);
nand U8130 (N_8130,N_8002,N_8032);
and U8131 (N_8131,N_8060,N_8021);
nand U8132 (N_8132,N_8043,N_8075);
and U8133 (N_8133,N_8040,N_8098);
nand U8134 (N_8134,N_8082,N_8037);
or U8135 (N_8135,N_8094,N_8077);
nor U8136 (N_8136,N_8091,N_8092);
and U8137 (N_8137,N_8074,N_8051);
or U8138 (N_8138,N_8062,N_8008);
and U8139 (N_8139,N_8026,N_8079);
or U8140 (N_8140,N_8081,N_8041);
nand U8141 (N_8141,N_8030,N_8042);
or U8142 (N_8142,N_8035,N_8019);
and U8143 (N_8143,N_8018,N_8036);
nor U8144 (N_8144,N_8089,N_8073);
and U8145 (N_8145,N_8022,N_8005);
nand U8146 (N_8146,N_8063,N_8083);
or U8147 (N_8147,N_8057,N_8048);
nor U8148 (N_8148,N_8014,N_8084);
nor U8149 (N_8149,N_8053,N_8046);
and U8150 (N_8150,N_8076,N_8083);
and U8151 (N_8151,N_8052,N_8056);
nand U8152 (N_8152,N_8096,N_8074);
nand U8153 (N_8153,N_8082,N_8025);
or U8154 (N_8154,N_8058,N_8054);
nand U8155 (N_8155,N_8088,N_8028);
nor U8156 (N_8156,N_8043,N_8008);
nand U8157 (N_8157,N_8030,N_8033);
or U8158 (N_8158,N_8007,N_8084);
or U8159 (N_8159,N_8012,N_8008);
or U8160 (N_8160,N_8059,N_8069);
nand U8161 (N_8161,N_8051,N_8042);
and U8162 (N_8162,N_8099,N_8021);
or U8163 (N_8163,N_8004,N_8031);
nand U8164 (N_8164,N_8005,N_8020);
or U8165 (N_8165,N_8081,N_8087);
or U8166 (N_8166,N_8068,N_8070);
or U8167 (N_8167,N_8045,N_8040);
and U8168 (N_8168,N_8096,N_8030);
and U8169 (N_8169,N_8086,N_8022);
nand U8170 (N_8170,N_8023,N_8016);
or U8171 (N_8171,N_8002,N_8089);
nor U8172 (N_8172,N_8042,N_8016);
nor U8173 (N_8173,N_8012,N_8089);
or U8174 (N_8174,N_8084,N_8058);
nor U8175 (N_8175,N_8036,N_8015);
or U8176 (N_8176,N_8085,N_8009);
and U8177 (N_8177,N_8066,N_8052);
nor U8178 (N_8178,N_8076,N_8007);
nor U8179 (N_8179,N_8054,N_8039);
and U8180 (N_8180,N_8008,N_8058);
nand U8181 (N_8181,N_8045,N_8095);
nand U8182 (N_8182,N_8049,N_8024);
nand U8183 (N_8183,N_8004,N_8089);
and U8184 (N_8184,N_8035,N_8071);
xnor U8185 (N_8185,N_8081,N_8061);
or U8186 (N_8186,N_8046,N_8076);
nor U8187 (N_8187,N_8030,N_8059);
nor U8188 (N_8188,N_8093,N_8092);
and U8189 (N_8189,N_8017,N_8041);
and U8190 (N_8190,N_8056,N_8028);
or U8191 (N_8191,N_8039,N_8027);
nor U8192 (N_8192,N_8012,N_8059);
nand U8193 (N_8193,N_8066,N_8094);
and U8194 (N_8194,N_8064,N_8097);
nor U8195 (N_8195,N_8033,N_8074);
nor U8196 (N_8196,N_8037,N_8094);
nand U8197 (N_8197,N_8059,N_8046);
and U8198 (N_8198,N_8076,N_8089);
nand U8199 (N_8199,N_8026,N_8063);
nor U8200 (N_8200,N_8102,N_8135);
and U8201 (N_8201,N_8186,N_8150);
nor U8202 (N_8202,N_8163,N_8119);
nor U8203 (N_8203,N_8155,N_8158);
or U8204 (N_8204,N_8118,N_8159);
or U8205 (N_8205,N_8107,N_8157);
and U8206 (N_8206,N_8162,N_8197);
or U8207 (N_8207,N_8183,N_8106);
and U8208 (N_8208,N_8109,N_8152);
and U8209 (N_8209,N_8101,N_8112);
nand U8210 (N_8210,N_8103,N_8129);
and U8211 (N_8211,N_8104,N_8156);
nor U8212 (N_8212,N_8153,N_8140);
or U8213 (N_8213,N_8169,N_8167);
or U8214 (N_8214,N_8185,N_8192);
nand U8215 (N_8215,N_8145,N_8124);
nor U8216 (N_8216,N_8164,N_8113);
or U8217 (N_8217,N_8138,N_8166);
and U8218 (N_8218,N_8126,N_8198);
and U8219 (N_8219,N_8137,N_8143);
or U8220 (N_8220,N_8184,N_8108);
nand U8221 (N_8221,N_8168,N_8146);
nand U8222 (N_8222,N_8176,N_8191);
or U8223 (N_8223,N_8195,N_8196);
nor U8224 (N_8224,N_8177,N_8100);
and U8225 (N_8225,N_8193,N_8133);
nor U8226 (N_8226,N_8160,N_8181);
nand U8227 (N_8227,N_8187,N_8139);
or U8228 (N_8228,N_8122,N_8173);
or U8229 (N_8229,N_8131,N_8171);
and U8230 (N_8230,N_8175,N_8144);
nor U8231 (N_8231,N_8174,N_8165);
nor U8232 (N_8232,N_8199,N_8142);
or U8233 (N_8233,N_8178,N_8148);
nand U8234 (N_8234,N_8130,N_8188);
nand U8235 (N_8235,N_8132,N_8179);
nand U8236 (N_8236,N_8161,N_8123);
or U8237 (N_8237,N_8125,N_8190);
nand U8238 (N_8238,N_8149,N_8147);
and U8239 (N_8239,N_8120,N_8136);
nor U8240 (N_8240,N_8105,N_8151);
nor U8241 (N_8241,N_8170,N_8182);
nor U8242 (N_8242,N_8116,N_8194);
nor U8243 (N_8243,N_8189,N_8154);
nand U8244 (N_8244,N_8114,N_8111);
or U8245 (N_8245,N_8141,N_8117);
nand U8246 (N_8246,N_8134,N_8121);
or U8247 (N_8247,N_8128,N_8180);
or U8248 (N_8248,N_8127,N_8115);
and U8249 (N_8249,N_8110,N_8172);
nand U8250 (N_8250,N_8176,N_8160);
and U8251 (N_8251,N_8186,N_8170);
or U8252 (N_8252,N_8185,N_8149);
nand U8253 (N_8253,N_8179,N_8121);
or U8254 (N_8254,N_8191,N_8182);
or U8255 (N_8255,N_8190,N_8164);
nor U8256 (N_8256,N_8107,N_8135);
and U8257 (N_8257,N_8120,N_8199);
or U8258 (N_8258,N_8127,N_8132);
nand U8259 (N_8259,N_8185,N_8151);
or U8260 (N_8260,N_8172,N_8137);
nor U8261 (N_8261,N_8151,N_8104);
nand U8262 (N_8262,N_8197,N_8158);
and U8263 (N_8263,N_8175,N_8170);
nand U8264 (N_8264,N_8130,N_8170);
nor U8265 (N_8265,N_8193,N_8102);
and U8266 (N_8266,N_8123,N_8178);
nand U8267 (N_8267,N_8138,N_8131);
nand U8268 (N_8268,N_8139,N_8133);
nor U8269 (N_8269,N_8101,N_8129);
or U8270 (N_8270,N_8195,N_8181);
nand U8271 (N_8271,N_8127,N_8109);
or U8272 (N_8272,N_8138,N_8175);
nand U8273 (N_8273,N_8199,N_8155);
or U8274 (N_8274,N_8104,N_8165);
and U8275 (N_8275,N_8199,N_8184);
nand U8276 (N_8276,N_8181,N_8169);
nor U8277 (N_8277,N_8111,N_8105);
nand U8278 (N_8278,N_8128,N_8172);
or U8279 (N_8279,N_8148,N_8158);
and U8280 (N_8280,N_8167,N_8152);
or U8281 (N_8281,N_8155,N_8197);
or U8282 (N_8282,N_8161,N_8107);
or U8283 (N_8283,N_8178,N_8101);
and U8284 (N_8284,N_8196,N_8187);
and U8285 (N_8285,N_8117,N_8136);
nand U8286 (N_8286,N_8143,N_8107);
and U8287 (N_8287,N_8125,N_8157);
or U8288 (N_8288,N_8149,N_8104);
or U8289 (N_8289,N_8174,N_8131);
nand U8290 (N_8290,N_8120,N_8164);
and U8291 (N_8291,N_8102,N_8156);
and U8292 (N_8292,N_8187,N_8164);
xor U8293 (N_8293,N_8155,N_8141);
nor U8294 (N_8294,N_8176,N_8139);
nand U8295 (N_8295,N_8167,N_8113);
nor U8296 (N_8296,N_8114,N_8182);
nor U8297 (N_8297,N_8165,N_8142);
nor U8298 (N_8298,N_8167,N_8174);
or U8299 (N_8299,N_8155,N_8145);
nor U8300 (N_8300,N_8273,N_8226);
and U8301 (N_8301,N_8231,N_8237);
or U8302 (N_8302,N_8269,N_8285);
or U8303 (N_8303,N_8239,N_8258);
nor U8304 (N_8304,N_8205,N_8241);
nor U8305 (N_8305,N_8233,N_8219);
nand U8306 (N_8306,N_8217,N_8209);
nand U8307 (N_8307,N_8281,N_8271);
and U8308 (N_8308,N_8254,N_8242);
or U8309 (N_8309,N_8287,N_8247);
nand U8310 (N_8310,N_8245,N_8223);
or U8311 (N_8311,N_8230,N_8296);
or U8312 (N_8312,N_8214,N_8275);
nand U8313 (N_8313,N_8268,N_8267);
xor U8314 (N_8314,N_8216,N_8298);
or U8315 (N_8315,N_8202,N_8284);
and U8316 (N_8316,N_8206,N_8261);
nor U8317 (N_8317,N_8204,N_8259);
nand U8318 (N_8318,N_8201,N_8256);
nor U8319 (N_8319,N_8211,N_8299);
nand U8320 (N_8320,N_8290,N_8236);
and U8321 (N_8321,N_8272,N_8224);
nand U8322 (N_8322,N_8291,N_8248);
nand U8323 (N_8323,N_8218,N_8213);
nand U8324 (N_8324,N_8215,N_8238);
or U8325 (N_8325,N_8270,N_8257);
nand U8326 (N_8326,N_8227,N_8246);
nand U8327 (N_8327,N_8278,N_8286);
or U8328 (N_8328,N_8279,N_8240);
and U8329 (N_8329,N_8282,N_8210);
nand U8330 (N_8330,N_8207,N_8274);
nor U8331 (N_8331,N_8250,N_8232);
nor U8332 (N_8332,N_8265,N_8277);
nor U8333 (N_8333,N_8292,N_8222);
nor U8334 (N_8334,N_8208,N_8244);
nor U8335 (N_8335,N_8276,N_8266);
nor U8336 (N_8336,N_8252,N_8212);
nor U8337 (N_8337,N_8203,N_8297);
and U8338 (N_8338,N_8225,N_8228);
and U8339 (N_8339,N_8283,N_8280);
nand U8340 (N_8340,N_8229,N_8235);
or U8341 (N_8341,N_8220,N_8234);
xnor U8342 (N_8342,N_8295,N_8263);
nand U8343 (N_8343,N_8288,N_8243);
and U8344 (N_8344,N_8293,N_8255);
and U8345 (N_8345,N_8251,N_8264);
nand U8346 (N_8346,N_8200,N_8289);
nand U8347 (N_8347,N_8221,N_8294);
or U8348 (N_8348,N_8249,N_8262);
and U8349 (N_8349,N_8253,N_8260);
nand U8350 (N_8350,N_8283,N_8277);
nor U8351 (N_8351,N_8242,N_8246);
and U8352 (N_8352,N_8221,N_8214);
and U8353 (N_8353,N_8224,N_8269);
nor U8354 (N_8354,N_8296,N_8298);
and U8355 (N_8355,N_8276,N_8216);
and U8356 (N_8356,N_8231,N_8275);
or U8357 (N_8357,N_8254,N_8263);
nor U8358 (N_8358,N_8264,N_8244);
nand U8359 (N_8359,N_8240,N_8259);
nor U8360 (N_8360,N_8265,N_8232);
or U8361 (N_8361,N_8219,N_8220);
nand U8362 (N_8362,N_8246,N_8231);
or U8363 (N_8363,N_8278,N_8295);
or U8364 (N_8364,N_8258,N_8282);
nor U8365 (N_8365,N_8214,N_8230);
nor U8366 (N_8366,N_8237,N_8235);
nand U8367 (N_8367,N_8222,N_8290);
and U8368 (N_8368,N_8252,N_8288);
and U8369 (N_8369,N_8217,N_8214);
nor U8370 (N_8370,N_8263,N_8244);
and U8371 (N_8371,N_8253,N_8232);
nand U8372 (N_8372,N_8211,N_8268);
or U8373 (N_8373,N_8265,N_8224);
and U8374 (N_8374,N_8240,N_8273);
nor U8375 (N_8375,N_8224,N_8251);
nand U8376 (N_8376,N_8286,N_8298);
nand U8377 (N_8377,N_8267,N_8262);
nor U8378 (N_8378,N_8204,N_8264);
nor U8379 (N_8379,N_8260,N_8265);
or U8380 (N_8380,N_8299,N_8279);
nor U8381 (N_8381,N_8297,N_8246);
and U8382 (N_8382,N_8252,N_8209);
nor U8383 (N_8383,N_8273,N_8278);
or U8384 (N_8384,N_8295,N_8248);
and U8385 (N_8385,N_8263,N_8221);
and U8386 (N_8386,N_8298,N_8269);
and U8387 (N_8387,N_8260,N_8259);
and U8388 (N_8388,N_8264,N_8206);
and U8389 (N_8389,N_8298,N_8241);
xnor U8390 (N_8390,N_8279,N_8232);
nand U8391 (N_8391,N_8284,N_8233);
and U8392 (N_8392,N_8247,N_8200);
or U8393 (N_8393,N_8227,N_8218);
and U8394 (N_8394,N_8275,N_8250);
or U8395 (N_8395,N_8266,N_8228);
or U8396 (N_8396,N_8223,N_8232);
and U8397 (N_8397,N_8276,N_8297);
or U8398 (N_8398,N_8245,N_8200);
and U8399 (N_8399,N_8270,N_8294);
or U8400 (N_8400,N_8339,N_8310);
and U8401 (N_8401,N_8362,N_8326);
and U8402 (N_8402,N_8314,N_8366);
and U8403 (N_8403,N_8341,N_8390);
or U8404 (N_8404,N_8300,N_8323);
nand U8405 (N_8405,N_8320,N_8364);
nor U8406 (N_8406,N_8351,N_8385);
nor U8407 (N_8407,N_8331,N_8306);
nor U8408 (N_8408,N_8376,N_8349);
and U8409 (N_8409,N_8361,N_8367);
and U8410 (N_8410,N_8399,N_8312);
or U8411 (N_8411,N_8379,N_8342);
nand U8412 (N_8412,N_8377,N_8384);
nand U8413 (N_8413,N_8386,N_8346);
nand U8414 (N_8414,N_8398,N_8308);
nand U8415 (N_8415,N_8389,N_8374);
or U8416 (N_8416,N_8387,N_8335);
nor U8417 (N_8417,N_8347,N_8397);
xnor U8418 (N_8418,N_8396,N_8337);
nand U8419 (N_8419,N_8345,N_8392);
nand U8420 (N_8420,N_8363,N_8378);
and U8421 (N_8421,N_8368,N_8356);
nor U8422 (N_8422,N_8358,N_8338);
and U8423 (N_8423,N_8327,N_8319);
nor U8424 (N_8424,N_8394,N_8344);
and U8425 (N_8425,N_8315,N_8330);
nor U8426 (N_8426,N_8360,N_8322);
nand U8427 (N_8427,N_8309,N_8371);
or U8428 (N_8428,N_8333,N_8381);
and U8429 (N_8429,N_8383,N_8321);
nand U8430 (N_8430,N_8304,N_8395);
or U8431 (N_8431,N_8307,N_8328);
nand U8432 (N_8432,N_8370,N_8365);
and U8433 (N_8433,N_8332,N_8353);
and U8434 (N_8434,N_8369,N_8329);
nor U8435 (N_8435,N_8372,N_8354);
nand U8436 (N_8436,N_8380,N_8334);
or U8437 (N_8437,N_8355,N_8391);
nand U8438 (N_8438,N_8302,N_8375);
nand U8439 (N_8439,N_8325,N_8316);
nand U8440 (N_8440,N_8393,N_8350);
nand U8441 (N_8441,N_8357,N_8317);
and U8442 (N_8442,N_8318,N_8336);
nand U8443 (N_8443,N_8348,N_8359);
nand U8444 (N_8444,N_8352,N_8340);
nand U8445 (N_8445,N_8388,N_8311);
and U8446 (N_8446,N_8313,N_8305);
and U8447 (N_8447,N_8324,N_8382);
nor U8448 (N_8448,N_8301,N_8373);
or U8449 (N_8449,N_8343,N_8303);
or U8450 (N_8450,N_8395,N_8331);
and U8451 (N_8451,N_8373,N_8328);
and U8452 (N_8452,N_8322,N_8306);
or U8453 (N_8453,N_8387,N_8301);
or U8454 (N_8454,N_8393,N_8398);
nor U8455 (N_8455,N_8338,N_8398);
nor U8456 (N_8456,N_8391,N_8326);
nand U8457 (N_8457,N_8347,N_8346);
and U8458 (N_8458,N_8346,N_8325);
and U8459 (N_8459,N_8335,N_8388);
nand U8460 (N_8460,N_8395,N_8366);
or U8461 (N_8461,N_8355,N_8393);
or U8462 (N_8462,N_8394,N_8361);
or U8463 (N_8463,N_8320,N_8331);
nor U8464 (N_8464,N_8362,N_8352);
or U8465 (N_8465,N_8328,N_8366);
and U8466 (N_8466,N_8335,N_8359);
or U8467 (N_8467,N_8396,N_8352);
and U8468 (N_8468,N_8339,N_8317);
or U8469 (N_8469,N_8333,N_8303);
nand U8470 (N_8470,N_8321,N_8311);
nand U8471 (N_8471,N_8351,N_8373);
nand U8472 (N_8472,N_8315,N_8380);
nor U8473 (N_8473,N_8344,N_8366);
and U8474 (N_8474,N_8391,N_8393);
nor U8475 (N_8475,N_8362,N_8396);
or U8476 (N_8476,N_8353,N_8343);
and U8477 (N_8477,N_8315,N_8336);
or U8478 (N_8478,N_8368,N_8339);
or U8479 (N_8479,N_8345,N_8368);
nand U8480 (N_8480,N_8379,N_8300);
or U8481 (N_8481,N_8350,N_8368);
nand U8482 (N_8482,N_8323,N_8319);
and U8483 (N_8483,N_8371,N_8377);
and U8484 (N_8484,N_8322,N_8340);
nor U8485 (N_8485,N_8344,N_8338);
nor U8486 (N_8486,N_8319,N_8315);
nor U8487 (N_8487,N_8344,N_8309);
or U8488 (N_8488,N_8371,N_8347);
and U8489 (N_8489,N_8398,N_8384);
or U8490 (N_8490,N_8344,N_8334);
nor U8491 (N_8491,N_8310,N_8321);
nor U8492 (N_8492,N_8381,N_8337);
or U8493 (N_8493,N_8373,N_8322);
nand U8494 (N_8494,N_8389,N_8367);
and U8495 (N_8495,N_8308,N_8386);
nor U8496 (N_8496,N_8385,N_8393);
and U8497 (N_8497,N_8316,N_8329);
and U8498 (N_8498,N_8391,N_8397);
and U8499 (N_8499,N_8307,N_8324);
or U8500 (N_8500,N_8425,N_8402);
and U8501 (N_8501,N_8405,N_8490);
nor U8502 (N_8502,N_8471,N_8420);
or U8503 (N_8503,N_8424,N_8462);
nor U8504 (N_8504,N_8457,N_8497);
nand U8505 (N_8505,N_8448,N_8427);
nand U8506 (N_8506,N_8418,N_8438);
or U8507 (N_8507,N_8439,N_8498);
nor U8508 (N_8508,N_8474,N_8466);
or U8509 (N_8509,N_8468,N_8432);
or U8510 (N_8510,N_8486,N_8461);
nor U8511 (N_8511,N_8417,N_8442);
and U8512 (N_8512,N_8499,N_8465);
nor U8513 (N_8513,N_8460,N_8437);
nor U8514 (N_8514,N_8409,N_8452);
or U8515 (N_8515,N_8400,N_8401);
nor U8516 (N_8516,N_8431,N_8426);
nor U8517 (N_8517,N_8434,N_8476);
and U8518 (N_8518,N_8483,N_8482);
and U8519 (N_8519,N_8433,N_8435);
nand U8520 (N_8520,N_8423,N_8406);
nand U8521 (N_8521,N_8444,N_8443);
nor U8522 (N_8522,N_8481,N_8404);
nor U8523 (N_8523,N_8489,N_8495);
nand U8524 (N_8524,N_8410,N_8416);
and U8525 (N_8525,N_8413,N_8441);
nor U8526 (N_8526,N_8494,N_8455);
nand U8527 (N_8527,N_8480,N_8421);
or U8528 (N_8528,N_8454,N_8458);
or U8529 (N_8529,N_8478,N_8470);
nor U8530 (N_8530,N_8456,N_8412);
and U8531 (N_8531,N_8403,N_8415);
nand U8532 (N_8532,N_8419,N_8436);
and U8533 (N_8533,N_8487,N_8429);
or U8534 (N_8534,N_8463,N_8428);
or U8535 (N_8535,N_8411,N_8488);
and U8536 (N_8536,N_8451,N_8491);
nor U8537 (N_8537,N_8479,N_8407);
nor U8538 (N_8538,N_8459,N_8469);
and U8539 (N_8539,N_8446,N_8414);
nor U8540 (N_8540,N_8467,N_8453);
nor U8541 (N_8541,N_8449,N_8477);
nor U8542 (N_8542,N_8422,N_8430);
and U8543 (N_8543,N_8493,N_8447);
nand U8544 (N_8544,N_8445,N_8472);
or U8545 (N_8545,N_8464,N_8485);
nor U8546 (N_8546,N_8496,N_8408);
or U8547 (N_8547,N_8450,N_8492);
nand U8548 (N_8548,N_8475,N_8484);
nor U8549 (N_8549,N_8473,N_8440);
and U8550 (N_8550,N_8419,N_8402);
and U8551 (N_8551,N_8410,N_8422);
nand U8552 (N_8552,N_8405,N_8492);
nand U8553 (N_8553,N_8492,N_8474);
and U8554 (N_8554,N_8467,N_8461);
and U8555 (N_8555,N_8488,N_8485);
nor U8556 (N_8556,N_8421,N_8487);
nor U8557 (N_8557,N_8414,N_8425);
and U8558 (N_8558,N_8439,N_8409);
and U8559 (N_8559,N_8474,N_8438);
nand U8560 (N_8560,N_8434,N_8497);
nor U8561 (N_8561,N_8414,N_8478);
nor U8562 (N_8562,N_8463,N_8439);
nand U8563 (N_8563,N_8405,N_8473);
and U8564 (N_8564,N_8482,N_8434);
nor U8565 (N_8565,N_8491,N_8466);
and U8566 (N_8566,N_8418,N_8484);
or U8567 (N_8567,N_8474,N_8421);
nor U8568 (N_8568,N_8492,N_8407);
and U8569 (N_8569,N_8482,N_8407);
or U8570 (N_8570,N_8454,N_8472);
or U8571 (N_8571,N_8407,N_8408);
nand U8572 (N_8572,N_8489,N_8428);
nand U8573 (N_8573,N_8407,N_8426);
and U8574 (N_8574,N_8463,N_8445);
nand U8575 (N_8575,N_8480,N_8496);
or U8576 (N_8576,N_8435,N_8426);
or U8577 (N_8577,N_8414,N_8491);
nand U8578 (N_8578,N_8492,N_8484);
nor U8579 (N_8579,N_8429,N_8412);
nand U8580 (N_8580,N_8435,N_8420);
nor U8581 (N_8581,N_8450,N_8420);
and U8582 (N_8582,N_8406,N_8439);
or U8583 (N_8583,N_8463,N_8478);
nor U8584 (N_8584,N_8459,N_8422);
nand U8585 (N_8585,N_8483,N_8466);
or U8586 (N_8586,N_8456,N_8424);
nand U8587 (N_8587,N_8433,N_8495);
nand U8588 (N_8588,N_8437,N_8462);
and U8589 (N_8589,N_8470,N_8484);
nand U8590 (N_8590,N_8404,N_8473);
nand U8591 (N_8591,N_8480,N_8490);
or U8592 (N_8592,N_8440,N_8459);
nor U8593 (N_8593,N_8426,N_8487);
nor U8594 (N_8594,N_8473,N_8479);
nand U8595 (N_8595,N_8416,N_8457);
nor U8596 (N_8596,N_8492,N_8410);
nor U8597 (N_8597,N_8413,N_8470);
or U8598 (N_8598,N_8457,N_8485);
nor U8599 (N_8599,N_8485,N_8441);
or U8600 (N_8600,N_8584,N_8554);
nand U8601 (N_8601,N_8558,N_8595);
nand U8602 (N_8602,N_8578,N_8540);
nand U8603 (N_8603,N_8504,N_8576);
or U8604 (N_8604,N_8511,N_8539);
nor U8605 (N_8605,N_8528,N_8500);
or U8606 (N_8606,N_8590,N_8547);
and U8607 (N_8607,N_8518,N_8535);
nor U8608 (N_8608,N_8510,N_8553);
xnor U8609 (N_8609,N_8561,N_8519);
nand U8610 (N_8610,N_8552,N_8524);
nor U8611 (N_8611,N_8573,N_8525);
or U8612 (N_8612,N_8507,N_8567);
and U8613 (N_8613,N_8502,N_8541);
and U8614 (N_8614,N_8522,N_8546);
or U8615 (N_8615,N_8588,N_8596);
or U8616 (N_8616,N_8563,N_8512);
or U8617 (N_8617,N_8572,N_8583);
nor U8618 (N_8618,N_8556,N_8569);
or U8619 (N_8619,N_8568,N_8562);
nor U8620 (N_8620,N_8594,N_8574);
nand U8621 (N_8621,N_8501,N_8542);
and U8622 (N_8622,N_8543,N_8538);
or U8623 (N_8623,N_8557,N_8533);
or U8624 (N_8624,N_8571,N_8506);
nand U8625 (N_8625,N_8555,N_8589);
and U8626 (N_8626,N_8551,N_8508);
and U8627 (N_8627,N_8566,N_8559);
nand U8628 (N_8628,N_8531,N_8544);
nand U8629 (N_8629,N_8526,N_8509);
or U8630 (N_8630,N_8534,N_8549);
and U8631 (N_8631,N_8577,N_8505);
and U8632 (N_8632,N_8581,N_8593);
nand U8633 (N_8633,N_8597,N_8503);
and U8634 (N_8634,N_8527,N_8520);
and U8635 (N_8635,N_8517,N_8591);
nand U8636 (N_8636,N_8570,N_8548);
nand U8637 (N_8637,N_8587,N_8514);
nor U8638 (N_8638,N_8585,N_8530);
nor U8639 (N_8639,N_8579,N_8513);
nand U8640 (N_8640,N_8592,N_8523);
or U8641 (N_8641,N_8516,N_8565);
and U8642 (N_8642,N_8564,N_8515);
and U8643 (N_8643,N_8575,N_8529);
nor U8644 (N_8644,N_8532,N_8580);
or U8645 (N_8645,N_8550,N_8537);
nor U8646 (N_8646,N_8586,N_8582);
nor U8647 (N_8647,N_8536,N_8560);
or U8648 (N_8648,N_8598,N_8545);
or U8649 (N_8649,N_8599,N_8521);
or U8650 (N_8650,N_8548,N_8529);
and U8651 (N_8651,N_8588,N_8585);
nor U8652 (N_8652,N_8533,N_8552);
nand U8653 (N_8653,N_8519,N_8548);
or U8654 (N_8654,N_8584,N_8548);
or U8655 (N_8655,N_8599,N_8588);
nor U8656 (N_8656,N_8549,N_8540);
or U8657 (N_8657,N_8568,N_8509);
nand U8658 (N_8658,N_8544,N_8533);
or U8659 (N_8659,N_8581,N_8579);
nor U8660 (N_8660,N_8502,N_8526);
nand U8661 (N_8661,N_8577,N_8568);
nor U8662 (N_8662,N_8554,N_8528);
nand U8663 (N_8663,N_8578,N_8524);
nor U8664 (N_8664,N_8529,N_8580);
nor U8665 (N_8665,N_8537,N_8538);
nand U8666 (N_8666,N_8586,N_8534);
and U8667 (N_8667,N_8573,N_8519);
nand U8668 (N_8668,N_8571,N_8593);
or U8669 (N_8669,N_8558,N_8539);
or U8670 (N_8670,N_8520,N_8526);
and U8671 (N_8671,N_8555,N_8542);
or U8672 (N_8672,N_8517,N_8514);
or U8673 (N_8673,N_8565,N_8576);
nand U8674 (N_8674,N_8582,N_8547);
nor U8675 (N_8675,N_8500,N_8568);
or U8676 (N_8676,N_8570,N_8567);
and U8677 (N_8677,N_8522,N_8586);
and U8678 (N_8678,N_8540,N_8534);
or U8679 (N_8679,N_8501,N_8523);
nor U8680 (N_8680,N_8584,N_8539);
nand U8681 (N_8681,N_8586,N_8599);
or U8682 (N_8682,N_8552,N_8506);
nor U8683 (N_8683,N_8572,N_8524);
nor U8684 (N_8684,N_8522,N_8576);
nor U8685 (N_8685,N_8564,N_8562);
nor U8686 (N_8686,N_8589,N_8529);
nand U8687 (N_8687,N_8553,N_8546);
nor U8688 (N_8688,N_8583,N_8552);
and U8689 (N_8689,N_8544,N_8507);
nand U8690 (N_8690,N_8599,N_8504);
and U8691 (N_8691,N_8512,N_8513);
or U8692 (N_8692,N_8566,N_8551);
nor U8693 (N_8693,N_8594,N_8559);
nor U8694 (N_8694,N_8579,N_8541);
nand U8695 (N_8695,N_8592,N_8541);
or U8696 (N_8696,N_8569,N_8597);
nor U8697 (N_8697,N_8556,N_8509);
nor U8698 (N_8698,N_8505,N_8580);
nor U8699 (N_8699,N_8596,N_8543);
nand U8700 (N_8700,N_8676,N_8667);
nand U8701 (N_8701,N_8678,N_8616);
nand U8702 (N_8702,N_8693,N_8688);
nand U8703 (N_8703,N_8658,N_8630);
or U8704 (N_8704,N_8602,N_8660);
and U8705 (N_8705,N_8686,N_8672);
nand U8706 (N_8706,N_8639,N_8666);
nor U8707 (N_8707,N_8631,N_8657);
or U8708 (N_8708,N_8662,N_8609);
and U8709 (N_8709,N_8668,N_8663);
or U8710 (N_8710,N_8612,N_8644);
or U8711 (N_8711,N_8617,N_8684);
or U8712 (N_8712,N_8622,N_8665);
or U8713 (N_8713,N_8611,N_8652);
or U8714 (N_8714,N_8603,N_8637);
nand U8715 (N_8715,N_8681,N_8600);
or U8716 (N_8716,N_8623,N_8669);
nand U8717 (N_8717,N_8692,N_8650);
and U8718 (N_8718,N_8634,N_8624);
nand U8719 (N_8719,N_8696,N_8641);
nor U8720 (N_8720,N_8689,N_8643);
nand U8721 (N_8721,N_8629,N_8677);
nand U8722 (N_8722,N_8649,N_8605);
nor U8723 (N_8723,N_8648,N_8654);
nand U8724 (N_8724,N_8620,N_8655);
nand U8725 (N_8725,N_8691,N_8604);
nand U8726 (N_8726,N_8679,N_8638);
nor U8727 (N_8727,N_8697,N_8633);
xnor U8728 (N_8728,N_8673,N_8601);
nand U8729 (N_8729,N_8640,N_8699);
or U8730 (N_8730,N_8656,N_8695);
or U8731 (N_8731,N_8614,N_8664);
or U8732 (N_8732,N_8698,N_8694);
or U8733 (N_8733,N_8627,N_8674);
nor U8734 (N_8734,N_8621,N_8635);
or U8735 (N_8735,N_8683,N_8625);
nand U8736 (N_8736,N_8642,N_8610);
and U8737 (N_8737,N_8670,N_8646);
or U8738 (N_8738,N_8619,N_8636);
nor U8739 (N_8739,N_8645,N_8682);
and U8740 (N_8740,N_8632,N_8647);
or U8741 (N_8741,N_8687,N_8675);
nor U8742 (N_8742,N_8685,N_8659);
nor U8743 (N_8743,N_8615,N_8618);
nand U8744 (N_8744,N_8608,N_8671);
or U8745 (N_8745,N_8626,N_8661);
nand U8746 (N_8746,N_8613,N_8653);
or U8747 (N_8747,N_8690,N_8607);
or U8748 (N_8748,N_8628,N_8606);
or U8749 (N_8749,N_8680,N_8651);
and U8750 (N_8750,N_8698,N_8693);
and U8751 (N_8751,N_8616,N_8661);
or U8752 (N_8752,N_8696,N_8688);
and U8753 (N_8753,N_8686,N_8668);
or U8754 (N_8754,N_8655,N_8623);
nand U8755 (N_8755,N_8634,N_8609);
nor U8756 (N_8756,N_8671,N_8621);
nor U8757 (N_8757,N_8659,N_8606);
nand U8758 (N_8758,N_8699,N_8647);
nand U8759 (N_8759,N_8675,N_8629);
or U8760 (N_8760,N_8610,N_8608);
or U8761 (N_8761,N_8676,N_8697);
or U8762 (N_8762,N_8645,N_8622);
and U8763 (N_8763,N_8627,N_8694);
or U8764 (N_8764,N_8676,N_8641);
or U8765 (N_8765,N_8653,N_8637);
and U8766 (N_8766,N_8640,N_8629);
or U8767 (N_8767,N_8685,N_8606);
and U8768 (N_8768,N_8693,N_8643);
and U8769 (N_8769,N_8613,N_8649);
nand U8770 (N_8770,N_8687,N_8612);
and U8771 (N_8771,N_8654,N_8664);
nand U8772 (N_8772,N_8685,N_8611);
or U8773 (N_8773,N_8625,N_8606);
nand U8774 (N_8774,N_8693,N_8649);
nand U8775 (N_8775,N_8611,N_8625);
nor U8776 (N_8776,N_8622,N_8606);
nor U8777 (N_8777,N_8681,N_8606);
nand U8778 (N_8778,N_8617,N_8634);
nand U8779 (N_8779,N_8650,N_8617);
or U8780 (N_8780,N_8688,N_8652);
nand U8781 (N_8781,N_8687,N_8604);
or U8782 (N_8782,N_8614,N_8662);
nand U8783 (N_8783,N_8670,N_8656);
and U8784 (N_8784,N_8613,N_8627);
nor U8785 (N_8785,N_8651,N_8670);
or U8786 (N_8786,N_8671,N_8616);
and U8787 (N_8787,N_8606,N_8698);
or U8788 (N_8788,N_8628,N_8630);
or U8789 (N_8789,N_8640,N_8697);
or U8790 (N_8790,N_8692,N_8686);
or U8791 (N_8791,N_8682,N_8688);
nor U8792 (N_8792,N_8646,N_8660);
nand U8793 (N_8793,N_8628,N_8686);
and U8794 (N_8794,N_8666,N_8640);
nand U8795 (N_8795,N_8674,N_8657);
nand U8796 (N_8796,N_8600,N_8606);
nand U8797 (N_8797,N_8657,N_8630);
nor U8798 (N_8798,N_8624,N_8668);
or U8799 (N_8799,N_8629,N_8680);
or U8800 (N_8800,N_8714,N_8759);
nor U8801 (N_8801,N_8727,N_8741);
and U8802 (N_8802,N_8777,N_8790);
and U8803 (N_8803,N_8760,N_8707);
and U8804 (N_8804,N_8746,N_8750);
and U8805 (N_8805,N_8775,N_8755);
nand U8806 (N_8806,N_8739,N_8751);
nand U8807 (N_8807,N_8743,N_8797);
nor U8808 (N_8808,N_8796,N_8791);
nand U8809 (N_8809,N_8736,N_8734);
or U8810 (N_8810,N_8798,N_8780);
nand U8811 (N_8811,N_8776,N_8769);
and U8812 (N_8812,N_8719,N_8704);
and U8813 (N_8813,N_8722,N_8799);
nand U8814 (N_8814,N_8781,N_8749);
or U8815 (N_8815,N_8758,N_8764);
or U8816 (N_8816,N_8752,N_8718);
and U8817 (N_8817,N_8783,N_8766);
nand U8818 (N_8818,N_8710,N_8779);
nand U8819 (N_8819,N_8772,N_8716);
and U8820 (N_8820,N_8706,N_8723);
or U8821 (N_8821,N_8711,N_8725);
or U8822 (N_8822,N_8782,N_8738);
or U8823 (N_8823,N_8768,N_8709);
nand U8824 (N_8824,N_8732,N_8701);
nor U8825 (N_8825,N_8733,N_8773);
nand U8826 (N_8826,N_8745,N_8715);
or U8827 (N_8827,N_8740,N_8712);
or U8828 (N_8828,N_8729,N_8705);
and U8829 (N_8829,N_8754,N_8765);
nand U8830 (N_8830,N_8737,N_8708);
nor U8831 (N_8831,N_8785,N_8744);
and U8832 (N_8832,N_8720,N_8786);
nor U8833 (N_8833,N_8795,N_8702);
nand U8834 (N_8834,N_8726,N_8700);
nor U8835 (N_8835,N_8771,N_8735);
nand U8836 (N_8836,N_8770,N_8788);
xnor U8837 (N_8837,N_8778,N_8703);
and U8838 (N_8838,N_8728,N_8792);
or U8839 (N_8839,N_8784,N_8767);
or U8840 (N_8840,N_8747,N_8730);
or U8841 (N_8841,N_8763,N_8787);
or U8842 (N_8842,N_8789,N_8717);
or U8843 (N_8843,N_8742,N_8774);
nand U8844 (N_8844,N_8753,N_8793);
or U8845 (N_8845,N_8748,N_8757);
nor U8846 (N_8846,N_8731,N_8724);
or U8847 (N_8847,N_8713,N_8756);
or U8848 (N_8848,N_8721,N_8761);
nor U8849 (N_8849,N_8762,N_8794);
and U8850 (N_8850,N_8771,N_8798);
and U8851 (N_8851,N_8724,N_8707);
and U8852 (N_8852,N_8791,N_8727);
and U8853 (N_8853,N_8781,N_8785);
nor U8854 (N_8854,N_8700,N_8762);
and U8855 (N_8855,N_8734,N_8700);
or U8856 (N_8856,N_8771,N_8708);
nor U8857 (N_8857,N_8786,N_8750);
and U8858 (N_8858,N_8764,N_8759);
or U8859 (N_8859,N_8753,N_8769);
nand U8860 (N_8860,N_8740,N_8724);
or U8861 (N_8861,N_8749,N_8754);
nand U8862 (N_8862,N_8709,N_8756);
and U8863 (N_8863,N_8745,N_8788);
nor U8864 (N_8864,N_8770,N_8758);
or U8865 (N_8865,N_8718,N_8788);
or U8866 (N_8866,N_8783,N_8768);
nor U8867 (N_8867,N_8735,N_8734);
nor U8868 (N_8868,N_8788,N_8763);
nor U8869 (N_8869,N_8708,N_8751);
nor U8870 (N_8870,N_8780,N_8713);
nand U8871 (N_8871,N_8772,N_8726);
or U8872 (N_8872,N_8702,N_8798);
or U8873 (N_8873,N_8764,N_8748);
nand U8874 (N_8874,N_8777,N_8787);
or U8875 (N_8875,N_8723,N_8758);
nor U8876 (N_8876,N_8754,N_8770);
and U8877 (N_8877,N_8748,N_8767);
nor U8878 (N_8878,N_8745,N_8784);
nand U8879 (N_8879,N_8758,N_8737);
or U8880 (N_8880,N_8780,N_8739);
nor U8881 (N_8881,N_8754,N_8720);
nor U8882 (N_8882,N_8731,N_8719);
nand U8883 (N_8883,N_8727,N_8717);
nor U8884 (N_8884,N_8785,N_8773);
nand U8885 (N_8885,N_8797,N_8708);
and U8886 (N_8886,N_8705,N_8715);
and U8887 (N_8887,N_8786,N_8751);
nand U8888 (N_8888,N_8706,N_8740);
nor U8889 (N_8889,N_8720,N_8745);
nand U8890 (N_8890,N_8778,N_8709);
and U8891 (N_8891,N_8752,N_8773);
nor U8892 (N_8892,N_8790,N_8749);
nand U8893 (N_8893,N_8728,N_8784);
nor U8894 (N_8894,N_8752,N_8729);
or U8895 (N_8895,N_8773,N_8772);
nor U8896 (N_8896,N_8721,N_8796);
or U8897 (N_8897,N_8705,N_8784);
nand U8898 (N_8898,N_8704,N_8713);
nand U8899 (N_8899,N_8760,N_8730);
nand U8900 (N_8900,N_8848,N_8884);
and U8901 (N_8901,N_8804,N_8839);
nand U8902 (N_8902,N_8802,N_8855);
and U8903 (N_8903,N_8856,N_8885);
nor U8904 (N_8904,N_8894,N_8811);
nor U8905 (N_8905,N_8863,N_8854);
and U8906 (N_8906,N_8897,N_8853);
and U8907 (N_8907,N_8898,N_8859);
nand U8908 (N_8908,N_8806,N_8846);
or U8909 (N_8909,N_8867,N_8823);
or U8910 (N_8910,N_8895,N_8824);
and U8911 (N_8911,N_8843,N_8887);
nand U8912 (N_8912,N_8876,N_8865);
or U8913 (N_8913,N_8814,N_8810);
and U8914 (N_8914,N_8857,N_8891);
and U8915 (N_8915,N_8808,N_8842);
and U8916 (N_8916,N_8819,N_8886);
or U8917 (N_8917,N_8869,N_8866);
nor U8918 (N_8918,N_8816,N_8851);
nand U8919 (N_8919,N_8892,N_8822);
nor U8920 (N_8920,N_8850,N_8880);
and U8921 (N_8921,N_8828,N_8807);
and U8922 (N_8922,N_8833,N_8815);
or U8923 (N_8923,N_8861,N_8831);
and U8924 (N_8924,N_8834,N_8847);
nor U8925 (N_8925,N_8829,N_8841);
nand U8926 (N_8926,N_8835,N_8871);
nand U8927 (N_8927,N_8862,N_8836);
or U8928 (N_8928,N_8893,N_8877);
or U8929 (N_8929,N_8870,N_8826);
nand U8930 (N_8930,N_8821,N_8817);
and U8931 (N_8931,N_8832,N_8858);
nor U8932 (N_8932,N_8852,N_8849);
and U8933 (N_8933,N_8874,N_8883);
and U8934 (N_8934,N_8801,N_8882);
xor U8935 (N_8935,N_8872,N_8890);
nor U8936 (N_8936,N_8805,N_8879);
or U8937 (N_8937,N_8840,N_8825);
nor U8938 (N_8938,N_8888,N_8889);
nor U8939 (N_8939,N_8844,N_8820);
or U8940 (N_8940,N_8896,N_8809);
or U8941 (N_8941,N_8873,N_8813);
and U8942 (N_8942,N_8827,N_8878);
or U8943 (N_8943,N_8899,N_8845);
or U8944 (N_8944,N_8800,N_8868);
and U8945 (N_8945,N_8818,N_8860);
or U8946 (N_8946,N_8838,N_8881);
and U8947 (N_8947,N_8837,N_8803);
and U8948 (N_8948,N_8864,N_8875);
xor U8949 (N_8949,N_8812,N_8830);
and U8950 (N_8950,N_8877,N_8807);
nor U8951 (N_8951,N_8874,N_8865);
xnor U8952 (N_8952,N_8871,N_8816);
nor U8953 (N_8953,N_8843,N_8861);
nand U8954 (N_8954,N_8881,N_8861);
nor U8955 (N_8955,N_8873,N_8883);
nor U8956 (N_8956,N_8873,N_8804);
xor U8957 (N_8957,N_8898,N_8832);
and U8958 (N_8958,N_8847,N_8821);
nand U8959 (N_8959,N_8804,N_8856);
nor U8960 (N_8960,N_8806,N_8821);
nor U8961 (N_8961,N_8886,N_8838);
nand U8962 (N_8962,N_8897,N_8874);
nor U8963 (N_8963,N_8878,N_8865);
nand U8964 (N_8964,N_8889,N_8870);
nor U8965 (N_8965,N_8827,N_8816);
or U8966 (N_8966,N_8819,N_8818);
or U8967 (N_8967,N_8841,N_8891);
nor U8968 (N_8968,N_8873,N_8891);
or U8969 (N_8969,N_8832,N_8857);
nor U8970 (N_8970,N_8803,N_8820);
and U8971 (N_8971,N_8861,N_8883);
nand U8972 (N_8972,N_8817,N_8884);
nand U8973 (N_8973,N_8835,N_8875);
nor U8974 (N_8974,N_8830,N_8877);
nor U8975 (N_8975,N_8859,N_8878);
nor U8976 (N_8976,N_8826,N_8892);
or U8977 (N_8977,N_8830,N_8869);
nor U8978 (N_8978,N_8811,N_8875);
nor U8979 (N_8979,N_8886,N_8851);
nand U8980 (N_8980,N_8892,N_8858);
and U8981 (N_8981,N_8818,N_8866);
and U8982 (N_8982,N_8846,N_8877);
nor U8983 (N_8983,N_8856,N_8834);
nor U8984 (N_8984,N_8859,N_8881);
nand U8985 (N_8985,N_8838,N_8816);
and U8986 (N_8986,N_8801,N_8845);
or U8987 (N_8987,N_8816,N_8802);
and U8988 (N_8988,N_8849,N_8840);
nor U8989 (N_8989,N_8825,N_8889);
or U8990 (N_8990,N_8857,N_8863);
or U8991 (N_8991,N_8836,N_8846);
and U8992 (N_8992,N_8824,N_8814);
and U8993 (N_8993,N_8863,N_8884);
or U8994 (N_8994,N_8894,N_8813);
and U8995 (N_8995,N_8898,N_8883);
nand U8996 (N_8996,N_8894,N_8812);
and U8997 (N_8997,N_8883,N_8837);
nand U8998 (N_8998,N_8899,N_8850);
nor U8999 (N_8999,N_8856,N_8853);
and U9000 (N_9000,N_8988,N_8945);
nor U9001 (N_9001,N_8997,N_8989);
or U9002 (N_9002,N_8911,N_8944);
or U9003 (N_9003,N_8904,N_8900);
nor U9004 (N_9004,N_8923,N_8943);
nor U9005 (N_9005,N_8968,N_8946);
and U9006 (N_9006,N_8920,N_8955);
nor U9007 (N_9007,N_8907,N_8986);
nand U9008 (N_9008,N_8921,N_8973);
or U9009 (N_9009,N_8980,N_8967);
nor U9010 (N_9010,N_8910,N_8931);
nor U9011 (N_9011,N_8970,N_8932);
nand U9012 (N_9012,N_8974,N_8924);
nor U9013 (N_9013,N_8965,N_8981);
and U9014 (N_9014,N_8982,N_8901);
or U9015 (N_9015,N_8971,N_8929);
nand U9016 (N_9016,N_8903,N_8952);
or U9017 (N_9017,N_8950,N_8998);
or U9018 (N_9018,N_8937,N_8947);
nor U9019 (N_9019,N_8956,N_8960);
nand U9020 (N_9020,N_8962,N_8948);
and U9021 (N_9021,N_8977,N_8963);
or U9022 (N_9022,N_8966,N_8939);
or U9023 (N_9023,N_8969,N_8938);
or U9024 (N_9024,N_8934,N_8908);
or U9025 (N_9025,N_8994,N_8916);
and U9026 (N_9026,N_8995,N_8959);
nor U9027 (N_9027,N_8919,N_8999);
or U9028 (N_9028,N_8978,N_8915);
and U9029 (N_9029,N_8925,N_8933);
and U9030 (N_9030,N_8913,N_8912);
or U9031 (N_9031,N_8964,N_8957);
and U9032 (N_9032,N_8985,N_8940);
or U9033 (N_9033,N_8975,N_8983);
xnor U9034 (N_9034,N_8935,N_8976);
and U9035 (N_9035,N_8987,N_8918);
and U9036 (N_9036,N_8941,N_8906);
or U9037 (N_9037,N_8936,N_8953);
nand U9038 (N_9038,N_8996,N_8954);
nor U9039 (N_9039,N_8922,N_8909);
and U9040 (N_9040,N_8914,N_8979);
or U9041 (N_9041,N_8961,N_8993);
nand U9042 (N_9042,N_8927,N_8984);
nand U9043 (N_9043,N_8990,N_8928);
nand U9044 (N_9044,N_8972,N_8917);
or U9045 (N_9045,N_8992,N_8951);
and U9046 (N_9046,N_8958,N_8949);
or U9047 (N_9047,N_8991,N_8930);
or U9048 (N_9048,N_8902,N_8942);
and U9049 (N_9049,N_8905,N_8926);
and U9050 (N_9050,N_8953,N_8968);
or U9051 (N_9051,N_8994,N_8950);
xor U9052 (N_9052,N_8953,N_8981);
or U9053 (N_9053,N_8988,N_8966);
or U9054 (N_9054,N_8982,N_8973);
and U9055 (N_9055,N_8957,N_8924);
nand U9056 (N_9056,N_8969,N_8926);
nand U9057 (N_9057,N_8937,N_8932);
or U9058 (N_9058,N_8919,N_8923);
nand U9059 (N_9059,N_8998,N_8981);
nand U9060 (N_9060,N_8914,N_8910);
nand U9061 (N_9061,N_8959,N_8974);
and U9062 (N_9062,N_8957,N_8918);
and U9063 (N_9063,N_8979,N_8960);
or U9064 (N_9064,N_8954,N_8950);
and U9065 (N_9065,N_8985,N_8934);
nand U9066 (N_9066,N_8976,N_8955);
and U9067 (N_9067,N_8912,N_8991);
and U9068 (N_9068,N_8960,N_8962);
nor U9069 (N_9069,N_8970,N_8955);
nand U9070 (N_9070,N_8997,N_8924);
or U9071 (N_9071,N_8953,N_8958);
nor U9072 (N_9072,N_8940,N_8969);
nor U9073 (N_9073,N_8922,N_8991);
and U9074 (N_9074,N_8909,N_8902);
or U9075 (N_9075,N_8900,N_8912);
nand U9076 (N_9076,N_8927,N_8999);
nand U9077 (N_9077,N_8970,N_8999);
nand U9078 (N_9078,N_8902,N_8934);
or U9079 (N_9079,N_8926,N_8914);
or U9080 (N_9080,N_8944,N_8901);
xor U9081 (N_9081,N_8997,N_8917);
or U9082 (N_9082,N_8922,N_8917);
nand U9083 (N_9083,N_8968,N_8917);
and U9084 (N_9084,N_8917,N_8930);
or U9085 (N_9085,N_8994,N_8914);
and U9086 (N_9086,N_8937,N_8994);
and U9087 (N_9087,N_8923,N_8967);
nand U9088 (N_9088,N_8955,N_8962);
and U9089 (N_9089,N_8901,N_8934);
or U9090 (N_9090,N_8926,N_8990);
and U9091 (N_9091,N_8920,N_8906);
nor U9092 (N_9092,N_8923,N_8916);
nand U9093 (N_9093,N_8917,N_8950);
and U9094 (N_9094,N_8995,N_8973);
nor U9095 (N_9095,N_8931,N_8918);
nor U9096 (N_9096,N_8914,N_8922);
nand U9097 (N_9097,N_8985,N_8954);
nand U9098 (N_9098,N_8908,N_8955);
or U9099 (N_9099,N_8933,N_8926);
and U9100 (N_9100,N_9001,N_9099);
nor U9101 (N_9101,N_9007,N_9071);
and U9102 (N_9102,N_9022,N_9021);
nand U9103 (N_9103,N_9050,N_9064);
or U9104 (N_9104,N_9082,N_9085);
nor U9105 (N_9105,N_9093,N_9024);
and U9106 (N_9106,N_9025,N_9033);
or U9107 (N_9107,N_9056,N_9074);
or U9108 (N_9108,N_9026,N_9004);
or U9109 (N_9109,N_9098,N_9047);
nor U9110 (N_9110,N_9058,N_9059);
nand U9111 (N_9111,N_9006,N_9072);
and U9112 (N_9112,N_9087,N_9018);
and U9113 (N_9113,N_9029,N_9015);
nand U9114 (N_9114,N_9063,N_9002);
and U9115 (N_9115,N_9016,N_9081);
and U9116 (N_9116,N_9048,N_9094);
or U9117 (N_9117,N_9070,N_9017);
and U9118 (N_9118,N_9075,N_9027);
or U9119 (N_9119,N_9068,N_9073);
and U9120 (N_9120,N_9010,N_9080);
or U9121 (N_9121,N_9020,N_9091);
nor U9122 (N_9122,N_9051,N_9088);
or U9123 (N_9123,N_9061,N_9036);
and U9124 (N_9124,N_9083,N_9039);
or U9125 (N_9125,N_9043,N_9078);
nor U9126 (N_9126,N_9079,N_9037);
nor U9127 (N_9127,N_9023,N_9012);
nor U9128 (N_9128,N_9000,N_9097);
nor U9129 (N_9129,N_9019,N_9057);
nand U9130 (N_9130,N_9038,N_9013);
nor U9131 (N_9131,N_9005,N_9003);
nand U9132 (N_9132,N_9041,N_9046);
and U9133 (N_9133,N_9034,N_9089);
and U9134 (N_9134,N_9011,N_9049);
and U9135 (N_9135,N_9008,N_9060);
nand U9136 (N_9136,N_9067,N_9069);
nand U9137 (N_9137,N_9052,N_9042);
and U9138 (N_9138,N_9054,N_9096);
nand U9139 (N_9139,N_9040,N_9062);
or U9140 (N_9140,N_9044,N_9009);
nor U9141 (N_9141,N_9092,N_9086);
and U9142 (N_9142,N_9077,N_9028);
or U9143 (N_9143,N_9032,N_9053);
nand U9144 (N_9144,N_9066,N_9035);
or U9145 (N_9145,N_9095,N_9014);
nor U9146 (N_9146,N_9055,N_9090);
nand U9147 (N_9147,N_9084,N_9045);
or U9148 (N_9148,N_9065,N_9076);
nor U9149 (N_9149,N_9031,N_9030);
nor U9150 (N_9150,N_9044,N_9073);
nand U9151 (N_9151,N_9048,N_9017);
nor U9152 (N_9152,N_9049,N_9065);
nand U9153 (N_9153,N_9023,N_9003);
nand U9154 (N_9154,N_9038,N_9016);
nand U9155 (N_9155,N_9015,N_9063);
or U9156 (N_9156,N_9094,N_9090);
nand U9157 (N_9157,N_9077,N_9058);
nor U9158 (N_9158,N_9013,N_9045);
xor U9159 (N_9159,N_9090,N_9009);
nor U9160 (N_9160,N_9073,N_9011);
and U9161 (N_9161,N_9047,N_9049);
and U9162 (N_9162,N_9096,N_9050);
or U9163 (N_9163,N_9053,N_9082);
and U9164 (N_9164,N_9069,N_9097);
nor U9165 (N_9165,N_9003,N_9059);
nor U9166 (N_9166,N_9034,N_9063);
and U9167 (N_9167,N_9051,N_9021);
or U9168 (N_9168,N_9020,N_9017);
and U9169 (N_9169,N_9048,N_9074);
nand U9170 (N_9170,N_9083,N_9089);
nor U9171 (N_9171,N_9095,N_9077);
nor U9172 (N_9172,N_9001,N_9046);
or U9173 (N_9173,N_9014,N_9080);
and U9174 (N_9174,N_9070,N_9098);
or U9175 (N_9175,N_9052,N_9087);
nand U9176 (N_9176,N_9030,N_9052);
and U9177 (N_9177,N_9064,N_9068);
and U9178 (N_9178,N_9074,N_9032);
and U9179 (N_9179,N_9093,N_9060);
and U9180 (N_9180,N_9095,N_9049);
nor U9181 (N_9181,N_9040,N_9060);
nor U9182 (N_9182,N_9023,N_9004);
or U9183 (N_9183,N_9059,N_9023);
nor U9184 (N_9184,N_9072,N_9011);
nor U9185 (N_9185,N_9063,N_9043);
nor U9186 (N_9186,N_9086,N_9025);
nand U9187 (N_9187,N_9052,N_9077);
nand U9188 (N_9188,N_9067,N_9025);
or U9189 (N_9189,N_9068,N_9054);
nor U9190 (N_9190,N_9018,N_9044);
or U9191 (N_9191,N_9095,N_9097);
and U9192 (N_9192,N_9013,N_9089);
and U9193 (N_9193,N_9091,N_9004);
and U9194 (N_9194,N_9081,N_9060);
or U9195 (N_9195,N_9024,N_9012);
and U9196 (N_9196,N_9056,N_9064);
or U9197 (N_9197,N_9089,N_9077);
nor U9198 (N_9198,N_9022,N_9072);
nand U9199 (N_9199,N_9070,N_9046);
nor U9200 (N_9200,N_9185,N_9158);
and U9201 (N_9201,N_9177,N_9102);
or U9202 (N_9202,N_9196,N_9100);
nor U9203 (N_9203,N_9126,N_9124);
and U9204 (N_9204,N_9164,N_9143);
nand U9205 (N_9205,N_9156,N_9195);
nand U9206 (N_9206,N_9190,N_9197);
or U9207 (N_9207,N_9169,N_9103);
or U9208 (N_9208,N_9175,N_9173);
and U9209 (N_9209,N_9199,N_9165);
or U9210 (N_9210,N_9117,N_9151);
or U9211 (N_9211,N_9183,N_9191);
or U9212 (N_9212,N_9178,N_9149);
nor U9213 (N_9213,N_9127,N_9128);
or U9214 (N_9214,N_9116,N_9188);
nand U9215 (N_9215,N_9181,N_9147);
nand U9216 (N_9216,N_9109,N_9110);
nand U9217 (N_9217,N_9137,N_9153);
nand U9218 (N_9218,N_9133,N_9154);
nand U9219 (N_9219,N_9138,N_9142);
nor U9220 (N_9220,N_9118,N_9112);
nor U9221 (N_9221,N_9123,N_9170);
nand U9222 (N_9222,N_9174,N_9150);
and U9223 (N_9223,N_9114,N_9182);
or U9224 (N_9224,N_9184,N_9193);
and U9225 (N_9225,N_9130,N_9145);
or U9226 (N_9226,N_9120,N_9125);
and U9227 (N_9227,N_9179,N_9172);
nor U9228 (N_9228,N_9111,N_9157);
nor U9229 (N_9229,N_9161,N_9163);
nand U9230 (N_9230,N_9171,N_9113);
nor U9231 (N_9231,N_9131,N_9122);
and U9232 (N_9232,N_9107,N_9167);
nand U9233 (N_9233,N_9155,N_9187);
and U9234 (N_9234,N_9136,N_9132);
and U9235 (N_9235,N_9194,N_9108);
or U9236 (N_9236,N_9104,N_9180);
nor U9237 (N_9237,N_9186,N_9159);
and U9238 (N_9238,N_9101,N_9135);
or U9239 (N_9239,N_9141,N_9119);
and U9240 (N_9240,N_9160,N_9144);
or U9241 (N_9241,N_9140,N_9115);
nand U9242 (N_9242,N_9168,N_9121);
or U9243 (N_9243,N_9134,N_9198);
nand U9244 (N_9244,N_9129,N_9105);
or U9245 (N_9245,N_9162,N_9176);
or U9246 (N_9246,N_9189,N_9148);
and U9247 (N_9247,N_9166,N_9146);
and U9248 (N_9248,N_9106,N_9152);
or U9249 (N_9249,N_9192,N_9139);
or U9250 (N_9250,N_9108,N_9138);
and U9251 (N_9251,N_9134,N_9148);
and U9252 (N_9252,N_9113,N_9180);
nor U9253 (N_9253,N_9174,N_9179);
or U9254 (N_9254,N_9119,N_9132);
and U9255 (N_9255,N_9171,N_9102);
nor U9256 (N_9256,N_9176,N_9166);
and U9257 (N_9257,N_9176,N_9148);
or U9258 (N_9258,N_9195,N_9139);
or U9259 (N_9259,N_9102,N_9147);
nand U9260 (N_9260,N_9193,N_9111);
nor U9261 (N_9261,N_9123,N_9136);
and U9262 (N_9262,N_9176,N_9109);
or U9263 (N_9263,N_9109,N_9194);
nand U9264 (N_9264,N_9181,N_9160);
nand U9265 (N_9265,N_9161,N_9108);
and U9266 (N_9266,N_9120,N_9136);
nand U9267 (N_9267,N_9191,N_9163);
and U9268 (N_9268,N_9198,N_9191);
and U9269 (N_9269,N_9127,N_9107);
nand U9270 (N_9270,N_9180,N_9116);
or U9271 (N_9271,N_9153,N_9176);
and U9272 (N_9272,N_9135,N_9152);
nand U9273 (N_9273,N_9188,N_9112);
nand U9274 (N_9274,N_9139,N_9110);
or U9275 (N_9275,N_9138,N_9164);
or U9276 (N_9276,N_9142,N_9190);
nand U9277 (N_9277,N_9129,N_9139);
and U9278 (N_9278,N_9141,N_9152);
nand U9279 (N_9279,N_9112,N_9176);
and U9280 (N_9280,N_9128,N_9107);
nand U9281 (N_9281,N_9171,N_9193);
and U9282 (N_9282,N_9176,N_9131);
nor U9283 (N_9283,N_9123,N_9115);
or U9284 (N_9284,N_9122,N_9124);
nor U9285 (N_9285,N_9143,N_9146);
and U9286 (N_9286,N_9106,N_9171);
nand U9287 (N_9287,N_9178,N_9101);
nand U9288 (N_9288,N_9190,N_9119);
or U9289 (N_9289,N_9120,N_9189);
and U9290 (N_9290,N_9139,N_9167);
nand U9291 (N_9291,N_9180,N_9179);
nand U9292 (N_9292,N_9131,N_9157);
nor U9293 (N_9293,N_9158,N_9198);
or U9294 (N_9294,N_9177,N_9182);
nand U9295 (N_9295,N_9135,N_9151);
or U9296 (N_9296,N_9102,N_9198);
nor U9297 (N_9297,N_9147,N_9177);
and U9298 (N_9298,N_9193,N_9182);
or U9299 (N_9299,N_9171,N_9140);
nor U9300 (N_9300,N_9281,N_9278);
nor U9301 (N_9301,N_9223,N_9231);
nand U9302 (N_9302,N_9277,N_9293);
or U9303 (N_9303,N_9259,N_9207);
and U9304 (N_9304,N_9225,N_9280);
nand U9305 (N_9305,N_9286,N_9244);
nand U9306 (N_9306,N_9284,N_9239);
nand U9307 (N_9307,N_9257,N_9227);
and U9308 (N_9308,N_9263,N_9200);
or U9309 (N_9309,N_9224,N_9233);
nand U9310 (N_9310,N_9218,N_9251);
nor U9311 (N_9311,N_9245,N_9241);
or U9312 (N_9312,N_9228,N_9209);
and U9313 (N_9313,N_9213,N_9220);
nand U9314 (N_9314,N_9237,N_9285);
nand U9315 (N_9315,N_9279,N_9282);
and U9316 (N_9316,N_9268,N_9214);
or U9317 (N_9317,N_9266,N_9270);
or U9318 (N_9318,N_9217,N_9248);
and U9319 (N_9319,N_9221,N_9273);
nand U9320 (N_9320,N_9205,N_9288);
nand U9321 (N_9321,N_9290,N_9272);
nor U9322 (N_9322,N_9222,N_9208);
or U9323 (N_9323,N_9256,N_9206);
nor U9324 (N_9324,N_9274,N_9238);
nand U9325 (N_9325,N_9276,N_9265);
nand U9326 (N_9326,N_9201,N_9295);
nor U9327 (N_9327,N_9287,N_9226);
and U9328 (N_9328,N_9230,N_9299);
and U9329 (N_9329,N_9262,N_9264);
and U9330 (N_9330,N_9249,N_9267);
or U9331 (N_9331,N_9243,N_9269);
nand U9332 (N_9332,N_9253,N_9212);
nand U9333 (N_9333,N_9204,N_9246);
or U9334 (N_9334,N_9234,N_9254);
nand U9335 (N_9335,N_9294,N_9211);
or U9336 (N_9336,N_9291,N_9240);
or U9337 (N_9337,N_9297,N_9202);
and U9338 (N_9338,N_9260,N_9232);
or U9339 (N_9339,N_9298,N_9215);
and U9340 (N_9340,N_9229,N_9296);
nand U9341 (N_9341,N_9216,N_9252);
and U9342 (N_9342,N_9258,N_9210);
nor U9343 (N_9343,N_9275,N_9203);
nor U9344 (N_9344,N_9283,N_9250);
nand U9345 (N_9345,N_9271,N_9255);
nor U9346 (N_9346,N_9236,N_9219);
or U9347 (N_9347,N_9261,N_9242);
nand U9348 (N_9348,N_9247,N_9289);
nor U9349 (N_9349,N_9292,N_9235);
and U9350 (N_9350,N_9227,N_9200);
or U9351 (N_9351,N_9228,N_9251);
or U9352 (N_9352,N_9283,N_9202);
nand U9353 (N_9353,N_9268,N_9230);
and U9354 (N_9354,N_9231,N_9249);
or U9355 (N_9355,N_9248,N_9220);
and U9356 (N_9356,N_9297,N_9203);
or U9357 (N_9357,N_9204,N_9294);
and U9358 (N_9358,N_9242,N_9263);
and U9359 (N_9359,N_9291,N_9288);
nand U9360 (N_9360,N_9284,N_9224);
nor U9361 (N_9361,N_9249,N_9233);
or U9362 (N_9362,N_9208,N_9256);
nand U9363 (N_9363,N_9216,N_9214);
nor U9364 (N_9364,N_9236,N_9265);
or U9365 (N_9365,N_9249,N_9296);
nand U9366 (N_9366,N_9252,N_9248);
and U9367 (N_9367,N_9282,N_9249);
and U9368 (N_9368,N_9255,N_9237);
xnor U9369 (N_9369,N_9264,N_9268);
nor U9370 (N_9370,N_9232,N_9272);
and U9371 (N_9371,N_9245,N_9294);
and U9372 (N_9372,N_9222,N_9261);
and U9373 (N_9373,N_9298,N_9210);
nand U9374 (N_9374,N_9240,N_9262);
or U9375 (N_9375,N_9295,N_9296);
nand U9376 (N_9376,N_9233,N_9270);
or U9377 (N_9377,N_9265,N_9251);
nand U9378 (N_9378,N_9206,N_9203);
or U9379 (N_9379,N_9233,N_9294);
nand U9380 (N_9380,N_9202,N_9271);
nand U9381 (N_9381,N_9286,N_9266);
and U9382 (N_9382,N_9294,N_9200);
and U9383 (N_9383,N_9291,N_9249);
or U9384 (N_9384,N_9200,N_9230);
nor U9385 (N_9385,N_9257,N_9264);
or U9386 (N_9386,N_9259,N_9220);
and U9387 (N_9387,N_9240,N_9227);
nor U9388 (N_9388,N_9252,N_9206);
nand U9389 (N_9389,N_9295,N_9227);
nor U9390 (N_9390,N_9273,N_9254);
and U9391 (N_9391,N_9258,N_9280);
nand U9392 (N_9392,N_9291,N_9204);
nand U9393 (N_9393,N_9285,N_9200);
nand U9394 (N_9394,N_9295,N_9228);
nand U9395 (N_9395,N_9225,N_9248);
nor U9396 (N_9396,N_9203,N_9295);
nor U9397 (N_9397,N_9223,N_9266);
and U9398 (N_9398,N_9241,N_9233);
or U9399 (N_9399,N_9219,N_9202);
and U9400 (N_9400,N_9354,N_9385);
nor U9401 (N_9401,N_9334,N_9342);
or U9402 (N_9402,N_9337,N_9318);
and U9403 (N_9403,N_9341,N_9368);
and U9404 (N_9404,N_9339,N_9352);
nand U9405 (N_9405,N_9358,N_9327);
and U9406 (N_9406,N_9335,N_9391);
and U9407 (N_9407,N_9393,N_9355);
or U9408 (N_9408,N_9367,N_9308);
or U9409 (N_9409,N_9311,N_9348);
and U9410 (N_9410,N_9300,N_9307);
or U9411 (N_9411,N_9374,N_9309);
or U9412 (N_9412,N_9366,N_9314);
or U9413 (N_9413,N_9330,N_9301);
xor U9414 (N_9414,N_9363,N_9323);
or U9415 (N_9415,N_9375,N_9353);
nor U9416 (N_9416,N_9395,N_9346);
and U9417 (N_9417,N_9361,N_9390);
nor U9418 (N_9418,N_9370,N_9382);
xnor U9419 (N_9419,N_9397,N_9356);
or U9420 (N_9420,N_9313,N_9324);
or U9421 (N_9421,N_9349,N_9321);
nand U9422 (N_9422,N_9359,N_9386);
nand U9423 (N_9423,N_9343,N_9317);
and U9424 (N_9424,N_9392,N_9365);
nand U9425 (N_9425,N_9340,N_9312);
nor U9426 (N_9426,N_9378,N_9399);
nor U9427 (N_9427,N_9364,N_9357);
nor U9428 (N_9428,N_9394,N_9331);
or U9429 (N_9429,N_9325,N_9302);
or U9430 (N_9430,N_9360,N_9388);
nor U9431 (N_9431,N_9338,N_9371);
nand U9432 (N_9432,N_9345,N_9319);
nor U9433 (N_9433,N_9379,N_9336);
nor U9434 (N_9434,N_9328,N_9373);
nor U9435 (N_9435,N_9383,N_9304);
or U9436 (N_9436,N_9347,N_9322);
and U9437 (N_9437,N_9305,N_9350);
or U9438 (N_9438,N_9315,N_9332);
and U9439 (N_9439,N_9387,N_9384);
nor U9440 (N_9440,N_9362,N_9381);
and U9441 (N_9441,N_9377,N_9316);
and U9442 (N_9442,N_9372,N_9376);
nor U9443 (N_9443,N_9389,N_9306);
or U9444 (N_9444,N_9380,N_9303);
or U9445 (N_9445,N_9369,N_9333);
nand U9446 (N_9446,N_9310,N_9351);
nor U9447 (N_9447,N_9320,N_9398);
nand U9448 (N_9448,N_9326,N_9344);
nor U9449 (N_9449,N_9396,N_9329);
and U9450 (N_9450,N_9319,N_9380);
or U9451 (N_9451,N_9310,N_9327);
or U9452 (N_9452,N_9376,N_9394);
and U9453 (N_9453,N_9380,N_9353);
nand U9454 (N_9454,N_9341,N_9354);
and U9455 (N_9455,N_9342,N_9394);
nand U9456 (N_9456,N_9372,N_9333);
nand U9457 (N_9457,N_9328,N_9319);
nor U9458 (N_9458,N_9380,N_9366);
and U9459 (N_9459,N_9390,N_9344);
or U9460 (N_9460,N_9337,N_9364);
and U9461 (N_9461,N_9354,N_9368);
and U9462 (N_9462,N_9306,N_9334);
and U9463 (N_9463,N_9377,N_9306);
nor U9464 (N_9464,N_9355,N_9326);
nor U9465 (N_9465,N_9329,N_9377);
nor U9466 (N_9466,N_9370,N_9362);
or U9467 (N_9467,N_9329,N_9312);
nor U9468 (N_9468,N_9394,N_9302);
nor U9469 (N_9469,N_9309,N_9362);
nor U9470 (N_9470,N_9338,N_9367);
or U9471 (N_9471,N_9372,N_9345);
and U9472 (N_9472,N_9382,N_9359);
or U9473 (N_9473,N_9373,N_9387);
or U9474 (N_9474,N_9308,N_9324);
and U9475 (N_9475,N_9336,N_9323);
and U9476 (N_9476,N_9342,N_9398);
or U9477 (N_9477,N_9384,N_9367);
nand U9478 (N_9478,N_9336,N_9364);
and U9479 (N_9479,N_9352,N_9375);
nor U9480 (N_9480,N_9375,N_9322);
and U9481 (N_9481,N_9342,N_9328);
or U9482 (N_9482,N_9346,N_9394);
or U9483 (N_9483,N_9367,N_9351);
or U9484 (N_9484,N_9362,N_9351);
nand U9485 (N_9485,N_9385,N_9340);
and U9486 (N_9486,N_9352,N_9300);
nand U9487 (N_9487,N_9368,N_9396);
and U9488 (N_9488,N_9382,N_9324);
nand U9489 (N_9489,N_9371,N_9353);
nand U9490 (N_9490,N_9342,N_9386);
nor U9491 (N_9491,N_9386,N_9355);
nand U9492 (N_9492,N_9322,N_9313);
nand U9493 (N_9493,N_9305,N_9360);
or U9494 (N_9494,N_9366,N_9335);
and U9495 (N_9495,N_9395,N_9336);
nor U9496 (N_9496,N_9319,N_9373);
and U9497 (N_9497,N_9390,N_9335);
nand U9498 (N_9498,N_9354,N_9330);
nor U9499 (N_9499,N_9350,N_9380);
nor U9500 (N_9500,N_9404,N_9427);
or U9501 (N_9501,N_9425,N_9466);
nand U9502 (N_9502,N_9492,N_9446);
nand U9503 (N_9503,N_9479,N_9423);
nand U9504 (N_9504,N_9429,N_9433);
or U9505 (N_9505,N_9449,N_9434);
nand U9506 (N_9506,N_9440,N_9421);
nand U9507 (N_9507,N_9412,N_9431);
nor U9508 (N_9508,N_9459,N_9467);
and U9509 (N_9509,N_9430,N_9444);
nor U9510 (N_9510,N_9435,N_9471);
nor U9511 (N_9511,N_9491,N_9438);
or U9512 (N_9512,N_9489,N_9483);
nand U9513 (N_9513,N_9481,N_9439);
nand U9514 (N_9514,N_9487,N_9484);
nand U9515 (N_9515,N_9402,N_9415);
nor U9516 (N_9516,N_9473,N_9443);
nand U9517 (N_9517,N_9441,N_9419);
nand U9518 (N_9518,N_9442,N_9445);
nand U9519 (N_9519,N_9410,N_9432);
nor U9520 (N_9520,N_9454,N_9496);
nor U9521 (N_9521,N_9428,N_9414);
nand U9522 (N_9522,N_9448,N_9405);
nor U9523 (N_9523,N_9436,N_9458);
and U9524 (N_9524,N_9453,N_9462);
nand U9525 (N_9525,N_9470,N_9499);
or U9526 (N_9526,N_9411,N_9424);
nand U9527 (N_9527,N_9472,N_9416);
or U9528 (N_9528,N_9408,N_9403);
nand U9529 (N_9529,N_9498,N_9460);
nand U9530 (N_9530,N_9455,N_9464);
nor U9531 (N_9531,N_9478,N_9486);
nor U9532 (N_9532,N_9409,N_9422);
xnor U9533 (N_9533,N_9463,N_9477);
nand U9534 (N_9534,N_9401,N_9493);
nand U9535 (N_9535,N_9474,N_9497);
or U9536 (N_9536,N_9456,N_9452);
nor U9537 (N_9537,N_9475,N_9468);
nand U9538 (N_9538,N_9420,N_9469);
nor U9539 (N_9539,N_9457,N_9495);
or U9540 (N_9540,N_9465,N_9451);
and U9541 (N_9541,N_9485,N_9482);
and U9542 (N_9542,N_9461,N_9407);
and U9543 (N_9543,N_9476,N_9488);
nor U9544 (N_9544,N_9490,N_9447);
and U9545 (N_9545,N_9417,N_9418);
and U9546 (N_9546,N_9450,N_9437);
nor U9547 (N_9547,N_9426,N_9494);
and U9548 (N_9548,N_9400,N_9480);
xnor U9549 (N_9549,N_9406,N_9413);
nand U9550 (N_9550,N_9420,N_9482);
nand U9551 (N_9551,N_9453,N_9455);
nor U9552 (N_9552,N_9497,N_9446);
nor U9553 (N_9553,N_9476,N_9403);
nand U9554 (N_9554,N_9429,N_9450);
or U9555 (N_9555,N_9445,N_9406);
and U9556 (N_9556,N_9415,N_9490);
and U9557 (N_9557,N_9421,N_9477);
or U9558 (N_9558,N_9470,N_9491);
or U9559 (N_9559,N_9414,N_9427);
or U9560 (N_9560,N_9497,N_9447);
nand U9561 (N_9561,N_9483,N_9462);
nor U9562 (N_9562,N_9493,N_9464);
nand U9563 (N_9563,N_9495,N_9413);
nand U9564 (N_9564,N_9449,N_9431);
nand U9565 (N_9565,N_9458,N_9459);
and U9566 (N_9566,N_9498,N_9476);
or U9567 (N_9567,N_9437,N_9422);
nor U9568 (N_9568,N_9445,N_9440);
nor U9569 (N_9569,N_9449,N_9401);
and U9570 (N_9570,N_9422,N_9465);
nand U9571 (N_9571,N_9415,N_9483);
nor U9572 (N_9572,N_9406,N_9468);
nor U9573 (N_9573,N_9428,N_9476);
nor U9574 (N_9574,N_9461,N_9438);
and U9575 (N_9575,N_9473,N_9416);
nor U9576 (N_9576,N_9402,N_9477);
nand U9577 (N_9577,N_9428,N_9411);
or U9578 (N_9578,N_9470,N_9444);
and U9579 (N_9579,N_9431,N_9447);
nor U9580 (N_9580,N_9478,N_9401);
or U9581 (N_9581,N_9493,N_9463);
nor U9582 (N_9582,N_9482,N_9496);
nor U9583 (N_9583,N_9469,N_9485);
nor U9584 (N_9584,N_9445,N_9401);
nor U9585 (N_9585,N_9426,N_9408);
or U9586 (N_9586,N_9496,N_9464);
nand U9587 (N_9587,N_9496,N_9474);
and U9588 (N_9588,N_9456,N_9422);
nand U9589 (N_9589,N_9453,N_9448);
or U9590 (N_9590,N_9425,N_9405);
or U9591 (N_9591,N_9449,N_9457);
nor U9592 (N_9592,N_9483,N_9412);
nand U9593 (N_9593,N_9428,N_9495);
nand U9594 (N_9594,N_9494,N_9443);
nor U9595 (N_9595,N_9441,N_9436);
or U9596 (N_9596,N_9435,N_9484);
nor U9597 (N_9597,N_9411,N_9416);
nand U9598 (N_9598,N_9426,N_9406);
and U9599 (N_9599,N_9409,N_9477);
or U9600 (N_9600,N_9523,N_9588);
nand U9601 (N_9601,N_9511,N_9570);
and U9602 (N_9602,N_9598,N_9577);
and U9603 (N_9603,N_9525,N_9581);
and U9604 (N_9604,N_9593,N_9555);
or U9605 (N_9605,N_9556,N_9596);
and U9606 (N_9606,N_9502,N_9595);
and U9607 (N_9607,N_9564,N_9584);
nor U9608 (N_9608,N_9582,N_9500);
nand U9609 (N_9609,N_9566,N_9513);
nand U9610 (N_9610,N_9547,N_9571);
nor U9611 (N_9611,N_9501,N_9552);
or U9612 (N_9612,N_9516,N_9515);
and U9613 (N_9613,N_9507,N_9548);
nor U9614 (N_9614,N_9569,N_9544);
and U9615 (N_9615,N_9509,N_9542);
nor U9616 (N_9616,N_9533,N_9559);
nand U9617 (N_9617,N_9560,N_9578);
and U9618 (N_9618,N_9554,N_9528);
and U9619 (N_9619,N_9541,N_9522);
and U9620 (N_9620,N_9535,N_9504);
or U9621 (N_9621,N_9532,N_9585);
or U9622 (N_9622,N_9565,N_9592);
nand U9623 (N_9623,N_9530,N_9583);
or U9624 (N_9624,N_9574,N_9568);
nor U9625 (N_9625,N_9540,N_9539);
nor U9626 (N_9626,N_9576,N_9520);
or U9627 (N_9627,N_9546,N_9567);
xnor U9628 (N_9628,N_9557,N_9517);
and U9629 (N_9629,N_9597,N_9537);
nand U9630 (N_9630,N_9586,N_9590);
or U9631 (N_9631,N_9503,N_9579);
nand U9632 (N_9632,N_9589,N_9550);
nor U9633 (N_9633,N_9587,N_9591);
nor U9634 (N_9634,N_9524,N_9562);
or U9635 (N_9635,N_9519,N_9512);
nand U9636 (N_9636,N_9506,N_9551);
nand U9637 (N_9637,N_9599,N_9531);
and U9638 (N_9638,N_9514,N_9573);
and U9639 (N_9639,N_9529,N_9575);
and U9640 (N_9640,N_9572,N_9545);
nand U9641 (N_9641,N_9536,N_9521);
and U9642 (N_9642,N_9510,N_9526);
nand U9643 (N_9643,N_9580,N_9508);
nand U9644 (N_9644,N_9549,N_9561);
xnor U9645 (N_9645,N_9518,N_9543);
and U9646 (N_9646,N_9534,N_9558);
and U9647 (N_9647,N_9527,N_9505);
nor U9648 (N_9648,N_9563,N_9538);
and U9649 (N_9649,N_9553,N_9594);
or U9650 (N_9650,N_9516,N_9548);
nand U9651 (N_9651,N_9551,N_9546);
nand U9652 (N_9652,N_9508,N_9567);
and U9653 (N_9653,N_9572,N_9501);
nand U9654 (N_9654,N_9591,N_9525);
or U9655 (N_9655,N_9576,N_9541);
and U9656 (N_9656,N_9542,N_9527);
nor U9657 (N_9657,N_9570,N_9578);
or U9658 (N_9658,N_9592,N_9507);
nand U9659 (N_9659,N_9570,N_9509);
nand U9660 (N_9660,N_9518,N_9547);
nand U9661 (N_9661,N_9594,N_9540);
nor U9662 (N_9662,N_9554,N_9589);
nor U9663 (N_9663,N_9526,N_9551);
and U9664 (N_9664,N_9563,N_9542);
or U9665 (N_9665,N_9531,N_9549);
or U9666 (N_9666,N_9566,N_9528);
or U9667 (N_9667,N_9513,N_9519);
nor U9668 (N_9668,N_9577,N_9590);
nor U9669 (N_9669,N_9533,N_9558);
nand U9670 (N_9670,N_9521,N_9595);
or U9671 (N_9671,N_9593,N_9542);
nand U9672 (N_9672,N_9500,N_9520);
nand U9673 (N_9673,N_9523,N_9508);
or U9674 (N_9674,N_9541,N_9564);
nand U9675 (N_9675,N_9506,N_9516);
or U9676 (N_9676,N_9539,N_9511);
nand U9677 (N_9677,N_9577,N_9571);
nor U9678 (N_9678,N_9525,N_9577);
or U9679 (N_9679,N_9595,N_9524);
and U9680 (N_9680,N_9580,N_9592);
nand U9681 (N_9681,N_9533,N_9564);
nor U9682 (N_9682,N_9550,N_9580);
nor U9683 (N_9683,N_9586,N_9553);
nand U9684 (N_9684,N_9556,N_9567);
and U9685 (N_9685,N_9509,N_9552);
and U9686 (N_9686,N_9553,N_9540);
or U9687 (N_9687,N_9565,N_9575);
nor U9688 (N_9688,N_9535,N_9580);
nand U9689 (N_9689,N_9577,N_9581);
or U9690 (N_9690,N_9502,N_9570);
nor U9691 (N_9691,N_9572,N_9534);
or U9692 (N_9692,N_9575,N_9571);
nand U9693 (N_9693,N_9591,N_9546);
nand U9694 (N_9694,N_9520,N_9509);
and U9695 (N_9695,N_9565,N_9579);
nand U9696 (N_9696,N_9573,N_9560);
and U9697 (N_9697,N_9537,N_9514);
nor U9698 (N_9698,N_9573,N_9547);
or U9699 (N_9699,N_9505,N_9535);
nor U9700 (N_9700,N_9681,N_9686);
nand U9701 (N_9701,N_9683,N_9699);
or U9702 (N_9702,N_9606,N_9632);
nand U9703 (N_9703,N_9688,N_9641);
and U9704 (N_9704,N_9690,N_9633);
and U9705 (N_9705,N_9660,N_9623);
and U9706 (N_9706,N_9685,N_9682);
or U9707 (N_9707,N_9616,N_9665);
nand U9708 (N_9708,N_9687,N_9671);
nand U9709 (N_9709,N_9658,N_9610);
nor U9710 (N_9710,N_9614,N_9611);
and U9711 (N_9711,N_9664,N_9675);
nor U9712 (N_9712,N_9629,N_9639);
and U9713 (N_9713,N_9692,N_9693);
nand U9714 (N_9714,N_9697,N_9654);
nand U9715 (N_9715,N_9627,N_9622);
and U9716 (N_9716,N_9646,N_9647);
nand U9717 (N_9717,N_9618,N_9684);
and U9718 (N_9718,N_9696,N_9670);
nor U9719 (N_9719,N_9676,N_9624);
nand U9720 (N_9720,N_9645,N_9640);
nand U9721 (N_9721,N_9636,N_9634);
nand U9722 (N_9722,N_9656,N_9638);
nor U9723 (N_9723,N_9642,N_9631);
or U9724 (N_9724,N_9678,N_9653);
and U9725 (N_9725,N_9619,N_9600);
and U9726 (N_9726,N_9628,N_9626);
or U9727 (N_9727,N_9609,N_9672);
nand U9728 (N_9728,N_9674,N_9635);
and U9729 (N_9729,N_9603,N_9637);
nor U9730 (N_9730,N_9602,N_9621);
and U9731 (N_9731,N_9607,N_9617);
nand U9732 (N_9732,N_9661,N_9650);
or U9733 (N_9733,N_9613,N_9698);
nor U9734 (N_9734,N_9657,N_9673);
and U9735 (N_9735,N_9677,N_9663);
nand U9736 (N_9736,N_9608,N_9648);
nand U9737 (N_9737,N_9666,N_9643);
nor U9738 (N_9738,N_9604,N_9605);
nor U9739 (N_9739,N_9669,N_9662);
and U9740 (N_9740,N_9644,N_9667);
nand U9741 (N_9741,N_9680,N_9630);
and U9742 (N_9742,N_9679,N_9659);
or U9743 (N_9743,N_9668,N_9649);
or U9744 (N_9744,N_9651,N_9655);
or U9745 (N_9745,N_9615,N_9601);
nand U9746 (N_9746,N_9694,N_9691);
nand U9747 (N_9747,N_9625,N_9689);
nor U9748 (N_9748,N_9652,N_9695);
or U9749 (N_9749,N_9612,N_9620);
or U9750 (N_9750,N_9663,N_9661);
nor U9751 (N_9751,N_9649,N_9685);
nand U9752 (N_9752,N_9650,N_9627);
and U9753 (N_9753,N_9640,N_9609);
nor U9754 (N_9754,N_9681,N_9689);
nor U9755 (N_9755,N_9673,N_9604);
nor U9756 (N_9756,N_9643,N_9694);
and U9757 (N_9757,N_9659,N_9670);
nand U9758 (N_9758,N_9698,N_9600);
nand U9759 (N_9759,N_9616,N_9606);
or U9760 (N_9760,N_9646,N_9682);
nand U9761 (N_9761,N_9618,N_9638);
nand U9762 (N_9762,N_9620,N_9622);
nor U9763 (N_9763,N_9630,N_9678);
nor U9764 (N_9764,N_9679,N_9687);
nand U9765 (N_9765,N_9698,N_9635);
nor U9766 (N_9766,N_9687,N_9635);
and U9767 (N_9767,N_9686,N_9602);
nand U9768 (N_9768,N_9613,N_9654);
nor U9769 (N_9769,N_9643,N_9685);
and U9770 (N_9770,N_9687,N_9623);
and U9771 (N_9771,N_9617,N_9638);
nor U9772 (N_9772,N_9618,N_9644);
or U9773 (N_9773,N_9634,N_9617);
nor U9774 (N_9774,N_9658,N_9611);
or U9775 (N_9775,N_9631,N_9656);
nor U9776 (N_9776,N_9655,N_9635);
nand U9777 (N_9777,N_9687,N_9673);
nor U9778 (N_9778,N_9691,N_9605);
nor U9779 (N_9779,N_9625,N_9631);
nand U9780 (N_9780,N_9676,N_9625);
nor U9781 (N_9781,N_9632,N_9652);
nor U9782 (N_9782,N_9603,N_9627);
nand U9783 (N_9783,N_9627,N_9684);
or U9784 (N_9784,N_9691,N_9624);
and U9785 (N_9785,N_9688,N_9610);
or U9786 (N_9786,N_9621,N_9613);
nand U9787 (N_9787,N_9645,N_9666);
nor U9788 (N_9788,N_9617,N_9682);
nor U9789 (N_9789,N_9627,N_9669);
and U9790 (N_9790,N_9628,N_9612);
nand U9791 (N_9791,N_9665,N_9698);
or U9792 (N_9792,N_9666,N_9676);
nand U9793 (N_9793,N_9623,N_9647);
nand U9794 (N_9794,N_9670,N_9618);
nand U9795 (N_9795,N_9686,N_9664);
nor U9796 (N_9796,N_9604,N_9648);
nand U9797 (N_9797,N_9673,N_9651);
nand U9798 (N_9798,N_9655,N_9647);
nand U9799 (N_9799,N_9684,N_9626);
or U9800 (N_9800,N_9765,N_9780);
and U9801 (N_9801,N_9710,N_9794);
nor U9802 (N_9802,N_9767,N_9729);
and U9803 (N_9803,N_9778,N_9733);
nor U9804 (N_9804,N_9738,N_9745);
or U9805 (N_9805,N_9726,N_9747);
and U9806 (N_9806,N_9749,N_9753);
nor U9807 (N_9807,N_9748,N_9713);
nor U9808 (N_9808,N_9793,N_9706);
or U9809 (N_9809,N_9740,N_9708);
nand U9810 (N_9810,N_9715,N_9762);
and U9811 (N_9811,N_9757,N_9755);
or U9812 (N_9812,N_9720,N_9707);
or U9813 (N_9813,N_9797,N_9776);
or U9814 (N_9814,N_9704,N_9705);
or U9815 (N_9815,N_9786,N_9773);
or U9816 (N_9816,N_9724,N_9790);
or U9817 (N_9817,N_9787,N_9791);
and U9818 (N_9818,N_9766,N_9744);
and U9819 (N_9819,N_9758,N_9752);
and U9820 (N_9820,N_9742,N_9711);
nand U9821 (N_9821,N_9741,N_9763);
nand U9822 (N_9822,N_9795,N_9727);
nand U9823 (N_9823,N_9764,N_9700);
nand U9824 (N_9824,N_9788,N_9712);
xor U9825 (N_9825,N_9723,N_9722);
and U9826 (N_9826,N_9734,N_9784);
or U9827 (N_9827,N_9731,N_9789);
and U9828 (N_9828,N_9701,N_9772);
or U9829 (N_9829,N_9768,N_9775);
and U9830 (N_9830,N_9702,N_9751);
and U9831 (N_9831,N_9779,N_9739);
or U9832 (N_9832,N_9756,N_9732);
and U9833 (N_9833,N_9716,N_9709);
nor U9834 (N_9834,N_9719,N_9777);
or U9835 (N_9835,N_9728,N_9730);
or U9836 (N_9836,N_9783,N_9714);
nor U9837 (N_9837,N_9759,N_9774);
and U9838 (N_9838,N_9781,N_9798);
nor U9839 (N_9839,N_9760,N_9769);
nor U9840 (N_9840,N_9721,N_9718);
nand U9841 (N_9841,N_9736,N_9771);
or U9842 (N_9842,N_9725,N_9717);
nor U9843 (N_9843,N_9754,N_9792);
and U9844 (N_9844,N_9782,N_9735);
and U9845 (N_9845,N_9703,N_9737);
nor U9846 (N_9846,N_9761,N_9799);
nand U9847 (N_9847,N_9796,N_9750);
and U9848 (N_9848,N_9785,N_9770);
nor U9849 (N_9849,N_9743,N_9746);
xnor U9850 (N_9850,N_9792,N_9751);
nand U9851 (N_9851,N_9720,N_9730);
and U9852 (N_9852,N_9784,N_9708);
nand U9853 (N_9853,N_9719,N_9754);
nor U9854 (N_9854,N_9795,N_9781);
or U9855 (N_9855,N_9770,N_9745);
nand U9856 (N_9856,N_9790,N_9747);
nor U9857 (N_9857,N_9715,N_9757);
nand U9858 (N_9858,N_9757,N_9710);
or U9859 (N_9859,N_9743,N_9768);
and U9860 (N_9860,N_9734,N_9711);
nor U9861 (N_9861,N_9782,N_9751);
nor U9862 (N_9862,N_9737,N_9716);
nand U9863 (N_9863,N_9741,N_9799);
nand U9864 (N_9864,N_9731,N_9777);
nand U9865 (N_9865,N_9747,N_9770);
and U9866 (N_9866,N_9749,N_9708);
nor U9867 (N_9867,N_9772,N_9775);
or U9868 (N_9868,N_9734,N_9760);
nor U9869 (N_9869,N_9709,N_9794);
or U9870 (N_9870,N_9716,N_9750);
and U9871 (N_9871,N_9754,N_9750);
nand U9872 (N_9872,N_9734,N_9793);
or U9873 (N_9873,N_9724,N_9762);
or U9874 (N_9874,N_9749,N_9710);
and U9875 (N_9875,N_9782,N_9778);
and U9876 (N_9876,N_9734,N_9792);
and U9877 (N_9877,N_9784,N_9781);
and U9878 (N_9878,N_9714,N_9737);
nand U9879 (N_9879,N_9792,N_9729);
nor U9880 (N_9880,N_9751,N_9799);
xor U9881 (N_9881,N_9796,N_9763);
nor U9882 (N_9882,N_9711,N_9704);
nand U9883 (N_9883,N_9727,N_9763);
or U9884 (N_9884,N_9752,N_9729);
nand U9885 (N_9885,N_9773,N_9798);
and U9886 (N_9886,N_9722,N_9792);
nor U9887 (N_9887,N_9749,N_9740);
and U9888 (N_9888,N_9737,N_9700);
nor U9889 (N_9889,N_9730,N_9710);
nand U9890 (N_9890,N_9786,N_9768);
or U9891 (N_9891,N_9784,N_9706);
nor U9892 (N_9892,N_9759,N_9724);
and U9893 (N_9893,N_9724,N_9764);
and U9894 (N_9894,N_9741,N_9797);
nand U9895 (N_9895,N_9714,N_9745);
nor U9896 (N_9896,N_9774,N_9712);
nor U9897 (N_9897,N_9731,N_9747);
or U9898 (N_9898,N_9731,N_9708);
nor U9899 (N_9899,N_9753,N_9786);
nor U9900 (N_9900,N_9835,N_9866);
nor U9901 (N_9901,N_9814,N_9826);
or U9902 (N_9902,N_9810,N_9854);
or U9903 (N_9903,N_9857,N_9892);
nand U9904 (N_9904,N_9894,N_9834);
nand U9905 (N_9905,N_9811,N_9885);
nand U9906 (N_9906,N_9816,N_9805);
nor U9907 (N_9907,N_9895,N_9869);
or U9908 (N_9908,N_9872,N_9846);
nand U9909 (N_9909,N_9878,N_9898);
nand U9910 (N_9910,N_9874,N_9877);
xor U9911 (N_9911,N_9882,N_9889);
nand U9912 (N_9912,N_9848,N_9838);
xnor U9913 (N_9913,N_9890,N_9815);
nand U9914 (N_9914,N_9853,N_9860);
nor U9915 (N_9915,N_9886,N_9803);
nor U9916 (N_9916,N_9808,N_9824);
or U9917 (N_9917,N_9847,N_9828);
or U9918 (N_9918,N_9812,N_9820);
and U9919 (N_9919,N_9855,N_9841);
nor U9920 (N_9920,N_9825,N_9842);
and U9921 (N_9921,N_9884,N_9821);
nor U9922 (N_9922,N_9896,N_9802);
nand U9923 (N_9923,N_9875,N_9862);
nand U9924 (N_9924,N_9806,N_9876);
nor U9925 (N_9925,N_9817,N_9888);
nor U9926 (N_9926,N_9840,N_9823);
and U9927 (N_9927,N_9809,N_9863);
or U9928 (N_9928,N_9883,N_9880);
and U9929 (N_9929,N_9856,N_9858);
xor U9930 (N_9930,N_9868,N_9851);
nand U9931 (N_9931,N_9800,N_9844);
and U9932 (N_9932,N_9870,N_9879);
and U9933 (N_9933,N_9801,N_9827);
nor U9934 (N_9934,N_9897,N_9832);
or U9935 (N_9935,N_9871,N_9813);
nor U9936 (N_9936,N_9887,N_9891);
and U9937 (N_9937,N_9833,N_9899);
nor U9938 (N_9938,N_9843,N_9836);
xor U9939 (N_9939,N_9861,N_9865);
nor U9940 (N_9940,N_9839,N_9804);
or U9941 (N_9941,N_9873,N_9831);
nor U9942 (N_9942,N_9837,N_9819);
nor U9943 (N_9943,N_9829,N_9850);
or U9944 (N_9944,N_9822,N_9859);
nand U9945 (N_9945,N_9807,N_9852);
xor U9946 (N_9946,N_9881,N_9845);
nand U9947 (N_9947,N_9867,N_9818);
nor U9948 (N_9948,N_9830,N_9893);
nor U9949 (N_9949,N_9849,N_9864);
and U9950 (N_9950,N_9867,N_9872);
nand U9951 (N_9951,N_9882,N_9802);
or U9952 (N_9952,N_9863,N_9893);
or U9953 (N_9953,N_9833,N_9839);
nand U9954 (N_9954,N_9803,N_9836);
xor U9955 (N_9955,N_9875,N_9866);
nor U9956 (N_9956,N_9881,N_9891);
nand U9957 (N_9957,N_9885,N_9829);
and U9958 (N_9958,N_9855,N_9835);
nor U9959 (N_9959,N_9865,N_9843);
nand U9960 (N_9960,N_9862,N_9803);
nand U9961 (N_9961,N_9883,N_9896);
nand U9962 (N_9962,N_9861,N_9825);
nor U9963 (N_9963,N_9889,N_9825);
nor U9964 (N_9964,N_9863,N_9816);
and U9965 (N_9965,N_9848,N_9822);
nor U9966 (N_9966,N_9899,N_9836);
or U9967 (N_9967,N_9840,N_9864);
nand U9968 (N_9968,N_9889,N_9810);
nand U9969 (N_9969,N_9850,N_9853);
nand U9970 (N_9970,N_9841,N_9852);
nor U9971 (N_9971,N_9825,N_9836);
and U9972 (N_9972,N_9819,N_9835);
xor U9973 (N_9973,N_9817,N_9827);
or U9974 (N_9974,N_9849,N_9800);
and U9975 (N_9975,N_9881,N_9841);
or U9976 (N_9976,N_9872,N_9842);
and U9977 (N_9977,N_9874,N_9873);
and U9978 (N_9978,N_9843,N_9862);
nand U9979 (N_9979,N_9875,N_9863);
nand U9980 (N_9980,N_9840,N_9854);
nor U9981 (N_9981,N_9832,N_9889);
and U9982 (N_9982,N_9893,N_9835);
nand U9983 (N_9983,N_9810,N_9804);
nor U9984 (N_9984,N_9849,N_9801);
nand U9985 (N_9985,N_9862,N_9871);
or U9986 (N_9986,N_9856,N_9860);
and U9987 (N_9987,N_9898,N_9825);
nor U9988 (N_9988,N_9814,N_9883);
nor U9989 (N_9989,N_9887,N_9805);
and U9990 (N_9990,N_9899,N_9840);
or U9991 (N_9991,N_9895,N_9814);
nand U9992 (N_9992,N_9858,N_9861);
nor U9993 (N_9993,N_9852,N_9879);
nand U9994 (N_9994,N_9831,N_9889);
nor U9995 (N_9995,N_9893,N_9853);
nor U9996 (N_9996,N_9808,N_9859);
nand U9997 (N_9997,N_9809,N_9839);
nand U9998 (N_9998,N_9804,N_9855);
nand U9999 (N_9999,N_9864,N_9848);
or UO_0 (O_0,N_9972,N_9930);
nand UO_1 (O_1,N_9988,N_9955);
or UO_2 (O_2,N_9941,N_9984);
nor UO_3 (O_3,N_9912,N_9938);
and UO_4 (O_4,N_9917,N_9973);
nor UO_5 (O_5,N_9965,N_9933);
and UO_6 (O_6,N_9991,N_9925);
nor UO_7 (O_7,N_9992,N_9944);
nor UO_8 (O_8,N_9952,N_9945);
nand UO_9 (O_9,N_9922,N_9910);
nand UO_10 (O_10,N_9985,N_9974);
or UO_11 (O_11,N_9977,N_9915);
nand UO_12 (O_12,N_9936,N_9964);
and UO_13 (O_13,N_9946,N_9975);
or UO_14 (O_14,N_9926,N_9932);
nand UO_15 (O_15,N_9949,N_9943);
nor UO_16 (O_16,N_9929,N_9923);
and UO_17 (O_17,N_9971,N_9942);
nor UO_18 (O_18,N_9914,N_9959);
nor UO_19 (O_19,N_9948,N_9968);
and UO_20 (O_20,N_9919,N_9905);
nor UO_21 (O_21,N_9913,N_9990);
nor UO_22 (O_22,N_9969,N_9983);
nor UO_23 (O_23,N_9993,N_9961);
and UO_24 (O_24,N_9994,N_9921);
nand UO_25 (O_25,N_9940,N_9934);
and UO_26 (O_26,N_9967,N_9957);
or UO_27 (O_27,N_9906,N_9997);
and UO_28 (O_28,N_9982,N_9995);
nand UO_29 (O_29,N_9978,N_9950);
or UO_30 (O_30,N_9962,N_9939);
and UO_31 (O_31,N_9947,N_9928);
or UO_32 (O_32,N_9903,N_9986);
and UO_33 (O_33,N_9902,N_9901);
or UO_34 (O_34,N_9920,N_9908);
nand UO_35 (O_35,N_9963,N_9907);
nand UO_36 (O_36,N_9911,N_9956);
nand UO_37 (O_37,N_9987,N_9998);
and UO_38 (O_38,N_9999,N_9953);
nor UO_39 (O_39,N_9951,N_9918);
nor UO_40 (O_40,N_9989,N_9979);
or UO_41 (O_41,N_9996,N_9909);
or UO_42 (O_42,N_9966,N_9935);
or UO_43 (O_43,N_9937,N_9976);
nor UO_44 (O_44,N_9960,N_9904);
nor UO_45 (O_45,N_9924,N_9931);
nand UO_46 (O_46,N_9954,N_9958);
and UO_47 (O_47,N_9900,N_9980);
and UO_48 (O_48,N_9927,N_9916);
nand UO_49 (O_49,N_9981,N_9970);
nand UO_50 (O_50,N_9966,N_9946);
or UO_51 (O_51,N_9991,N_9958);
nor UO_52 (O_52,N_9983,N_9920);
or UO_53 (O_53,N_9927,N_9921);
or UO_54 (O_54,N_9932,N_9967);
nand UO_55 (O_55,N_9958,N_9900);
nand UO_56 (O_56,N_9979,N_9954);
or UO_57 (O_57,N_9971,N_9907);
and UO_58 (O_58,N_9937,N_9936);
nand UO_59 (O_59,N_9932,N_9909);
nor UO_60 (O_60,N_9943,N_9914);
nor UO_61 (O_61,N_9938,N_9910);
or UO_62 (O_62,N_9978,N_9934);
nand UO_63 (O_63,N_9975,N_9935);
and UO_64 (O_64,N_9911,N_9965);
nand UO_65 (O_65,N_9928,N_9966);
nand UO_66 (O_66,N_9966,N_9975);
nor UO_67 (O_67,N_9942,N_9922);
nor UO_68 (O_68,N_9985,N_9952);
or UO_69 (O_69,N_9900,N_9911);
nand UO_70 (O_70,N_9944,N_9993);
nor UO_71 (O_71,N_9967,N_9901);
nand UO_72 (O_72,N_9972,N_9969);
nand UO_73 (O_73,N_9998,N_9954);
or UO_74 (O_74,N_9924,N_9918);
nand UO_75 (O_75,N_9919,N_9927);
nand UO_76 (O_76,N_9906,N_9931);
nor UO_77 (O_77,N_9913,N_9960);
nand UO_78 (O_78,N_9909,N_9931);
nor UO_79 (O_79,N_9960,N_9959);
and UO_80 (O_80,N_9977,N_9949);
nor UO_81 (O_81,N_9941,N_9983);
or UO_82 (O_82,N_9973,N_9954);
xor UO_83 (O_83,N_9903,N_9909);
or UO_84 (O_84,N_9960,N_9928);
nor UO_85 (O_85,N_9954,N_9911);
nand UO_86 (O_86,N_9987,N_9989);
nand UO_87 (O_87,N_9956,N_9975);
or UO_88 (O_88,N_9914,N_9993);
or UO_89 (O_89,N_9971,N_9925);
nand UO_90 (O_90,N_9966,N_9909);
or UO_91 (O_91,N_9923,N_9915);
nor UO_92 (O_92,N_9931,N_9997);
xor UO_93 (O_93,N_9924,N_9903);
nand UO_94 (O_94,N_9924,N_9913);
or UO_95 (O_95,N_9903,N_9947);
and UO_96 (O_96,N_9949,N_9961);
and UO_97 (O_97,N_9923,N_9920);
nor UO_98 (O_98,N_9921,N_9967);
nor UO_99 (O_99,N_9917,N_9953);
or UO_100 (O_100,N_9960,N_9927);
nor UO_101 (O_101,N_9902,N_9946);
and UO_102 (O_102,N_9964,N_9946);
nand UO_103 (O_103,N_9914,N_9977);
nand UO_104 (O_104,N_9967,N_9935);
nor UO_105 (O_105,N_9937,N_9962);
or UO_106 (O_106,N_9963,N_9902);
and UO_107 (O_107,N_9965,N_9914);
nand UO_108 (O_108,N_9949,N_9956);
and UO_109 (O_109,N_9902,N_9976);
or UO_110 (O_110,N_9917,N_9940);
nand UO_111 (O_111,N_9941,N_9958);
and UO_112 (O_112,N_9934,N_9933);
or UO_113 (O_113,N_9985,N_9975);
nor UO_114 (O_114,N_9932,N_9942);
nor UO_115 (O_115,N_9999,N_9963);
or UO_116 (O_116,N_9949,N_9918);
and UO_117 (O_117,N_9912,N_9999);
nor UO_118 (O_118,N_9985,N_9940);
nand UO_119 (O_119,N_9945,N_9918);
and UO_120 (O_120,N_9914,N_9970);
nand UO_121 (O_121,N_9999,N_9930);
nor UO_122 (O_122,N_9998,N_9931);
or UO_123 (O_123,N_9940,N_9933);
nor UO_124 (O_124,N_9992,N_9947);
or UO_125 (O_125,N_9961,N_9957);
nand UO_126 (O_126,N_9959,N_9955);
or UO_127 (O_127,N_9968,N_9913);
or UO_128 (O_128,N_9991,N_9941);
or UO_129 (O_129,N_9966,N_9924);
or UO_130 (O_130,N_9903,N_9945);
nor UO_131 (O_131,N_9918,N_9914);
and UO_132 (O_132,N_9945,N_9941);
nor UO_133 (O_133,N_9914,N_9979);
nand UO_134 (O_134,N_9960,N_9985);
or UO_135 (O_135,N_9998,N_9910);
and UO_136 (O_136,N_9933,N_9926);
and UO_137 (O_137,N_9907,N_9999);
nor UO_138 (O_138,N_9927,N_9957);
or UO_139 (O_139,N_9918,N_9965);
or UO_140 (O_140,N_9940,N_9984);
nand UO_141 (O_141,N_9903,N_9910);
or UO_142 (O_142,N_9974,N_9956);
and UO_143 (O_143,N_9967,N_9991);
and UO_144 (O_144,N_9929,N_9993);
nor UO_145 (O_145,N_9967,N_9913);
or UO_146 (O_146,N_9930,N_9954);
or UO_147 (O_147,N_9934,N_9941);
and UO_148 (O_148,N_9924,N_9939);
nand UO_149 (O_149,N_9925,N_9977);
and UO_150 (O_150,N_9961,N_9918);
or UO_151 (O_151,N_9957,N_9985);
and UO_152 (O_152,N_9971,N_9951);
and UO_153 (O_153,N_9904,N_9934);
and UO_154 (O_154,N_9984,N_9950);
and UO_155 (O_155,N_9946,N_9900);
nand UO_156 (O_156,N_9948,N_9956);
nor UO_157 (O_157,N_9964,N_9976);
nor UO_158 (O_158,N_9941,N_9970);
and UO_159 (O_159,N_9991,N_9959);
nor UO_160 (O_160,N_9971,N_9984);
nor UO_161 (O_161,N_9989,N_9983);
nor UO_162 (O_162,N_9926,N_9920);
and UO_163 (O_163,N_9937,N_9998);
nand UO_164 (O_164,N_9926,N_9978);
or UO_165 (O_165,N_9983,N_9934);
nand UO_166 (O_166,N_9940,N_9944);
or UO_167 (O_167,N_9902,N_9986);
and UO_168 (O_168,N_9957,N_9901);
or UO_169 (O_169,N_9984,N_9923);
and UO_170 (O_170,N_9940,N_9981);
nand UO_171 (O_171,N_9930,N_9990);
and UO_172 (O_172,N_9996,N_9952);
or UO_173 (O_173,N_9950,N_9998);
and UO_174 (O_174,N_9988,N_9939);
nand UO_175 (O_175,N_9980,N_9975);
nor UO_176 (O_176,N_9968,N_9964);
and UO_177 (O_177,N_9905,N_9984);
nand UO_178 (O_178,N_9945,N_9986);
nand UO_179 (O_179,N_9980,N_9983);
xnor UO_180 (O_180,N_9999,N_9968);
nand UO_181 (O_181,N_9915,N_9963);
nand UO_182 (O_182,N_9996,N_9959);
nor UO_183 (O_183,N_9969,N_9913);
and UO_184 (O_184,N_9970,N_9924);
nor UO_185 (O_185,N_9908,N_9989);
and UO_186 (O_186,N_9930,N_9953);
or UO_187 (O_187,N_9901,N_9996);
nand UO_188 (O_188,N_9989,N_9929);
xor UO_189 (O_189,N_9911,N_9972);
nand UO_190 (O_190,N_9965,N_9940);
nor UO_191 (O_191,N_9945,N_9937);
or UO_192 (O_192,N_9955,N_9929);
nor UO_193 (O_193,N_9930,N_9945);
nor UO_194 (O_194,N_9951,N_9974);
or UO_195 (O_195,N_9959,N_9994);
or UO_196 (O_196,N_9984,N_9987);
nand UO_197 (O_197,N_9918,N_9931);
nand UO_198 (O_198,N_9932,N_9976);
nand UO_199 (O_199,N_9987,N_9944);
nor UO_200 (O_200,N_9914,N_9934);
nor UO_201 (O_201,N_9943,N_9944);
and UO_202 (O_202,N_9985,N_9991);
or UO_203 (O_203,N_9913,N_9958);
or UO_204 (O_204,N_9990,N_9989);
or UO_205 (O_205,N_9967,N_9951);
nor UO_206 (O_206,N_9912,N_9985);
and UO_207 (O_207,N_9947,N_9948);
or UO_208 (O_208,N_9909,N_9916);
or UO_209 (O_209,N_9984,N_9915);
nand UO_210 (O_210,N_9993,N_9950);
nor UO_211 (O_211,N_9933,N_9990);
or UO_212 (O_212,N_9966,N_9976);
nand UO_213 (O_213,N_9957,N_9995);
nor UO_214 (O_214,N_9938,N_9916);
and UO_215 (O_215,N_9942,N_9984);
nor UO_216 (O_216,N_9991,N_9976);
nand UO_217 (O_217,N_9953,N_9944);
nor UO_218 (O_218,N_9917,N_9944);
nand UO_219 (O_219,N_9923,N_9925);
nor UO_220 (O_220,N_9979,N_9923);
or UO_221 (O_221,N_9963,N_9939);
nand UO_222 (O_222,N_9918,N_9997);
nand UO_223 (O_223,N_9916,N_9991);
nor UO_224 (O_224,N_9961,N_9906);
xor UO_225 (O_225,N_9900,N_9955);
and UO_226 (O_226,N_9901,N_9952);
nor UO_227 (O_227,N_9969,N_9921);
and UO_228 (O_228,N_9967,N_9948);
or UO_229 (O_229,N_9921,N_9992);
nand UO_230 (O_230,N_9916,N_9963);
and UO_231 (O_231,N_9965,N_9931);
nor UO_232 (O_232,N_9923,N_9994);
nand UO_233 (O_233,N_9994,N_9905);
nor UO_234 (O_234,N_9950,N_9915);
nand UO_235 (O_235,N_9944,N_9984);
nand UO_236 (O_236,N_9939,N_9990);
nand UO_237 (O_237,N_9909,N_9971);
nand UO_238 (O_238,N_9943,N_9919);
or UO_239 (O_239,N_9953,N_9966);
and UO_240 (O_240,N_9984,N_9989);
nand UO_241 (O_241,N_9913,N_9939);
and UO_242 (O_242,N_9952,N_9934);
and UO_243 (O_243,N_9913,N_9938);
or UO_244 (O_244,N_9966,N_9952);
nand UO_245 (O_245,N_9948,N_9990);
or UO_246 (O_246,N_9952,N_9911);
and UO_247 (O_247,N_9915,N_9941);
and UO_248 (O_248,N_9915,N_9974);
and UO_249 (O_249,N_9904,N_9976);
or UO_250 (O_250,N_9977,N_9955);
nor UO_251 (O_251,N_9992,N_9934);
nand UO_252 (O_252,N_9901,N_9956);
or UO_253 (O_253,N_9905,N_9973);
nor UO_254 (O_254,N_9922,N_9955);
nand UO_255 (O_255,N_9929,N_9976);
nand UO_256 (O_256,N_9976,N_9923);
and UO_257 (O_257,N_9938,N_9930);
and UO_258 (O_258,N_9905,N_9902);
nand UO_259 (O_259,N_9946,N_9924);
or UO_260 (O_260,N_9986,N_9956);
and UO_261 (O_261,N_9999,N_9996);
or UO_262 (O_262,N_9972,N_9998);
and UO_263 (O_263,N_9941,N_9909);
and UO_264 (O_264,N_9976,N_9984);
nand UO_265 (O_265,N_9993,N_9947);
and UO_266 (O_266,N_9917,N_9983);
or UO_267 (O_267,N_9994,N_9952);
nor UO_268 (O_268,N_9945,N_9933);
nor UO_269 (O_269,N_9996,N_9908);
or UO_270 (O_270,N_9943,N_9986);
or UO_271 (O_271,N_9933,N_9957);
or UO_272 (O_272,N_9927,N_9981);
or UO_273 (O_273,N_9931,N_9915);
and UO_274 (O_274,N_9913,N_9980);
or UO_275 (O_275,N_9986,N_9915);
or UO_276 (O_276,N_9945,N_9922);
or UO_277 (O_277,N_9911,N_9957);
nor UO_278 (O_278,N_9942,N_9967);
and UO_279 (O_279,N_9919,N_9930);
or UO_280 (O_280,N_9921,N_9964);
or UO_281 (O_281,N_9902,N_9964);
and UO_282 (O_282,N_9956,N_9995);
nor UO_283 (O_283,N_9930,N_9927);
and UO_284 (O_284,N_9933,N_9960);
nor UO_285 (O_285,N_9920,N_9917);
or UO_286 (O_286,N_9960,N_9984);
and UO_287 (O_287,N_9954,N_9929);
nor UO_288 (O_288,N_9960,N_9901);
or UO_289 (O_289,N_9919,N_9970);
and UO_290 (O_290,N_9964,N_9972);
and UO_291 (O_291,N_9919,N_9980);
or UO_292 (O_292,N_9940,N_9987);
xor UO_293 (O_293,N_9911,N_9994);
and UO_294 (O_294,N_9969,N_9928);
nor UO_295 (O_295,N_9975,N_9917);
or UO_296 (O_296,N_9921,N_9922);
nand UO_297 (O_297,N_9957,N_9919);
nand UO_298 (O_298,N_9932,N_9955);
nor UO_299 (O_299,N_9910,N_9990);
and UO_300 (O_300,N_9930,N_9903);
and UO_301 (O_301,N_9949,N_9914);
or UO_302 (O_302,N_9951,N_9929);
nor UO_303 (O_303,N_9975,N_9950);
nand UO_304 (O_304,N_9935,N_9969);
nor UO_305 (O_305,N_9953,N_9965);
or UO_306 (O_306,N_9912,N_9976);
nor UO_307 (O_307,N_9936,N_9919);
nand UO_308 (O_308,N_9937,N_9966);
or UO_309 (O_309,N_9915,N_9934);
nand UO_310 (O_310,N_9912,N_9908);
and UO_311 (O_311,N_9921,N_9977);
or UO_312 (O_312,N_9992,N_9989);
nand UO_313 (O_313,N_9915,N_9932);
and UO_314 (O_314,N_9947,N_9973);
and UO_315 (O_315,N_9971,N_9945);
nand UO_316 (O_316,N_9916,N_9933);
and UO_317 (O_317,N_9962,N_9971);
or UO_318 (O_318,N_9928,N_9997);
or UO_319 (O_319,N_9980,N_9927);
or UO_320 (O_320,N_9968,N_9903);
and UO_321 (O_321,N_9919,N_9952);
nand UO_322 (O_322,N_9989,N_9997);
nand UO_323 (O_323,N_9917,N_9942);
nor UO_324 (O_324,N_9986,N_9946);
or UO_325 (O_325,N_9919,N_9926);
and UO_326 (O_326,N_9984,N_9901);
nand UO_327 (O_327,N_9958,N_9977);
nand UO_328 (O_328,N_9998,N_9926);
or UO_329 (O_329,N_9966,N_9987);
nor UO_330 (O_330,N_9989,N_9935);
and UO_331 (O_331,N_9940,N_9947);
nor UO_332 (O_332,N_9971,N_9957);
nor UO_333 (O_333,N_9916,N_9926);
or UO_334 (O_334,N_9912,N_9990);
or UO_335 (O_335,N_9999,N_9977);
nor UO_336 (O_336,N_9907,N_9942);
and UO_337 (O_337,N_9959,N_9911);
nor UO_338 (O_338,N_9955,N_9905);
nor UO_339 (O_339,N_9935,N_9947);
or UO_340 (O_340,N_9920,N_9944);
or UO_341 (O_341,N_9904,N_9986);
and UO_342 (O_342,N_9941,N_9985);
nor UO_343 (O_343,N_9965,N_9909);
and UO_344 (O_344,N_9902,N_9987);
nand UO_345 (O_345,N_9915,N_9940);
and UO_346 (O_346,N_9993,N_9978);
nand UO_347 (O_347,N_9926,N_9997);
nor UO_348 (O_348,N_9969,N_9997);
or UO_349 (O_349,N_9959,N_9981);
or UO_350 (O_350,N_9934,N_9909);
nor UO_351 (O_351,N_9998,N_9929);
nor UO_352 (O_352,N_9901,N_9940);
nor UO_353 (O_353,N_9910,N_9946);
nor UO_354 (O_354,N_9941,N_9952);
nand UO_355 (O_355,N_9962,N_9997);
or UO_356 (O_356,N_9997,N_9967);
and UO_357 (O_357,N_9961,N_9907);
and UO_358 (O_358,N_9986,N_9962);
and UO_359 (O_359,N_9999,N_9989);
or UO_360 (O_360,N_9918,N_9907);
nand UO_361 (O_361,N_9937,N_9933);
nor UO_362 (O_362,N_9966,N_9921);
or UO_363 (O_363,N_9984,N_9918);
or UO_364 (O_364,N_9995,N_9946);
nor UO_365 (O_365,N_9967,N_9911);
nand UO_366 (O_366,N_9962,N_9901);
nand UO_367 (O_367,N_9926,N_9985);
nor UO_368 (O_368,N_9959,N_9930);
nor UO_369 (O_369,N_9980,N_9948);
and UO_370 (O_370,N_9955,N_9970);
nand UO_371 (O_371,N_9954,N_9961);
and UO_372 (O_372,N_9923,N_9960);
nand UO_373 (O_373,N_9968,N_9989);
nor UO_374 (O_374,N_9949,N_9916);
nor UO_375 (O_375,N_9998,N_9986);
and UO_376 (O_376,N_9985,N_9983);
nor UO_377 (O_377,N_9978,N_9941);
nand UO_378 (O_378,N_9939,N_9979);
nor UO_379 (O_379,N_9989,N_9947);
or UO_380 (O_380,N_9927,N_9933);
or UO_381 (O_381,N_9919,N_9924);
nand UO_382 (O_382,N_9965,N_9980);
and UO_383 (O_383,N_9967,N_9962);
nor UO_384 (O_384,N_9922,N_9956);
or UO_385 (O_385,N_9946,N_9962);
nor UO_386 (O_386,N_9958,N_9978);
and UO_387 (O_387,N_9945,N_9909);
and UO_388 (O_388,N_9958,N_9976);
nand UO_389 (O_389,N_9910,N_9925);
nand UO_390 (O_390,N_9966,N_9961);
nor UO_391 (O_391,N_9955,N_9939);
nor UO_392 (O_392,N_9957,N_9928);
or UO_393 (O_393,N_9966,N_9992);
nor UO_394 (O_394,N_9959,N_9926);
or UO_395 (O_395,N_9958,N_9926);
nand UO_396 (O_396,N_9974,N_9977);
or UO_397 (O_397,N_9963,N_9981);
or UO_398 (O_398,N_9935,N_9945);
or UO_399 (O_399,N_9969,N_9987);
and UO_400 (O_400,N_9948,N_9946);
nor UO_401 (O_401,N_9948,N_9975);
and UO_402 (O_402,N_9992,N_9988);
or UO_403 (O_403,N_9980,N_9993);
nand UO_404 (O_404,N_9900,N_9922);
nand UO_405 (O_405,N_9913,N_9997);
nand UO_406 (O_406,N_9909,N_9960);
or UO_407 (O_407,N_9963,N_9955);
or UO_408 (O_408,N_9970,N_9905);
nor UO_409 (O_409,N_9935,N_9951);
or UO_410 (O_410,N_9981,N_9929);
nand UO_411 (O_411,N_9978,N_9930);
nand UO_412 (O_412,N_9994,N_9928);
and UO_413 (O_413,N_9932,N_9901);
nand UO_414 (O_414,N_9932,N_9933);
and UO_415 (O_415,N_9984,N_9981);
or UO_416 (O_416,N_9926,N_9930);
nor UO_417 (O_417,N_9995,N_9922);
or UO_418 (O_418,N_9951,N_9993);
or UO_419 (O_419,N_9920,N_9929);
and UO_420 (O_420,N_9969,N_9909);
xnor UO_421 (O_421,N_9971,N_9970);
or UO_422 (O_422,N_9968,N_9939);
and UO_423 (O_423,N_9985,N_9998);
nor UO_424 (O_424,N_9997,N_9919);
nand UO_425 (O_425,N_9978,N_9949);
or UO_426 (O_426,N_9919,N_9953);
or UO_427 (O_427,N_9953,N_9979);
nand UO_428 (O_428,N_9954,N_9997);
nand UO_429 (O_429,N_9954,N_9943);
nand UO_430 (O_430,N_9921,N_9997);
and UO_431 (O_431,N_9950,N_9948);
or UO_432 (O_432,N_9998,N_9966);
nor UO_433 (O_433,N_9908,N_9929);
nand UO_434 (O_434,N_9982,N_9972);
and UO_435 (O_435,N_9916,N_9953);
or UO_436 (O_436,N_9979,N_9943);
and UO_437 (O_437,N_9989,N_9980);
or UO_438 (O_438,N_9933,N_9964);
nand UO_439 (O_439,N_9930,N_9932);
and UO_440 (O_440,N_9989,N_9936);
or UO_441 (O_441,N_9914,N_9997);
nand UO_442 (O_442,N_9975,N_9958);
nand UO_443 (O_443,N_9970,N_9931);
and UO_444 (O_444,N_9992,N_9905);
and UO_445 (O_445,N_9979,N_9987);
xnor UO_446 (O_446,N_9910,N_9924);
or UO_447 (O_447,N_9993,N_9953);
nor UO_448 (O_448,N_9939,N_9943);
and UO_449 (O_449,N_9947,N_9908);
nor UO_450 (O_450,N_9933,N_9924);
or UO_451 (O_451,N_9955,N_9949);
nor UO_452 (O_452,N_9937,N_9963);
and UO_453 (O_453,N_9956,N_9998);
and UO_454 (O_454,N_9924,N_9909);
nor UO_455 (O_455,N_9961,N_9902);
or UO_456 (O_456,N_9989,N_9976);
nor UO_457 (O_457,N_9946,N_9968);
nor UO_458 (O_458,N_9953,N_9922);
and UO_459 (O_459,N_9951,N_9942);
nor UO_460 (O_460,N_9928,N_9927);
and UO_461 (O_461,N_9992,N_9912);
and UO_462 (O_462,N_9989,N_9960);
and UO_463 (O_463,N_9945,N_9964);
nand UO_464 (O_464,N_9929,N_9931);
or UO_465 (O_465,N_9981,N_9998);
or UO_466 (O_466,N_9913,N_9991);
or UO_467 (O_467,N_9919,N_9981);
nand UO_468 (O_468,N_9907,N_9906);
nand UO_469 (O_469,N_9933,N_9952);
nor UO_470 (O_470,N_9918,N_9971);
nor UO_471 (O_471,N_9941,N_9963);
nand UO_472 (O_472,N_9987,N_9960);
or UO_473 (O_473,N_9912,N_9910);
or UO_474 (O_474,N_9970,N_9943);
nor UO_475 (O_475,N_9977,N_9956);
nand UO_476 (O_476,N_9958,N_9911);
nand UO_477 (O_477,N_9989,N_9991);
and UO_478 (O_478,N_9977,N_9971);
nand UO_479 (O_479,N_9917,N_9947);
and UO_480 (O_480,N_9906,N_9925);
nand UO_481 (O_481,N_9977,N_9997);
or UO_482 (O_482,N_9955,N_9915);
and UO_483 (O_483,N_9965,N_9952);
nor UO_484 (O_484,N_9908,N_9978);
or UO_485 (O_485,N_9959,N_9949);
and UO_486 (O_486,N_9953,N_9957);
nor UO_487 (O_487,N_9999,N_9949);
nor UO_488 (O_488,N_9992,N_9938);
nor UO_489 (O_489,N_9926,N_9983);
nand UO_490 (O_490,N_9994,N_9968);
and UO_491 (O_491,N_9920,N_9959);
and UO_492 (O_492,N_9922,N_9938);
or UO_493 (O_493,N_9949,N_9986);
or UO_494 (O_494,N_9959,N_9985);
and UO_495 (O_495,N_9932,N_9939);
nor UO_496 (O_496,N_9968,N_9988);
nor UO_497 (O_497,N_9942,N_9998);
and UO_498 (O_498,N_9972,N_9939);
and UO_499 (O_499,N_9975,N_9973);
nand UO_500 (O_500,N_9916,N_9920);
and UO_501 (O_501,N_9991,N_9912);
nand UO_502 (O_502,N_9901,N_9982);
nor UO_503 (O_503,N_9955,N_9938);
or UO_504 (O_504,N_9969,N_9959);
or UO_505 (O_505,N_9900,N_9962);
nand UO_506 (O_506,N_9964,N_9919);
or UO_507 (O_507,N_9971,N_9946);
or UO_508 (O_508,N_9983,N_9984);
nand UO_509 (O_509,N_9921,N_9938);
nand UO_510 (O_510,N_9934,N_9921);
and UO_511 (O_511,N_9983,N_9908);
or UO_512 (O_512,N_9940,N_9977);
nor UO_513 (O_513,N_9980,N_9955);
or UO_514 (O_514,N_9903,N_9966);
or UO_515 (O_515,N_9900,N_9933);
and UO_516 (O_516,N_9911,N_9969);
nor UO_517 (O_517,N_9953,N_9961);
and UO_518 (O_518,N_9919,N_9965);
nand UO_519 (O_519,N_9918,N_9911);
nand UO_520 (O_520,N_9959,N_9988);
nand UO_521 (O_521,N_9914,N_9978);
and UO_522 (O_522,N_9900,N_9982);
nor UO_523 (O_523,N_9974,N_9996);
nor UO_524 (O_524,N_9907,N_9914);
nand UO_525 (O_525,N_9902,N_9922);
nand UO_526 (O_526,N_9904,N_9991);
or UO_527 (O_527,N_9943,N_9972);
nor UO_528 (O_528,N_9943,N_9951);
nor UO_529 (O_529,N_9905,N_9983);
nand UO_530 (O_530,N_9917,N_9904);
and UO_531 (O_531,N_9995,N_9965);
and UO_532 (O_532,N_9932,N_9951);
or UO_533 (O_533,N_9900,N_9984);
or UO_534 (O_534,N_9907,N_9969);
nor UO_535 (O_535,N_9946,N_9930);
and UO_536 (O_536,N_9987,N_9971);
and UO_537 (O_537,N_9989,N_9902);
and UO_538 (O_538,N_9968,N_9954);
and UO_539 (O_539,N_9929,N_9994);
or UO_540 (O_540,N_9901,N_9917);
or UO_541 (O_541,N_9973,N_9922);
nor UO_542 (O_542,N_9965,N_9938);
or UO_543 (O_543,N_9977,N_9928);
or UO_544 (O_544,N_9900,N_9977);
or UO_545 (O_545,N_9931,N_9986);
and UO_546 (O_546,N_9979,N_9906);
and UO_547 (O_547,N_9927,N_9937);
nand UO_548 (O_548,N_9989,N_9917);
nor UO_549 (O_549,N_9920,N_9910);
nand UO_550 (O_550,N_9959,N_9941);
or UO_551 (O_551,N_9913,N_9949);
nand UO_552 (O_552,N_9939,N_9914);
nand UO_553 (O_553,N_9916,N_9965);
or UO_554 (O_554,N_9976,N_9945);
or UO_555 (O_555,N_9952,N_9943);
nor UO_556 (O_556,N_9947,N_9988);
or UO_557 (O_557,N_9915,N_9954);
nand UO_558 (O_558,N_9950,N_9936);
or UO_559 (O_559,N_9998,N_9930);
and UO_560 (O_560,N_9955,N_9997);
nand UO_561 (O_561,N_9973,N_9953);
nor UO_562 (O_562,N_9909,N_9959);
and UO_563 (O_563,N_9922,N_9978);
nor UO_564 (O_564,N_9907,N_9988);
nor UO_565 (O_565,N_9953,N_9925);
and UO_566 (O_566,N_9995,N_9967);
nor UO_567 (O_567,N_9909,N_9937);
and UO_568 (O_568,N_9958,N_9998);
or UO_569 (O_569,N_9981,N_9912);
nand UO_570 (O_570,N_9929,N_9937);
or UO_571 (O_571,N_9928,N_9908);
nor UO_572 (O_572,N_9956,N_9926);
and UO_573 (O_573,N_9956,N_9954);
nand UO_574 (O_574,N_9907,N_9903);
nand UO_575 (O_575,N_9931,N_9972);
and UO_576 (O_576,N_9909,N_9963);
or UO_577 (O_577,N_9930,N_9904);
nand UO_578 (O_578,N_9962,N_9917);
nand UO_579 (O_579,N_9950,N_9902);
or UO_580 (O_580,N_9956,N_9964);
nand UO_581 (O_581,N_9926,N_9903);
nand UO_582 (O_582,N_9926,N_9913);
and UO_583 (O_583,N_9924,N_9974);
nand UO_584 (O_584,N_9999,N_9997);
and UO_585 (O_585,N_9985,N_9956);
or UO_586 (O_586,N_9958,N_9901);
nand UO_587 (O_587,N_9918,N_9946);
and UO_588 (O_588,N_9974,N_9969);
or UO_589 (O_589,N_9972,N_9929);
nor UO_590 (O_590,N_9913,N_9918);
and UO_591 (O_591,N_9972,N_9992);
nand UO_592 (O_592,N_9985,N_9986);
and UO_593 (O_593,N_9947,N_9925);
and UO_594 (O_594,N_9916,N_9959);
nor UO_595 (O_595,N_9957,N_9962);
and UO_596 (O_596,N_9938,N_9988);
and UO_597 (O_597,N_9910,N_9950);
and UO_598 (O_598,N_9950,N_9967);
nor UO_599 (O_599,N_9943,N_9913);
nor UO_600 (O_600,N_9998,N_9955);
and UO_601 (O_601,N_9999,N_9957);
or UO_602 (O_602,N_9964,N_9952);
or UO_603 (O_603,N_9920,N_9933);
nand UO_604 (O_604,N_9969,N_9954);
nand UO_605 (O_605,N_9967,N_9916);
or UO_606 (O_606,N_9951,N_9933);
nand UO_607 (O_607,N_9912,N_9963);
and UO_608 (O_608,N_9988,N_9967);
and UO_609 (O_609,N_9907,N_9992);
nand UO_610 (O_610,N_9958,N_9980);
nand UO_611 (O_611,N_9966,N_9978);
and UO_612 (O_612,N_9925,N_9997);
nor UO_613 (O_613,N_9981,N_9928);
nor UO_614 (O_614,N_9971,N_9993);
and UO_615 (O_615,N_9903,N_9960);
nor UO_616 (O_616,N_9949,N_9925);
nand UO_617 (O_617,N_9921,N_9986);
or UO_618 (O_618,N_9970,N_9977);
nor UO_619 (O_619,N_9903,N_9913);
nor UO_620 (O_620,N_9904,N_9990);
nor UO_621 (O_621,N_9923,N_9922);
or UO_622 (O_622,N_9927,N_9971);
and UO_623 (O_623,N_9931,N_9990);
and UO_624 (O_624,N_9972,N_9922);
or UO_625 (O_625,N_9918,N_9906);
or UO_626 (O_626,N_9964,N_9987);
and UO_627 (O_627,N_9995,N_9929);
or UO_628 (O_628,N_9973,N_9987);
nor UO_629 (O_629,N_9941,N_9918);
and UO_630 (O_630,N_9901,N_9978);
nand UO_631 (O_631,N_9991,N_9957);
nor UO_632 (O_632,N_9903,N_9934);
and UO_633 (O_633,N_9948,N_9902);
xor UO_634 (O_634,N_9990,N_9973);
nand UO_635 (O_635,N_9907,N_9981);
and UO_636 (O_636,N_9955,N_9948);
nand UO_637 (O_637,N_9961,N_9975);
or UO_638 (O_638,N_9976,N_9987);
nor UO_639 (O_639,N_9924,N_9935);
nand UO_640 (O_640,N_9988,N_9990);
and UO_641 (O_641,N_9925,N_9933);
and UO_642 (O_642,N_9911,N_9983);
nand UO_643 (O_643,N_9939,N_9958);
or UO_644 (O_644,N_9913,N_9957);
nor UO_645 (O_645,N_9945,N_9907);
or UO_646 (O_646,N_9976,N_9943);
or UO_647 (O_647,N_9990,N_9907);
and UO_648 (O_648,N_9976,N_9930);
nor UO_649 (O_649,N_9922,N_9982);
nor UO_650 (O_650,N_9938,N_9956);
or UO_651 (O_651,N_9998,N_9952);
or UO_652 (O_652,N_9977,N_9947);
or UO_653 (O_653,N_9984,N_9931);
nand UO_654 (O_654,N_9907,N_9953);
or UO_655 (O_655,N_9937,N_9908);
nor UO_656 (O_656,N_9935,N_9910);
and UO_657 (O_657,N_9975,N_9908);
and UO_658 (O_658,N_9969,N_9976);
nand UO_659 (O_659,N_9906,N_9901);
or UO_660 (O_660,N_9944,N_9989);
nor UO_661 (O_661,N_9979,N_9991);
nor UO_662 (O_662,N_9913,N_9919);
nor UO_663 (O_663,N_9955,N_9993);
and UO_664 (O_664,N_9999,N_9954);
or UO_665 (O_665,N_9920,N_9939);
nor UO_666 (O_666,N_9944,N_9912);
nand UO_667 (O_667,N_9908,N_9923);
nand UO_668 (O_668,N_9956,N_9963);
nand UO_669 (O_669,N_9979,N_9911);
nand UO_670 (O_670,N_9913,N_9963);
and UO_671 (O_671,N_9900,N_9951);
and UO_672 (O_672,N_9943,N_9909);
nor UO_673 (O_673,N_9911,N_9966);
or UO_674 (O_674,N_9988,N_9996);
and UO_675 (O_675,N_9931,N_9914);
or UO_676 (O_676,N_9941,N_9914);
or UO_677 (O_677,N_9960,N_9919);
and UO_678 (O_678,N_9902,N_9982);
nor UO_679 (O_679,N_9934,N_9991);
and UO_680 (O_680,N_9915,N_9980);
nand UO_681 (O_681,N_9981,N_9999);
and UO_682 (O_682,N_9996,N_9948);
and UO_683 (O_683,N_9959,N_9932);
nand UO_684 (O_684,N_9978,N_9905);
nand UO_685 (O_685,N_9973,N_9911);
nor UO_686 (O_686,N_9956,N_9934);
nand UO_687 (O_687,N_9983,N_9946);
nand UO_688 (O_688,N_9943,N_9963);
and UO_689 (O_689,N_9983,N_9945);
and UO_690 (O_690,N_9955,N_9942);
nor UO_691 (O_691,N_9974,N_9936);
nor UO_692 (O_692,N_9942,N_9980);
or UO_693 (O_693,N_9980,N_9959);
nor UO_694 (O_694,N_9908,N_9973);
or UO_695 (O_695,N_9985,N_9937);
and UO_696 (O_696,N_9950,N_9989);
and UO_697 (O_697,N_9952,N_9942);
and UO_698 (O_698,N_9957,N_9932);
nor UO_699 (O_699,N_9976,N_9931);
or UO_700 (O_700,N_9983,N_9944);
nor UO_701 (O_701,N_9957,N_9908);
xnor UO_702 (O_702,N_9976,N_9900);
or UO_703 (O_703,N_9981,N_9954);
and UO_704 (O_704,N_9951,N_9997);
or UO_705 (O_705,N_9903,N_9991);
nand UO_706 (O_706,N_9902,N_9956);
nand UO_707 (O_707,N_9940,N_9941);
nand UO_708 (O_708,N_9974,N_9957);
or UO_709 (O_709,N_9991,N_9970);
or UO_710 (O_710,N_9982,N_9965);
and UO_711 (O_711,N_9949,N_9929);
or UO_712 (O_712,N_9988,N_9940);
or UO_713 (O_713,N_9920,N_9968);
nand UO_714 (O_714,N_9910,N_9995);
nor UO_715 (O_715,N_9950,N_9982);
or UO_716 (O_716,N_9912,N_9902);
nor UO_717 (O_717,N_9910,N_9975);
nand UO_718 (O_718,N_9925,N_9975);
or UO_719 (O_719,N_9953,N_9983);
or UO_720 (O_720,N_9908,N_9915);
or UO_721 (O_721,N_9984,N_9913);
or UO_722 (O_722,N_9945,N_9902);
nand UO_723 (O_723,N_9979,N_9959);
nor UO_724 (O_724,N_9918,N_9934);
nand UO_725 (O_725,N_9908,N_9906);
nand UO_726 (O_726,N_9911,N_9991);
nand UO_727 (O_727,N_9963,N_9932);
or UO_728 (O_728,N_9947,N_9913);
nand UO_729 (O_729,N_9955,N_9926);
nand UO_730 (O_730,N_9913,N_9945);
and UO_731 (O_731,N_9964,N_9943);
nor UO_732 (O_732,N_9922,N_9917);
nand UO_733 (O_733,N_9980,N_9982);
or UO_734 (O_734,N_9905,N_9964);
nand UO_735 (O_735,N_9944,N_9933);
and UO_736 (O_736,N_9991,N_9922);
nor UO_737 (O_737,N_9951,N_9903);
or UO_738 (O_738,N_9966,N_9943);
or UO_739 (O_739,N_9937,N_9919);
or UO_740 (O_740,N_9990,N_9922);
nor UO_741 (O_741,N_9923,N_9930);
nand UO_742 (O_742,N_9932,N_9949);
nand UO_743 (O_743,N_9948,N_9994);
nor UO_744 (O_744,N_9920,N_9973);
nand UO_745 (O_745,N_9932,N_9934);
or UO_746 (O_746,N_9932,N_9962);
nand UO_747 (O_747,N_9959,N_9907);
or UO_748 (O_748,N_9927,N_9929);
and UO_749 (O_749,N_9928,N_9942);
nand UO_750 (O_750,N_9982,N_9987);
nor UO_751 (O_751,N_9959,N_9942);
or UO_752 (O_752,N_9915,N_9976);
or UO_753 (O_753,N_9920,N_9948);
xor UO_754 (O_754,N_9962,N_9955);
nor UO_755 (O_755,N_9911,N_9938);
and UO_756 (O_756,N_9988,N_9957);
or UO_757 (O_757,N_9994,N_9983);
nor UO_758 (O_758,N_9994,N_9917);
nor UO_759 (O_759,N_9973,N_9963);
nor UO_760 (O_760,N_9972,N_9926);
and UO_761 (O_761,N_9944,N_9942);
nand UO_762 (O_762,N_9973,N_9979);
nand UO_763 (O_763,N_9938,N_9909);
and UO_764 (O_764,N_9970,N_9995);
or UO_765 (O_765,N_9998,N_9939);
and UO_766 (O_766,N_9967,N_9941);
and UO_767 (O_767,N_9906,N_9989);
and UO_768 (O_768,N_9932,N_9929);
or UO_769 (O_769,N_9989,N_9920);
nand UO_770 (O_770,N_9994,N_9937);
or UO_771 (O_771,N_9978,N_9990);
or UO_772 (O_772,N_9970,N_9917);
or UO_773 (O_773,N_9965,N_9989);
and UO_774 (O_774,N_9959,N_9908);
and UO_775 (O_775,N_9996,N_9902);
or UO_776 (O_776,N_9988,N_9961);
and UO_777 (O_777,N_9932,N_9966);
and UO_778 (O_778,N_9901,N_9999);
and UO_779 (O_779,N_9923,N_9943);
or UO_780 (O_780,N_9940,N_9948);
nand UO_781 (O_781,N_9988,N_9976);
or UO_782 (O_782,N_9967,N_9989);
or UO_783 (O_783,N_9972,N_9936);
nor UO_784 (O_784,N_9931,N_9967);
nor UO_785 (O_785,N_9913,N_9976);
xnor UO_786 (O_786,N_9916,N_9979);
nand UO_787 (O_787,N_9992,N_9952);
or UO_788 (O_788,N_9943,N_9947);
nor UO_789 (O_789,N_9994,N_9947);
or UO_790 (O_790,N_9943,N_9968);
xor UO_791 (O_791,N_9905,N_9920);
nand UO_792 (O_792,N_9934,N_9936);
nor UO_793 (O_793,N_9957,N_9929);
nor UO_794 (O_794,N_9950,N_9994);
nor UO_795 (O_795,N_9958,N_9923);
nor UO_796 (O_796,N_9942,N_9934);
nand UO_797 (O_797,N_9901,N_9983);
and UO_798 (O_798,N_9936,N_9979);
nor UO_799 (O_799,N_9904,N_9956);
nand UO_800 (O_800,N_9926,N_9954);
xnor UO_801 (O_801,N_9967,N_9924);
nor UO_802 (O_802,N_9903,N_9936);
or UO_803 (O_803,N_9901,N_9943);
and UO_804 (O_804,N_9934,N_9994);
and UO_805 (O_805,N_9955,N_9935);
nand UO_806 (O_806,N_9935,N_9902);
xor UO_807 (O_807,N_9954,N_9984);
nor UO_808 (O_808,N_9914,N_9916);
nand UO_809 (O_809,N_9990,N_9964);
nor UO_810 (O_810,N_9944,N_9958);
nand UO_811 (O_811,N_9990,N_9934);
nor UO_812 (O_812,N_9999,N_9915);
nand UO_813 (O_813,N_9957,N_9968);
and UO_814 (O_814,N_9982,N_9994);
nand UO_815 (O_815,N_9951,N_9987);
or UO_816 (O_816,N_9986,N_9950);
nor UO_817 (O_817,N_9902,N_9925);
or UO_818 (O_818,N_9918,N_9936);
nor UO_819 (O_819,N_9989,N_9901);
nand UO_820 (O_820,N_9955,N_9979);
nand UO_821 (O_821,N_9900,N_9949);
nor UO_822 (O_822,N_9936,N_9991);
nor UO_823 (O_823,N_9948,N_9965);
and UO_824 (O_824,N_9945,N_9932);
or UO_825 (O_825,N_9927,N_9905);
nor UO_826 (O_826,N_9953,N_9984);
nand UO_827 (O_827,N_9947,N_9966);
or UO_828 (O_828,N_9995,N_9977);
and UO_829 (O_829,N_9909,N_9935);
nor UO_830 (O_830,N_9968,N_9934);
and UO_831 (O_831,N_9935,N_9912);
and UO_832 (O_832,N_9910,N_9977);
or UO_833 (O_833,N_9924,N_9922);
nor UO_834 (O_834,N_9987,N_9934);
and UO_835 (O_835,N_9929,N_9919);
nand UO_836 (O_836,N_9945,N_9992);
and UO_837 (O_837,N_9905,N_9912);
nand UO_838 (O_838,N_9903,N_9940);
or UO_839 (O_839,N_9931,N_9994);
and UO_840 (O_840,N_9927,N_9907);
or UO_841 (O_841,N_9966,N_9968);
and UO_842 (O_842,N_9957,N_9904);
nor UO_843 (O_843,N_9954,N_9949);
and UO_844 (O_844,N_9979,N_9985);
or UO_845 (O_845,N_9970,N_9972);
nor UO_846 (O_846,N_9968,N_9960);
and UO_847 (O_847,N_9952,N_9973);
nand UO_848 (O_848,N_9988,N_9965);
nor UO_849 (O_849,N_9963,N_9946);
or UO_850 (O_850,N_9924,N_9983);
or UO_851 (O_851,N_9927,N_9976);
nand UO_852 (O_852,N_9947,N_9915);
nand UO_853 (O_853,N_9902,N_9910);
or UO_854 (O_854,N_9999,N_9974);
nor UO_855 (O_855,N_9919,N_9972);
nand UO_856 (O_856,N_9995,N_9951);
and UO_857 (O_857,N_9964,N_9982);
and UO_858 (O_858,N_9905,N_9995);
nor UO_859 (O_859,N_9958,N_9973);
nor UO_860 (O_860,N_9930,N_9937);
nor UO_861 (O_861,N_9993,N_9917);
nor UO_862 (O_862,N_9950,N_9962);
nand UO_863 (O_863,N_9969,N_9956);
and UO_864 (O_864,N_9948,N_9943);
or UO_865 (O_865,N_9936,N_9900);
nand UO_866 (O_866,N_9903,N_9901);
or UO_867 (O_867,N_9978,N_9953);
or UO_868 (O_868,N_9914,N_9983);
nand UO_869 (O_869,N_9940,N_9990);
nand UO_870 (O_870,N_9951,N_9969);
nor UO_871 (O_871,N_9973,N_9944);
or UO_872 (O_872,N_9920,N_9919);
nand UO_873 (O_873,N_9922,N_9926);
or UO_874 (O_874,N_9913,N_9936);
and UO_875 (O_875,N_9973,N_9970);
nor UO_876 (O_876,N_9962,N_9968);
or UO_877 (O_877,N_9920,N_9936);
nor UO_878 (O_878,N_9907,N_9955);
nand UO_879 (O_879,N_9951,N_9913);
nand UO_880 (O_880,N_9965,N_9968);
nand UO_881 (O_881,N_9945,N_9947);
or UO_882 (O_882,N_9956,N_9953);
xor UO_883 (O_883,N_9923,N_9963);
or UO_884 (O_884,N_9951,N_9985);
xor UO_885 (O_885,N_9959,N_9956);
or UO_886 (O_886,N_9909,N_9925);
or UO_887 (O_887,N_9994,N_9900);
or UO_888 (O_888,N_9920,N_9928);
and UO_889 (O_889,N_9953,N_9950);
nand UO_890 (O_890,N_9947,N_9934);
and UO_891 (O_891,N_9982,N_9959);
and UO_892 (O_892,N_9921,N_9930);
nor UO_893 (O_893,N_9914,N_9900);
and UO_894 (O_894,N_9965,N_9910);
or UO_895 (O_895,N_9942,N_9969);
or UO_896 (O_896,N_9939,N_9916);
or UO_897 (O_897,N_9965,N_9976);
nor UO_898 (O_898,N_9983,N_9960);
or UO_899 (O_899,N_9966,N_9977);
and UO_900 (O_900,N_9925,N_9968);
or UO_901 (O_901,N_9958,N_9963);
nand UO_902 (O_902,N_9910,N_9936);
or UO_903 (O_903,N_9983,N_9981);
nor UO_904 (O_904,N_9960,N_9915);
and UO_905 (O_905,N_9961,N_9996);
and UO_906 (O_906,N_9935,N_9908);
and UO_907 (O_907,N_9971,N_9986);
and UO_908 (O_908,N_9960,N_9950);
nand UO_909 (O_909,N_9918,N_9989);
or UO_910 (O_910,N_9956,N_9929);
nor UO_911 (O_911,N_9970,N_9959);
or UO_912 (O_912,N_9981,N_9924);
nor UO_913 (O_913,N_9988,N_9987);
nand UO_914 (O_914,N_9957,N_9952);
nor UO_915 (O_915,N_9933,N_9996);
xor UO_916 (O_916,N_9909,N_9917);
and UO_917 (O_917,N_9942,N_9941);
and UO_918 (O_918,N_9981,N_9980);
and UO_919 (O_919,N_9935,N_9905);
or UO_920 (O_920,N_9966,N_9954);
nand UO_921 (O_921,N_9915,N_9913);
or UO_922 (O_922,N_9943,N_9962);
nand UO_923 (O_923,N_9931,N_9950);
and UO_924 (O_924,N_9954,N_9902);
nand UO_925 (O_925,N_9979,N_9976);
nor UO_926 (O_926,N_9990,N_9944);
or UO_927 (O_927,N_9960,N_9935);
or UO_928 (O_928,N_9917,N_9978);
and UO_929 (O_929,N_9919,N_9915);
and UO_930 (O_930,N_9956,N_9955);
nand UO_931 (O_931,N_9974,N_9952);
or UO_932 (O_932,N_9963,N_9940);
nand UO_933 (O_933,N_9912,N_9904);
and UO_934 (O_934,N_9901,N_9991);
and UO_935 (O_935,N_9938,N_9971);
and UO_936 (O_936,N_9927,N_9970);
and UO_937 (O_937,N_9949,N_9950);
nand UO_938 (O_938,N_9928,N_9993);
nor UO_939 (O_939,N_9955,N_9986);
and UO_940 (O_940,N_9901,N_9990);
nor UO_941 (O_941,N_9997,N_9944);
or UO_942 (O_942,N_9955,N_9973);
nand UO_943 (O_943,N_9981,N_9996);
nor UO_944 (O_944,N_9998,N_9969);
and UO_945 (O_945,N_9976,N_9981);
and UO_946 (O_946,N_9953,N_9980);
nand UO_947 (O_947,N_9931,N_9963);
and UO_948 (O_948,N_9920,N_9903);
and UO_949 (O_949,N_9949,N_9982);
and UO_950 (O_950,N_9927,N_9910);
nand UO_951 (O_951,N_9917,N_9939);
or UO_952 (O_952,N_9976,N_9916);
nor UO_953 (O_953,N_9935,N_9981);
or UO_954 (O_954,N_9979,N_9963);
and UO_955 (O_955,N_9966,N_9919);
or UO_956 (O_956,N_9953,N_9948);
or UO_957 (O_957,N_9977,N_9945);
and UO_958 (O_958,N_9957,N_9905);
nand UO_959 (O_959,N_9986,N_9935);
nor UO_960 (O_960,N_9937,N_9997);
or UO_961 (O_961,N_9952,N_9980);
and UO_962 (O_962,N_9966,N_9969);
and UO_963 (O_963,N_9913,N_9942);
nand UO_964 (O_964,N_9920,N_9974);
nor UO_965 (O_965,N_9902,N_9965);
nor UO_966 (O_966,N_9901,N_9951);
and UO_967 (O_967,N_9930,N_9989);
nand UO_968 (O_968,N_9985,N_9903);
and UO_969 (O_969,N_9912,N_9918);
nand UO_970 (O_970,N_9963,N_9970);
nor UO_971 (O_971,N_9922,N_9988);
or UO_972 (O_972,N_9900,N_9924);
nand UO_973 (O_973,N_9936,N_9998);
and UO_974 (O_974,N_9912,N_9958);
or UO_975 (O_975,N_9914,N_9905);
nor UO_976 (O_976,N_9974,N_9993);
nand UO_977 (O_977,N_9995,N_9901);
or UO_978 (O_978,N_9907,N_9986);
or UO_979 (O_979,N_9922,N_9962);
and UO_980 (O_980,N_9901,N_9900);
or UO_981 (O_981,N_9990,N_9920);
nand UO_982 (O_982,N_9917,N_9926);
or UO_983 (O_983,N_9903,N_9973);
nand UO_984 (O_984,N_9993,N_9904);
nand UO_985 (O_985,N_9914,N_9919);
or UO_986 (O_986,N_9988,N_9924);
and UO_987 (O_987,N_9928,N_9967);
and UO_988 (O_988,N_9965,N_9979);
nand UO_989 (O_989,N_9939,N_9944);
nand UO_990 (O_990,N_9976,N_9940);
nand UO_991 (O_991,N_9973,N_9916);
or UO_992 (O_992,N_9980,N_9962);
or UO_993 (O_993,N_9910,N_9948);
nor UO_994 (O_994,N_9987,N_9950);
nand UO_995 (O_995,N_9920,N_9940);
nand UO_996 (O_996,N_9995,N_9916);
nor UO_997 (O_997,N_9905,N_9928);
or UO_998 (O_998,N_9908,N_9997);
nor UO_999 (O_999,N_9918,N_9932);
nand UO_1000 (O_1000,N_9973,N_9998);
or UO_1001 (O_1001,N_9912,N_9975);
nor UO_1002 (O_1002,N_9902,N_9979);
or UO_1003 (O_1003,N_9940,N_9957);
and UO_1004 (O_1004,N_9934,N_9966);
nand UO_1005 (O_1005,N_9950,N_9957);
nor UO_1006 (O_1006,N_9993,N_9988);
or UO_1007 (O_1007,N_9950,N_9913);
or UO_1008 (O_1008,N_9932,N_9944);
and UO_1009 (O_1009,N_9951,N_9954);
and UO_1010 (O_1010,N_9986,N_9989);
or UO_1011 (O_1011,N_9929,N_9943);
nor UO_1012 (O_1012,N_9908,N_9905);
or UO_1013 (O_1013,N_9991,N_9978);
or UO_1014 (O_1014,N_9947,N_9998);
or UO_1015 (O_1015,N_9969,N_9929);
and UO_1016 (O_1016,N_9961,N_9983);
or UO_1017 (O_1017,N_9933,N_9930);
and UO_1018 (O_1018,N_9920,N_9964);
and UO_1019 (O_1019,N_9907,N_9989);
and UO_1020 (O_1020,N_9962,N_9963);
or UO_1021 (O_1021,N_9979,N_9934);
nand UO_1022 (O_1022,N_9909,N_9974);
or UO_1023 (O_1023,N_9910,N_9921);
or UO_1024 (O_1024,N_9925,N_9981);
and UO_1025 (O_1025,N_9989,N_9955);
nand UO_1026 (O_1026,N_9912,N_9909);
nor UO_1027 (O_1027,N_9970,N_9961);
nand UO_1028 (O_1028,N_9905,N_9997);
nor UO_1029 (O_1029,N_9941,N_9962);
or UO_1030 (O_1030,N_9923,N_9916);
or UO_1031 (O_1031,N_9997,N_9949);
and UO_1032 (O_1032,N_9984,N_9992);
or UO_1033 (O_1033,N_9991,N_9981);
and UO_1034 (O_1034,N_9927,N_9973);
nand UO_1035 (O_1035,N_9971,N_9911);
nand UO_1036 (O_1036,N_9992,N_9959);
nand UO_1037 (O_1037,N_9933,N_9980);
nor UO_1038 (O_1038,N_9963,N_9952);
and UO_1039 (O_1039,N_9983,N_9913);
nand UO_1040 (O_1040,N_9932,N_9921);
nand UO_1041 (O_1041,N_9916,N_9925);
or UO_1042 (O_1042,N_9922,N_9935);
or UO_1043 (O_1043,N_9939,N_9959);
and UO_1044 (O_1044,N_9928,N_9985);
nor UO_1045 (O_1045,N_9983,N_9958);
nand UO_1046 (O_1046,N_9921,N_9902);
or UO_1047 (O_1047,N_9937,N_9950);
nor UO_1048 (O_1048,N_9930,N_9924);
or UO_1049 (O_1049,N_9943,N_9945);
and UO_1050 (O_1050,N_9921,N_9913);
nand UO_1051 (O_1051,N_9906,N_9923);
nand UO_1052 (O_1052,N_9999,N_9943);
nand UO_1053 (O_1053,N_9906,N_9977);
or UO_1054 (O_1054,N_9937,N_9995);
nand UO_1055 (O_1055,N_9962,N_9953);
nand UO_1056 (O_1056,N_9927,N_9906);
nand UO_1057 (O_1057,N_9996,N_9965);
and UO_1058 (O_1058,N_9993,N_9907);
nand UO_1059 (O_1059,N_9949,N_9981);
and UO_1060 (O_1060,N_9988,N_9964);
nor UO_1061 (O_1061,N_9955,N_9978);
nor UO_1062 (O_1062,N_9934,N_9988);
and UO_1063 (O_1063,N_9960,N_9942);
nand UO_1064 (O_1064,N_9981,N_9994);
nand UO_1065 (O_1065,N_9918,N_9958);
or UO_1066 (O_1066,N_9962,N_9979);
nand UO_1067 (O_1067,N_9912,N_9951);
and UO_1068 (O_1068,N_9973,N_9994);
nand UO_1069 (O_1069,N_9931,N_9945);
nand UO_1070 (O_1070,N_9976,N_9993);
or UO_1071 (O_1071,N_9998,N_9900);
nor UO_1072 (O_1072,N_9944,N_9914);
nand UO_1073 (O_1073,N_9943,N_9925);
nand UO_1074 (O_1074,N_9945,N_9946);
and UO_1075 (O_1075,N_9925,N_9931);
or UO_1076 (O_1076,N_9979,N_9931);
nor UO_1077 (O_1077,N_9991,N_9948);
nor UO_1078 (O_1078,N_9960,N_9907);
nor UO_1079 (O_1079,N_9936,N_9931);
nor UO_1080 (O_1080,N_9918,N_9922);
nand UO_1081 (O_1081,N_9978,N_9912);
or UO_1082 (O_1082,N_9970,N_9949);
nor UO_1083 (O_1083,N_9938,N_9904);
and UO_1084 (O_1084,N_9990,N_9991);
nand UO_1085 (O_1085,N_9941,N_9961);
nor UO_1086 (O_1086,N_9958,N_9916);
and UO_1087 (O_1087,N_9960,N_9957);
and UO_1088 (O_1088,N_9928,N_9901);
nand UO_1089 (O_1089,N_9964,N_9989);
nor UO_1090 (O_1090,N_9999,N_9921);
or UO_1091 (O_1091,N_9916,N_9900);
or UO_1092 (O_1092,N_9989,N_9977);
or UO_1093 (O_1093,N_9990,N_9965);
xnor UO_1094 (O_1094,N_9985,N_9943);
or UO_1095 (O_1095,N_9947,N_9984);
or UO_1096 (O_1096,N_9943,N_9935);
and UO_1097 (O_1097,N_9937,N_9981);
and UO_1098 (O_1098,N_9976,N_9954);
or UO_1099 (O_1099,N_9963,N_9992);
nand UO_1100 (O_1100,N_9964,N_9949);
nor UO_1101 (O_1101,N_9998,N_9945);
nand UO_1102 (O_1102,N_9974,N_9919);
nand UO_1103 (O_1103,N_9936,N_9941);
nand UO_1104 (O_1104,N_9907,N_9940);
or UO_1105 (O_1105,N_9946,N_9937);
and UO_1106 (O_1106,N_9968,N_9906);
nand UO_1107 (O_1107,N_9956,N_9962);
and UO_1108 (O_1108,N_9978,N_9915);
nand UO_1109 (O_1109,N_9977,N_9936);
or UO_1110 (O_1110,N_9979,N_9933);
and UO_1111 (O_1111,N_9964,N_9970);
nor UO_1112 (O_1112,N_9958,N_9919);
nand UO_1113 (O_1113,N_9977,N_9996);
and UO_1114 (O_1114,N_9929,N_9978);
or UO_1115 (O_1115,N_9975,N_9969);
or UO_1116 (O_1116,N_9979,N_9952);
nor UO_1117 (O_1117,N_9973,N_9948);
nor UO_1118 (O_1118,N_9971,N_9992);
and UO_1119 (O_1119,N_9917,N_9902);
and UO_1120 (O_1120,N_9942,N_9979);
and UO_1121 (O_1121,N_9928,N_9964);
or UO_1122 (O_1122,N_9912,N_9945);
nor UO_1123 (O_1123,N_9984,N_9998);
and UO_1124 (O_1124,N_9902,N_9993);
and UO_1125 (O_1125,N_9929,N_9913);
nor UO_1126 (O_1126,N_9929,N_9903);
and UO_1127 (O_1127,N_9950,N_9988);
or UO_1128 (O_1128,N_9943,N_9912);
or UO_1129 (O_1129,N_9961,N_9982);
and UO_1130 (O_1130,N_9952,N_9953);
or UO_1131 (O_1131,N_9985,N_9999);
nand UO_1132 (O_1132,N_9941,N_9994);
and UO_1133 (O_1133,N_9906,N_9913);
or UO_1134 (O_1134,N_9995,N_9958);
or UO_1135 (O_1135,N_9996,N_9903);
and UO_1136 (O_1136,N_9932,N_9993);
and UO_1137 (O_1137,N_9979,N_9924);
nor UO_1138 (O_1138,N_9904,N_9947);
nand UO_1139 (O_1139,N_9963,N_9997);
or UO_1140 (O_1140,N_9954,N_9946);
nor UO_1141 (O_1141,N_9920,N_9957);
or UO_1142 (O_1142,N_9927,N_9952);
nor UO_1143 (O_1143,N_9964,N_9900);
nand UO_1144 (O_1144,N_9996,N_9976);
nor UO_1145 (O_1145,N_9974,N_9900);
nor UO_1146 (O_1146,N_9949,N_9942);
and UO_1147 (O_1147,N_9963,N_9930);
and UO_1148 (O_1148,N_9988,N_9911);
nor UO_1149 (O_1149,N_9915,N_9952);
nand UO_1150 (O_1150,N_9981,N_9988);
and UO_1151 (O_1151,N_9988,N_9973);
xor UO_1152 (O_1152,N_9953,N_9915);
and UO_1153 (O_1153,N_9974,N_9987);
nor UO_1154 (O_1154,N_9946,N_9942);
nor UO_1155 (O_1155,N_9948,N_9941);
nor UO_1156 (O_1156,N_9983,N_9903);
and UO_1157 (O_1157,N_9951,N_9984);
and UO_1158 (O_1158,N_9946,N_9973);
nand UO_1159 (O_1159,N_9941,N_9929);
or UO_1160 (O_1160,N_9959,N_9993);
or UO_1161 (O_1161,N_9965,N_9907);
nand UO_1162 (O_1162,N_9960,N_9994);
or UO_1163 (O_1163,N_9913,N_9982);
nand UO_1164 (O_1164,N_9903,N_9976);
nor UO_1165 (O_1165,N_9953,N_9900);
nand UO_1166 (O_1166,N_9954,N_9990);
nor UO_1167 (O_1167,N_9984,N_9991);
and UO_1168 (O_1168,N_9933,N_9948);
or UO_1169 (O_1169,N_9978,N_9959);
nand UO_1170 (O_1170,N_9954,N_9995);
and UO_1171 (O_1171,N_9986,N_9916);
or UO_1172 (O_1172,N_9969,N_9968);
and UO_1173 (O_1173,N_9976,N_9942);
or UO_1174 (O_1174,N_9973,N_9912);
or UO_1175 (O_1175,N_9967,N_9958);
or UO_1176 (O_1176,N_9962,N_9929);
nor UO_1177 (O_1177,N_9931,N_9966);
nor UO_1178 (O_1178,N_9939,N_9992);
nor UO_1179 (O_1179,N_9922,N_9964);
nand UO_1180 (O_1180,N_9947,N_9949);
nor UO_1181 (O_1181,N_9918,N_9966);
nor UO_1182 (O_1182,N_9965,N_9926);
nor UO_1183 (O_1183,N_9918,N_9947);
nand UO_1184 (O_1184,N_9949,N_9924);
nand UO_1185 (O_1185,N_9963,N_9926);
nor UO_1186 (O_1186,N_9960,N_9934);
and UO_1187 (O_1187,N_9982,N_9986);
nor UO_1188 (O_1188,N_9951,N_9998);
or UO_1189 (O_1189,N_9932,N_9931);
nand UO_1190 (O_1190,N_9961,N_9936);
nor UO_1191 (O_1191,N_9916,N_9931);
and UO_1192 (O_1192,N_9945,N_9985);
nor UO_1193 (O_1193,N_9989,N_9923);
and UO_1194 (O_1194,N_9989,N_9926);
and UO_1195 (O_1195,N_9969,N_9912);
nand UO_1196 (O_1196,N_9921,N_9937);
or UO_1197 (O_1197,N_9963,N_9938);
nand UO_1198 (O_1198,N_9924,N_9958);
and UO_1199 (O_1199,N_9975,N_9943);
nor UO_1200 (O_1200,N_9904,N_9949);
and UO_1201 (O_1201,N_9944,N_9949);
and UO_1202 (O_1202,N_9982,N_9989);
and UO_1203 (O_1203,N_9978,N_9979);
or UO_1204 (O_1204,N_9914,N_9989);
and UO_1205 (O_1205,N_9930,N_9947);
nor UO_1206 (O_1206,N_9944,N_9918);
nand UO_1207 (O_1207,N_9997,N_9986);
nand UO_1208 (O_1208,N_9933,N_9972);
and UO_1209 (O_1209,N_9922,N_9977);
nor UO_1210 (O_1210,N_9950,N_9938);
nor UO_1211 (O_1211,N_9937,N_9999);
and UO_1212 (O_1212,N_9932,N_9968);
or UO_1213 (O_1213,N_9988,N_9919);
or UO_1214 (O_1214,N_9996,N_9990);
and UO_1215 (O_1215,N_9931,N_9973);
nor UO_1216 (O_1216,N_9979,N_9990);
or UO_1217 (O_1217,N_9933,N_9963);
nand UO_1218 (O_1218,N_9909,N_9970);
or UO_1219 (O_1219,N_9987,N_9935);
nor UO_1220 (O_1220,N_9913,N_9977);
nor UO_1221 (O_1221,N_9931,N_9975);
and UO_1222 (O_1222,N_9934,N_9955);
nand UO_1223 (O_1223,N_9982,N_9975);
nand UO_1224 (O_1224,N_9929,N_9900);
and UO_1225 (O_1225,N_9944,N_9904);
nor UO_1226 (O_1226,N_9979,N_9935);
and UO_1227 (O_1227,N_9978,N_9964);
xor UO_1228 (O_1228,N_9968,N_9924);
and UO_1229 (O_1229,N_9990,N_9985);
and UO_1230 (O_1230,N_9903,N_9961);
or UO_1231 (O_1231,N_9959,N_9986);
or UO_1232 (O_1232,N_9953,N_9959);
or UO_1233 (O_1233,N_9921,N_9988);
xnor UO_1234 (O_1234,N_9954,N_9970);
and UO_1235 (O_1235,N_9909,N_9939);
or UO_1236 (O_1236,N_9932,N_9952);
nand UO_1237 (O_1237,N_9971,N_9978);
xnor UO_1238 (O_1238,N_9996,N_9997);
nand UO_1239 (O_1239,N_9967,N_9993);
and UO_1240 (O_1240,N_9957,N_9922);
nand UO_1241 (O_1241,N_9906,N_9958);
nand UO_1242 (O_1242,N_9954,N_9957);
nand UO_1243 (O_1243,N_9947,N_9980);
or UO_1244 (O_1244,N_9926,N_9970);
nand UO_1245 (O_1245,N_9912,N_9972);
nor UO_1246 (O_1246,N_9967,N_9952);
or UO_1247 (O_1247,N_9958,N_9959);
or UO_1248 (O_1248,N_9923,N_9901);
and UO_1249 (O_1249,N_9910,N_9943);
and UO_1250 (O_1250,N_9942,N_9975);
and UO_1251 (O_1251,N_9909,N_9956);
and UO_1252 (O_1252,N_9975,N_9929);
and UO_1253 (O_1253,N_9950,N_9919);
or UO_1254 (O_1254,N_9931,N_9982);
or UO_1255 (O_1255,N_9979,N_9949);
and UO_1256 (O_1256,N_9905,N_9990);
and UO_1257 (O_1257,N_9933,N_9918);
nor UO_1258 (O_1258,N_9945,N_9957);
xnor UO_1259 (O_1259,N_9974,N_9980);
nor UO_1260 (O_1260,N_9950,N_9904);
or UO_1261 (O_1261,N_9902,N_9966);
and UO_1262 (O_1262,N_9907,N_9964);
nand UO_1263 (O_1263,N_9970,N_9930);
and UO_1264 (O_1264,N_9926,N_9984);
nand UO_1265 (O_1265,N_9976,N_9998);
and UO_1266 (O_1266,N_9964,N_9938);
nor UO_1267 (O_1267,N_9927,N_9949);
nor UO_1268 (O_1268,N_9907,N_9913);
nor UO_1269 (O_1269,N_9929,N_9906);
nor UO_1270 (O_1270,N_9944,N_9916);
and UO_1271 (O_1271,N_9901,N_9985);
and UO_1272 (O_1272,N_9944,N_9995);
and UO_1273 (O_1273,N_9959,N_9998);
nor UO_1274 (O_1274,N_9944,N_9955);
and UO_1275 (O_1275,N_9929,N_9910);
nor UO_1276 (O_1276,N_9983,N_9902);
nor UO_1277 (O_1277,N_9992,N_9974);
or UO_1278 (O_1278,N_9933,N_9935);
nor UO_1279 (O_1279,N_9939,N_9902);
or UO_1280 (O_1280,N_9936,N_9904);
or UO_1281 (O_1281,N_9907,N_9900);
and UO_1282 (O_1282,N_9931,N_9921);
and UO_1283 (O_1283,N_9906,N_9930);
or UO_1284 (O_1284,N_9909,N_9950);
nor UO_1285 (O_1285,N_9910,N_9963);
nor UO_1286 (O_1286,N_9946,N_9921);
nand UO_1287 (O_1287,N_9999,N_9933);
and UO_1288 (O_1288,N_9991,N_9937);
and UO_1289 (O_1289,N_9931,N_9977);
nor UO_1290 (O_1290,N_9967,N_9919);
and UO_1291 (O_1291,N_9953,N_9947);
and UO_1292 (O_1292,N_9921,N_9971);
or UO_1293 (O_1293,N_9916,N_9913);
nand UO_1294 (O_1294,N_9960,N_9991);
nand UO_1295 (O_1295,N_9982,N_9990);
or UO_1296 (O_1296,N_9996,N_9964);
nor UO_1297 (O_1297,N_9950,N_9999);
nand UO_1298 (O_1298,N_9917,N_9965);
nor UO_1299 (O_1299,N_9907,N_9936);
nor UO_1300 (O_1300,N_9951,N_9940);
and UO_1301 (O_1301,N_9963,N_9908);
nand UO_1302 (O_1302,N_9957,N_9973);
nor UO_1303 (O_1303,N_9995,N_9921);
and UO_1304 (O_1304,N_9915,N_9925);
nor UO_1305 (O_1305,N_9907,N_9939);
or UO_1306 (O_1306,N_9907,N_9919);
nand UO_1307 (O_1307,N_9990,N_9943);
nand UO_1308 (O_1308,N_9965,N_9966);
nor UO_1309 (O_1309,N_9907,N_9985);
nand UO_1310 (O_1310,N_9932,N_9983);
or UO_1311 (O_1311,N_9988,N_9977);
or UO_1312 (O_1312,N_9964,N_9934);
or UO_1313 (O_1313,N_9930,N_9939);
and UO_1314 (O_1314,N_9925,N_9920);
nor UO_1315 (O_1315,N_9986,N_9901);
or UO_1316 (O_1316,N_9997,N_9998);
nor UO_1317 (O_1317,N_9912,N_9928);
and UO_1318 (O_1318,N_9929,N_9990);
and UO_1319 (O_1319,N_9924,N_9925);
or UO_1320 (O_1320,N_9935,N_9942);
nand UO_1321 (O_1321,N_9976,N_9975);
nand UO_1322 (O_1322,N_9998,N_9980);
or UO_1323 (O_1323,N_9904,N_9948);
or UO_1324 (O_1324,N_9908,N_9925);
nor UO_1325 (O_1325,N_9972,N_9942);
nand UO_1326 (O_1326,N_9925,N_9982);
nor UO_1327 (O_1327,N_9953,N_9974);
and UO_1328 (O_1328,N_9969,N_9916);
or UO_1329 (O_1329,N_9937,N_9989);
and UO_1330 (O_1330,N_9931,N_9981);
or UO_1331 (O_1331,N_9904,N_9925);
nor UO_1332 (O_1332,N_9949,N_9935);
or UO_1333 (O_1333,N_9961,N_9928);
and UO_1334 (O_1334,N_9943,N_9973);
and UO_1335 (O_1335,N_9969,N_9977);
nor UO_1336 (O_1336,N_9986,N_9979);
nand UO_1337 (O_1337,N_9944,N_9951);
nand UO_1338 (O_1338,N_9963,N_9927);
nand UO_1339 (O_1339,N_9939,N_9936);
and UO_1340 (O_1340,N_9945,N_9936);
nor UO_1341 (O_1341,N_9924,N_9953);
nand UO_1342 (O_1342,N_9953,N_9996);
or UO_1343 (O_1343,N_9982,N_9988);
nor UO_1344 (O_1344,N_9977,N_9938);
or UO_1345 (O_1345,N_9942,N_9953);
nor UO_1346 (O_1346,N_9937,N_9993);
or UO_1347 (O_1347,N_9908,N_9986);
and UO_1348 (O_1348,N_9987,N_9928);
nand UO_1349 (O_1349,N_9950,N_9952);
nor UO_1350 (O_1350,N_9904,N_9929);
nand UO_1351 (O_1351,N_9981,N_9977);
or UO_1352 (O_1352,N_9980,N_9945);
nand UO_1353 (O_1353,N_9957,N_9955);
and UO_1354 (O_1354,N_9931,N_9900);
nor UO_1355 (O_1355,N_9953,N_9909);
nand UO_1356 (O_1356,N_9966,N_9956);
or UO_1357 (O_1357,N_9944,N_9934);
or UO_1358 (O_1358,N_9980,N_9902);
nor UO_1359 (O_1359,N_9975,N_9944);
nand UO_1360 (O_1360,N_9994,N_9963);
and UO_1361 (O_1361,N_9992,N_9962);
nor UO_1362 (O_1362,N_9913,N_9911);
and UO_1363 (O_1363,N_9975,N_9972);
and UO_1364 (O_1364,N_9904,N_9923);
and UO_1365 (O_1365,N_9903,N_9993);
nand UO_1366 (O_1366,N_9937,N_9920);
nand UO_1367 (O_1367,N_9942,N_9940);
and UO_1368 (O_1368,N_9909,N_9951);
nor UO_1369 (O_1369,N_9973,N_9986);
nor UO_1370 (O_1370,N_9933,N_9943);
nor UO_1371 (O_1371,N_9976,N_9928);
or UO_1372 (O_1372,N_9911,N_9909);
nor UO_1373 (O_1373,N_9914,N_9998);
nor UO_1374 (O_1374,N_9915,N_9987);
nor UO_1375 (O_1375,N_9946,N_9960);
or UO_1376 (O_1376,N_9982,N_9970);
nor UO_1377 (O_1377,N_9982,N_9985);
nor UO_1378 (O_1378,N_9933,N_9969);
and UO_1379 (O_1379,N_9995,N_9993);
nand UO_1380 (O_1380,N_9960,N_9906);
nand UO_1381 (O_1381,N_9975,N_9914);
or UO_1382 (O_1382,N_9964,N_9991);
and UO_1383 (O_1383,N_9968,N_9973);
and UO_1384 (O_1384,N_9998,N_9932);
and UO_1385 (O_1385,N_9949,N_9946);
or UO_1386 (O_1386,N_9952,N_9978);
nor UO_1387 (O_1387,N_9904,N_9913);
nor UO_1388 (O_1388,N_9941,N_9993);
nand UO_1389 (O_1389,N_9964,N_9950);
or UO_1390 (O_1390,N_9964,N_9912);
nor UO_1391 (O_1391,N_9905,N_9981);
or UO_1392 (O_1392,N_9964,N_9993);
nand UO_1393 (O_1393,N_9996,N_9912);
and UO_1394 (O_1394,N_9982,N_9907);
nand UO_1395 (O_1395,N_9959,N_9983);
or UO_1396 (O_1396,N_9941,N_9919);
nand UO_1397 (O_1397,N_9908,N_9954);
or UO_1398 (O_1398,N_9904,N_9999);
or UO_1399 (O_1399,N_9968,N_9942);
and UO_1400 (O_1400,N_9986,N_9957);
or UO_1401 (O_1401,N_9928,N_9978);
nand UO_1402 (O_1402,N_9974,N_9997);
and UO_1403 (O_1403,N_9928,N_9970);
or UO_1404 (O_1404,N_9922,N_9928);
or UO_1405 (O_1405,N_9920,N_9993);
and UO_1406 (O_1406,N_9915,N_9970);
nor UO_1407 (O_1407,N_9907,N_9984);
or UO_1408 (O_1408,N_9997,N_9970);
nand UO_1409 (O_1409,N_9955,N_9910);
or UO_1410 (O_1410,N_9900,N_9963);
and UO_1411 (O_1411,N_9941,N_9995);
or UO_1412 (O_1412,N_9933,N_9905);
xor UO_1413 (O_1413,N_9968,N_9915);
and UO_1414 (O_1414,N_9914,N_9968);
and UO_1415 (O_1415,N_9993,N_9938);
nand UO_1416 (O_1416,N_9924,N_9999);
nand UO_1417 (O_1417,N_9958,N_9905);
or UO_1418 (O_1418,N_9980,N_9928);
and UO_1419 (O_1419,N_9947,N_9999);
nand UO_1420 (O_1420,N_9999,N_9938);
or UO_1421 (O_1421,N_9935,N_9936);
and UO_1422 (O_1422,N_9961,N_9989);
nor UO_1423 (O_1423,N_9937,N_9923);
nor UO_1424 (O_1424,N_9970,N_9935);
or UO_1425 (O_1425,N_9987,N_9925);
and UO_1426 (O_1426,N_9900,N_9969);
nor UO_1427 (O_1427,N_9937,N_9902);
nand UO_1428 (O_1428,N_9985,N_9978);
or UO_1429 (O_1429,N_9904,N_9980);
nor UO_1430 (O_1430,N_9944,N_9964);
nand UO_1431 (O_1431,N_9921,N_9973);
and UO_1432 (O_1432,N_9905,N_9940);
or UO_1433 (O_1433,N_9988,N_9986);
nand UO_1434 (O_1434,N_9940,N_9909);
nor UO_1435 (O_1435,N_9982,N_9933);
nor UO_1436 (O_1436,N_9914,N_9951);
nand UO_1437 (O_1437,N_9906,N_9920);
or UO_1438 (O_1438,N_9978,N_9983);
or UO_1439 (O_1439,N_9923,N_9990);
nand UO_1440 (O_1440,N_9996,N_9978);
and UO_1441 (O_1441,N_9927,N_9959);
and UO_1442 (O_1442,N_9960,N_9925);
nand UO_1443 (O_1443,N_9983,N_9979);
nand UO_1444 (O_1444,N_9946,N_9976);
or UO_1445 (O_1445,N_9935,N_9918);
and UO_1446 (O_1446,N_9934,N_9939);
or UO_1447 (O_1447,N_9950,N_9939);
nor UO_1448 (O_1448,N_9984,N_9922);
and UO_1449 (O_1449,N_9997,N_9933);
or UO_1450 (O_1450,N_9970,N_9904);
and UO_1451 (O_1451,N_9925,N_9928);
nand UO_1452 (O_1452,N_9921,N_9960);
nand UO_1453 (O_1453,N_9921,N_9908);
nand UO_1454 (O_1454,N_9997,N_9953);
nand UO_1455 (O_1455,N_9933,N_9991);
or UO_1456 (O_1456,N_9902,N_9936);
nand UO_1457 (O_1457,N_9926,N_9914);
nor UO_1458 (O_1458,N_9988,N_9909);
nand UO_1459 (O_1459,N_9948,N_9987);
or UO_1460 (O_1460,N_9965,N_9941);
nand UO_1461 (O_1461,N_9966,N_9951);
or UO_1462 (O_1462,N_9923,N_9910);
nand UO_1463 (O_1463,N_9950,N_9935);
and UO_1464 (O_1464,N_9936,N_9952);
and UO_1465 (O_1465,N_9933,N_9971);
nor UO_1466 (O_1466,N_9993,N_9954);
and UO_1467 (O_1467,N_9972,N_9948);
nand UO_1468 (O_1468,N_9940,N_9945);
and UO_1469 (O_1469,N_9992,N_9903);
and UO_1470 (O_1470,N_9969,N_9973);
xor UO_1471 (O_1471,N_9924,N_9905);
nor UO_1472 (O_1472,N_9913,N_9994);
or UO_1473 (O_1473,N_9915,N_9973);
nor UO_1474 (O_1474,N_9908,N_9974);
and UO_1475 (O_1475,N_9922,N_9939);
and UO_1476 (O_1476,N_9990,N_9986);
nand UO_1477 (O_1477,N_9977,N_9904);
nor UO_1478 (O_1478,N_9978,N_9925);
or UO_1479 (O_1479,N_9967,N_9963);
or UO_1480 (O_1480,N_9982,N_9906);
nand UO_1481 (O_1481,N_9944,N_9950);
nand UO_1482 (O_1482,N_9970,N_9958);
nor UO_1483 (O_1483,N_9995,N_9969);
nand UO_1484 (O_1484,N_9916,N_9978);
and UO_1485 (O_1485,N_9931,N_9968);
and UO_1486 (O_1486,N_9947,N_9983);
nor UO_1487 (O_1487,N_9941,N_9949);
nor UO_1488 (O_1488,N_9901,N_9910);
nor UO_1489 (O_1489,N_9970,N_9957);
nor UO_1490 (O_1490,N_9940,N_9964);
or UO_1491 (O_1491,N_9962,N_9933);
or UO_1492 (O_1492,N_9905,N_9913);
nand UO_1493 (O_1493,N_9960,N_9969);
nand UO_1494 (O_1494,N_9908,N_9952);
and UO_1495 (O_1495,N_9997,N_9984);
nand UO_1496 (O_1496,N_9947,N_9924);
and UO_1497 (O_1497,N_9907,N_9910);
and UO_1498 (O_1498,N_9999,N_9965);
and UO_1499 (O_1499,N_9946,N_9916);
endmodule