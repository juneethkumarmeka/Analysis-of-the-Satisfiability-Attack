module basic_1500_15000_2000_30_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_715,In_818);
xnor U1 (N_1,In_231,In_849);
nand U2 (N_2,In_1113,In_124);
and U3 (N_3,In_1088,In_1216);
xnor U4 (N_4,In_352,In_114);
nor U5 (N_5,In_1299,In_1364);
nand U6 (N_6,In_462,In_50);
nand U7 (N_7,In_932,In_1473);
xnor U8 (N_8,In_996,In_831);
xnor U9 (N_9,In_1097,In_890);
nand U10 (N_10,In_269,In_1380);
nor U11 (N_11,In_125,In_493);
and U12 (N_12,In_11,In_395);
and U13 (N_13,In_116,In_0);
and U14 (N_14,In_1213,In_931);
nor U15 (N_15,In_1076,In_596);
nand U16 (N_16,In_320,In_633);
xnor U17 (N_17,In_180,In_1203);
or U18 (N_18,In_323,In_1198);
xor U19 (N_19,In_214,In_693);
nand U20 (N_20,In_168,In_1145);
and U21 (N_21,In_1115,In_461);
xor U22 (N_22,In_452,In_432);
nor U23 (N_23,In_1008,In_1469);
nand U24 (N_24,In_1067,In_1383);
or U25 (N_25,In_193,In_1238);
xnor U26 (N_26,In_799,In_1495);
or U27 (N_27,In_1459,In_296);
nor U28 (N_28,In_1189,In_120);
nor U29 (N_29,In_143,In_920);
and U30 (N_30,In_601,In_979);
nand U31 (N_31,In_328,In_454);
or U32 (N_32,In_83,In_367);
xnor U33 (N_33,In_271,In_638);
and U34 (N_34,In_1241,In_872);
xnor U35 (N_35,In_413,In_962);
or U36 (N_36,In_1131,In_665);
nor U37 (N_37,In_43,In_924);
xnor U38 (N_38,In_1389,In_527);
and U39 (N_39,In_115,In_986);
and U40 (N_40,In_769,In_933);
or U41 (N_41,In_541,In_1298);
xor U42 (N_42,In_1318,In_426);
nand U43 (N_43,In_412,In_772);
nand U44 (N_44,In_1490,In_1212);
and U45 (N_45,In_163,In_128);
xnor U46 (N_46,In_257,In_105);
nand U47 (N_47,In_443,In_36);
nor U48 (N_48,In_842,In_347);
or U49 (N_49,In_1056,In_1262);
xnor U50 (N_50,In_20,In_1043);
xor U51 (N_51,In_390,In_976);
nor U52 (N_52,In_262,In_91);
and U53 (N_53,In_546,In_1351);
nor U54 (N_54,In_167,In_247);
and U55 (N_55,In_189,In_1379);
xor U56 (N_56,In_1227,In_1183);
xnor U57 (N_57,In_978,In_716);
nand U58 (N_58,In_1108,In_683);
and U59 (N_59,In_204,In_1423);
nand U60 (N_60,In_349,In_343);
nand U61 (N_61,In_1005,In_302);
and U62 (N_62,In_1020,In_261);
nand U63 (N_63,In_833,In_748);
or U64 (N_64,In_1180,In_1271);
nand U65 (N_65,In_1051,In_297);
or U66 (N_66,In_642,In_1498);
xnor U67 (N_67,In_1477,In_1416);
nand U68 (N_68,In_511,In_517);
xor U69 (N_69,In_687,In_942);
nand U70 (N_70,In_844,In_1362);
xor U71 (N_71,In_1480,In_441);
xnor U72 (N_72,In_1047,In_709);
nor U73 (N_73,In_1392,In_1059);
or U74 (N_74,In_508,In_1060);
and U75 (N_75,In_640,In_937);
and U76 (N_76,In_578,In_795);
nor U77 (N_77,In_170,In_492);
nand U78 (N_78,In_593,In_202);
and U79 (N_79,In_1363,In_156);
or U80 (N_80,In_55,In_308);
or U81 (N_81,In_845,In_641);
nand U82 (N_82,In_568,In_1019);
nor U83 (N_83,In_1100,In_628);
and U84 (N_84,In_377,In_1329);
xor U85 (N_85,In_474,In_782);
xnor U86 (N_86,In_67,In_957);
nand U87 (N_87,In_1127,In_538);
and U88 (N_88,In_57,In_1280);
and U89 (N_89,In_736,In_1099);
or U90 (N_90,In_817,In_65);
nor U91 (N_91,In_164,In_1120);
or U92 (N_92,In_659,In_564);
or U93 (N_93,In_526,In_109);
nand U94 (N_94,In_188,In_652);
nand U95 (N_95,In_1319,In_900);
nor U96 (N_96,In_1058,In_543);
and U97 (N_97,In_1201,In_371);
or U98 (N_98,In_569,In_958);
nor U99 (N_99,In_1394,In_746);
and U100 (N_100,In_1235,In_944);
nand U101 (N_101,In_1309,In_518);
xor U102 (N_102,In_1007,In_960);
nor U103 (N_103,In_397,In_745);
nor U104 (N_104,In_1234,In_419);
or U105 (N_105,In_1179,In_949);
xnor U106 (N_106,In_1103,In_350);
nand U107 (N_107,In_1378,In_557);
or U108 (N_108,In_74,In_941);
nand U109 (N_109,In_704,In_485);
or U110 (N_110,In_946,In_206);
nand U111 (N_111,In_528,In_322);
xor U112 (N_112,In_1288,In_353);
nand U113 (N_113,In_759,In_918);
nand U114 (N_114,In_467,In_574);
nand U115 (N_115,In_1429,In_737);
and U116 (N_116,In_1455,In_1426);
xnor U117 (N_117,In_270,In_1432);
or U118 (N_118,In_398,In_1149);
or U119 (N_119,In_649,In_815);
nand U120 (N_120,In_1037,In_1221);
xnor U121 (N_121,In_103,In_32);
or U122 (N_122,In_314,In_263);
xnor U123 (N_123,In_827,In_486);
nand U124 (N_124,In_436,In_161);
and U125 (N_125,In_331,In_404);
nand U126 (N_126,In_977,In_893);
nand U127 (N_127,In_101,In_1320);
nor U128 (N_128,In_273,In_1018);
and U129 (N_129,In_1011,In_51);
xnor U130 (N_130,In_916,In_137);
xor U131 (N_131,In_1292,In_555);
or U132 (N_132,In_494,In_1031);
nor U133 (N_133,In_7,In_1286);
or U134 (N_134,In_1489,In_1200);
nor U135 (N_135,In_1461,In_656);
or U136 (N_136,In_104,In_368);
nand U137 (N_137,In_1285,In_1369);
or U138 (N_138,In_1410,In_847);
xnor U139 (N_139,In_1282,In_973);
and U140 (N_140,In_1358,In_1366);
xnor U141 (N_141,In_39,In_18);
xnor U142 (N_142,In_1193,In_293);
and U143 (N_143,In_165,In_282);
xor U144 (N_144,In_325,In_1014);
or U145 (N_145,In_340,In_1417);
nor U146 (N_146,In_27,In_95);
and U147 (N_147,In_657,In_599);
xor U148 (N_148,In_773,In_972);
and U149 (N_149,In_1090,In_295);
xor U150 (N_150,In_850,In_1481);
xnor U151 (N_151,In_778,In_1162);
nand U152 (N_152,In_1470,In_1028);
xor U153 (N_153,In_46,In_765);
or U154 (N_154,In_283,In_1073);
or U155 (N_155,In_1025,In_917);
xor U156 (N_156,In_1077,In_252);
xor U157 (N_157,In_1098,In_97);
xnor U158 (N_158,In_739,In_240);
nor U159 (N_159,In_524,In_460);
xnor U160 (N_160,In_1419,In_581);
and U161 (N_161,In_808,In_249);
and U162 (N_162,In_729,In_311);
nor U163 (N_163,In_255,In_1096);
nor U164 (N_164,In_768,In_667);
nand U165 (N_165,In_1012,In_663);
xor U166 (N_166,In_44,In_1451);
or U167 (N_167,In_854,In_330);
xnor U168 (N_168,In_1085,In_786);
or U169 (N_169,In_459,In_1218);
nor U170 (N_170,In_926,In_600);
and U171 (N_171,In_439,In_38);
or U172 (N_172,In_747,In_911);
xor U173 (N_173,In_1258,In_514);
or U174 (N_174,In_939,In_1377);
and U175 (N_175,In_619,In_157);
or U176 (N_176,In_691,In_732);
xor U177 (N_177,In_530,In_411);
or U178 (N_178,In_521,In_199);
and U179 (N_179,In_807,In_981);
nor U180 (N_180,In_315,In_1340);
or U181 (N_181,In_562,In_1348);
xor U182 (N_182,In_1121,In_914);
nand U183 (N_183,In_1424,In_212);
and U184 (N_184,In_242,In_93);
or U185 (N_185,In_658,In_1317);
nor U186 (N_186,In_1467,In_783);
xnor U187 (N_187,In_185,In_25);
nand U188 (N_188,In_119,In_66);
or U189 (N_189,In_561,In_87);
and U190 (N_190,In_1443,In_402);
nor U191 (N_191,In_162,In_999);
nor U192 (N_192,In_724,In_618);
or U193 (N_193,In_1324,In_805);
or U194 (N_194,In_1344,In_1223);
nor U195 (N_195,In_1204,In_130);
xnor U196 (N_196,In_552,In_396);
or U197 (N_197,In_1386,In_545);
xor U198 (N_198,In_1341,In_1261);
xnor U199 (N_199,In_415,In_1174);
and U200 (N_200,In_1370,In_1035);
or U201 (N_201,In_146,In_586);
xnor U202 (N_202,In_339,In_1045);
nor U203 (N_203,In_582,In_414);
or U204 (N_204,In_158,In_1231);
nor U205 (N_205,In_626,In_1185);
or U206 (N_206,In_810,In_757);
and U207 (N_207,In_305,In_1316);
xnor U208 (N_208,In_1297,In_13);
nor U209 (N_209,In_312,In_338);
nor U210 (N_210,In_1214,In_653);
nand U211 (N_211,In_356,In_394);
or U212 (N_212,In_708,In_896);
nor U213 (N_213,In_536,In_1175);
nand U214 (N_214,In_506,In_442);
xnor U215 (N_215,In_49,In_664);
xor U216 (N_216,In_1034,In_381);
and U217 (N_217,In_1053,In_1273);
nand U218 (N_218,In_673,In_151);
and U219 (N_219,In_1301,In_1430);
or U220 (N_220,In_479,In_15);
and U221 (N_221,In_42,In_1491);
nor U222 (N_222,In_1163,In_567);
nand U223 (N_223,In_672,In_852);
or U224 (N_224,In_31,In_1474);
nor U225 (N_225,In_816,In_1);
nor U226 (N_226,In_1146,In_478);
nor U227 (N_227,In_1381,In_28);
nor U228 (N_228,In_868,In_47);
nor U229 (N_229,In_1006,In_1478);
or U230 (N_230,In_970,In_217);
nor U231 (N_231,In_856,In_1062);
nor U232 (N_232,In_440,In_329);
nor U233 (N_233,In_1119,In_286);
nand U234 (N_234,In_76,In_264);
and U235 (N_235,In_1251,In_630);
xor U236 (N_236,In_294,In_621);
nor U237 (N_237,In_908,In_209);
nor U238 (N_238,In_370,In_1061);
xor U239 (N_239,In_1281,In_316);
or U240 (N_240,In_826,In_1448);
nor U241 (N_241,In_602,In_989);
and U242 (N_242,In_554,In_435);
or U243 (N_243,In_1173,In_1194);
nand U244 (N_244,In_186,In_821);
and U245 (N_245,In_71,In_1274);
and U246 (N_246,In_935,In_1052);
and U247 (N_247,In_741,In_1220);
and U248 (N_248,In_1009,In_288);
and U249 (N_249,In_1303,In_1411);
or U250 (N_250,In_1081,In_605);
xnor U251 (N_251,In_752,In_934);
nor U252 (N_252,In_738,In_1326);
or U253 (N_253,In_1456,In_1249);
nand U254 (N_254,In_481,In_496);
nand U255 (N_255,In_207,In_225);
and U256 (N_256,In_6,In_532);
nand U257 (N_257,In_614,In_1256);
and U258 (N_258,In_1078,In_1315);
xnor U259 (N_259,In_111,In_690);
or U260 (N_260,In_874,In_1476);
xnor U261 (N_261,In_409,In_516);
and U262 (N_262,In_774,In_112);
nor U263 (N_263,In_1265,In_851);
and U264 (N_264,In_505,In_1391);
nand U265 (N_265,In_434,In_155);
or U266 (N_266,In_985,In_837);
xor U267 (N_267,In_80,In_1295);
xor U268 (N_268,In_813,In_1493);
nand U269 (N_269,In_455,In_603);
xnor U270 (N_270,In_451,In_430);
and U271 (N_271,In_686,In_241);
xnor U272 (N_272,In_1046,In_775);
and U273 (N_273,In_1475,In_1217);
nor U274 (N_274,In_950,In_814);
nand U275 (N_275,In_332,In_131);
nand U276 (N_276,In_210,In_141);
nand U277 (N_277,In_902,In_608);
nor U278 (N_278,In_533,In_859);
or U279 (N_279,In_871,In_123);
and U280 (N_280,In_1016,In_401);
or U281 (N_281,In_488,In_268);
nand U282 (N_282,In_750,In_246);
nand U283 (N_283,In_1437,In_853);
nor U284 (N_284,In_1130,In_243);
and U285 (N_285,In_895,In_1397);
xor U286 (N_286,In_174,In_735);
nor U287 (N_287,In_1433,In_706);
xor U288 (N_288,In_346,In_565);
and U289 (N_289,In_607,In_366);
or U290 (N_290,In_54,In_1404);
nor U291 (N_291,In_21,In_983);
xor U292 (N_292,In_731,In_1065);
or U293 (N_293,In_969,In_1118);
nand U294 (N_294,In_433,In_287);
or U295 (N_295,In_1134,In_1486);
nor U296 (N_296,In_1278,In_1312);
and U297 (N_297,In_56,In_139);
xor U298 (N_298,In_583,In_447);
nor U299 (N_299,In_1070,In_472);
xnor U300 (N_300,In_1346,In_509);
nor U301 (N_301,In_364,In_1359);
xnor U302 (N_302,In_1188,In_613);
or U303 (N_303,In_1181,In_437);
or U304 (N_304,In_444,In_360);
nor U305 (N_305,In_448,In_113);
nand U306 (N_306,In_886,In_830);
nand U307 (N_307,In_232,In_936);
xnor U308 (N_308,In_1440,In_881);
or U309 (N_309,In_326,In_1004);
and U310 (N_310,In_839,In_682);
or U311 (N_311,In_1355,In_635);
nand U312 (N_312,In_779,In_1393);
nor U313 (N_313,In_726,In_542);
or U314 (N_314,In_449,In_727);
nand U315 (N_315,In_1465,In_1349);
or U316 (N_316,In_882,In_1087);
or U317 (N_317,In_3,In_354);
and U318 (N_318,In_1039,In_375);
or U319 (N_319,In_1139,In_1350);
nor U320 (N_320,In_655,In_1205);
xnor U321 (N_321,In_1029,In_947);
xor U322 (N_322,In_766,In_1157);
and U323 (N_323,In_846,In_878);
xor U324 (N_324,In_1387,In_1409);
xor U325 (N_325,In_798,In_389);
or U326 (N_326,In_840,In_843);
nand U327 (N_327,In_169,In_913);
nor U328 (N_328,In_1184,In_1372);
nand U329 (N_329,In_1026,In_34);
xnor U330 (N_330,In_1352,In_387);
and U331 (N_331,In_1401,In_597);
nand U332 (N_332,In_61,In_645);
nor U333 (N_333,In_12,In_1255);
nand U334 (N_334,In_560,In_800);
nand U335 (N_335,In_928,In_1178);
and U336 (N_336,In_258,In_1164);
nand U337 (N_337,In_733,In_1044);
nor U338 (N_338,In_1225,In_1343);
nand U339 (N_339,In_964,In_1445);
and U340 (N_340,In_1150,In_1027);
nor U341 (N_341,In_577,In_259);
and U342 (N_342,In_860,In_1311);
or U343 (N_343,In_617,In_1290);
nand U344 (N_344,In_889,In_198);
or U345 (N_345,In_749,In_281);
xor U346 (N_346,In_877,In_1017);
and U347 (N_347,In_1237,In_227);
nand U348 (N_348,In_1219,In_1243);
xor U349 (N_349,In_876,In_224);
nand U350 (N_350,In_1226,In_905);
and U351 (N_351,In_1142,In_388);
nand U352 (N_352,In_811,In_927);
or U353 (N_353,In_802,In_1293);
or U354 (N_354,In_147,In_1095);
nor U355 (N_355,In_719,In_1291);
nand U356 (N_356,In_723,In_78);
and U357 (N_357,In_420,In_1335);
xnor U358 (N_358,In_812,In_4);
nand U359 (N_359,In_674,In_68);
or U360 (N_360,In_1159,In_176);
nand U361 (N_361,In_535,In_668);
xor U362 (N_362,In_179,In_776);
or U363 (N_363,In_1123,In_471);
or U364 (N_364,In_804,In_963);
nor U365 (N_365,In_1487,In_1483);
and U366 (N_366,In_1013,In_1384);
xnor U367 (N_367,In_828,In_1395);
nand U368 (N_368,In_337,In_152);
or U369 (N_369,In_1327,In_1105);
or U370 (N_370,In_987,In_292);
and U371 (N_371,In_943,In_575);
and U372 (N_372,In_1257,In_1460);
xor U373 (N_373,In_760,In_457);
xnor U374 (N_374,In_205,In_961);
nor U375 (N_375,In_37,In_196);
nor U376 (N_376,In_498,In_429);
and U377 (N_377,In_1038,In_1289);
or U378 (N_378,In_159,In_675);
and U379 (N_379,In_679,In_1406);
nor U380 (N_380,In_373,In_763);
or U381 (N_381,In_1252,In_1064);
nor U382 (N_382,In_797,In_1434);
nand U383 (N_383,In_938,In_787);
nor U384 (N_384,In_1233,In_740);
and U385 (N_385,In_317,In_265);
xor U386 (N_386,In_698,In_1023);
or U387 (N_387,In_299,In_559);
nand U388 (N_388,In_507,In_90);
and U389 (N_389,In_476,In_278);
xor U390 (N_390,In_1403,In_475);
xor U391 (N_391,In_721,In_873);
nand U392 (N_392,In_445,In_1361);
nand U393 (N_393,In_399,In_275);
xor U394 (N_394,In_324,In_149);
and U395 (N_395,In_707,In_1463);
and U396 (N_396,In_1464,In_688);
xor U397 (N_397,In_1144,In_615);
xnor U398 (N_398,In_1439,In_362);
nand U399 (N_399,In_1151,In_2);
nand U400 (N_400,In_1496,In_997);
or U401 (N_401,In_450,In_660);
nor U402 (N_402,In_1137,In_758);
nand U403 (N_403,In_525,In_885);
xor U404 (N_404,In_702,In_801);
nand U405 (N_405,In_579,In_512);
xnor U406 (N_406,In_1072,In_24);
or U407 (N_407,In_796,In_534);
nor U408 (N_408,In_1453,In_138);
nand U409 (N_409,In_611,In_1328);
nand U410 (N_410,In_922,In_117);
or U411 (N_411,In_883,In_1068);
nand U412 (N_412,In_753,In_233);
xor U413 (N_413,In_629,In_197);
xnor U414 (N_414,In_403,In_1360);
and U415 (N_415,In_866,In_235);
and U416 (N_416,In_1152,In_1240);
nor U417 (N_417,In_1066,In_1356);
or U418 (N_418,In_428,In_1172);
nand U419 (N_419,In_650,In_248);
or U420 (N_420,In_1040,In_284);
nand U421 (N_421,In_697,In_728);
nand U422 (N_422,In_722,In_19);
and U423 (N_423,In_572,In_72);
and U424 (N_424,In_393,In_245);
nand U425 (N_425,In_10,In_861);
nand U426 (N_426,In_648,In_834);
nand U427 (N_427,In_1260,In_971);
and U428 (N_428,In_118,In_1420);
xnor U429 (N_429,In_544,In_1024);
nand U430 (N_430,In_540,In_888);
nor U431 (N_431,In_819,In_624);
nor U432 (N_432,In_784,In_504);
nor U433 (N_433,In_487,In_1306);
nor U434 (N_434,In_1075,In_73);
nor U435 (N_435,In_1171,In_953);
nand U436 (N_436,In_495,In_1375);
or U437 (N_437,In_107,In_792);
nor U438 (N_438,In_1135,In_345);
nand U439 (N_439,In_1036,In_154);
or U440 (N_440,In_1147,In_580);
and U441 (N_441,In_1071,In_1484);
nand U442 (N_442,In_267,In_955);
xor U443 (N_443,In_190,In_134);
xnor U444 (N_444,In_1266,In_1457);
and U445 (N_445,In_453,In_1472);
nand U446 (N_446,In_1000,In_374);
xnor U447 (N_447,In_695,In_576);
or U448 (N_448,In_14,In_636);
xnor U449 (N_449,In_178,In_994);
nor U450 (N_450,In_385,In_662);
or U451 (N_451,In_1229,In_623);
xor U452 (N_452,In_1143,In_216);
or U453 (N_453,In_1048,In_1167);
xor U454 (N_454,In_952,In_993);
nand U455 (N_455,In_1405,In_1055);
xnor U456 (N_456,In_1471,In_677);
xor U457 (N_457,In_1452,In_898);
nor U458 (N_458,In_1094,In_1368);
xor U459 (N_459,In_725,In_408);
and U460 (N_460,In_670,In_1160);
nand U461 (N_461,In_86,In_372);
nand U462 (N_462,In_1435,In_145);
and U463 (N_463,In_1425,In_1371);
and U464 (N_464,In_836,In_1187);
xor U465 (N_465,In_771,In_627);
nor U466 (N_466,In_1248,In_22);
or U467 (N_467,In_761,In_502);
nand U468 (N_468,In_809,In_1365);
xor U469 (N_469,In_1296,In_785);
nand U470 (N_470,In_465,In_1140);
xnor U471 (N_471,In_1279,In_228);
nor U472 (N_472,In_604,In_1331);
nand U473 (N_473,In_975,In_200);
nor U474 (N_474,In_1110,In_1268);
nand U475 (N_475,In_201,In_678);
nand U476 (N_476,In_1314,In_589);
xor U477 (N_477,In_1101,In_220);
or U478 (N_478,In_864,In_857);
xnor U479 (N_479,In_260,In_710);
nand U480 (N_480,In_718,In_274);
xnor U481 (N_481,In_469,In_218);
and U482 (N_482,In_754,In_1333);
and U483 (N_483,In_1126,In_48);
or U484 (N_484,In_223,In_907);
nand U485 (N_485,In_82,In_912);
xor U486 (N_486,In_192,In_1148);
nor U487 (N_487,In_1414,In_643);
or U488 (N_488,In_1186,In_229);
nand U489 (N_489,In_239,In_215);
and U490 (N_490,In_53,In_1427);
xnor U491 (N_491,In_714,In_1367);
or U492 (N_492,In_1116,In_696);
nand U493 (N_493,In_171,In_187);
xor U494 (N_494,In_887,In_684);
nor U495 (N_495,In_1211,In_26);
nand U496 (N_496,In_751,In_1128);
or U497 (N_497,In_1267,In_1089);
or U498 (N_498,In_135,In_1402);
nor U499 (N_499,In_1165,In_803);
nand U500 (N_500,N_448,N_328);
or U501 (N_501,In_1300,N_14);
nor U502 (N_502,In_1057,In_822);
nor U503 (N_503,In_276,N_199);
xnor U504 (N_504,In_1373,In_921);
and U505 (N_505,In_23,N_467);
and U506 (N_506,N_116,In_1376);
nand U507 (N_507,N_281,N_206);
nand U508 (N_508,In_1276,N_287);
and U509 (N_509,N_490,In_92);
nand U510 (N_510,In_1250,In_427);
xor U511 (N_511,N_275,In_29);
and U512 (N_512,In_1155,In_5);
nand U513 (N_513,N_369,In_790);
xnor U514 (N_514,In_237,N_355);
or U515 (N_515,In_81,In_341);
nor U516 (N_516,In_637,In_1499);
and U517 (N_517,In_129,In_184);
nand U518 (N_518,N_412,In_1308);
nand U519 (N_519,N_175,In_304);
nand U520 (N_520,N_115,In_909);
nor U521 (N_521,In_1353,In_342);
and U522 (N_522,In_625,N_273);
xnor U523 (N_523,In_333,N_141);
nand U524 (N_524,In_906,N_26);
nand U525 (N_525,In_551,N_425);
or U526 (N_526,N_395,N_112);
or U527 (N_527,N_219,N_2);
nand U528 (N_528,In_318,In_558);
and U529 (N_529,In_1228,N_233);
or U530 (N_530,N_479,In_140);
xnor U531 (N_531,N_41,In_418);
nand U532 (N_532,In_894,In_421);
nor U533 (N_533,N_133,N_27);
or U534 (N_534,N_209,N_13);
or U535 (N_535,N_295,N_347);
and U536 (N_536,In_1136,In_301);
nor U537 (N_537,In_1153,In_1283);
or U538 (N_538,N_52,N_452);
or U539 (N_539,In_182,N_53);
nor U540 (N_540,In_1001,In_954);
and U541 (N_541,N_57,N_393);
or U542 (N_542,N_335,N_284);
xnor U543 (N_543,In_556,N_407);
nand U544 (N_544,In_392,In_319);
and U545 (N_545,N_414,N_247);
and U546 (N_546,In_483,In_221);
nand U547 (N_547,In_1449,N_211);
nand U548 (N_548,N_391,In_386);
nand U549 (N_549,N_110,In_272);
or U550 (N_550,N_411,N_362);
and U551 (N_551,In_794,In_666);
or U552 (N_552,N_82,In_929);
xor U553 (N_553,In_1330,In_948);
or U554 (N_554,N_92,N_270);
and U555 (N_555,N_150,N_371);
nand U556 (N_556,In_309,N_152);
or U557 (N_557,N_188,In_1454);
nand U558 (N_558,N_450,N_221);
or U559 (N_559,In_835,N_288);
or U560 (N_560,N_75,In_510);
and U561 (N_561,N_471,N_195);
or U562 (N_562,N_239,In_620);
or U563 (N_563,N_103,In_1015);
xnor U564 (N_564,N_144,In_40);
and U565 (N_565,N_40,N_336);
xor U566 (N_566,N_317,N_132);
or U567 (N_567,N_79,N_463);
and U568 (N_568,N_334,In_334);
and U569 (N_569,N_482,N_404);
and U570 (N_570,N_260,N_280);
nand U571 (N_571,In_405,In_1422);
xnor U572 (N_572,In_1342,In_69);
nand U573 (N_573,In_1245,N_217);
or U574 (N_574,In_838,In_355);
nand U575 (N_575,N_55,N_315);
or U576 (N_576,In_1442,N_262);
nand U577 (N_577,In_606,In_1458);
xnor U578 (N_578,In_148,N_227);
and U579 (N_579,In_501,N_164);
or U580 (N_580,N_86,N_166);
nand U581 (N_581,In_891,In_1177);
xnor U582 (N_582,N_396,In_1322);
nand U583 (N_583,N_7,In_1041);
nor U584 (N_584,In_689,N_184);
or U585 (N_585,N_171,N_392);
nand U586 (N_586,In_897,In_1338);
and U587 (N_587,N_87,In_595);
xor U588 (N_588,In_1206,In_1441);
nor U589 (N_589,In_965,N_248);
or U590 (N_590,N_470,N_366);
nor U591 (N_591,In_351,N_201);
xnor U592 (N_592,In_244,N_240);
or U593 (N_593,N_465,In_256);
nor U594 (N_594,In_869,N_76);
nand U595 (N_595,In_122,N_230);
or U596 (N_596,N_106,In_1166);
and U597 (N_597,N_89,In_1310);
and U598 (N_598,N_121,N_160);
nand U599 (N_599,N_486,In_213);
or U600 (N_600,N_489,In_644);
nor U601 (N_601,In_1158,In_855);
and U602 (N_602,In_307,N_337);
and U603 (N_603,N_36,N_378);
nand U604 (N_604,In_862,In_175);
nand U605 (N_605,N_182,In_410);
nor U606 (N_606,N_309,N_491);
nand U607 (N_607,In_1138,N_462);
and U608 (N_608,In_500,N_135);
xnor U609 (N_609,In_1450,In_407);
xnor U610 (N_610,N_481,In_880);
nand U611 (N_611,In_548,N_173);
or U612 (N_612,N_72,N_15);
xor U613 (N_613,N_29,N_226);
and U614 (N_614,N_460,In_132);
and U615 (N_615,In_160,In_858);
nand U616 (N_616,N_348,N_494);
xor U617 (N_617,In_925,In_1446);
or U618 (N_618,N_267,N_332);
nor U619 (N_619,In_669,N_360);
and U620 (N_620,In_376,N_314);
and U621 (N_621,N_350,In_1197);
nand U622 (N_622,N_299,In_98);
nor U623 (N_623,In_1385,N_399);
or U624 (N_624,N_11,N_458);
and U625 (N_625,N_220,In_1284);
and U626 (N_626,N_422,In_96);
and U627 (N_627,In_1002,N_138);
nand U628 (N_628,N_434,N_415);
nand U629 (N_629,N_157,In_1334);
or U630 (N_630,In_519,In_357);
nor U631 (N_631,N_456,N_397);
nor U632 (N_632,N_234,In_875);
or U633 (N_633,N_134,N_214);
nor U634 (N_634,In_1468,N_18);
or U635 (N_635,In_742,N_418);
xor U636 (N_636,In_1191,In_100);
xnor U637 (N_637,N_60,In_219);
xnor U638 (N_638,In_1253,In_867);
and U639 (N_639,In_191,N_417);
nand U640 (N_640,In_289,N_105);
nor U641 (N_641,In_870,In_1054);
nand U642 (N_642,In_503,In_75);
nor U643 (N_643,In_959,In_425);
xor U644 (N_644,N_437,N_96);
and U645 (N_645,In_1347,N_374);
nand U646 (N_646,In_590,In_651);
and U647 (N_647,In_121,N_194);
or U648 (N_648,In_923,N_68);
and U649 (N_649,N_421,N_438);
nand U650 (N_650,N_322,N_444);
xnor U651 (N_651,N_114,In_150);
and U652 (N_652,N_3,In_1208);
nor U653 (N_653,N_236,In_1270);
nand U654 (N_654,In_1337,In_609);
xnor U655 (N_655,In_458,N_99);
xor U656 (N_656,In_730,In_254);
and U657 (N_657,In_1325,N_216);
xor U658 (N_658,N_1,In_1438);
nor U659 (N_659,N_210,N_222);
or U660 (N_660,N_340,In_464);
or U661 (N_661,In_1336,N_232);
and U662 (N_662,In_904,In_181);
nor U663 (N_663,In_1156,In_195);
xor U664 (N_664,N_451,In_823);
xor U665 (N_665,In_41,In_1003);
nor U666 (N_666,N_376,In_1345);
nand U667 (N_667,In_711,In_285);
xnor U668 (N_668,N_163,N_388);
nor U669 (N_669,In_832,In_1091);
nand U670 (N_670,In_685,N_282);
nand U671 (N_671,In_764,In_344);
nor U672 (N_672,In_8,In_358);
or U673 (N_673,N_442,In_1321);
nor U674 (N_674,In_1125,In_1112);
and U675 (N_675,N_174,N_276);
nor U676 (N_676,In_592,N_148);
or U677 (N_677,N_263,In_1210);
xnor U678 (N_678,In_491,N_413);
or U679 (N_679,N_384,In_133);
and U680 (N_680,N_145,In_1170);
and U681 (N_681,In_136,N_101);
nand U682 (N_682,In_1354,In_522);
or U683 (N_683,N_58,In_1244);
nand U684 (N_684,N_264,In_701);
or U685 (N_685,In_879,N_454);
or U686 (N_686,N_126,In_829);
and U687 (N_687,N_139,In_253);
nand U688 (N_688,N_176,N_303);
or U689 (N_689,N_290,N_375);
or U690 (N_690,N_237,N_429);
nor U691 (N_691,In_379,In_88);
xnor U692 (N_692,N_402,N_159);
and U693 (N_693,In_1161,In_984);
nor U694 (N_694,In_1107,In_1010);
and U695 (N_695,N_44,In_369);
nand U696 (N_696,In_313,N_178);
and U697 (N_697,In_99,In_661);
or U698 (N_698,N_202,N_56);
xnor U699 (N_699,N_50,In_303);
xor U700 (N_700,N_488,N_377);
or U701 (N_701,N_311,N_153);
nand U702 (N_702,In_30,In_468);
xor U703 (N_703,In_1242,N_365);
nand U704 (N_704,N_228,N_351);
xnor U705 (N_705,In_52,N_266);
or U706 (N_706,N_468,In_234);
xor U707 (N_707,In_1421,N_107);
and U708 (N_708,N_190,N_88);
or U709 (N_709,In_1083,N_416);
nand U710 (N_710,N_243,In_1398);
and U711 (N_711,N_66,In_788);
and U712 (N_712,In_365,N_231);
xnor U713 (N_713,In_820,In_1129);
nor U714 (N_714,N_492,N_272);
or U715 (N_715,N_238,In_824);
or U716 (N_716,N_331,In_1169);
xor U717 (N_717,In_734,In_1462);
nand U718 (N_718,In_335,N_394);
nor U719 (N_719,N_131,N_271);
and U720 (N_720,In_529,N_123);
nor U721 (N_721,N_119,N_93);
or U722 (N_722,N_136,N_358);
or U723 (N_723,In_1399,In_1132);
nand U724 (N_724,In_300,N_324);
nand U725 (N_725,In_1492,N_95);
nor U726 (N_726,N_251,In_990);
xor U727 (N_727,In_489,In_612);
xor U728 (N_728,N_191,N_496);
xnor U729 (N_729,In_1497,N_155);
xnor U730 (N_730,In_35,In_473);
and U731 (N_731,N_212,N_170);
xor U732 (N_732,In_646,In_238);
nor U733 (N_733,N_10,In_378);
nor U734 (N_734,N_330,In_1190);
and U735 (N_735,N_17,N_80);
xnor U736 (N_736,N_229,N_71);
or U737 (N_737,In_361,N_23);
nand U738 (N_738,In_1154,In_585);
nor U739 (N_739,In_1133,N_363);
nor U740 (N_740,N_449,In_59);
and U741 (N_741,In_632,In_676);
xor U742 (N_742,N_25,In_951);
nand U743 (N_743,N_278,In_762);
nor U744 (N_744,In_417,N_259);
or U745 (N_745,In_520,N_424);
or U746 (N_746,N_147,In_1049);
xnor U747 (N_747,N_8,In_1408);
nor U748 (N_748,N_167,In_1230);
or U749 (N_749,N_300,N_297);
nand U750 (N_750,In_848,In_1199);
nor U751 (N_751,In_1259,In_1141);
and U752 (N_752,N_59,In_424);
and U753 (N_753,In_1323,N_91);
nor U754 (N_754,N_258,In_1114);
nor U755 (N_755,N_69,N_30);
nand U756 (N_756,N_84,In_639);
nor U757 (N_757,In_974,In_982);
and U758 (N_758,N_51,In_781);
nor U759 (N_759,In_968,N_398);
nor U760 (N_760,N_325,In_482);
xnor U761 (N_761,N_341,In_910);
xnor U762 (N_762,N_24,In_102);
or U763 (N_763,N_291,In_703);
and U764 (N_764,In_566,In_1222);
or U765 (N_765,In_1168,In_1224);
and U766 (N_766,N_447,In_166);
and U767 (N_767,In_85,N_129);
or U768 (N_768,N_373,In_380);
or U769 (N_769,In_1428,In_110);
or U770 (N_770,N_380,In_172);
nor U771 (N_771,N_181,In_1232);
and U772 (N_772,N_361,N_39);
nand U773 (N_773,N_254,N_130);
nand U774 (N_774,In_446,N_98);
nor U775 (N_775,N_323,In_60);
or U776 (N_776,N_345,In_456);
and U777 (N_777,In_1415,N_480);
nor U778 (N_778,N_446,In_327);
and U779 (N_779,N_9,In_865);
or U780 (N_780,N_484,N_168);
and U781 (N_781,N_339,In_1122);
nand U782 (N_782,N_242,In_1307);
or U783 (N_783,N_349,N_149);
nor U784 (N_784,In_634,In_694);
nand U785 (N_785,In_549,In_1215);
and U786 (N_786,N_277,In_251);
and U787 (N_787,In_1272,N_257);
nand U788 (N_788,In_1079,In_1413);
or U789 (N_789,N_35,N_83);
nor U790 (N_790,In_903,N_62);
or U791 (N_791,In_1069,N_285);
xnor U792 (N_792,N_74,N_370);
nor U793 (N_793,N_180,N_473);
nor U794 (N_794,In_967,N_70);
or U795 (N_795,In_142,In_1332);
xor U796 (N_796,In_919,N_431);
and U797 (N_797,N_120,In_1080);
nor U798 (N_798,In_539,In_553);
or U799 (N_799,In_126,In_584);
and U800 (N_800,In_692,In_1304);
and U801 (N_801,In_1275,In_789);
or U802 (N_802,N_198,N_124);
nand U803 (N_803,In_884,N_61);
xnor U804 (N_804,N_78,In_610);
nand U805 (N_805,N_102,N_165);
and U806 (N_806,N_476,In_966);
xor U807 (N_807,N_483,N_307);
xnor U808 (N_808,N_357,In_194);
or U809 (N_809,N_122,In_523);
and U810 (N_810,N_256,In_1022);
nand U811 (N_811,N_296,N_321);
and U812 (N_812,N_205,N_162);
or U813 (N_813,In_1313,N_245);
nor U814 (N_814,N_31,N_386);
and U815 (N_815,N_372,N_241);
xnor U816 (N_816,In_290,N_493);
nand U817 (N_817,In_713,N_22);
nor U818 (N_818,N_77,N_464);
nand U819 (N_819,N_499,N_32);
nand U820 (N_820,N_128,In_998);
and U821 (N_821,In_631,N_403);
xor U822 (N_822,In_306,N_200);
nand U823 (N_823,N_364,In_1418);
xor U824 (N_824,In_1196,In_1396);
or U825 (N_825,In_1466,N_37);
and U826 (N_826,In_1074,In_348);
nor U827 (N_827,N_253,N_154);
nand U828 (N_828,In_230,In_63);
xor U829 (N_829,In_1182,In_1269);
nor U830 (N_830,In_956,In_1412);
nor U831 (N_831,N_192,N_65);
xor U832 (N_832,In_108,In_1192);
or U833 (N_833,In_1106,N_189);
xor U834 (N_834,N_85,N_432);
xnor U835 (N_835,N_118,N_109);
and U836 (N_836,N_433,In_321);
xor U837 (N_837,In_515,In_980);
xor U838 (N_838,N_410,N_383);
nand U839 (N_839,N_430,N_343);
nor U840 (N_840,In_277,N_283);
and U841 (N_841,In_743,In_298);
nor U842 (N_842,In_470,In_1082);
and U843 (N_843,N_104,In_384);
and U844 (N_844,In_945,N_354);
and U845 (N_845,In_563,N_252);
nand U846 (N_846,In_431,N_63);
and U847 (N_847,In_1479,N_409);
nand U848 (N_848,In_571,N_218);
and U849 (N_849,N_169,N_387);
nand U850 (N_850,In_1236,In_222);
xnor U851 (N_851,In_863,N_111);
nor U852 (N_852,N_320,In_591);
xnor U853 (N_853,In_1263,In_777);
and U854 (N_854,N_440,N_156);
and U855 (N_855,In_587,N_466);
nor U856 (N_856,N_33,In_17);
xor U857 (N_857,N_367,N_47);
and U858 (N_858,N_478,In_1050);
and U859 (N_859,In_1287,N_151);
xor U860 (N_860,N_474,N_203);
and U861 (N_861,In_1388,N_475);
nand U862 (N_862,In_1494,N_34);
or U863 (N_863,N_261,N_333);
nand U864 (N_864,N_183,In_1374);
nand U865 (N_865,N_196,N_289);
or U866 (N_866,In_477,N_45);
and U867 (N_867,N_389,In_767);
or U868 (N_868,In_1339,N_305);
xnor U869 (N_869,N_319,In_363);
and U870 (N_870,In_310,N_477);
nor U871 (N_871,N_326,In_780);
or U872 (N_872,In_588,In_423);
xor U873 (N_873,N_274,N_301);
nor U874 (N_874,In_484,In_416);
and U875 (N_875,N_406,N_143);
and U876 (N_876,In_1209,N_423);
nor U877 (N_877,N_279,N_381);
or U878 (N_878,In_279,In_79);
or U879 (N_879,N_441,N_304);
and U880 (N_880,N_64,N_485);
xor U881 (N_881,N_385,N_428);
or U882 (N_882,N_81,In_1447);
and U883 (N_883,N_461,In_988);
or U884 (N_884,N_28,In_1431);
nand U885 (N_885,N_400,N_265);
and U886 (N_886,N_137,In_992);
xnor U887 (N_887,In_654,In_570);
nor U888 (N_888,In_899,N_46);
and U889 (N_889,In_94,N_408);
xnor U890 (N_890,N_187,N_308);
nor U891 (N_891,N_67,N_353);
or U892 (N_892,N_140,N_439);
or U893 (N_893,In_1195,In_62);
nand U894 (N_894,N_435,N_459);
and U895 (N_895,N_292,N_312);
and U896 (N_896,N_207,N_329);
nand U897 (N_897,N_249,In_1436);
xnor U898 (N_898,In_756,N_38);
nand U899 (N_899,In_236,In_1086);
nand U900 (N_900,N_4,In_1390);
nand U901 (N_901,N_177,In_1117);
or U902 (N_902,N_204,In_466);
or U903 (N_903,In_400,N_108);
xnor U904 (N_904,In_173,N_498);
and U905 (N_905,In_699,In_1111);
nor U906 (N_906,N_294,N_172);
and U907 (N_907,In_744,In_995);
xnor U908 (N_908,N_0,In_717);
xor U909 (N_909,In_1032,In_1246);
xor U910 (N_910,In_1109,N_495);
or U911 (N_911,In_291,N_223);
nor U912 (N_912,In_1302,N_401);
and U913 (N_913,N_338,In_594);
xnor U914 (N_914,N_94,In_70);
xnor U915 (N_915,In_671,In_382);
and U916 (N_916,In_1239,In_892);
and U917 (N_917,N_235,N_146);
xor U918 (N_918,In_622,N_193);
xor U919 (N_919,N_73,N_359);
or U920 (N_920,In_1444,N_352);
and U921 (N_921,In_1294,In_1030);
or U922 (N_922,N_327,N_250);
or U923 (N_923,In_106,In_1207);
or U924 (N_924,In_901,In_755);
and U925 (N_925,N_100,In_841);
nor U926 (N_926,In_647,In_16);
xnor U927 (N_927,In_1104,N_342);
or U928 (N_928,In_1176,In_770);
or U929 (N_929,In_1254,N_19);
and U930 (N_930,N_286,N_346);
and U931 (N_931,In_1400,N_298);
and U932 (N_932,N_472,In_705);
and U933 (N_933,In_1021,N_208);
xnor U934 (N_934,In_127,N_127);
and U935 (N_935,In_359,In_208);
or U936 (N_936,In_406,In_712);
and U937 (N_937,N_246,N_268);
nor U938 (N_938,N_43,In_1482);
xor U939 (N_939,In_1305,N_419);
nor U940 (N_940,In_720,N_269);
nor U941 (N_941,N_318,N_213);
and U942 (N_942,N_469,In_203);
and U943 (N_943,In_680,N_427);
xor U944 (N_944,In_700,N_186);
nand U945 (N_945,In_177,N_445);
xnor U946 (N_946,In_463,In_383);
nand U947 (N_947,In_1247,N_405);
or U948 (N_948,In_33,In_1277);
xnor U949 (N_949,In_537,In_499);
or U950 (N_950,N_90,In_211);
and U951 (N_951,In_1033,In_183);
nor U952 (N_952,N_443,In_1382);
nand U953 (N_953,In_573,In_144);
or U954 (N_954,N_16,N_197);
nor U955 (N_955,In_1092,N_225);
or U956 (N_956,N_158,N_215);
nand U957 (N_957,N_390,In_915);
or U958 (N_958,In_1093,N_306);
or U959 (N_959,N_244,In_422);
nor U960 (N_960,N_54,In_84);
or U961 (N_961,N_42,N_21);
and U962 (N_962,N_379,In_1488);
nor U963 (N_963,N_316,In_598);
nor U964 (N_964,N_436,In_64);
and U965 (N_965,N_457,N_310);
and U966 (N_966,In_550,In_497);
xnor U967 (N_967,In_438,N_455);
and U968 (N_968,N_497,In_480);
nor U969 (N_969,In_940,In_250);
nand U970 (N_970,In_1485,In_1357);
or U971 (N_971,N_356,In_513);
and U972 (N_972,In_266,N_185);
and U973 (N_973,In_1102,N_302);
or U974 (N_974,N_487,N_113);
nor U975 (N_975,N_224,In_531);
xor U976 (N_976,N_20,In_806);
xnor U977 (N_977,N_344,N_12);
nand U978 (N_978,In_1407,In_547);
or U979 (N_979,In_45,In_681);
nor U980 (N_980,N_6,In_226);
nor U981 (N_981,N_48,In_930);
xor U982 (N_982,N_142,In_791);
nor U983 (N_983,N_179,In_58);
xnor U984 (N_984,N_255,In_1042);
nand U985 (N_985,In_280,N_161);
nand U986 (N_986,N_5,In_153);
and U987 (N_987,N_125,In_991);
nor U988 (N_988,N_313,N_368);
nand U989 (N_989,In_1202,N_382);
or U990 (N_990,N_420,In_1124);
xor U991 (N_991,In_391,In_793);
and U992 (N_992,In_9,In_825);
xnor U993 (N_993,N_117,In_490);
nand U994 (N_994,In_616,In_89);
nand U995 (N_995,N_426,N_97);
nor U996 (N_996,In_1084,In_1264);
nand U997 (N_997,N_49,In_77);
nor U998 (N_998,N_453,In_336);
xor U999 (N_999,In_1063,N_293);
nor U1000 (N_1000,N_938,N_555);
nand U1001 (N_1001,N_830,N_846);
nand U1002 (N_1002,N_918,N_585);
nand U1003 (N_1003,N_863,N_602);
nand U1004 (N_1004,N_685,N_996);
xor U1005 (N_1005,N_536,N_875);
nand U1006 (N_1006,N_777,N_856);
nand U1007 (N_1007,N_772,N_642);
xnor U1008 (N_1008,N_668,N_535);
and U1009 (N_1009,N_864,N_519);
or U1010 (N_1010,N_925,N_929);
xor U1011 (N_1011,N_596,N_537);
and U1012 (N_1012,N_647,N_865);
or U1013 (N_1013,N_747,N_968);
nand U1014 (N_1014,N_569,N_713);
nand U1015 (N_1015,N_898,N_505);
xnor U1016 (N_1016,N_852,N_890);
nor U1017 (N_1017,N_802,N_581);
and U1018 (N_1018,N_733,N_708);
nand U1019 (N_1019,N_711,N_834);
xor U1020 (N_1020,N_832,N_965);
nor U1021 (N_1021,N_945,N_994);
xnor U1022 (N_1022,N_526,N_667);
nor U1023 (N_1023,N_690,N_600);
nor U1024 (N_1024,N_648,N_958);
xor U1025 (N_1025,N_880,N_934);
xor U1026 (N_1026,N_551,N_946);
and U1027 (N_1027,N_807,N_594);
nand U1028 (N_1028,N_528,N_847);
or U1029 (N_1029,N_913,N_513);
nor U1030 (N_1030,N_564,N_984);
nand U1031 (N_1031,N_557,N_988);
and U1032 (N_1032,N_921,N_666);
nor U1033 (N_1033,N_631,N_952);
and U1034 (N_1034,N_565,N_768);
or U1035 (N_1035,N_756,N_656);
nor U1036 (N_1036,N_509,N_781);
and U1037 (N_1037,N_607,N_917);
and U1038 (N_1038,N_548,N_974);
and U1039 (N_1039,N_858,N_961);
and U1040 (N_1040,N_637,N_819);
xor U1041 (N_1041,N_811,N_997);
and U1042 (N_1042,N_905,N_910);
nor U1043 (N_1043,N_661,N_771);
xnor U1044 (N_1044,N_823,N_870);
nand U1045 (N_1045,N_599,N_533);
nand U1046 (N_1046,N_887,N_953);
and U1047 (N_1047,N_680,N_609);
xnor U1048 (N_1048,N_833,N_787);
xnor U1049 (N_1049,N_963,N_543);
and U1050 (N_1050,N_757,N_588);
nor U1051 (N_1051,N_818,N_545);
nor U1052 (N_1052,N_684,N_542);
xnor U1053 (N_1053,N_553,N_576);
nor U1054 (N_1054,N_877,N_512);
and U1055 (N_1055,N_665,N_595);
xor U1056 (N_1056,N_770,N_794);
nor U1057 (N_1057,N_605,N_638);
nor U1058 (N_1058,N_897,N_891);
or U1059 (N_1059,N_980,N_502);
or U1060 (N_1060,N_730,N_698);
nor U1061 (N_1061,N_854,N_696);
nand U1062 (N_1062,N_704,N_939);
nand U1063 (N_1063,N_981,N_635);
or U1064 (N_1064,N_957,N_892);
or U1065 (N_1065,N_866,N_650);
nor U1066 (N_1066,N_759,N_572);
nor U1067 (N_1067,N_644,N_790);
and U1068 (N_1068,N_949,N_702);
nor U1069 (N_1069,N_669,N_797);
nand U1070 (N_1070,N_828,N_804);
nand U1071 (N_1071,N_796,N_641);
and U1072 (N_1072,N_950,N_738);
nand U1073 (N_1073,N_568,N_710);
xnor U1074 (N_1074,N_622,N_620);
xnor U1075 (N_1075,N_932,N_752);
nand U1076 (N_1076,N_853,N_560);
and U1077 (N_1077,N_817,N_839);
and U1078 (N_1078,N_829,N_671);
xor U1079 (N_1079,N_709,N_989);
xnor U1080 (N_1080,N_900,N_619);
and U1081 (N_1081,N_598,N_908);
xnor U1082 (N_1082,N_612,N_523);
and U1083 (N_1083,N_753,N_646);
nor U1084 (N_1084,N_906,N_559);
and U1085 (N_1085,N_538,N_597);
xnor U1086 (N_1086,N_792,N_960);
nor U1087 (N_1087,N_741,N_601);
xnor U1088 (N_1088,N_577,N_675);
nor U1089 (N_1089,N_987,N_860);
xor U1090 (N_1090,N_527,N_774);
nor U1091 (N_1091,N_888,N_783);
nand U1092 (N_1092,N_521,N_937);
or U1093 (N_1093,N_979,N_697);
or U1094 (N_1094,N_746,N_922);
xnor U1095 (N_1095,N_676,N_862);
and U1096 (N_1096,N_649,N_517);
or U1097 (N_1097,N_975,N_861);
or U1098 (N_1098,N_558,N_749);
and U1099 (N_1099,N_972,N_782);
nand U1100 (N_1100,N_687,N_820);
or U1101 (N_1101,N_885,N_943);
and U1102 (N_1102,N_844,N_552);
or U1103 (N_1103,N_522,N_529);
xor U1104 (N_1104,N_876,N_789);
nor U1105 (N_1105,N_948,N_688);
nor U1106 (N_1106,N_745,N_580);
xnor U1107 (N_1107,N_705,N_769);
nand U1108 (N_1108,N_652,N_567);
xnor U1109 (N_1109,N_714,N_775);
and U1110 (N_1110,N_902,N_767);
nor U1111 (N_1111,N_813,N_742);
nor U1112 (N_1112,N_722,N_840);
and U1113 (N_1113,N_928,N_663);
or U1114 (N_1114,N_779,N_983);
nor U1115 (N_1115,N_806,N_843);
nand U1116 (N_1116,N_603,N_848);
or U1117 (N_1117,N_748,N_682);
nand U1118 (N_1118,N_679,N_608);
and U1119 (N_1119,N_563,N_624);
nand U1120 (N_1120,N_578,N_626);
and U1121 (N_1121,N_546,N_604);
nor U1122 (N_1122,N_901,N_985);
or U1123 (N_1123,N_850,N_993);
xnor U1124 (N_1124,N_579,N_916);
xnor U1125 (N_1125,N_694,N_801);
and U1126 (N_1126,N_867,N_911);
xor U1127 (N_1127,N_732,N_670);
nor U1128 (N_1128,N_912,N_630);
nor U1129 (N_1129,N_763,N_808);
nand U1130 (N_1130,N_785,N_821);
nor U1131 (N_1131,N_969,N_971);
xnor U1132 (N_1132,N_510,N_758);
nand U1133 (N_1133,N_584,N_793);
nand U1134 (N_1134,N_762,N_628);
nand U1135 (N_1135,N_524,N_904);
nor U1136 (N_1136,N_532,N_959);
or U1137 (N_1137,N_681,N_511);
and U1138 (N_1138,N_838,N_723);
xnor U1139 (N_1139,N_506,N_837);
nor U1140 (N_1140,N_926,N_719);
nor U1141 (N_1141,N_999,N_909);
or U1142 (N_1142,N_773,N_991);
nor U1143 (N_1143,N_566,N_924);
nand U1144 (N_1144,N_692,N_973);
and U1145 (N_1145,N_874,N_664);
xor U1146 (N_1146,N_835,N_695);
nand U1147 (N_1147,N_586,N_618);
or U1148 (N_1148,N_734,N_990);
nand U1149 (N_1149,N_872,N_744);
xor U1150 (N_1150,N_977,N_556);
nand U1151 (N_1151,N_970,N_955);
nor U1152 (N_1152,N_729,N_583);
nor U1153 (N_1153,N_855,N_776);
nand U1154 (N_1154,N_658,N_549);
or U1155 (N_1155,N_755,N_851);
nor U1156 (N_1156,N_815,N_613);
or U1157 (N_1157,N_919,N_589);
xnor U1158 (N_1158,N_899,N_896);
xnor U1159 (N_1159,N_812,N_700);
and U1160 (N_1160,N_824,N_992);
or U1161 (N_1161,N_822,N_800);
nor U1162 (N_1162,N_761,N_716);
and U1163 (N_1163,N_998,N_873);
nor U1164 (N_1164,N_930,N_544);
nand U1165 (N_1165,N_515,N_814);
nor U1166 (N_1166,N_884,N_582);
and U1167 (N_1167,N_942,N_726);
or U1168 (N_1168,N_751,N_691);
nand U1169 (N_1169,N_606,N_501);
nor U1170 (N_1170,N_657,N_780);
nand U1171 (N_1171,N_660,N_640);
nor U1172 (N_1172,N_720,N_889);
xor U1173 (N_1173,N_736,N_786);
nand U1174 (N_1174,N_575,N_615);
and U1175 (N_1175,N_805,N_743);
or U1176 (N_1176,N_827,N_740);
or U1177 (N_1177,N_520,N_845);
nor U1178 (N_1178,N_868,N_857);
nor U1179 (N_1179,N_735,N_718);
or U1180 (N_1180,N_571,N_914);
nor U1181 (N_1181,N_895,N_784);
nor U1182 (N_1182,N_616,N_662);
or U1183 (N_1183,N_707,N_962);
nor U1184 (N_1184,N_915,N_645);
and U1185 (N_1185,N_689,N_659);
and U1186 (N_1186,N_803,N_504);
nand U1187 (N_1187,N_530,N_500);
xor U1188 (N_1188,N_514,N_636);
and U1189 (N_1189,N_653,N_570);
or U1190 (N_1190,N_825,N_561);
and U1191 (N_1191,N_923,N_715);
xor U1192 (N_1192,N_587,N_655);
nand U1193 (N_1193,N_701,N_550);
or U1194 (N_1194,N_964,N_764);
nor U1195 (N_1195,N_788,N_562);
xnor U1196 (N_1196,N_778,N_826);
and U1197 (N_1197,N_677,N_810);
nand U1198 (N_1198,N_731,N_739);
nor U1199 (N_1199,N_750,N_590);
xnor U1200 (N_1200,N_886,N_651);
xnor U1201 (N_1201,N_927,N_816);
or U1202 (N_1202,N_516,N_634);
nand U1203 (N_1203,N_693,N_956);
and U1204 (N_1204,N_933,N_686);
or U1205 (N_1205,N_920,N_712);
xor U1206 (N_1206,N_754,N_760);
xnor U1207 (N_1207,N_869,N_625);
or U1208 (N_1208,N_508,N_944);
nand U1209 (N_1209,N_976,N_507);
nor U1210 (N_1210,N_765,N_831);
xnor U1211 (N_1211,N_931,N_672);
or U1212 (N_1212,N_525,N_725);
or U1213 (N_1213,N_639,N_881);
nor U1214 (N_1214,N_574,N_503);
and U1215 (N_1215,N_699,N_982);
xnor U1216 (N_1216,N_614,N_703);
xor U1217 (N_1217,N_883,N_683);
nand U1218 (N_1218,N_632,N_842);
nor U1219 (N_1219,N_841,N_654);
nand U1220 (N_1220,N_541,N_809);
or U1221 (N_1221,N_629,N_593);
and U1222 (N_1222,N_967,N_592);
nor U1223 (N_1223,N_947,N_728);
nor U1224 (N_1224,N_978,N_554);
nand U1225 (N_1225,N_706,N_617);
nand U1226 (N_1226,N_951,N_791);
xor U1227 (N_1227,N_941,N_986);
xor U1228 (N_1228,N_795,N_633);
and U1229 (N_1229,N_627,N_966);
and U1230 (N_1230,N_766,N_621);
or U1231 (N_1231,N_674,N_531);
nand U1232 (N_1232,N_610,N_879);
xor U1233 (N_1233,N_935,N_678);
nand U1234 (N_1234,N_727,N_894);
xnor U1235 (N_1235,N_540,N_954);
and U1236 (N_1236,N_799,N_903);
or U1237 (N_1237,N_907,N_547);
nand U1238 (N_1238,N_623,N_643);
or U1239 (N_1239,N_859,N_995);
nand U1240 (N_1240,N_940,N_573);
nor U1241 (N_1241,N_611,N_673);
or U1242 (N_1242,N_721,N_878);
nand U1243 (N_1243,N_591,N_717);
and U1244 (N_1244,N_893,N_882);
and U1245 (N_1245,N_836,N_737);
and U1246 (N_1246,N_849,N_518);
or U1247 (N_1247,N_936,N_871);
or U1248 (N_1248,N_539,N_534);
nor U1249 (N_1249,N_798,N_724);
and U1250 (N_1250,N_731,N_536);
nor U1251 (N_1251,N_857,N_905);
or U1252 (N_1252,N_728,N_861);
and U1253 (N_1253,N_650,N_579);
and U1254 (N_1254,N_840,N_739);
or U1255 (N_1255,N_735,N_542);
and U1256 (N_1256,N_570,N_871);
xor U1257 (N_1257,N_651,N_797);
nand U1258 (N_1258,N_782,N_779);
xor U1259 (N_1259,N_983,N_882);
xor U1260 (N_1260,N_741,N_897);
and U1261 (N_1261,N_717,N_884);
nand U1262 (N_1262,N_712,N_506);
xnor U1263 (N_1263,N_680,N_959);
xor U1264 (N_1264,N_566,N_739);
and U1265 (N_1265,N_810,N_947);
nand U1266 (N_1266,N_886,N_696);
nand U1267 (N_1267,N_925,N_878);
xor U1268 (N_1268,N_938,N_945);
nand U1269 (N_1269,N_579,N_878);
nand U1270 (N_1270,N_643,N_600);
and U1271 (N_1271,N_520,N_987);
xor U1272 (N_1272,N_510,N_531);
and U1273 (N_1273,N_718,N_884);
nand U1274 (N_1274,N_516,N_922);
nor U1275 (N_1275,N_934,N_839);
nand U1276 (N_1276,N_650,N_566);
and U1277 (N_1277,N_761,N_934);
xnor U1278 (N_1278,N_892,N_852);
or U1279 (N_1279,N_796,N_936);
nor U1280 (N_1280,N_706,N_643);
nand U1281 (N_1281,N_771,N_759);
and U1282 (N_1282,N_734,N_717);
nor U1283 (N_1283,N_558,N_768);
nand U1284 (N_1284,N_976,N_710);
xnor U1285 (N_1285,N_779,N_732);
or U1286 (N_1286,N_967,N_593);
or U1287 (N_1287,N_798,N_733);
nand U1288 (N_1288,N_674,N_880);
nand U1289 (N_1289,N_834,N_649);
or U1290 (N_1290,N_543,N_806);
nor U1291 (N_1291,N_884,N_522);
nor U1292 (N_1292,N_812,N_598);
xnor U1293 (N_1293,N_963,N_780);
or U1294 (N_1294,N_780,N_743);
nand U1295 (N_1295,N_807,N_735);
or U1296 (N_1296,N_560,N_503);
nor U1297 (N_1297,N_964,N_736);
and U1298 (N_1298,N_978,N_572);
nor U1299 (N_1299,N_505,N_895);
and U1300 (N_1300,N_622,N_669);
and U1301 (N_1301,N_896,N_912);
xor U1302 (N_1302,N_689,N_629);
nand U1303 (N_1303,N_763,N_936);
or U1304 (N_1304,N_753,N_828);
and U1305 (N_1305,N_805,N_824);
nor U1306 (N_1306,N_579,N_765);
xnor U1307 (N_1307,N_912,N_971);
nand U1308 (N_1308,N_792,N_534);
or U1309 (N_1309,N_783,N_535);
nor U1310 (N_1310,N_593,N_530);
nand U1311 (N_1311,N_942,N_701);
xnor U1312 (N_1312,N_633,N_656);
xor U1313 (N_1313,N_548,N_783);
nor U1314 (N_1314,N_934,N_624);
and U1315 (N_1315,N_819,N_880);
or U1316 (N_1316,N_772,N_921);
nor U1317 (N_1317,N_958,N_840);
nor U1318 (N_1318,N_931,N_502);
xnor U1319 (N_1319,N_856,N_768);
nand U1320 (N_1320,N_916,N_886);
or U1321 (N_1321,N_615,N_897);
and U1322 (N_1322,N_991,N_538);
or U1323 (N_1323,N_623,N_942);
or U1324 (N_1324,N_931,N_678);
nand U1325 (N_1325,N_748,N_773);
or U1326 (N_1326,N_860,N_637);
xor U1327 (N_1327,N_704,N_968);
nor U1328 (N_1328,N_602,N_581);
or U1329 (N_1329,N_664,N_681);
xor U1330 (N_1330,N_863,N_961);
nor U1331 (N_1331,N_916,N_532);
xor U1332 (N_1332,N_882,N_539);
or U1333 (N_1333,N_739,N_855);
nor U1334 (N_1334,N_967,N_872);
xnor U1335 (N_1335,N_903,N_936);
xor U1336 (N_1336,N_949,N_696);
nand U1337 (N_1337,N_698,N_764);
or U1338 (N_1338,N_684,N_547);
xnor U1339 (N_1339,N_942,N_893);
nor U1340 (N_1340,N_511,N_667);
nand U1341 (N_1341,N_801,N_516);
nor U1342 (N_1342,N_700,N_704);
xor U1343 (N_1343,N_684,N_672);
nand U1344 (N_1344,N_770,N_955);
nor U1345 (N_1345,N_896,N_709);
or U1346 (N_1346,N_981,N_949);
or U1347 (N_1347,N_787,N_912);
nor U1348 (N_1348,N_841,N_562);
or U1349 (N_1349,N_816,N_929);
or U1350 (N_1350,N_707,N_900);
xnor U1351 (N_1351,N_729,N_853);
or U1352 (N_1352,N_843,N_746);
nor U1353 (N_1353,N_880,N_670);
nand U1354 (N_1354,N_654,N_722);
xor U1355 (N_1355,N_739,N_910);
nor U1356 (N_1356,N_797,N_556);
or U1357 (N_1357,N_998,N_715);
and U1358 (N_1358,N_675,N_786);
nor U1359 (N_1359,N_772,N_507);
xor U1360 (N_1360,N_796,N_989);
and U1361 (N_1361,N_912,N_870);
nor U1362 (N_1362,N_526,N_911);
and U1363 (N_1363,N_514,N_545);
xnor U1364 (N_1364,N_501,N_920);
xor U1365 (N_1365,N_631,N_511);
nand U1366 (N_1366,N_840,N_756);
or U1367 (N_1367,N_897,N_841);
and U1368 (N_1368,N_546,N_509);
or U1369 (N_1369,N_878,N_824);
or U1370 (N_1370,N_962,N_576);
xnor U1371 (N_1371,N_733,N_616);
and U1372 (N_1372,N_636,N_633);
xor U1373 (N_1373,N_668,N_633);
or U1374 (N_1374,N_966,N_526);
or U1375 (N_1375,N_983,N_652);
and U1376 (N_1376,N_775,N_594);
nor U1377 (N_1377,N_784,N_658);
and U1378 (N_1378,N_614,N_873);
nand U1379 (N_1379,N_855,N_634);
or U1380 (N_1380,N_781,N_960);
nor U1381 (N_1381,N_646,N_724);
nand U1382 (N_1382,N_956,N_524);
nor U1383 (N_1383,N_503,N_716);
nor U1384 (N_1384,N_520,N_858);
and U1385 (N_1385,N_566,N_974);
nand U1386 (N_1386,N_507,N_817);
and U1387 (N_1387,N_607,N_577);
or U1388 (N_1388,N_504,N_824);
and U1389 (N_1389,N_847,N_999);
xnor U1390 (N_1390,N_695,N_597);
or U1391 (N_1391,N_660,N_688);
and U1392 (N_1392,N_584,N_742);
nand U1393 (N_1393,N_898,N_862);
and U1394 (N_1394,N_958,N_751);
nor U1395 (N_1395,N_920,N_711);
and U1396 (N_1396,N_725,N_562);
nor U1397 (N_1397,N_882,N_768);
and U1398 (N_1398,N_770,N_525);
xor U1399 (N_1399,N_509,N_917);
or U1400 (N_1400,N_510,N_727);
or U1401 (N_1401,N_510,N_516);
and U1402 (N_1402,N_766,N_828);
nor U1403 (N_1403,N_855,N_544);
nand U1404 (N_1404,N_678,N_860);
nand U1405 (N_1405,N_907,N_539);
nor U1406 (N_1406,N_804,N_863);
xor U1407 (N_1407,N_754,N_815);
and U1408 (N_1408,N_974,N_829);
nor U1409 (N_1409,N_928,N_587);
nor U1410 (N_1410,N_520,N_938);
and U1411 (N_1411,N_910,N_914);
nor U1412 (N_1412,N_528,N_562);
or U1413 (N_1413,N_814,N_784);
and U1414 (N_1414,N_616,N_894);
and U1415 (N_1415,N_953,N_922);
nor U1416 (N_1416,N_609,N_620);
or U1417 (N_1417,N_677,N_842);
or U1418 (N_1418,N_894,N_858);
nor U1419 (N_1419,N_647,N_984);
nor U1420 (N_1420,N_872,N_823);
xnor U1421 (N_1421,N_678,N_623);
nand U1422 (N_1422,N_730,N_814);
nor U1423 (N_1423,N_985,N_567);
or U1424 (N_1424,N_681,N_553);
nand U1425 (N_1425,N_984,N_638);
and U1426 (N_1426,N_517,N_604);
xor U1427 (N_1427,N_746,N_968);
nor U1428 (N_1428,N_579,N_859);
xor U1429 (N_1429,N_564,N_978);
nand U1430 (N_1430,N_764,N_554);
and U1431 (N_1431,N_623,N_713);
nor U1432 (N_1432,N_884,N_777);
nor U1433 (N_1433,N_694,N_865);
nand U1434 (N_1434,N_827,N_770);
and U1435 (N_1435,N_837,N_598);
nor U1436 (N_1436,N_536,N_559);
nand U1437 (N_1437,N_863,N_678);
nor U1438 (N_1438,N_509,N_652);
nor U1439 (N_1439,N_848,N_846);
or U1440 (N_1440,N_635,N_994);
nand U1441 (N_1441,N_502,N_576);
nand U1442 (N_1442,N_699,N_871);
or U1443 (N_1443,N_516,N_793);
nand U1444 (N_1444,N_744,N_746);
nand U1445 (N_1445,N_554,N_821);
and U1446 (N_1446,N_573,N_894);
nor U1447 (N_1447,N_931,N_831);
or U1448 (N_1448,N_782,N_936);
nor U1449 (N_1449,N_974,N_725);
nor U1450 (N_1450,N_986,N_683);
and U1451 (N_1451,N_653,N_652);
xor U1452 (N_1452,N_856,N_959);
or U1453 (N_1453,N_853,N_929);
or U1454 (N_1454,N_796,N_651);
xor U1455 (N_1455,N_693,N_919);
nor U1456 (N_1456,N_908,N_650);
or U1457 (N_1457,N_774,N_675);
nand U1458 (N_1458,N_599,N_546);
or U1459 (N_1459,N_929,N_926);
nor U1460 (N_1460,N_526,N_555);
and U1461 (N_1461,N_785,N_909);
or U1462 (N_1462,N_609,N_795);
nor U1463 (N_1463,N_978,N_929);
and U1464 (N_1464,N_982,N_619);
xor U1465 (N_1465,N_531,N_717);
nor U1466 (N_1466,N_914,N_698);
nand U1467 (N_1467,N_983,N_738);
or U1468 (N_1468,N_664,N_938);
and U1469 (N_1469,N_624,N_979);
or U1470 (N_1470,N_592,N_586);
nor U1471 (N_1471,N_683,N_830);
nor U1472 (N_1472,N_851,N_665);
xnor U1473 (N_1473,N_624,N_929);
or U1474 (N_1474,N_641,N_646);
and U1475 (N_1475,N_567,N_861);
xnor U1476 (N_1476,N_512,N_897);
or U1477 (N_1477,N_809,N_655);
nor U1478 (N_1478,N_573,N_549);
nand U1479 (N_1479,N_565,N_984);
and U1480 (N_1480,N_993,N_950);
nand U1481 (N_1481,N_673,N_834);
nand U1482 (N_1482,N_800,N_720);
and U1483 (N_1483,N_644,N_730);
and U1484 (N_1484,N_938,N_812);
xor U1485 (N_1485,N_601,N_999);
and U1486 (N_1486,N_794,N_932);
and U1487 (N_1487,N_509,N_576);
xnor U1488 (N_1488,N_933,N_745);
nor U1489 (N_1489,N_960,N_966);
and U1490 (N_1490,N_996,N_736);
nand U1491 (N_1491,N_888,N_900);
or U1492 (N_1492,N_739,N_761);
and U1493 (N_1493,N_691,N_741);
nand U1494 (N_1494,N_940,N_576);
nand U1495 (N_1495,N_862,N_514);
and U1496 (N_1496,N_543,N_624);
nor U1497 (N_1497,N_791,N_663);
or U1498 (N_1498,N_693,N_717);
and U1499 (N_1499,N_879,N_764);
nor U1500 (N_1500,N_1437,N_1073);
nand U1501 (N_1501,N_1328,N_1166);
or U1502 (N_1502,N_1462,N_1101);
xor U1503 (N_1503,N_1093,N_1032);
xnor U1504 (N_1504,N_1120,N_1132);
and U1505 (N_1505,N_1096,N_1390);
xor U1506 (N_1506,N_1426,N_1196);
and U1507 (N_1507,N_1237,N_1065);
nand U1508 (N_1508,N_1180,N_1001);
or U1509 (N_1509,N_1159,N_1052);
or U1510 (N_1510,N_1171,N_1023);
or U1511 (N_1511,N_1025,N_1195);
nand U1512 (N_1512,N_1402,N_1369);
xor U1513 (N_1513,N_1385,N_1264);
nand U1514 (N_1514,N_1499,N_1388);
and U1515 (N_1515,N_1313,N_1213);
xnor U1516 (N_1516,N_1004,N_1478);
nor U1517 (N_1517,N_1245,N_1394);
nand U1518 (N_1518,N_1080,N_1401);
and U1519 (N_1519,N_1044,N_1365);
nor U1520 (N_1520,N_1290,N_1179);
and U1521 (N_1521,N_1235,N_1293);
xor U1522 (N_1522,N_1410,N_1185);
and U1523 (N_1523,N_1493,N_1461);
or U1524 (N_1524,N_1027,N_1123);
xor U1525 (N_1525,N_1323,N_1434);
or U1526 (N_1526,N_1307,N_1095);
or U1527 (N_1527,N_1042,N_1090);
nor U1528 (N_1528,N_1194,N_1294);
and U1529 (N_1529,N_1189,N_1429);
nor U1530 (N_1530,N_1361,N_1452);
or U1531 (N_1531,N_1176,N_1445);
or U1532 (N_1532,N_1260,N_1136);
and U1533 (N_1533,N_1366,N_1404);
xor U1534 (N_1534,N_1269,N_1126);
or U1535 (N_1535,N_1251,N_1305);
or U1536 (N_1536,N_1480,N_1053);
nand U1537 (N_1537,N_1484,N_1270);
nor U1538 (N_1538,N_1284,N_1283);
nor U1539 (N_1539,N_1041,N_1201);
xnor U1540 (N_1540,N_1376,N_1464);
and U1541 (N_1541,N_1377,N_1068);
nand U1542 (N_1542,N_1121,N_1471);
or U1543 (N_1543,N_1038,N_1277);
xnor U1544 (N_1544,N_1491,N_1084);
nand U1545 (N_1545,N_1474,N_1497);
nor U1546 (N_1546,N_1064,N_1415);
and U1547 (N_1547,N_1314,N_1011);
nor U1548 (N_1548,N_1476,N_1382);
and U1549 (N_1549,N_1431,N_1240);
or U1550 (N_1550,N_1303,N_1048);
and U1551 (N_1551,N_1302,N_1066);
nor U1552 (N_1552,N_1133,N_1250);
or U1553 (N_1553,N_1435,N_1083);
xnor U1554 (N_1554,N_1425,N_1422);
nand U1555 (N_1555,N_1420,N_1359);
or U1556 (N_1556,N_1168,N_1383);
nand U1557 (N_1557,N_1172,N_1308);
nor U1558 (N_1558,N_1450,N_1049);
nand U1559 (N_1559,N_1267,N_1028);
and U1560 (N_1560,N_1242,N_1012);
or U1561 (N_1561,N_1490,N_1131);
and U1562 (N_1562,N_1396,N_1291);
nor U1563 (N_1563,N_1035,N_1442);
xnor U1564 (N_1564,N_1127,N_1163);
nor U1565 (N_1565,N_1333,N_1218);
and U1566 (N_1566,N_1373,N_1288);
or U1567 (N_1567,N_1386,N_1063);
xnor U1568 (N_1568,N_1204,N_1322);
nor U1569 (N_1569,N_1088,N_1424);
xnor U1570 (N_1570,N_1321,N_1263);
or U1571 (N_1571,N_1433,N_1114);
and U1572 (N_1572,N_1051,N_1329);
nor U1573 (N_1573,N_1183,N_1393);
xnor U1574 (N_1574,N_1246,N_1406);
or U1575 (N_1575,N_1444,N_1129);
xnor U1576 (N_1576,N_1432,N_1379);
nor U1577 (N_1577,N_1273,N_1258);
nor U1578 (N_1578,N_1036,N_1353);
nand U1579 (N_1579,N_1453,N_1178);
nand U1580 (N_1580,N_1468,N_1400);
and U1581 (N_1581,N_1363,N_1262);
nand U1582 (N_1582,N_1206,N_1230);
and U1583 (N_1583,N_1463,N_1152);
nor U1584 (N_1584,N_1309,N_1482);
or U1585 (N_1585,N_1078,N_1031);
nor U1586 (N_1586,N_1219,N_1224);
nand U1587 (N_1587,N_1020,N_1413);
and U1588 (N_1588,N_1352,N_1456);
and U1589 (N_1589,N_1334,N_1356);
nor U1590 (N_1590,N_1100,N_1197);
nand U1591 (N_1591,N_1207,N_1017);
nand U1592 (N_1592,N_1203,N_1466);
and U1593 (N_1593,N_1222,N_1327);
nand U1594 (N_1594,N_1370,N_1335);
nand U1595 (N_1595,N_1339,N_1254);
or U1596 (N_1596,N_1261,N_1289);
or U1597 (N_1597,N_1002,N_1311);
xor U1598 (N_1598,N_1153,N_1043);
and U1599 (N_1599,N_1330,N_1142);
xor U1600 (N_1600,N_1138,N_1029);
nand U1601 (N_1601,N_1488,N_1387);
xor U1602 (N_1602,N_1244,N_1326);
nand U1603 (N_1603,N_1010,N_1086);
or U1604 (N_1604,N_1058,N_1107);
nand U1605 (N_1605,N_1037,N_1033);
nand U1606 (N_1606,N_1380,N_1440);
nand U1607 (N_1607,N_1416,N_1475);
xor U1608 (N_1608,N_1117,N_1319);
nor U1609 (N_1609,N_1407,N_1310);
xor U1610 (N_1610,N_1439,N_1128);
and U1611 (N_1611,N_1248,N_1438);
xnor U1612 (N_1612,N_1274,N_1104);
nand U1613 (N_1613,N_1000,N_1211);
and U1614 (N_1614,N_1124,N_1423);
nor U1615 (N_1615,N_1018,N_1430);
or U1616 (N_1616,N_1072,N_1443);
nor U1617 (N_1617,N_1249,N_1479);
nand U1618 (N_1618,N_1102,N_1143);
nand U1619 (N_1619,N_1216,N_1300);
nand U1620 (N_1620,N_1292,N_1316);
xnor U1621 (N_1621,N_1351,N_1287);
and U1622 (N_1622,N_1061,N_1193);
nand U1623 (N_1623,N_1074,N_1336);
or U1624 (N_1624,N_1278,N_1364);
or U1625 (N_1625,N_1286,N_1059);
xnor U1626 (N_1626,N_1003,N_1014);
and U1627 (N_1627,N_1360,N_1485);
nand U1628 (N_1628,N_1460,N_1381);
nor U1629 (N_1629,N_1113,N_1115);
xnor U1630 (N_1630,N_1495,N_1325);
or U1631 (N_1631,N_1355,N_1349);
or U1632 (N_1632,N_1455,N_1079);
nor U1633 (N_1633,N_1296,N_1186);
nand U1634 (N_1634,N_1040,N_1141);
xor U1635 (N_1635,N_1362,N_1441);
or U1636 (N_1636,N_1275,N_1021);
xnor U1637 (N_1637,N_1492,N_1165);
nand U1638 (N_1638,N_1060,N_1105);
or U1639 (N_1639,N_1050,N_1496);
nand U1640 (N_1640,N_1076,N_1081);
or U1641 (N_1641,N_1162,N_1144);
nor U1642 (N_1642,N_1170,N_1226);
xnor U1643 (N_1643,N_1421,N_1007);
xnor U1644 (N_1644,N_1089,N_1331);
nand U1645 (N_1645,N_1232,N_1174);
nor U1646 (N_1646,N_1409,N_1215);
and U1647 (N_1647,N_1221,N_1054);
nand U1648 (N_1648,N_1139,N_1257);
and U1649 (N_1649,N_1006,N_1070);
nor U1650 (N_1650,N_1239,N_1454);
xor U1651 (N_1651,N_1408,N_1446);
nand U1652 (N_1652,N_1135,N_1469);
xnor U1653 (N_1653,N_1371,N_1259);
nor U1654 (N_1654,N_1116,N_1158);
xnor U1655 (N_1655,N_1087,N_1134);
xor U1656 (N_1656,N_1008,N_1367);
and U1657 (N_1657,N_1298,N_1137);
nand U1658 (N_1658,N_1494,N_1392);
and U1659 (N_1659,N_1071,N_1013);
nor U1660 (N_1660,N_1005,N_1299);
or U1661 (N_1661,N_1253,N_1405);
nand U1662 (N_1662,N_1487,N_1481);
nor U1663 (N_1663,N_1091,N_1057);
and U1664 (N_1664,N_1110,N_1009);
and U1665 (N_1665,N_1149,N_1338);
xor U1666 (N_1666,N_1094,N_1473);
nor U1667 (N_1667,N_1412,N_1202);
and U1668 (N_1668,N_1034,N_1119);
nand U1669 (N_1669,N_1342,N_1111);
nor U1670 (N_1670,N_1247,N_1148);
nand U1671 (N_1671,N_1103,N_1175);
nor U1672 (N_1672,N_1276,N_1085);
and U1673 (N_1673,N_1345,N_1045);
xnor U1674 (N_1674,N_1169,N_1205);
nor U1675 (N_1675,N_1428,N_1268);
xnor U1676 (N_1676,N_1055,N_1122);
and U1677 (N_1677,N_1243,N_1295);
or U1678 (N_1678,N_1324,N_1395);
and U1679 (N_1679,N_1318,N_1209);
nor U1680 (N_1680,N_1157,N_1448);
and U1681 (N_1681,N_1457,N_1200);
nand U1682 (N_1682,N_1458,N_1164);
nand U1683 (N_1683,N_1236,N_1467);
or U1684 (N_1684,N_1154,N_1252);
nor U1685 (N_1685,N_1282,N_1181);
or U1686 (N_1686,N_1372,N_1411);
and U1687 (N_1687,N_1398,N_1198);
nor U1688 (N_1688,N_1150,N_1312);
and U1689 (N_1689,N_1056,N_1419);
xor U1690 (N_1690,N_1161,N_1069);
or U1691 (N_1691,N_1403,N_1384);
and U1692 (N_1692,N_1399,N_1341);
xnor U1693 (N_1693,N_1156,N_1024);
xor U1694 (N_1694,N_1486,N_1317);
nor U1695 (N_1695,N_1229,N_1378);
xor U1696 (N_1696,N_1098,N_1470);
nor U1697 (N_1697,N_1212,N_1173);
xnor U1698 (N_1698,N_1227,N_1348);
nand U1699 (N_1699,N_1271,N_1192);
nor U1700 (N_1700,N_1146,N_1026);
or U1701 (N_1701,N_1374,N_1489);
nor U1702 (N_1702,N_1459,N_1417);
and U1703 (N_1703,N_1332,N_1280);
nand U1704 (N_1704,N_1389,N_1220);
xnor U1705 (N_1705,N_1344,N_1281);
nand U1706 (N_1706,N_1075,N_1099);
nor U1707 (N_1707,N_1155,N_1320);
nand U1708 (N_1708,N_1272,N_1483);
and U1709 (N_1709,N_1279,N_1077);
xnor U1710 (N_1710,N_1357,N_1375);
nor U1711 (N_1711,N_1062,N_1167);
xor U1712 (N_1712,N_1151,N_1285);
or U1713 (N_1713,N_1190,N_1304);
or U1714 (N_1714,N_1418,N_1414);
xor U1715 (N_1715,N_1238,N_1231);
xnor U1716 (N_1716,N_1097,N_1182);
nand U1717 (N_1717,N_1125,N_1368);
or U1718 (N_1718,N_1199,N_1145);
nand U1719 (N_1719,N_1358,N_1067);
nand U1720 (N_1720,N_1015,N_1451);
xnor U1721 (N_1721,N_1046,N_1019);
nor U1722 (N_1722,N_1177,N_1022);
and U1723 (N_1723,N_1447,N_1108);
or U1724 (N_1724,N_1147,N_1160);
or U1725 (N_1725,N_1346,N_1228);
xnor U1726 (N_1726,N_1255,N_1112);
nand U1727 (N_1727,N_1234,N_1436);
nor U1728 (N_1728,N_1350,N_1266);
or U1729 (N_1729,N_1047,N_1397);
or U1730 (N_1730,N_1477,N_1187);
xor U1731 (N_1731,N_1472,N_1109);
and U1732 (N_1732,N_1188,N_1016);
xor U1733 (N_1733,N_1039,N_1347);
xnor U1734 (N_1734,N_1210,N_1217);
xnor U1735 (N_1735,N_1106,N_1082);
or U1736 (N_1736,N_1498,N_1337);
or U1737 (N_1737,N_1449,N_1191);
and U1738 (N_1738,N_1301,N_1256);
xnor U1739 (N_1739,N_1214,N_1184);
and U1740 (N_1740,N_1306,N_1208);
nor U1741 (N_1741,N_1225,N_1092);
nand U1742 (N_1742,N_1340,N_1130);
or U1743 (N_1743,N_1297,N_1265);
nor U1744 (N_1744,N_1118,N_1223);
and U1745 (N_1745,N_1465,N_1233);
nand U1746 (N_1746,N_1354,N_1343);
nor U1747 (N_1747,N_1140,N_1241);
nor U1748 (N_1748,N_1030,N_1391);
xnor U1749 (N_1749,N_1315,N_1427);
or U1750 (N_1750,N_1234,N_1038);
xnor U1751 (N_1751,N_1004,N_1308);
and U1752 (N_1752,N_1343,N_1218);
and U1753 (N_1753,N_1283,N_1009);
and U1754 (N_1754,N_1499,N_1166);
and U1755 (N_1755,N_1143,N_1410);
and U1756 (N_1756,N_1192,N_1005);
or U1757 (N_1757,N_1169,N_1077);
and U1758 (N_1758,N_1395,N_1233);
nand U1759 (N_1759,N_1294,N_1293);
or U1760 (N_1760,N_1421,N_1445);
nand U1761 (N_1761,N_1115,N_1304);
xor U1762 (N_1762,N_1484,N_1032);
nor U1763 (N_1763,N_1407,N_1079);
and U1764 (N_1764,N_1395,N_1255);
or U1765 (N_1765,N_1354,N_1228);
or U1766 (N_1766,N_1186,N_1312);
xor U1767 (N_1767,N_1142,N_1456);
nor U1768 (N_1768,N_1089,N_1368);
nor U1769 (N_1769,N_1307,N_1014);
and U1770 (N_1770,N_1150,N_1203);
and U1771 (N_1771,N_1476,N_1335);
or U1772 (N_1772,N_1346,N_1166);
or U1773 (N_1773,N_1423,N_1472);
and U1774 (N_1774,N_1401,N_1171);
and U1775 (N_1775,N_1355,N_1378);
or U1776 (N_1776,N_1129,N_1468);
nor U1777 (N_1777,N_1256,N_1361);
nor U1778 (N_1778,N_1196,N_1471);
xnor U1779 (N_1779,N_1454,N_1410);
nand U1780 (N_1780,N_1061,N_1068);
nand U1781 (N_1781,N_1085,N_1038);
or U1782 (N_1782,N_1370,N_1338);
nor U1783 (N_1783,N_1353,N_1131);
xnor U1784 (N_1784,N_1011,N_1085);
and U1785 (N_1785,N_1340,N_1021);
nor U1786 (N_1786,N_1316,N_1235);
or U1787 (N_1787,N_1141,N_1240);
xnor U1788 (N_1788,N_1215,N_1382);
xor U1789 (N_1789,N_1319,N_1255);
nand U1790 (N_1790,N_1415,N_1233);
nor U1791 (N_1791,N_1207,N_1433);
xnor U1792 (N_1792,N_1034,N_1399);
and U1793 (N_1793,N_1457,N_1141);
or U1794 (N_1794,N_1069,N_1259);
nand U1795 (N_1795,N_1227,N_1080);
nor U1796 (N_1796,N_1235,N_1253);
nand U1797 (N_1797,N_1310,N_1031);
and U1798 (N_1798,N_1179,N_1090);
nor U1799 (N_1799,N_1001,N_1468);
or U1800 (N_1800,N_1338,N_1040);
or U1801 (N_1801,N_1284,N_1406);
or U1802 (N_1802,N_1118,N_1121);
or U1803 (N_1803,N_1029,N_1083);
nand U1804 (N_1804,N_1190,N_1049);
or U1805 (N_1805,N_1012,N_1265);
nor U1806 (N_1806,N_1162,N_1470);
nor U1807 (N_1807,N_1025,N_1473);
nor U1808 (N_1808,N_1474,N_1183);
and U1809 (N_1809,N_1197,N_1018);
xnor U1810 (N_1810,N_1070,N_1488);
nand U1811 (N_1811,N_1039,N_1047);
or U1812 (N_1812,N_1458,N_1374);
nor U1813 (N_1813,N_1082,N_1114);
and U1814 (N_1814,N_1455,N_1063);
nand U1815 (N_1815,N_1091,N_1112);
xor U1816 (N_1816,N_1391,N_1058);
and U1817 (N_1817,N_1218,N_1423);
or U1818 (N_1818,N_1390,N_1377);
and U1819 (N_1819,N_1157,N_1279);
nor U1820 (N_1820,N_1263,N_1081);
or U1821 (N_1821,N_1089,N_1241);
xnor U1822 (N_1822,N_1075,N_1484);
nand U1823 (N_1823,N_1394,N_1067);
nand U1824 (N_1824,N_1491,N_1296);
or U1825 (N_1825,N_1209,N_1004);
or U1826 (N_1826,N_1133,N_1232);
and U1827 (N_1827,N_1177,N_1351);
and U1828 (N_1828,N_1494,N_1269);
or U1829 (N_1829,N_1041,N_1181);
and U1830 (N_1830,N_1275,N_1491);
nand U1831 (N_1831,N_1212,N_1301);
nand U1832 (N_1832,N_1181,N_1130);
nor U1833 (N_1833,N_1333,N_1226);
xnor U1834 (N_1834,N_1251,N_1320);
xnor U1835 (N_1835,N_1150,N_1241);
nand U1836 (N_1836,N_1351,N_1054);
nand U1837 (N_1837,N_1419,N_1172);
nor U1838 (N_1838,N_1480,N_1313);
nor U1839 (N_1839,N_1031,N_1186);
nor U1840 (N_1840,N_1337,N_1038);
nor U1841 (N_1841,N_1061,N_1021);
nor U1842 (N_1842,N_1141,N_1038);
and U1843 (N_1843,N_1472,N_1373);
or U1844 (N_1844,N_1273,N_1475);
nand U1845 (N_1845,N_1337,N_1471);
and U1846 (N_1846,N_1327,N_1397);
and U1847 (N_1847,N_1461,N_1034);
nor U1848 (N_1848,N_1104,N_1391);
and U1849 (N_1849,N_1097,N_1433);
nor U1850 (N_1850,N_1136,N_1268);
nor U1851 (N_1851,N_1135,N_1448);
and U1852 (N_1852,N_1247,N_1423);
or U1853 (N_1853,N_1067,N_1270);
and U1854 (N_1854,N_1187,N_1133);
nor U1855 (N_1855,N_1147,N_1433);
nor U1856 (N_1856,N_1021,N_1407);
or U1857 (N_1857,N_1418,N_1313);
and U1858 (N_1858,N_1494,N_1247);
and U1859 (N_1859,N_1151,N_1100);
xor U1860 (N_1860,N_1291,N_1186);
nor U1861 (N_1861,N_1379,N_1257);
nor U1862 (N_1862,N_1071,N_1359);
nor U1863 (N_1863,N_1022,N_1081);
or U1864 (N_1864,N_1137,N_1481);
nor U1865 (N_1865,N_1419,N_1278);
or U1866 (N_1866,N_1413,N_1177);
nor U1867 (N_1867,N_1336,N_1031);
nor U1868 (N_1868,N_1497,N_1256);
nand U1869 (N_1869,N_1005,N_1032);
nor U1870 (N_1870,N_1301,N_1406);
or U1871 (N_1871,N_1473,N_1270);
xnor U1872 (N_1872,N_1406,N_1254);
and U1873 (N_1873,N_1247,N_1035);
and U1874 (N_1874,N_1311,N_1029);
and U1875 (N_1875,N_1292,N_1049);
and U1876 (N_1876,N_1138,N_1197);
and U1877 (N_1877,N_1476,N_1079);
nor U1878 (N_1878,N_1327,N_1001);
and U1879 (N_1879,N_1342,N_1166);
and U1880 (N_1880,N_1196,N_1353);
and U1881 (N_1881,N_1250,N_1126);
and U1882 (N_1882,N_1133,N_1135);
nand U1883 (N_1883,N_1366,N_1465);
xnor U1884 (N_1884,N_1264,N_1136);
xor U1885 (N_1885,N_1058,N_1244);
xnor U1886 (N_1886,N_1465,N_1192);
nand U1887 (N_1887,N_1176,N_1377);
nand U1888 (N_1888,N_1423,N_1329);
xor U1889 (N_1889,N_1143,N_1125);
xor U1890 (N_1890,N_1352,N_1054);
xnor U1891 (N_1891,N_1088,N_1394);
nor U1892 (N_1892,N_1101,N_1263);
nor U1893 (N_1893,N_1169,N_1420);
nor U1894 (N_1894,N_1116,N_1040);
and U1895 (N_1895,N_1018,N_1044);
xnor U1896 (N_1896,N_1335,N_1061);
nand U1897 (N_1897,N_1150,N_1475);
or U1898 (N_1898,N_1338,N_1023);
or U1899 (N_1899,N_1288,N_1319);
xor U1900 (N_1900,N_1443,N_1259);
nand U1901 (N_1901,N_1326,N_1298);
and U1902 (N_1902,N_1393,N_1299);
and U1903 (N_1903,N_1114,N_1061);
xnor U1904 (N_1904,N_1228,N_1291);
nor U1905 (N_1905,N_1010,N_1091);
nor U1906 (N_1906,N_1244,N_1233);
or U1907 (N_1907,N_1369,N_1230);
nor U1908 (N_1908,N_1288,N_1219);
nand U1909 (N_1909,N_1439,N_1321);
xnor U1910 (N_1910,N_1415,N_1086);
xnor U1911 (N_1911,N_1282,N_1339);
and U1912 (N_1912,N_1335,N_1398);
or U1913 (N_1913,N_1079,N_1158);
nand U1914 (N_1914,N_1283,N_1141);
nand U1915 (N_1915,N_1082,N_1237);
xor U1916 (N_1916,N_1249,N_1041);
or U1917 (N_1917,N_1353,N_1411);
xor U1918 (N_1918,N_1133,N_1347);
xnor U1919 (N_1919,N_1335,N_1365);
nand U1920 (N_1920,N_1445,N_1459);
and U1921 (N_1921,N_1372,N_1356);
and U1922 (N_1922,N_1174,N_1277);
and U1923 (N_1923,N_1407,N_1322);
nand U1924 (N_1924,N_1069,N_1020);
nand U1925 (N_1925,N_1333,N_1417);
xnor U1926 (N_1926,N_1438,N_1417);
or U1927 (N_1927,N_1478,N_1281);
nor U1928 (N_1928,N_1164,N_1330);
nor U1929 (N_1929,N_1020,N_1350);
or U1930 (N_1930,N_1067,N_1006);
or U1931 (N_1931,N_1499,N_1403);
nor U1932 (N_1932,N_1077,N_1019);
xor U1933 (N_1933,N_1090,N_1005);
and U1934 (N_1934,N_1198,N_1417);
and U1935 (N_1935,N_1102,N_1198);
nand U1936 (N_1936,N_1196,N_1448);
xor U1937 (N_1937,N_1312,N_1388);
or U1938 (N_1938,N_1201,N_1247);
nor U1939 (N_1939,N_1456,N_1464);
xnor U1940 (N_1940,N_1254,N_1115);
and U1941 (N_1941,N_1033,N_1050);
xor U1942 (N_1942,N_1356,N_1115);
nand U1943 (N_1943,N_1330,N_1450);
and U1944 (N_1944,N_1470,N_1028);
nand U1945 (N_1945,N_1217,N_1321);
or U1946 (N_1946,N_1398,N_1032);
or U1947 (N_1947,N_1142,N_1367);
and U1948 (N_1948,N_1341,N_1329);
nand U1949 (N_1949,N_1261,N_1054);
nand U1950 (N_1950,N_1150,N_1263);
nand U1951 (N_1951,N_1281,N_1122);
or U1952 (N_1952,N_1373,N_1202);
or U1953 (N_1953,N_1159,N_1025);
and U1954 (N_1954,N_1275,N_1045);
nor U1955 (N_1955,N_1270,N_1080);
or U1956 (N_1956,N_1347,N_1491);
or U1957 (N_1957,N_1343,N_1482);
or U1958 (N_1958,N_1319,N_1415);
nand U1959 (N_1959,N_1260,N_1343);
nor U1960 (N_1960,N_1180,N_1220);
xnor U1961 (N_1961,N_1138,N_1417);
nor U1962 (N_1962,N_1183,N_1020);
and U1963 (N_1963,N_1391,N_1494);
and U1964 (N_1964,N_1206,N_1393);
nand U1965 (N_1965,N_1083,N_1147);
nor U1966 (N_1966,N_1177,N_1108);
nand U1967 (N_1967,N_1304,N_1110);
and U1968 (N_1968,N_1155,N_1252);
xor U1969 (N_1969,N_1356,N_1391);
nor U1970 (N_1970,N_1268,N_1315);
nor U1971 (N_1971,N_1288,N_1374);
or U1972 (N_1972,N_1244,N_1454);
nand U1973 (N_1973,N_1026,N_1441);
xor U1974 (N_1974,N_1226,N_1100);
and U1975 (N_1975,N_1008,N_1209);
nor U1976 (N_1976,N_1375,N_1413);
nand U1977 (N_1977,N_1281,N_1114);
xor U1978 (N_1978,N_1063,N_1135);
xnor U1979 (N_1979,N_1317,N_1176);
nand U1980 (N_1980,N_1477,N_1432);
or U1981 (N_1981,N_1406,N_1438);
and U1982 (N_1982,N_1371,N_1229);
nor U1983 (N_1983,N_1214,N_1272);
or U1984 (N_1984,N_1328,N_1036);
and U1985 (N_1985,N_1129,N_1234);
nand U1986 (N_1986,N_1449,N_1275);
and U1987 (N_1987,N_1001,N_1494);
nand U1988 (N_1988,N_1148,N_1296);
nand U1989 (N_1989,N_1429,N_1049);
and U1990 (N_1990,N_1396,N_1177);
nand U1991 (N_1991,N_1056,N_1359);
and U1992 (N_1992,N_1296,N_1254);
xor U1993 (N_1993,N_1187,N_1422);
or U1994 (N_1994,N_1010,N_1258);
nand U1995 (N_1995,N_1255,N_1118);
and U1996 (N_1996,N_1149,N_1005);
nand U1997 (N_1997,N_1026,N_1271);
xnor U1998 (N_1998,N_1249,N_1049);
or U1999 (N_1999,N_1434,N_1006);
and U2000 (N_2000,N_1832,N_1942);
or U2001 (N_2001,N_1643,N_1862);
nor U2002 (N_2002,N_1994,N_1707);
nand U2003 (N_2003,N_1745,N_1959);
xor U2004 (N_2004,N_1888,N_1816);
nor U2005 (N_2005,N_1814,N_1540);
nand U2006 (N_2006,N_1833,N_1756);
or U2007 (N_2007,N_1658,N_1851);
and U2008 (N_2008,N_1843,N_1501);
xor U2009 (N_2009,N_1790,N_1515);
nand U2010 (N_2010,N_1989,N_1892);
nand U2011 (N_2011,N_1673,N_1688);
or U2012 (N_2012,N_1677,N_1736);
nor U2013 (N_2013,N_1693,N_1624);
nor U2014 (N_2014,N_1772,N_1992);
and U2015 (N_2015,N_1689,N_1977);
nand U2016 (N_2016,N_1825,N_1823);
xnor U2017 (N_2017,N_1993,N_1670);
xor U2018 (N_2018,N_1605,N_1742);
or U2019 (N_2019,N_1741,N_1676);
nand U2020 (N_2020,N_1958,N_1848);
nand U2021 (N_2021,N_1762,N_1854);
nor U2022 (N_2022,N_1530,N_1627);
or U2023 (N_2023,N_1713,N_1903);
or U2024 (N_2024,N_1894,N_1522);
nor U2025 (N_2025,N_1671,N_1821);
xor U2026 (N_2026,N_1793,N_1866);
and U2027 (N_2027,N_1682,N_1811);
xor U2028 (N_2028,N_1754,N_1509);
or U2029 (N_2029,N_1571,N_1512);
or U2030 (N_2030,N_1615,N_1808);
nor U2031 (N_2031,N_1973,N_1988);
and U2032 (N_2032,N_1621,N_1697);
xor U2033 (N_2033,N_1572,N_1828);
or U2034 (N_2034,N_1990,N_1529);
and U2035 (N_2035,N_1961,N_1696);
xnor U2036 (N_2036,N_1794,N_1776);
nor U2037 (N_2037,N_1545,N_1863);
and U2038 (N_2038,N_1698,N_1724);
nor U2039 (N_2039,N_1651,N_1806);
nor U2040 (N_2040,N_1800,N_1637);
and U2041 (N_2041,N_1907,N_1983);
and U2042 (N_2042,N_1830,N_1604);
and U2043 (N_2043,N_1887,N_1998);
nor U2044 (N_2044,N_1886,N_1779);
xnor U2045 (N_2045,N_1568,N_1967);
nand U2046 (N_2046,N_1946,N_1686);
or U2047 (N_2047,N_1955,N_1739);
and U2048 (N_2048,N_1516,N_1985);
or U2049 (N_2049,N_1553,N_1582);
and U2050 (N_2050,N_1934,N_1896);
nand U2051 (N_2051,N_1921,N_1917);
or U2052 (N_2052,N_1839,N_1660);
nor U2053 (N_2053,N_1653,N_1623);
xor U2054 (N_2054,N_1902,N_1703);
and U2055 (N_2055,N_1928,N_1730);
xnor U2056 (N_2056,N_1565,N_1581);
and U2057 (N_2057,N_1710,N_1836);
xor U2058 (N_2058,N_1687,N_1751);
nand U2059 (N_2059,N_1978,N_1858);
nand U2060 (N_2060,N_1891,N_1504);
nor U2061 (N_2061,N_1592,N_1879);
nand U2062 (N_2062,N_1838,N_1878);
xor U2063 (N_2063,N_1603,N_1655);
or U2064 (N_2064,N_1997,N_1783);
or U2065 (N_2065,N_1586,N_1564);
and U2066 (N_2066,N_1727,N_1717);
or U2067 (N_2067,N_1585,N_1949);
or U2068 (N_2068,N_1746,N_1923);
nor U2069 (N_2069,N_1780,N_1867);
nor U2070 (N_2070,N_1890,N_1555);
and U2071 (N_2071,N_1922,N_1726);
nor U2072 (N_2072,N_1781,N_1588);
and U2073 (N_2073,N_1953,N_1721);
nor U2074 (N_2074,N_1778,N_1506);
or U2075 (N_2075,N_1803,N_1812);
xor U2076 (N_2076,N_1981,N_1680);
or U2077 (N_2077,N_1583,N_1593);
nor U2078 (N_2078,N_1744,N_1749);
nand U2079 (N_2079,N_1633,N_1574);
xor U2080 (N_2080,N_1587,N_1578);
and U2081 (N_2081,N_1602,N_1943);
or U2082 (N_2082,N_1791,N_1711);
or U2083 (N_2083,N_1813,N_1523);
nor U2084 (N_2084,N_1667,N_1514);
and U2085 (N_2085,N_1700,N_1982);
or U2086 (N_2086,N_1884,N_1809);
or U2087 (N_2087,N_1659,N_1984);
xnor U2088 (N_2088,N_1834,N_1556);
nand U2089 (N_2089,N_1566,N_1526);
nor U2090 (N_2090,N_1999,N_1580);
xnor U2091 (N_2091,N_1827,N_1541);
or U2092 (N_2092,N_1718,N_1906);
nand U2093 (N_2093,N_1563,N_1964);
and U2094 (N_2094,N_1511,N_1951);
xnor U2095 (N_2095,N_1757,N_1962);
xnor U2096 (N_2096,N_1939,N_1844);
or U2097 (N_2097,N_1842,N_1738);
or U2098 (N_2098,N_1665,N_1557);
or U2099 (N_2099,N_1678,N_1770);
nor U2100 (N_2100,N_1639,N_1974);
and U2101 (N_2101,N_1775,N_1972);
xor U2102 (N_2102,N_1532,N_1976);
xor U2103 (N_2103,N_1782,N_1877);
or U2104 (N_2104,N_1647,N_1542);
nor U2105 (N_2105,N_1761,N_1785);
nor U2106 (N_2106,N_1620,N_1747);
nor U2107 (N_2107,N_1788,N_1648);
xnor U2108 (N_2108,N_1908,N_1699);
nand U2109 (N_2109,N_1692,N_1634);
xnor U2110 (N_2110,N_1929,N_1570);
nor U2111 (N_2111,N_1644,N_1801);
nand U2112 (N_2112,N_1594,N_1966);
or U2113 (N_2113,N_1763,N_1549);
or U2114 (N_2114,N_1599,N_1715);
nor U2115 (N_2115,N_1712,N_1737);
nand U2116 (N_2116,N_1933,N_1753);
and U2117 (N_2117,N_1547,N_1690);
or U2118 (N_2118,N_1940,N_1871);
xor U2119 (N_2119,N_1952,N_1614);
or U2120 (N_2120,N_1740,N_1635);
or U2121 (N_2121,N_1668,N_1610);
nand U2122 (N_2122,N_1666,N_1956);
nand U2123 (N_2123,N_1915,N_1799);
nor U2124 (N_2124,N_1840,N_1607);
xor U2125 (N_2125,N_1550,N_1706);
xnor U2126 (N_2126,N_1641,N_1861);
nand U2127 (N_2127,N_1792,N_1979);
or U2128 (N_2128,N_1817,N_1971);
xnor U2129 (N_2129,N_1649,N_1598);
nand U2130 (N_2130,N_1846,N_1748);
and U2131 (N_2131,N_1880,N_1849);
nand U2132 (N_2132,N_1657,N_1650);
xor U2133 (N_2133,N_1938,N_1960);
nand U2134 (N_2134,N_1510,N_1517);
xnor U2135 (N_2135,N_1954,N_1534);
nand U2136 (N_2136,N_1609,N_1525);
nand U2137 (N_2137,N_1968,N_1784);
and U2138 (N_2138,N_1819,N_1760);
nand U2139 (N_2139,N_1787,N_1694);
xor U2140 (N_2140,N_1732,N_1991);
nor U2141 (N_2141,N_1552,N_1656);
xnor U2142 (N_2142,N_1767,N_1619);
xor U2143 (N_2143,N_1935,N_1875);
xor U2144 (N_2144,N_1764,N_1868);
or U2145 (N_2145,N_1683,N_1654);
nor U2146 (N_2146,N_1546,N_1904);
or U2147 (N_2147,N_1898,N_1562);
nor U2148 (N_2148,N_1796,N_1963);
nand U2149 (N_2149,N_1729,N_1535);
nand U2150 (N_2150,N_1618,N_1554);
xnor U2151 (N_2151,N_1669,N_1743);
nor U2152 (N_2152,N_1629,N_1810);
nor U2153 (N_2153,N_1925,N_1558);
or U2154 (N_2154,N_1590,N_1857);
or U2155 (N_2155,N_1714,N_1543);
xnor U2156 (N_2156,N_1860,N_1987);
or U2157 (N_2157,N_1835,N_1941);
nor U2158 (N_2158,N_1705,N_1573);
nand U2159 (N_2159,N_1759,N_1895);
nand U2160 (N_2160,N_1822,N_1652);
xor U2161 (N_2161,N_1548,N_1765);
nor U2162 (N_2162,N_1521,N_1613);
or U2163 (N_2163,N_1595,N_1872);
and U2164 (N_2164,N_1897,N_1533);
and U2165 (N_2165,N_1539,N_1576);
nor U2166 (N_2166,N_1575,N_1752);
nand U2167 (N_2167,N_1559,N_1845);
nand U2168 (N_2168,N_1519,N_1750);
nand U2169 (N_2169,N_1617,N_1640);
xor U2170 (N_2170,N_1758,N_1913);
or U2171 (N_2171,N_1709,N_1926);
and U2172 (N_2172,N_1642,N_1662);
or U2173 (N_2173,N_1537,N_1569);
nand U2174 (N_2174,N_1685,N_1612);
or U2175 (N_2175,N_1975,N_1719);
nor U2176 (N_2176,N_1931,N_1970);
nand U2177 (N_2177,N_1536,N_1859);
nand U2178 (N_2178,N_1735,N_1731);
or U2179 (N_2179,N_1606,N_1734);
or U2180 (N_2180,N_1957,N_1513);
and U2181 (N_2181,N_1919,N_1538);
nor U2182 (N_2182,N_1725,N_1881);
or U2183 (N_2183,N_1824,N_1518);
xnor U2184 (N_2184,N_1560,N_1531);
or U2185 (N_2185,N_1632,N_1722);
or U2186 (N_2186,N_1625,N_1996);
nand U2187 (N_2187,N_1589,N_1950);
nor U2188 (N_2188,N_1507,N_1918);
nand U2189 (N_2189,N_1829,N_1684);
xnor U2190 (N_2190,N_1841,N_1723);
and U2191 (N_2191,N_1755,N_1505);
xnor U2192 (N_2192,N_1936,N_1969);
or U2193 (N_2193,N_1597,N_1807);
xor U2194 (N_2194,N_1932,N_1873);
or U2195 (N_2195,N_1773,N_1716);
and U2196 (N_2196,N_1870,N_1503);
nor U2197 (N_2197,N_1672,N_1630);
or U2198 (N_2198,N_1865,N_1551);
and U2199 (N_2199,N_1733,N_1986);
xor U2200 (N_2200,N_1804,N_1852);
xor U2201 (N_2201,N_1616,N_1826);
and U2202 (N_2202,N_1528,N_1622);
nor U2203 (N_2203,N_1577,N_1789);
or U2204 (N_2204,N_1820,N_1774);
and U2205 (N_2205,N_1916,N_1885);
nand U2206 (N_2206,N_1771,N_1853);
or U2207 (N_2207,N_1708,N_1695);
and U2208 (N_2208,N_1720,N_1701);
xor U2209 (N_2209,N_1837,N_1909);
or U2210 (N_2210,N_1944,N_1914);
nand U2211 (N_2211,N_1930,N_1636);
nand U2212 (N_2212,N_1646,N_1910);
nand U2213 (N_2213,N_1675,N_1945);
or U2214 (N_2214,N_1664,N_1638);
nor U2215 (N_2215,N_1769,N_1912);
and U2216 (N_2216,N_1901,N_1626);
nand U2217 (N_2217,N_1567,N_1856);
xnor U2218 (N_2218,N_1900,N_1786);
and U2219 (N_2219,N_1795,N_1608);
xnor U2220 (N_2220,N_1502,N_1527);
xor U2221 (N_2221,N_1869,N_1899);
xor U2222 (N_2222,N_1850,N_1704);
xor U2223 (N_2223,N_1797,N_1831);
xor U2224 (N_2224,N_1855,N_1584);
nand U2225 (N_2225,N_1520,N_1847);
and U2226 (N_2226,N_1691,N_1815);
xor U2227 (N_2227,N_1920,N_1777);
nand U2228 (N_2228,N_1600,N_1663);
nor U2229 (N_2229,N_1874,N_1728);
xor U2230 (N_2230,N_1524,N_1702);
and U2231 (N_2231,N_1679,N_1661);
xnor U2232 (N_2232,N_1611,N_1674);
nor U2233 (N_2233,N_1805,N_1995);
xor U2234 (N_2234,N_1561,N_1927);
nor U2235 (N_2235,N_1508,N_1591);
xor U2236 (N_2236,N_1905,N_1628);
and U2237 (N_2237,N_1911,N_1876);
or U2238 (N_2238,N_1948,N_1883);
xnor U2239 (N_2239,N_1864,N_1882);
xor U2240 (N_2240,N_1544,N_1766);
nand U2241 (N_2241,N_1768,N_1596);
and U2242 (N_2242,N_1937,N_1798);
and U2243 (N_2243,N_1802,N_1645);
xor U2244 (N_2244,N_1601,N_1579);
nor U2245 (N_2245,N_1500,N_1924);
xnor U2246 (N_2246,N_1980,N_1889);
nor U2247 (N_2247,N_1681,N_1631);
xnor U2248 (N_2248,N_1965,N_1947);
nand U2249 (N_2249,N_1818,N_1893);
nor U2250 (N_2250,N_1925,N_1639);
and U2251 (N_2251,N_1856,N_1564);
or U2252 (N_2252,N_1622,N_1637);
nor U2253 (N_2253,N_1566,N_1530);
nand U2254 (N_2254,N_1726,N_1927);
and U2255 (N_2255,N_1944,N_1852);
or U2256 (N_2256,N_1671,N_1717);
xor U2257 (N_2257,N_1636,N_1773);
nand U2258 (N_2258,N_1954,N_1938);
xor U2259 (N_2259,N_1547,N_1916);
and U2260 (N_2260,N_1667,N_1574);
nand U2261 (N_2261,N_1916,N_1682);
nand U2262 (N_2262,N_1850,N_1697);
nand U2263 (N_2263,N_1774,N_1586);
nand U2264 (N_2264,N_1628,N_1911);
nand U2265 (N_2265,N_1841,N_1743);
nor U2266 (N_2266,N_1511,N_1837);
and U2267 (N_2267,N_1595,N_1545);
nor U2268 (N_2268,N_1780,N_1826);
or U2269 (N_2269,N_1757,N_1854);
xnor U2270 (N_2270,N_1878,N_1931);
nand U2271 (N_2271,N_1744,N_1669);
or U2272 (N_2272,N_1557,N_1632);
nand U2273 (N_2273,N_1810,N_1625);
and U2274 (N_2274,N_1842,N_1947);
nor U2275 (N_2275,N_1641,N_1713);
nor U2276 (N_2276,N_1552,N_1505);
xor U2277 (N_2277,N_1791,N_1889);
and U2278 (N_2278,N_1771,N_1868);
nor U2279 (N_2279,N_1761,N_1845);
nand U2280 (N_2280,N_1887,N_1791);
xnor U2281 (N_2281,N_1882,N_1584);
or U2282 (N_2282,N_1863,N_1668);
xnor U2283 (N_2283,N_1921,N_1731);
and U2284 (N_2284,N_1941,N_1821);
nand U2285 (N_2285,N_1890,N_1833);
nand U2286 (N_2286,N_1641,N_1523);
xor U2287 (N_2287,N_1626,N_1573);
or U2288 (N_2288,N_1799,N_1566);
and U2289 (N_2289,N_1703,N_1997);
xor U2290 (N_2290,N_1973,N_1698);
nor U2291 (N_2291,N_1570,N_1637);
nor U2292 (N_2292,N_1683,N_1639);
and U2293 (N_2293,N_1587,N_1521);
nor U2294 (N_2294,N_1676,N_1977);
and U2295 (N_2295,N_1874,N_1625);
or U2296 (N_2296,N_1627,N_1616);
and U2297 (N_2297,N_1593,N_1904);
and U2298 (N_2298,N_1810,N_1905);
nor U2299 (N_2299,N_1699,N_1930);
xnor U2300 (N_2300,N_1936,N_1721);
nor U2301 (N_2301,N_1700,N_1608);
and U2302 (N_2302,N_1878,N_1952);
or U2303 (N_2303,N_1664,N_1703);
nor U2304 (N_2304,N_1696,N_1957);
nor U2305 (N_2305,N_1837,N_1757);
xor U2306 (N_2306,N_1639,N_1843);
nand U2307 (N_2307,N_1769,N_1768);
xor U2308 (N_2308,N_1839,N_1856);
nand U2309 (N_2309,N_1772,N_1783);
xnor U2310 (N_2310,N_1630,N_1775);
or U2311 (N_2311,N_1612,N_1872);
nand U2312 (N_2312,N_1694,N_1804);
and U2313 (N_2313,N_1504,N_1519);
nor U2314 (N_2314,N_1761,N_1689);
or U2315 (N_2315,N_1797,N_1537);
xor U2316 (N_2316,N_1594,N_1890);
xnor U2317 (N_2317,N_1821,N_1733);
or U2318 (N_2318,N_1824,N_1670);
and U2319 (N_2319,N_1643,N_1954);
and U2320 (N_2320,N_1752,N_1527);
nor U2321 (N_2321,N_1926,N_1901);
nand U2322 (N_2322,N_1992,N_1754);
nor U2323 (N_2323,N_1559,N_1699);
and U2324 (N_2324,N_1697,N_1712);
or U2325 (N_2325,N_1517,N_1930);
and U2326 (N_2326,N_1879,N_1958);
and U2327 (N_2327,N_1930,N_1842);
nand U2328 (N_2328,N_1768,N_1594);
xor U2329 (N_2329,N_1702,N_1986);
xnor U2330 (N_2330,N_1657,N_1861);
or U2331 (N_2331,N_1715,N_1923);
and U2332 (N_2332,N_1910,N_1786);
xor U2333 (N_2333,N_1916,N_1929);
nand U2334 (N_2334,N_1634,N_1600);
xnor U2335 (N_2335,N_1571,N_1513);
or U2336 (N_2336,N_1899,N_1901);
nand U2337 (N_2337,N_1654,N_1671);
and U2338 (N_2338,N_1830,N_1954);
or U2339 (N_2339,N_1970,N_1536);
xnor U2340 (N_2340,N_1512,N_1726);
and U2341 (N_2341,N_1603,N_1556);
or U2342 (N_2342,N_1778,N_1566);
and U2343 (N_2343,N_1976,N_1551);
or U2344 (N_2344,N_1853,N_1558);
or U2345 (N_2345,N_1904,N_1863);
or U2346 (N_2346,N_1825,N_1899);
nor U2347 (N_2347,N_1565,N_1861);
nand U2348 (N_2348,N_1605,N_1801);
and U2349 (N_2349,N_1563,N_1818);
and U2350 (N_2350,N_1984,N_1609);
nand U2351 (N_2351,N_1776,N_1823);
nand U2352 (N_2352,N_1877,N_1898);
nand U2353 (N_2353,N_1840,N_1784);
and U2354 (N_2354,N_1647,N_1723);
xor U2355 (N_2355,N_1543,N_1604);
nand U2356 (N_2356,N_1621,N_1663);
and U2357 (N_2357,N_1848,N_1908);
and U2358 (N_2358,N_1833,N_1640);
xor U2359 (N_2359,N_1644,N_1785);
nor U2360 (N_2360,N_1503,N_1782);
and U2361 (N_2361,N_1830,N_1514);
or U2362 (N_2362,N_1789,N_1754);
nand U2363 (N_2363,N_1853,N_1549);
xnor U2364 (N_2364,N_1827,N_1797);
or U2365 (N_2365,N_1509,N_1915);
or U2366 (N_2366,N_1907,N_1883);
nand U2367 (N_2367,N_1788,N_1721);
and U2368 (N_2368,N_1994,N_1951);
or U2369 (N_2369,N_1759,N_1683);
nand U2370 (N_2370,N_1765,N_1777);
nand U2371 (N_2371,N_1692,N_1597);
and U2372 (N_2372,N_1704,N_1530);
and U2373 (N_2373,N_1901,N_1830);
nand U2374 (N_2374,N_1897,N_1940);
or U2375 (N_2375,N_1868,N_1557);
or U2376 (N_2376,N_1665,N_1800);
or U2377 (N_2377,N_1652,N_1747);
nor U2378 (N_2378,N_1736,N_1503);
or U2379 (N_2379,N_1748,N_1679);
and U2380 (N_2380,N_1878,N_1724);
nand U2381 (N_2381,N_1659,N_1885);
nand U2382 (N_2382,N_1536,N_1640);
nor U2383 (N_2383,N_1673,N_1834);
nor U2384 (N_2384,N_1523,N_1898);
nor U2385 (N_2385,N_1603,N_1682);
and U2386 (N_2386,N_1876,N_1916);
and U2387 (N_2387,N_1857,N_1699);
and U2388 (N_2388,N_1955,N_1764);
nand U2389 (N_2389,N_1547,N_1824);
or U2390 (N_2390,N_1572,N_1647);
or U2391 (N_2391,N_1668,N_1532);
nor U2392 (N_2392,N_1643,N_1911);
xor U2393 (N_2393,N_1513,N_1601);
and U2394 (N_2394,N_1729,N_1611);
and U2395 (N_2395,N_1631,N_1740);
nand U2396 (N_2396,N_1797,N_1564);
xnor U2397 (N_2397,N_1534,N_1662);
and U2398 (N_2398,N_1610,N_1867);
or U2399 (N_2399,N_1654,N_1979);
xnor U2400 (N_2400,N_1675,N_1565);
nor U2401 (N_2401,N_1790,N_1947);
nor U2402 (N_2402,N_1929,N_1707);
or U2403 (N_2403,N_1559,N_1533);
nor U2404 (N_2404,N_1503,N_1569);
xor U2405 (N_2405,N_1733,N_1550);
nor U2406 (N_2406,N_1610,N_1805);
nor U2407 (N_2407,N_1871,N_1651);
or U2408 (N_2408,N_1936,N_1548);
nand U2409 (N_2409,N_1989,N_1965);
nor U2410 (N_2410,N_1719,N_1805);
and U2411 (N_2411,N_1921,N_1636);
nor U2412 (N_2412,N_1823,N_1643);
nor U2413 (N_2413,N_1719,N_1832);
nor U2414 (N_2414,N_1555,N_1625);
nor U2415 (N_2415,N_1967,N_1676);
or U2416 (N_2416,N_1791,N_1835);
nor U2417 (N_2417,N_1583,N_1500);
nand U2418 (N_2418,N_1871,N_1729);
or U2419 (N_2419,N_1713,N_1756);
nand U2420 (N_2420,N_1592,N_1722);
and U2421 (N_2421,N_1748,N_1675);
nand U2422 (N_2422,N_1869,N_1916);
nor U2423 (N_2423,N_1592,N_1560);
and U2424 (N_2424,N_1928,N_1843);
nand U2425 (N_2425,N_1828,N_1610);
or U2426 (N_2426,N_1577,N_1859);
and U2427 (N_2427,N_1541,N_1675);
nor U2428 (N_2428,N_1758,N_1668);
xor U2429 (N_2429,N_1571,N_1818);
or U2430 (N_2430,N_1588,N_1563);
or U2431 (N_2431,N_1937,N_1689);
nand U2432 (N_2432,N_1894,N_1694);
or U2433 (N_2433,N_1672,N_1745);
nor U2434 (N_2434,N_1837,N_1945);
and U2435 (N_2435,N_1828,N_1889);
or U2436 (N_2436,N_1776,N_1878);
or U2437 (N_2437,N_1991,N_1931);
or U2438 (N_2438,N_1854,N_1964);
nor U2439 (N_2439,N_1923,N_1861);
xor U2440 (N_2440,N_1888,N_1680);
and U2441 (N_2441,N_1982,N_1625);
xnor U2442 (N_2442,N_1870,N_1628);
or U2443 (N_2443,N_1743,N_1625);
and U2444 (N_2444,N_1657,N_1773);
xor U2445 (N_2445,N_1710,N_1957);
nor U2446 (N_2446,N_1837,N_1500);
xnor U2447 (N_2447,N_1786,N_1854);
or U2448 (N_2448,N_1834,N_1735);
and U2449 (N_2449,N_1550,N_1731);
xnor U2450 (N_2450,N_1875,N_1763);
or U2451 (N_2451,N_1658,N_1687);
nor U2452 (N_2452,N_1808,N_1865);
nand U2453 (N_2453,N_1819,N_1944);
xor U2454 (N_2454,N_1838,N_1929);
nor U2455 (N_2455,N_1799,N_1643);
xor U2456 (N_2456,N_1672,N_1517);
nand U2457 (N_2457,N_1941,N_1932);
and U2458 (N_2458,N_1727,N_1594);
nand U2459 (N_2459,N_1862,N_1821);
xor U2460 (N_2460,N_1919,N_1639);
or U2461 (N_2461,N_1869,N_1561);
and U2462 (N_2462,N_1616,N_1927);
nand U2463 (N_2463,N_1602,N_1976);
xnor U2464 (N_2464,N_1808,N_1896);
and U2465 (N_2465,N_1677,N_1975);
or U2466 (N_2466,N_1521,N_1731);
or U2467 (N_2467,N_1900,N_1635);
nor U2468 (N_2468,N_1532,N_1704);
and U2469 (N_2469,N_1572,N_1963);
nor U2470 (N_2470,N_1824,N_1938);
nand U2471 (N_2471,N_1917,N_1625);
xor U2472 (N_2472,N_1676,N_1770);
nor U2473 (N_2473,N_1991,N_1995);
or U2474 (N_2474,N_1737,N_1840);
or U2475 (N_2475,N_1861,N_1579);
nor U2476 (N_2476,N_1894,N_1506);
nor U2477 (N_2477,N_1552,N_1731);
nand U2478 (N_2478,N_1642,N_1961);
xor U2479 (N_2479,N_1577,N_1642);
nand U2480 (N_2480,N_1802,N_1556);
and U2481 (N_2481,N_1904,N_1525);
xnor U2482 (N_2482,N_1823,N_1672);
nor U2483 (N_2483,N_1524,N_1802);
and U2484 (N_2484,N_1736,N_1628);
nand U2485 (N_2485,N_1997,N_1934);
and U2486 (N_2486,N_1914,N_1545);
xnor U2487 (N_2487,N_1755,N_1918);
xnor U2488 (N_2488,N_1893,N_1623);
nor U2489 (N_2489,N_1982,N_1927);
xor U2490 (N_2490,N_1620,N_1881);
or U2491 (N_2491,N_1824,N_1975);
and U2492 (N_2492,N_1578,N_1996);
xor U2493 (N_2493,N_1934,N_1736);
nor U2494 (N_2494,N_1557,N_1654);
nand U2495 (N_2495,N_1881,N_1961);
xor U2496 (N_2496,N_1881,N_1717);
or U2497 (N_2497,N_1570,N_1872);
xnor U2498 (N_2498,N_1672,N_1737);
nand U2499 (N_2499,N_1730,N_1884);
nor U2500 (N_2500,N_2376,N_2401);
nand U2501 (N_2501,N_2373,N_2490);
nand U2502 (N_2502,N_2218,N_2379);
and U2503 (N_2503,N_2112,N_2035);
or U2504 (N_2504,N_2247,N_2458);
xnor U2505 (N_2505,N_2446,N_2282);
nor U2506 (N_2506,N_2382,N_2414);
nor U2507 (N_2507,N_2014,N_2452);
or U2508 (N_2508,N_2354,N_2496);
nand U2509 (N_2509,N_2450,N_2211);
nor U2510 (N_2510,N_2063,N_2200);
nor U2511 (N_2511,N_2321,N_2111);
or U2512 (N_2512,N_2428,N_2342);
and U2513 (N_2513,N_2015,N_2089);
nor U2514 (N_2514,N_2029,N_2206);
xor U2515 (N_2515,N_2148,N_2327);
and U2516 (N_2516,N_2067,N_2236);
nor U2517 (N_2517,N_2136,N_2171);
or U2518 (N_2518,N_2389,N_2030);
or U2519 (N_2519,N_2051,N_2073);
and U2520 (N_2520,N_2176,N_2351);
xnor U2521 (N_2521,N_2037,N_2469);
nor U2522 (N_2522,N_2040,N_2476);
or U2523 (N_2523,N_2170,N_2495);
or U2524 (N_2524,N_2307,N_2092);
nor U2525 (N_2525,N_2058,N_2241);
or U2526 (N_2526,N_2483,N_2437);
nor U2527 (N_2527,N_2477,N_2021);
or U2528 (N_2528,N_2315,N_2185);
nor U2529 (N_2529,N_2480,N_2479);
and U2530 (N_2530,N_2138,N_2086);
nor U2531 (N_2531,N_2120,N_2059);
nand U2532 (N_2532,N_2337,N_2292);
nor U2533 (N_2533,N_2155,N_2362);
or U2534 (N_2534,N_2046,N_2130);
nand U2535 (N_2535,N_2064,N_2262);
nand U2536 (N_2536,N_2287,N_2277);
nand U2537 (N_2537,N_2183,N_2137);
and U2538 (N_2538,N_2203,N_2334);
nor U2539 (N_2539,N_2234,N_2028);
and U2540 (N_2540,N_2426,N_2209);
and U2541 (N_2541,N_2072,N_2325);
xnor U2542 (N_2542,N_2433,N_2018);
nor U2543 (N_2543,N_2365,N_2377);
nor U2544 (N_2544,N_2177,N_2027);
and U2545 (N_2545,N_2164,N_2444);
xnor U2546 (N_2546,N_2356,N_2473);
nor U2547 (N_2547,N_2381,N_2098);
nor U2548 (N_2548,N_2181,N_2126);
nand U2549 (N_2549,N_2332,N_2099);
and U2550 (N_2550,N_2095,N_2424);
nor U2551 (N_2551,N_2188,N_2363);
nor U2552 (N_2552,N_2047,N_2187);
and U2553 (N_2553,N_2397,N_2281);
nand U2554 (N_2554,N_2215,N_2494);
and U2555 (N_2555,N_2470,N_2115);
nand U2556 (N_2556,N_2201,N_2260);
nand U2557 (N_2557,N_2278,N_2109);
xnor U2558 (N_2558,N_2113,N_2061);
or U2559 (N_2559,N_2129,N_2145);
and U2560 (N_2560,N_2198,N_2172);
nor U2561 (N_2561,N_2141,N_2492);
or U2562 (N_2562,N_2335,N_2229);
or U2563 (N_2563,N_2383,N_2256);
and U2564 (N_2564,N_2418,N_2268);
nand U2565 (N_2565,N_2220,N_2313);
xnor U2566 (N_2566,N_2182,N_2107);
xnor U2567 (N_2567,N_2340,N_2317);
xor U2568 (N_2568,N_2068,N_2008);
or U2569 (N_2569,N_2165,N_2336);
nor U2570 (N_2570,N_2116,N_2415);
xor U2571 (N_2571,N_2269,N_2294);
xnor U2572 (N_2572,N_2216,N_2104);
xnor U2573 (N_2573,N_2425,N_2349);
and U2574 (N_2574,N_2387,N_2066);
or U2575 (N_2575,N_2189,N_2244);
nand U2576 (N_2576,N_2467,N_2261);
xnor U2577 (N_2577,N_2108,N_2497);
nand U2578 (N_2578,N_2297,N_2443);
nor U2579 (N_2579,N_2195,N_2346);
xnor U2580 (N_2580,N_2253,N_2360);
and U2581 (N_2581,N_2402,N_2166);
nor U2582 (N_2582,N_2284,N_2408);
and U2583 (N_2583,N_2259,N_2150);
nor U2584 (N_2584,N_2295,N_2273);
and U2585 (N_2585,N_2135,N_2392);
nor U2586 (N_2586,N_2318,N_2413);
nand U2587 (N_2587,N_2090,N_2006);
nand U2588 (N_2588,N_2167,N_2353);
nor U2589 (N_2589,N_2175,N_2239);
and U2590 (N_2590,N_2065,N_2097);
nand U2591 (N_2591,N_2235,N_2403);
nand U2592 (N_2592,N_2289,N_2328);
or U2593 (N_2593,N_2157,N_2255);
nand U2594 (N_2594,N_2053,N_2398);
or U2595 (N_2595,N_2440,N_2404);
and U2596 (N_2596,N_2173,N_2184);
nand U2597 (N_2597,N_2412,N_2326);
xnor U2598 (N_2598,N_2079,N_2096);
nand U2599 (N_2599,N_2482,N_2314);
and U2600 (N_2600,N_2478,N_2463);
nand U2601 (N_2601,N_2462,N_2248);
nor U2602 (N_2602,N_2055,N_2430);
and U2603 (N_2603,N_2464,N_2405);
xor U2604 (N_2604,N_2355,N_2219);
nor U2605 (N_2605,N_2118,N_2227);
and U2606 (N_2606,N_2084,N_2213);
or U2607 (N_2607,N_2320,N_2266);
xnor U2608 (N_2608,N_2400,N_2013);
nand U2609 (N_2609,N_2385,N_2132);
xnor U2610 (N_2610,N_2019,N_2105);
nand U2611 (N_2611,N_2125,N_2017);
nand U2612 (N_2612,N_2484,N_2069);
or U2613 (N_2613,N_2323,N_2222);
xnor U2614 (N_2614,N_2384,N_2368);
nand U2615 (N_2615,N_2214,N_2386);
or U2616 (N_2616,N_2243,N_2488);
and U2617 (N_2617,N_2279,N_2455);
nor U2618 (N_2618,N_2267,N_2094);
xor U2619 (N_2619,N_2204,N_2232);
nand U2620 (N_2620,N_2251,N_2350);
xnor U2621 (N_2621,N_2309,N_2436);
nand U2622 (N_2622,N_2038,N_2169);
nor U2623 (N_2623,N_2160,N_2357);
nand U2624 (N_2624,N_2308,N_2449);
nor U2625 (N_2625,N_2103,N_2192);
or U2626 (N_2626,N_2264,N_2190);
nand U2627 (N_2627,N_2205,N_2472);
xnor U2628 (N_2628,N_2471,N_2186);
xor U2629 (N_2629,N_2466,N_2147);
xor U2630 (N_2630,N_2311,N_2212);
xnor U2631 (N_2631,N_2146,N_2022);
nor U2632 (N_2632,N_2310,N_2304);
nand U2633 (N_2633,N_2475,N_2034);
and U2634 (N_2634,N_2396,N_2366);
xnor U2635 (N_2635,N_2423,N_2272);
and U2636 (N_2636,N_2249,N_2343);
nor U2637 (N_2637,N_2143,N_2399);
xor U2638 (N_2638,N_2486,N_2161);
nor U2639 (N_2639,N_2372,N_2179);
and U2640 (N_2640,N_2296,N_2339);
and U2641 (N_2641,N_2207,N_2240);
nand U2642 (N_2642,N_2001,N_2331);
and U2643 (N_2643,N_2049,N_2411);
xnor U2644 (N_2644,N_2316,N_2276);
nor U2645 (N_2645,N_2417,N_2230);
xor U2646 (N_2646,N_2039,N_2454);
nand U2647 (N_2647,N_2265,N_2071);
nand U2648 (N_2648,N_2238,N_2100);
or U2649 (N_2649,N_2481,N_2416);
nor U2650 (N_2650,N_2083,N_2299);
nand U2651 (N_2651,N_2274,N_2300);
and U2652 (N_2652,N_2062,N_2052);
nor U2653 (N_2653,N_2395,N_2431);
nor U2654 (N_2654,N_2298,N_2461);
nand U2655 (N_2655,N_2361,N_2093);
xnor U2656 (N_2656,N_2081,N_2144);
nor U2657 (N_2657,N_2162,N_2142);
or U2658 (N_2658,N_2033,N_2110);
xnor U2659 (N_2659,N_2114,N_2054);
nand U2660 (N_2660,N_2131,N_2448);
or U2661 (N_2661,N_2283,N_2427);
or U2662 (N_2662,N_2223,N_2288);
or U2663 (N_2663,N_2441,N_2158);
or U2664 (N_2664,N_2102,N_2286);
nand U2665 (N_2665,N_2026,N_2487);
xnor U2666 (N_2666,N_2004,N_2237);
nor U2667 (N_2667,N_2371,N_2333);
xnor U2668 (N_2668,N_2010,N_2154);
nor U2669 (N_2669,N_2250,N_2152);
nor U2670 (N_2670,N_2036,N_2041);
and U2671 (N_2671,N_2406,N_2293);
xnor U2672 (N_2672,N_2388,N_2194);
and U2673 (N_2673,N_2302,N_2045);
and U2674 (N_2674,N_2139,N_2375);
nor U2675 (N_2675,N_2499,N_2390);
or U2676 (N_2676,N_2270,N_2048);
nor U2677 (N_2677,N_2348,N_2078);
xor U2678 (N_2678,N_2319,N_2465);
nor U2679 (N_2679,N_2149,N_2391);
nor U2680 (N_2680,N_2134,N_2074);
or U2681 (N_2681,N_2280,N_2101);
or U2682 (N_2682,N_2271,N_2208);
xnor U2683 (N_2683,N_2445,N_2031);
or U2684 (N_2684,N_2221,N_2493);
and U2685 (N_2685,N_2224,N_2023);
and U2686 (N_2686,N_2303,N_2060);
and U2687 (N_2687,N_2202,N_2491);
nor U2688 (N_2688,N_2329,N_2106);
nor U2689 (N_2689,N_2070,N_2024);
and U2690 (N_2690,N_2210,N_2453);
xnor U2691 (N_2691,N_2245,N_2057);
and U2692 (N_2692,N_2410,N_2422);
xor U2693 (N_2693,N_2257,N_2254);
and U2694 (N_2694,N_2447,N_2291);
xnor U2695 (N_2695,N_2011,N_2085);
or U2696 (N_2696,N_2258,N_2474);
nor U2697 (N_2697,N_2124,N_2352);
or U2698 (N_2698,N_2393,N_2380);
nand U2699 (N_2699,N_2228,N_2364);
xor U2700 (N_2700,N_2242,N_2407);
xor U2701 (N_2701,N_2438,N_2312);
and U2702 (N_2702,N_2044,N_2080);
xor U2703 (N_2703,N_2128,N_2002);
and U2704 (N_2704,N_2442,N_2020);
xnor U2705 (N_2705,N_2088,N_2468);
nand U2706 (N_2706,N_2370,N_2077);
or U2707 (N_2707,N_2153,N_2435);
nand U2708 (N_2708,N_2330,N_2075);
and U2709 (N_2709,N_2421,N_2459);
nand U2710 (N_2710,N_2032,N_2003);
nor U2711 (N_2711,N_2180,N_2123);
or U2712 (N_2712,N_2217,N_2140);
or U2713 (N_2713,N_2025,N_2306);
nand U2714 (N_2714,N_2485,N_2199);
xnor U2715 (N_2715,N_2009,N_2082);
nor U2716 (N_2716,N_2344,N_2087);
or U2717 (N_2717,N_2358,N_2275);
xnor U2718 (N_2718,N_2451,N_2174);
xnor U2719 (N_2719,N_2056,N_2434);
or U2720 (N_2720,N_2341,N_2050);
or U2721 (N_2721,N_2409,N_2498);
or U2722 (N_2722,N_2133,N_2305);
nand U2723 (N_2723,N_2012,N_2117);
xor U2724 (N_2724,N_2439,N_2000);
or U2725 (N_2725,N_2159,N_2196);
nand U2726 (N_2726,N_2043,N_2007);
and U2727 (N_2727,N_2460,N_2121);
nor U2728 (N_2728,N_2178,N_2419);
and U2729 (N_2729,N_2225,N_2091);
and U2730 (N_2730,N_2394,N_2322);
or U2731 (N_2731,N_2191,N_2016);
nor U2732 (N_2732,N_2163,N_2119);
nor U2733 (N_2733,N_2156,N_2429);
nand U2734 (N_2734,N_2226,N_2168);
nor U2735 (N_2735,N_2324,N_2263);
nand U2736 (N_2736,N_2290,N_2369);
nor U2737 (N_2737,N_2246,N_2122);
xnor U2738 (N_2738,N_2151,N_2076);
or U2739 (N_2739,N_2489,N_2359);
nor U2740 (N_2740,N_2420,N_2285);
and U2741 (N_2741,N_2378,N_2345);
nor U2742 (N_2742,N_2367,N_2231);
and U2743 (N_2743,N_2347,N_2252);
nor U2744 (N_2744,N_2042,N_2005);
nand U2745 (N_2745,N_2456,N_2432);
and U2746 (N_2746,N_2338,N_2127);
or U2747 (N_2747,N_2233,N_2193);
nor U2748 (N_2748,N_2197,N_2301);
or U2749 (N_2749,N_2374,N_2457);
or U2750 (N_2750,N_2009,N_2309);
or U2751 (N_2751,N_2448,N_2066);
nor U2752 (N_2752,N_2315,N_2074);
xor U2753 (N_2753,N_2216,N_2375);
and U2754 (N_2754,N_2169,N_2056);
xor U2755 (N_2755,N_2495,N_2173);
nor U2756 (N_2756,N_2037,N_2081);
nand U2757 (N_2757,N_2151,N_2056);
nor U2758 (N_2758,N_2060,N_2470);
xnor U2759 (N_2759,N_2328,N_2142);
xor U2760 (N_2760,N_2335,N_2205);
xnor U2761 (N_2761,N_2120,N_2058);
nand U2762 (N_2762,N_2208,N_2450);
nor U2763 (N_2763,N_2426,N_2482);
or U2764 (N_2764,N_2376,N_2331);
nand U2765 (N_2765,N_2253,N_2424);
or U2766 (N_2766,N_2344,N_2112);
or U2767 (N_2767,N_2236,N_2106);
xor U2768 (N_2768,N_2302,N_2021);
nor U2769 (N_2769,N_2433,N_2195);
or U2770 (N_2770,N_2223,N_2264);
or U2771 (N_2771,N_2310,N_2461);
and U2772 (N_2772,N_2006,N_2436);
nor U2773 (N_2773,N_2138,N_2220);
xor U2774 (N_2774,N_2052,N_2094);
and U2775 (N_2775,N_2019,N_2456);
xnor U2776 (N_2776,N_2138,N_2178);
xnor U2777 (N_2777,N_2065,N_2165);
nand U2778 (N_2778,N_2283,N_2314);
and U2779 (N_2779,N_2396,N_2223);
and U2780 (N_2780,N_2182,N_2350);
nor U2781 (N_2781,N_2213,N_2140);
or U2782 (N_2782,N_2287,N_2477);
and U2783 (N_2783,N_2059,N_2210);
nand U2784 (N_2784,N_2170,N_2254);
or U2785 (N_2785,N_2298,N_2104);
nand U2786 (N_2786,N_2383,N_2419);
xnor U2787 (N_2787,N_2395,N_2422);
nand U2788 (N_2788,N_2353,N_2026);
nor U2789 (N_2789,N_2350,N_2275);
nand U2790 (N_2790,N_2265,N_2417);
and U2791 (N_2791,N_2291,N_2063);
or U2792 (N_2792,N_2057,N_2032);
and U2793 (N_2793,N_2168,N_2265);
xnor U2794 (N_2794,N_2309,N_2204);
and U2795 (N_2795,N_2167,N_2387);
nor U2796 (N_2796,N_2240,N_2308);
nor U2797 (N_2797,N_2174,N_2017);
nor U2798 (N_2798,N_2273,N_2388);
nor U2799 (N_2799,N_2373,N_2464);
nand U2800 (N_2800,N_2098,N_2389);
nand U2801 (N_2801,N_2158,N_2382);
and U2802 (N_2802,N_2497,N_2215);
and U2803 (N_2803,N_2046,N_2188);
or U2804 (N_2804,N_2449,N_2141);
or U2805 (N_2805,N_2152,N_2409);
xnor U2806 (N_2806,N_2048,N_2483);
nand U2807 (N_2807,N_2160,N_2106);
and U2808 (N_2808,N_2286,N_2012);
or U2809 (N_2809,N_2457,N_2334);
and U2810 (N_2810,N_2441,N_2014);
and U2811 (N_2811,N_2444,N_2397);
or U2812 (N_2812,N_2168,N_2072);
nand U2813 (N_2813,N_2231,N_2149);
xor U2814 (N_2814,N_2254,N_2043);
nor U2815 (N_2815,N_2061,N_2063);
xnor U2816 (N_2816,N_2065,N_2213);
nand U2817 (N_2817,N_2196,N_2389);
or U2818 (N_2818,N_2047,N_2057);
nor U2819 (N_2819,N_2405,N_2100);
nand U2820 (N_2820,N_2339,N_2107);
nand U2821 (N_2821,N_2089,N_2459);
and U2822 (N_2822,N_2153,N_2091);
nor U2823 (N_2823,N_2028,N_2494);
and U2824 (N_2824,N_2357,N_2323);
xnor U2825 (N_2825,N_2146,N_2013);
nor U2826 (N_2826,N_2388,N_2268);
nor U2827 (N_2827,N_2456,N_2400);
nand U2828 (N_2828,N_2058,N_2099);
nor U2829 (N_2829,N_2449,N_2002);
and U2830 (N_2830,N_2478,N_2354);
and U2831 (N_2831,N_2130,N_2158);
nand U2832 (N_2832,N_2078,N_2302);
and U2833 (N_2833,N_2043,N_2369);
or U2834 (N_2834,N_2003,N_2062);
nand U2835 (N_2835,N_2299,N_2381);
nor U2836 (N_2836,N_2272,N_2050);
nand U2837 (N_2837,N_2195,N_2351);
nor U2838 (N_2838,N_2331,N_2158);
or U2839 (N_2839,N_2290,N_2494);
xnor U2840 (N_2840,N_2219,N_2151);
xnor U2841 (N_2841,N_2354,N_2278);
xnor U2842 (N_2842,N_2371,N_2071);
nor U2843 (N_2843,N_2380,N_2235);
xnor U2844 (N_2844,N_2352,N_2010);
nor U2845 (N_2845,N_2335,N_2310);
xor U2846 (N_2846,N_2039,N_2214);
nand U2847 (N_2847,N_2068,N_2112);
and U2848 (N_2848,N_2018,N_2354);
nor U2849 (N_2849,N_2013,N_2432);
nand U2850 (N_2850,N_2262,N_2044);
nand U2851 (N_2851,N_2210,N_2446);
nand U2852 (N_2852,N_2467,N_2236);
and U2853 (N_2853,N_2339,N_2284);
and U2854 (N_2854,N_2084,N_2142);
nor U2855 (N_2855,N_2116,N_2471);
and U2856 (N_2856,N_2451,N_2322);
or U2857 (N_2857,N_2445,N_2287);
or U2858 (N_2858,N_2166,N_2101);
xor U2859 (N_2859,N_2490,N_2277);
nand U2860 (N_2860,N_2287,N_2118);
and U2861 (N_2861,N_2046,N_2105);
or U2862 (N_2862,N_2125,N_2471);
or U2863 (N_2863,N_2176,N_2373);
or U2864 (N_2864,N_2443,N_2268);
nand U2865 (N_2865,N_2269,N_2449);
and U2866 (N_2866,N_2004,N_2133);
xnor U2867 (N_2867,N_2282,N_2478);
nand U2868 (N_2868,N_2265,N_2084);
xor U2869 (N_2869,N_2083,N_2064);
nand U2870 (N_2870,N_2267,N_2482);
or U2871 (N_2871,N_2491,N_2026);
or U2872 (N_2872,N_2293,N_2337);
or U2873 (N_2873,N_2348,N_2334);
nand U2874 (N_2874,N_2373,N_2106);
xor U2875 (N_2875,N_2289,N_2265);
nor U2876 (N_2876,N_2126,N_2142);
or U2877 (N_2877,N_2364,N_2074);
nor U2878 (N_2878,N_2090,N_2241);
and U2879 (N_2879,N_2411,N_2150);
nand U2880 (N_2880,N_2499,N_2067);
nand U2881 (N_2881,N_2277,N_2325);
or U2882 (N_2882,N_2011,N_2091);
xnor U2883 (N_2883,N_2183,N_2211);
nor U2884 (N_2884,N_2140,N_2444);
nand U2885 (N_2885,N_2433,N_2006);
and U2886 (N_2886,N_2499,N_2163);
and U2887 (N_2887,N_2175,N_2300);
nor U2888 (N_2888,N_2160,N_2297);
and U2889 (N_2889,N_2136,N_2063);
xnor U2890 (N_2890,N_2460,N_2286);
and U2891 (N_2891,N_2404,N_2449);
or U2892 (N_2892,N_2308,N_2111);
and U2893 (N_2893,N_2336,N_2257);
nand U2894 (N_2894,N_2036,N_2475);
and U2895 (N_2895,N_2307,N_2324);
nand U2896 (N_2896,N_2024,N_2484);
nand U2897 (N_2897,N_2168,N_2437);
nor U2898 (N_2898,N_2430,N_2151);
nand U2899 (N_2899,N_2444,N_2370);
xnor U2900 (N_2900,N_2390,N_2003);
xor U2901 (N_2901,N_2246,N_2217);
xor U2902 (N_2902,N_2378,N_2431);
or U2903 (N_2903,N_2365,N_2122);
xnor U2904 (N_2904,N_2453,N_2493);
or U2905 (N_2905,N_2475,N_2282);
and U2906 (N_2906,N_2052,N_2109);
nand U2907 (N_2907,N_2238,N_2004);
and U2908 (N_2908,N_2099,N_2401);
or U2909 (N_2909,N_2351,N_2419);
and U2910 (N_2910,N_2100,N_2305);
and U2911 (N_2911,N_2290,N_2250);
nand U2912 (N_2912,N_2012,N_2032);
and U2913 (N_2913,N_2388,N_2282);
nand U2914 (N_2914,N_2399,N_2179);
nor U2915 (N_2915,N_2183,N_2452);
and U2916 (N_2916,N_2056,N_2215);
xor U2917 (N_2917,N_2217,N_2437);
or U2918 (N_2918,N_2390,N_2264);
nand U2919 (N_2919,N_2300,N_2374);
nand U2920 (N_2920,N_2076,N_2437);
xnor U2921 (N_2921,N_2241,N_2034);
xor U2922 (N_2922,N_2112,N_2197);
or U2923 (N_2923,N_2370,N_2302);
or U2924 (N_2924,N_2353,N_2060);
and U2925 (N_2925,N_2241,N_2222);
nor U2926 (N_2926,N_2434,N_2156);
nor U2927 (N_2927,N_2326,N_2209);
or U2928 (N_2928,N_2219,N_2468);
or U2929 (N_2929,N_2229,N_2308);
nor U2930 (N_2930,N_2353,N_2023);
nor U2931 (N_2931,N_2076,N_2283);
or U2932 (N_2932,N_2090,N_2478);
nand U2933 (N_2933,N_2115,N_2338);
or U2934 (N_2934,N_2341,N_2310);
xnor U2935 (N_2935,N_2023,N_2286);
or U2936 (N_2936,N_2119,N_2074);
nand U2937 (N_2937,N_2490,N_2439);
and U2938 (N_2938,N_2106,N_2477);
or U2939 (N_2939,N_2371,N_2236);
nor U2940 (N_2940,N_2064,N_2390);
xnor U2941 (N_2941,N_2365,N_2103);
and U2942 (N_2942,N_2265,N_2368);
or U2943 (N_2943,N_2317,N_2234);
xor U2944 (N_2944,N_2029,N_2162);
and U2945 (N_2945,N_2096,N_2153);
xor U2946 (N_2946,N_2434,N_2037);
xnor U2947 (N_2947,N_2454,N_2470);
xor U2948 (N_2948,N_2405,N_2303);
nand U2949 (N_2949,N_2314,N_2275);
or U2950 (N_2950,N_2099,N_2345);
xor U2951 (N_2951,N_2239,N_2176);
xnor U2952 (N_2952,N_2049,N_2317);
nor U2953 (N_2953,N_2197,N_2414);
and U2954 (N_2954,N_2014,N_2167);
xor U2955 (N_2955,N_2368,N_2375);
xnor U2956 (N_2956,N_2206,N_2480);
and U2957 (N_2957,N_2080,N_2444);
nand U2958 (N_2958,N_2017,N_2197);
nor U2959 (N_2959,N_2079,N_2221);
nor U2960 (N_2960,N_2280,N_2172);
nor U2961 (N_2961,N_2254,N_2268);
or U2962 (N_2962,N_2264,N_2033);
xnor U2963 (N_2963,N_2359,N_2002);
nand U2964 (N_2964,N_2335,N_2379);
or U2965 (N_2965,N_2421,N_2132);
and U2966 (N_2966,N_2402,N_2420);
and U2967 (N_2967,N_2083,N_2045);
and U2968 (N_2968,N_2434,N_2187);
nor U2969 (N_2969,N_2313,N_2221);
xor U2970 (N_2970,N_2184,N_2030);
and U2971 (N_2971,N_2368,N_2377);
nand U2972 (N_2972,N_2144,N_2486);
nor U2973 (N_2973,N_2398,N_2346);
nor U2974 (N_2974,N_2332,N_2228);
or U2975 (N_2975,N_2012,N_2128);
and U2976 (N_2976,N_2265,N_2142);
xor U2977 (N_2977,N_2395,N_2201);
or U2978 (N_2978,N_2204,N_2244);
nor U2979 (N_2979,N_2151,N_2232);
xnor U2980 (N_2980,N_2034,N_2060);
xor U2981 (N_2981,N_2309,N_2227);
and U2982 (N_2982,N_2093,N_2183);
xnor U2983 (N_2983,N_2496,N_2355);
and U2984 (N_2984,N_2012,N_2499);
nand U2985 (N_2985,N_2220,N_2036);
or U2986 (N_2986,N_2356,N_2112);
and U2987 (N_2987,N_2015,N_2467);
nand U2988 (N_2988,N_2277,N_2009);
xor U2989 (N_2989,N_2453,N_2448);
and U2990 (N_2990,N_2228,N_2456);
or U2991 (N_2991,N_2179,N_2311);
and U2992 (N_2992,N_2037,N_2429);
nand U2993 (N_2993,N_2388,N_2030);
nand U2994 (N_2994,N_2083,N_2231);
or U2995 (N_2995,N_2174,N_2474);
xnor U2996 (N_2996,N_2146,N_2199);
nand U2997 (N_2997,N_2124,N_2125);
nor U2998 (N_2998,N_2152,N_2324);
and U2999 (N_2999,N_2132,N_2304);
or U3000 (N_3000,N_2970,N_2761);
or U3001 (N_3001,N_2561,N_2788);
nor U3002 (N_3002,N_2839,N_2612);
or U3003 (N_3003,N_2724,N_2908);
nand U3004 (N_3004,N_2840,N_2722);
and U3005 (N_3005,N_2917,N_2637);
or U3006 (N_3006,N_2543,N_2711);
nand U3007 (N_3007,N_2736,N_2662);
xor U3008 (N_3008,N_2720,N_2525);
and U3009 (N_3009,N_2687,N_2732);
xnor U3010 (N_3010,N_2654,N_2815);
or U3011 (N_3011,N_2857,N_2795);
and U3012 (N_3012,N_2876,N_2506);
nand U3013 (N_3013,N_2709,N_2733);
and U3014 (N_3014,N_2865,N_2877);
xnor U3015 (N_3015,N_2640,N_2534);
xor U3016 (N_3016,N_2820,N_2671);
and U3017 (N_3017,N_2993,N_2901);
xnor U3018 (N_3018,N_2717,N_2558);
and U3019 (N_3019,N_2953,N_2578);
and U3020 (N_3020,N_2962,N_2951);
nand U3021 (N_3021,N_2582,N_2816);
or U3022 (N_3022,N_2676,N_2811);
nand U3023 (N_3023,N_2950,N_2926);
nand U3024 (N_3024,N_2505,N_2801);
and U3025 (N_3025,N_2531,N_2763);
nand U3026 (N_3026,N_2939,N_2862);
nand U3027 (N_3027,N_2828,N_2764);
nand U3028 (N_3028,N_2725,N_2686);
nor U3029 (N_3029,N_2872,N_2672);
nor U3030 (N_3030,N_2988,N_2976);
or U3031 (N_3031,N_2690,N_2907);
nor U3032 (N_3032,N_2704,N_2797);
nor U3033 (N_3033,N_2632,N_2739);
nand U3034 (N_3034,N_2581,N_2730);
nor U3035 (N_3035,N_2875,N_2874);
or U3036 (N_3036,N_2835,N_2842);
nor U3037 (N_3037,N_2997,N_2963);
nor U3038 (N_3038,N_2501,N_2870);
nand U3039 (N_3039,N_2579,N_2802);
xor U3040 (N_3040,N_2555,N_2848);
nor U3041 (N_3041,N_2734,N_2931);
and U3042 (N_3042,N_2775,N_2933);
nand U3043 (N_3043,N_2726,N_2718);
nand U3044 (N_3044,N_2861,N_2985);
nand U3045 (N_3045,N_2992,N_2750);
nand U3046 (N_3046,N_2616,N_2751);
and U3047 (N_3047,N_2667,N_2510);
nand U3048 (N_3048,N_2943,N_2559);
nor U3049 (N_3049,N_2879,N_2834);
and U3050 (N_3050,N_2833,N_2871);
and U3051 (N_3051,N_2584,N_2526);
xor U3052 (N_3052,N_2844,N_2785);
nand U3053 (N_3053,N_2883,N_2841);
nand U3054 (N_3054,N_2850,N_2509);
nor U3055 (N_3055,N_2999,N_2779);
or U3056 (N_3056,N_2629,N_2602);
or U3057 (N_3057,N_2758,N_2936);
nor U3058 (N_3058,N_2888,N_2500);
nor U3059 (N_3059,N_2530,N_2817);
and U3060 (N_3060,N_2603,N_2836);
and U3061 (N_3061,N_2956,N_2716);
xnor U3062 (N_3062,N_2681,N_2896);
xnor U3063 (N_3063,N_2884,N_2567);
nor U3064 (N_3064,N_2787,N_2575);
or U3065 (N_3065,N_2967,N_2913);
xor U3066 (N_3066,N_2646,N_2903);
nor U3067 (N_3067,N_2929,N_2891);
or U3068 (N_3068,N_2606,N_2807);
nor U3069 (N_3069,N_2854,N_2916);
nor U3070 (N_3070,N_2539,N_2631);
xnor U3071 (N_3071,N_2564,N_2762);
nor U3072 (N_3072,N_2759,N_2705);
and U3073 (N_3073,N_2623,N_2904);
nor U3074 (N_3074,N_2978,N_2957);
or U3075 (N_3075,N_2927,N_2975);
or U3076 (N_3076,N_2952,N_2912);
or U3077 (N_3077,N_2695,N_2812);
or U3078 (N_3078,N_2626,N_2678);
and U3079 (N_3079,N_2809,N_2987);
and U3080 (N_3080,N_2565,N_2982);
and U3081 (N_3081,N_2691,N_2521);
xnor U3082 (N_3082,N_2906,N_2799);
and U3083 (N_3083,N_2911,N_2885);
nand U3084 (N_3084,N_2659,N_2635);
or U3085 (N_3085,N_2921,N_2878);
nor U3086 (N_3086,N_2557,N_2601);
nor U3087 (N_3087,N_2728,N_2591);
or U3088 (N_3088,N_2533,N_2778);
nor U3089 (N_3089,N_2965,N_2658);
nand U3090 (N_3090,N_2648,N_2998);
nand U3091 (N_3091,N_2502,N_2666);
xor U3092 (N_3092,N_2613,N_2556);
or U3093 (N_3093,N_2715,N_2846);
nor U3094 (N_3094,N_2618,N_2580);
nor U3095 (N_3095,N_2627,N_2856);
xnor U3096 (N_3096,N_2511,N_2949);
nand U3097 (N_3097,N_2808,N_2860);
nand U3098 (N_3098,N_2920,N_2643);
xnor U3099 (N_3099,N_2925,N_2712);
and U3100 (N_3100,N_2864,N_2609);
or U3101 (N_3101,N_2889,N_2593);
nand U3102 (N_3102,N_2919,N_2605);
nand U3103 (N_3103,N_2589,N_2744);
nor U3104 (N_3104,N_2905,N_2610);
xor U3105 (N_3105,N_2914,N_2946);
or U3106 (N_3106,N_2973,N_2628);
nand U3107 (N_3107,N_2524,N_2600);
or U3108 (N_3108,N_2981,N_2882);
nor U3109 (N_3109,N_2657,N_2831);
and U3110 (N_3110,N_2624,N_2818);
xor U3111 (N_3111,N_2793,N_2881);
xnor U3112 (N_3112,N_2650,N_2832);
and U3113 (N_3113,N_2587,N_2960);
and U3114 (N_3114,N_2858,N_2958);
xnor U3115 (N_3115,N_2644,N_2607);
nand U3116 (N_3116,N_2670,N_2701);
xnor U3117 (N_3117,N_2642,N_2548);
nand U3118 (N_3118,N_2886,N_2512);
nand U3119 (N_3119,N_2697,N_2867);
or U3120 (N_3120,N_2824,N_2772);
xnor U3121 (N_3121,N_2576,N_2677);
xor U3122 (N_3122,N_2934,N_2549);
and U3123 (N_3123,N_2866,N_2767);
nand U3124 (N_3124,N_2868,N_2566);
and U3125 (N_3125,N_2852,N_2710);
nand U3126 (N_3126,N_2892,N_2663);
or U3127 (N_3127,N_2898,N_2563);
nor U3128 (N_3128,N_2942,N_2765);
or U3129 (N_3129,N_2518,N_2741);
nor U3130 (N_3130,N_2777,N_2544);
nor U3131 (N_3131,N_2928,N_2621);
nand U3132 (N_3132,N_2887,N_2966);
nand U3133 (N_3133,N_2800,N_2707);
nor U3134 (N_3134,N_2829,N_2656);
or U3135 (N_3135,N_2682,N_2989);
nor U3136 (N_3136,N_2652,N_2814);
nor U3137 (N_3137,N_2838,N_2837);
nor U3138 (N_3138,N_2507,N_2645);
nor U3139 (N_3139,N_2994,N_2774);
xor U3140 (N_3140,N_2937,N_2855);
xor U3141 (N_3141,N_2708,N_2536);
nor U3142 (N_3142,N_2508,N_2542);
and U3143 (N_3143,N_2968,N_2633);
and U3144 (N_3144,N_2940,N_2743);
nand U3145 (N_3145,N_2528,N_2696);
nor U3146 (N_3146,N_2519,N_2504);
and U3147 (N_3147,N_2714,N_2706);
xor U3148 (N_3148,N_2932,N_2794);
nor U3149 (N_3149,N_2685,N_2611);
or U3150 (N_3150,N_2661,N_2964);
nor U3151 (N_3151,N_2770,N_2537);
nor U3152 (N_3152,N_2747,N_2959);
or U3153 (N_3153,N_2547,N_2798);
nor U3154 (N_3154,N_2822,N_2955);
nor U3155 (N_3155,N_2604,N_2550);
and U3156 (N_3156,N_2961,N_2853);
and U3157 (N_3157,N_2740,N_2782);
and U3158 (N_3158,N_2698,N_2748);
and U3159 (N_3159,N_2620,N_2583);
xor U3160 (N_3160,N_2649,N_2938);
or U3161 (N_3161,N_2595,N_2894);
xor U3162 (N_3162,N_2986,N_2538);
and U3163 (N_3163,N_2909,N_2630);
and U3164 (N_3164,N_2599,N_2684);
nor U3165 (N_3165,N_2945,N_2766);
or U3166 (N_3166,N_2980,N_2924);
and U3167 (N_3167,N_2796,N_2668);
xor U3168 (N_3168,N_2689,N_2810);
nand U3169 (N_3169,N_2893,N_2863);
xor U3170 (N_3170,N_2664,N_2520);
or U3171 (N_3171,N_2890,N_2948);
xor U3172 (N_3172,N_2673,N_2830);
nand U3173 (N_3173,N_2918,N_2615);
xnor U3174 (N_3174,N_2574,N_2760);
nor U3175 (N_3175,N_2780,N_2895);
xor U3176 (N_3176,N_2523,N_2922);
and U3177 (N_3177,N_2639,N_2634);
nor U3178 (N_3178,N_2803,N_2827);
or U3179 (N_3179,N_2843,N_2745);
nor U3180 (N_3180,N_2823,N_2608);
xnor U3181 (N_3181,N_2713,N_2572);
and U3182 (N_3182,N_2791,N_2983);
xor U3183 (N_3183,N_2915,N_2619);
and U3184 (N_3184,N_2792,N_2923);
or U3185 (N_3185,N_2516,N_2776);
nor U3186 (N_3186,N_2617,N_2503);
xnor U3187 (N_3187,N_2995,N_2757);
xnor U3188 (N_3188,N_2790,N_2969);
nand U3189 (N_3189,N_2804,N_2522);
and U3190 (N_3190,N_2996,N_2692);
or U3191 (N_3191,N_2570,N_2674);
nand U3192 (N_3192,N_2641,N_2694);
nor U3193 (N_3193,N_2753,N_2586);
and U3194 (N_3194,N_2669,N_2727);
nand U3195 (N_3195,N_2910,N_2573);
nand U3196 (N_3196,N_2768,N_2821);
and U3197 (N_3197,N_2665,N_2638);
or U3198 (N_3198,N_2897,N_2781);
and U3199 (N_3199,N_2755,N_2954);
or U3200 (N_3200,N_2545,N_2974);
and U3201 (N_3201,N_2699,N_2568);
and U3202 (N_3202,N_2742,N_2683);
or U3203 (N_3203,N_2622,N_2737);
or U3204 (N_3204,N_2902,N_2571);
nand U3205 (N_3205,N_2752,N_2806);
nand U3206 (N_3206,N_2845,N_2731);
xor U3207 (N_3207,N_2693,N_2721);
xor U3208 (N_3208,N_2977,N_2513);
and U3209 (N_3209,N_2554,N_2813);
xor U3210 (N_3210,N_2738,N_2562);
or U3211 (N_3211,N_2851,N_2700);
and U3212 (N_3212,N_2746,N_2947);
nand U3213 (N_3213,N_2535,N_2703);
xnor U3214 (N_3214,N_2979,N_2869);
and U3215 (N_3215,N_2756,N_2551);
or U3216 (N_3216,N_2873,N_2517);
and U3217 (N_3217,N_2679,N_2552);
and U3218 (N_3218,N_2651,N_2546);
xor U3219 (N_3219,N_2729,N_2749);
and U3220 (N_3220,N_2688,N_2636);
xor U3221 (N_3221,N_2569,N_2675);
and U3222 (N_3222,N_2597,N_2719);
or U3223 (N_3223,N_2585,N_2805);
nand U3224 (N_3224,N_2930,N_2577);
xor U3225 (N_3225,N_2614,N_2984);
or U3226 (N_3226,N_2527,N_2847);
nor U3227 (N_3227,N_2900,N_2769);
or U3228 (N_3228,N_2849,N_2596);
xnor U3229 (N_3229,N_2592,N_2944);
or U3230 (N_3230,N_2941,N_2541);
nor U3231 (N_3231,N_2625,N_2825);
and U3232 (N_3232,N_2789,N_2723);
or U3233 (N_3233,N_2783,N_2972);
nor U3234 (N_3234,N_2532,N_2819);
and U3235 (N_3235,N_2588,N_2647);
and U3236 (N_3236,N_2660,N_2702);
xnor U3237 (N_3237,N_2529,N_2655);
or U3238 (N_3238,N_2990,N_2773);
xor U3239 (N_3239,N_2680,N_2971);
and U3240 (N_3240,N_2515,N_2653);
xnor U3241 (N_3241,N_2594,N_2754);
nand U3242 (N_3242,N_2560,N_2553);
or U3243 (N_3243,N_2771,N_2540);
nor U3244 (N_3244,N_2899,N_2514);
nor U3245 (N_3245,N_2935,N_2598);
or U3246 (N_3246,N_2784,N_2859);
nor U3247 (N_3247,N_2590,N_2786);
nor U3248 (N_3248,N_2735,N_2991);
nor U3249 (N_3249,N_2880,N_2826);
or U3250 (N_3250,N_2745,N_2610);
or U3251 (N_3251,N_2929,N_2782);
xor U3252 (N_3252,N_2844,N_2597);
and U3253 (N_3253,N_2595,N_2995);
or U3254 (N_3254,N_2658,N_2859);
and U3255 (N_3255,N_2927,N_2896);
nand U3256 (N_3256,N_2736,N_2764);
nand U3257 (N_3257,N_2606,N_2828);
nor U3258 (N_3258,N_2652,N_2801);
nor U3259 (N_3259,N_2834,N_2864);
xnor U3260 (N_3260,N_2566,N_2530);
nand U3261 (N_3261,N_2788,N_2647);
nand U3262 (N_3262,N_2871,N_2781);
nor U3263 (N_3263,N_2712,N_2834);
xor U3264 (N_3264,N_2507,N_2983);
or U3265 (N_3265,N_2637,N_2689);
xor U3266 (N_3266,N_2505,N_2951);
or U3267 (N_3267,N_2603,N_2769);
or U3268 (N_3268,N_2962,N_2810);
xnor U3269 (N_3269,N_2535,N_2866);
nor U3270 (N_3270,N_2702,N_2841);
nor U3271 (N_3271,N_2595,N_2535);
nor U3272 (N_3272,N_2520,N_2696);
or U3273 (N_3273,N_2512,N_2609);
xor U3274 (N_3274,N_2755,N_2556);
nand U3275 (N_3275,N_2786,N_2872);
xnor U3276 (N_3276,N_2628,N_2862);
nor U3277 (N_3277,N_2773,N_2944);
or U3278 (N_3278,N_2957,N_2958);
xnor U3279 (N_3279,N_2695,N_2611);
and U3280 (N_3280,N_2625,N_2626);
nand U3281 (N_3281,N_2945,N_2991);
and U3282 (N_3282,N_2547,N_2736);
nand U3283 (N_3283,N_2540,N_2588);
xor U3284 (N_3284,N_2613,N_2854);
xor U3285 (N_3285,N_2986,N_2890);
or U3286 (N_3286,N_2642,N_2711);
xnor U3287 (N_3287,N_2900,N_2889);
nor U3288 (N_3288,N_2790,N_2723);
and U3289 (N_3289,N_2740,N_2829);
and U3290 (N_3290,N_2555,N_2962);
nand U3291 (N_3291,N_2708,N_2857);
or U3292 (N_3292,N_2990,N_2850);
or U3293 (N_3293,N_2729,N_2936);
xor U3294 (N_3294,N_2525,N_2999);
or U3295 (N_3295,N_2777,N_2704);
and U3296 (N_3296,N_2947,N_2998);
and U3297 (N_3297,N_2892,N_2912);
and U3298 (N_3298,N_2569,N_2651);
xor U3299 (N_3299,N_2556,N_2858);
xnor U3300 (N_3300,N_2792,N_2655);
or U3301 (N_3301,N_2553,N_2725);
xor U3302 (N_3302,N_2646,N_2652);
and U3303 (N_3303,N_2650,N_2600);
nand U3304 (N_3304,N_2632,N_2836);
and U3305 (N_3305,N_2625,N_2597);
nand U3306 (N_3306,N_2701,N_2630);
and U3307 (N_3307,N_2508,N_2774);
xor U3308 (N_3308,N_2847,N_2538);
xnor U3309 (N_3309,N_2814,N_2582);
nor U3310 (N_3310,N_2593,N_2936);
or U3311 (N_3311,N_2630,N_2929);
nand U3312 (N_3312,N_2947,N_2634);
nor U3313 (N_3313,N_2627,N_2733);
or U3314 (N_3314,N_2887,N_2766);
nand U3315 (N_3315,N_2599,N_2514);
or U3316 (N_3316,N_2793,N_2918);
nor U3317 (N_3317,N_2724,N_2973);
xnor U3318 (N_3318,N_2565,N_2507);
nor U3319 (N_3319,N_2825,N_2530);
or U3320 (N_3320,N_2762,N_2955);
nand U3321 (N_3321,N_2733,N_2968);
nand U3322 (N_3322,N_2861,N_2730);
xnor U3323 (N_3323,N_2985,N_2804);
nand U3324 (N_3324,N_2777,N_2670);
nor U3325 (N_3325,N_2820,N_2738);
or U3326 (N_3326,N_2805,N_2788);
xnor U3327 (N_3327,N_2568,N_2987);
xor U3328 (N_3328,N_2889,N_2726);
nand U3329 (N_3329,N_2538,N_2962);
and U3330 (N_3330,N_2985,N_2942);
xor U3331 (N_3331,N_2553,N_2637);
or U3332 (N_3332,N_2518,N_2856);
nand U3333 (N_3333,N_2769,N_2692);
xor U3334 (N_3334,N_2744,N_2796);
nor U3335 (N_3335,N_2976,N_2539);
or U3336 (N_3336,N_2746,N_2724);
and U3337 (N_3337,N_2770,N_2834);
nand U3338 (N_3338,N_2933,N_2797);
nand U3339 (N_3339,N_2735,N_2705);
nor U3340 (N_3340,N_2680,N_2833);
xnor U3341 (N_3341,N_2796,N_2736);
or U3342 (N_3342,N_2767,N_2921);
and U3343 (N_3343,N_2557,N_2794);
or U3344 (N_3344,N_2532,N_2510);
or U3345 (N_3345,N_2895,N_2685);
or U3346 (N_3346,N_2620,N_2702);
xnor U3347 (N_3347,N_2813,N_2961);
xnor U3348 (N_3348,N_2765,N_2763);
nand U3349 (N_3349,N_2683,N_2694);
nand U3350 (N_3350,N_2575,N_2629);
and U3351 (N_3351,N_2647,N_2666);
xnor U3352 (N_3352,N_2956,N_2609);
and U3353 (N_3353,N_2713,N_2596);
nand U3354 (N_3354,N_2591,N_2524);
or U3355 (N_3355,N_2528,N_2730);
nor U3356 (N_3356,N_2627,N_2846);
or U3357 (N_3357,N_2962,N_2707);
or U3358 (N_3358,N_2671,N_2504);
and U3359 (N_3359,N_2585,N_2848);
nor U3360 (N_3360,N_2863,N_2917);
xnor U3361 (N_3361,N_2501,N_2839);
or U3362 (N_3362,N_2862,N_2951);
and U3363 (N_3363,N_2808,N_2505);
xnor U3364 (N_3364,N_2737,N_2547);
or U3365 (N_3365,N_2874,N_2566);
nand U3366 (N_3366,N_2980,N_2762);
xor U3367 (N_3367,N_2955,N_2704);
nor U3368 (N_3368,N_2593,N_2899);
and U3369 (N_3369,N_2850,N_2855);
or U3370 (N_3370,N_2620,N_2672);
or U3371 (N_3371,N_2519,N_2699);
or U3372 (N_3372,N_2655,N_2806);
nand U3373 (N_3373,N_2580,N_2935);
xor U3374 (N_3374,N_2940,N_2690);
xnor U3375 (N_3375,N_2757,N_2791);
nor U3376 (N_3376,N_2872,N_2537);
and U3377 (N_3377,N_2624,N_2700);
xnor U3378 (N_3378,N_2888,N_2538);
nor U3379 (N_3379,N_2983,N_2922);
xnor U3380 (N_3380,N_2513,N_2972);
nand U3381 (N_3381,N_2655,N_2840);
or U3382 (N_3382,N_2811,N_2860);
nand U3383 (N_3383,N_2580,N_2505);
nor U3384 (N_3384,N_2652,N_2636);
nor U3385 (N_3385,N_2905,N_2760);
nor U3386 (N_3386,N_2936,N_2889);
or U3387 (N_3387,N_2877,N_2643);
and U3388 (N_3388,N_2534,N_2768);
nor U3389 (N_3389,N_2932,N_2636);
and U3390 (N_3390,N_2567,N_2500);
xor U3391 (N_3391,N_2564,N_2947);
or U3392 (N_3392,N_2765,N_2962);
nor U3393 (N_3393,N_2510,N_2557);
nor U3394 (N_3394,N_2604,N_2933);
and U3395 (N_3395,N_2953,N_2807);
nand U3396 (N_3396,N_2639,N_2626);
xnor U3397 (N_3397,N_2995,N_2748);
xnor U3398 (N_3398,N_2969,N_2932);
nand U3399 (N_3399,N_2855,N_2732);
nor U3400 (N_3400,N_2972,N_2680);
or U3401 (N_3401,N_2714,N_2746);
nand U3402 (N_3402,N_2654,N_2630);
or U3403 (N_3403,N_2724,N_2807);
nand U3404 (N_3404,N_2779,N_2802);
or U3405 (N_3405,N_2639,N_2727);
or U3406 (N_3406,N_2903,N_2533);
and U3407 (N_3407,N_2996,N_2781);
xnor U3408 (N_3408,N_2827,N_2792);
or U3409 (N_3409,N_2926,N_2647);
nand U3410 (N_3410,N_2886,N_2593);
xnor U3411 (N_3411,N_2541,N_2915);
nor U3412 (N_3412,N_2797,N_2855);
nor U3413 (N_3413,N_2762,N_2847);
nor U3414 (N_3414,N_2796,N_2714);
nand U3415 (N_3415,N_2960,N_2746);
xnor U3416 (N_3416,N_2994,N_2723);
nand U3417 (N_3417,N_2533,N_2670);
nand U3418 (N_3418,N_2611,N_2963);
and U3419 (N_3419,N_2919,N_2723);
nand U3420 (N_3420,N_2936,N_2894);
xor U3421 (N_3421,N_2654,N_2993);
nand U3422 (N_3422,N_2659,N_2797);
nor U3423 (N_3423,N_2887,N_2620);
nor U3424 (N_3424,N_2626,N_2569);
nor U3425 (N_3425,N_2973,N_2529);
nor U3426 (N_3426,N_2532,N_2773);
and U3427 (N_3427,N_2889,N_2789);
xnor U3428 (N_3428,N_2986,N_2781);
nor U3429 (N_3429,N_2738,N_2550);
nand U3430 (N_3430,N_2844,N_2581);
nor U3431 (N_3431,N_2597,N_2865);
or U3432 (N_3432,N_2659,N_2693);
nand U3433 (N_3433,N_2897,N_2649);
and U3434 (N_3434,N_2619,N_2648);
nor U3435 (N_3435,N_2723,N_2892);
nor U3436 (N_3436,N_2784,N_2552);
and U3437 (N_3437,N_2799,N_2582);
nand U3438 (N_3438,N_2729,N_2533);
xnor U3439 (N_3439,N_2661,N_2580);
nor U3440 (N_3440,N_2686,N_2855);
xnor U3441 (N_3441,N_2969,N_2890);
or U3442 (N_3442,N_2608,N_2846);
nand U3443 (N_3443,N_2570,N_2918);
xor U3444 (N_3444,N_2620,N_2693);
nand U3445 (N_3445,N_2816,N_2921);
nand U3446 (N_3446,N_2938,N_2953);
nand U3447 (N_3447,N_2640,N_2518);
nand U3448 (N_3448,N_2875,N_2933);
nand U3449 (N_3449,N_2647,N_2978);
or U3450 (N_3450,N_2625,N_2920);
or U3451 (N_3451,N_2723,N_2616);
xor U3452 (N_3452,N_2651,N_2506);
or U3453 (N_3453,N_2877,N_2921);
nor U3454 (N_3454,N_2988,N_2596);
nor U3455 (N_3455,N_2613,N_2759);
nand U3456 (N_3456,N_2688,N_2947);
or U3457 (N_3457,N_2540,N_2800);
or U3458 (N_3458,N_2585,N_2588);
nand U3459 (N_3459,N_2558,N_2659);
nand U3460 (N_3460,N_2611,N_2529);
nand U3461 (N_3461,N_2573,N_2623);
and U3462 (N_3462,N_2575,N_2545);
nand U3463 (N_3463,N_2937,N_2814);
nand U3464 (N_3464,N_2864,N_2655);
nand U3465 (N_3465,N_2554,N_2812);
xor U3466 (N_3466,N_2755,N_2699);
xor U3467 (N_3467,N_2583,N_2578);
nor U3468 (N_3468,N_2678,N_2683);
nor U3469 (N_3469,N_2916,N_2856);
nand U3470 (N_3470,N_2813,N_2508);
or U3471 (N_3471,N_2769,N_2748);
nand U3472 (N_3472,N_2844,N_2624);
nor U3473 (N_3473,N_2618,N_2742);
and U3474 (N_3474,N_2649,N_2761);
nor U3475 (N_3475,N_2711,N_2639);
or U3476 (N_3476,N_2823,N_2578);
nor U3477 (N_3477,N_2615,N_2733);
or U3478 (N_3478,N_2776,N_2967);
nor U3479 (N_3479,N_2792,N_2813);
or U3480 (N_3480,N_2606,N_2763);
nor U3481 (N_3481,N_2504,N_2788);
xnor U3482 (N_3482,N_2712,N_2939);
or U3483 (N_3483,N_2710,N_2542);
and U3484 (N_3484,N_2727,N_2894);
or U3485 (N_3485,N_2554,N_2567);
or U3486 (N_3486,N_2510,N_2695);
xor U3487 (N_3487,N_2551,N_2959);
xor U3488 (N_3488,N_2596,N_2676);
or U3489 (N_3489,N_2541,N_2866);
nand U3490 (N_3490,N_2603,N_2913);
nand U3491 (N_3491,N_2699,N_2708);
nand U3492 (N_3492,N_2785,N_2958);
and U3493 (N_3493,N_2921,N_2585);
xor U3494 (N_3494,N_2560,N_2884);
nand U3495 (N_3495,N_2808,N_2938);
nor U3496 (N_3496,N_2683,N_2793);
or U3497 (N_3497,N_2879,N_2734);
nand U3498 (N_3498,N_2956,N_2822);
or U3499 (N_3499,N_2965,N_2523);
nor U3500 (N_3500,N_3262,N_3157);
nand U3501 (N_3501,N_3216,N_3356);
nand U3502 (N_3502,N_3219,N_3451);
and U3503 (N_3503,N_3105,N_3231);
or U3504 (N_3504,N_3286,N_3166);
nand U3505 (N_3505,N_3028,N_3236);
and U3506 (N_3506,N_3131,N_3283);
nor U3507 (N_3507,N_3434,N_3189);
nand U3508 (N_3508,N_3387,N_3490);
nor U3509 (N_3509,N_3246,N_3017);
nor U3510 (N_3510,N_3056,N_3297);
nor U3511 (N_3511,N_3104,N_3433);
or U3512 (N_3512,N_3372,N_3335);
nor U3513 (N_3513,N_3315,N_3051);
xor U3514 (N_3514,N_3244,N_3429);
or U3515 (N_3515,N_3467,N_3369);
xnor U3516 (N_3516,N_3426,N_3247);
nand U3517 (N_3517,N_3079,N_3025);
nor U3518 (N_3518,N_3242,N_3052);
nand U3519 (N_3519,N_3156,N_3403);
or U3520 (N_3520,N_3260,N_3305);
or U3521 (N_3521,N_3319,N_3098);
nand U3522 (N_3522,N_3078,N_3340);
nor U3523 (N_3523,N_3459,N_3243);
nor U3524 (N_3524,N_3053,N_3210);
nor U3525 (N_3525,N_3087,N_3313);
nand U3526 (N_3526,N_3148,N_3227);
nand U3527 (N_3527,N_3392,N_3018);
nor U3528 (N_3528,N_3465,N_3034);
xnor U3529 (N_3529,N_3419,N_3456);
and U3530 (N_3530,N_3149,N_3327);
nand U3531 (N_3531,N_3442,N_3365);
nor U3532 (N_3532,N_3486,N_3291);
and U3533 (N_3533,N_3310,N_3440);
xnor U3534 (N_3534,N_3274,N_3135);
or U3535 (N_3535,N_3094,N_3101);
nand U3536 (N_3536,N_3499,N_3031);
nor U3537 (N_3537,N_3000,N_3437);
nor U3538 (N_3538,N_3288,N_3237);
nand U3539 (N_3539,N_3133,N_3136);
nand U3540 (N_3540,N_3225,N_3108);
xnor U3541 (N_3541,N_3151,N_3004);
nand U3542 (N_3542,N_3479,N_3117);
nand U3543 (N_3543,N_3386,N_3468);
or U3544 (N_3544,N_3081,N_3047);
nor U3545 (N_3545,N_3044,N_3445);
xnor U3546 (N_3546,N_3383,N_3495);
and U3547 (N_3547,N_3185,N_3298);
or U3548 (N_3548,N_3009,N_3010);
or U3549 (N_3549,N_3245,N_3399);
xor U3550 (N_3550,N_3099,N_3295);
or U3551 (N_3551,N_3269,N_3045);
and U3552 (N_3552,N_3406,N_3436);
and U3553 (N_3553,N_3141,N_3464);
nor U3554 (N_3554,N_3088,N_3027);
nand U3555 (N_3555,N_3316,N_3040);
xor U3556 (N_3556,N_3175,N_3152);
and U3557 (N_3557,N_3171,N_3324);
nor U3558 (N_3558,N_3270,N_3444);
nand U3559 (N_3559,N_3443,N_3475);
xor U3560 (N_3560,N_3458,N_3455);
nor U3561 (N_3561,N_3007,N_3235);
nand U3562 (N_3562,N_3390,N_3402);
and U3563 (N_3563,N_3375,N_3147);
nor U3564 (N_3564,N_3089,N_3348);
or U3565 (N_3565,N_3124,N_3418);
nand U3566 (N_3566,N_3222,N_3041);
and U3567 (N_3567,N_3153,N_3005);
or U3568 (N_3568,N_3112,N_3284);
nor U3569 (N_3569,N_3302,N_3215);
xnor U3570 (N_3570,N_3042,N_3071);
or U3571 (N_3571,N_3179,N_3414);
xor U3572 (N_3572,N_3329,N_3203);
and U3573 (N_3573,N_3318,N_3218);
nand U3574 (N_3574,N_3158,N_3366);
nand U3575 (N_3575,N_3176,N_3038);
nand U3576 (N_3576,N_3427,N_3223);
nand U3577 (N_3577,N_3014,N_3363);
or U3578 (N_3578,N_3100,N_3300);
nor U3579 (N_3579,N_3065,N_3116);
or U3580 (N_3580,N_3320,N_3069);
nand U3581 (N_3581,N_3473,N_3015);
and U3582 (N_3582,N_3165,N_3022);
and U3583 (N_3583,N_3020,N_3354);
nor U3584 (N_3584,N_3368,N_3252);
nor U3585 (N_3585,N_3067,N_3396);
and U3586 (N_3586,N_3251,N_3257);
xnor U3587 (N_3587,N_3453,N_3123);
nand U3588 (N_3588,N_3199,N_3491);
and U3589 (N_3589,N_3212,N_3357);
nand U3590 (N_3590,N_3439,N_3481);
xnor U3591 (N_3591,N_3476,N_3161);
and U3592 (N_3592,N_3238,N_3328);
and U3593 (N_3593,N_3169,N_3285);
nor U3594 (N_3594,N_3194,N_3201);
and U3595 (N_3595,N_3400,N_3030);
nor U3596 (N_3596,N_3226,N_3113);
or U3597 (N_3597,N_3039,N_3466);
nor U3598 (N_3598,N_3118,N_3084);
nor U3599 (N_3599,N_3351,N_3377);
nor U3600 (N_3600,N_3205,N_3177);
xor U3601 (N_3601,N_3186,N_3170);
xor U3602 (N_3602,N_3046,N_3191);
xor U3603 (N_3603,N_3125,N_3435);
or U3604 (N_3604,N_3208,N_3085);
xnor U3605 (N_3605,N_3379,N_3266);
or U3606 (N_3606,N_3401,N_3114);
and U3607 (N_3607,N_3268,N_3095);
or U3608 (N_3608,N_3342,N_3430);
and U3609 (N_3609,N_3492,N_3425);
nor U3610 (N_3610,N_3281,N_3282);
xor U3611 (N_3611,N_3144,N_3415);
and U3612 (N_3612,N_3193,N_3217);
nand U3613 (N_3613,N_3146,N_3160);
nand U3614 (N_3614,N_3248,N_3280);
nand U3615 (N_3615,N_3164,N_3331);
and U3616 (N_3616,N_3301,N_3011);
xor U3617 (N_3617,N_3360,N_3076);
nor U3618 (N_3618,N_3241,N_3367);
nor U3619 (N_3619,N_3312,N_3323);
nor U3620 (N_3620,N_3353,N_3178);
xnor U3621 (N_3621,N_3192,N_3111);
and U3622 (N_3622,N_3134,N_3438);
and U3623 (N_3623,N_3265,N_3424);
and U3624 (N_3624,N_3447,N_3371);
nand U3625 (N_3625,N_3240,N_3024);
or U3626 (N_3626,N_3068,N_3279);
and U3627 (N_3627,N_3063,N_3330);
nand U3628 (N_3628,N_3143,N_3023);
xnor U3629 (N_3629,N_3322,N_3431);
xor U3630 (N_3630,N_3446,N_3332);
or U3631 (N_3631,N_3168,N_3132);
xnor U3632 (N_3632,N_3493,N_3304);
nor U3633 (N_3633,N_3423,N_3083);
xor U3634 (N_3634,N_3259,N_3461);
nand U3635 (N_3635,N_3066,N_3350);
nand U3636 (N_3636,N_3278,N_3352);
nand U3637 (N_3637,N_3130,N_3033);
and U3638 (N_3638,N_3232,N_3140);
and U3639 (N_3639,N_3277,N_3333);
nand U3640 (N_3640,N_3092,N_3059);
nand U3641 (N_3641,N_3263,N_3489);
xnor U3642 (N_3642,N_3373,N_3119);
or U3643 (N_3643,N_3110,N_3482);
nor U3644 (N_3644,N_3093,N_3128);
nor U3645 (N_3645,N_3485,N_3097);
or U3646 (N_3646,N_3082,N_3254);
or U3647 (N_3647,N_3197,N_3224);
xnor U3648 (N_3648,N_3389,N_3211);
nor U3649 (N_3649,N_3397,N_3016);
xor U3650 (N_3650,N_3306,N_3006);
nand U3651 (N_3651,N_3432,N_3173);
nand U3652 (N_3652,N_3345,N_3384);
xnor U3653 (N_3653,N_3196,N_3388);
or U3654 (N_3654,N_3347,N_3086);
or U3655 (N_3655,N_3487,N_3376);
or U3656 (N_3656,N_3391,N_3058);
and U3657 (N_3657,N_3472,N_3394);
or U3658 (N_3658,N_3250,N_3463);
nand U3659 (N_3659,N_3405,N_3221);
and U3660 (N_3660,N_3019,N_3370);
xnor U3661 (N_3661,N_3209,N_3129);
xor U3662 (N_3662,N_3336,N_3072);
and U3663 (N_3663,N_3115,N_3050);
nand U3664 (N_3664,N_3404,N_3230);
nor U3665 (N_3665,N_3122,N_3273);
and U3666 (N_3666,N_3035,N_3393);
or U3667 (N_3667,N_3183,N_3207);
nand U3668 (N_3668,N_3229,N_3337);
nand U3669 (N_3669,N_3159,N_3362);
or U3670 (N_3670,N_3441,N_3471);
xnor U3671 (N_3671,N_3299,N_3296);
nor U3672 (N_3672,N_3075,N_3417);
nand U3673 (N_3673,N_3395,N_3325);
nor U3674 (N_3674,N_3339,N_3061);
nand U3675 (N_3675,N_3150,N_3013);
xnor U3676 (N_3676,N_3261,N_3074);
and U3677 (N_3677,N_3102,N_3091);
xor U3678 (N_3678,N_3062,N_3303);
nand U3679 (N_3679,N_3460,N_3498);
and U3680 (N_3680,N_3139,N_3204);
and U3681 (N_3681,N_3137,N_3054);
and U3682 (N_3682,N_3162,N_3073);
nor U3683 (N_3683,N_3450,N_3349);
and U3684 (N_3684,N_3256,N_3145);
and U3685 (N_3685,N_3154,N_3308);
xnor U3686 (N_3686,N_3452,N_3195);
nor U3687 (N_3687,N_3172,N_3334);
nand U3688 (N_3688,N_3483,N_3180);
and U3689 (N_3689,N_3293,N_3364);
nor U3690 (N_3690,N_3214,N_3142);
nand U3691 (N_3691,N_3480,N_3309);
nor U3692 (N_3692,N_3289,N_3341);
or U3693 (N_3693,N_3060,N_3478);
or U3694 (N_3694,N_3381,N_3190);
xor U3695 (N_3695,N_3412,N_3421);
xnor U3696 (N_3696,N_3021,N_3198);
nor U3697 (N_3697,N_3344,N_3077);
xor U3698 (N_3698,N_3271,N_3321);
and U3699 (N_3699,N_3003,N_3167);
and U3700 (N_3700,N_3413,N_3338);
nor U3701 (N_3701,N_3361,N_3385);
and U3702 (N_3702,N_3294,N_3276);
nand U3703 (N_3703,N_3290,N_3382);
or U3704 (N_3704,N_3200,N_3008);
nand U3705 (N_3705,N_3233,N_3457);
or U3706 (N_3706,N_3267,N_3036);
or U3707 (N_3707,N_3080,N_3055);
nand U3708 (N_3708,N_3462,N_3001);
or U3709 (N_3709,N_3127,N_3380);
nand U3710 (N_3710,N_3307,N_3121);
and U3711 (N_3711,N_3378,N_3420);
or U3712 (N_3712,N_3264,N_3497);
and U3713 (N_3713,N_3188,N_3416);
xnor U3714 (N_3714,N_3049,N_3181);
xnor U3715 (N_3715,N_3407,N_3428);
xor U3716 (N_3716,N_3469,N_3070);
nand U3717 (N_3717,N_3410,N_3002);
and U3718 (N_3718,N_3103,N_3258);
or U3719 (N_3719,N_3474,N_3012);
xor U3720 (N_3720,N_3494,N_3109);
and U3721 (N_3721,N_3120,N_3155);
or U3722 (N_3722,N_3496,N_3228);
nor U3723 (N_3723,N_3355,N_3346);
nand U3724 (N_3724,N_3359,N_3343);
and U3725 (N_3725,N_3126,N_3107);
nand U3726 (N_3726,N_3488,N_3311);
or U3727 (N_3727,N_3096,N_3043);
or U3728 (N_3728,N_3409,N_3253);
nand U3729 (N_3729,N_3206,N_3484);
and U3730 (N_3730,N_3029,N_3326);
or U3731 (N_3731,N_3272,N_3090);
nor U3732 (N_3732,N_3234,N_3448);
nand U3733 (N_3733,N_3026,N_3249);
and U3734 (N_3734,N_3477,N_3408);
and U3735 (N_3735,N_3202,N_3106);
or U3736 (N_3736,N_3187,N_3220);
or U3737 (N_3737,N_3032,N_3411);
nor U3738 (N_3738,N_3255,N_3182);
and U3739 (N_3739,N_3057,N_3454);
nand U3740 (N_3740,N_3287,N_3422);
and U3741 (N_3741,N_3048,N_3213);
and U3742 (N_3742,N_3314,N_3292);
or U3743 (N_3743,N_3037,N_3358);
nor U3744 (N_3744,N_3163,N_3470);
nand U3745 (N_3745,N_3138,N_3184);
nand U3746 (N_3746,N_3174,N_3398);
and U3747 (N_3747,N_3449,N_3275);
xnor U3748 (N_3748,N_3064,N_3374);
and U3749 (N_3749,N_3239,N_3317);
or U3750 (N_3750,N_3244,N_3041);
and U3751 (N_3751,N_3464,N_3126);
nand U3752 (N_3752,N_3478,N_3280);
nor U3753 (N_3753,N_3229,N_3175);
and U3754 (N_3754,N_3417,N_3390);
nand U3755 (N_3755,N_3205,N_3087);
and U3756 (N_3756,N_3389,N_3349);
and U3757 (N_3757,N_3181,N_3433);
nor U3758 (N_3758,N_3396,N_3344);
nand U3759 (N_3759,N_3255,N_3370);
and U3760 (N_3760,N_3427,N_3360);
nand U3761 (N_3761,N_3215,N_3220);
or U3762 (N_3762,N_3038,N_3408);
nand U3763 (N_3763,N_3017,N_3076);
nand U3764 (N_3764,N_3182,N_3273);
xnor U3765 (N_3765,N_3350,N_3121);
nor U3766 (N_3766,N_3288,N_3359);
and U3767 (N_3767,N_3044,N_3039);
and U3768 (N_3768,N_3423,N_3081);
or U3769 (N_3769,N_3308,N_3108);
or U3770 (N_3770,N_3314,N_3336);
nor U3771 (N_3771,N_3373,N_3191);
nand U3772 (N_3772,N_3379,N_3374);
nand U3773 (N_3773,N_3134,N_3201);
nor U3774 (N_3774,N_3067,N_3430);
and U3775 (N_3775,N_3468,N_3397);
xor U3776 (N_3776,N_3493,N_3163);
or U3777 (N_3777,N_3184,N_3353);
and U3778 (N_3778,N_3310,N_3011);
or U3779 (N_3779,N_3099,N_3186);
and U3780 (N_3780,N_3354,N_3456);
nor U3781 (N_3781,N_3296,N_3083);
and U3782 (N_3782,N_3212,N_3057);
xor U3783 (N_3783,N_3151,N_3344);
nand U3784 (N_3784,N_3089,N_3065);
xor U3785 (N_3785,N_3047,N_3073);
nor U3786 (N_3786,N_3305,N_3301);
or U3787 (N_3787,N_3214,N_3212);
xnor U3788 (N_3788,N_3373,N_3282);
or U3789 (N_3789,N_3139,N_3335);
nor U3790 (N_3790,N_3164,N_3219);
nand U3791 (N_3791,N_3281,N_3338);
or U3792 (N_3792,N_3430,N_3167);
and U3793 (N_3793,N_3018,N_3033);
nand U3794 (N_3794,N_3036,N_3357);
or U3795 (N_3795,N_3089,N_3048);
nor U3796 (N_3796,N_3395,N_3476);
or U3797 (N_3797,N_3042,N_3185);
nor U3798 (N_3798,N_3272,N_3080);
xnor U3799 (N_3799,N_3454,N_3026);
and U3800 (N_3800,N_3292,N_3347);
xnor U3801 (N_3801,N_3217,N_3268);
or U3802 (N_3802,N_3147,N_3331);
or U3803 (N_3803,N_3257,N_3282);
nor U3804 (N_3804,N_3003,N_3114);
and U3805 (N_3805,N_3133,N_3110);
and U3806 (N_3806,N_3479,N_3192);
and U3807 (N_3807,N_3194,N_3039);
or U3808 (N_3808,N_3164,N_3206);
xor U3809 (N_3809,N_3058,N_3394);
nor U3810 (N_3810,N_3350,N_3272);
or U3811 (N_3811,N_3245,N_3296);
and U3812 (N_3812,N_3466,N_3315);
nand U3813 (N_3813,N_3124,N_3338);
nor U3814 (N_3814,N_3390,N_3055);
nand U3815 (N_3815,N_3338,N_3248);
nor U3816 (N_3816,N_3063,N_3424);
xor U3817 (N_3817,N_3188,N_3303);
and U3818 (N_3818,N_3091,N_3131);
nand U3819 (N_3819,N_3109,N_3103);
and U3820 (N_3820,N_3168,N_3217);
xnor U3821 (N_3821,N_3048,N_3252);
xor U3822 (N_3822,N_3403,N_3186);
nor U3823 (N_3823,N_3461,N_3400);
nor U3824 (N_3824,N_3198,N_3108);
nand U3825 (N_3825,N_3275,N_3481);
nor U3826 (N_3826,N_3291,N_3411);
nor U3827 (N_3827,N_3033,N_3021);
xnor U3828 (N_3828,N_3168,N_3170);
and U3829 (N_3829,N_3044,N_3189);
nand U3830 (N_3830,N_3353,N_3430);
and U3831 (N_3831,N_3080,N_3001);
nor U3832 (N_3832,N_3224,N_3225);
and U3833 (N_3833,N_3484,N_3410);
xor U3834 (N_3834,N_3023,N_3484);
nand U3835 (N_3835,N_3307,N_3365);
nor U3836 (N_3836,N_3261,N_3302);
or U3837 (N_3837,N_3432,N_3370);
or U3838 (N_3838,N_3152,N_3174);
xnor U3839 (N_3839,N_3441,N_3496);
xnor U3840 (N_3840,N_3376,N_3192);
nor U3841 (N_3841,N_3290,N_3210);
nand U3842 (N_3842,N_3079,N_3089);
xnor U3843 (N_3843,N_3169,N_3405);
nor U3844 (N_3844,N_3177,N_3086);
nand U3845 (N_3845,N_3314,N_3006);
xor U3846 (N_3846,N_3493,N_3143);
nand U3847 (N_3847,N_3271,N_3403);
and U3848 (N_3848,N_3121,N_3066);
nand U3849 (N_3849,N_3203,N_3082);
xor U3850 (N_3850,N_3041,N_3206);
xor U3851 (N_3851,N_3222,N_3306);
nand U3852 (N_3852,N_3105,N_3478);
nor U3853 (N_3853,N_3347,N_3144);
nand U3854 (N_3854,N_3271,N_3280);
nand U3855 (N_3855,N_3271,N_3430);
nand U3856 (N_3856,N_3099,N_3471);
nand U3857 (N_3857,N_3166,N_3039);
or U3858 (N_3858,N_3269,N_3117);
and U3859 (N_3859,N_3246,N_3272);
nor U3860 (N_3860,N_3318,N_3451);
xor U3861 (N_3861,N_3459,N_3489);
and U3862 (N_3862,N_3077,N_3341);
or U3863 (N_3863,N_3464,N_3051);
and U3864 (N_3864,N_3113,N_3439);
nor U3865 (N_3865,N_3074,N_3183);
nor U3866 (N_3866,N_3132,N_3309);
nand U3867 (N_3867,N_3373,N_3367);
or U3868 (N_3868,N_3437,N_3335);
nor U3869 (N_3869,N_3305,N_3449);
or U3870 (N_3870,N_3184,N_3095);
nor U3871 (N_3871,N_3135,N_3133);
xnor U3872 (N_3872,N_3051,N_3200);
nand U3873 (N_3873,N_3472,N_3156);
xnor U3874 (N_3874,N_3243,N_3007);
or U3875 (N_3875,N_3090,N_3391);
or U3876 (N_3876,N_3283,N_3476);
nand U3877 (N_3877,N_3374,N_3089);
and U3878 (N_3878,N_3339,N_3294);
nand U3879 (N_3879,N_3170,N_3036);
and U3880 (N_3880,N_3363,N_3101);
and U3881 (N_3881,N_3157,N_3119);
nor U3882 (N_3882,N_3090,N_3498);
nand U3883 (N_3883,N_3166,N_3448);
or U3884 (N_3884,N_3296,N_3332);
or U3885 (N_3885,N_3033,N_3040);
and U3886 (N_3886,N_3069,N_3259);
xor U3887 (N_3887,N_3130,N_3022);
xnor U3888 (N_3888,N_3127,N_3023);
nor U3889 (N_3889,N_3431,N_3137);
xor U3890 (N_3890,N_3183,N_3278);
and U3891 (N_3891,N_3052,N_3205);
nor U3892 (N_3892,N_3368,N_3412);
xnor U3893 (N_3893,N_3288,N_3405);
nand U3894 (N_3894,N_3472,N_3272);
or U3895 (N_3895,N_3388,N_3444);
or U3896 (N_3896,N_3008,N_3326);
nor U3897 (N_3897,N_3135,N_3243);
xnor U3898 (N_3898,N_3141,N_3495);
and U3899 (N_3899,N_3076,N_3083);
and U3900 (N_3900,N_3131,N_3453);
or U3901 (N_3901,N_3251,N_3181);
xor U3902 (N_3902,N_3099,N_3134);
nand U3903 (N_3903,N_3113,N_3340);
or U3904 (N_3904,N_3077,N_3420);
nand U3905 (N_3905,N_3172,N_3268);
and U3906 (N_3906,N_3043,N_3464);
or U3907 (N_3907,N_3080,N_3374);
nor U3908 (N_3908,N_3318,N_3276);
nor U3909 (N_3909,N_3096,N_3049);
xnor U3910 (N_3910,N_3303,N_3202);
xnor U3911 (N_3911,N_3106,N_3381);
nand U3912 (N_3912,N_3062,N_3480);
xnor U3913 (N_3913,N_3205,N_3328);
and U3914 (N_3914,N_3318,N_3022);
xnor U3915 (N_3915,N_3241,N_3116);
and U3916 (N_3916,N_3406,N_3041);
and U3917 (N_3917,N_3061,N_3013);
and U3918 (N_3918,N_3176,N_3194);
and U3919 (N_3919,N_3471,N_3465);
or U3920 (N_3920,N_3344,N_3204);
nand U3921 (N_3921,N_3042,N_3432);
or U3922 (N_3922,N_3060,N_3375);
xnor U3923 (N_3923,N_3318,N_3235);
nand U3924 (N_3924,N_3164,N_3318);
xor U3925 (N_3925,N_3384,N_3307);
nor U3926 (N_3926,N_3086,N_3451);
nand U3927 (N_3927,N_3417,N_3096);
xor U3928 (N_3928,N_3239,N_3257);
nor U3929 (N_3929,N_3059,N_3490);
and U3930 (N_3930,N_3300,N_3231);
or U3931 (N_3931,N_3432,N_3100);
xor U3932 (N_3932,N_3401,N_3202);
nor U3933 (N_3933,N_3333,N_3155);
nand U3934 (N_3934,N_3169,N_3095);
nand U3935 (N_3935,N_3006,N_3315);
nor U3936 (N_3936,N_3473,N_3188);
nand U3937 (N_3937,N_3229,N_3103);
nand U3938 (N_3938,N_3496,N_3016);
nand U3939 (N_3939,N_3312,N_3051);
nor U3940 (N_3940,N_3240,N_3464);
nor U3941 (N_3941,N_3435,N_3315);
nor U3942 (N_3942,N_3106,N_3326);
xnor U3943 (N_3943,N_3451,N_3404);
or U3944 (N_3944,N_3307,N_3478);
xor U3945 (N_3945,N_3407,N_3236);
and U3946 (N_3946,N_3155,N_3475);
and U3947 (N_3947,N_3032,N_3466);
nor U3948 (N_3948,N_3155,N_3121);
and U3949 (N_3949,N_3426,N_3323);
xnor U3950 (N_3950,N_3117,N_3136);
nor U3951 (N_3951,N_3433,N_3078);
nand U3952 (N_3952,N_3371,N_3345);
and U3953 (N_3953,N_3028,N_3320);
nor U3954 (N_3954,N_3309,N_3024);
and U3955 (N_3955,N_3137,N_3369);
nor U3956 (N_3956,N_3167,N_3397);
nor U3957 (N_3957,N_3341,N_3431);
nand U3958 (N_3958,N_3059,N_3079);
and U3959 (N_3959,N_3307,N_3236);
nand U3960 (N_3960,N_3218,N_3245);
or U3961 (N_3961,N_3300,N_3298);
nor U3962 (N_3962,N_3100,N_3222);
xnor U3963 (N_3963,N_3488,N_3107);
and U3964 (N_3964,N_3413,N_3369);
nor U3965 (N_3965,N_3245,N_3435);
nor U3966 (N_3966,N_3431,N_3127);
nor U3967 (N_3967,N_3312,N_3215);
nor U3968 (N_3968,N_3229,N_3299);
nor U3969 (N_3969,N_3148,N_3313);
nand U3970 (N_3970,N_3064,N_3442);
or U3971 (N_3971,N_3345,N_3258);
and U3972 (N_3972,N_3063,N_3392);
nand U3973 (N_3973,N_3110,N_3068);
xnor U3974 (N_3974,N_3333,N_3486);
or U3975 (N_3975,N_3380,N_3360);
nor U3976 (N_3976,N_3475,N_3409);
nand U3977 (N_3977,N_3014,N_3296);
nor U3978 (N_3978,N_3097,N_3077);
xnor U3979 (N_3979,N_3118,N_3354);
or U3980 (N_3980,N_3385,N_3422);
nor U3981 (N_3981,N_3167,N_3168);
and U3982 (N_3982,N_3064,N_3194);
nand U3983 (N_3983,N_3348,N_3314);
nand U3984 (N_3984,N_3447,N_3298);
nand U3985 (N_3985,N_3127,N_3354);
nand U3986 (N_3986,N_3151,N_3142);
xor U3987 (N_3987,N_3054,N_3025);
nor U3988 (N_3988,N_3116,N_3259);
nor U3989 (N_3989,N_3309,N_3239);
nor U3990 (N_3990,N_3081,N_3397);
and U3991 (N_3991,N_3329,N_3489);
nor U3992 (N_3992,N_3079,N_3034);
xor U3993 (N_3993,N_3322,N_3267);
xnor U3994 (N_3994,N_3376,N_3068);
nand U3995 (N_3995,N_3336,N_3460);
xor U3996 (N_3996,N_3292,N_3146);
xnor U3997 (N_3997,N_3170,N_3470);
xnor U3998 (N_3998,N_3264,N_3009);
nor U3999 (N_3999,N_3022,N_3355);
nand U4000 (N_4000,N_3778,N_3594);
or U4001 (N_4001,N_3549,N_3983);
or U4002 (N_4002,N_3690,N_3502);
xnor U4003 (N_4003,N_3981,N_3923);
nand U4004 (N_4004,N_3819,N_3897);
nor U4005 (N_4005,N_3913,N_3921);
nand U4006 (N_4006,N_3583,N_3917);
or U4007 (N_4007,N_3808,N_3753);
xnor U4008 (N_4008,N_3516,N_3947);
nor U4009 (N_4009,N_3810,N_3795);
or U4010 (N_4010,N_3912,N_3843);
nor U4011 (N_4011,N_3679,N_3847);
and U4012 (N_4012,N_3554,N_3946);
xor U4013 (N_4013,N_3576,N_3669);
or U4014 (N_4014,N_3855,N_3556);
nor U4015 (N_4015,N_3738,N_3850);
and U4016 (N_4016,N_3513,N_3541);
and U4017 (N_4017,N_3641,N_3900);
nor U4018 (N_4018,N_3870,N_3942);
xor U4019 (N_4019,N_3938,N_3729);
nor U4020 (N_4020,N_3857,N_3812);
xnor U4021 (N_4021,N_3998,N_3539);
or U4022 (N_4022,N_3538,N_3561);
nor U4023 (N_4023,N_3834,N_3560);
nor U4024 (N_4024,N_3929,N_3658);
and U4025 (N_4025,N_3547,N_3809);
and U4026 (N_4026,N_3905,N_3572);
nand U4027 (N_4027,N_3600,N_3545);
nand U4028 (N_4028,N_3979,N_3704);
nor U4029 (N_4029,N_3707,N_3780);
or U4030 (N_4030,N_3884,N_3699);
nand U4031 (N_4031,N_3644,N_3893);
or U4032 (N_4032,N_3828,N_3761);
xnor U4033 (N_4033,N_3649,N_3526);
nand U4034 (N_4034,N_3973,N_3933);
xor U4035 (N_4035,N_3728,N_3614);
or U4036 (N_4036,N_3646,N_3841);
nor U4037 (N_4037,N_3524,N_3694);
or U4038 (N_4038,N_3798,N_3675);
nor U4039 (N_4039,N_3967,N_3939);
nand U4040 (N_4040,N_3667,N_3747);
and U4041 (N_4041,N_3741,N_3661);
nor U4042 (N_4042,N_3501,N_3980);
and U4043 (N_4043,N_3719,N_3793);
or U4044 (N_4044,N_3889,N_3581);
or U4045 (N_4045,N_3557,N_3832);
xor U4046 (N_4046,N_3711,N_3823);
and U4047 (N_4047,N_3901,N_3678);
xor U4048 (N_4048,N_3735,N_3925);
nor U4049 (N_4049,N_3971,N_3598);
and U4050 (N_4050,N_3818,N_3910);
xor U4051 (N_4051,N_3687,N_3977);
nand U4052 (N_4052,N_3589,N_3805);
xor U4053 (N_4053,N_3908,N_3764);
xnor U4054 (N_4054,N_3505,N_3886);
xnor U4055 (N_4055,N_3584,N_3800);
or U4056 (N_4056,N_3715,N_3759);
nand U4057 (N_4057,N_3708,N_3858);
or U4058 (N_4058,N_3882,N_3914);
or U4059 (N_4059,N_3571,N_3776);
and U4060 (N_4060,N_3622,N_3978);
nand U4061 (N_4061,N_3628,N_3582);
xnor U4062 (N_4062,N_3794,N_3639);
nor U4063 (N_4063,N_3559,N_3875);
and U4064 (N_4064,N_3540,N_3573);
nand U4065 (N_4065,N_3535,N_3878);
xor U4066 (N_4066,N_3617,N_3602);
and U4067 (N_4067,N_3999,N_3907);
nor U4068 (N_4068,N_3955,N_3743);
nand U4069 (N_4069,N_3763,N_3960);
xor U4070 (N_4070,N_3500,N_3948);
nand U4071 (N_4071,N_3902,N_3846);
nand U4072 (N_4072,N_3799,N_3990);
and U4073 (N_4073,N_3997,N_3773);
or U4074 (N_4074,N_3896,N_3625);
nor U4075 (N_4075,N_3922,N_3777);
or U4076 (N_4076,N_3888,N_3721);
and U4077 (N_4077,N_3710,N_3944);
and U4078 (N_4078,N_3883,N_3957);
nand U4079 (N_4079,N_3636,N_3749);
and U4080 (N_4080,N_3592,N_3564);
or U4081 (N_4081,N_3926,N_3558);
xnor U4082 (N_4082,N_3987,N_3631);
and U4083 (N_4083,N_3781,N_3731);
xor U4084 (N_4084,N_3839,N_3697);
xnor U4085 (N_4085,N_3612,N_3624);
and U4086 (N_4086,N_3989,N_3924);
nand U4087 (N_4087,N_3531,N_3804);
and U4088 (N_4088,N_3705,N_3525);
and U4089 (N_4089,N_3919,N_3765);
nor U4090 (N_4090,N_3730,N_3873);
or U4091 (N_4091,N_3899,N_3542);
or U4092 (N_4092,N_3567,N_3643);
nand U4093 (N_4093,N_3941,N_3827);
or U4094 (N_4094,N_3634,N_3806);
nand U4095 (N_4095,N_3797,N_3609);
xor U4096 (N_4096,N_3654,N_3666);
xnor U4097 (N_4097,N_3943,N_3618);
and U4098 (N_4098,N_3685,N_3537);
nor U4099 (N_4099,N_3740,N_3551);
nor U4100 (N_4100,N_3783,N_3637);
xnor U4101 (N_4101,N_3752,N_3648);
or U4102 (N_4102,N_3803,N_3934);
or U4103 (N_4103,N_3845,N_3726);
and U4104 (N_4104,N_3503,N_3891);
nand U4105 (N_4105,N_3782,N_3959);
xnor U4106 (N_4106,N_3853,N_3595);
nand U4107 (N_4107,N_3758,N_3991);
nand U4108 (N_4108,N_3536,N_3826);
nor U4109 (N_4109,N_3930,N_3709);
nor U4110 (N_4110,N_3528,N_3664);
nor U4111 (N_4111,N_3651,N_3771);
and U4112 (N_4112,N_3543,N_3652);
xnor U4113 (N_4113,N_3993,N_3577);
nor U4114 (N_4114,N_3848,N_3779);
or U4115 (N_4115,N_3769,N_3824);
and U4116 (N_4116,N_3831,N_3518);
xnor U4117 (N_4117,N_3898,N_3623);
xnor U4118 (N_4118,N_3787,N_3670);
nor U4119 (N_4119,N_3746,N_3613);
nand U4120 (N_4120,N_3890,N_3723);
or U4121 (N_4121,N_3750,N_3653);
or U4122 (N_4122,N_3995,N_3916);
and U4123 (N_4123,N_3885,N_3548);
nor U4124 (N_4124,N_3701,N_3963);
and U4125 (N_4125,N_3876,N_3590);
or U4126 (N_4126,N_3785,N_3727);
nor U4127 (N_4127,N_3868,N_3504);
or U4128 (N_4128,N_3837,N_3932);
nand U4129 (N_4129,N_3951,N_3881);
nand U4130 (N_4130,N_3520,N_3970);
nor U4131 (N_4131,N_3838,N_3903);
xor U4132 (N_4132,N_3877,N_3574);
nor U4133 (N_4133,N_3615,N_3863);
nor U4134 (N_4134,N_3736,N_3770);
and U4135 (N_4135,N_3596,N_3610);
nor U4136 (N_4136,N_3660,N_3680);
nand U4137 (N_4137,N_3587,N_3620);
or U4138 (N_4138,N_3673,N_3994);
and U4139 (N_4139,N_3533,N_3969);
nor U4140 (N_4140,N_3755,N_3645);
xnor U4141 (N_4141,N_3760,N_3691);
and U4142 (N_4142,N_3920,N_3861);
xor U4143 (N_4143,N_3936,N_3703);
nor U4144 (N_4144,N_3786,N_3801);
nor U4145 (N_4145,N_3796,N_3717);
or U4146 (N_4146,N_3742,N_3608);
nand U4147 (N_4147,N_3909,N_3956);
nand U4148 (N_4148,N_3714,N_3976);
or U4149 (N_4149,N_3689,N_3580);
nor U4150 (N_4150,N_3553,N_3972);
and U4151 (N_4151,N_3880,N_3966);
nor U4152 (N_4152,N_3734,N_3964);
or U4153 (N_4153,N_3968,N_3836);
nand U4154 (N_4154,N_3864,N_3874);
and U4155 (N_4155,N_3950,N_3522);
or U4156 (N_4156,N_3725,N_3958);
and U4157 (N_4157,N_3546,N_3511);
nand U4158 (N_4158,N_3982,N_3720);
nor U4159 (N_4159,N_3816,N_3811);
xnor U4160 (N_4160,N_3862,N_3974);
or U4161 (N_4161,N_3892,N_3737);
xor U4162 (N_4162,N_3601,N_3702);
nand U4163 (N_4163,N_3928,N_3813);
nor U4164 (N_4164,N_3854,N_3568);
or U4165 (N_4165,N_3512,N_3683);
nand U4166 (N_4166,N_3599,N_3565);
nand U4167 (N_4167,N_3869,N_3851);
nand U4168 (N_4168,N_3510,N_3790);
or U4169 (N_4169,N_3681,N_3593);
xor U4170 (N_4170,N_3650,N_3616);
and U4171 (N_4171,N_3586,N_3867);
or U4172 (N_4172,N_3591,N_3784);
nor U4173 (N_4173,N_3521,N_3918);
xnor U4174 (N_4174,N_3856,N_3911);
nand U4175 (N_4175,N_3835,N_3684);
nor U4176 (N_4176,N_3775,N_3751);
or U4177 (N_4177,N_3544,N_3509);
nor U4178 (N_4178,N_3605,N_3692);
xnor U4179 (N_4179,N_3927,N_3904);
nor U4180 (N_4180,N_3633,N_3527);
and U4181 (N_4181,N_3830,N_3579);
xor U4182 (N_4182,N_3887,N_3671);
nor U4183 (N_4183,N_3603,N_3865);
or U4184 (N_4184,N_3791,N_3829);
and U4185 (N_4185,N_3988,N_3852);
nor U4186 (N_4186,N_3849,N_3820);
and U4187 (N_4187,N_3588,N_3844);
xnor U4188 (N_4188,N_3517,N_3663);
xor U4189 (N_4189,N_3662,N_3514);
nor U4190 (N_4190,N_3570,N_3712);
xnor U4191 (N_4191,N_3986,N_3996);
xnor U4192 (N_4192,N_3745,N_3682);
nor U4193 (N_4193,N_3984,N_3985);
nand U4194 (N_4194,N_3621,N_3647);
xnor U4195 (N_4195,N_3744,N_3693);
and U4196 (N_4196,N_3945,N_3722);
and U4197 (N_4197,N_3965,N_3935);
nand U4198 (N_4198,N_3706,N_3508);
nor U4199 (N_4199,N_3552,N_3724);
xor U4200 (N_4200,N_3562,N_3802);
nand U4201 (N_4201,N_3550,N_3774);
or U4202 (N_4202,N_3638,N_3688);
nand U4203 (N_4203,N_3627,N_3871);
xor U4204 (N_4204,N_3506,N_3676);
nand U4205 (N_4205,N_3733,N_3677);
xnor U4206 (N_4206,N_3629,N_3519);
or U4207 (N_4207,N_3906,N_3772);
or U4208 (N_4208,N_3949,N_3672);
and U4209 (N_4209,N_3700,N_3767);
xor U4210 (N_4210,N_3515,N_3732);
and U4211 (N_4211,N_3665,N_3768);
nand U4212 (N_4212,N_3630,N_3842);
or U4213 (N_4213,N_3659,N_3597);
xor U4214 (N_4214,N_3756,N_3815);
nor U4215 (N_4215,N_3825,N_3894);
and U4216 (N_4216,N_3530,N_3833);
and U4217 (N_4217,N_3569,N_3817);
and U4218 (N_4218,N_3762,N_3686);
and U4219 (N_4219,N_3563,N_3961);
nor U4220 (N_4220,N_3859,N_3895);
xnor U4221 (N_4221,N_3822,N_3792);
nand U4222 (N_4222,N_3695,N_3789);
nand U4223 (N_4223,N_3534,N_3642);
nand U4224 (N_4224,N_3814,N_3915);
nor U4225 (N_4225,N_3529,N_3716);
or U4226 (N_4226,N_3674,N_3655);
xor U4227 (N_4227,N_3640,N_3788);
xor U4228 (N_4228,N_3931,N_3606);
xnor U4229 (N_4229,N_3748,N_3635);
or U4230 (N_4230,N_3879,N_3992);
and U4231 (N_4231,N_3754,N_3668);
nand U4232 (N_4232,N_3807,N_3566);
and U4233 (N_4233,N_3698,N_3507);
xor U4234 (N_4234,N_3611,N_3954);
or U4235 (N_4235,N_3975,N_3607);
xnor U4236 (N_4236,N_3696,N_3555);
or U4237 (N_4237,N_3860,N_3766);
xnor U4238 (N_4238,N_3866,N_3619);
nand U4239 (N_4239,N_3739,N_3713);
and U4240 (N_4240,N_3575,N_3656);
or U4241 (N_4241,N_3840,N_3532);
xor U4242 (N_4242,N_3952,N_3872);
nor U4243 (N_4243,N_3604,N_3962);
nand U4244 (N_4244,N_3585,N_3657);
nor U4245 (N_4245,N_3821,N_3626);
nand U4246 (N_4246,N_3523,N_3937);
nand U4247 (N_4247,N_3718,N_3632);
nor U4248 (N_4248,N_3953,N_3757);
nor U4249 (N_4249,N_3578,N_3940);
or U4250 (N_4250,N_3511,N_3640);
xnor U4251 (N_4251,N_3680,N_3681);
nand U4252 (N_4252,N_3763,N_3559);
nor U4253 (N_4253,N_3676,N_3775);
nand U4254 (N_4254,N_3821,N_3779);
nand U4255 (N_4255,N_3781,N_3522);
nor U4256 (N_4256,N_3692,N_3932);
nor U4257 (N_4257,N_3666,N_3790);
or U4258 (N_4258,N_3797,N_3971);
and U4259 (N_4259,N_3961,N_3801);
xnor U4260 (N_4260,N_3903,N_3779);
or U4261 (N_4261,N_3691,N_3960);
or U4262 (N_4262,N_3500,N_3837);
nand U4263 (N_4263,N_3533,N_3677);
xor U4264 (N_4264,N_3749,N_3909);
nand U4265 (N_4265,N_3581,N_3828);
nand U4266 (N_4266,N_3506,N_3637);
or U4267 (N_4267,N_3728,N_3955);
or U4268 (N_4268,N_3644,N_3764);
xor U4269 (N_4269,N_3984,N_3596);
and U4270 (N_4270,N_3689,N_3844);
or U4271 (N_4271,N_3758,N_3894);
nand U4272 (N_4272,N_3673,N_3894);
and U4273 (N_4273,N_3945,N_3728);
and U4274 (N_4274,N_3929,N_3824);
nand U4275 (N_4275,N_3558,N_3713);
nand U4276 (N_4276,N_3678,N_3677);
nand U4277 (N_4277,N_3795,N_3837);
nor U4278 (N_4278,N_3631,N_3971);
nor U4279 (N_4279,N_3995,N_3643);
and U4280 (N_4280,N_3773,N_3865);
xnor U4281 (N_4281,N_3580,N_3881);
xor U4282 (N_4282,N_3633,N_3703);
and U4283 (N_4283,N_3661,N_3871);
nor U4284 (N_4284,N_3684,N_3713);
or U4285 (N_4285,N_3539,N_3690);
nand U4286 (N_4286,N_3819,N_3749);
nor U4287 (N_4287,N_3802,N_3756);
nand U4288 (N_4288,N_3584,N_3631);
nor U4289 (N_4289,N_3581,N_3561);
nor U4290 (N_4290,N_3835,N_3918);
and U4291 (N_4291,N_3619,N_3973);
nand U4292 (N_4292,N_3527,N_3718);
nand U4293 (N_4293,N_3965,N_3602);
nor U4294 (N_4294,N_3806,N_3510);
nor U4295 (N_4295,N_3572,N_3993);
xor U4296 (N_4296,N_3688,N_3861);
xor U4297 (N_4297,N_3786,N_3959);
nand U4298 (N_4298,N_3606,N_3856);
xor U4299 (N_4299,N_3751,N_3901);
and U4300 (N_4300,N_3576,N_3675);
and U4301 (N_4301,N_3735,N_3890);
xor U4302 (N_4302,N_3640,N_3683);
xnor U4303 (N_4303,N_3861,N_3633);
nand U4304 (N_4304,N_3644,N_3836);
xor U4305 (N_4305,N_3939,N_3998);
and U4306 (N_4306,N_3603,N_3626);
nor U4307 (N_4307,N_3983,N_3607);
nor U4308 (N_4308,N_3637,N_3702);
nor U4309 (N_4309,N_3984,N_3986);
nor U4310 (N_4310,N_3888,N_3549);
xnor U4311 (N_4311,N_3826,N_3582);
and U4312 (N_4312,N_3778,N_3512);
nand U4313 (N_4313,N_3805,N_3835);
and U4314 (N_4314,N_3830,N_3628);
xor U4315 (N_4315,N_3775,N_3666);
xnor U4316 (N_4316,N_3884,N_3757);
and U4317 (N_4317,N_3893,N_3512);
xnor U4318 (N_4318,N_3886,N_3879);
nand U4319 (N_4319,N_3590,N_3834);
nor U4320 (N_4320,N_3770,N_3603);
nand U4321 (N_4321,N_3881,N_3945);
and U4322 (N_4322,N_3899,N_3513);
nor U4323 (N_4323,N_3721,N_3930);
xnor U4324 (N_4324,N_3509,N_3928);
nor U4325 (N_4325,N_3858,N_3592);
and U4326 (N_4326,N_3545,N_3573);
nor U4327 (N_4327,N_3780,N_3667);
or U4328 (N_4328,N_3772,N_3940);
nand U4329 (N_4329,N_3719,N_3992);
nand U4330 (N_4330,N_3693,N_3827);
nand U4331 (N_4331,N_3764,N_3993);
and U4332 (N_4332,N_3541,N_3596);
xnor U4333 (N_4333,N_3962,N_3883);
nor U4334 (N_4334,N_3970,N_3647);
nand U4335 (N_4335,N_3731,N_3904);
and U4336 (N_4336,N_3801,N_3927);
and U4337 (N_4337,N_3642,N_3805);
xor U4338 (N_4338,N_3827,N_3951);
or U4339 (N_4339,N_3558,N_3980);
or U4340 (N_4340,N_3972,N_3993);
xor U4341 (N_4341,N_3652,N_3599);
xnor U4342 (N_4342,N_3907,N_3542);
nor U4343 (N_4343,N_3767,N_3732);
xnor U4344 (N_4344,N_3800,N_3761);
or U4345 (N_4345,N_3869,N_3776);
and U4346 (N_4346,N_3995,N_3863);
nand U4347 (N_4347,N_3893,N_3682);
nor U4348 (N_4348,N_3548,N_3794);
xor U4349 (N_4349,N_3877,N_3673);
or U4350 (N_4350,N_3568,N_3978);
nand U4351 (N_4351,N_3523,N_3679);
nand U4352 (N_4352,N_3562,N_3654);
or U4353 (N_4353,N_3922,N_3500);
or U4354 (N_4354,N_3847,N_3774);
nand U4355 (N_4355,N_3941,N_3974);
xor U4356 (N_4356,N_3953,N_3796);
or U4357 (N_4357,N_3957,N_3899);
xnor U4358 (N_4358,N_3670,N_3821);
xor U4359 (N_4359,N_3961,N_3516);
nor U4360 (N_4360,N_3852,N_3789);
or U4361 (N_4361,N_3556,N_3663);
and U4362 (N_4362,N_3860,N_3948);
xor U4363 (N_4363,N_3944,N_3914);
nand U4364 (N_4364,N_3932,N_3511);
or U4365 (N_4365,N_3811,N_3743);
nor U4366 (N_4366,N_3531,N_3963);
xnor U4367 (N_4367,N_3763,N_3505);
xnor U4368 (N_4368,N_3801,N_3654);
nor U4369 (N_4369,N_3870,N_3864);
or U4370 (N_4370,N_3652,N_3650);
and U4371 (N_4371,N_3985,N_3899);
xnor U4372 (N_4372,N_3797,N_3866);
or U4373 (N_4373,N_3869,N_3544);
and U4374 (N_4374,N_3868,N_3526);
and U4375 (N_4375,N_3655,N_3569);
nor U4376 (N_4376,N_3775,N_3641);
or U4377 (N_4377,N_3770,N_3624);
xor U4378 (N_4378,N_3831,N_3537);
nand U4379 (N_4379,N_3744,N_3671);
and U4380 (N_4380,N_3686,N_3962);
and U4381 (N_4381,N_3791,N_3534);
and U4382 (N_4382,N_3990,N_3665);
xnor U4383 (N_4383,N_3792,N_3929);
and U4384 (N_4384,N_3697,N_3628);
xnor U4385 (N_4385,N_3800,N_3726);
nand U4386 (N_4386,N_3994,N_3755);
or U4387 (N_4387,N_3867,N_3846);
and U4388 (N_4388,N_3688,N_3720);
nor U4389 (N_4389,N_3764,N_3760);
xnor U4390 (N_4390,N_3744,N_3779);
xnor U4391 (N_4391,N_3591,N_3884);
or U4392 (N_4392,N_3500,N_3877);
nor U4393 (N_4393,N_3613,N_3554);
nor U4394 (N_4394,N_3756,N_3710);
and U4395 (N_4395,N_3857,N_3652);
nor U4396 (N_4396,N_3607,N_3664);
nand U4397 (N_4397,N_3742,N_3666);
xor U4398 (N_4398,N_3866,N_3720);
nand U4399 (N_4399,N_3533,N_3706);
or U4400 (N_4400,N_3797,N_3546);
xnor U4401 (N_4401,N_3724,N_3962);
xnor U4402 (N_4402,N_3697,N_3906);
xnor U4403 (N_4403,N_3654,N_3940);
or U4404 (N_4404,N_3839,N_3517);
and U4405 (N_4405,N_3874,N_3764);
nand U4406 (N_4406,N_3833,N_3778);
nand U4407 (N_4407,N_3642,N_3524);
or U4408 (N_4408,N_3611,N_3730);
xnor U4409 (N_4409,N_3637,N_3899);
nand U4410 (N_4410,N_3940,N_3728);
nand U4411 (N_4411,N_3857,N_3713);
nor U4412 (N_4412,N_3699,N_3747);
xor U4413 (N_4413,N_3988,N_3811);
and U4414 (N_4414,N_3675,N_3508);
xor U4415 (N_4415,N_3612,N_3688);
or U4416 (N_4416,N_3648,N_3745);
nand U4417 (N_4417,N_3560,N_3768);
nor U4418 (N_4418,N_3729,N_3617);
or U4419 (N_4419,N_3782,N_3937);
or U4420 (N_4420,N_3876,N_3554);
and U4421 (N_4421,N_3700,N_3934);
xnor U4422 (N_4422,N_3632,N_3854);
xor U4423 (N_4423,N_3964,N_3534);
or U4424 (N_4424,N_3912,N_3527);
nor U4425 (N_4425,N_3802,N_3937);
and U4426 (N_4426,N_3513,N_3956);
or U4427 (N_4427,N_3610,N_3960);
nand U4428 (N_4428,N_3703,N_3810);
nand U4429 (N_4429,N_3538,N_3973);
and U4430 (N_4430,N_3595,N_3846);
nand U4431 (N_4431,N_3551,N_3768);
nor U4432 (N_4432,N_3862,N_3650);
nor U4433 (N_4433,N_3917,N_3817);
or U4434 (N_4434,N_3520,N_3544);
or U4435 (N_4435,N_3608,N_3875);
or U4436 (N_4436,N_3577,N_3819);
xnor U4437 (N_4437,N_3905,N_3536);
xor U4438 (N_4438,N_3957,N_3640);
and U4439 (N_4439,N_3970,N_3861);
nand U4440 (N_4440,N_3906,N_3677);
or U4441 (N_4441,N_3683,N_3725);
nor U4442 (N_4442,N_3896,N_3690);
nor U4443 (N_4443,N_3531,N_3876);
nand U4444 (N_4444,N_3986,N_3583);
nand U4445 (N_4445,N_3787,N_3878);
nand U4446 (N_4446,N_3555,N_3609);
xnor U4447 (N_4447,N_3797,N_3603);
and U4448 (N_4448,N_3846,N_3910);
and U4449 (N_4449,N_3799,N_3695);
nor U4450 (N_4450,N_3632,N_3901);
and U4451 (N_4451,N_3748,N_3847);
xnor U4452 (N_4452,N_3561,N_3516);
xor U4453 (N_4453,N_3702,N_3900);
or U4454 (N_4454,N_3825,N_3500);
nor U4455 (N_4455,N_3700,N_3892);
and U4456 (N_4456,N_3611,N_3508);
nand U4457 (N_4457,N_3572,N_3701);
nor U4458 (N_4458,N_3810,N_3888);
nand U4459 (N_4459,N_3563,N_3650);
nand U4460 (N_4460,N_3919,N_3547);
xor U4461 (N_4461,N_3561,N_3507);
nor U4462 (N_4462,N_3664,N_3975);
and U4463 (N_4463,N_3984,N_3603);
xor U4464 (N_4464,N_3548,N_3618);
or U4465 (N_4465,N_3735,N_3810);
nor U4466 (N_4466,N_3759,N_3852);
or U4467 (N_4467,N_3610,N_3655);
and U4468 (N_4468,N_3524,N_3606);
nor U4469 (N_4469,N_3708,N_3795);
nand U4470 (N_4470,N_3768,N_3880);
xnor U4471 (N_4471,N_3865,N_3891);
nand U4472 (N_4472,N_3538,N_3639);
nor U4473 (N_4473,N_3735,N_3532);
or U4474 (N_4474,N_3842,N_3516);
and U4475 (N_4475,N_3775,N_3529);
nand U4476 (N_4476,N_3529,N_3887);
or U4477 (N_4477,N_3739,N_3621);
xor U4478 (N_4478,N_3816,N_3630);
and U4479 (N_4479,N_3989,N_3611);
and U4480 (N_4480,N_3679,N_3559);
or U4481 (N_4481,N_3950,N_3766);
and U4482 (N_4482,N_3958,N_3707);
xor U4483 (N_4483,N_3596,N_3705);
nand U4484 (N_4484,N_3828,N_3805);
nand U4485 (N_4485,N_3505,N_3923);
nor U4486 (N_4486,N_3836,N_3585);
nand U4487 (N_4487,N_3894,N_3563);
nor U4488 (N_4488,N_3951,N_3576);
xor U4489 (N_4489,N_3624,N_3515);
and U4490 (N_4490,N_3881,N_3864);
or U4491 (N_4491,N_3525,N_3760);
nand U4492 (N_4492,N_3827,N_3789);
xor U4493 (N_4493,N_3818,N_3678);
xnor U4494 (N_4494,N_3672,N_3821);
nand U4495 (N_4495,N_3956,N_3641);
nand U4496 (N_4496,N_3831,N_3959);
or U4497 (N_4497,N_3915,N_3698);
xor U4498 (N_4498,N_3903,N_3941);
nor U4499 (N_4499,N_3976,N_3987);
or U4500 (N_4500,N_4074,N_4406);
nor U4501 (N_4501,N_4470,N_4227);
or U4502 (N_4502,N_4361,N_4004);
or U4503 (N_4503,N_4363,N_4120);
or U4504 (N_4504,N_4332,N_4371);
nor U4505 (N_4505,N_4108,N_4310);
xor U4506 (N_4506,N_4170,N_4494);
nand U4507 (N_4507,N_4401,N_4482);
and U4508 (N_4508,N_4005,N_4015);
nand U4509 (N_4509,N_4404,N_4391);
or U4510 (N_4510,N_4331,N_4422);
nand U4511 (N_4511,N_4408,N_4014);
nor U4512 (N_4512,N_4385,N_4091);
and U4513 (N_4513,N_4233,N_4127);
nor U4514 (N_4514,N_4119,N_4435);
nand U4515 (N_4515,N_4180,N_4319);
and U4516 (N_4516,N_4322,N_4380);
or U4517 (N_4517,N_4265,N_4316);
or U4518 (N_4518,N_4354,N_4295);
xnor U4519 (N_4519,N_4365,N_4036);
nand U4520 (N_4520,N_4344,N_4444);
xor U4521 (N_4521,N_4343,N_4457);
nor U4522 (N_4522,N_4258,N_4166);
nand U4523 (N_4523,N_4135,N_4184);
nand U4524 (N_4524,N_4273,N_4282);
nor U4525 (N_4525,N_4025,N_4461);
nand U4526 (N_4526,N_4023,N_4008);
nand U4527 (N_4527,N_4414,N_4205);
nand U4528 (N_4528,N_4255,N_4153);
xor U4529 (N_4529,N_4218,N_4424);
and U4530 (N_4530,N_4341,N_4381);
and U4531 (N_4531,N_4201,N_4202);
and U4532 (N_4532,N_4474,N_4433);
nor U4533 (N_4533,N_4021,N_4421);
xor U4534 (N_4534,N_4291,N_4378);
xnor U4535 (N_4535,N_4191,N_4017);
xnor U4536 (N_4536,N_4056,N_4204);
or U4537 (N_4537,N_4309,N_4146);
nand U4538 (N_4538,N_4054,N_4376);
nor U4539 (N_4539,N_4216,N_4425);
nor U4540 (N_4540,N_4210,N_4219);
and U4541 (N_4541,N_4411,N_4050);
xor U4542 (N_4542,N_4304,N_4045);
nand U4543 (N_4543,N_4415,N_4386);
or U4544 (N_4544,N_4040,N_4167);
nand U4545 (N_4545,N_4278,N_4335);
nand U4546 (N_4546,N_4149,N_4181);
or U4547 (N_4547,N_4007,N_4152);
nand U4548 (N_4548,N_4075,N_4061);
nor U4549 (N_4549,N_4031,N_4193);
xnor U4550 (N_4550,N_4360,N_4409);
nand U4551 (N_4551,N_4147,N_4397);
or U4552 (N_4552,N_4093,N_4122);
xor U4553 (N_4553,N_4456,N_4328);
xnor U4554 (N_4554,N_4028,N_4038);
or U4555 (N_4555,N_4246,N_4215);
xnor U4556 (N_4556,N_4357,N_4434);
or U4557 (N_4557,N_4418,N_4020);
nand U4558 (N_4558,N_4275,N_4116);
or U4559 (N_4559,N_4262,N_4329);
and U4560 (N_4560,N_4213,N_4492);
nor U4561 (N_4561,N_4398,N_4057);
nand U4562 (N_4562,N_4009,N_4067);
xnor U4563 (N_4563,N_4000,N_4231);
nor U4564 (N_4564,N_4345,N_4419);
nand U4565 (N_4565,N_4128,N_4268);
or U4566 (N_4566,N_4438,N_4251);
nand U4567 (N_4567,N_4445,N_4306);
nand U4568 (N_4568,N_4078,N_4163);
xor U4569 (N_4569,N_4129,N_4261);
nand U4570 (N_4570,N_4035,N_4179);
and U4571 (N_4571,N_4252,N_4307);
nor U4572 (N_4572,N_4452,N_4432);
and U4573 (N_4573,N_4175,N_4157);
and U4574 (N_4574,N_4214,N_4041);
or U4575 (N_4575,N_4126,N_4292);
xor U4576 (N_4576,N_4393,N_4467);
or U4577 (N_4577,N_4182,N_4453);
or U4578 (N_4578,N_4177,N_4185);
nor U4579 (N_4579,N_4373,N_4294);
and U4580 (N_4580,N_4440,N_4417);
xor U4581 (N_4581,N_4480,N_4084);
nand U4582 (N_4582,N_4264,N_4188);
xnor U4583 (N_4583,N_4387,N_4172);
nor U4584 (N_4584,N_4465,N_4248);
nor U4585 (N_4585,N_4109,N_4475);
or U4586 (N_4586,N_4018,N_4131);
or U4587 (N_4587,N_4199,N_4187);
xor U4588 (N_4588,N_4276,N_4263);
nand U4589 (N_4589,N_4374,N_4174);
nand U4590 (N_4590,N_4266,N_4337);
xnor U4591 (N_4591,N_4159,N_4256);
and U4592 (N_4592,N_4220,N_4441);
nand U4593 (N_4593,N_4479,N_4290);
or U4594 (N_4594,N_4112,N_4383);
nand U4595 (N_4595,N_4455,N_4446);
nand U4596 (N_4596,N_4469,N_4229);
and U4597 (N_4597,N_4176,N_4064);
nand U4598 (N_4598,N_4019,N_4171);
nand U4599 (N_4599,N_4254,N_4058);
nor U4600 (N_4600,N_4087,N_4250);
and U4601 (N_4601,N_4355,N_4285);
or U4602 (N_4602,N_4339,N_4097);
xnor U4603 (N_4603,N_4013,N_4267);
or U4604 (N_4604,N_4002,N_4110);
or U4605 (N_4605,N_4208,N_4001);
nand U4606 (N_4606,N_4423,N_4113);
and U4607 (N_4607,N_4403,N_4111);
nor U4608 (N_4608,N_4142,N_4428);
or U4609 (N_4609,N_4103,N_4396);
nand U4610 (N_4610,N_4079,N_4346);
nand U4611 (N_4611,N_4379,N_4407);
and U4612 (N_4612,N_4338,N_4459);
nor U4613 (N_4613,N_4235,N_4194);
nand U4614 (N_4614,N_4493,N_4160);
xor U4615 (N_4615,N_4249,N_4144);
nand U4616 (N_4616,N_4260,N_4301);
xnor U4617 (N_4617,N_4240,N_4454);
and U4618 (N_4618,N_4431,N_4281);
or U4619 (N_4619,N_4311,N_4498);
nor U4620 (N_4620,N_4137,N_4302);
or U4621 (N_4621,N_4083,N_4101);
nand U4622 (N_4622,N_4359,N_4217);
xor U4623 (N_4623,N_4351,N_4037);
and U4624 (N_4624,N_4450,N_4155);
and U4625 (N_4625,N_4165,N_4464);
nor U4626 (N_4626,N_4222,N_4226);
xor U4627 (N_4627,N_4118,N_4062);
xor U4628 (N_4628,N_4297,N_4388);
xnor U4629 (N_4629,N_4224,N_4347);
or U4630 (N_4630,N_4169,N_4089);
and U4631 (N_4631,N_4390,N_4121);
or U4632 (N_4632,N_4148,N_4203);
xnor U4633 (N_4633,N_4490,N_4139);
nor U4634 (N_4634,N_4211,N_4032);
or U4635 (N_4635,N_4356,N_4162);
xnor U4636 (N_4636,N_4313,N_4367);
and U4637 (N_4637,N_4234,N_4195);
nor U4638 (N_4638,N_4033,N_4027);
nand U4639 (N_4639,N_4186,N_4238);
nor U4640 (N_4640,N_4189,N_4039);
nand U4641 (N_4641,N_4065,N_4197);
and U4642 (N_4642,N_4140,N_4134);
and U4643 (N_4643,N_4099,N_4049);
xnor U4644 (N_4644,N_4342,N_4308);
or U4645 (N_4645,N_4236,N_4198);
and U4646 (N_4646,N_4042,N_4353);
or U4647 (N_4647,N_4427,N_4068);
nand U4648 (N_4648,N_4420,N_4066);
and U4649 (N_4649,N_4447,N_4488);
nand U4650 (N_4650,N_4491,N_4340);
xor U4651 (N_4651,N_4489,N_4468);
or U4652 (N_4652,N_4105,N_4053);
or U4653 (N_4653,N_4288,N_4048);
xor U4654 (N_4654,N_4471,N_4326);
nand U4655 (N_4655,N_4026,N_4259);
nor U4656 (N_4656,N_4085,N_4496);
or U4657 (N_4657,N_4164,N_4003);
nand U4658 (N_4658,N_4283,N_4375);
nand U4659 (N_4659,N_4449,N_4034);
xnor U4660 (N_4660,N_4270,N_4377);
xor U4661 (N_4661,N_4130,N_4124);
xor U4662 (N_4662,N_4429,N_4368);
nor U4663 (N_4663,N_4138,N_4312);
nand U4664 (N_4664,N_4132,N_4253);
xor U4665 (N_4665,N_4069,N_4389);
nor U4666 (N_4666,N_4392,N_4463);
nor U4667 (N_4667,N_4272,N_4296);
and U4668 (N_4668,N_4333,N_4209);
and U4669 (N_4669,N_4060,N_4245);
xor U4670 (N_4670,N_4030,N_4466);
or U4671 (N_4671,N_4200,N_4369);
and U4672 (N_4672,N_4237,N_4416);
and U4673 (N_4673,N_4104,N_4293);
xor U4674 (N_4674,N_4358,N_4076);
and U4675 (N_4675,N_4451,N_4043);
or U4676 (N_4676,N_4145,N_4046);
and U4677 (N_4677,N_4228,N_4320);
and U4678 (N_4678,N_4442,N_4168);
nand U4679 (N_4679,N_4289,N_4044);
xnor U4680 (N_4680,N_4114,N_4458);
xor U4681 (N_4681,N_4484,N_4269);
and U4682 (N_4682,N_4239,N_4192);
or U4683 (N_4683,N_4151,N_4395);
and U4684 (N_4684,N_4212,N_4399);
or U4685 (N_4685,N_4221,N_4412);
and U4686 (N_4686,N_4115,N_4400);
nand U4687 (N_4687,N_4277,N_4321);
xor U4688 (N_4688,N_4315,N_4052);
nand U4689 (N_4689,N_4225,N_4095);
nand U4690 (N_4690,N_4318,N_4323);
nor U4691 (N_4691,N_4244,N_4125);
nand U4692 (N_4692,N_4497,N_4370);
or U4693 (N_4693,N_4081,N_4232);
nor U4694 (N_4694,N_4243,N_4071);
xnor U4695 (N_4695,N_4372,N_4107);
nand U4696 (N_4696,N_4055,N_4051);
or U4697 (N_4697,N_4460,N_4499);
nand U4698 (N_4698,N_4394,N_4024);
or U4699 (N_4699,N_4047,N_4082);
or U4700 (N_4700,N_4366,N_4156);
nor U4701 (N_4701,N_4063,N_4348);
or U4702 (N_4702,N_4206,N_4336);
nand U4703 (N_4703,N_4384,N_4006);
xor U4704 (N_4704,N_4413,N_4059);
xnor U4705 (N_4705,N_4223,N_4092);
or U4706 (N_4706,N_4257,N_4314);
or U4707 (N_4707,N_4280,N_4305);
and U4708 (N_4708,N_4477,N_4010);
nand U4709 (N_4709,N_4136,N_4462);
xor U4710 (N_4710,N_4405,N_4102);
nand U4711 (N_4711,N_4382,N_4196);
or U4712 (N_4712,N_4173,N_4011);
and U4713 (N_4713,N_4443,N_4016);
and U4714 (N_4714,N_4247,N_4486);
xor U4715 (N_4715,N_4284,N_4086);
or U4716 (N_4716,N_4279,N_4100);
xnor U4717 (N_4717,N_4271,N_4487);
xnor U4718 (N_4718,N_4436,N_4094);
xor U4719 (N_4719,N_4352,N_4241);
and U4720 (N_4720,N_4299,N_4349);
xnor U4721 (N_4721,N_4481,N_4154);
nand U4722 (N_4722,N_4077,N_4230);
and U4723 (N_4723,N_4426,N_4090);
or U4724 (N_4724,N_4096,N_4287);
and U4725 (N_4725,N_4473,N_4012);
nor U4726 (N_4726,N_4073,N_4158);
xnor U4727 (N_4727,N_4483,N_4123);
or U4728 (N_4728,N_4303,N_4410);
nor U4729 (N_4729,N_4350,N_4324);
or U4730 (N_4730,N_4133,N_4242);
xnor U4731 (N_4731,N_4317,N_4286);
and U4732 (N_4732,N_4080,N_4476);
nor U4733 (N_4733,N_4495,N_4106);
xnor U4734 (N_4734,N_4448,N_4143);
and U4735 (N_4735,N_4088,N_4274);
xor U4736 (N_4736,N_4485,N_4141);
or U4737 (N_4737,N_4439,N_4298);
and U4738 (N_4738,N_4364,N_4022);
nand U4739 (N_4739,N_4183,N_4029);
nand U4740 (N_4740,N_4437,N_4207);
xnor U4741 (N_4741,N_4362,N_4327);
xnor U4742 (N_4742,N_4178,N_4161);
xor U4743 (N_4743,N_4330,N_4072);
and U4744 (N_4744,N_4117,N_4325);
nand U4745 (N_4745,N_4430,N_4070);
nand U4746 (N_4746,N_4478,N_4190);
and U4747 (N_4747,N_4402,N_4300);
nor U4748 (N_4748,N_4472,N_4334);
and U4749 (N_4749,N_4098,N_4150);
or U4750 (N_4750,N_4372,N_4357);
xnor U4751 (N_4751,N_4218,N_4304);
nor U4752 (N_4752,N_4391,N_4224);
nand U4753 (N_4753,N_4428,N_4450);
xor U4754 (N_4754,N_4444,N_4111);
and U4755 (N_4755,N_4163,N_4324);
or U4756 (N_4756,N_4276,N_4482);
xor U4757 (N_4757,N_4291,N_4157);
xnor U4758 (N_4758,N_4244,N_4375);
nand U4759 (N_4759,N_4096,N_4100);
and U4760 (N_4760,N_4366,N_4078);
nand U4761 (N_4761,N_4043,N_4495);
xor U4762 (N_4762,N_4402,N_4045);
and U4763 (N_4763,N_4436,N_4366);
nor U4764 (N_4764,N_4208,N_4377);
xnor U4765 (N_4765,N_4467,N_4263);
and U4766 (N_4766,N_4301,N_4083);
nor U4767 (N_4767,N_4067,N_4203);
or U4768 (N_4768,N_4310,N_4460);
xor U4769 (N_4769,N_4280,N_4010);
and U4770 (N_4770,N_4209,N_4499);
and U4771 (N_4771,N_4126,N_4398);
xnor U4772 (N_4772,N_4369,N_4250);
nor U4773 (N_4773,N_4339,N_4166);
nand U4774 (N_4774,N_4167,N_4262);
nand U4775 (N_4775,N_4071,N_4372);
xor U4776 (N_4776,N_4352,N_4129);
nor U4777 (N_4777,N_4000,N_4133);
nand U4778 (N_4778,N_4021,N_4293);
nand U4779 (N_4779,N_4321,N_4440);
or U4780 (N_4780,N_4185,N_4049);
or U4781 (N_4781,N_4210,N_4361);
nor U4782 (N_4782,N_4267,N_4294);
and U4783 (N_4783,N_4183,N_4390);
xor U4784 (N_4784,N_4341,N_4143);
and U4785 (N_4785,N_4001,N_4481);
xnor U4786 (N_4786,N_4005,N_4266);
nor U4787 (N_4787,N_4298,N_4218);
nand U4788 (N_4788,N_4472,N_4407);
or U4789 (N_4789,N_4308,N_4274);
nor U4790 (N_4790,N_4039,N_4090);
nand U4791 (N_4791,N_4171,N_4292);
xnor U4792 (N_4792,N_4046,N_4271);
nand U4793 (N_4793,N_4105,N_4163);
or U4794 (N_4794,N_4480,N_4170);
and U4795 (N_4795,N_4409,N_4154);
and U4796 (N_4796,N_4422,N_4297);
nor U4797 (N_4797,N_4162,N_4292);
and U4798 (N_4798,N_4383,N_4095);
xor U4799 (N_4799,N_4491,N_4294);
and U4800 (N_4800,N_4232,N_4277);
nand U4801 (N_4801,N_4353,N_4440);
nor U4802 (N_4802,N_4171,N_4000);
and U4803 (N_4803,N_4185,N_4200);
xnor U4804 (N_4804,N_4311,N_4353);
xnor U4805 (N_4805,N_4432,N_4060);
or U4806 (N_4806,N_4049,N_4379);
and U4807 (N_4807,N_4457,N_4238);
xor U4808 (N_4808,N_4405,N_4263);
or U4809 (N_4809,N_4239,N_4466);
or U4810 (N_4810,N_4190,N_4493);
nand U4811 (N_4811,N_4160,N_4459);
or U4812 (N_4812,N_4425,N_4445);
or U4813 (N_4813,N_4023,N_4069);
xnor U4814 (N_4814,N_4133,N_4322);
nor U4815 (N_4815,N_4185,N_4088);
and U4816 (N_4816,N_4478,N_4150);
xnor U4817 (N_4817,N_4256,N_4374);
nor U4818 (N_4818,N_4489,N_4142);
and U4819 (N_4819,N_4441,N_4125);
or U4820 (N_4820,N_4317,N_4045);
xnor U4821 (N_4821,N_4111,N_4224);
nor U4822 (N_4822,N_4447,N_4090);
and U4823 (N_4823,N_4387,N_4380);
xnor U4824 (N_4824,N_4088,N_4047);
and U4825 (N_4825,N_4468,N_4333);
xor U4826 (N_4826,N_4403,N_4491);
nand U4827 (N_4827,N_4457,N_4416);
nand U4828 (N_4828,N_4177,N_4388);
and U4829 (N_4829,N_4244,N_4138);
and U4830 (N_4830,N_4154,N_4202);
or U4831 (N_4831,N_4071,N_4064);
xnor U4832 (N_4832,N_4195,N_4439);
and U4833 (N_4833,N_4204,N_4389);
nand U4834 (N_4834,N_4269,N_4477);
xor U4835 (N_4835,N_4063,N_4389);
and U4836 (N_4836,N_4074,N_4120);
xor U4837 (N_4837,N_4072,N_4021);
nand U4838 (N_4838,N_4430,N_4254);
nand U4839 (N_4839,N_4092,N_4356);
or U4840 (N_4840,N_4473,N_4172);
or U4841 (N_4841,N_4394,N_4343);
xnor U4842 (N_4842,N_4448,N_4365);
or U4843 (N_4843,N_4151,N_4118);
and U4844 (N_4844,N_4399,N_4403);
and U4845 (N_4845,N_4261,N_4284);
nand U4846 (N_4846,N_4226,N_4166);
and U4847 (N_4847,N_4406,N_4316);
nand U4848 (N_4848,N_4107,N_4077);
nor U4849 (N_4849,N_4133,N_4197);
nand U4850 (N_4850,N_4061,N_4042);
nand U4851 (N_4851,N_4430,N_4022);
and U4852 (N_4852,N_4379,N_4312);
and U4853 (N_4853,N_4480,N_4389);
nand U4854 (N_4854,N_4406,N_4486);
nor U4855 (N_4855,N_4450,N_4426);
and U4856 (N_4856,N_4368,N_4353);
xnor U4857 (N_4857,N_4165,N_4366);
nor U4858 (N_4858,N_4205,N_4088);
xnor U4859 (N_4859,N_4086,N_4486);
and U4860 (N_4860,N_4062,N_4387);
xnor U4861 (N_4861,N_4312,N_4173);
xnor U4862 (N_4862,N_4347,N_4165);
nor U4863 (N_4863,N_4199,N_4122);
and U4864 (N_4864,N_4039,N_4422);
nor U4865 (N_4865,N_4042,N_4080);
and U4866 (N_4866,N_4067,N_4395);
nor U4867 (N_4867,N_4223,N_4456);
xnor U4868 (N_4868,N_4069,N_4226);
nor U4869 (N_4869,N_4264,N_4491);
xor U4870 (N_4870,N_4272,N_4338);
nor U4871 (N_4871,N_4366,N_4000);
nand U4872 (N_4872,N_4380,N_4489);
nand U4873 (N_4873,N_4110,N_4174);
nand U4874 (N_4874,N_4334,N_4387);
nand U4875 (N_4875,N_4166,N_4005);
xor U4876 (N_4876,N_4358,N_4455);
and U4877 (N_4877,N_4307,N_4288);
nor U4878 (N_4878,N_4438,N_4222);
xnor U4879 (N_4879,N_4003,N_4292);
xnor U4880 (N_4880,N_4249,N_4465);
and U4881 (N_4881,N_4097,N_4069);
nor U4882 (N_4882,N_4044,N_4262);
or U4883 (N_4883,N_4179,N_4336);
nand U4884 (N_4884,N_4053,N_4433);
nor U4885 (N_4885,N_4327,N_4046);
xnor U4886 (N_4886,N_4418,N_4345);
and U4887 (N_4887,N_4145,N_4028);
nand U4888 (N_4888,N_4468,N_4454);
and U4889 (N_4889,N_4033,N_4431);
or U4890 (N_4890,N_4360,N_4219);
and U4891 (N_4891,N_4133,N_4428);
nor U4892 (N_4892,N_4012,N_4168);
nor U4893 (N_4893,N_4418,N_4430);
nand U4894 (N_4894,N_4468,N_4444);
xnor U4895 (N_4895,N_4118,N_4274);
xnor U4896 (N_4896,N_4477,N_4313);
nor U4897 (N_4897,N_4473,N_4091);
nand U4898 (N_4898,N_4105,N_4055);
xor U4899 (N_4899,N_4191,N_4237);
or U4900 (N_4900,N_4161,N_4482);
nand U4901 (N_4901,N_4248,N_4070);
nor U4902 (N_4902,N_4019,N_4365);
xor U4903 (N_4903,N_4326,N_4364);
nor U4904 (N_4904,N_4387,N_4492);
or U4905 (N_4905,N_4494,N_4324);
and U4906 (N_4906,N_4075,N_4119);
nor U4907 (N_4907,N_4281,N_4237);
nor U4908 (N_4908,N_4262,N_4196);
xnor U4909 (N_4909,N_4000,N_4415);
and U4910 (N_4910,N_4312,N_4412);
xor U4911 (N_4911,N_4386,N_4265);
nor U4912 (N_4912,N_4461,N_4070);
or U4913 (N_4913,N_4240,N_4077);
xnor U4914 (N_4914,N_4212,N_4273);
or U4915 (N_4915,N_4489,N_4473);
or U4916 (N_4916,N_4040,N_4110);
nand U4917 (N_4917,N_4117,N_4167);
xor U4918 (N_4918,N_4251,N_4465);
nor U4919 (N_4919,N_4365,N_4030);
nand U4920 (N_4920,N_4214,N_4429);
nor U4921 (N_4921,N_4020,N_4382);
or U4922 (N_4922,N_4413,N_4289);
nand U4923 (N_4923,N_4402,N_4266);
nor U4924 (N_4924,N_4059,N_4437);
nand U4925 (N_4925,N_4311,N_4025);
and U4926 (N_4926,N_4078,N_4340);
nor U4927 (N_4927,N_4301,N_4038);
or U4928 (N_4928,N_4306,N_4061);
and U4929 (N_4929,N_4316,N_4407);
nor U4930 (N_4930,N_4417,N_4032);
nor U4931 (N_4931,N_4241,N_4440);
nand U4932 (N_4932,N_4009,N_4024);
or U4933 (N_4933,N_4104,N_4389);
nand U4934 (N_4934,N_4264,N_4184);
nand U4935 (N_4935,N_4318,N_4241);
nor U4936 (N_4936,N_4464,N_4390);
or U4937 (N_4937,N_4457,N_4381);
nor U4938 (N_4938,N_4445,N_4175);
or U4939 (N_4939,N_4374,N_4100);
nor U4940 (N_4940,N_4269,N_4341);
xor U4941 (N_4941,N_4355,N_4087);
and U4942 (N_4942,N_4247,N_4040);
nor U4943 (N_4943,N_4281,N_4319);
nor U4944 (N_4944,N_4042,N_4363);
nor U4945 (N_4945,N_4420,N_4021);
or U4946 (N_4946,N_4035,N_4437);
nand U4947 (N_4947,N_4180,N_4493);
nand U4948 (N_4948,N_4314,N_4095);
xnor U4949 (N_4949,N_4222,N_4338);
xor U4950 (N_4950,N_4142,N_4337);
nand U4951 (N_4951,N_4359,N_4145);
xnor U4952 (N_4952,N_4456,N_4246);
nand U4953 (N_4953,N_4348,N_4389);
nand U4954 (N_4954,N_4381,N_4224);
or U4955 (N_4955,N_4306,N_4014);
and U4956 (N_4956,N_4362,N_4454);
xor U4957 (N_4957,N_4323,N_4093);
nand U4958 (N_4958,N_4145,N_4067);
or U4959 (N_4959,N_4408,N_4481);
xor U4960 (N_4960,N_4027,N_4140);
nor U4961 (N_4961,N_4427,N_4214);
xnor U4962 (N_4962,N_4159,N_4390);
nand U4963 (N_4963,N_4437,N_4156);
or U4964 (N_4964,N_4421,N_4276);
xnor U4965 (N_4965,N_4019,N_4490);
nor U4966 (N_4966,N_4108,N_4454);
nand U4967 (N_4967,N_4136,N_4024);
nand U4968 (N_4968,N_4246,N_4024);
and U4969 (N_4969,N_4035,N_4076);
nand U4970 (N_4970,N_4127,N_4031);
xnor U4971 (N_4971,N_4042,N_4215);
and U4972 (N_4972,N_4108,N_4235);
nand U4973 (N_4973,N_4282,N_4264);
nor U4974 (N_4974,N_4492,N_4397);
or U4975 (N_4975,N_4453,N_4135);
nand U4976 (N_4976,N_4026,N_4201);
or U4977 (N_4977,N_4110,N_4293);
nand U4978 (N_4978,N_4340,N_4045);
nor U4979 (N_4979,N_4160,N_4166);
and U4980 (N_4980,N_4087,N_4377);
xnor U4981 (N_4981,N_4435,N_4410);
xnor U4982 (N_4982,N_4497,N_4248);
nor U4983 (N_4983,N_4108,N_4013);
or U4984 (N_4984,N_4029,N_4237);
or U4985 (N_4985,N_4410,N_4295);
or U4986 (N_4986,N_4153,N_4194);
and U4987 (N_4987,N_4023,N_4411);
xor U4988 (N_4988,N_4043,N_4361);
or U4989 (N_4989,N_4196,N_4066);
xnor U4990 (N_4990,N_4123,N_4337);
nor U4991 (N_4991,N_4331,N_4100);
nand U4992 (N_4992,N_4280,N_4379);
and U4993 (N_4993,N_4354,N_4462);
and U4994 (N_4994,N_4223,N_4396);
xor U4995 (N_4995,N_4001,N_4199);
xnor U4996 (N_4996,N_4428,N_4211);
or U4997 (N_4997,N_4323,N_4422);
and U4998 (N_4998,N_4131,N_4061);
and U4999 (N_4999,N_4420,N_4032);
nor U5000 (N_5000,N_4632,N_4510);
or U5001 (N_5001,N_4720,N_4509);
nand U5002 (N_5002,N_4679,N_4542);
or U5003 (N_5003,N_4746,N_4996);
nor U5004 (N_5004,N_4858,N_4845);
or U5005 (N_5005,N_4979,N_4687);
xor U5006 (N_5006,N_4909,N_4520);
nor U5007 (N_5007,N_4659,N_4837);
xor U5008 (N_5008,N_4727,N_4886);
or U5009 (N_5009,N_4770,N_4622);
or U5010 (N_5010,N_4648,N_4818);
nand U5011 (N_5011,N_4904,N_4983);
or U5012 (N_5012,N_4950,N_4742);
or U5013 (N_5013,N_4824,N_4676);
nand U5014 (N_5014,N_4829,N_4760);
or U5015 (N_5015,N_4800,N_4876);
or U5016 (N_5016,N_4976,N_4893);
and U5017 (N_5017,N_4888,N_4777);
nand U5018 (N_5018,N_4743,N_4568);
and U5019 (N_5019,N_4582,N_4629);
xor U5020 (N_5020,N_4724,N_4719);
or U5021 (N_5021,N_4994,N_4600);
or U5022 (N_5022,N_4998,N_4645);
nand U5023 (N_5023,N_4710,N_4534);
xnor U5024 (N_5024,N_4574,N_4641);
and U5025 (N_5025,N_4736,N_4847);
xnor U5026 (N_5026,N_4682,N_4587);
xor U5027 (N_5027,N_4821,N_4572);
or U5028 (N_5028,N_4913,N_4581);
nor U5029 (N_5029,N_4541,N_4854);
or U5030 (N_5030,N_4717,N_4855);
and U5031 (N_5031,N_4563,N_4506);
nor U5032 (N_5032,N_4671,N_4741);
xor U5033 (N_5033,N_4834,N_4929);
nand U5034 (N_5034,N_4969,N_4851);
or U5035 (N_5035,N_4762,N_4898);
or U5036 (N_5036,N_4623,N_4519);
xor U5037 (N_5037,N_4780,N_4795);
or U5038 (N_5038,N_4840,N_4995);
xor U5039 (N_5039,N_4726,N_4778);
nand U5040 (N_5040,N_4836,N_4814);
nor U5041 (N_5041,N_4784,N_4722);
or U5042 (N_5042,N_4993,N_4702);
nor U5043 (N_5043,N_4941,N_4947);
nand U5044 (N_5044,N_4966,N_4763);
nand U5045 (N_5045,N_4677,N_4816);
xor U5046 (N_5046,N_4889,N_4959);
nand U5047 (N_5047,N_4631,N_4859);
nor U5048 (N_5048,N_4723,N_4967);
nor U5049 (N_5049,N_4644,N_4903);
xor U5050 (N_5050,N_4711,N_4612);
or U5051 (N_5051,N_4865,N_4730);
or U5052 (N_5052,N_4557,N_4655);
and U5053 (N_5053,N_4954,N_4672);
nand U5054 (N_5054,N_4789,N_4828);
nor U5055 (N_5055,N_4586,N_4508);
or U5056 (N_5056,N_4921,N_4625);
nand U5057 (N_5057,N_4968,N_4652);
nand U5058 (N_5058,N_4850,N_4963);
nand U5059 (N_5059,N_4565,N_4566);
xor U5060 (N_5060,N_4986,N_4887);
or U5061 (N_5061,N_4694,N_4708);
xor U5062 (N_5062,N_4755,N_4779);
nor U5063 (N_5063,N_4759,N_4635);
and U5064 (N_5064,N_4756,N_4598);
xor U5065 (N_5065,N_4788,N_4806);
and U5066 (N_5066,N_4626,N_4826);
nor U5067 (N_5067,N_4924,N_4656);
nor U5068 (N_5068,N_4750,N_4544);
xor U5069 (N_5069,N_4856,N_4670);
and U5070 (N_5070,N_4545,N_4513);
or U5071 (N_5071,N_4906,N_4945);
nor U5072 (N_5072,N_4658,N_4879);
and U5073 (N_5073,N_4901,N_4864);
and U5074 (N_5074,N_4737,N_4897);
xnor U5075 (N_5075,N_4857,N_4740);
or U5076 (N_5076,N_4604,N_4504);
or U5077 (N_5077,N_4646,N_4522);
nor U5078 (N_5078,N_4827,N_4546);
xnor U5079 (N_5079,N_4914,N_4628);
nor U5080 (N_5080,N_4621,N_4819);
or U5081 (N_5081,N_4804,N_4744);
xor U5082 (N_5082,N_4558,N_4503);
nor U5083 (N_5083,N_4601,N_4877);
xor U5084 (N_5084,N_4961,N_4787);
nand U5085 (N_5085,N_4725,N_4946);
and U5086 (N_5086,N_4807,N_4982);
xor U5087 (N_5087,N_4577,N_4922);
nor U5088 (N_5088,N_4585,N_4505);
nand U5089 (N_5089,N_4823,N_4507);
and U5090 (N_5090,N_4665,N_4956);
and U5091 (N_5091,N_4797,N_4521);
and U5092 (N_5092,N_4987,N_4799);
and U5093 (N_5093,N_4562,N_4543);
xnor U5094 (N_5094,N_4874,N_4917);
and U5095 (N_5095,N_4928,N_4860);
nor U5096 (N_5096,N_4576,N_4637);
nor U5097 (N_5097,N_4617,N_4571);
and U5098 (N_5098,N_4932,N_4761);
and U5099 (N_5099,N_4939,N_4943);
and U5100 (N_5100,N_4796,N_4841);
nor U5101 (N_5101,N_4531,N_4697);
nor U5102 (N_5102,N_4844,N_4957);
and U5103 (N_5103,N_4811,N_4525);
nand U5104 (N_5104,N_4692,N_4530);
nand U5105 (N_5105,N_4989,N_4822);
nand U5106 (N_5106,N_4684,N_4942);
or U5107 (N_5107,N_4579,N_4925);
nor U5108 (N_5108,N_4895,N_4552);
nand U5109 (N_5109,N_4920,N_4892);
nor U5110 (N_5110,N_4547,N_4614);
xor U5111 (N_5111,N_4825,N_4935);
nand U5112 (N_5112,N_4607,N_4754);
nor U5113 (N_5113,N_4785,N_4907);
nand U5114 (N_5114,N_4790,N_4870);
nor U5115 (N_5115,N_4634,N_4685);
and U5116 (N_5116,N_4872,N_4638);
xor U5117 (N_5117,N_4538,N_4540);
or U5118 (N_5118,N_4820,N_4782);
or U5119 (N_5119,N_4813,N_4731);
and U5120 (N_5120,N_4700,N_4657);
or U5121 (N_5121,N_4846,N_4765);
xor U5122 (N_5122,N_4919,N_4690);
and U5123 (N_5123,N_4709,N_4523);
or U5124 (N_5124,N_4798,N_4931);
xor U5125 (N_5125,N_4609,N_4599);
and U5126 (N_5126,N_4596,N_4535);
or U5127 (N_5127,N_4583,N_4771);
nor U5128 (N_5128,N_4866,N_4647);
or U5129 (N_5129,N_4526,N_4564);
xor U5130 (N_5130,N_4593,N_4990);
nor U5131 (N_5131,N_4516,N_4749);
nand U5132 (N_5132,N_4615,N_4616);
or U5133 (N_5133,N_4733,N_4960);
and U5134 (N_5134,N_4686,N_4934);
and U5135 (N_5135,N_4680,N_4775);
nand U5136 (N_5136,N_4970,N_4768);
or U5137 (N_5137,N_4611,N_4654);
xor U5138 (N_5138,N_4958,N_4649);
nand U5139 (N_5139,N_4691,N_4550);
nor U5140 (N_5140,N_4774,N_4630);
and U5141 (N_5141,N_4606,N_4643);
and U5142 (N_5142,N_4529,N_4739);
nand U5143 (N_5143,N_4962,N_4938);
or U5144 (N_5144,N_4991,N_4964);
or U5145 (N_5145,N_4885,N_4537);
xor U5146 (N_5146,N_4512,N_4908);
xnor U5147 (N_5147,N_4764,N_4704);
nand U5148 (N_5148,N_4642,N_4873);
xor U5149 (N_5149,N_4910,N_4891);
and U5150 (N_5150,N_4911,N_4619);
nand U5151 (N_5151,N_4718,N_4666);
xnor U5152 (N_5152,N_4703,N_4899);
nor U5153 (N_5153,N_4861,N_4772);
nand U5154 (N_5154,N_4830,N_4668);
xnor U5155 (N_5155,N_4636,N_4849);
and U5156 (N_5156,N_4949,N_4548);
nor U5157 (N_5157,N_4735,N_4862);
and U5158 (N_5158,N_4902,N_4868);
or U5159 (N_5159,N_4975,N_4624);
nor U5160 (N_5160,N_4751,N_4580);
and U5161 (N_5161,N_4984,N_4882);
nor U5162 (N_5162,N_4588,N_4595);
and U5163 (N_5163,N_4878,N_4705);
nor U5164 (N_5164,N_4992,N_4880);
nand U5165 (N_5165,N_4732,N_4524);
nand U5166 (N_5166,N_4613,N_4940);
nor U5167 (N_5167,N_4890,N_4675);
and U5168 (N_5168,N_4663,N_4618);
nand U5169 (N_5169,N_4933,N_4955);
and U5170 (N_5170,N_4833,N_4681);
or U5171 (N_5171,N_4783,N_4867);
nor U5172 (N_5172,N_4747,N_4594);
xnor U5173 (N_5173,N_4673,N_4721);
xnor U5174 (N_5174,N_4660,N_4729);
and U5175 (N_5175,N_4786,N_4997);
xor U5176 (N_5176,N_4769,N_4951);
and U5177 (N_5177,N_4669,N_4999);
or U5178 (N_5178,N_4808,N_4570);
nor U5179 (N_5179,N_4894,N_4839);
nor U5180 (N_5180,N_4712,N_4640);
nand U5181 (N_5181,N_4633,N_4835);
or U5182 (N_5182,N_4842,N_4812);
xnor U5183 (N_5183,N_4936,N_4728);
or U5184 (N_5184,N_4533,N_4794);
or U5185 (N_5185,N_4781,N_4674);
nand U5186 (N_5186,N_4884,N_4831);
nor U5187 (N_5187,N_4667,N_4918);
nand U5188 (N_5188,N_4916,N_4590);
or U5189 (N_5189,N_4793,N_4539);
nand U5190 (N_5190,N_4896,N_4650);
or U5191 (N_5191,N_4639,N_4561);
xnor U5192 (N_5192,N_4852,N_4926);
or U5193 (N_5193,N_4589,N_4688);
xor U5194 (N_5194,N_4514,N_4853);
nand U5195 (N_5195,N_4532,N_4575);
and U5196 (N_5196,N_4555,N_4701);
xor U5197 (N_5197,N_4602,N_4651);
or U5198 (N_5198,N_4802,N_4713);
and U5199 (N_5199,N_4944,N_4567);
and U5200 (N_5200,N_4815,N_4773);
xor U5201 (N_5201,N_4863,N_4883);
nand U5202 (N_5202,N_4905,N_4559);
nand U5203 (N_5203,N_4683,N_4734);
nor U5204 (N_5204,N_4714,N_4554);
xnor U5205 (N_5205,N_4930,N_4985);
nor U5206 (N_5206,N_4502,N_4556);
nand U5207 (N_5207,N_4832,N_4745);
nor U5208 (N_5208,N_4766,N_4965);
xor U5209 (N_5209,N_4707,N_4753);
xor U5210 (N_5210,N_4678,N_4695);
or U5211 (N_5211,N_4517,N_4776);
xnor U5212 (N_5212,N_4974,N_4980);
nand U5213 (N_5213,N_4923,N_4757);
xor U5214 (N_5214,N_4518,N_4699);
and U5215 (N_5215,N_4696,N_4952);
xor U5216 (N_5216,N_4551,N_4698);
nand U5217 (N_5217,N_4805,N_4597);
nor U5218 (N_5218,N_4767,N_4900);
nand U5219 (N_5219,N_4515,N_4848);
nand U5220 (N_5220,N_4948,N_4527);
or U5221 (N_5221,N_4809,N_4578);
nor U5222 (N_5222,N_4758,N_4988);
and U5223 (N_5223,N_4752,N_4792);
or U5224 (N_5224,N_4972,N_4843);
nor U5225 (N_5225,N_4810,N_4592);
or U5226 (N_5226,N_4501,N_4801);
nor U5227 (N_5227,N_4803,N_4511);
and U5228 (N_5228,N_4738,N_4608);
and U5229 (N_5229,N_4653,N_4915);
xor U5230 (N_5230,N_4912,N_4549);
or U5231 (N_5231,N_4661,N_4528);
and U5232 (N_5232,N_4605,N_4748);
and U5233 (N_5233,N_4627,N_4591);
nor U5234 (N_5234,N_4971,N_4937);
xor U5235 (N_5235,N_4662,N_4553);
nor U5236 (N_5236,N_4610,N_4871);
and U5237 (N_5237,N_4881,N_4584);
nand U5238 (N_5238,N_4977,N_4603);
nor U5239 (N_5239,N_4953,N_4560);
xnor U5240 (N_5240,N_4569,N_4978);
nand U5241 (N_5241,N_4706,N_4664);
nor U5242 (N_5242,N_4620,N_4927);
or U5243 (N_5243,N_4973,N_4693);
xor U5244 (N_5244,N_4715,N_4869);
xnor U5245 (N_5245,N_4838,N_4500);
nor U5246 (N_5246,N_4791,N_4716);
xnor U5247 (N_5247,N_4981,N_4875);
xor U5248 (N_5248,N_4689,N_4536);
or U5249 (N_5249,N_4817,N_4573);
nor U5250 (N_5250,N_4875,N_4738);
or U5251 (N_5251,N_4665,N_4952);
and U5252 (N_5252,N_4993,N_4570);
or U5253 (N_5253,N_4576,N_4621);
xnor U5254 (N_5254,N_4760,N_4951);
and U5255 (N_5255,N_4823,N_4548);
or U5256 (N_5256,N_4668,N_4710);
nor U5257 (N_5257,N_4824,N_4589);
nor U5258 (N_5258,N_4752,N_4547);
nand U5259 (N_5259,N_4965,N_4753);
nand U5260 (N_5260,N_4790,N_4725);
and U5261 (N_5261,N_4708,N_4862);
or U5262 (N_5262,N_4995,N_4768);
or U5263 (N_5263,N_4931,N_4872);
nor U5264 (N_5264,N_4999,N_4608);
xor U5265 (N_5265,N_4929,N_4776);
or U5266 (N_5266,N_4969,N_4857);
nor U5267 (N_5267,N_4985,N_4850);
xor U5268 (N_5268,N_4783,N_4937);
nor U5269 (N_5269,N_4949,N_4860);
and U5270 (N_5270,N_4955,N_4510);
nand U5271 (N_5271,N_4672,N_4759);
or U5272 (N_5272,N_4691,N_4769);
and U5273 (N_5273,N_4737,N_4859);
xnor U5274 (N_5274,N_4564,N_4981);
nand U5275 (N_5275,N_4787,N_4574);
or U5276 (N_5276,N_4568,N_4869);
nor U5277 (N_5277,N_4884,N_4869);
xnor U5278 (N_5278,N_4529,N_4569);
or U5279 (N_5279,N_4868,N_4808);
or U5280 (N_5280,N_4511,N_4651);
nand U5281 (N_5281,N_4864,N_4775);
and U5282 (N_5282,N_4763,N_4953);
xnor U5283 (N_5283,N_4769,N_4654);
xnor U5284 (N_5284,N_4779,N_4683);
or U5285 (N_5285,N_4709,N_4701);
nor U5286 (N_5286,N_4708,N_4879);
nor U5287 (N_5287,N_4842,N_4658);
nor U5288 (N_5288,N_4955,N_4897);
or U5289 (N_5289,N_4690,N_4610);
nor U5290 (N_5290,N_4974,N_4981);
nor U5291 (N_5291,N_4593,N_4628);
or U5292 (N_5292,N_4685,N_4623);
xor U5293 (N_5293,N_4737,N_4772);
or U5294 (N_5294,N_4861,N_4985);
and U5295 (N_5295,N_4901,N_4943);
xnor U5296 (N_5296,N_4719,N_4944);
and U5297 (N_5297,N_4824,N_4924);
nor U5298 (N_5298,N_4587,N_4962);
xnor U5299 (N_5299,N_4893,N_4989);
nand U5300 (N_5300,N_4657,N_4597);
or U5301 (N_5301,N_4648,N_4981);
xnor U5302 (N_5302,N_4992,N_4731);
nor U5303 (N_5303,N_4744,N_4797);
nor U5304 (N_5304,N_4866,N_4642);
or U5305 (N_5305,N_4945,N_4991);
xnor U5306 (N_5306,N_4814,N_4978);
or U5307 (N_5307,N_4748,N_4757);
xor U5308 (N_5308,N_4817,N_4508);
and U5309 (N_5309,N_4519,N_4895);
nand U5310 (N_5310,N_4627,N_4609);
xor U5311 (N_5311,N_4929,N_4980);
or U5312 (N_5312,N_4938,N_4854);
and U5313 (N_5313,N_4757,N_4640);
and U5314 (N_5314,N_4941,N_4810);
nor U5315 (N_5315,N_4792,N_4886);
nor U5316 (N_5316,N_4806,N_4666);
nor U5317 (N_5317,N_4673,N_4992);
nand U5318 (N_5318,N_4874,N_4771);
nor U5319 (N_5319,N_4864,N_4852);
xnor U5320 (N_5320,N_4944,N_4632);
or U5321 (N_5321,N_4861,N_4522);
or U5322 (N_5322,N_4803,N_4982);
nand U5323 (N_5323,N_4650,N_4866);
or U5324 (N_5324,N_4627,N_4594);
or U5325 (N_5325,N_4512,N_4565);
xnor U5326 (N_5326,N_4756,N_4785);
and U5327 (N_5327,N_4927,N_4629);
or U5328 (N_5328,N_4844,N_4551);
and U5329 (N_5329,N_4503,N_4848);
and U5330 (N_5330,N_4553,N_4668);
and U5331 (N_5331,N_4620,N_4576);
nor U5332 (N_5332,N_4916,N_4730);
or U5333 (N_5333,N_4843,N_4620);
or U5334 (N_5334,N_4775,N_4989);
xor U5335 (N_5335,N_4875,N_4782);
nor U5336 (N_5336,N_4945,N_4652);
xor U5337 (N_5337,N_4980,N_4682);
or U5338 (N_5338,N_4729,N_4949);
nand U5339 (N_5339,N_4910,N_4780);
xor U5340 (N_5340,N_4969,N_4971);
nand U5341 (N_5341,N_4544,N_4721);
xnor U5342 (N_5342,N_4670,N_4839);
xnor U5343 (N_5343,N_4815,N_4721);
xnor U5344 (N_5344,N_4920,N_4623);
nand U5345 (N_5345,N_4769,N_4843);
or U5346 (N_5346,N_4750,N_4675);
or U5347 (N_5347,N_4619,N_4913);
xor U5348 (N_5348,N_4848,N_4828);
nor U5349 (N_5349,N_4693,N_4997);
nand U5350 (N_5350,N_4962,N_4514);
xnor U5351 (N_5351,N_4899,N_4737);
nor U5352 (N_5352,N_4657,N_4998);
and U5353 (N_5353,N_4946,N_4548);
nand U5354 (N_5354,N_4804,N_4617);
nand U5355 (N_5355,N_4542,N_4825);
nor U5356 (N_5356,N_4639,N_4837);
nand U5357 (N_5357,N_4787,N_4963);
or U5358 (N_5358,N_4911,N_4768);
nor U5359 (N_5359,N_4758,N_4718);
or U5360 (N_5360,N_4768,N_4791);
or U5361 (N_5361,N_4746,N_4519);
and U5362 (N_5362,N_4523,N_4975);
xor U5363 (N_5363,N_4864,N_4969);
nor U5364 (N_5364,N_4960,N_4609);
or U5365 (N_5365,N_4976,N_4546);
xnor U5366 (N_5366,N_4731,N_4542);
nand U5367 (N_5367,N_4570,N_4891);
nand U5368 (N_5368,N_4816,N_4566);
xnor U5369 (N_5369,N_4744,N_4569);
nand U5370 (N_5370,N_4707,N_4695);
nand U5371 (N_5371,N_4512,N_4887);
or U5372 (N_5372,N_4868,N_4500);
or U5373 (N_5373,N_4618,N_4814);
or U5374 (N_5374,N_4760,N_4629);
and U5375 (N_5375,N_4634,N_4974);
and U5376 (N_5376,N_4513,N_4681);
nand U5377 (N_5377,N_4813,N_4725);
or U5378 (N_5378,N_4943,N_4810);
xnor U5379 (N_5379,N_4769,N_4889);
xnor U5380 (N_5380,N_4987,N_4927);
or U5381 (N_5381,N_4950,N_4733);
nand U5382 (N_5382,N_4911,N_4942);
or U5383 (N_5383,N_4851,N_4603);
or U5384 (N_5384,N_4858,N_4881);
nand U5385 (N_5385,N_4958,N_4674);
nand U5386 (N_5386,N_4613,N_4803);
or U5387 (N_5387,N_4591,N_4956);
or U5388 (N_5388,N_4743,N_4646);
xnor U5389 (N_5389,N_4965,N_4869);
nor U5390 (N_5390,N_4718,N_4668);
nand U5391 (N_5391,N_4921,N_4962);
and U5392 (N_5392,N_4826,N_4993);
nand U5393 (N_5393,N_4513,N_4658);
nor U5394 (N_5394,N_4770,N_4608);
or U5395 (N_5395,N_4891,N_4758);
nor U5396 (N_5396,N_4831,N_4625);
nand U5397 (N_5397,N_4881,N_4995);
or U5398 (N_5398,N_4817,N_4949);
and U5399 (N_5399,N_4730,N_4812);
nand U5400 (N_5400,N_4650,N_4794);
nand U5401 (N_5401,N_4507,N_4737);
nand U5402 (N_5402,N_4988,N_4573);
nand U5403 (N_5403,N_4877,N_4965);
nand U5404 (N_5404,N_4832,N_4953);
nor U5405 (N_5405,N_4696,N_4699);
and U5406 (N_5406,N_4757,N_4643);
xor U5407 (N_5407,N_4755,N_4856);
nor U5408 (N_5408,N_4974,N_4730);
nand U5409 (N_5409,N_4564,N_4576);
nand U5410 (N_5410,N_4974,N_4624);
or U5411 (N_5411,N_4520,N_4878);
xor U5412 (N_5412,N_4540,N_4594);
xnor U5413 (N_5413,N_4974,N_4940);
or U5414 (N_5414,N_4785,N_4771);
xor U5415 (N_5415,N_4750,N_4843);
and U5416 (N_5416,N_4638,N_4632);
nor U5417 (N_5417,N_4744,N_4559);
or U5418 (N_5418,N_4711,N_4678);
and U5419 (N_5419,N_4799,N_4577);
and U5420 (N_5420,N_4508,N_4979);
and U5421 (N_5421,N_4567,N_4971);
nand U5422 (N_5422,N_4793,N_4794);
xnor U5423 (N_5423,N_4663,N_4959);
or U5424 (N_5424,N_4500,N_4823);
xnor U5425 (N_5425,N_4621,N_4857);
or U5426 (N_5426,N_4657,N_4563);
xnor U5427 (N_5427,N_4536,N_4941);
or U5428 (N_5428,N_4942,N_4598);
xnor U5429 (N_5429,N_4866,N_4909);
xor U5430 (N_5430,N_4570,N_4696);
or U5431 (N_5431,N_4816,N_4660);
and U5432 (N_5432,N_4883,N_4747);
nand U5433 (N_5433,N_4992,N_4609);
or U5434 (N_5434,N_4854,N_4861);
nor U5435 (N_5435,N_4870,N_4588);
nor U5436 (N_5436,N_4894,N_4668);
and U5437 (N_5437,N_4946,N_4972);
xor U5438 (N_5438,N_4864,N_4806);
nand U5439 (N_5439,N_4597,N_4945);
or U5440 (N_5440,N_4552,N_4822);
or U5441 (N_5441,N_4841,N_4524);
xor U5442 (N_5442,N_4667,N_4837);
xnor U5443 (N_5443,N_4665,N_4502);
or U5444 (N_5444,N_4978,N_4597);
or U5445 (N_5445,N_4744,N_4878);
nand U5446 (N_5446,N_4772,N_4547);
nand U5447 (N_5447,N_4915,N_4843);
nand U5448 (N_5448,N_4593,N_4713);
nor U5449 (N_5449,N_4863,N_4678);
nand U5450 (N_5450,N_4801,N_4609);
and U5451 (N_5451,N_4641,N_4555);
xnor U5452 (N_5452,N_4914,N_4878);
or U5453 (N_5453,N_4581,N_4705);
or U5454 (N_5454,N_4703,N_4900);
or U5455 (N_5455,N_4827,N_4522);
nand U5456 (N_5456,N_4962,N_4561);
nor U5457 (N_5457,N_4657,N_4799);
or U5458 (N_5458,N_4868,N_4539);
and U5459 (N_5459,N_4859,N_4975);
nor U5460 (N_5460,N_4660,N_4724);
and U5461 (N_5461,N_4952,N_4736);
and U5462 (N_5462,N_4945,N_4604);
and U5463 (N_5463,N_4627,N_4726);
nor U5464 (N_5464,N_4727,N_4729);
or U5465 (N_5465,N_4534,N_4567);
nand U5466 (N_5466,N_4515,N_4649);
nor U5467 (N_5467,N_4707,N_4963);
or U5468 (N_5468,N_4787,N_4918);
nand U5469 (N_5469,N_4995,N_4892);
nand U5470 (N_5470,N_4616,N_4967);
xnor U5471 (N_5471,N_4892,N_4575);
xor U5472 (N_5472,N_4887,N_4653);
nand U5473 (N_5473,N_4830,N_4735);
or U5474 (N_5474,N_4872,N_4516);
nor U5475 (N_5475,N_4695,N_4680);
and U5476 (N_5476,N_4521,N_4734);
and U5477 (N_5477,N_4639,N_4973);
and U5478 (N_5478,N_4837,N_4651);
nand U5479 (N_5479,N_4529,N_4951);
nor U5480 (N_5480,N_4572,N_4764);
nand U5481 (N_5481,N_4832,N_4721);
nand U5482 (N_5482,N_4916,N_4656);
nor U5483 (N_5483,N_4647,N_4635);
nand U5484 (N_5484,N_4789,N_4649);
nand U5485 (N_5485,N_4531,N_4735);
nor U5486 (N_5486,N_4605,N_4732);
and U5487 (N_5487,N_4795,N_4641);
nor U5488 (N_5488,N_4646,N_4782);
or U5489 (N_5489,N_4971,N_4651);
or U5490 (N_5490,N_4816,N_4828);
nor U5491 (N_5491,N_4881,N_4898);
nor U5492 (N_5492,N_4633,N_4640);
nand U5493 (N_5493,N_4523,N_4533);
nor U5494 (N_5494,N_4813,N_4745);
and U5495 (N_5495,N_4661,N_4724);
nand U5496 (N_5496,N_4947,N_4971);
and U5497 (N_5497,N_4995,N_4794);
xnor U5498 (N_5498,N_4749,N_4672);
and U5499 (N_5499,N_4680,N_4557);
and U5500 (N_5500,N_5143,N_5290);
or U5501 (N_5501,N_5428,N_5295);
and U5502 (N_5502,N_5230,N_5485);
nand U5503 (N_5503,N_5455,N_5311);
xor U5504 (N_5504,N_5426,N_5142);
and U5505 (N_5505,N_5083,N_5403);
nand U5506 (N_5506,N_5364,N_5436);
nor U5507 (N_5507,N_5082,N_5237);
nand U5508 (N_5508,N_5238,N_5487);
nor U5509 (N_5509,N_5366,N_5358);
nand U5510 (N_5510,N_5379,N_5398);
nand U5511 (N_5511,N_5216,N_5175);
or U5512 (N_5512,N_5271,N_5400);
nand U5513 (N_5513,N_5224,N_5367);
nand U5514 (N_5514,N_5039,N_5222);
xnor U5515 (N_5515,N_5460,N_5267);
or U5516 (N_5516,N_5419,N_5458);
and U5517 (N_5517,N_5075,N_5192);
nor U5518 (N_5518,N_5446,N_5088);
or U5519 (N_5519,N_5332,N_5371);
and U5520 (N_5520,N_5242,N_5103);
and U5521 (N_5521,N_5424,N_5063);
xor U5522 (N_5522,N_5359,N_5119);
nor U5523 (N_5523,N_5155,N_5148);
nand U5524 (N_5524,N_5264,N_5244);
or U5525 (N_5525,N_5227,N_5183);
and U5526 (N_5526,N_5125,N_5369);
or U5527 (N_5527,N_5442,N_5262);
or U5528 (N_5528,N_5343,N_5489);
xor U5529 (N_5529,N_5429,N_5173);
and U5530 (N_5530,N_5225,N_5462);
xor U5531 (N_5531,N_5117,N_5065);
and U5532 (N_5532,N_5049,N_5093);
xor U5533 (N_5533,N_5282,N_5395);
nand U5534 (N_5534,N_5029,N_5360);
and U5535 (N_5535,N_5002,N_5010);
nand U5536 (N_5536,N_5060,N_5185);
or U5537 (N_5537,N_5337,N_5381);
nor U5538 (N_5538,N_5272,N_5133);
xor U5539 (N_5539,N_5350,N_5077);
nor U5540 (N_5540,N_5368,N_5132);
or U5541 (N_5541,N_5466,N_5273);
or U5542 (N_5542,N_5461,N_5146);
nand U5543 (N_5543,N_5152,N_5382);
or U5544 (N_5544,N_5416,N_5294);
nand U5545 (N_5545,N_5336,N_5247);
or U5546 (N_5546,N_5048,N_5390);
and U5547 (N_5547,N_5086,N_5300);
nand U5548 (N_5548,N_5085,N_5109);
xor U5549 (N_5549,N_5445,N_5014);
nor U5550 (N_5550,N_5318,N_5313);
or U5551 (N_5551,N_5404,N_5035);
and U5552 (N_5552,N_5432,N_5134);
nand U5553 (N_5553,N_5389,N_5456);
and U5554 (N_5554,N_5101,N_5055);
nor U5555 (N_5555,N_5494,N_5129);
or U5556 (N_5556,N_5087,N_5452);
nand U5557 (N_5557,N_5098,N_5120);
or U5558 (N_5558,N_5321,N_5154);
xor U5559 (N_5559,N_5444,N_5030);
nor U5560 (N_5560,N_5484,N_5316);
nor U5561 (N_5561,N_5032,N_5474);
nand U5562 (N_5562,N_5396,N_5451);
nor U5563 (N_5563,N_5127,N_5160);
nor U5564 (N_5564,N_5195,N_5254);
nor U5565 (N_5565,N_5062,N_5393);
and U5566 (N_5566,N_5205,N_5328);
xor U5567 (N_5567,N_5374,N_5326);
and U5568 (N_5568,N_5165,N_5331);
and U5569 (N_5569,N_5453,N_5415);
nor U5570 (N_5570,N_5301,N_5033);
nand U5571 (N_5571,N_5115,N_5110);
and U5572 (N_5572,N_5181,N_5344);
and U5573 (N_5573,N_5169,N_5219);
nor U5574 (N_5574,N_5402,N_5268);
or U5575 (N_5575,N_5011,N_5009);
nor U5576 (N_5576,N_5199,N_5186);
nand U5577 (N_5577,N_5001,N_5397);
and U5578 (N_5578,N_5182,N_5376);
nand U5579 (N_5579,N_5283,N_5214);
or U5580 (N_5580,N_5138,N_5118);
nor U5581 (N_5581,N_5293,N_5215);
xnor U5582 (N_5582,N_5307,N_5027);
or U5583 (N_5583,N_5433,N_5174);
and U5584 (N_5584,N_5299,N_5399);
nor U5585 (N_5585,N_5236,N_5303);
and U5586 (N_5586,N_5220,N_5347);
or U5587 (N_5587,N_5476,N_5051);
nand U5588 (N_5588,N_5255,N_5380);
nor U5589 (N_5589,N_5208,N_5217);
xnor U5590 (N_5590,N_5486,N_5206);
nand U5591 (N_5591,N_5274,N_5427);
or U5592 (N_5592,N_5228,N_5100);
or U5593 (N_5593,N_5210,N_5161);
nand U5594 (N_5594,N_5090,N_5006);
xnor U5595 (N_5595,N_5412,N_5123);
and U5596 (N_5596,N_5309,N_5018);
xnor U5597 (N_5597,N_5270,N_5322);
xnor U5598 (N_5598,N_5437,N_5067);
xor U5599 (N_5599,N_5354,N_5459);
or U5600 (N_5600,N_5052,N_5166);
xnor U5601 (N_5601,N_5450,N_5481);
xor U5602 (N_5602,N_5031,N_5339);
or U5603 (N_5603,N_5479,N_5340);
xnor U5604 (N_5604,N_5286,N_5207);
or U5605 (N_5605,N_5408,N_5324);
and U5606 (N_5606,N_5187,N_5080);
nor U5607 (N_5607,N_5068,N_5044);
and U5608 (N_5608,N_5259,N_5258);
and U5609 (N_5609,N_5246,N_5095);
nor U5610 (N_5610,N_5266,N_5353);
xor U5611 (N_5611,N_5020,N_5441);
or U5612 (N_5612,N_5047,N_5289);
nor U5613 (N_5613,N_5457,N_5036);
and U5614 (N_5614,N_5064,N_5025);
nand U5615 (N_5615,N_5463,N_5054);
or U5616 (N_5616,N_5305,N_5257);
nor U5617 (N_5617,N_5378,N_5156);
xnor U5618 (N_5618,N_5016,N_5363);
and U5619 (N_5619,N_5245,N_5140);
nor U5620 (N_5620,N_5291,N_5464);
xor U5621 (N_5621,N_5388,N_5172);
xor U5622 (N_5622,N_5356,N_5112);
nand U5623 (N_5623,N_5162,N_5406);
and U5624 (N_5624,N_5059,N_5066);
or U5625 (N_5625,N_5015,N_5202);
xor U5626 (N_5626,N_5285,N_5349);
nor U5627 (N_5627,N_5221,N_5251);
nand U5628 (N_5628,N_5041,N_5443);
xnor U5629 (N_5629,N_5203,N_5385);
xnor U5630 (N_5630,N_5003,N_5361);
and U5631 (N_5631,N_5315,N_5421);
nor U5632 (N_5632,N_5204,N_5078);
nor U5633 (N_5633,N_5200,N_5448);
or U5634 (N_5634,N_5394,N_5284);
or U5635 (N_5635,N_5423,N_5277);
or U5636 (N_5636,N_5212,N_5038);
nand U5637 (N_5637,N_5004,N_5239);
xor U5638 (N_5638,N_5157,N_5298);
nand U5639 (N_5639,N_5113,N_5050);
and U5640 (N_5640,N_5072,N_5334);
nand U5641 (N_5641,N_5076,N_5124);
nand U5642 (N_5642,N_5056,N_5040);
or U5643 (N_5643,N_5126,N_5229);
nor U5644 (N_5644,N_5231,N_5306);
nor U5645 (N_5645,N_5176,N_5482);
or U5646 (N_5646,N_5053,N_5387);
or U5647 (N_5647,N_5330,N_5159);
xor U5648 (N_5648,N_5304,N_5104);
nand U5649 (N_5649,N_5470,N_5116);
xnor U5650 (N_5650,N_5121,N_5495);
xor U5651 (N_5651,N_5308,N_5241);
xnor U5652 (N_5652,N_5407,N_5130);
and U5653 (N_5653,N_5499,N_5073);
and U5654 (N_5654,N_5475,N_5310);
and U5655 (N_5655,N_5269,N_5043);
or U5656 (N_5656,N_5177,N_5420);
nor U5657 (N_5657,N_5136,N_5401);
and U5658 (N_5658,N_5431,N_5278);
or U5659 (N_5659,N_5034,N_5213);
xnor U5660 (N_5660,N_5493,N_5106);
and U5661 (N_5661,N_5471,N_5345);
nor U5662 (N_5662,N_5144,N_5317);
xor U5663 (N_5663,N_5355,N_5197);
or U5664 (N_5664,N_5496,N_5449);
nor U5665 (N_5665,N_5467,N_5000);
xor U5666 (N_5666,N_5352,N_5058);
nand U5667 (N_5667,N_5296,N_5483);
nor U5668 (N_5668,N_5179,N_5440);
xnor U5669 (N_5669,N_5417,N_5097);
nand U5670 (N_5670,N_5386,N_5373);
xor U5671 (N_5671,N_5218,N_5488);
nor U5672 (N_5672,N_5265,N_5434);
xor U5673 (N_5673,N_5365,N_5362);
nand U5674 (N_5674,N_5193,N_5094);
xor U5675 (N_5675,N_5418,N_5131);
nand U5676 (N_5676,N_5105,N_5348);
nand U5677 (N_5677,N_5092,N_5191);
nand U5678 (N_5678,N_5081,N_5492);
and U5679 (N_5679,N_5201,N_5149);
and U5680 (N_5680,N_5026,N_5171);
and U5681 (N_5681,N_5383,N_5249);
and U5682 (N_5682,N_5069,N_5280);
nor U5683 (N_5683,N_5021,N_5107);
nor U5684 (N_5684,N_5335,N_5012);
or U5685 (N_5685,N_5079,N_5276);
and U5686 (N_5686,N_5468,N_5137);
or U5687 (N_5687,N_5430,N_5287);
xnor U5688 (N_5688,N_5375,N_5226);
and U5689 (N_5689,N_5319,N_5384);
and U5690 (N_5690,N_5498,N_5141);
nand U5691 (N_5691,N_5042,N_5045);
nand U5692 (N_5692,N_5410,N_5111);
xnor U5693 (N_5693,N_5454,N_5477);
nor U5694 (N_5694,N_5250,N_5323);
xnor U5695 (N_5695,N_5439,N_5211);
nand U5696 (N_5696,N_5370,N_5252);
nand U5697 (N_5697,N_5235,N_5469);
and U5698 (N_5698,N_5405,N_5114);
and U5699 (N_5699,N_5377,N_5099);
and U5700 (N_5700,N_5473,N_5263);
nor U5701 (N_5701,N_5028,N_5338);
or U5702 (N_5702,N_5178,N_5153);
and U5703 (N_5703,N_5438,N_5122);
nand U5704 (N_5704,N_5346,N_5167);
and U5705 (N_5705,N_5070,N_5071);
xnor U5706 (N_5706,N_5281,N_5102);
nand U5707 (N_5707,N_5435,N_5297);
nor U5708 (N_5708,N_5312,N_5325);
nand U5709 (N_5709,N_5253,N_5413);
or U5710 (N_5710,N_5372,N_5209);
and U5711 (N_5711,N_5279,N_5327);
and U5712 (N_5712,N_5096,N_5008);
xor U5713 (N_5713,N_5411,N_5248);
and U5714 (N_5714,N_5472,N_5168);
nand U5715 (N_5715,N_5163,N_5147);
and U5716 (N_5716,N_5170,N_5314);
nor U5717 (N_5717,N_5333,N_5091);
nand U5718 (N_5718,N_5184,N_5046);
nand U5719 (N_5719,N_5128,N_5261);
xor U5720 (N_5720,N_5158,N_5320);
nor U5721 (N_5721,N_5108,N_5135);
nand U5722 (N_5722,N_5391,N_5357);
nand U5723 (N_5723,N_5022,N_5232);
xor U5724 (N_5724,N_5233,N_5414);
and U5725 (N_5725,N_5190,N_5422);
or U5726 (N_5726,N_5409,N_5341);
and U5727 (N_5727,N_5139,N_5240);
xor U5728 (N_5728,N_5491,N_5005);
and U5729 (N_5729,N_5275,N_5013);
nor U5730 (N_5730,N_5061,N_5302);
xor U5731 (N_5731,N_5198,N_5196);
xor U5732 (N_5732,N_5164,N_5342);
and U5733 (N_5733,N_5084,N_5188);
or U5734 (N_5734,N_5425,N_5194);
and U5735 (N_5735,N_5260,N_5074);
xor U5736 (N_5736,N_5490,N_5256);
xnor U5737 (N_5737,N_5007,N_5189);
nor U5738 (N_5738,N_5480,N_5351);
and U5739 (N_5739,N_5023,N_5288);
nand U5740 (N_5740,N_5234,N_5223);
and U5741 (N_5741,N_5243,N_5329);
or U5742 (N_5742,N_5037,N_5478);
nor U5743 (N_5743,N_5057,N_5180);
nor U5744 (N_5744,N_5024,N_5089);
xnor U5745 (N_5745,N_5447,N_5392);
nand U5746 (N_5746,N_5017,N_5465);
xnor U5747 (N_5747,N_5497,N_5150);
nand U5748 (N_5748,N_5145,N_5019);
xnor U5749 (N_5749,N_5151,N_5292);
and U5750 (N_5750,N_5126,N_5262);
nor U5751 (N_5751,N_5408,N_5148);
or U5752 (N_5752,N_5045,N_5221);
nor U5753 (N_5753,N_5131,N_5410);
or U5754 (N_5754,N_5355,N_5089);
xnor U5755 (N_5755,N_5494,N_5032);
nor U5756 (N_5756,N_5263,N_5018);
nand U5757 (N_5757,N_5330,N_5145);
nand U5758 (N_5758,N_5035,N_5189);
or U5759 (N_5759,N_5122,N_5425);
or U5760 (N_5760,N_5027,N_5478);
nor U5761 (N_5761,N_5073,N_5018);
or U5762 (N_5762,N_5051,N_5334);
and U5763 (N_5763,N_5289,N_5113);
nor U5764 (N_5764,N_5431,N_5003);
or U5765 (N_5765,N_5318,N_5069);
and U5766 (N_5766,N_5273,N_5193);
or U5767 (N_5767,N_5214,N_5103);
xnor U5768 (N_5768,N_5446,N_5340);
and U5769 (N_5769,N_5345,N_5222);
nand U5770 (N_5770,N_5146,N_5314);
nand U5771 (N_5771,N_5392,N_5231);
and U5772 (N_5772,N_5498,N_5107);
nor U5773 (N_5773,N_5012,N_5259);
and U5774 (N_5774,N_5196,N_5253);
or U5775 (N_5775,N_5176,N_5134);
xnor U5776 (N_5776,N_5497,N_5054);
xnor U5777 (N_5777,N_5007,N_5157);
nand U5778 (N_5778,N_5431,N_5178);
and U5779 (N_5779,N_5045,N_5199);
and U5780 (N_5780,N_5276,N_5054);
nand U5781 (N_5781,N_5179,N_5160);
nand U5782 (N_5782,N_5115,N_5108);
xor U5783 (N_5783,N_5377,N_5013);
or U5784 (N_5784,N_5457,N_5298);
or U5785 (N_5785,N_5308,N_5493);
nor U5786 (N_5786,N_5310,N_5397);
and U5787 (N_5787,N_5042,N_5382);
and U5788 (N_5788,N_5111,N_5344);
nand U5789 (N_5789,N_5438,N_5262);
nor U5790 (N_5790,N_5274,N_5230);
and U5791 (N_5791,N_5406,N_5438);
xor U5792 (N_5792,N_5060,N_5485);
xor U5793 (N_5793,N_5001,N_5131);
nor U5794 (N_5794,N_5231,N_5005);
nand U5795 (N_5795,N_5427,N_5119);
xnor U5796 (N_5796,N_5014,N_5178);
xnor U5797 (N_5797,N_5397,N_5481);
xor U5798 (N_5798,N_5300,N_5438);
and U5799 (N_5799,N_5328,N_5130);
xnor U5800 (N_5800,N_5434,N_5411);
nand U5801 (N_5801,N_5475,N_5391);
nand U5802 (N_5802,N_5442,N_5450);
nand U5803 (N_5803,N_5161,N_5241);
xor U5804 (N_5804,N_5076,N_5448);
nor U5805 (N_5805,N_5205,N_5422);
nor U5806 (N_5806,N_5375,N_5491);
nor U5807 (N_5807,N_5177,N_5433);
xnor U5808 (N_5808,N_5131,N_5076);
or U5809 (N_5809,N_5252,N_5011);
xor U5810 (N_5810,N_5379,N_5417);
and U5811 (N_5811,N_5132,N_5238);
nor U5812 (N_5812,N_5040,N_5455);
or U5813 (N_5813,N_5115,N_5070);
or U5814 (N_5814,N_5160,N_5002);
xor U5815 (N_5815,N_5458,N_5243);
xor U5816 (N_5816,N_5222,N_5371);
or U5817 (N_5817,N_5336,N_5105);
nand U5818 (N_5818,N_5308,N_5180);
nand U5819 (N_5819,N_5230,N_5308);
xor U5820 (N_5820,N_5148,N_5371);
and U5821 (N_5821,N_5054,N_5305);
xor U5822 (N_5822,N_5465,N_5095);
nand U5823 (N_5823,N_5192,N_5084);
or U5824 (N_5824,N_5051,N_5372);
and U5825 (N_5825,N_5422,N_5049);
xnor U5826 (N_5826,N_5278,N_5418);
or U5827 (N_5827,N_5327,N_5487);
nand U5828 (N_5828,N_5446,N_5300);
xnor U5829 (N_5829,N_5174,N_5341);
nand U5830 (N_5830,N_5146,N_5116);
and U5831 (N_5831,N_5470,N_5362);
xnor U5832 (N_5832,N_5025,N_5403);
nand U5833 (N_5833,N_5438,N_5446);
xnor U5834 (N_5834,N_5195,N_5274);
nand U5835 (N_5835,N_5203,N_5265);
and U5836 (N_5836,N_5347,N_5445);
xnor U5837 (N_5837,N_5299,N_5157);
xor U5838 (N_5838,N_5165,N_5477);
nand U5839 (N_5839,N_5156,N_5070);
xor U5840 (N_5840,N_5292,N_5185);
and U5841 (N_5841,N_5235,N_5447);
nand U5842 (N_5842,N_5146,N_5413);
xor U5843 (N_5843,N_5076,N_5252);
and U5844 (N_5844,N_5306,N_5204);
xnor U5845 (N_5845,N_5188,N_5146);
nor U5846 (N_5846,N_5444,N_5075);
nor U5847 (N_5847,N_5074,N_5275);
xor U5848 (N_5848,N_5276,N_5226);
nand U5849 (N_5849,N_5361,N_5062);
nand U5850 (N_5850,N_5317,N_5208);
nand U5851 (N_5851,N_5081,N_5406);
xor U5852 (N_5852,N_5051,N_5468);
nor U5853 (N_5853,N_5156,N_5005);
and U5854 (N_5854,N_5394,N_5280);
xor U5855 (N_5855,N_5278,N_5268);
nor U5856 (N_5856,N_5321,N_5322);
nor U5857 (N_5857,N_5030,N_5122);
xnor U5858 (N_5858,N_5447,N_5048);
nor U5859 (N_5859,N_5219,N_5099);
nand U5860 (N_5860,N_5382,N_5468);
nand U5861 (N_5861,N_5170,N_5222);
nand U5862 (N_5862,N_5007,N_5323);
nor U5863 (N_5863,N_5009,N_5245);
nor U5864 (N_5864,N_5039,N_5282);
or U5865 (N_5865,N_5315,N_5115);
or U5866 (N_5866,N_5440,N_5299);
nand U5867 (N_5867,N_5084,N_5028);
nand U5868 (N_5868,N_5322,N_5212);
nor U5869 (N_5869,N_5443,N_5400);
and U5870 (N_5870,N_5321,N_5092);
nor U5871 (N_5871,N_5102,N_5077);
xor U5872 (N_5872,N_5341,N_5007);
xnor U5873 (N_5873,N_5317,N_5034);
xnor U5874 (N_5874,N_5019,N_5373);
nand U5875 (N_5875,N_5368,N_5181);
nand U5876 (N_5876,N_5023,N_5155);
nor U5877 (N_5877,N_5219,N_5168);
nor U5878 (N_5878,N_5036,N_5423);
or U5879 (N_5879,N_5211,N_5491);
and U5880 (N_5880,N_5376,N_5320);
nor U5881 (N_5881,N_5294,N_5269);
and U5882 (N_5882,N_5227,N_5284);
nor U5883 (N_5883,N_5311,N_5481);
and U5884 (N_5884,N_5465,N_5076);
or U5885 (N_5885,N_5333,N_5497);
and U5886 (N_5886,N_5336,N_5442);
xor U5887 (N_5887,N_5400,N_5423);
nor U5888 (N_5888,N_5254,N_5343);
nand U5889 (N_5889,N_5396,N_5119);
nand U5890 (N_5890,N_5041,N_5347);
nor U5891 (N_5891,N_5207,N_5497);
xor U5892 (N_5892,N_5011,N_5283);
and U5893 (N_5893,N_5292,N_5453);
or U5894 (N_5894,N_5374,N_5030);
and U5895 (N_5895,N_5218,N_5377);
nand U5896 (N_5896,N_5024,N_5446);
xor U5897 (N_5897,N_5100,N_5294);
nand U5898 (N_5898,N_5362,N_5084);
and U5899 (N_5899,N_5252,N_5024);
nand U5900 (N_5900,N_5211,N_5278);
nor U5901 (N_5901,N_5244,N_5141);
nor U5902 (N_5902,N_5135,N_5123);
or U5903 (N_5903,N_5453,N_5444);
nor U5904 (N_5904,N_5119,N_5050);
or U5905 (N_5905,N_5053,N_5072);
nand U5906 (N_5906,N_5347,N_5414);
xnor U5907 (N_5907,N_5227,N_5015);
or U5908 (N_5908,N_5458,N_5352);
nand U5909 (N_5909,N_5135,N_5311);
xnor U5910 (N_5910,N_5050,N_5085);
and U5911 (N_5911,N_5175,N_5091);
nand U5912 (N_5912,N_5058,N_5131);
nor U5913 (N_5913,N_5330,N_5087);
xnor U5914 (N_5914,N_5475,N_5454);
or U5915 (N_5915,N_5272,N_5412);
nor U5916 (N_5916,N_5377,N_5199);
xnor U5917 (N_5917,N_5412,N_5215);
or U5918 (N_5918,N_5274,N_5042);
and U5919 (N_5919,N_5119,N_5220);
xor U5920 (N_5920,N_5077,N_5272);
xnor U5921 (N_5921,N_5380,N_5348);
xnor U5922 (N_5922,N_5422,N_5385);
or U5923 (N_5923,N_5497,N_5384);
nor U5924 (N_5924,N_5168,N_5463);
nor U5925 (N_5925,N_5346,N_5383);
nor U5926 (N_5926,N_5349,N_5256);
or U5927 (N_5927,N_5462,N_5001);
and U5928 (N_5928,N_5144,N_5379);
or U5929 (N_5929,N_5421,N_5454);
nand U5930 (N_5930,N_5340,N_5430);
and U5931 (N_5931,N_5111,N_5063);
or U5932 (N_5932,N_5113,N_5348);
or U5933 (N_5933,N_5444,N_5308);
or U5934 (N_5934,N_5244,N_5358);
or U5935 (N_5935,N_5478,N_5290);
xnor U5936 (N_5936,N_5115,N_5287);
nand U5937 (N_5937,N_5401,N_5058);
or U5938 (N_5938,N_5371,N_5011);
xnor U5939 (N_5939,N_5259,N_5280);
or U5940 (N_5940,N_5454,N_5374);
nor U5941 (N_5941,N_5279,N_5173);
nor U5942 (N_5942,N_5048,N_5153);
xor U5943 (N_5943,N_5355,N_5264);
nor U5944 (N_5944,N_5429,N_5270);
or U5945 (N_5945,N_5430,N_5475);
nor U5946 (N_5946,N_5143,N_5012);
and U5947 (N_5947,N_5359,N_5411);
or U5948 (N_5948,N_5252,N_5175);
xnor U5949 (N_5949,N_5184,N_5487);
xnor U5950 (N_5950,N_5348,N_5415);
nand U5951 (N_5951,N_5307,N_5044);
or U5952 (N_5952,N_5359,N_5230);
xor U5953 (N_5953,N_5116,N_5353);
nand U5954 (N_5954,N_5346,N_5382);
nor U5955 (N_5955,N_5425,N_5069);
nor U5956 (N_5956,N_5335,N_5030);
and U5957 (N_5957,N_5200,N_5381);
or U5958 (N_5958,N_5370,N_5238);
or U5959 (N_5959,N_5073,N_5145);
xor U5960 (N_5960,N_5098,N_5203);
xnor U5961 (N_5961,N_5375,N_5352);
nand U5962 (N_5962,N_5246,N_5458);
xnor U5963 (N_5963,N_5168,N_5444);
and U5964 (N_5964,N_5213,N_5284);
and U5965 (N_5965,N_5116,N_5435);
nand U5966 (N_5966,N_5373,N_5008);
or U5967 (N_5967,N_5173,N_5211);
nand U5968 (N_5968,N_5259,N_5043);
or U5969 (N_5969,N_5460,N_5094);
nor U5970 (N_5970,N_5287,N_5033);
and U5971 (N_5971,N_5197,N_5432);
and U5972 (N_5972,N_5340,N_5173);
or U5973 (N_5973,N_5316,N_5371);
nand U5974 (N_5974,N_5145,N_5010);
or U5975 (N_5975,N_5320,N_5488);
xor U5976 (N_5976,N_5483,N_5096);
xnor U5977 (N_5977,N_5139,N_5155);
nand U5978 (N_5978,N_5465,N_5186);
and U5979 (N_5979,N_5495,N_5024);
or U5980 (N_5980,N_5250,N_5473);
and U5981 (N_5981,N_5478,N_5008);
nor U5982 (N_5982,N_5387,N_5149);
or U5983 (N_5983,N_5032,N_5081);
and U5984 (N_5984,N_5226,N_5365);
nor U5985 (N_5985,N_5056,N_5416);
or U5986 (N_5986,N_5163,N_5035);
or U5987 (N_5987,N_5243,N_5074);
nand U5988 (N_5988,N_5163,N_5305);
nor U5989 (N_5989,N_5496,N_5084);
xor U5990 (N_5990,N_5026,N_5456);
and U5991 (N_5991,N_5297,N_5020);
xor U5992 (N_5992,N_5142,N_5445);
or U5993 (N_5993,N_5061,N_5320);
nor U5994 (N_5994,N_5459,N_5375);
xor U5995 (N_5995,N_5253,N_5000);
or U5996 (N_5996,N_5041,N_5094);
and U5997 (N_5997,N_5483,N_5191);
xnor U5998 (N_5998,N_5095,N_5266);
xnor U5999 (N_5999,N_5045,N_5411);
nor U6000 (N_6000,N_5930,N_5500);
nor U6001 (N_6001,N_5835,N_5876);
xor U6002 (N_6002,N_5808,N_5526);
nor U6003 (N_6003,N_5965,N_5867);
nand U6004 (N_6004,N_5865,N_5860);
nand U6005 (N_6005,N_5823,N_5825);
nor U6006 (N_6006,N_5506,N_5810);
or U6007 (N_6007,N_5912,N_5542);
xor U6008 (N_6008,N_5780,N_5770);
or U6009 (N_6009,N_5661,N_5693);
xor U6010 (N_6010,N_5749,N_5772);
nor U6011 (N_6011,N_5667,N_5826);
and U6012 (N_6012,N_5995,N_5522);
or U6013 (N_6013,N_5901,N_5634);
nand U6014 (N_6014,N_5552,N_5791);
nor U6015 (N_6015,N_5978,N_5730);
nor U6016 (N_6016,N_5723,N_5899);
nor U6017 (N_6017,N_5537,N_5747);
or U6018 (N_6018,N_5902,N_5805);
or U6019 (N_6019,N_5685,N_5960);
and U6020 (N_6020,N_5618,N_5888);
nor U6021 (N_6021,N_5656,N_5696);
and U6022 (N_6022,N_5907,N_5962);
nor U6023 (N_6023,N_5933,N_5520);
or U6024 (N_6024,N_5732,N_5528);
or U6025 (N_6025,N_5869,N_5561);
nand U6026 (N_6026,N_5556,N_5894);
nor U6027 (N_6027,N_5841,N_5569);
and U6028 (N_6028,N_5690,N_5983);
nand U6029 (N_6029,N_5640,N_5748);
or U6030 (N_6030,N_5813,N_5928);
nor U6031 (N_6031,N_5776,N_5824);
nand U6032 (N_6032,N_5982,N_5967);
xor U6033 (N_6033,N_5775,N_5757);
and U6034 (N_6034,N_5535,N_5692);
nor U6035 (N_6035,N_5746,N_5647);
and U6036 (N_6036,N_5670,N_5992);
xor U6037 (N_6037,N_5855,N_5553);
and U6038 (N_6038,N_5501,N_5691);
and U6039 (N_6039,N_5760,N_5633);
nor U6040 (N_6040,N_5873,N_5815);
nor U6041 (N_6041,N_5905,N_5991);
and U6042 (N_6042,N_5650,N_5801);
xnor U6043 (N_6043,N_5517,N_5559);
or U6044 (N_6044,N_5931,N_5877);
xor U6045 (N_6045,N_5684,N_5726);
and U6046 (N_6046,N_5927,N_5729);
or U6047 (N_6047,N_5508,N_5716);
nand U6048 (N_6048,N_5623,N_5534);
and U6049 (N_6049,N_5733,N_5602);
or U6050 (N_6050,N_5703,N_5745);
and U6051 (N_6051,N_5679,N_5792);
nand U6052 (N_6052,N_5574,N_5900);
nand U6053 (N_6053,N_5799,N_5505);
nand U6054 (N_6054,N_5840,N_5822);
nor U6055 (N_6055,N_5663,N_5964);
xor U6056 (N_6056,N_5645,N_5849);
xnor U6057 (N_6057,N_5625,N_5707);
nand U6058 (N_6058,N_5611,N_5953);
and U6059 (N_6059,N_5934,N_5919);
xnor U6060 (N_6060,N_5916,N_5641);
or U6061 (N_6061,N_5655,N_5728);
and U6062 (N_6062,N_5794,N_5986);
xnor U6063 (N_6063,N_5845,N_5563);
nor U6064 (N_6064,N_5713,N_5543);
xor U6065 (N_6065,N_5999,N_5853);
and U6066 (N_6066,N_5512,N_5642);
nor U6067 (N_6067,N_5756,N_5584);
nand U6068 (N_6068,N_5949,N_5632);
xnor U6069 (N_6069,N_5718,N_5544);
or U6070 (N_6070,N_5887,N_5631);
or U6071 (N_6071,N_5509,N_5638);
and U6072 (N_6072,N_5752,N_5886);
nand U6073 (N_6073,N_5596,N_5626);
nand U6074 (N_6074,N_5976,N_5959);
nor U6075 (N_6075,N_5737,N_5968);
or U6076 (N_6076,N_5809,N_5669);
xor U6077 (N_6077,N_5938,N_5981);
or U6078 (N_6078,N_5606,N_5697);
nor U6079 (N_6079,N_5832,N_5654);
nor U6080 (N_6080,N_5781,N_5831);
or U6081 (N_6081,N_5778,N_5513);
or U6082 (N_6082,N_5514,N_5954);
nand U6083 (N_6083,N_5951,N_5699);
nor U6084 (N_6084,N_5795,N_5765);
and U6085 (N_6085,N_5568,N_5593);
or U6086 (N_6086,N_5751,N_5687);
nor U6087 (N_6087,N_5635,N_5947);
and U6088 (N_6088,N_5646,N_5578);
or U6089 (N_6089,N_5767,N_5896);
or U6090 (N_6090,N_5777,N_5811);
nand U6091 (N_6091,N_5936,N_5895);
nor U6092 (N_6092,N_5579,N_5963);
nor U6093 (N_6093,N_5892,N_5711);
or U6094 (N_6094,N_5893,N_5980);
or U6095 (N_6095,N_5612,N_5782);
xnor U6096 (N_6096,N_5819,N_5616);
nand U6097 (N_6097,N_5603,N_5935);
and U6098 (N_6098,N_5989,N_5750);
nand U6099 (N_6099,N_5743,N_5678);
and U6100 (N_6100,N_5830,N_5939);
xnor U6101 (N_6101,N_5725,N_5820);
nor U6102 (N_6102,N_5977,N_5871);
or U6103 (N_6103,N_5613,N_5779);
nor U6104 (N_6104,N_5605,N_5624);
or U6105 (N_6105,N_5839,N_5971);
nor U6106 (N_6106,N_5628,N_5769);
nand U6107 (N_6107,N_5838,N_5619);
nor U6108 (N_6108,N_5940,N_5878);
nand U6109 (N_6109,N_5666,N_5975);
nor U6110 (N_6110,N_5979,N_5904);
and U6111 (N_6111,N_5861,N_5852);
or U6112 (N_6112,N_5507,N_5829);
or U6113 (N_6113,N_5538,N_5648);
or U6114 (N_6114,N_5798,N_5575);
and U6115 (N_6115,N_5994,N_5620);
xor U6116 (N_6116,N_5818,N_5547);
nand U6117 (N_6117,N_5758,N_5681);
xor U6118 (N_6118,N_5741,N_5583);
and U6119 (N_6119,N_5848,N_5519);
and U6120 (N_6120,N_5662,N_5854);
nor U6121 (N_6121,N_5555,N_5680);
or U6122 (N_6122,N_5639,N_5889);
nor U6123 (N_6123,N_5636,N_5615);
and U6124 (N_6124,N_5683,N_5511);
nand U6125 (N_6125,N_5875,N_5870);
nand U6126 (N_6126,N_5571,N_5796);
and U6127 (N_6127,N_5708,N_5577);
or U6128 (N_6128,N_5665,N_5945);
nand U6129 (N_6129,N_5806,N_5521);
and U6130 (N_6130,N_5570,N_5759);
nor U6131 (N_6131,N_5533,N_5793);
nand U6132 (N_6132,N_5701,N_5503);
xnor U6133 (N_6133,N_5993,N_5937);
nor U6134 (N_6134,N_5609,N_5597);
nand U6135 (N_6135,N_5686,N_5958);
nor U6136 (N_6136,N_5859,N_5689);
nor U6137 (N_6137,N_5649,N_5607);
nor U6138 (N_6138,N_5785,N_5744);
or U6139 (N_6139,N_5972,N_5948);
nand U6140 (N_6140,N_5688,N_5952);
and U6141 (N_6141,N_5846,N_5973);
xnor U6142 (N_6142,N_5531,N_5910);
nor U6143 (N_6143,N_5600,N_5722);
nand U6144 (N_6144,N_5591,N_5572);
nor U6145 (N_6145,N_5890,N_5518);
and U6146 (N_6146,N_5807,N_5786);
nand U6147 (N_6147,N_5643,N_5816);
nor U6148 (N_6148,N_5885,N_5550);
xor U6149 (N_6149,N_5671,N_5587);
or U6150 (N_6150,N_5814,N_5714);
nand U6151 (N_6151,N_5585,N_5709);
and U6152 (N_6152,N_5724,N_5630);
xnor U6153 (N_6153,N_5515,N_5863);
or U6154 (N_6154,N_5712,N_5546);
xnor U6155 (N_6155,N_5704,N_5657);
or U6156 (N_6156,N_5944,N_5987);
xor U6157 (N_6157,N_5644,N_5943);
nor U6158 (N_6158,N_5906,N_5766);
nand U6159 (N_6159,N_5851,N_5592);
xor U6160 (N_6160,N_5803,N_5549);
xnor U6161 (N_6161,N_5755,N_5560);
xnor U6162 (N_6162,N_5788,N_5998);
nor U6163 (N_6163,N_5957,N_5817);
and U6164 (N_6164,N_5874,N_5719);
and U6165 (N_6165,N_5698,N_5921);
and U6166 (N_6166,N_5768,N_5946);
xor U6167 (N_6167,N_5588,N_5567);
nand U6168 (N_6168,N_5834,N_5598);
nand U6169 (N_6169,N_5627,N_5705);
xor U6170 (N_6170,N_5674,N_5797);
nand U6171 (N_6171,N_5926,N_5844);
xnor U6172 (N_6172,N_5884,N_5727);
or U6173 (N_6173,N_5675,N_5922);
nand U6174 (N_6174,N_5984,N_5883);
and U6175 (N_6175,N_5622,N_5988);
xor U6176 (N_6176,N_5653,N_5558);
or U6177 (N_6177,N_5610,N_5706);
nand U6178 (N_6178,N_5918,N_5858);
nor U6179 (N_6179,N_5710,N_5827);
and U6180 (N_6180,N_5763,N_5668);
xnor U6181 (N_6181,N_5909,N_5908);
nand U6182 (N_6182,N_5771,N_5586);
and U6183 (N_6183,N_5997,N_5557);
nand U6184 (N_6184,N_5738,N_5527);
and U6185 (N_6185,N_5897,N_5614);
xor U6186 (N_6186,N_5721,N_5659);
xor U6187 (N_6187,N_5955,N_5651);
or U6188 (N_6188,N_5784,N_5545);
or U6189 (N_6189,N_5565,N_5966);
and U6190 (N_6190,N_5695,N_5974);
xnor U6191 (N_6191,N_5736,N_5821);
nor U6192 (N_6192,N_5595,N_5842);
or U6193 (N_6193,N_5608,N_5637);
nor U6194 (N_6194,N_5594,N_5864);
nand U6195 (N_6195,N_5925,N_5857);
nor U6196 (N_6196,N_5720,N_5911);
nand U6197 (N_6197,N_5554,N_5540);
and U6198 (N_6198,N_5802,N_5790);
xor U6199 (N_6199,N_5682,N_5516);
and U6200 (N_6200,N_5970,N_5532);
nor U6201 (N_6201,N_5694,N_5836);
nand U6202 (N_6202,N_5879,N_5621);
nor U6203 (N_6203,N_5917,N_5920);
xor U6204 (N_6204,N_5580,N_5856);
or U6205 (N_6205,N_5862,N_5996);
nor U6206 (N_6206,N_5739,N_5812);
or U6207 (N_6207,N_5702,N_5504);
nor U6208 (N_6208,N_5941,N_5589);
or U6209 (N_6209,N_5617,N_5833);
or U6210 (N_6210,N_5753,N_5658);
xor U6211 (N_6211,N_5581,N_5789);
or U6212 (N_6212,N_5664,N_5898);
nor U6213 (N_6213,N_5525,N_5562);
and U6214 (N_6214,N_5956,N_5881);
nor U6215 (N_6215,N_5676,N_5915);
nand U6216 (N_6216,N_5715,N_5573);
and U6217 (N_6217,N_5800,N_5660);
nor U6218 (N_6218,N_5843,N_5740);
or U6219 (N_6219,N_5564,N_5524);
xnor U6220 (N_6220,N_5903,N_5523);
nor U6221 (N_6221,N_5783,N_5929);
nor U6222 (N_6222,N_5985,N_5891);
or U6223 (N_6223,N_5590,N_5541);
or U6224 (N_6224,N_5731,N_5990);
or U6225 (N_6225,N_5762,N_5551);
nor U6226 (N_6226,N_5828,N_5672);
or U6227 (N_6227,N_5868,N_5804);
xnor U6228 (N_6228,N_5529,N_5582);
xnor U6229 (N_6229,N_5761,N_5764);
or U6230 (N_6230,N_5913,N_5961);
or U6231 (N_6231,N_5950,N_5774);
or U6232 (N_6232,N_5742,N_5734);
nand U6233 (N_6233,N_5652,N_5872);
nor U6234 (N_6234,N_5882,N_5787);
and U6235 (N_6235,N_5866,N_5837);
xnor U6236 (N_6236,N_5850,N_5914);
and U6237 (N_6237,N_5539,N_5754);
or U6238 (N_6238,N_5629,N_5548);
and U6239 (N_6239,N_5677,N_5673);
or U6240 (N_6240,N_5880,N_5717);
nand U6241 (N_6241,N_5502,N_5942);
or U6242 (N_6242,N_5510,N_5604);
and U6243 (N_6243,N_5536,N_5735);
nand U6244 (N_6244,N_5932,N_5924);
or U6245 (N_6245,N_5923,N_5566);
or U6246 (N_6246,N_5700,N_5601);
nand U6247 (N_6247,N_5773,N_5530);
and U6248 (N_6248,N_5847,N_5576);
and U6249 (N_6249,N_5969,N_5599);
nand U6250 (N_6250,N_5866,N_5682);
or U6251 (N_6251,N_5794,N_5868);
nand U6252 (N_6252,N_5649,N_5669);
or U6253 (N_6253,N_5641,N_5953);
xor U6254 (N_6254,N_5527,N_5730);
and U6255 (N_6255,N_5577,N_5947);
nand U6256 (N_6256,N_5880,N_5710);
or U6257 (N_6257,N_5664,N_5962);
xnor U6258 (N_6258,N_5989,N_5521);
nor U6259 (N_6259,N_5801,N_5722);
and U6260 (N_6260,N_5593,N_5523);
nand U6261 (N_6261,N_5856,N_5596);
xnor U6262 (N_6262,N_5547,N_5762);
xor U6263 (N_6263,N_5984,N_5567);
and U6264 (N_6264,N_5586,N_5642);
and U6265 (N_6265,N_5882,N_5747);
and U6266 (N_6266,N_5989,N_5715);
or U6267 (N_6267,N_5554,N_5603);
nand U6268 (N_6268,N_5901,N_5833);
or U6269 (N_6269,N_5630,N_5772);
xnor U6270 (N_6270,N_5729,N_5887);
and U6271 (N_6271,N_5916,N_5853);
nor U6272 (N_6272,N_5647,N_5992);
nand U6273 (N_6273,N_5988,N_5784);
xnor U6274 (N_6274,N_5674,N_5625);
nor U6275 (N_6275,N_5823,N_5867);
nor U6276 (N_6276,N_5509,N_5883);
and U6277 (N_6277,N_5721,N_5511);
nand U6278 (N_6278,N_5716,N_5975);
nor U6279 (N_6279,N_5905,N_5868);
and U6280 (N_6280,N_5819,N_5519);
or U6281 (N_6281,N_5703,N_5540);
nor U6282 (N_6282,N_5648,N_5740);
and U6283 (N_6283,N_5927,N_5619);
nor U6284 (N_6284,N_5663,N_5662);
nor U6285 (N_6285,N_5522,N_5519);
xor U6286 (N_6286,N_5608,N_5590);
or U6287 (N_6287,N_5688,N_5781);
nand U6288 (N_6288,N_5590,N_5506);
nand U6289 (N_6289,N_5618,N_5584);
xor U6290 (N_6290,N_5653,N_5554);
nor U6291 (N_6291,N_5996,N_5557);
and U6292 (N_6292,N_5842,N_5559);
or U6293 (N_6293,N_5728,N_5517);
nand U6294 (N_6294,N_5652,N_5608);
xnor U6295 (N_6295,N_5977,N_5834);
nand U6296 (N_6296,N_5824,N_5585);
or U6297 (N_6297,N_5821,N_5962);
or U6298 (N_6298,N_5517,N_5883);
nand U6299 (N_6299,N_5547,N_5730);
nor U6300 (N_6300,N_5632,N_5692);
xor U6301 (N_6301,N_5979,N_5796);
nor U6302 (N_6302,N_5535,N_5677);
and U6303 (N_6303,N_5612,N_5895);
and U6304 (N_6304,N_5954,N_5733);
and U6305 (N_6305,N_5509,N_5783);
xor U6306 (N_6306,N_5678,N_5763);
nand U6307 (N_6307,N_5595,N_5661);
nand U6308 (N_6308,N_5828,N_5601);
xor U6309 (N_6309,N_5743,N_5703);
nor U6310 (N_6310,N_5840,N_5512);
and U6311 (N_6311,N_5798,N_5720);
or U6312 (N_6312,N_5991,N_5801);
xor U6313 (N_6313,N_5795,N_5523);
xnor U6314 (N_6314,N_5655,N_5890);
xor U6315 (N_6315,N_5708,N_5526);
xor U6316 (N_6316,N_5824,N_5723);
and U6317 (N_6317,N_5775,N_5505);
or U6318 (N_6318,N_5891,N_5677);
nor U6319 (N_6319,N_5566,N_5823);
nand U6320 (N_6320,N_5838,N_5865);
or U6321 (N_6321,N_5881,N_5972);
and U6322 (N_6322,N_5790,N_5518);
nor U6323 (N_6323,N_5646,N_5650);
and U6324 (N_6324,N_5750,N_5683);
xor U6325 (N_6325,N_5607,N_5825);
nand U6326 (N_6326,N_5659,N_5584);
and U6327 (N_6327,N_5898,N_5531);
or U6328 (N_6328,N_5898,N_5783);
or U6329 (N_6329,N_5624,N_5826);
or U6330 (N_6330,N_5537,N_5580);
xnor U6331 (N_6331,N_5523,N_5835);
or U6332 (N_6332,N_5804,N_5954);
xnor U6333 (N_6333,N_5929,N_5955);
nor U6334 (N_6334,N_5972,N_5903);
nor U6335 (N_6335,N_5526,N_5919);
or U6336 (N_6336,N_5703,N_5794);
or U6337 (N_6337,N_5535,N_5588);
nor U6338 (N_6338,N_5714,N_5556);
nor U6339 (N_6339,N_5752,N_5610);
nand U6340 (N_6340,N_5750,N_5912);
xor U6341 (N_6341,N_5932,N_5516);
or U6342 (N_6342,N_5832,N_5734);
nand U6343 (N_6343,N_5714,N_5529);
or U6344 (N_6344,N_5652,N_5532);
xor U6345 (N_6345,N_5813,N_5671);
xor U6346 (N_6346,N_5571,N_5833);
and U6347 (N_6347,N_5865,N_5524);
nand U6348 (N_6348,N_5862,N_5737);
xor U6349 (N_6349,N_5583,N_5668);
xor U6350 (N_6350,N_5754,N_5519);
nor U6351 (N_6351,N_5952,N_5915);
xor U6352 (N_6352,N_5994,N_5986);
nand U6353 (N_6353,N_5554,N_5693);
nor U6354 (N_6354,N_5819,N_5583);
nand U6355 (N_6355,N_5552,N_5931);
nor U6356 (N_6356,N_5815,N_5968);
or U6357 (N_6357,N_5868,N_5651);
nand U6358 (N_6358,N_5835,N_5543);
nand U6359 (N_6359,N_5884,N_5910);
or U6360 (N_6360,N_5679,N_5678);
nand U6361 (N_6361,N_5883,N_5770);
nand U6362 (N_6362,N_5661,N_5569);
and U6363 (N_6363,N_5637,N_5842);
xnor U6364 (N_6364,N_5514,N_5832);
and U6365 (N_6365,N_5825,N_5892);
or U6366 (N_6366,N_5808,N_5734);
xor U6367 (N_6367,N_5593,N_5935);
or U6368 (N_6368,N_5936,N_5721);
xor U6369 (N_6369,N_5850,N_5643);
nand U6370 (N_6370,N_5816,N_5966);
and U6371 (N_6371,N_5615,N_5538);
and U6372 (N_6372,N_5978,N_5781);
and U6373 (N_6373,N_5748,N_5787);
or U6374 (N_6374,N_5754,N_5945);
and U6375 (N_6375,N_5732,N_5686);
or U6376 (N_6376,N_5878,N_5556);
or U6377 (N_6377,N_5658,N_5723);
or U6378 (N_6378,N_5738,N_5676);
or U6379 (N_6379,N_5791,N_5547);
and U6380 (N_6380,N_5556,N_5885);
xnor U6381 (N_6381,N_5749,N_5885);
xor U6382 (N_6382,N_5509,N_5649);
nor U6383 (N_6383,N_5996,N_5878);
and U6384 (N_6384,N_5815,N_5961);
nor U6385 (N_6385,N_5959,N_5941);
xor U6386 (N_6386,N_5934,N_5711);
and U6387 (N_6387,N_5897,N_5766);
and U6388 (N_6388,N_5739,N_5717);
and U6389 (N_6389,N_5876,N_5531);
xor U6390 (N_6390,N_5756,N_5868);
nand U6391 (N_6391,N_5654,N_5707);
xor U6392 (N_6392,N_5768,N_5559);
nor U6393 (N_6393,N_5771,N_5547);
nand U6394 (N_6394,N_5706,N_5953);
and U6395 (N_6395,N_5853,N_5637);
and U6396 (N_6396,N_5676,N_5955);
nand U6397 (N_6397,N_5550,N_5850);
or U6398 (N_6398,N_5646,N_5805);
xor U6399 (N_6399,N_5517,N_5986);
and U6400 (N_6400,N_5559,N_5769);
or U6401 (N_6401,N_5915,N_5656);
or U6402 (N_6402,N_5692,N_5528);
nand U6403 (N_6403,N_5708,N_5662);
xor U6404 (N_6404,N_5675,N_5644);
and U6405 (N_6405,N_5839,N_5871);
and U6406 (N_6406,N_5748,N_5602);
nor U6407 (N_6407,N_5741,N_5626);
nand U6408 (N_6408,N_5995,N_5584);
nor U6409 (N_6409,N_5596,N_5809);
or U6410 (N_6410,N_5624,N_5744);
nor U6411 (N_6411,N_5907,N_5729);
and U6412 (N_6412,N_5503,N_5838);
and U6413 (N_6413,N_5872,N_5625);
or U6414 (N_6414,N_5601,N_5615);
or U6415 (N_6415,N_5806,N_5529);
nand U6416 (N_6416,N_5784,N_5880);
or U6417 (N_6417,N_5667,N_5857);
nand U6418 (N_6418,N_5869,N_5752);
xnor U6419 (N_6419,N_5790,N_5556);
xor U6420 (N_6420,N_5808,N_5692);
nor U6421 (N_6421,N_5802,N_5907);
nor U6422 (N_6422,N_5533,N_5945);
or U6423 (N_6423,N_5882,N_5538);
xor U6424 (N_6424,N_5965,N_5833);
nand U6425 (N_6425,N_5615,N_5713);
nand U6426 (N_6426,N_5788,N_5805);
and U6427 (N_6427,N_5615,N_5870);
and U6428 (N_6428,N_5768,N_5840);
or U6429 (N_6429,N_5521,N_5829);
or U6430 (N_6430,N_5671,N_5852);
nand U6431 (N_6431,N_5914,N_5807);
nor U6432 (N_6432,N_5992,N_5552);
nand U6433 (N_6433,N_5891,N_5579);
nor U6434 (N_6434,N_5756,N_5763);
nor U6435 (N_6435,N_5684,N_5747);
nand U6436 (N_6436,N_5715,N_5798);
xor U6437 (N_6437,N_5822,N_5884);
or U6438 (N_6438,N_5602,N_5502);
xor U6439 (N_6439,N_5721,N_5575);
nand U6440 (N_6440,N_5628,N_5990);
or U6441 (N_6441,N_5975,N_5617);
nor U6442 (N_6442,N_5925,N_5865);
and U6443 (N_6443,N_5501,N_5903);
xnor U6444 (N_6444,N_5586,N_5735);
nor U6445 (N_6445,N_5891,N_5978);
nor U6446 (N_6446,N_5671,N_5843);
nor U6447 (N_6447,N_5974,N_5823);
nor U6448 (N_6448,N_5565,N_5810);
xor U6449 (N_6449,N_5832,N_5913);
and U6450 (N_6450,N_5769,N_5617);
and U6451 (N_6451,N_5976,N_5908);
nor U6452 (N_6452,N_5712,N_5904);
xnor U6453 (N_6453,N_5526,N_5684);
nand U6454 (N_6454,N_5561,N_5883);
or U6455 (N_6455,N_5541,N_5857);
and U6456 (N_6456,N_5687,N_5542);
and U6457 (N_6457,N_5768,N_5774);
or U6458 (N_6458,N_5689,N_5785);
or U6459 (N_6459,N_5869,N_5588);
nand U6460 (N_6460,N_5962,N_5542);
nand U6461 (N_6461,N_5863,N_5909);
nand U6462 (N_6462,N_5636,N_5775);
and U6463 (N_6463,N_5835,N_5927);
or U6464 (N_6464,N_5541,N_5775);
nand U6465 (N_6465,N_5795,N_5516);
nor U6466 (N_6466,N_5918,N_5692);
xor U6467 (N_6467,N_5514,N_5671);
and U6468 (N_6468,N_5960,N_5575);
nand U6469 (N_6469,N_5554,N_5500);
xor U6470 (N_6470,N_5945,N_5991);
nand U6471 (N_6471,N_5628,N_5832);
nor U6472 (N_6472,N_5858,N_5787);
xor U6473 (N_6473,N_5681,N_5977);
or U6474 (N_6474,N_5605,N_5823);
and U6475 (N_6475,N_5589,N_5636);
or U6476 (N_6476,N_5558,N_5500);
xor U6477 (N_6477,N_5801,N_5540);
nand U6478 (N_6478,N_5639,N_5767);
and U6479 (N_6479,N_5523,N_5864);
nand U6480 (N_6480,N_5959,N_5831);
xor U6481 (N_6481,N_5899,N_5930);
nor U6482 (N_6482,N_5610,N_5540);
nor U6483 (N_6483,N_5817,N_5861);
and U6484 (N_6484,N_5966,N_5520);
or U6485 (N_6485,N_5502,N_5891);
nor U6486 (N_6486,N_5964,N_5792);
or U6487 (N_6487,N_5728,N_5984);
xor U6488 (N_6488,N_5521,N_5828);
or U6489 (N_6489,N_5946,N_5616);
nor U6490 (N_6490,N_5675,N_5608);
xor U6491 (N_6491,N_5783,N_5775);
nor U6492 (N_6492,N_5675,N_5555);
or U6493 (N_6493,N_5613,N_5803);
or U6494 (N_6494,N_5913,N_5641);
xor U6495 (N_6495,N_5917,N_5709);
nand U6496 (N_6496,N_5936,N_5824);
nand U6497 (N_6497,N_5805,N_5764);
xnor U6498 (N_6498,N_5855,N_5766);
xnor U6499 (N_6499,N_5714,N_5864);
or U6500 (N_6500,N_6162,N_6197);
nor U6501 (N_6501,N_6059,N_6307);
and U6502 (N_6502,N_6318,N_6286);
and U6503 (N_6503,N_6013,N_6329);
nand U6504 (N_6504,N_6422,N_6038);
and U6505 (N_6505,N_6484,N_6259);
nor U6506 (N_6506,N_6423,N_6102);
nor U6507 (N_6507,N_6475,N_6135);
xnor U6508 (N_6508,N_6409,N_6127);
nor U6509 (N_6509,N_6031,N_6463);
or U6510 (N_6510,N_6296,N_6284);
xnor U6511 (N_6511,N_6223,N_6327);
and U6512 (N_6512,N_6216,N_6430);
nor U6513 (N_6513,N_6361,N_6129);
xor U6514 (N_6514,N_6078,N_6432);
or U6515 (N_6515,N_6191,N_6247);
nor U6516 (N_6516,N_6260,N_6351);
nand U6517 (N_6517,N_6410,N_6195);
xnor U6518 (N_6518,N_6248,N_6087);
and U6519 (N_6519,N_6388,N_6072);
nor U6520 (N_6520,N_6320,N_6266);
nor U6521 (N_6521,N_6219,N_6280);
xor U6522 (N_6522,N_6016,N_6198);
and U6523 (N_6523,N_6451,N_6364);
or U6524 (N_6524,N_6261,N_6147);
and U6525 (N_6525,N_6112,N_6084);
xnor U6526 (N_6526,N_6499,N_6406);
nand U6527 (N_6527,N_6371,N_6257);
nor U6528 (N_6528,N_6455,N_6480);
xnor U6529 (N_6529,N_6160,N_6113);
and U6530 (N_6530,N_6048,N_6435);
nor U6531 (N_6531,N_6051,N_6477);
xor U6532 (N_6532,N_6218,N_6085);
nand U6533 (N_6533,N_6495,N_6073);
nor U6534 (N_6534,N_6097,N_6464);
and U6535 (N_6535,N_6452,N_6133);
nand U6536 (N_6536,N_6447,N_6496);
nor U6537 (N_6537,N_6028,N_6044);
and U6538 (N_6538,N_6145,N_6263);
xor U6539 (N_6539,N_6489,N_6148);
nor U6540 (N_6540,N_6377,N_6277);
and U6541 (N_6541,N_6458,N_6478);
xor U6542 (N_6542,N_6319,N_6335);
and U6543 (N_6543,N_6104,N_6490);
and U6544 (N_6544,N_6333,N_6360);
or U6545 (N_6545,N_6159,N_6368);
xnor U6546 (N_6546,N_6056,N_6253);
or U6547 (N_6547,N_6125,N_6256);
xor U6548 (N_6548,N_6356,N_6065);
nand U6549 (N_6549,N_6397,N_6365);
and U6550 (N_6550,N_6267,N_6394);
nand U6551 (N_6551,N_6220,N_6355);
or U6552 (N_6552,N_6354,N_6153);
xor U6553 (N_6553,N_6245,N_6173);
or U6554 (N_6554,N_6214,N_6025);
nand U6555 (N_6555,N_6460,N_6168);
xor U6556 (N_6556,N_6311,N_6299);
xor U6557 (N_6557,N_6081,N_6110);
nand U6558 (N_6558,N_6212,N_6251);
nor U6559 (N_6559,N_6066,N_6120);
nor U6560 (N_6560,N_6021,N_6448);
nor U6561 (N_6561,N_6004,N_6165);
or U6562 (N_6562,N_6033,N_6177);
and U6563 (N_6563,N_6002,N_6313);
or U6564 (N_6564,N_6249,N_6005);
xor U6565 (N_6565,N_6264,N_6389);
nor U6566 (N_6566,N_6121,N_6017);
nand U6567 (N_6567,N_6193,N_6374);
and U6568 (N_6568,N_6180,N_6433);
xor U6569 (N_6569,N_6239,N_6288);
nor U6570 (N_6570,N_6283,N_6396);
nand U6571 (N_6571,N_6080,N_6301);
or U6572 (N_6572,N_6092,N_6428);
nand U6573 (N_6573,N_6407,N_6449);
nor U6574 (N_6574,N_6014,N_6238);
nor U6575 (N_6575,N_6471,N_6134);
or U6576 (N_6576,N_6182,N_6481);
and U6577 (N_6577,N_6415,N_6470);
and U6578 (N_6578,N_6128,N_6010);
or U6579 (N_6579,N_6137,N_6466);
or U6580 (N_6580,N_6187,N_6071);
or U6581 (N_6581,N_6414,N_6184);
nor U6582 (N_6582,N_6403,N_6139);
or U6583 (N_6583,N_6332,N_6457);
nand U6584 (N_6584,N_6109,N_6090);
nor U6585 (N_6585,N_6438,N_6486);
xor U6586 (N_6586,N_6281,N_6348);
nand U6587 (N_6587,N_6459,N_6098);
and U6588 (N_6588,N_6023,N_6209);
nand U6589 (N_6589,N_6210,N_6154);
or U6590 (N_6590,N_6419,N_6379);
or U6591 (N_6591,N_6158,N_6237);
and U6592 (N_6592,N_6330,N_6290);
nor U6593 (N_6593,N_6367,N_6363);
or U6594 (N_6594,N_6445,N_6221);
nand U6595 (N_6595,N_6231,N_6429);
xor U6596 (N_6596,N_6054,N_6254);
nand U6597 (N_6597,N_6342,N_6172);
xnor U6598 (N_6598,N_6352,N_6305);
xnor U6599 (N_6599,N_6234,N_6293);
and U6600 (N_6600,N_6175,N_6310);
or U6601 (N_6601,N_6443,N_6385);
or U6602 (N_6602,N_6456,N_6115);
nor U6603 (N_6603,N_6009,N_6323);
or U6604 (N_6604,N_6094,N_6244);
and U6605 (N_6605,N_6183,N_6316);
and U6606 (N_6606,N_6304,N_6383);
xnor U6607 (N_6607,N_6226,N_6022);
and U6608 (N_6608,N_6019,N_6297);
nor U6609 (N_6609,N_6375,N_6328);
and U6610 (N_6610,N_6292,N_6192);
and U6611 (N_6611,N_6099,N_6105);
or U6612 (N_6612,N_6287,N_6344);
and U6613 (N_6613,N_6298,N_6376);
or U6614 (N_6614,N_6326,N_6049);
or U6615 (N_6615,N_6107,N_6431);
or U6616 (N_6616,N_6207,N_6426);
xor U6617 (N_6617,N_6061,N_6395);
xor U6618 (N_6618,N_6369,N_6140);
or U6619 (N_6619,N_6346,N_6268);
and U6620 (N_6620,N_6041,N_6117);
or U6621 (N_6621,N_6189,N_6294);
or U6622 (N_6622,N_6026,N_6272);
or U6623 (N_6623,N_6164,N_6163);
xor U6624 (N_6624,N_6350,N_6075);
nand U6625 (N_6625,N_6349,N_6390);
xor U6626 (N_6626,N_6181,N_6076);
or U6627 (N_6627,N_6215,N_6067);
nand U6628 (N_6628,N_6161,N_6201);
xor U6629 (N_6629,N_6345,N_6074);
or U6630 (N_6630,N_6408,N_6392);
nand U6631 (N_6631,N_6089,N_6384);
nor U6632 (N_6632,N_6034,N_6483);
xor U6633 (N_6633,N_6402,N_6274);
xnor U6634 (N_6634,N_6252,N_6232);
xnor U6635 (N_6635,N_6086,N_6289);
nor U6636 (N_6636,N_6230,N_6391);
and U6637 (N_6637,N_6169,N_6042);
nor U6638 (N_6638,N_6040,N_6123);
nand U6639 (N_6639,N_6424,N_6303);
or U6640 (N_6640,N_6088,N_6050);
nor U6641 (N_6641,N_6491,N_6425);
nand U6642 (N_6642,N_6058,N_6227);
or U6643 (N_6643,N_6434,N_6273);
nor U6644 (N_6644,N_6100,N_6416);
or U6645 (N_6645,N_6068,N_6082);
and U6646 (N_6646,N_6037,N_6324);
nand U6647 (N_6647,N_6093,N_6242);
nand U6648 (N_6648,N_6453,N_6494);
nand U6649 (N_6649,N_6450,N_6468);
xor U6650 (N_6650,N_6053,N_6208);
xor U6651 (N_6651,N_6150,N_6498);
xnor U6652 (N_6652,N_6308,N_6096);
and U6653 (N_6653,N_6171,N_6046);
and U6654 (N_6654,N_6091,N_6012);
nand U6655 (N_6655,N_6411,N_6029);
nand U6656 (N_6656,N_6217,N_6236);
nand U6657 (N_6657,N_6497,N_6482);
or U6658 (N_6658,N_6176,N_6250);
nor U6659 (N_6659,N_6178,N_6341);
nor U6660 (N_6660,N_6157,N_6462);
or U6661 (N_6661,N_6131,N_6138);
nor U6662 (N_6662,N_6126,N_6243);
nor U6663 (N_6663,N_6132,N_6278);
xor U6664 (N_6664,N_6204,N_6461);
nand U6665 (N_6665,N_6312,N_6473);
nor U6666 (N_6666,N_6108,N_6151);
xnor U6667 (N_6667,N_6295,N_6030);
nor U6668 (N_6668,N_6142,N_6358);
or U6669 (N_6669,N_6321,N_6469);
or U6670 (N_6670,N_6020,N_6202);
or U6671 (N_6671,N_6467,N_6440);
nor U6672 (N_6672,N_6008,N_6106);
nand U6673 (N_6673,N_6413,N_6205);
xor U6674 (N_6674,N_6079,N_6336);
and U6675 (N_6675,N_6225,N_6141);
nor U6676 (N_6676,N_6258,N_6255);
xor U6677 (N_6677,N_6246,N_6186);
and U6678 (N_6678,N_6043,N_6437);
or U6679 (N_6679,N_6386,N_6130);
or U6680 (N_6680,N_6347,N_6339);
or U6681 (N_6681,N_6317,N_6271);
nand U6682 (N_6682,N_6156,N_6062);
nand U6683 (N_6683,N_6229,N_6439);
nand U6684 (N_6684,N_6185,N_6170);
nand U6685 (N_6685,N_6275,N_6338);
xor U6686 (N_6686,N_6291,N_6279);
xnor U6687 (N_6687,N_6362,N_6444);
nor U6688 (N_6688,N_6493,N_6372);
nand U6689 (N_6689,N_6114,N_6136);
xnor U6690 (N_6690,N_6155,N_6331);
nor U6691 (N_6691,N_6003,N_6069);
or U6692 (N_6692,N_6213,N_6045);
xnor U6693 (N_6693,N_6337,N_6276);
or U6694 (N_6694,N_6196,N_6064);
xor U6695 (N_6695,N_6047,N_6378);
nor U6696 (N_6696,N_6488,N_6119);
nand U6697 (N_6697,N_6001,N_6101);
xor U6698 (N_6698,N_6400,N_6306);
and U6699 (N_6699,N_6472,N_6083);
or U6700 (N_6700,N_6179,N_6035);
xnor U6701 (N_6701,N_6190,N_6007);
and U6702 (N_6702,N_6095,N_6366);
nand U6703 (N_6703,N_6373,N_6359);
nor U6704 (N_6704,N_6436,N_6353);
nand U6705 (N_6705,N_6404,N_6036);
or U6706 (N_6706,N_6055,N_6124);
or U6707 (N_6707,N_6152,N_6262);
nand U6708 (N_6708,N_6070,N_6325);
nor U6709 (N_6709,N_6188,N_6027);
and U6710 (N_6710,N_6111,N_6060);
and U6711 (N_6711,N_6006,N_6300);
and U6712 (N_6712,N_6315,N_6492);
nor U6713 (N_6713,N_6167,N_6011);
nand U6714 (N_6714,N_6420,N_6314);
and U6715 (N_6715,N_6199,N_6340);
nand U6716 (N_6716,N_6454,N_6146);
xnor U6717 (N_6717,N_6343,N_6270);
and U6718 (N_6718,N_6144,N_6421);
xnor U6719 (N_6719,N_6398,N_6309);
nor U6720 (N_6720,N_6476,N_6334);
and U6721 (N_6721,N_6322,N_6233);
nand U6722 (N_6722,N_6015,N_6052);
nor U6723 (N_6723,N_6143,N_6166);
nand U6724 (N_6724,N_6285,N_6370);
xor U6725 (N_6725,N_6174,N_6057);
nand U6726 (N_6726,N_6103,N_6487);
nor U6727 (N_6727,N_6401,N_6063);
or U6728 (N_6728,N_6024,N_6442);
nand U6729 (N_6729,N_6077,N_6194);
xnor U6730 (N_6730,N_6265,N_6399);
and U6731 (N_6731,N_6441,N_6418);
or U6732 (N_6732,N_6417,N_6118);
nand U6733 (N_6733,N_6381,N_6479);
or U6734 (N_6734,N_6393,N_6039);
or U6735 (N_6735,N_6122,N_6224);
xnor U6736 (N_6736,N_6412,N_6405);
or U6737 (N_6737,N_6235,N_6228);
nand U6738 (N_6738,N_6387,N_6446);
nor U6739 (N_6739,N_6222,N_6240);
or U6740 (N_6740,N_6382,N_6211);
nor U6741 (N_6741,N_6206,N_6465);
nor U6742 (N_6742,N_6200,N_6427);
xnor U6743 (N_6743,N_6241,N_6380);
nand U6744 (N_6744,N_6203,N_6302);
nand U6745 (N_6745,N_6032,N_6000);
and U6746 (N_6746,N_6018,N_6149);
nand U6747 (N_6747,N_6282,N_6474);
and U6748 (N_6748,N_6485,N_6357);
xnor U6749 (N_6749,N_6269,N_6116);
or U6750 (N_6750,N_6240,N_6143);
xnor U6751 (N_6751,N_6445,N_6222);
and U6752 (N_6752,N_6213,N_6263);
nand U6753 (N_6753,N_6257,N_6201);
and U6754 (N_6754,N_6015,N_6061);
nor U6755 (N_6755,N_6107,N_6082);
and U6756 (N_6756,N_6352,N_6121);
or U6757 (N_6757,N_6437,N_6366);
nor U6758 (N_6758,N_6457,N_6360);
or U6759 (N_6759,N_6227,N_6140);
xor U6760 (N_6760,N_6462,N_6325);
nor U6761 (N_6761,N_6277,N_6147);
nor U6762 (N_6762,N_6451,N_6489);
nor U6763 (N_6763,N_6394,N_6246);
nor U6764 (N_6764,N_6379,N_6438);
and U6765 (N_6765,N_6253,N_6005);
and U6766 (N_6766,N_6284,N_6488);
and U6767 (N_6767,N_6079,N_6234);
xnor U6768 (N_6768,N_6349,N_6469);
and U6769 (N_6769,N_6174,N_6202);
nand U6770 (N_6770,N_6467,N_6269);
xnor U6771 (N_6771,N_6015,N_6225);
xnor U6772 (N_6772,N_6494,N_6254);
nor U6773 (N_6773,N_6149,N_6293);
xnor U6774 (N_6774,N_6418,N_6336);
or U6775 (N_6775,N_6353,N_6134);
or U6776 (N_6776,N_6427,N_6371);
nand U6777 (N_6777,N_6026,N_6054);
nand U6778 (N_6778,N_6128,N_6247);
xnor U6779 (N_6779,N_6433,N_6165);
nand U6780 (N_6780,N_6395,N_6183);
xor U6781 (N_6781,N_6352,N_6048);
or U6782 (N_6782,N_6194,N_6479);
xor U6783 (N_6783,N_6023,N_6219);
nor U6784 (N_6784,N_6321,N_6365);
xnor U6785 (N_6785,N_6181,N_6174);
nor U6786 (N_6786,N_6395,N_6085);
and U6787 (N_6787,N_6049,N_6469);
or U6788 (N_6788,N_6407,N_6363);
xnor U6789 (N_6789,N_6496,N_6499);
nand U6790 (N_6790,N_6284,N_6159);
xnor U6791 (N_6791,N_6097,N_6102);
nand U6792 (N_6792,N_6322,N_6305);
nand U6793 (N_6793,N_6162,N_6013);
xnor U6794 (N_6794,N_6102,N_6261);
nor U6795 (N_6795,N_6179,N_6300);
and U6796 (N_6796,N_6208,N_6249);
xor U6797 (N_6797,N_6058,N_6449);
or U6798 (N_6798,N_6198,N_6136);
nand U6799 (N_6799,N_6482,N_6066);
xnor U6800 (N_6800,N_6111,N_6039);
nand U6801 (N_6801,N_6399,N_6109);
nand U6802 (N_6802,N_6254,N_6296);
xor U6803 (N_6803,N_6332,N_6068);
or U6804 (N_6804,N_6208,N_6343);
and U6805 (N_6805,N_6093,N_6122);
xor U6806 (N_6806,N_6366,N_6039);
nor U6807 (N_6807,N_6429,N_6403);
xor U6808 (N_6808,N_6208,N_6307);
xnor U6809 (N_6809,N_6069,N_6047);
and U6810 (N_6810,N_6489,N_6247);
and U6811 (N_6811,N_6495,N_6431);
and U6812 (N_6812,N_6130,N_6072);
nor U6813 (N_6813,N_6170,N_6246);
nand U6814 (N_6814,N_6326,N_6352);
nor U6815 (N_6815,N_6057,N_6232);
xor U6816 (N_6816,N_6072,N_6440);
nor U6817 (N_6817,N_6432,N_6422);
nand U6818 (N_6818,N_6326,N_6365);
or U6819 (N_6819,N_6344,N_6104);
and U6820 (N_6820,N_6269,N_6424);
and U6821 (N_6821,N_6497,N_6036);
nor U6822 (N_6822,N_6133,N_6305);
and U6823 (N_6823,N_6332,N_6161);
xor U6824 (N_6824,N_6160,N_6141);
nand U6825 (N_6825,N_6450,N_6112);
and U6826 (N_6826,N_6409,N_6362);
and U6827 (N_6827,N_6347,N_6458);
xor U6828 (N_6828,N_6443,N_6431);
nor U6829 (N_6829,N_6069,N_6005);
xnor U6830 (N_6830,N_6302,N_6094);
and U6831 (N_6831,N_6002,N_6060);
nand U6832 (N_6832,N_6117,N_6022);
or U6833 (N_6833,N_6081,N_6079);
nand U6834 (N_6834,N_6262,N_6331);
nand U6835 (N_6835,N_6103,N_6353);
xor U6836 (N_6836,N_6326,N_6363);
or U6837 (N_6837,N_6477,N_6259);
or U6838 (N_6838,N_6333,N_6116);
or U6839 (N_6839,N_6227,N_6319);
xor U6840 (N_6840,N_6194,N_6224);
nand U6841 (N_6841,N_6059,N_6464);
nand U6842 (N_6842,N_6026,N_6310);
nor U6843 (N_6843,N_6275,N_6437);
or U6844 (N_6844,N_6250,N_6321);
and U6845 (N_6845,N_6283,N_6116);
or U6846 (N_6846,N_6110,N_6222);
xnor U6847 (N_6847,N_6182,N_6367);
nor U6848 (N_6848,N_6227,N_6187);
nor U6849 (N_6849,N_6256,N_6249);
or U6850 (N_6850,N_6013,N_6284);
nand U6851 (N_6851,N_6397,N_6439);
xor U6852 (N_6852,N_6476,N_6322);
xnor U6853 (N_6853,N_6143,N_6286);
nand U6854 (N_6854,N_6117,N_6060);
and U6855 (N_6855,N_6244,N_6291);
xor U6856 (N_6856,N_6205,N_6486);
nor U6857 (N_6857,N_6420,N_6140);
xnor U6858 (N_6858,N_6417,N_6239);
nand U6859 (N_6859,N_6476,N_6389);
xnor U6860 (N_6860,N_6425,N_6199);
and U6861 (N_6861,N_6491,N_6304);
and U6862 (N_6862,N_6480,N_6258);
nand U6863 (N_6863,N_6425,N_6414);
xnor U6864 (N_6864,N_6269,N_6230);
nand U6865 (N_6865,N_6105,N_6243);
nor U6866 (N_6866,N_6128,N_6237);
nor U6867 (N_6867,N_6091,N_6309);
xor U6868 (N_6868,N_6049,N_6262);
and U6869 (N_6869,N_6268,N_6470);
and U6870 (N_6870,N_6171,N_6272);
or U6871 (N_6871,N_6137,N_6418);
nand U6872 (N_6872,N_6461,N_6271);
and U6873 (N_6873,N_6260,N_6134);
nand U6874 (N_6874,N_6141,N_6336);
and U6875 (N_6875,N_6238,N_6352);
or U6876 (N_6876,N_6429,N_6337);
or U6877 (N_6877,N_6462,N_6397);
or U6878 (N_6878,N_6186,N_6251);
xor U6879 (N_6879,N_6133,N_6366);
xnor U6880 (N_6880,N_6235,N_6275);
or U6881 (N_6881,N_6116,N_6181);
xnor U6882 (N_6882,N_6052,N_6245);
or U6883 (N_6883,N_6467,N_6404);
and U6884 (N_6884,N_6403,N_6143);
xor U6885 (N_6885,N_6150,N_6374);
nor U6886 (N_6886,N_6291,N_6464);
nand U6887 (N_6887,N_6249,N_6065);
nor U6888 (N_6888,N_6469,N_6409);
nor U6889 (N_6889,N_6278,N_6407);
or U6890 (N_6890,N_6276,N_6434);
nor U6891 (N_6891,N_6329,N_6221);
xnor U6892 (N_6892,N_6227,N_6316);
nor U6893 (N_6893,N_6077,N_6464);
nor U6894 (N_6894,N_6157,N_6080);
xor U6895 (N_6895,N_6206,N_6238);
or U6896 (N_6896,N_6443,N_6445);
nand U6897 (N_6897,N_6290,N_6495);
and U6898 (N_6898,N_6199,N_6253);
or U6899 (N_6899,N_6224,N_6333);
nor U6900 (N_6900,N_6426,N_6398);
or U6901 (N_6901,N_6016,N_6000);
and U6902 (N_6902,N_6227,N_6089);
xor U6903 (N_6903,N_6293,N_6062);
nand U6904 (N_6904,N_6425,N_6299);
and U6905 (N_6905,N_6201,N_6245);
nand U6906 (N_6906,N_6414,N_6409);
nor U6907 (N_6907,N_6411,N_6380);
or U6908 (N_6908,N_6162,N_6318);
nor U6909 (N_6909,N_6386,N_6365);
nor U6910 (N_6910,N_6424,N_6006);
xnor U6911 (N_6911,N_6038,N_6168);
or U6912 (N_6912,N_6406,N_6274);
xnor U6913 (N_6913,N_6001,N_6493);
xnor U6914 (N_6914,N_6238,N_6228);
and U6915 (N_6915,N_6489,N_6238);
or U6916 (N_6916,N_6001,N_6267);
and U6917 (N_6917,N_6061,N_6153);
nand U6918 (N_6918,N_6489,N_6433);
nand U6919 (N_6919,N_6414,N_6058);
and U6920 (N_6920,N_6089,N_6165);
xnor U6921 (N_6921,N_6258,N_6250);
nor U6922 (N_6922,N_6120,N_6455);
nand U6923 (N_6923,N_6027,N_6105);
xnor U6924 (N_6924,N_6297,N_6239);
or U6925 (N_6925,N_6103,N_6026);
nand U6926 (N_6926,N_6220,N_6191);
and U6927 (N_6927,N_6180,N_6382);
nand U6928 (N_6928,N_6287,N_6020);
nor U6929 (N_6929,N_6495,N_6216);
xnor U6930 (N_6930,N_6185,N_6419);
or U6931 (N_6931,N_6120,N_6449);
and U6932 (N_6932,N_6258,N_6360);
xor U6933 (N_6933,N_6035,N_6216);
xnor U6934 (N_6934,N_6105,N_6048);
and U6935 (N_6935,N_6263,N_6216);
or U6936 (N_6936,N_6021,N_6249);
and U6937 (N_6937,N_6179,N_6212);
nand U6938 (N_6938,N_6081,N_6397);
or U6939 (N_6939,N_6279,N_6177);
nand U6940 (N_6940,N_6347,N_6340);
or U6941 (N_6941,N_6288,N_6479);
and U6942 (N_6942,N_6418,N_6167);
xnor U6943 (N_6943,N_6274,N_6142);
or U6944 (N_6944,N_6000,N_6020);
nor U6945 (N_6945,N_6242,N_6226);
nand U6946 (N_6946,N_6214,N_6382);
and U6947 (N_6947,N_6452,N_6063);
nor U6948 (N_6948,N_6340,N_6049);
xnor U6949 (N_6949,N_6003,N_6180);
nand U6950 (N_6950,N_6144,N_6420);
and U6951 (N_6951,N_6368,N_6358);
and U6952 (N_6952,N_6424,N_6387);
and U6953 (N_6953,N_6498,N_6229);
or U6954 (N_6954,N_6188,N_6159);
xnor U6955 (N_6955,N_6286,N_6240);
xor U6956 (N_6956,N_6168,N_6283);
or U6957 (N_6957,N_6128,N_6330);
nand U6958 (N_6958,N_6482,N_6362);
or U6959 (N_6959,N_6096,N_6465);
xor U6960 (N_6960,N_6031,N_6069);
nor U6961 (N_6961,N_6224,N_6485);
nand U6962 (N_6962,N_6492,N_6273);
or U6963 (N_6963,N_6255,N_6108);
and U6964 (N_6964,N_6440,N_6171);
xor U6965 (N_6965,N_6322,N_6392);
nor U6966 (N_6966,N_6258,N_6295);
and U6967 (N_6967,N_6339,N_6244);
and U6968 (N_6968,N_6378,N_6104);
and U6969 (N_6969,N_6355,N_6200);
and U6970 (N_6970,N_6207,N_6054);
nand U6971 (N_6971,N_6036,N_6158);
nand U6972 (N_6972,N_6451,N_6177);
nand U6973 (N_6973,N_6313,N_6076);
nand U6974 (N_6974,N_6454,N_6343);
or U6975 (N_6975,N_6045,N_6393);
xor U6976 (N_6976,N_6072,N_6447);
and U6977 (N_6977,N_6119,N_6311);
xor U6978 (N_6978,N_6012,N_6183);
nand U6979 (N_6979,N_6037,N_6256);
and U6980 (N_6980,N_6084,N_6406);
nor U6981 (N_6981,N_6299,N_6070);
xor U6982 (N_6982,N_6422,N_6464);
nor U6983 (N_6983,N_6030,N_6379);
xnor U6984 (N_6984,N_6310,N_6226);
or U6985 (N_6985,N_6487,N_6148);
nand U6986 (N_6986,N_6241,N_6459);
nor U6987 (N_6987,N_6115,N_6365);
nand U6988 (N_6988,N_6478,N_6077);
nor U6989 (N_6989,N_6282,N_6128);
nor U6990 (N_6990,N_6484,N_6173);
or U6991 (N_6991,N_6002,N_6498);
and U6992 (N_6992,N_6450,N_6251);
nand U6993 (N_6993,N_6079,N_6323);
nand U6994 (N_6994,N_6435,N_6361);
xor U6995 (N_6995,N_6179,N_6233);
or U6996 (N_6996,N_6320,N_6129);
and U6997 (N_6997,N_6460,N_6094);
nand U6998 (N_6998,N_6071,N_6487);
nor U6999 (N_6999,N_6282,N_6396);
or U7000 (N_7000,N_6518,N_6886);
nor U7001 (N_7001,N_6536,N_6627);
and U7002 (N_7002,N_6789,N_6846);
nand U7003 (N_7003,N_6618,N_6844);
xor U7004 (N_7004,N_6630,N_6828);
xnor U7005 (N_7005,N_6504,N_6832);
nand U7006 (N_7006,N_6756,N_6685);
or U7007 (N_7007,N_6523,N_6739);
nand U7008 (N_7008,N_6644,N_6717);
and U7009 (N_7009,N_6767,N_6532);
nand U7010 (N_7010,N_6897,N_6623);
and U7011 (N_7011,N_6976,N_6850);
xnor U7012 (N_7012,N_6662,N_6744);
xor U7013 (N_7013,N_6791,N_6859);
xnor U7014 (N_7014,N_6902,N_6629);
nand U7015 (N_7015,N_6787,N_6928);
or U7016 (N_7016,N_6936,N_6697);
and U7017 (N_7017,N_6683,N_6593);
nor U7018 (N_7018,N_6605,N_6815);
nor U7019 (N_7019,N_6544,N_6993);
or U7020 (N_7020,N_6777,N_6917);
and U7021 (N_7021,N_6770,N_6707);
nand U7022 (N_7022,N_6616,N_6748);
nand U7023 (N_7023,N_6669,N_6804);
nor U7024 (N_7024,N_6933,N_6582);
or U7025 (N_7025,N_6614,N_6915);
or U7026 (N_7026,N_6866,N_6619);
nand U7027 (N_7027,N_6860,N_6842);
nor U7028 (N_7028,N_6913,N_6723);
and U7029 (N_7029,N_6914,N_6573);
xor U7030 (N_7030,N_6758,N_6769);
and U7031 (N_7031,N_6564,N_6575);
xor U7032 (N_7032,N_6525,N_6870);
or U7033 (N_7033,N_6740,N_6505);
nand U7034 (N_7034,N_6706,N_6595);
and U7035 (N_7035,N_6910,N_6974);
or U7036 (N_7036,N_6854,N_6786);
or U7037 (N_7037,N_6882,N_6983);
nor U7038 (N_7038,N_6800,N_6552);
nand U7039 (N_7039,N_6782,N_6898);
and U7040 (N_7040,N_6531,N_6676);
or U7041 (N_7041,N_6780,N_6999);
or U7042 (N_7042,N_6736,N_6773);
xor U7043 (N_7043,N_6576,N_6660);
and U7044 (N_7044,N_6608,N_6817);
nor U7045 (N_7045,N_6514,N_6588);
or U7046 (N_7046,N_6749,N_6925);
nand U7047 (N_7047,N_6597,N_6829);
nand U7048 (N_7048,N_6708,N_6907);
nand U7049 (N_7049,N_6643,N_6524);
nand U7050 (N_7050,N_6964,N_6994);
xnor U7051 (N_7051,N_6764,N_6811);
and U7052 (N_7052,N_6835,N_6931);
xnor U7053 (N_7053,N_6534,N_6672);
nand U7054 (N_7054,N_6788,N_6684);
nor U7055 (N_7055,N_6890,N_6819);
xor U7056 (N_7056,N_6746,N_6851);
or U7057 (N_7057,N_6624,N_6664);
xor U7058 (N_7058,N_6906,N_6986);
xor U7059 (N_7059,N_6973,N_6583);
xnor U7060 (N_7060,N_6603,N_6852);
nor U7061 (N_7061,N_6939,N_6995);
nor U7062 (N_7062,N_6937,N_6803);
xor U7063 (N_7063,N_6935,N_6533);
nand U7064 (N_7064,N_6901,N_6691);
nand U7065 (N_7065,N_6961,N_6923);
nor U7066 (N_7066,N_6857,N_6871);
nor U7067 (N_7067,N_6631,N_6674);
or U7068 (N_7068,N_6659,N_6668);
and U7069 (N_7069,N_6600,N_6895);
and U7070 (N_7070,N_6511,N_6899);
or U7071 (N_7071,N_6700,N_6801);
nor U7072 (N_7072,N_6727,N_6848);
and U7073 (N_7073,N_6927,N_6962);
xor U7074 (N_7074,N_6725,N_6891);
nand U7075 (N_7075,N_6922,N_6806);
or U7076 (N_7076,N_6904,N_6502);
or U7077 (N_7077,N_6594,N_6825);
or U7078 (N_7078,N_6989,N_6509);
nor U7079 (N_7079,N_6953,N_6837);
and U7080 (N_7080,N_6753,N_6952);
or U7081 (N_7081,N_6759,N_6526);
and U7082 (N_7082,N_6881,N_6555);
and U7083 (N_7083,N_6581,N_6887);
xor U7084 (N_7084,N_6985,N_6620);
or U7085 (N_7085,N_6527,N_6947);
nor U7086 (N_7086,N_6641,N_6940);
and U7087 (N_7087,N_6709,N_6823);
xor U7088 (N_7088,N_6734,N_6550);
nor U7089 (N_7089,N_6768,N_6816);
or U7090 (N_7090,N_6716,N_6546);
or U7091 (N_7091,N_6840,N_6506);
and U7092 (N_7092,N_6834,N_6742);
and U7093 (N_7093,N_6889,N_6635);
nor U7094 (N_7094,N_6699,N_6761);
nand U7095 (N_7095,N_6776,N_6554);
nor U7096 (N_7096,N_6984,N_6833);
nand U7097 (N_7097,N_6869,N_6880);
nor U7098 (N_7098,N_6892,N_6675);
and U7099 (N_7099,N_6818,N_6578);
and U7100 (N_7100,N_6515,N_6519);
nand U7101 (N_7101,N_6867,N_6562);
nor U7102 (N_7102,N_6918,N_6778);
nor U7103 (N_7103,N_6948,N_6598);
xnor U7104 (N_7104,N_6980,N_6657);
and U7105 (N_7105,N_6903,N_6843);
and U7106 (N_7106,N_6566,N_6704);
xor U7107 (N_7107,N_6855,N_6858);
nor U7108 (N_7108,N_6567,N_6754);
nor U7109 (N_7109,N_6990,N_6760);
and U7110 (N_7110,N_6971,N_6591);
xnor U7111 (N_7111,N_6522,N_6545);
and U7112 (N_7112,N_6521,N_6720);
and U7113 (N_7113,N_6912,N_6998);
nor U7114 (N_7114,N_6938,N_6563);
nor U7115 (N_7115,N_6571,N_6694);
xor U7116 (N_7116,N_6655,N_6549);
nand U7117 (N_7117,N_6826,N_6879);
xnor U7118 (N_7118,N_6951,N_6649);
nor U7119 (N_7119,N_6693,N_6670);
and U7120 (N_7120,N_6959,N_6680);
xnor U7121 (N_7121,N_6875,N_6654);
nor U7122 (N_7122,N_6622,N_6508);
xnor U7123 (N_7123,N_6596,N_6696);
or U7124 (N_7124,N_6745,N_6666);
or U7125 (N_7125,N_6589,N_6909);
xnor U7126 (N_7126,N_6609,N_6540);
nand U7127 (N_7127,N_6710,N_6743);
and U7128 (N_7128,N_6967,N_6796);
xor U7129 (N_7129,N_6751,N_6868);
nor U7130 (N_7130,N_6920,N_6698);
and U7131 (N_7131,N_6501,N_6516);
nor U7132 (N_7132,N_6645,N_6528);
nor U7133 (N_7133,N_6997,N_6726);
xor U7134 (N_7134,N_6814,N_6812);
and U7135 (N_7135,N_6945,N_6638);
and U7136 (N_7136,N_6601,N_6960);
or U7137 (N_7137,N_6561,N_6689);
nand U7138 (N_7138,N_6982,N_6604);
nor U7139 (N_7139,N_6827,N_6975);
xor U7140 (N_7140,N_6741,N_6580);
and U7141 (N_7141,N_6981,N_6548);
nand U7142 (N_7142,N_6648,N_6547);
or U7143 (N_7143,N_6893,N_6977);
nand U7144 (N_7144,N_6681,N_6957);
xor U7145 (N_7145,N_6729,N_6721);
and U7146 (N_7146,N_6678,N_6690);
nand U7147 (N_7147,N_6763,N_6781);
or U7148 (N_7148,N_6820,N_6877);
and U7149 (N_7149,N_6894,N_6647);
or U7150 (N_7150,N_6577,N_6507);
and U7151 (N_7151,N_6941,N_6530);
nand U7152 (N_7152,N_6830,N_6865);
nor U7153 (N_7153,N_6771,N_6625);
and U7154 (N_7154,N_6752,N_6632);
nand U7155 (N_7155,N_6884,N_6946);
nor U7156 (N_7156,N_6956,N_6838);
nand U7157 (N_7157,N_6772,N_6926);
nor U7158 (N_7158,N_6905,N_6539);
and U7159 (N_7159,N_6799,N_6701);
nand U7160 (N_7160,N_6878,N_6730);
and U7161 (N_7161,N_6841,N_6615);
and U7162 (N_7162,N_6663,N_6757);
or U7163 (N_7163,N_6774,N_6731);
xor U7164 (N_7164,N_6510,N_6541);
xnor U7165 (N_7165,N_6590,N_6612);
or U7166 (N_7166,N_6711,N_6996);
and U7167 (N_7167,N_6813,N_6944);
or U7168 (N_7168,N_6682,N_6610);
xor U7169 (N_7169,N_6568,N_6824);
and U7170 (N_7170,N_6574,N_6686);
or U7171 (N_7171,N_6847,N_6599);
and U7172 (N_7172,N_6738,N_6978);
nor U7173 (N_7173,N_6930,N_6919);
or U7174 (N_7174,N_6908,N_6942);
or U7175 (N_7175,N_6888,N_6652);
or U7176 (N_7176,N_6979,N_6606);
or U7177 (N_7177,N_6535,N_6621);
nand U7178 (N_7178,N_6988,N_6766);
xnor U7179 (N_7179,N_6992,N_6537);
nand U7180 (N_7180,N_6950,N_6633);
and U7181 (N_7181,N_6667,N_6797);
nor U7182 (N_7182,N_6853,N_6737);
nor U7183 (N_7183,N_6517,N_6765);
nand U7184 (N_7184,N_6943,N_6934);
or U7185 (N_7185,N_6790,N_6642);
nand U7186 (N_7186,N_6873,N_6966);
and U7187 (N_7187,N_6714,N_6949);
nor U7188 (N_7188,N_6779,N_6836);
nor U7189 (N_7189,N_6775,N_6512);
nor U7190 (N_7190,N_6969,N_6585);
nand U7191 (N_7191,N_6559,N_6658);
and U7192 (N_7192,N_6570,N_6712);
or U7193 (N_7193,N_6785,N_6965);
nand U7194 (N_7194,N_6713,N_6661);
or U7195 (N_7195,N_6874,N_6687);
nand U7196 (N_7196,N_6883,N_6795);
nand U7197 (N_7197,N_6885,N_6924);
or U7198 (N_7198,N_6958,N_6503);
and U7199 (N_7199,N_6876,N_6560);
nand U7200 (N_7200,N_6861,N_6640);
xnor U7201 (N_7201,N_6972,N_6735);
or U7202 (N_7202,N_6929,N_6695);
and U7203 (N_7203,N_6705,N_6558);
or U7204 (N_7204,N_6702,N_6955);
or U7205 (N_7205,N_6586,N_6565);
or U7206 (N_7206,N_6677,N_6724);
and U7207 (N_7207,N_6513,N_6807);
xnor U7208 (N_7208,N_6794,N_6792);
or U7209 (N_7209,N_6636,N_6613);
nor U7210 (N_7210,N_6520,N_6602);
or U7211 (N_7211,N_6656,N_6968);
nor U7212 (N_7212,N_6932,N_6650);
or U7213 (N_7213,N_6607,N_6728);
xnor U7214 (N_7214,N_6688,N_6849);
xor U7215 (N_7215,N_6862,N_6719);
and U7216 (N_7216,N_6553,N_6572);
nor U7217 (N_7217,N_6808,N_6872);
nor U7218 (N_7218,N_6831,N_6784);
nand U7219 (N_7219,N_6921,N_6911);
nand U7220 (N_7220,N_6856,N_6805);
nor U7221 (N_7221,N_6991,N_6617);
nor U7222 (N_7222,N_6798,N_6543);
nand U7223 (N_7223,N_6755,N_6671);
xor U7224 (N_7224,N_6673,N_6732);
xnor U7225 (N_7225,N_6750,N_6611);
xor U7226 (N_7226,N_6637,N_6802);
or U7227 (N_7227,N_6793,N_6747);
xor U7228 (N_7228,N_6584,N_6557);
or U7229 (N_7229,N_6556,N_6722);
nand U7230 (N_7230,N_6587,N_6500);
nor U7231 (N_7231,N_6703,N_6592);
nand U7232 (N_7232,N_6529,N_6987);
xor U7233 (N_7233,N_6864,N_6718);
nand U7234 (N_7234,N_6651,N_6542);
nand U7235 (N_7235,N_6679,N_6715);
and U7236 (N_7236,N_6845,N_6551);
xnor U7237 (N_7237,N_6954,N_6821);
nand U7238 (N_7238,N_6692,N_6665);
nand U7239 (N_7239,N_6653,N_6809);
nand U7240 (N_7240,N_6783,N_6916);
nor U7241 (N_7241,N_6970,N_6822);
xnor U7242 (N_7242,N_6810,N_6569);
and U7243 (N_7243,N_6896,N_6963);
nor U7244 (N_7244,N_6863,N_6900);
and U7245 (N_7245,N_6579,N_6626);
or U7246 (N_7246,N_6634,N_6628);
nand U7247 (N_7247,N_6733,N_6646);
or U7248 (N_7248,N_6639,N_6839);
and U7249 (N_7249,N_6538,N_6762);
or U7250 (N_7250,N_6591,N_6588);
nor U7251 (N_7251,N_6939,N_6859);
nor U7252 (N_7252,N_6862,N_6626);
xnor U7253 (N_7253,N_6929,N_6934);
nand U7254 (N_7254,N_6586,N_6892);
and U7255 (N_7255,N_6688,N_6927);
nand U7256 (N_7256,N_6766,N_6581);
nor U7257 (N_7257,N_6768,N_6999);
xnor U7258 (N_7258,N_6677,N_6828);
nand U7259 (N_7259,N_6977,N_6962);
or U7260 (N_7260,N_6619,N_6671);
nand U7261 (N_7261,N_6582,N_6788);
and U7262 (N_7262,N_6721,N_6651);
or U7263 (N_7263,N_6575,N_6646);
nor U7264 (N_7264,N_6907,N_6538);
or U7265 (N_7265,N_6638,N_6682);
or U7266 (N_7266,N_6987,N_6623);
or U7267 (N_7267,N_6617,N_6675);
xnor U7268 (N_7268,N_6890,N_6668);
nand U7269 (N_7269,N_6926,N_6800);
and U7270 (N_7270,N_6631,N_6677);
or U7271 (N_7271,N_6824,N_6834);
or U7272 (N_7272,N_6580,N_6925);
and U7273 (N_7273,N_6732,N_6657);
xnor U7274 (N_7274,N_6900,N_6549);
and U7275 (N_7275,N_6511,N_6804);
or U7276 (N_7276,N_6501,N_6574);
or U7277 (N_7277,N_6566,N_6636);
nand U7278 (N_7278,N_6881,N_6776);
and U7279 (N_7279,N_6755,N_6718);
nand U7280 (N_7280,N_6775,N_6811);
nand U7281 (N_7281,N_6513,N_6537);
nand U7282 (N_7282,N_6881,N_6526);
xor U7283 (N_7283,N_6672,N_6952);
nand U7284 (N_7284,N_6592,N_6576);
nand U7285 (N_7285,N_6566,N_6754);
nand U7286 (N_7286,N_6619,N_6768);
nand U7287 (N_7287,N_6965,N_6727);
and U7288 (N_7288,N_6889,N_6690);
or U7289 (N_7289,N_6753,N_6552);
and U7290 (N_7290,N_6646,N_6919);
or U7291 (N_7291,N_6773,N_6666);
nand U7292 (N_7292,N_6933,N_6998);
nor U7293 (N_7293,N_6594,N_6906);
nand U7294 (N_7294,N_6654,N_6896);
and U7295 (N_7295,N_6922,N_6520);
or U7296 (N_7296,N_6533,N_6582);
nand U7297 (N_7297,N_6877,N_6644);
or U7298 (N_7298,N_6708,N_6532);
xnor U7299 (N_7299,N_6715,N_6552);
nor U7300 (N_7300,N_6683,N_6857);
and U7301 (N_7301,N_6625,N_6881);
xnor U7302 (N_7302,N_6674,N_6662);
nor U7303 (N_7303,N_6806,N_6670);
nand U7304 (N_7304,N_6872,N_6680);
nand U7305 (N_7305,N_6761,N_6643);
nor U7306 (N_7306,N_6998,N_6843);
and U7307 (N_7307,N_6830,N_6883);
nand U7308 (N_7308,N_6943,N_6563);
and U7309 (N_7309,N_6786,N_6621);
nor U7310 (N_7310,N_6658,N_6783);
nor U7311 (N_7311,N_6974,N_6836);
and U7312 (N_7312,N_6794,N_6738);
and U7313 (N_7313,N_6592,N_6549);
and U7314 (N_7314,N_6802,N_6601);
nor U7315 (N_7315,N_6882,N_6926);
or U7316 (N_7316,N_6820,N_6894);
or U7317 (N_7317,N_6940,N_6963);
nor U7318 (N_7318,N_6638,N_6718);
nand U7319 (N_7319,N_6828,N_6860);
xor U7320 (N_7320,N_6852,N_6608);
or U7321 (N_7321,N_6565,N_6582);
or U7322 (N_7322,N_6978,N_6526);
or U7323 (N_7323,N_6976,N_6712);
nor U7324 (N_7324,N_6781,N_6787);
nor U7325 (N_7325,N_6944,N_6668);
nand U7326 (N_7326,N_6850,N_6534);
xnor U7327 (N_7327,N_6914,N_6549);
xnor U7328 (N_7328,N_6673,N_6861);
xnor U7329 (N_7329,N_6750,N_6894);
and U7330 (N_7330,N_6804,N_6839);
nor U7331 (N_7331,N_6979,N_6579);
or U7332 (N_7332,N_6697,N_6540);
xor U7333 (N_7333,N_6727,N_6683);
nor U7334 (N_7334,N_6913,N_6672);
nor U7335 (N_7335,N_6557,N_6559);
nand U7336 (N_7336,N_6960,N_6824);
and U7337 (N_7337,N_6811,N_6739);
and U7338 (N_7338,N_6782,N_6561);
nor U7339 (N_7339,N_6934,N_6548);
nor U7340 (N_7340,N_6589,N_6801);
nor U7341 (N_7341,N_6663,N_6584);
xor U7342 (N_7342,N_6628,N_6708);
nor U7343 (N_7343,N_6819,N_6793);
xnor U7344 (N_7344,N_6841,N_6697);
and U7345 (N_7345,N_6923,N_6561);
nor U7346 (N_7346,N_6684,N_6833);
nand U7347 (N_7347,N_6851,N_6908);
xor U7348 (N_7348,N_6636,N_6666);
nor U7349 (N_7349,N_6976,N_6563);
xnor U7350 (N_7350,N_6688,N_6704);
and U7351 (N_7351,N_6802,N_6978);
xnor U7352 (N_7352,N_6788,N_6980);
and U7353 (N_7353,N_6801,N_6547);
xor U7354 (N_7354,N_6626,N_6675);
or U7355 (N_7355,N_6806,N_6803);
xnor U7356 (N_7356,N_6993,N_6798);
nand U7357 (N_7357,N_6544,N_6684);
and U7358 (N_7358,N_6573,N_6960);
xnor U7359 (N_7359,N_6642,N_6860);
and U7360 (N_7360,N_6569,N_6509);
xnor U7361 (N_7361,N_6561,N_6758);
nor U7362 (N_7362,N_6956,N_6863);
xor U7363 (N_7363,N_6997,N_6785);
and U7364 (N_7364,N_6557,N_6833);
and U7365 (N_7365,N_6814,N_6624);
and U7366 (N_7366,N_6858,N_6886);
nand U7367 (N_7367,N_6603,N_6654);
nor U7368 (N_7368,N_6806,N_6832);
or U7369 (N_7369,N_6624,N_6776);
and U7370 (N_7370,N_6733,N_6567);
xnor U7371 (N_7371,N_6996,N_6505);
xor U7372 (N_7372,N_6998,N_6951);
and U7373 (N_7373,N_6535,N_6662);
or U7374 (N_7374,N_6880,N_6530);
and U7375 (N_7375,N_6644,N_6729);
and U7376 (N_7376,N_6562,N_6667);
nand U7377 (N_7377,N_6740,N_6777);
nor U7378 (N_7378,N_6508,N_6631);
nand U7379 (N_7379,N_6923,N_6506);
and U7380 (N_7380,N_6777,N_6951);
xnor U7381 (N_7381,N_6818,N_6598);
nand U7382 (N_7382,N_6827,N_6882);
or U7383 (N_7383,N_6506,N_6798);
xnor U7384 (N_7384,N_6673,N_6543);
nor U7385 (N_7385,N_6701,N_6995);
xor U7386 (N_7386,N_6962,N_6832);
or U7387 (N_7387,N_6702,N_6786);
or U7388 (N_7388,N_6510,N_6913);
nand U7389 (N_7389,N_6925,N_6846);
xnor U7390 (N_7390,N_6570,N_6901);
and U7391 (N_7391,N_6503,N_6640);
and U7392 (N_7392,N_6944,N_6758);
and U7393 (N_7393,N_6540,N_6615);
and U7394 (N_7394,N_6908,N_6880);
nand U7395 (N_7395,N_6861,N_6518);
or U7396 (N_7396,N_6660,N_6609);
nand U7397 (N_7397,N_6858,N_6503);
nor U7398 (N_7398,N_6764,N_6871);
xnor U7399 (N_7399,N_6682,N_6576);
nor U7400 (N_7400,N_6671,N_6950);
nand U7401 (N_7401,N_6649,N_6662);
and U7402 (N_7402,N_6560,N_6533);
xnor U7403 (N_7403,N_6796,N_6573);
and U7404 (N_7404,N_6786,N_6535);
xor U7405 (N_7405,N_6771,N_6557);
or U7406 (N_7406,N_6602,N_6697);
nor U7407 (N_7407,N_6603,N_6516);
and U7408 (N_7408,N_6617,N_6800);
nor U7409 (N_7409,N_6887,N_6826);
nand U7410 (N_7410,N_6985,N_6642);
or U7411 (N_7411,N_6813,N_6895);
or U7412 (N_7412,N_6523,N_6541);
nor U7413 (N_7413,N_6933,N_6517);
nand U7414 (N_7414,N_6726,N_6887);
or U7415 (N_7415,N_6637,N_6750);
nand U7416 (N_7416,N_6546,N_6719);
nor U7417 (N_7417,N_6827,N_6578);
and U7418 (N_7418,N_6805,N_6806);
and U7419 (N_7419,N_6996,N_6649);
and U7420 (N_7420,N_6530,N_6942);
nor U7421 (N_7421,N_6556,N_6708);
nand U7422 (N_7422,N_6821,N_6576);
xnor U7423 (N_7423,N_6631,N_6923);
and U7424 (N_7424,N_6683,N_6591);
nand U7425 (N_7425,N_6954,N_6918);
or U7426 (N_7426,N_6620,N_6635);
and U7427 (N_7427,N_6808,N_6718);
nand U7428 (N_7428,N_6725,N_6512);
xor U7429 (N_7429,N_6683,N_6990);
or U7430 (N_7430,N_6548,N_6980);
nand U7431 (N_7431,N_6847,N_6694);
nor U7432 (N_7432,N_6920,N_6722);
nand U7433 (N_7433,N_6746,N_6848);
nor U7434 (N_7434,N_6523,N_6630);
and U7435 (N_7435,N_6918,N_6519);
nor U7436 (N_7436,N_6902,N_6927);
xnor U7437 (N_7437,N_6701,N_6711);
and U7438 (N_7438,N_6721,N_6831);
xnor U7439 (N_7439,N_6798,N_6672);
nor U7440 (N_7440,N_6941,N_6557);
xnor U7441 (N_7441,N_6549,N_6983);
xor U7442 (N_7442,N_6944,N_6817);
xnor U7443 (N_7443,N_6712,N_6943);
xor U7444 (N_7444,N_6675,N_6659);
nand U7445 (N_7445,N_6699,N_6532);
or U7446 (N_7446,N_6972,N_6653);
xor U7447 (N_7447,N_6509,N_6939);
nor U7448 (N_7448,N_6669,N_6771);
or U7449 (N_7449,N_6981,N_6627);
or U7450 (N_7450,N_6508,N_6833);
and U7451 (N_7451,N_6833,N_6998);
or U7452 (N_7452,N_6549,N_6830);
nor U7453 (N_7453,N_6713,N_6915);
xnor U7454 (N_7454,N_6933,N_6785);
xor U7455 (N_7455,N_6923,N_6781);
nor U7456 (N_7456,N_6880,N_6511);
nor U7457 (N_7457,N_6571,N_6847);
and U7458 (N_7458,N_6727,N_6969);
nand U7459 (N_7459,N_6969,N_6958);
xor U7460 (N_7460,N_6728,N_6651);
nand U7461 (N_7461,N_6653,N_6861);
and U7462 (N_7462,N_6897,N_6884);
xor U7463 (N_7463,N_6542,N_6827);
nand U7464 (N_7464,N_6638,N_6692);
nand U7465 (N_7465,N_6883,N_6731);
nand U7466 (N_7466,N_6717,N_6933);
or U7467 (N_7467,N_6895,N_6659);
and U7468 (N_7468,N_6890,N_6521);
nand U7469 (N_7469,N_6643,N_6886);
or U7470 (N_7470,N_6768,N_6685);
nor U7471 (N_7471,N_6937,N_6840);
or U7472 (N_7472,N_6556,N_6614);
nand U7473 (N_7473,N_6665,N_6929);
nand U7474 (N_7474,N_6876,N_6921);
nor U7475 (N_7475,N_6767,N_6668);
and U7476 (N_7476,N_6622,N_6966);
or U7477 (N_7477,N_6723,N_6934);
nor U7478 (N_7478,N_6560,N_6896);
xnor U7479 (N_7479,N_6707,N_6820);
or U7480 (N_7480,N_6744,N_6582);
nor U7481 (N_7481,N_6565,N_6796);
nor U7482 (N_7482,N_6766,N_6805);
and U7483 (N_7483,N_6808,N_6881);
nor U7484 (N_7484,N_6566,N_6948);
nand U7485 (N_7485,N_6757,N_6533);
nor U7486 (N_7486,N_6906,N_6827);
nand U7487 (N_7487,N_6905,N_6613);
nand U7488 (N_7488,N_6562,N_6502);
and U7489 (N_7489,N_6628,N_6832);
or U7490 (N_7490,N_6968,N_6561);
or U7491 (N_7491,N_6935,N_6516);
nand U7492 (N_7492,N_6544,N_6545);
nor U7493 (N_7493,N_6548,N_6597);
or U7494 (N_7494,N_6748,N_6532);
and U7495 (N_7495,N_6652,N_6620);
nor U7496 (N_7496,N_6809,N_6775);
or U7497 (N_7497,N_6953,N_6684);
nand U7498 (N_7498,N_6752,N_6661);
nor U7499 (N_7499,N_6925,N_6629);
nor U7500 (N_7500,N_7143,N_7036);
nand U7501 (N_7501,N_7354,N_7366);
and U7502 (N_7502,N_7356,N_7003);
xnor U7503 (N_7503,N_7397,N_7473);
or U7504 (N_7504,N_7442,N_7447);
nand U7505 (N_7505,N_7131,N_7172);
nor U7506 (N_7506,N_7492,N_7082);
or U7507 (N_7507,N_7414,N_7048);
and U7508 (N_7508,N_7054,N_7062);
xor U7509 (N_7509,N_7471,N_7495);
xor U7510 (N_7510,N_7437,N_7417);
and U7511 (N_7511,N_7137,N_7141);
or U7512 (N_7512,N_7402,N_7390);
and U7513 (N_7513,N_7215,N_7005);
nor U7514 (N_7514,N_7053,N_7433);
nor U7515 (N_7515,N_7247,N_7256);
nor U7516 (N_7516,N_7330,N_7420);
or U7517 (N_7517,N_7357,N_7446);
or U7518 (N_7518,N_7068,N_7423);
xnor U7519 (N_7519,N_7378,N_7223);
nor U7520 (N_7520,N_7123,N_7008);
xnor U7521 (N_7521,N_7409,N_7004);
nor U7522 (N_7522,N_7193,N_7252);
xor U7523 (N_7523,N_7029,N_7148);
nand U7524 (N_7524,N_7092,N_7147);
nand U7525 (N_7525,N_7311,N_7001);
or U7526 (N_7526,N_7071,N_7466);
nor U7527 (N_7527,N_7216,N_7445);
nor U7528 (N_7528,N_7388,N_7499);
xnor U7529 (N_7529,N_7056,N_7144);
nand U7530 (N_7530,N_7284,N_7482);
nand U7531 (N_7531,N_7343,N_7463);
and U7532 (N_7532,N_7051,N_7305);
xor U7533 (N_7533,N_7323,N_7006);
or U7534 (N_7534,N_7077,N_7010);
and U7535 (N_7535,N_7194,N_7465);
or U7536 (N_7536,N_7220,N_7307);
or U7537 (N_7537,N_7204,N_7134);
xnor U7538 (N_7538,N_7023,N_7325);
nor U7539 (N_7539,N_7327,N_7316);
and U7540 (N_7540,N_7235,N_7116);
or U7541 (N_7541,N_7269,N_7239);
and U7542 (N_7542,N_7274,N_7254);
xnor U7543 (N_7543,N_7488,N_7364);
and U7544 (N_7544,N_7341,N_7047);
xnor U7545 (N_7545,N_7493,N_7360);
nand U7546 (N_7546,N_7335,N_7177);
xor U7547 (N_7547,N_7486,N_7314);
and U7548 (N_7548,N_7014,N_7175);
and U7549 (N_7549,N_7200,N_7210);
and U7550 (N_7550,N_7340,N_7146);
and U7551 (N_7551,N_7227,N_7065);
and U7552 (N_7552,N_7035,N_7407);
or U7553 (N_7553,N_7236,N_7368);
xor U7554 (N_7554,N_7369,N_7348);
xnor U7555 (N_7555,N_7233,N_7179);
nor U7556 (N_7556,N_7483,N_7095);
nand U7557 (N_7557,N_7472,N_7454);
xnor U7558 (N_7558,N_7059,N_7101);
xnor U7559 (N_7559,N_7007,N_7067);
or U7560 (N_7560,N_7430,N_7034);
nor U7561 (N_7561,N_7055,N_7453);
or U7562 (N_7562,N_7221,N_7374);
xor U7563 (N_7563,N_7191,N_7279);
nand U7564 (N_7564,N_7289,N_7481);
nand U7565 (N_7565,N_7324,N_7322);
nand U7566 (N_7566,N_7183,N_7196);
xnor U7567 (N_7567,N_7404,N_7461);
nor U7568 (N_7568,N_7353,N_7302);
xor U7569 (N_7569,N_7057,N_7460);
nor U7570 (N_7570,N_7312,N_7443);
and U7571 (N_7571,N_7208,N_7087);
nand U7572 (N_7572,N_7372,N_7180);
and U7573 (N_7573,N_7344,N_7290);
xor U7574 (N_7574,N_7273,N_7153);
or U7575 (N_7575,N_7242,N_7106);
and U7576 (N_7576,N_7070,N_7283);
nor U7577 (N_7577,N_7432,N_7350);
and U7578 (N_7578,N_7399,N_7099);
nor U7579 (N_7579,N_7020,N_7250);
xor U7580 (N_7580,N_7406,N_7219);
nand U7581 (N_7581,N_7231,N_7209);
xnor U7582 (N_7582,N_7394,N_7145);
and U7583 (N_7583,N_7039,N_7117);
or U7584 (N_7584,N_7464,N_7258);
and U7585 (N_7585,N_7228,N_7450);
or U7586 (N_7586,N_7294,N_7011);
or U7587 (N_7587,N_7142,N_7091);
and U7588 (N_7588,N_7296,N_7139);
nand U7589 (N_7589,N_7136,N_7352);
nor U7590 (N_7590,N_7052,N_7428);
nand U7591 (N_7591,N_7112,N_7469);
xnor U7592 (N_7592,N_7094,N_7458);
and U7593 (N_7593,N_7021,N_7476);
nand U7594 (N_7594,N_7074,N_7484);
or U7595 (N_7595,N_7061,N_7113);
or U7596 (N_7596,N_7028,N_7127);
nand U7597 (N_7597,N_7206,N_7022);
xnor U7598 (N_7598,N_7224,N_7122);
and U7599 (N_7599,N_7395,N_7214);
nor U7600 (N_7600,N_7181,N_7096);
nand U7601 (N_7601,N_7009,N_7104);
nand U7602 (N_7602,N_7226,N_7434);
xor U7603 (N_7603,N_7285,N_7346);
and U7604 (N_7604,N_7411,N_7410);
xor U7605 (N_7605,N_7243,N_7040);
xor U7606 (N_7606,N_7336,N_7467);
xor U7607 (N_7607,N_7081,N_7151);
xnor U7608 (N_7608,N_7287,N_7083);
xor U7609 (N_7609,N_7415,N_7046);
and U7610 (N_7610,N_7462,N_7377);
nand U7611 (N_7611,N_7103,N_7187);
nor U7612 (N_7612,N_7255,N_7363);
nor U7613 (N_7613,N_7381,N_7436);
nand U7614 (N_7614,N_7184,N_7358);
xor U7615 (N_7615,N_7159,N_7063);
xor U7616 (N_7616,N_7424,N_7114);
nor U7617 (N_7617,N_7192,N_7315);
nor U7618 (N_7618,N_7199,N_7490);
nand U7619 (N_7619,N_7129,N_7319);
nor U7620 (N_7620,N_7111,N_7165);
nand U7621 (N_7621,N_7244,N_7419);
and U7622 (N_7622,N_7253,N_7263);
and U7623 (N_7623,N_7173,N_7457);
nand U7624 (N_7624,N_7002,N_7421);
xnor U7625 (N_7625,N_7174,N_7291);
xnor U7626 (N_7626,N_7078,N_7297);
and U7627 (N_7627,N_7408,N_7249);
and U7628 (N_7628,N_7198,N_7286);
nand U7629 (N_7629,N_7386,N_7238);
or U7630 (N_7630,N_7088,N_7361);
nor U7631 (N_7631,N_7079,N_7392);
nand U7632 (N_7632,N_7313,N_7158);
xnor U7633 (N_7633,N_7396,N_7245);
and U7634 (N_7634,N_7119,N_7405);
or U7635 (N_7635,N_7468,N_7485);
and U7636 (N_7636,N_7212,N_7045);
xor U7637 (N_7637,N_7042,N_7265);
nor U7638 (N_7638,N_7037,N_7248);
and U7639 (N_7639,N_7189,N_7050);
and U7640 (N_7640,N_7132,N_7422);
nor U7641 (N_7641,N_7477,N_7060);
nand U7642 (N_7642,N_7229,N_7303);
xor U7643 (N_7643,N_7275,N_7293);
or U7644 (N_7644,N_7202,N_7351);
xor U7645 (N_7645,N_7098,N_7292);
or U7646 (N_7646,N_7225,N_7321);
xor U7647 (N_7647,N_7076,N_7439);
or U7648 (N_7648,N_7403,N_7138);
nor U7649 (N_7649,N_7496,N_7018);
xor U7650 (N_7650,N_7000,N_7261);
or U7651 (N_7651,N_7349,N_7093);
and U7652 (N_7652,N_7170,N_7389);
and U7653 (N_7653,N_7331,N_7387);
xor U7654 (N_7654,N_7272,N_7367);
xor U7655 (N_7655,N_7478,N_7282);
xnor U7656 (N_7656,N_7133,N_7044);
nor U7657 (N_7657,N_7498,N_7125);
or U7658 (N_7658,N_7073,N_7075);
or U7659 (N_7659,N_7120,N_7479);
and U7660 (N_7660,N_7109,N_7418);
nand U7661 (N_7661,N_7298,N_7295);
or U7662 (N_7662,N_7033,N_7385);
and U7663 (N_7663,N_7218,N_7126);
nor U7664 (N_7664,N_7426,N_7066);
nand U7665 (N_7665,N_7130,N_7474);
nor U7666 (N_7666,N_7329,N_7013);
xor U7667 (N_7667,N_7102,N_7080);
nor U7668 (N_7668,N_7201,N_7032);
xnor U7669 (N_7669,N_7085,N_7154);
nor U7670 (N_7670,N_7149,N_7301);
nor U7671 (N_7671,N_7260,N_7449);
and U7672 (N_7672,N_7382,N_7267);
or U7673 (N_7673,N_7240,N_7376);
nor U7674 (N_7674,N_7176,N_7169);
or U7675 (N_7675,N_7299,N_7064);
xnor U7676 (N_7676,N_7487,N_7168);
and U7677 (N_7677,N_7310,N_7379);
xor U7678 (N_7678,N_7456,N_7320);
or U7679 (N_7679,N_7086,N_7049);
xnor U7680 (N_7680,N_7345,N_7280);
nor U7681 (N_7681,N_7425,N_7398);
or U7682 (N_7682,N_7391,N_7203);
and U7683 (N_7683,N_7401,N_7150);
and U7684 (N_7684,N_7207,N_7309);
nand U7685 (N_7685,N_7370,N_7452);
xnor U7686 (N_7686,N_7217,N_7326);
and U7687 (N_7687,N_7304,N_7030);
or U7688 (N_7688,N_7470,N_7015);
or U7689 (N_7689,N_7429,N_7140);
xnor U7690 (N_7690,N_7431,N_7234);
nand U7691 (N_7691,N_7270,N_7246);
xor U7692 (N_7692,N_7166,N_7118);
and U7693 (N_7693,N_7097,N_7268);
and U7694 (N_7694,N_7342,N_7105);
nor U7695 (N_7695,N_7237,N_7412);
or U7696 (N_7696,N_7384,N_7161);
and U7697 (N_7697,N_7160,N_7038);
xnor U7698 (N_7698,N_7383,N_7222);
xnor U7699 (N_7699,N_7251,N_7332);
nand U7700 (N_7700,N_7306,N_7012);
nor U7701 (N_7701,N_7355,N_7089);
and U7702 (N_7702,N_7300,N_7281);
or U7703 (N_7703,N_7259,N_7190);
xor U7704 (N_7704,N_7115,N_7441);
nand U7705 (N_7705,N_7156,N_7277);
xnor U7706 (N_7706,N_7152,N_7416);
xnor U7707 (N_7707,N_7257,N_7164);
nand U7708 (N_7708,N_7359,N_7338);
nor U7709 (N_7709,N_7016,N_7163);
nor U7710 (N_7710,N_7318,N_7027);
and U7711 (N_7711,N_7195,N_7121);
nor U7712 (N_7712,N_7017,N_7438);
and U7713 (N_7713,N_7264,N_7317);
and U7714 (N_7714,N_7019,N_7167);
and U7715 (N_7715,N_7241,N_7440);
xnor U7716 (N_7716,N_7185,N_7084);
and U7717 (N_7717,N_7373,N_7072);
nor U7718 (N_7718,N_7266,N_7024);
nor U7719 (N_7719,N_7171,N_7393);
nor U7720 (N_7720,N_7230,N_7339);
xor U7721 (N_7721,N_7155,N_7491);
nand U7722 (N_7722,N_7026,N_7413);
xnor U7723 (N_7723,N_7178,N_7380);
and U7724 (N_7724,N_7157,N_7110);
nor U7725 (N_7725,N_7435,N_7334);
or U7726 (N_7726,N_7205,N_7276);
nand U7727 (N_7727,N_7232,N_7288);
and U7728 (N_7728,N_7128,N_7375);
and U7729 (N_7729,N_7058,N_7427);
and U7730 (N_7730,N_7480,N_7371);
nor U7731 (N_7731,N_7124,N_7489);
or U7732 (N_7732,N_7262,N_7162);
nor U7733 (N_7733,N_7211,N_7494);
xnor U7734 (N_7734,N_7362,N_7328);
or U7735 (N_7735,N_7337,N_7182);
nor U7736 (N_7736,N_7100,N_7271);
and U7737 (N_7737,N_7459,N_7031);
xor U7738 (N_7738,N_7041,N_7455);
nand U7739 (N_7739,N_7043,N_7451);
xnor U7740 (N_7740,N_7108,N_7278);
or U7741 (N_7741,N_7400,N_7213);
xor U7742 (N_7742,N_7333,N_7107);
nor U7743 (N_7743,N_7186,N_7444);
and U7744 (N_7744,N_7188,N_7197);
xnor U7745 (N_7745,N_7308,N_7497);
nor U7746 (N_7746,N_7347,N_7025);
nor U7747 (N_7747,N_7135,N_7069);
or U7748 (N_7748,N_7365,N_7090);
nand U7749 (N_7749,N_7475,N_7448);
xnor U7750 (N_7750,N_7296,N_7115);
nor U7751 (N_7751,N_7422,N_7361);
nand U7752 (N_7752,N_7108,N_7016);
or U7753 (N_7753,N_7039,N_7171);
nand U7754 (N_7754,N_7195,N_7107);
nand U7755 (N_7755,N_7347,N_7417);
nor U7756 (N_7756,N_7051,N_7375);
or U7757 (N_7757,N_7060,N_7497);
and U7758 (N_7758,N_7124,N_7401);
nor U7759 (N_7759,N_7466,N_7084);
nand U7760 (N_7760,N_7314,N_7302);
xnor U7761 (N_7761,N_7176,N_7186);
nand U7762 (N_7762,N_7189,N_7499);
nor U7763 (N_7763,N_7069,N_7047);
nand U7764 (N_7764,N_7227,N_7075);
nand U7765 (N_7765,N_7222,N_7107);
or U7766 (N_7766,N_7274,N_7339);
xor U7767 (N_7767,N_7321,N_7234);
nand U7768 (N_7768,N_7148,N_7084);
nor U7769 (N_7769,N_7336,N_7021);
nor U7770 (N_7770,N_7210,N_7180);
nand U7771 (N_7771,N_7425,N_7426);
or U7772 (N_7772,N_7316,N_7418);
xor U7773 (N_7773,N_7287,N_7288);
xor U7774 (N_7774,N_7196,N_7455);
and U7775 (N_7775,N_7231,N_7037);
or U7776 (N_7776,N_7364,N_7348);
nand U7777 (N_7777,N_7260,N_7042);
or U7778 (N_7778,N_7103,N_7186);
and U7779 (N_7779,N_7104,N_7225);
xor U7780 (N_7780,N_7282,N_7083);
xnor U7781 (N_7781,N_7025,N_7104);
nor U7782 (N_7782,N_7075,N_7437);
nor U7783 (N_7783,N_7155,N_7097);
or U7784 (N_7784,N_7471,N_7300);
and U7785 (N_7785,N_7101,N_7369);
xnor U7786 (N_7786,N_7130,N_7253);
and U7787 (N_7787,N_7471,N_7474);
and U7788 (N_7788,N_7406,N_7390);
xnor U7789 (N_7789,N_7045,N_7369);
or U7790 (N_7790,N_7442,N_7250);
nor U7791 (N_7791,N_7141,N_7494);
nor U7792 (N_7792,N_7470,N_7482);
and U7793 (N_7793,N_7149,N_7283);
nor U7794 (N_7794,N_7036,N_7249);
and U7795 (N_7795,N_7478,N_7116);
nor U7796 (N_7796,N_7346,N_7484);
or U7797 (N_7797,N_7475,N_7380);
or U7798 (N_7798,N_7206,N_7427);
and U7799 (N_7799,N_7117,N_7205);
nand U7800 (N_7800,N_7089,N_7319);
and U7801 (N_7801,N_7339,N_7163);
or U7802 (N_7802,N_7203,N_7366);
nor U7803 (N_7803,N_7357,N_7265);
xnor U7804 (N_7804,N_7294,N_7062);
xor U7805 (N_7805,N_7345,N_7362);
xnor U7806 (N_7806,N_7266,N_7332);
or U7807 (N_7807,N_7425,N_7310);
nand U7808 (N_7808,N_7393,N_7052);
and U7809 (N_7809,N_7321,N_7343);
nor U7810 (N_7810,N_7454,N_7074);
and U7811 (N_7811,N_7090,N_7017);
nor U7812 (N_7812,N_7418,N_7155);
or U7813 (N_7813,N_7360,N_7296);
nor U7814 (N_7814,N_7210,N_7295);
nor U7815 (N_7815,N_7214,N_7162);
and U7816 (N_7816,N_7184,N_7494);
and U7817 (N_7817,N_7167,N_7264);
or U7818 (N_7818,N_7310,N_7369);
xnor U7819 (N_7819,N_7327,N_7110);
nor U7820 (N_7820,N_7438,N_7190);
xor U7821 (N_7821,N_7401,N_7018);
nor U7822 (N_7822,N_7380,N_7415);
nor U7823 (N_7823,N_7449,N_7372);
xor U7824 (N_7824,N_7002,N_7163);
and U7825 (N_7825,N_7346,N_7417);
nor U7826 (N_7826,N_7159,N_7309);
nand U7827 (N_7827,N_7178,N_7008);
xor U7828 (N_7828,N_7399,N_7432);
nand U7829 (N_7829,N_7303,N_7441);
nand U7830 (N_7830,N_7179,N_7266);
xor U7831 (N_7831,N_7458,N_7452);
nor U7832 (N_7832,N_7113,N_7052);
nand U7833 (N_7833,N_7289,N_7034);
or U7834 (N_7834,N_7050,N_7109);
xnor U7835 (N_7835,N_7222,N_7456);
nand U7836 (N_7836,N_7186,N_7395);
and U7837 (N_7837,N_7352,N_7462);
nand U7838 (N_7838,N_7433,N_7481);
nand U7839 (N_7839,N_7335,N_7197);
nor U7840 (N_7840,N_7116,N_7300);
or U7841 (N_7841,N_7019,N_7171);
and U7842 (N_7842,N_7206,N_7060);
and U7843 (N_7843,N_7266,N_7454);
and U7844 (N_7844,N_7385,N_7471);
and U7845 (N_7845,N_7014,N_7171);
xnor U7846 (N_7846,N_7206,N_7146);
or U7847 (N_7847,N_7385,N_7035);
xnor U7848 (N_7848,N_7122,N_7467);
xnor U7849 (N_7849,N_7213,N_7391);
xnor U7850 (N_7850,N_7492,N_7437);
nor U7851 (N_7851,N_7386,N_7461);
and U7852 (N_7852,N_7044,N_7128);
xnor U7853 (N_7853,N_7055,N_7257);
and U7854 (N_7854,N_7054,N_7097);
nor U7855 (N_7855,N_7368,N_7337);
or U7856 (N_7856,N_7188,N_7410);
or U7857 (N_7857,N_7275,N_7173);
and U7858 (N_7858,N_7016,N_7020);
and U7859 (N_7859,N_7229,N_7306);
xnor U7860 (N_7860,N_7433,N_7440);
xnor U7861 (N_7861,N_7113,N_7264);
or U7862 (N_7862,N_7082,N_7172);
or U7863 (N_7863,N_7431,N_7246);
and U7864 (N_7864,N_7285,N_7128);
nand U7865 (N_7865,N_7109,N_7285);
nor U7866 (N_7866,N_7479,N_7135);
or U7867 (N_7867,N_7024,N_7475);
nor U7868 (N_7868,N_7039,N_7209);
or U7869 (N_7869,N_7428,N_7305);
nor U7870 (N_7870,N_7107,N_7310);
and U7871 (N_7871,N_7068,N_7041);
nand U7872 (N_7872,N_7373,N_7205);
xnor U7873 (N_7873,N_7429,N_7389);
xor U7874 (N_7874,N_7164,N_7237);
and U7875 (N_7875,N_7310,N_7478);
nor U7876 (N_7876,N_7084,N_7261);
nor U7877 (N_7877,N_7098,N_7486);
xnor U7878 (N_7878,N_7422,N_7490);
nor U7879 (N_7879,N_7197,N_7424);
or U7880 (N_7880,N_7102,N_7248);
or U7881 (N_7881,N_7035,N_7033);
nor U7882 (N_7882,N_7111,N_7385);
nor U7883 (N_7883,N_7218,N_7172);
xnor U7884 (N_7884,N_7390,N_7356);
nor U7885 (N_7885,N_7090,N_7101);
xnor U7886 (N_7886,N_7151,N_7264);
nand U7887 (N_7887,N_7293,N_7406);
nand U7888 (N_7888,N_7386,N_7025);
nor U7889 (N_7889,N_7057,N_7378);
or U7890 (N_7890,N_7442,N_7463);
xnor U7891 (N_7891,N_7334,N_7042);
or U7892 (N_7892,N_7399,N_7102);
and U7893 (N_7893,N_7441,N_7200);
and U7894 (N_7894,N_7036,N_7066);
or U7895 (N_7895,N_7413,N_7124);
or U7896 (N_7896,N_7464,N_7271);
nor U7897 (N_7897,N_7099,N_7307);
or U7898 (N_7898,N_7482,N_7229);
and U7899 (N_7899,N_7098,N_7131);
xnor U7900 (N_7900,N_7177,N_7477);
or U7901 (N_7901,N_7340,N_7048);
nand U7902 (N_7902,N_7131,N_7233);
or U7903 (N_7903,N_7161,N_7396);
xor U7904 (N_7904,N_7266,N_7296);
xnor U7905 (N_7905,N_7234,N_7198);
or U7906 (N_7906,N_7333,N_7441);
xor U7907 (N_7907,N_7302,N_7338);
or U7908 (N_7908,N_7366,N_7301);
or U7909 (N_7909,N_7187,N_7299);
or U7910 (N_7910,N_7490,N_7079);
nor U7911 (N_7911,N_7423,N_7027);
nor U7912 (N_7912,N_7000,N_7467);
and U7913 (N_7913,N_7278,N_7181);
or U7914 (N_7914,N_7392,N_7218);
nand U7915 (N_7915,N_7358,N_7393);
and U7916 (N_7916,N_7305,N_7476);
or U7917 (N_7917,N_7466,N_7101);
or U7918 (N_7918,N_7369,N_7393);
and U7919 (N_7919,N_7251,N_7135);
nor U7920 (N_7920,N_7135,N_7165);
nor U7921 (N_7921,N_7086,N_7452);
nor U7922 (N_7922,N_7275,N_7413);
xnor U7923 (N_7923,N_7173,N_7000);
and U7924 (N_7924,N_7350,N_7317);
xor U7925 (N_7925,N_7339,N_7047);
or U7926 (N_7926,N_7039,N_7431);
nor U7927 (N_7927,N_7063,N_7475);
and U7928 (N_7928,N_7070,N_7077);
xnor U7929 (N_7929,N_7168,N_7149);
xnor U7930 (N_7930,N_7021,N_7164);
nor U7931 (N_7931,N_7248,N_7341);
and U7932 (N_7932,N_7487,N_7160);
nor U7933 (N_7933,N_7263,N_7455);
nand U7934 (N_7934,N_7128,N_7325);
or U7935 (N_7935,N_7295,N_7383);
nor U7936 (N_7936,N_7083,N_7034);
nand U7937 (N_7937,N_7099,N_7157);
nand U7938 (N_7938,N_7362,N_7000);
xnor U7939 (N_7939,N_7430,N_7301);
nor U7940 (N_7940,N_7489,N_7184);
nand U7941 (N_7941,N_7208,N_7214);
or U7942 (N_7942,N_7106,N_7263);
xor U7943 (N_7943,N_7194,N_7025);
xor U7944 (N_7944,N_7323,N_7257);
and U7945 (N_7945,N_7146,N_7179);
or U7946 (N_7946,N_7218,N_7202);
nor U7947 (N_7947,N_7350,N_7252);
nand U7948 (N_7948,N_7164,N_7254);
or U7949 (N_7949,N_7185,N_7202);
xor U7950 (N_7950,N_7135,N_7152);
xnor U7951 (N_7951,N_7107,N_7021);
nor U7952 (N_7952,N_7159,N_7270);
or U7953 (N_7953,N_7152,N_7330);
nor U7954 (N_7954,N_7108,N_7072);
nor U7955 (N_7955,N_7429,N_7147);
and U7956 (N_7956,N_7059,N_7247);
xnor U7957 (N_7957,N_7031,N_7359);
nor U7958 (N_7958,N_7127,N_7450);
nand U7959 (N_7959,N_7260,N_7469);
and U7960 (N_7960,N_7052,N_7047);
nor U7961 (N_7961,N_7322,N_7233);
nand U7962 (N_7962,N_7196,N_7388);
nor U7963 (N_7963,N_7225,N_7295);
nor U7964 (N_7964,N_7142,N_7037);
or U7965 (N_7965,N_7054,N_7170);
or U7966 (N_7966,N_7222,N_7282);
nor U7967 (N_7967,N_7044,N_7433);
or U7968 (N_7968,N_7035,N_7146);
and U7969 (N_7969,N_7041,N_7478);
xnor U7970 (N_7970,N_7407,N_7401);
nor U7971 (N_7971,N_7148,N_7277);
nand U7972 (N_7972,N_7396,N_7033);
nand U7973 (N_7973,N_7007,N_7251);
and U7974 (N_7974,N_7492,N_7430);
nand U7975 (N_7975,N_7450,N_7091);
xnor U7976 (N_7976,N_7185,N_7300);
nand U7977 (N_7977,N_7485,N_7354);
nor U7978 (N_7978,N_7035,N_7065);
or U7979 (N_7979,N_7052,N_7356);
or U7980 (N_7980,N_7454,N_7115);
nor U7981 (N_7981,N_7333,N_7494);
and U7982 (N_7982,N_7358,N_7316);
or U7983 (N_7983,N_7334,N_7215);
nor U7984 (N_7984,N_7481,N_7262);
and U7985 (N_7985,N_7315,N_7274);
nor U7986 (N_7986,N_7456,N_7180);
and U7987 (N_7987,N_7236,N_7332);
nor U7988 (N_7988,N_7033,N_7192);
or U7989 (N_7989,N_7128,N_7041);
or U7990 (N_7990,N_7070,N_7367);
or U7991 (N_7991,N_7223,N_7461);
nand U7992 (N_7992,N_7208,N_7105);
and U7993 (N_7993,N_7037,N_7378);
nor U7994 (N_7994,N_7365,N_7173);
xnor U7995 (N_7995,N_7239,N_7106);
or U7996 (N_7996,N_7061,N_7225);
and U7997 (N_7997,N_7193,N_7329);
nor U7998 (N_7998,N_7197,N_7155);
or U7999 (N_7999,N_7160,N_7484);
or U8000 (N_8000,N_7695,N_7864);
nor U8001 (N_8001,N_7880,N_7720);
nand U8002 (N_8002,N_7932,N_7573);
nor U8003 (N_8003,N_7751,N_7830);
nor U8004 (N_8004,N_7536,N_7507);
or U8005 (N_8005,N_7846,N_7651);
xnor U8006 (N_8006,N_7972,N_7577);
or U8007 (N_8007,N_7733,N_7627);
nor U8008 (N_8008,N_7780,N_7735);
and U8009 (N_8009,N_7660,N_7851);
nor U8010 (N_8010,N_7801,N_7689);
and U8011 (N_8011,N_7915,N_7844);
nor U8012 (N_8012,N_7638,N_7973);
or U8013 (N_8013,N_7685,N_7575);
nand U8014 (N_8014,N_7617,N_7517);
or U8015 (N_8015,N_7853,N_7582);
xor U8016 (N_8016,N_7555,N_7825);
and U8017 (N_8017,N_7603,N_7670);
and U8018 (N_8018,N_7522,N_7701);
and U8019 (N_8019,N_7659,N_7841);
and U8020 (N_8020,N_7643,N_7752);
or U8021 (N_8021,N_7871,N_7840);
or U8022 (N_8022,N_7988,N_7703);
nand U8023 (N_8023,N_7585,N_7712);
and U8024 (N_8024,N_7726,N_7762);
nand U8025 (N_8025,N_7583,N_7766);
nand U8026 (N_8026,N_7737,N_7615);
and U8027 (N_8027,N_7919,N_7686);
and U8028 (N_8028,N_7734,N_7745);
and U8029 (N_8029,N_7708,N_7792);
or U8030 (N_8030,N_7635,N_7781);
nand U8031 (N_8031,N_7794,N_7934);
nand U8032 (N_8032,N_7997,N_7796);
or U8033 (N_8033,N_7933,N_7764);
xnor U8034 (N_8034,N_7661,N_7899);
and U8035 (N_8035,N_7967,N_7868);
or U8036 (N_8036,N_7674,N_7984);
xor U8037 (N_8037,N_7918,N_7608);
or U8038 (N_8038,N_7539,N_7977);
nor U8039 (N_8039,N_7858,N_7598);
or U8040 (N_8040,N_7620,N_7525);
and U8041 (N_8041,N_7892,N_7518);
or U8042 (N_8042,N_7818,N_7785);
and U8043 (N_8043,N_7879,N_7609);
nand U8044 (N_8044,N_7537,N_7610);
nor U8045 (N_8045,N_7602,N_7527);
and U8046 (N_8046,N_7787,N_7877);
and U8047 (N_8047,N_7758,N_7628);
nor U8048 (N_8048,N_7748,N_7849);
xnor U8049 (N_8049,N_7778,N_7633);
nor U8050 (N_8050,N_7993,N_7999);
or U8051 (N_8051,N_7510,N_7672);
nand U8052 (N_8052,N_7746,N_7980);
xor U8053 (N_8053,N_7958,N_7731);
or U8054 (N_8054,N_7770,N_7524);
or U8055 (N_8055,N_7508,N_7554);
nor U8056 (N_8056,N_7775,N_7966);
xor U8057 (N_8057,N_7882,N_7538);
xor U8058 (N_8058,N_7957,N_7719);
and U8059 (N_8059,N_7970,N_7631);
nor U8060 (N_8060,N_7543,N_7870);
and U8061 (N_8061,N_7811,N_7978);
xnor U8062 (N_8062,N_7684,N_7898);
nor U8063 (N_8063,N_7855,N_7634);
xnor U8064 (N_8064,N_7904,N_7588);
xor U8065 (N_8065,N_7579,N_7845);
nor U8066 (N_8066,N_7878,N_7905);
or U8067 (N_8067,N_7803,N_7928);
or U8068 (N_8068,N_7856,N_7860);
nand U8069 (N_8069,N_7618,N_7560);
xnor U8070 (N_8070,N_7534,N_7850);
nand U8071 (N_8071,N_7837,N_7549);
nand U8072 (N_8072,N_7697,N_7813);
xor U8073 (N_8073,N_7551,N_7863);
nor U8074 (N_8074,N_7922,N_7971);
nand U8075 (N_8075,N_7506,N_7625);
xor U8076 (N_8076,N_7614,N_7929);
nor U8077 (N_8077,N_7676,N_7753);
nand U8078 (N_8078,N_7663,N_7902);
nand U8079 (N_8079,N_7611,N_7909);
nand U8080 (N_8080,N_7895,N_7657);
nor U8081 (N_8081,N_7713,N_7949);
and U8082 (N_8082,N_7744,N_7831);
xnor U8083 (N_8083,N_7519,N_7976);
nand U8084 (N_8084,N_7710,N_7716);
nor U8085 (N_8085,N_7891,N_7835);
nand U8086 (N_8086,N_7561,N_7662);
xnor U8087 (N_8087,N_7696,N_7694);
nor U8088 (N_8088,N_7606,N_7616);
or U8089 (N_8089,N_7718,N_7702);
nor U8090 (N_8090,N_7668,N_7848);
nor U8091 (N_8091,N_7649,N_7773);
nand U8092 (N_8092,N_7910,N_7869);
nand U8093 (N_8093,N_7693,N_7930);
nor U8094 (N_8094,N_7812,N_7866);
or U8095 (N_8095,N_7884,N_7816);
or U8096 (N_8096,N_7520,N_7673);
or U8097 (N_8097,N_7777,N_7564);
and U8098 (N_8098,N_7962,N_7505);
nor U8099 (N_8099,N_7822,N_7562);
and U8100 (N_8100,N_7671,N_7817);
nor U8101 (N_8101,N_7920,N_7942);
nor U8102 (N_8102,N_7730,N_7998);
nor U8103 (N_8103,N_7772,N_7595);
nand U8104 (N_8104,N_7503,N_7636);
or U8105 (N_8105,N_7945,N_7897);
nand U8106 (N_8106,N_7722,N_7826);
or U8107 (N_8107,N_7600,N_7509);
or U8108 (N_8108,N_7943,N_7688);
nor U8109 (N_8109,N_7883,N_7593);
nand U8110 (N_8110,N_7641,N_7607);
or U8111 (N_8111,N_7950,N_7691);
nand U8112 (N_8112,N_7647,N_7632);
nand U8113 (N_8113,N_7768,N_7911);
or U8114 (N_8114,N_7664,N_7798);
and U8115 (N_8115,N_7836,N_7568);
and U8116 (N_8116,N_7815,N_7605);
or U8117 (N_8117,N_7501,N_7592);
xor U8118 (N_8118,N_7834,N_7747);
nand U8119 (N_8119,N_7574,N_7621);
xnor U8120 (N_8120,N_7665,N_7760);
xnor U8121 (N_8121,N_7797,N_7968);
xor U8122 (N_8122,N_7888,N_7724);
nor U8123 (N_8123,N_7854,N_7556);
xor U8124 (N_8124,N_7799,N_7529);
or U8125 (N_8125,N_7901,N_7623);
nand U8126 (N_8126,N_7547,N_7808);
and U8127 (N_8127,N_7893,N_7533);
or U8128 (N_8128,N_7894,N_7924);
nor U8129 (N_8129,N_7829,N_7738);
or U8130 (N_8130,N_7994,N_7552);
nand U8131 (N_8131,N_7591,N_7907);
and U8132 (N_8132,N_7941,N_7742);
and U8133 (N_8133,N_7776,N_7947);
and U8134 (N_8134,N_7626,N_7927);
nand U8135 (N_8135,N_7754,N_7975);
or U8136 (N_8136,N_7824,N_7546);
xnor U8137 (N_8137,N_7959,N_7956);
nand U8138 (N_8138,N_7655,N_7586);
nand U8139 (N_8139,N_7532,N_7590);
or U8140 (N_8140,N_7881,N_7926);
nand U8141 (N_8141,N_7828,N_7658);
xnor U8142 (N_8142,N_7667,N_7743);
nor U8143 (N_8143,N_7514,N_7596);
nand U8144 (N_8144,N_7523,N_7639);
or U8145 (N_8145,N_7587,N_7875);
nor U8146 (N_8146,N_7951,N_7584);
xnor U8147 (N_8147,N_7791,N_7706);
or U8148 (N_8148,N_7896,N_7675);
and U8149 (N_8149,N_7714,N_7717);
nor U8150 (N_8150,N_7974,N_7707);
or U8151 (N_8151,N_7515,N_7862);
nor U8152 (N_8152,N_7867,N_7982);
xor U8153 (N_8153,N_7653,N_7885);
xor U8154 (N_8154,N_7946,N_7983);
and U8155 (N_8155,N_7755,N_7948);
or U8156 (N_8156,N_7727,N_7557);
xnor U8157 (N_8157,N_7541,N_7839);
and U8158 (N_8158,N_7802,N_7771);
xnor U8159 (N_8159,N_7843,N_7669);
and U8160 (N_8160,N_7680,N_7642);
or U8161 (N_8161,N_7521,N_7783);
or U8162 (N_8162,N_7767,N_7576);
or U8163 (N_8163,N_7936,N_7876);
xor U8164 (N_8164,N_7995,N_7757);
or U8165 (N_8165,N_7728,N_7938);
nand U8166 (N_8166,N_7810,N_7699);
and U8167 (N_8167,N_7961,N_7900);
nand U8168 (N_8168,N_7567,N_7804);
xor U8169 (N_8169,N_7645,N_7559);
xor U8170 (N_8170,N_7566,N_7739);
xor U8171 (N_8171,N_7571,N_7624);
or U8172 (N_8172,N_7935,N_7709);
xor U8173 (N_8173,N_7542,N_7544);
and U8174 (N_8174,N_7916,N_7729);
xor U8175 (N_8175,N_7814,N_7931);
nor U8176 (N_8176,N_7581,N_7923);
xor U8177 (N_8177,N_7989,N_7504);
nand U8178 (N_8178,N_7887,N_7682);
xnor U8179 (N_8179,N_7807,N_7652);
xor U8180 (N_8180,N_7687,N_7819);
nand U8181 (N_8181,N_7741,N_7865);
nor U8182 (N_8182,N_7761,N_7654);
or U8183 (N_8183,N_7612,N_7502);
and U8184 (N_8184,N_7650,N_7784);
xnor U8185 (N_8185,N_7679,N_7805);
xor U8186 (N_8186,N_7553,N_7550);
or U8187 (N_8187,N_7763,N_7530);
or U8188 (N_8188,N_7604,N_7666);
and U8189 (N_8189,N_7512,N_7921);
xnor U8190 (N_8190,N_7789,N_7700);
and U8191 (N_8191,N_7889,N_7913);
nand U8192 (N_8192,N_7622,N_7721);
xor U8193 (N_8193,N_7558,N_7578);
xnor U8194 (N_8194,N_7528,N_7969);
or U8195 (N_8195,N_7692,N_7996);
nor U8196 (N_8196,N_7890,N_7859);
nor U8197 (N_8197,N_7756,N_7725);
or U8198 (N_8198,N_7873,N_7823);
xnor U8199 (N_8199,N_7677,N_7981);
nor U8200 (N_8200,N_7991,N_7992);
nand U8201 (N_8201,N_7809,N_7861);
nor U8202 (N_8202,N_7917,N_7912);
nor U8203 (N_8203,N_7795,N_7872);
xnor U8204 (N_8204,N_7903,N_7779);
nor U8205 (N_8205,N_7800,N_7704);
nand U8206 (N_8206,N_7513,N_7852);
nand U8207 (N_8207,N_7678,N_7630);
and U8208 (N_8208,N_7833,N_7545);
nand U8209 (N_8209,N_7987,N_7986);
nand U8210 (N_8210,N_7925,N_7601);
nor U8211 (N_8211,N_7847,N_7540);
and U8212 (N_8212,N_7765,N_7939);
or U8213 (N_8213,N_7953,N_7820);
nand U8214 (N_8214,N_7711,N_7500);
or U8215 (N_8215,N_7535,N_7736);
or U8216 (N_8216,N_7985,N_7690);
and U8217 (N_8217,N_7786,N_7759);
and U8218 (N_8218,N_7944,N_7965);
xnor U8219 (N_8219,N_7580,N_7740);
nand U8220 (N_8220,N_7511,N_7698);
nand U8221 (N_8221,N_7572,N_7656);
nor U8222 (N_8222,N_7937,N_7749);
nor U8223 (N_8223,N_7648,N_7908);
xor U8224 (N_8224,N_7640,N_7832);
xnor U8225 (N_8225,N_7806,N_7715);
xor U8226 (N_8226,N_7599,N_7613);
or U8227 (N_8227,N_7644,N_7594);
xnor U8228 (N_8228,N_7838,N_7793);
nor U8229 (N_8229,N_7954,N_7723);
nor U8230 (N_8230,N_7548,N_7788);
xor U8231 (N_8231,N_7827,N_7569);
xnor U8232 (N_8232,N_7565,N_7646);
nor U8233 (N_8233,N_7952,N_7821);
xnor U8234 (N_8234,N_7906,N_7842);
xor U8235 (N_8235,N_7769,N_7782);
xnor U8236 (N_8236,N_7629,N_7589);
nor U8237 (N_8237,N_7570,N_7526);
nand U8238 (N_8238,N_7963,N_7790);
and U8239 (N_8239,N_7979,N_7531);
nor U8240 (N_8240,N_7637,N_7597);
xnor U8241 (N_8241,N_7681,N_7940);
nor U8242 (N_8242,N_7990,N_7732);
or U8243 (N_8243,N_7774,N_7964);
and U8244 (N_8244,N_7563,N_7955);
nor U8245 (N_8245,N_7914,N_7705);
nand U8246 (N_8246,N_7516,N_7683);
and U8247 (N_8247,N_7857,N_7960);
nand U8248 (N_8248,N_7874,N_7619);
or U8249 (N_8249,N_7886,N_7750);
and U8250 (N_8250,N_7816,N_7969);
xor U8251 (N_8251,N_7923,N_7502);
and U8252 (N_8252,N_7648,N_7626);
xnor U8253 (N_8253,N_7743,N_7807);
or U8254 (N_8254,N_7799,N_7685);
nor U8255 (N_8255,N_7967,N_7589);
or U8256 (N_8256,N_7614,N_7592);
or U8257 (N_8257,N_7723,N_7851);
nand U8258 (N_8258,N_7765,N_7681);
nor U8259 (N_8259,N_7909,N_7835);
xnor U8260 (N_8260,N_7574,N_7877);
and U8261 (N_8261,N_7827,N_7796);
nor U8262 (N_8262,N_7950,N_7762);
nor U8263 (N_8263,N_7632,N_7878);
nor U8264 (N_8264,N_7939,N_7630);
and U8265 (N_8265,N_7987,N_7820);
and U8266 (N_8266,N_7939,N_7745);
nand U8267 (N_8267,N_7848,N_7946);
or U8268 (N_8268,N_7967,N_7582);
xnor U8269 (N_8269,N_7803,N_7742);
and U8270 (N_8270,N_7979,N_7616);
nor U8271 (N_8271,N_7551,N_7814);
xor U8272 (N_8272,N_7672,N_7919);
and U8273 (N_8273,N_7678,N_7749);
xnor U8274 (N_8274,N_7802,N_7957);
nor U8275 (N_8275,N_7967,N_7973);
and U8276 (N_8276,N_7885,N_7538);
nand U8277 (N_8277,N_7516,N_7636);
xor U8278 (N_8278,N_7637,N_7961);
and U8279 (N_8279,N_7577,N_7982);
xnor U8280 (N_8280,N_7674,N_7739);
or U8281 (N_8281,N_7686,N_7642);
and U8282 (N_8282,N_7641,N_7545);
xnor U8283 (N_8283,N_7619,N_7679);
nor U8284 (N_8284,N_7867,N_7848);
and U8285 (N_8285,N_7514,N_7912);
xnor U8286 (N_8286,N_7798,N_7701);
or U8287 (N_8287,N_7784,N_7737);
nand U8288 (N_8288,N_7961,N_7862);
or U8289 (N_8289,N_7705,N_7986);
and U8290 (N_8290,N_7718,N_7601);
and U8291 (N_8291,N_7804,N_7991);
xnor U8292 (N_8292,N_7808,N_7615);
and U8293 (N_8293,N_7541,N_7673);
nor U8294 (N_8294,N_7914,N_7927);
nor U8295 (N_8295,N_7838,N_7902);
nor U8296 (N_8296,N_7674,N_7573);
or U8297 (N_8297,N_7739,N_7933);
and U8298 (N_8298,N_7651,N_7704);
or U8299 (N_8299,N_7798,N_7960);
and U8300 (N_8300,N_7767,N_7624);
or U8301 (N_8301,N_7745,N_7796);
nor U8302 (N_8302,N_7630,N_7731);
and U8303 (N_8303,N_7765,N_7966);
or U8304 (N_8304,N_7947,N_7561);
and U8305 (N_8305,N_7984,N_7903);
or U8306 (N_8306,N_7803,N_7639);
nand U8307 (N_8307,N_7767,N_7805);
and U8308 (N_8308,N_7892,N_7681);
and U8309 (N_8309,N_7510,N_7663);
nor U8310 (N_8310,N_7814,N_7918);
and U8311 (N_8311,N_7862,N_7576);
and U8312 (N_8312,N_7849,N_7961);
nand U8313 (N_8313,N_7850,N_7678);
nor U8314 (N_8314,N_7908,N_7665);
nor U8315 (N_8315,N_7976,N_7731);
and U8316 (N_8316,N_7804,N_7759);
xnor U8317 (N_8317,N_7880,N_7601);
or U8318 (N_8318,N_7774,N_7568);
or U8319 (N_8319,N_7689,N_7948);
xor U8320 (N_8320,N_7722,N_7589);
and U8321 (N_8321,N_7903,N_7898);
and U8322 (N_8322,N_7867,N_7664);
and U8323 (N_8323,N_7557,N_7859);
nor U8324 (N_8324,N_7750,N_7795);
nor U8325 (N_8325,N_7508,N_7876);
nand U8326 (N_8326,N_7636,N_7979);
xor U8327 (N_8327,N_7824,N_7555);
or U8328 (N_8328,N_7983,N_7780);
or U8329 (N_8329,N_7647,N_7585);
xor U8330 (N_8330,N_7706,N_7570);
nand U8331 (N_8331,N_7819,N_7878);
and U8332 (N_8332,N_7705,N_7569);
nand U8333 (N_8333,N_7547,N_7828);
or U8334 (N_8334,N_7741,N_7889);
xor U8335 (N_8335,N_7753,N_7806);
nand U8336 (N_8336,N_7712,N_7632);
nor U8337 (N_8337,N_7962,N_7742);
and U8338 (N_8338,N_7822,N_7901);
and U8339 (N_8339,N_7849,N_7614);
nand U8340 (N_8340,N_7985,N_7940);
xor U8341 (N_8341,N_7903,N_7881);
nor U8342 (N_8342,N_7982,N_7936);
xor U8343 (N_8343,N_7643,N_7560);
nor U8344 (N_8344,N_7619,N_7576);
and U8345 (N_8345,N_7542,N_7744);
or U8346 (N_8346,N_7755,N_7958);
and U8347 (N_8347,N_7958,N_7639);
nand U8348 (N_8348,N_7537,N_7970);
nand U8349 (N_8349,N_7581,N_7794);
xnor U8350 (N_8350,N_7613,N_7835);
nor U8351 (N_8351,N_7551,N_7892);
xnor U8352 (N_8352,N_7934,N_7938);
nand U8353 (N_8353,N_7986,N_7642);
or U8354 (N_8354,N_7676,N_7921);
nand U8355 (N_8355,N_7751,N_7523);
nor U8356 (N_8356,N_7653,N_7843);
nand U8357 (N_8357,N_7642,N_7631);
nor U8358 (N_8358,N_7928,N_7953);
and U8359 (N_8359,N_7911,N_7965);
nor U8360 (N_8360,N_7951,N_7999);
or U8361 (N_8361,N_7676,N_7733);
xor U8362 (N_8362,N_7672,N_7797);
and U8363 (N_8363,N_7786,N_7616);
xnor U8364 (N_8364,N_7854,N_7511);
nor U8365 (N_8365,N_7818,N_7677);
nor U8366 (N_8366,N_7823,N_7643);
xnor U8367 (N_8367,N_7755,N_7744);
and U8368 (N_8368,N_7600,N_7775);
and U8369 (N_8369,N_7922,N_7665);
or U8370 (N_8370,N_7540,N_7797);
nor U8371 (N_8371,N_7553,N_7629);
or U8372 (N_8372,N_7842,N_7919);
nor U8373 (N_8373,N_7612,N_7856);
or U8374 (N_8374,N_7848,N_7799);
and U8375 (N_8375,N_7602,N_7992);
nor U8376 (N_8376,N_7725,N_7576);
nor U8377 (N_8377,N_7511,N_7764);
nand U8378 (N_8378,N_7933,N_7801);
xnor U8379 (N_8379,N_7822,N_7820);
xor U8380 (N_8380,N_7758,N_7929);
and U8381 (N_8381,N_7685,N_7730);
nor U8382 (N_8382,N_7634,N_7953);
nand U8383 (N_8383,N_7711,N_7576);
and U8384 (N_8384,N_7795,N_7952);
and U8385 (N_8385,N_7783,N_7529);
nand U8386 (N_8386,N_7839,N_7613);
nand U8387 (N_8387,N_7556,N_7593);
and U8388 (N_8388,N_7964,N_7798);
xor U8389 (N_8389,N_7838,N_7798);
and U8390 (N_8390,N_7775,N_7864);
nor U8391 (N_8391,N_7503,N_7559);
and U8392 (N_8392,N_7877,N_7806);
xor U8393 (N_8393,N_7640,N_7991);
xor U8394 (N_8394,N_7708,N_7989);
and U8395 (N_8395,N_7999,N_7578);
xor U8396 (N_8396,N_7647,N_7529);
or U8397 (N_8397,N_7572,N_7667);
nor U8398 (N_8398,N_7907,N_7991);
nand U8399 (N_8399,N_7836,N_7643);
xor U8400 (N_8400,N_7650,N_7513);
nand U8401 (N_8401,N_7650,N_7992);
nor U8402 (N_8402,N_7978,N_7798);
nand U8403 (N_8403,N_7581,N_7786);
xnor U8404 (N_8404,N_7585,N_7759);
and U8405 (N_8405,N_7565,N_7910);
nor U8406 (N_8406,N_7816,N_7794);
or U8407 (N_8407,N_7737,N_7646);
xor U8408 (N_8408,N_7700,N_7648);
or U8409 (N_8409,N_7932,N_7529);
nand U8410 (N_8410,N_7622,N_7695);
nand U8411 (N_8411,N_7928,N_7502);
nor U8412 (N_8412,N_7502,N_7733);
or U8413 (N_8413,N_7693,N_7594);
and U8414 (N_8414,N_7991,N_7936);
nor U8415 (N_8415,N_7622,N_7893);
nand U8416 (N_8416,N_7563,N_7965);
or U8417 (N_8417,N_7884,N_7535);
nand U8418 (N_8418,N_7886,N_7708);
nor U8419 (N_8419,N_7864,N_7856);
nand U8420 (N_8420,N_7647,N_7773);
and U8421 (N_8421,N_7664,N_7693);
xnor U8422 (N_8422,N_7856,N_7507);
nand U8423 (N_8423,N_7918,N_7832);
nor U8424 (N_8424,N_7649,N_7850);
nand U8425 (N_8425,N_7652,N_7971);
nor U8426 (N_8426,N_7636,N_7572);
xnor U8427 (N_8427,N_7925,N_7958);
or U8428 (N_8428,N_7593,N_7522);
nor U8429 (N_8429,N_7687,N_7605);
xor U8430 (N_8430,N_7775,N_7663);
xnor U8431 (N_8431,N_7950,N_7695);
nor U8432 (N_8432,N_7531,N_7870);
xnor U8433 (N_8433,N_7506,N_7662);
or U8434 (N_8434,N_7712,N_7983);
nand U8435 (N_8435,N_7969,N_7959);
xor U8436 (N_8436,N_7715,N_7779);
and U8437 (N_8437,N_7972,N_7562);
and U8438 (N_8438,N_7579,N_7586);
or U8439 (N_8439,N_7571,N_7846);
xnor U8440 (N_8440,N_7941,N_7961);
nor U8441 (N_8441,N_7746,N_7920);
or U8442 (N_8442,N_7622,N_7975);
xnor U8443 (N_8443,N_7652,N_7667);
or U8444 (N_8444,N_7856,N_7976);
nand U8445 (N_8445,N_7614,N_7829);
nand U8446 (N_8446,N_7830,N_7685);
xnor U8447 (N_8447,N_7927,N_7827);
and U8448 (N_8448,N_7916,N_7972);
nor U8449 (N_8449,N_7821,N_7602);
or U8450 (N_8450,N_7769,N_7800);
nor U8451 (N_8451,N_7540,N_7994);
or U8452 (N_8452,N_7718,N_7515);
nand U8453 (N_8453,N_7517,N_7756);
and U8454 (N_8454,N_7947,N_7801);
nand U8455 (N_8455,N_7812,N_7748);
nand U8456 (N_8456,N_7973,N_7632);
or U8457 (N_8457,N_7823,N_7560);
nand U8458 (N_8458,N_7615,N_7606);
xnor U8459 (N_8459,N_7780,N_7688);
nand U8460 (N_8460,N_7530,N_7984);
or U8461 (N_8461,N_7593,N_7844);
nor U8462 (N_8462,N_7897,N_7979);
nor U8463 (N_8463,N_7798,N_7918);
nand U8464 (N_8464,N_7552,N_7755);
and U8465 (N_8465,N_7679,N_7728);
or U8466 (N_8466,N_7677,N_7953);
and U8467 (N_8467,N_7953,N_7881);
or U8468 (N_8468,N_7961,N_7734);
and U8469 (N_8469,N_7934,N_7741);
nand U8470 (N_8470,N_7967,N_7845);
nand U8471 (N_8471,N_7712,N_7874);
xor U8472 (N_8472,N_7724,N_7986);
nand U8473 (N_8473,N_7601,N_7575);
xor U8474 (N_8474,N_7502,N_7852);
nor U8475 (N_8475,N_7671,N_7795);
nor U8476 (N_8476,N_7835,N_7870);
xnor U8477 (N_8477,N_7991,N_7764);
or U8478 (N_8478,N_7824,N_7876);
nand U8479 (N_8479,N_7666,N_7571);
nor U8480 (N_8480,N_7691,N_7772);
xnor U8481 (N_8481,N_7648,N_7632);
and U8482 (N_8482,N_7752,N_7741);
or U8483 (N_8483,N_7575,N_7582);
nor U8484 (N_8484,N_7640,N_7952);
or U8485 (N_8485,N_7604,N_7929);
or U8486 (N_8486,N_7891,N_7857);
nor U8487 (N_8487,N_7865,N_7851);
nand U8488 (N_8488,N_7844,N_7552);
nand U8489 (N_8489,N_7544,N_7989);
or U8490 (N_8490,N_7797,N_7690);
xor U8491 (N_8491,N_7922,N_7605);
xor U8492 (N_8492,N_7909,N_7512);
xor U8493 (N_8493,N_7913,N_7735);
and U8494 (N_8494,N_7580,N_7531);
and U8495 (N_8495,N_7910,N_7930);
or U8496 (N_8496,N_7587,N_7853);
xnor U8497 (N_8497,N_7966,N_7827);
nor U8498 (N_8498,N_7917,N_7835);
and U8499 (N_8499,N_7672,N_7785);
nor U8500 (N_8500,N_8168,N_8086);
and U8501 (N_8501,N_8176,N_8367);
nor U8502 (N_8502,N_8330,N_8184);
or U8503 (N_8503,N_8045,N_8326);
xor U8504 (N_8504,N_8424,N_8122);
nand U8505 (N_8505,N_8169,N_8419);
nand U8506 (N_8506,N_8136,N_8365);
or U8507 (N_8507,N_8213,N_8148);
or U8508 (N_8508,N_8220,N_8327);
nor U8509 (N_8509,N_8091,N_8199);
nand U8510 (N_8510,N_8123,N_8234);
nand U8511 (N_8511,N_8138,N_8301);
and U8512 (N_8512,N_8294,N_8076);
nor U8513 (N_8513,N_8224,N_8054);
xnor U8514 (N_8514,N_8156,N_8111);
nand U8515 (N_8515,N_8238,N_8484);
and U8516 (N_8516,N_8228,N_8012);
xnor U8517 (N_8517,N_8347,N_8428);
or U8518 (N_8518,N_8312,N_8488);
nand U8519 (N_8519,N_8097,N_8172);
and U8520 (N_8520,N_8265,N_8048);
nor U8521 (N_8521,N_8165,N_8426);
and U8522 (N_8522,N_8406,N_8034);
nor U8523 (N_8523,N_8167,N_8134);
or U8524 (N_8524,N_8062,N_8436);
and U8525 (N_8525,N_8246,N_8018);
and U8526 (N_8526,N_8236,N_8103);
or U8527 (N_8527,N_8116,N_8493);
and U8528 (N_8528,N_8047,N_8314);
nor U8529 (N_8529,N_8447,N_8371);
nand U8530 (N_8530,N_8117,N_8458);
xor U8531 (N_8531,N_8140,N_8363);
xor U8532 (N_8532,N_8015,N_8029);
xor U8533 (N_8533,N_8207,N_8074);
xor U8534 (N_8534,N_8453,N_8262);
nand U8535 (N_8535,N_8162,N_8152);
xor U8536 (N_8536,N_8450,N_8397);
and U8537 (N_8537,N_8359,N_8325);
and U8538 (N_8538,N_8470,N_8252);
or U8539 (N_8539,N_8385,N_8042);
nor U8540 (N_8540,N_8124,N_8019);
xnor U8541 (N_8541,N_8126,N_8380);
nor U8542 (N_8542,N_8455,N_8250);
nor U8543 (N_8543,N_8104,N_8376);
and U8544 (N_8544,N_8283,N_8336);
nor U8545 (N_8545,N_8084,N_8320);
xor U8546 (N_8546,N_8316,N_8435);
or U8547 (N_8547,N_8101,N_8090);
or U8548 (N_8548,N_8313,N_8203);
xor U8549 (N_8549,N_8041,N_8171);
and U8550 (N_8550,N_8442,N_8159);
nor U8551 (N_8551,N_8473,N_8415);
or U8552 (N_8552,N_8417,N_8464);
nor U8553 (N_8553,N_8217,N_8348);
xnor U8554 (N_8554,N_8170,N_8269);
and U8555 (N_8555,N_8108,N_8379);
or U8556 (N_8556,N_8078,N_8418);
or U8557 (N_8557,N_8288,N_8248);
and U8558 (N_8558,N_8043,N_8174);
or U8559 (N_8559,N_8334,N_8085);
xor U8560 (N_8560,N_8235,N_8144);
nand U8561 (N_8561,N_8191,N_8155);
nor U8562 (N_8562,N_8185,N_8410);
nand U8563 (N_8563,N_8486,N_8438);
or U8564 (N_8564,N_8149,N_8130);
or U8565 (N_8565,N_8281,N_8016);
nand U8566 (N_8566,N_8182,N_8321);
xnor U8567 (N_8567,N_8193,N_8020);
nor U8568 (N_8568,N_8200,N_8343);
nor U8569 (N_8569,N_8245,N_8386);
and U8570 (N_8570,N_8340,N_8432);
xor U8571 (N_8571,N_8256,N_8364);
xor U8572 (N_8572,N_8231,N_8011);
xor U8573 (N_8573,N_8033,N_8405);
xnor U8574 (N_8574,N_8444,N_8295);
or U8575 (N_8575,N_8333,N_8487);
or U8576 (N_8576,N_8192,N_8287);
xnor U8577 (N_8577,N_8081,N_8163);
or U8578 (N_8578,N_8206,N_8361);
nand U8579 (N_8579,N_8096,N_8142);
nor U8580 (N_8580,N_8490,N_8087);
nand U8581 (N_8581,N_8215,N_8050);
nor U8582 (N_8582,N_8446,N_8300);
or U8583 (N_8583,N_8399,N_8329);
or U8584 (N_8584,N_8483,N_8489);
and U8585 (N_8585,N_8083,N_8175);
or U8586 (N_8586,N_8402,N_8056);
nor U8587 (N_8587,N_8390,N_8431);
nor U8588 (N_8588,N_8279,N_8494);
nand U8589 (N_8589,N_8382,N_8061);
nand U8590 (N_8590,N_8055,N_8059);
and U8591 (N_8591,N_8197,N_8482);
and U8592 (N_8592,N_8388,N_8044);
nand U8593 (N_8593,N_8384,N_8210);
nor U8594 (N_8594,N_8065,N_8244);
and U8595 (N_8595,N_8237,N_8195);
and U8596 (N_8596,N_8060,N_8350);
xnor U8597 (N_8597,N_8378,N_8434);
nand U8598 (N_8598,N_8151,N_8098);
nor U8599 (N_8599,N_8289,N_8064);
nand U8600 (N_8600,N_8357,N_8392);
or U8601 (N_8601,N_8369,N_8120);
nand U8602 (N_8602,N_8221,N_8253);
nor U8603 (N_8603,N_8129,N_8227);
xnor U8604 (N_8604,N_8139,N_8346);
or U8605 (N_8605,N_8258,N_8010);
and U8606 (N_8606,N_8344,N_8499);
or U8607 (N_8607,N_8131,N_8389);
or U8608 (N_8608,N_8299,N_8186);
nor U8609 (N_8609,N_8077,N_8472);
nand U8610 (N_8610,N_8286,N_8107);
and U8611 (N_8611,N_8268,N_8356);
or U8612 (N_8612,N_8179,N_8180);
xor U8613 (N_8613,N_8441,N_8292);
nor U8614 (N_8614,N_8110,N_8260);
and U8615 (N_8615,N_8479,N_8498);
xnor U8616 (N_8616,N_8454,N_8478);
and U8617 (N_8617,N_8310,N_8133);
nor U8618 (N_8618,N_8063,N_8467);
or U8619 (N_8619,N_8323,N_8395);
nor U8620 (N_8620,N_8035,N_8368);
nor U8621 (N_8621,N_8072,N_8353);
or U8622 (N_8622,N_8208,N_8480);
xnor U8623 (N_8623,N_8177,N_8457);
nor U8624 (N_8624,N_8051,N_8004);
nand U8625 (N_8625,N_8427,N_8451);
xnor U8626 (N_8626,N_8093,N_8115);
nor U8627 (N_8627,N_8154,N_8251);
xor U8628 (N_8628,N_8031,N_8423);
nand U8629 (N_8629,N_8311,N_8099);
xnor U8630 (N_8630,N_8461,N_8337);
nor U8631 (N_8631,N_8375,N_8471);
nor U8632 (N_8632,N_8342,N_8293);
and U8633 (N_8633,N_8135,N_8481);
nand U8634 (N_8634,N_8408,N_8317);
xnor U8635 (N_8635,N_8302,N_8223);
nor U8636 (N_8636,N_8025,N_8088);
nand U8637 (N_8637,N_8291,N_8497);
nor U8638 (N_8638,N_8264,N_8421);
xnor U8639 (N_8639,N_8073,N_8194);
nand U8640 (N_8640,N_8053,N_8411);
xor U8641 (N_8641,N_8014,N_8396);
nand U8642 (N_8642,N_8400,N_8021);
or U8643 (N_8643,N_8491,N_8358);
and U8644 (N_8644,N_8324,N_8017);
xnor U8645 (N_8645,N_8121,N_8259);
and U8646 (N_8646,N_8066,N_8146);
or U8647 (N_8647,N_8092,N_8230);
xor U8648 (N_8648,N_8370,N_8173);
nand U8649 (N_8649,N_8404,N_8332);
xnor U8650 (N_8650,N_8331,N_8459);
xnor U8651 (N_8651,N_8443,N_8005);
nor U8652 (N_8652,N_8039,N_8475);
or U8653 (N_8653,N_8437,N_8212);
nor U8654 (N_8654,N_8373,N_8339);
and U8655 (N_8655,N_8449,N_8413);
or U8656 (N_8656,N_8425,N_8150);
xor U8657 (N_8657,N_8477,N_8094);
nand U8658 (N_8658,N_8026,N_8240);
nand U8659 (N_8659,N_8102,N_8469);
nor U8660 (N_8660,N_8335,N_8229);
nand U8661 (N_8661,N_8394,N_8440);
xor U8662 (N_8662,N_8205,N_8328);
and U8663 (N_8663,N_8273,N_8001);
and U8664 (N_8664,N_8307,N_8409);
and U8665 (N_8665,N_8257,N_8222);
nor U8666 (N_8666,N_8218,N_8374);
or U8667 (N_8667,N_8381,N_8495);
or U8668 (N_8668,N_8398,N_8322);
and U8669 (N_8669,N_8351,N_8009);
xor U8670 (N_8670,N_8040,N_8002);
nor U8671 (N_8671,N_8401,N_8249);
and U8672 (N_8672,N_8118,N_8297);
nor U8673 (N_8673,N_8306,N_8341);
nand U8674 (N_8674,N_8100,N_8315);
nor U8675 (N_8675,N_8067,N_8393);
nor U8676 (N_8676,N_8429,N_8080);
nor U8677 (N_8677,N_8158,N_8190);
nand U8678 (N_8678,N_8153,N_8204);
nor U8679 (N_8679,N_8303,N_8391);
nor U8680 (N_8680,N_8119,N_8030);
nand U8681 (N_8681,N_8280,N_8095);
and U8682 (N_8682,N_8105,N_8338);
nand U8683 (N_8683,N_8414,N_8052);
nand U8684 (N_8684,N_8226,N_8112);
or U8685 (N_8685,N_8366,N_8183);
xor U8686 (N_8686,N_8319,N_8233);
xor U8687 (N_8687,N_8492,N_8188);
xor U8688 (N_8688,N_8113,N_8046);
and U8689 (N_8689,N_8032,N_8189);
xor U8690 (N_8690,N_8008,N_8211);
xnor U8691 (N_8691,N_8285,N_8027);
nor U8692 (N_8692,N_8468,N_8164);
and U8693 (N_8693,N_8242,N_8145);
nand U8694 (N_8694,N_8377,N_8079);
nand U8695 (N_8695,N_8352,N_8354);
nand U8696 (N_8696,N_8383,N_8128);
and U8697 (N_8697,N_8345,N_8460);
or U8698 (N_8698,N_8439,N_8267);
and U8699 (N_8699,N_8075,N_8082);
nand U8700 (N_8700,N_8304,N_8462);
nand U8701 (N_8701,N_8201,N_8476);
nor U8702 (N_8702,N_8024,N_8232);
and U8703 (N_8703,N_8003,N_8387);
xnor U8704 (N_8704,N_8127,N_8255);
nor U8705 (N_8705,N_8308,N_8125);
nor U8706 (N_8706,N_8013,N_8407);
xnor U8707 (N_8707,N_8372,N_8070);
or U8708 (N_8708,N_8254,N_8278);
and U8709 (N_8709,N_8272,N_8277);
nor U8710 (N_8710,N_8036,N_8141);
nor U8711 (N_8711,N_8028,N_8412);
nor U8712 (N_8712,N_8037,N_8355);
nand U8713 (N_8713,N_8496,N_8196);
and U8714 (N_8714,N_8187,N_8465);
nor U8715 (N_8715,N_8166,N_8219);
xor U8716 (N_8716,N_8143,N_8261);
or U8717 (N_8717,N_8057,N_8023);
xor U8718 (N_8718,N_8058,N_8474);
xnor U8719 (N_8719,N_8071,N_8147);
nand U8720 (N_8720,N_8270,N_8305);
nor U8721 (N_8721,N_8000,N_8445);
and U8722 (N_8722,N_8038,N_8068);
nand U8723 (N_8723,N_8296,N_8178);
nand U8724 (N_8724,N_8137,N_8318);
nor U8725 (N_8725,N_8225,N_8430);
and U8726 (N_8726,N_8007,N_8241);
xnor U8727 (N_8727,N_8214,N_8161);
and U8728 (N_8728,N_8360,N_8022);
nand U8729 (N_8729,N_8284,N_8157);
xor U8730 (N_8730,N_8239,N_8349);
or U8731 (N_8731,N_8416,N_8448);
nor U8732 (N_8732,N_8181,N_8132);
or U8733 (N_8733,N_8106,N_8463);
or U8734 (N_8734,N_8309,N_8109);
xor U8735 (N_8735,N_8247,N_8271);
xor U8736 (N_8736,N_8216,N_8466);
nor U8737 (N_8737,N_8202,N_8114);
and U8738 (N_8738,N_8276,N_8089);
or U8739 (N_8739,N_8243,N_8362);
nand U8740 (N_8740,N_8160,N_8485);
nand U8741 (N_8741,N_8006,N_8263);
nand U8742 (N_8742,N_8298,N_8282);
xor U8743 (N_8743,N_8452,N_8198);
nor U8744 (N_8744,N_8422,N_8049);
and U8745 (N_8745,N_8069,N_8209);
or U8746 (N_8746,N_8266,N_8456);
or U8747 (N_8747,N_8290,N_8274);
xor U8748 (N_8748,N_8403,N_8275);
or U8749 (N_8749,N_8433,N_8420);
xor U8750 (N_8750,N_8272,N_8336);
or U8751 (N_8751,N_8481,N_8044);
xor U8752 (N_8752,N_8052,N_8239);
or U8753 (N_8753,N_8226,N_8368);
xnor U8754 (N_8754,N_8299,N_8254);
and U8755 (N_8755,N_8233,N_8060);
xor U8756 (N_8756,N_8153,N_8426);
nand U8757 (N_8757,N_8246,N_8374);
nor U8758 (N_8758,N_8271,N_8055);
nor U8759 (N_8759,N_8245,N_8155);
nand U8760 (N_8760,N_8446,N_8402);
nor U8761 (N_8761,N_8153,N_8110);
xnor U8762 (N_8762,N_8307,N_8209);
nand U8763 (N_8763,N_8468,N_8175);
nand U8764 (N_8764,N_8325,N_8285);
xor U8765 (N_8765,N_8344,N_8052);
nand U8766 (N_8766,N_8002,N_8045);
nand U8767 (N_8767,N_8062,N_8066);
nand U8768 (N_8768,N_8314,N_8100);
xor U8769 (N_8769,N_8087,N_8259);
nand U8770 (N_8770,N_8215,N_8391);
xor U8771 (N_8771,N_8019,N_8165);
xor U8772 (N_8772,N_8078,N_8426);
nand U8773 (N_8773,N_8408,N_8319);
and U8774 (N_8774,N_8207,N_8221);
nand U8775 (N_8775,N_8319,N_8086);
xor U8776 (N_8776,N_8358,N_8000);
or U8777 (N_8777,N_8153,N_8259);
nor U8778 (N_8778,N_8056,N_8067);
nor U8779 (N_8779,N_8134,N_8103);
nor U8780 (N_8780,N_8259,N_8240);
and U8781 (N_8781,N_8484,N_8011);
and U8782 (N_8782,N_8248,N_8029);
nand U8783 (N_8783,N_8165,N_8011);
or U8784 (N_8784,N_8310,N_8159);
or U8785 (N_8785,N_8214,N_8131);
or U8786 (N_8786,N_8445,N_8268);
and U8787 (N_8787,N_8256,N_8465);
or U8788 (N_8788,N_8314,N_8470);
and U8789 (N_8789,N_8185,N_8199);
xor U8790 (N_8790,N_8002,N_8095);
nor U8791 (N_8791,N_8203,N_8491);
nor U8792 (N_8792,N_8119,N_8464);
nand U8793 (N_8793,N_8170,N_8305);
xnor U8794 (N_8794,N_8116,N_8216);
or U8795 (N_8795,N_8060,N_8399);
and U8796 (N_8796,N_8114,N_8020);
xnor U8797 (N_8797,N_8036,N_8313);
xor U8798 (N_8798,N_8150,N_8434);
or U8799 (N_8799,N_8097,N_8408);
nand U8800 (N_8800,N_8391,N_8130);
xnor U8801 (N_8801,N_8014,N_8062);
or U8802 (N_8802,N_8378,N_8361);
and U8803 (N_8803,N_8315,N_8445);
nor U8804 (N_8804,N_8460,N_8063);
nor U8805 (N_8805,N_8459,N_8075);
and U8806 (N_8806,N_8316,N_8382);
nor U8807 (N_8807,N_8000,N_8091);
xnor U8808 (N_8808,N_8427,N_8367);
nor U8809 (N_8809,N_8036,N_8072);
and U8810 (N_8810,N_8029,N_8396);
nand U8811 (N_8811,N_8236,N_8183);
nor U8812 (N_8812,N_8174,N_8170);
or U8813 (N_8813,N_8421,N_8338);
nand U8814 (N_8814,N_8401,N_8017);
or U8815 (N_8815,N_8135,N_8225);
xnor U8816 (N_8816,N_8111,N_8144);
nor U8817 (N_8817,N_8035,N_8416);
or U8818 (N_8818,N_8206,N_8264);
and U8819 (N_8819,N_8406,N_8294);
nor U8820 (N_8820,N_8097,N_8084);
and U8821 (N_8821,N_8396,N_8304);
nand U8822 (N_8822,N_8193,N_8474);
nand U8823 (N_8823,N_8036,N_8430);
and U8824 (N_8824,N_8381,N_8372);
xnor U8825 (N_8825,N_8003,N_8025);
or U8826 (N_8826,N_8418,N_8213);
xor U8827 (N_8827,N_8307,N_8318);
xor U8828 (N_8828,N_8279,N_8182);
or U8829 (N_8829,N_8122,N_8419);
xor U8830 (N_8830,N_8299,N_8212);
or U8831 (N_8831,N_8309,N_8363);
or U8832 (N_8832,N_8458,N_8012);
nand U8833 (N_8833,N_8189,N_8277);
and U8834 (N_8834,N_8156,N_8224);
nor U8835 (N_8835,N_8057,N_8148);
nor U8836 (N_8836,N_8416,N_8141);
nor U8837 (N_8837,N_8430,N_8070);
xor U8838 (N_8838,N_8233,N_8016);
and U8839 (N_8839,N_8208,N_8198);
or U8840 (N_8840,N_8458,N_8017);
nand U8841 (N_8841,N_8191,N_8011);
and U8842 (N_8842,N_8024,N_8385);
nand U8843 (N_8843,N_8403,N_8383);
nand U8844 (N_8844,N_8028,N_8279);
nor U8845 (N_8845,N_8038,N_8343);
or U8846 (N_8846,N_8286,N_8132);
xnor U8847 (N_8847,N_8273,N_8375);
or U8848 (N_8848,N_8299,N_8435);
nand U8849 (N_8849,N_8286,N_8290);
and U8850 (N_8850,N_8192,N_8370);
and U8851 (N_8851,N_8371,N_8452);
and U8852 (N_8852,N_8421,N_8076);
and U8853 (N_8853,N_8452,N_8312);
xnor U8854 (N_8854,N_8001,N_8205);
nand U8855 (N_8855,N_8402,N_8078);
and U8856 (N_8856,N_8463,N_8250);
and U8857 (N_8857,N_8034,N_8279);
xor U8858 (N_8858,N_8366,N_8077);
or U8859 (N_8859,N_8209,N_8012);
nand U8860 (N_8860,N_8050,N_8185);
nor U8861 (N_8861,N_8074,N_8020);
nor U8862 (N_8862,N_8134,N_8335);
or U8863 (N_8863,N_8454,N_8402);
and U8864 (N_8864,N_8296,N_8027);
nor U8865 (N_8865,N_8032,N_8358);
xnor U8866 (N_8866,N_8199,N_8418);
xor U8867 (N_8867,N_8297,N_8131);
and U8868 (N_8868,N_8339,N_8459);
and U8869 (N_8869,N_8154,N_8239);
nand U8870 (N_8870,N_8275,N_8268);
and U8871 (N_8871,N_8247,N_8059);
or U8872 (N_8872,N_8105,N_8091);
xnor U8873 (N_8873,N_8228,N_8277);
or U8874 (N_8874,N_8103,N_8449);
xnor U8875 (N_8875,N_8317,N_8223);
nor U8876 (N_8876,N_8281,N_8139);
xnor U8877 (N_8877,N_8219,N_8021);
or U8878 (N_8878,N_8397,N_8312);
and U8879 (N_8879,N_8421,N_8449);
xor U8880 (N_8880,N_8400,N_8177);
nand U8881 (N_8881,N_8184,N_8061);
nand U8882 (N_8882,N_8269,N_8390);
nor U8883 (N_8883,N_8408,N_8370);
nor U8884 (N_8884,N_8180,N_8121);
or U8885 (N_8885,N_8064,N_8097);
or U8886 (N_8886,N_8447,N_8162);
xnor U8887 (N_8887,N_8395,N_8204);
nor U8888 (N_8888,N_8032,N_8062);
or U8889 (N_8889,N_8389,N_8346);
xnor U8890 (N_8890,N_8273,N_8075);
nand U8891 (N_8891,N_8270,N_8350);
or U8892 (N_8892,N_8009,N_8327);
or U8893 (N_8893,N_8413,N_8136);
or U8894 (N_8894,N_8336,N_8087);
and U8895 (N_8895,N_8223,N_8171);
xor U8896 (N_8896,N_8392,N_8130);
or U8897 (N_8897,N_8445,N_8396);
nand U8898 (N_8898,N_8188,N_8467);
nor U8899 (N_8899,N_8276,N_8016);
nor U8900 (N_8900,N_8416,N_8107);
xor U8901 (N_8901,N_8310,N_8135);
nor U8902 (N_8902,N_8476,N_8121);
xnor U8903 (N_8903,N_8050,N_8378);
nand U8904 (N_8904,N_8449,N_8191);
or U8905 (N_8905,N_8079,N_8299);
nand U8906 (N_8906,N_8266,N_8355);
or U8907 (N_8907,N_8318,N_8006);
nor U8908 (N_8908,N_8036,N_8334);
and U8909 (N_8909,N_8079,N_8176);
nor U8910 (N_8910,N_8400,N_8439);
nand U8911 (N_8911,N_8153,N_8285);
xnor U8912 (N_8912,N_8013,N_8369);
xnor U8913 (N_8913,N_8169,N_8143);
nand U8914 (N_8914,N_8052,N_8040);
nor U8915 (N_8915,N_8228,N_8033);
xnor U8916 (N_8916,N_8212,N_8012);
nor U8917 (N_8917,N_8219,N_8287);
nor U8918 (N_8918,N_8386,N_8191);
xnor U8919 (N_8919,N_8364,N_8173);
nor U8920 (N_8920,N_8101,N_8346);
xnor U8921 (N_8921,N_8171,N_8366);
or U8922 (N_8922,N_8243,N_8268);
nand U8923 (N_8923,N_8121,N_8462);
nor U8924 (N_8924,N_8142,N_8109);
nor U8925 (N_8925,N_8044,N_8045);
nand U8926 (N_8926,N_8187,N_8466);
nor U8927 (N_8927,N_8267,N_8344);
nand U8928 (N_8928,N_8230,N_8355);
nor U8929 (N_8929,N_8117,N_8260);
or U8930 (N_8930,N_8385,N_8083);
or U8931 (N_8931,N_8417,N_8421);
or U8932 (N_8932,N_8237,N_8272);
and U8933 (N_8933,N_8393,N_8247);
xor U8934 (N_8934,N_8003,N_8219);
xnor U8935 (N_8935,N_8238,N_8110);
nand U8936 (N_8936,N_8230,N_8239);
and U8937 (N_8937,N_8131,N_8338);
nand U8938 (N_8938,N_8194,N_8074);
xor U8939 (N_8939,N_8217,N_8384);
nor U8940 (N_8940,N_8096,N_8056);
nor U8941 (N_8941,N_8402,N_8109);
and U8942 (N_8942,N_8009,N_8477);
nand U8943 (N_8943,N_8099,N_8428);
nand U8944 (N_8944,N_8251,N_8397);
nor U8945 (N_8945,N_8129,N_8171);
and U8946 (N_8946,N_8037,N_8295);
nor U8947 (N_8947,N_8405,N_8406);
nand U8948 (N_8948,N_8199,N_8443);
and U8949 (N_8949,N_8220,N_8055);
xor U8950 (N_8950,N_8243,N_8165);
nor U8951 (N_8951,N_8472,N_8123);
or U8952 (N_8952,N_8206,N_8239);
nand U8953 (N_8953,N_8258,N_8418);
nand U8954 (N_8954,N_8445,N_8245);
xnor U8955 (N_8955,N_8293,N_8292);
xnor U8956 (N_8956,N_8280,N_8146);
and U8957 (N_8957,N_8113,N_8462);
nor U8958 (N_8958,N_8226,N_8498);
xnor U8959 (N_8959,N_8464,N_8266);
xor U8960 (N_8960,N_8243,N_8416);
or U8961 (N_8961,N_8226,N_8341);
xnor U8962 (N_8962,N_8065,N_8214);
xor U8963 (N_8963,N_8345,N_8397);
and U8964 (N_8964,N_8495,N_8239);
or U8965 (N_8965,N_8250,N_8039);
xor U8966 (N_8966,N_8079,N_8254);
nand U8967 (N_8967,N_8232,N_8068);
nor U8968 (N_8968,N_8112,N_8315);
xor U8969 (N_8969,N_8067,N_8388);
xor U8970 (N_8970,N_8390,N_8194);
xor U8971 (N_8971,N_8044,N_8404);
and U8972 (N_8972,N_8426,N_8092);
nand U8973 (N_8973,N_8270,N_8166);
nor U8974 (N_8974,N_8023,N_8145);
or U8975 (N_8975,N_8118,N_8157);
nor U8976 (N_8976,N_8414,N_8346);
nand U8977 (N_8977,N_8424,N_8025);
nor U8978 (N_8978,N_8403,N_8283);
or U8979 (N_8979,N_8382,N_8131);
or U8980 (N_8980,N_8329,N_8025);
xor U8981 (N_8981,N_8327,N_8092);
or U8982 (N_8982,N_8294,N_8444);
or U8983 (N_8983,N_8262,N_8079);
and U8984 (N_8984,N_8184,N_8177);
nand U8985 (N_8985,N_8109,N_8465);
or U8986 (N_8986,N_8267,N_8443);
nand U8987 (N_8987,N_8210,N_8025);
and U8988 (N_8988,N_8310,N_8262);
nor U8989 (N_8989,N_8251,N_8178);
or U8990 (N_8990,N_8036,N_8241);
xor U8991 (N_8991,N_8207,N_8445);
xor U8992 (N_8992,N_8134,N_8338);
and U8993 (N_8993,N_8227,N_8455);
nand U8994 (N_8994,N_8115,N_8353);
nor U8995 (N_8995,N_8479,N_8281);
nor U8996 (N_8996,N_8036,N_8465);
xnor U8997 (N_8997,N_8220,N_8185);
or U8998 (N_8998,N_8493,N_8165);
nand U8999 (N_8999,N_8432,N_8195);
xnor U9000 (N_9000,N_8919,N_8921);
or U9001 (N_9001,N_8874,N_8848);
or U9002 (N_9002,N_8953,N_8998);
or U9003 (N_9003,N_8963,N_8712);
and U9004 (N_9004,N_8657,N_8689);
nand U9005 (N_9005,N_8508,N_8965);
nor U9006 (N_9006,N_8853,N_8969);
nor U9007 (N_9007,N_8534,N_8753);
xnor U9008 (N_9008,N_8602,N_8554);
and U9009 (N_9009,N_8995,N_8833);
or U9010 (N_9010,N_8793,N_8807);
xor U9011 (N_9011,N_8530,N_8962);
nor U9012 (N_9012,N_8682,N_8935);
and U9013 (N_9013,N_8529,N_8822);
or U9014 (N_9014,N_8887,N_8715);
nand U9015 (N_9015,N_8590,N_8844);
or U9016 (N_9016,N_8842,N_8597);
or U9017 (N_9017,N_8619,N_8889);
or U9018 (N_9018,N_8851,N_8852);
nor U9019 (N_9019,N_8829,N_8687);
and U9020 (N_9020,N_8605,N_8952);
xnor U9021 (N_9021,N_8629,N_8884);
or U9022 (N_9022,N_8573,N_8881);
and U9023 (N_9023,N_8947,N_8517);
and U9024 (N_9024,N_8731,N_8817);
nor U9025 (N_9025,N_8612,N_8911);
nand U9026 (N_9026,N_8631,N_8836);
nand U9027 (N_9027,N_8797,N_8885);
xor U9028 (N_9028,N_8946,N_8796);
nand U9029 (N_9029,N_8511,N_8599);
or U9030 (N_9030,N_8669,N_8788);
or U9031 (N_9031,N_8973,N_8616);
xnor U9032 (N_9032,N_8834,N_8943);
nand U9033 (N_9033,N_8985,N_8835);
and U9034 (N_9034,N_8642,N_8522);
nor U9035 (N_9035,N_8883,N_8580);
nor U9036 (N_9036,N_8592,N_8572);
and U9037 (N_9037,N_8533,N_8798);
or U9038 (N_9038,N_8724,N_8830);
nor U9039 (N_9039,N_8691,N_8979);
or U9040 (N_9040,N_8507,N_8902);
nand U9041 (N_9041,N_8795,N_8639);
xnor U9042 (N_9042,N_8941,N_8688);
nand U9043 (N_9043,N_8920,N_8536);
and U9044 (N_9044,N_8564,N_8557);
xnor U9045 (N_9045,N_8500,N_8974);
nor U9046 (N_9046,N_8879,N_8526);
and U9047 (N_9047,N_8664,N_8790);
nand U9048 (N_9048,N_8825,N_8742);
nand U9049 (N_9049,N_8655,N_8726);
or U9050 (N_9050,N_8800,N_8578);
and U9051 (N_9051,N_8741,N_8686);
nor U9052 (N_9052,N_8558,N_8782);
xor U9053 (N_9053,N_8586,N_8737);
xnor U9054 (N_9054,N_8721,N_8992);
nor U9055 (N_9055,N_8865,N_8934);
nor U9056 (N_9056,N_8542,N_8923);
nand U9057 (N_9057,N_8735,N_8914);
and U9058 (N_9058,N_8990,N_8815);
nand U9059 (N_9059,N_8520,N_8634);
xor U9060 (N_9060,N_8984,N_8703);
and U9061 (N_9061,N_8770,N_8701);
or U9062 (N_9062,N_8824,N_8860);
xnor U9063 (N_9063,N_8804,N_8603);
nor U9064 (N_9064,N_8899,N_8579);
and U9065 (N_9065,N_8736,N_8838);
nand U9066 (N_9066,N_8549,N_8762);
and U9067 (N_9067,N_8751,N_8681);
nand U9068 (N_9068,N_8863,N_8928);
xnor U9069 (N_9069,N_8818,N_8760);
nor U9070 (N_9070,N_8613,N_8819);
or U9071 (N_9071,N_8933,N_8778);
xor U9072 (N_9072,N_8596,N_8978);
and U9073 (N_9073,N_8506,N_8886);
and U9074 (N_9074,N_8684,N_8729);
nand U9075 (N_9075,N_8845,N_8545);
nor U9076 (N_9076,N_8803,N_8570);
xor U9077 (N_9077,N_8810,N_8734);
nor U9078 (N_9078,N_8826,N_8621);
and U9079 (N_9079,N_8768,N_8537);
and U9080 (N_9080,N_8872,N_8502);
nand U9081 (N_9081,N_8954,N_8509);
nand U9082 (N_9082,N_8695,N_8843);
nor U9083 (N_9083,N_8662,N_8764);
and U9084 (N_9084,N_8783,N_8666);
nand U9085 (N_9085,N_8917,N_8660);
nand U9086 (N_9086,N_8707,N_8513);
nand U9087 (N_9087,N_8746,N_8577);
nor U9088 (N_9088,N_8926,N_8606);
nand U9089 (N_9089,N_8988,N_8630);
xnor U9090 (N_9090,N_8591,N_8780);
and U9091 (N_9091,N_8993,N_8991);
and U9092 (N_9092,N_8747,N_8527);
nor U9093 (N_9093,N_8870,N_8980);
and U9094 (N_9094,N_8907,N_8651);
and U9095 (N_9095,N_8582,N_8620);
or U9096 (N_9096,N_8541,N_8938);
nand U9097 (N_9097,N_8722,N_8544);
nand U9098 (N_9098,N_8784,N_8725);
xor U9099 (N_9099,N_8940,N_8752);
xnor U9100 (N_9100,N_8891,N_8813);
nor U9101 (N_9101,N_8565,N_8769);
and U9102 (N_9102,N_8994,N_8659);
nor U9103 (N_9103,N_8799,N_8937);
nor U9104 (N_9104,N_8972,N_8540);
nor U9105 (N_9105,N_8515,N_8647);
nand U9106 (N_9106,N_8588,N_8975);
or U9107 (N_9107,N_8611,N_8525);
nor U9108 (N_9108,N_8854,N_8915);
or U9109 (N_9109,N_8786,N_8608);
nand U9110 (N_9110,N_8906,N_8773);
xor U9111 (N_9111,N_8524,N_8821);
xnor U9112 (N_9112,N_8600,N_8574);
xor U9113 (N_9113,N_8718,N_8971);
or U9114 (N_9114,N_8702,N_8699);
or U9115 (N_9115,N_8837,N_8679);
nor U9116 (N_9116,N_8663,N_8999);
and U9117 (N_9117,N_8705,N_8581);
or U9118 (N_9118,N_8932,N_8716);
nand U9119 (N_9119,N_8623,N_8945);
or U9120 (N_9120,N_8922,N_8615);
xnor U9121 (N_9121,N_8589,N_8868);
nor U9122 (N_9122,N_8996,N_8958);
nand U9123 (N_9123,N_8547,N_8505);
nor U9124 (N_9124,N_8811,N_8567);
nor U9125 (N_9125,N_8950,N_8649);
and U9126 (N_9126,N_8646,N_8949);
or U9127 (N_9127,N_8601,N_8744);
and U9128 (N_9128,N_8670,N_8614);
xor U9129 (N_9129,N_8528,N_8693);
nand U9130 (N_9130,N_8787,N_8882);
nand U9131 (N_9131,N_8568,N_8896);
and U9132 (N_9132,N_8708,N_8624);
or U9133 (N_9133,N_8794,N_8774);
xor U9134 (N_9134,N_8698,N_8931);
nand U9135 (N_9135,N_8755,N_8968);
or U9136 (N_9136,N_8959,N_8839);
or U9137 (N_9137,N_8673,N_8903);
xor U9138 (N_9138,N_8862,N_8641);
or U9139 (N_9139,N_8514,N_8503);
or U9140 (N_9140,N_8849,N_8640);
xor U9141 (N_9141,N_8504,N_8587);
and U9142 (N_9142,N_8987,N_8633);
xor U9143 (N_9143,N_8925,N_8743);
and U9144 (N_9144,N_8680,N_8981);
and U9145 (N_9145,N_8677,N_8964);
nor U9146 (N_9146,N_8519,N_8924);
nor U9147 (N_9147,N_8694,N_8977);
nand U9148 (N_9148,N_8713,N_8888);
xor U9149 (N_9149,N_8719,N_8535);
xor U9150 (N_9150,N_8665,N_8692);
xnor U9151 (N_9151,N_8538,N_8957);
nor U9152 (N_9152,N_8775,N_8880);
or U9153 (N_9153,N_8892,N_8635);
nor U9154 (N_9154,N_8717,N_8856);
nor U9155 (N_9155,N_8823,N_8518);
nand U9156 (N_9156,N_8900,N_8555);
or U9157 (N_9157,N_8767,N_8727);
nand U9158 (N_9158,N_8850,N_8548);
or U9159 (N_9159,N_8711,N_8696);
or U9160 (N_9160,N_8864,N_8930);
nand U9161 (N_9161,N_8918,N_8714);
or U9162 (N_9162,N_8948,N_8622);
nand U9163 (N_9163,N_8913,N_8551);
or U9164 (N_9164,N_8857,N_8643);
and U9165 (N_9165,N_8970,N_8671);
nand U9166 (N_9166,N_8560,N_8967);
and U9167 (N_9167,N_8531,N_8654);
and U9168 (N_9168,N_8831,N_8674);
and U9169 (N_9169,N_8912,N_8576);
and U9170 (N_9170,N_8706,N_8709);
and U9171 (N_9171,N_8607,N_8512);
or U9172 (N_9172,N_8598,N_8986);
and U9173 (N_9173,N_8861,N_8828);
nor U9174 (N_9174,N_8909,N_8672);
nand U9175 (N_9175,N_8552,N_8792);
xnor U9176 (N_9176,N_8583,N_8869);
or U9177 (N_9177,N_8789,N_8748);
nor U9178 (N_9178,N_8894,N_8756);
nor U9179 (N_9179,N_8876,N_8816);
nor U9180 (N_9180,N_8739,N_8728);
xor U9181 (N_9181,N_8546,N_8791);
nor U9182 (N_9182,N_8650,N_8771);
nor U9183 (N_9183,N_8627,N_8750);
xor U9184 (N_9184,N_8895,N_8827);
nand U9185 (N_9185,N_8539,N_8961);
xnor U9186 (N_9186,N_8936,N_8730);
and U9187 (N_9187,N_8955,N_8690);
and U9188 (N_9188,N_8841,N_8510);
and U9189 (N_9189,N_8806,N_8820);
and U9190 (N_9190,N_8997,N_8625);
nand U9191 (N_9191,N_8569,N_8749);
nor U9192 (N_9192,N_8553,N_8571);
nor U9193 (N_9193,N_8563,N_8929);
nor U9194 (N_9194,N_8983,N_8982);
nor U9195 (N_9195,N_8704,N_8575);
nor U9196 (N_9196,N_8858,N_8556);
nand U9197 (N_9197,N_8676,N_8758);
and U9198 (N_9198,N_8904,N_8532);
or U9199 (N_9199,N_8989,N_8916);
nand U9200 (N_9200,N_8594,N_8808);
and U9201 (N_9201,N_8638,N_8584);
and U9202 (N_9202,N_8772,N_8840);
nand U9203 (N_9203,N_8814,N_8628);
nor U9204 (N_9204,N_8785,N_8781);
and U9205 (N_9205,N_8637,N_8652);
nand U9206 (N_9206,N_8846,N_8543);
nor U9207 (N_9207,N_8897,N_8878);
nor U9208 (N_9208,N_8875,N_8966);
and U9209 (N_9209,N_8832,N_8697);
and U9210 (N_9210,N_8761,N_8626);
and U9211 (N_9211,N_8661,N_8779);
xnor U9212 (N_9212,N_8710,N_8595);
or U9213 (N_9213,N_8956,N_8667);
nor U9214 (N_9214,N_8723,N_8593);
nor U9215 (N_9215,N_8910,N_8683);
nor U9216 (N_9216,N_8720,N_8908);
or U9217 (N_9217,N_8890,N_8675);
or U9218 (N_9218,N_8559,N_8653);
nand U9219 (N_9219,N_8658,N_8648);
and U9220 (N_9220,N_8740,N_8636);
nor U9221 (N_9221,N_8733,N_8898);
nand U9222 (N_9222,N_8927,N_8604);
nand U9223 (N_9223,N_8668,N_8801);
and U9224 (N_9224,N_8516,N_8805);
xor U9225 (N_9225,N_8759,N_8754);
nand U9226 (N_9226,N_8566,N_8732);
or U9227 (N_9227,N_8960,N_8766);
and U9228 (N_9228,N_8644,N_8777);
and U9229 (N_9229,N_8859,N_8521);
xor U9230 (N_9230,N_8501,N_8812);
nor U9231 (N_9231,N_8562,N_8809);
nand U9232 (N_9232,N_8685,N_8738);
nor U9233 (N_9233,N_8745,N_8905);
or U9234 (N_9234,N_8976,N_8523);
or U9235 (N_9235,N_8765,N_8873);
or U9236 (N_9236,N_8678,N_8867);
nor U9237 (N_9237,N_8550,N_8610);
and U9238 (N_9238,N_8951,N_8763);
nor U9239 (N_9239,N_8855,N_8871);
nor U9240 (N_9240,N_8942,N_8877);
nor U9241 (N_9241,N_8656,N_8618);
nor U9242 (N_9242,N_8561,N_8700);
nand U9243 (N_9243,N_8609,N_8632);
xnor U9244 (N_9244,N_8944,N_8645);
nand U9245 (N_9245,N_8757,N_8802);
and U9246 (N_9246,N_8939,N_8617);
or U9247 (N_9247,N_8866,N_8776);
and U9248 (N_9248,N_8893,N_8847);
and U9249 (N_9249,N_8901,N_8585);
xnor U9250 (N_9250,N_8914,N_8910);
nor U9251 (N_9251,N_8995,N_8916);
nand U9252 (N_9252,N_8714,N_8804);
or U9253 (N_9253,N_8698,N_8758);
nand U9254 (N_9254,N_8756,N_8981);
or U9255 (N_9255,N_8924,N_8959);
xnor U9256 (N_9256,N_8740,N_8878);
nor U9257 (N_9257,N_8616,N_8655);
nor U9258 (N_9258,N_8769,N_8707);
and U9259 (N_9259,N_8773,N_8656);
and U9260 (N_9260,N_8524,N_8892);
nor U9261 (N_9261,N_8565,N_8522);
or U9262 (N_9262,N_8828,N_8979);
or U9263 (N_9263,N_8668,N_8591);
xor U9264 (N_9264,N_8748,N_8974);
and U9265 (N_9265,N_8784,N_8976);
or U9266 (N_9266,N_8738,N_8915);
xor U9267 (N_9267,N_8992,N_8631);
xnor U9268 (N_9268,N_8605,N_8650);
xor U9269 (N_9269,N_8650,N_8612);
and U9270 (N_9270,N_8889,N_8545);
xnor U9271 (N_9271,N_8518,N_8625);
nand U9272 (N_9272,N_8551,N_8995);
nor U9273 (N_9273,N_8931,N_8788);
or U9274 (N_9274,N_8776,N_8957);
and U9275 (N_9275,N_8901,N_8501);
nor U9276 (N_9276,N_8855,N_8849);
and U9277 (N_9277,N_8803,N_8688);
nor U9278 (N_9278,N_8943,N_8681);
and U9279 (N_9279,N_8749,N_8748);
nor U9280 (N_9280,N_8526,N_8930);
nor U9281 (N_9281,N_8948,N_8981);
and U9282 (N_9282,N_8962,N_8607);
and U9283 (N_9283,N_8566,N_8695);
and U9284 (N_9284,N_8874,N_8852);
xor U9285 (N_9285,N_8672,N_8971);
xnor U9286 (N_9286,N_8695,N_8883);
nor U9287 (N_9287,N_8788,N_8874);
nand U9288 (N_9288,N_8649,N_8821);
xor U9289 (N_9289,N_8727,N_8563);
nor U9290 (N_9290,N_8896,N_8637);
and U9291 (N_9291,N_8526,N_8622);
nand U9292 (N_9292,N_8659,N_8911);
xnor U9293 (N_9293,N_8725,N_8602);
and U9294 (N_9294,N_8791,N_8640);
nor U9295 (N_9295,N_8743,N_8520);
and U9296 (N_9296,N_8784,N_8809);
and U9297 (N_9297,N_8530,N_8643);
xnor U9298 (N_9298,N_8696,N_8806);
xnor U9299 (N_9299,N_8555,N_8570);
and U9300 (N_9300,N_8873,N_8595);
nor U9301 (N_9301,N_8648,N_8601);
nand U9302 (N_9302,N_8815,N_8605);
or U9303 (N_9303,N_8610,N_8723);
and U9304 (N_9304,N_8947,N_8759);
nand U9305 (N_9305,N_8512,N_8533);
nor U9306 (N_9306,N_8852,N_8967);
xnor U9307 (N_9307,N_8848,N_8521);
and U9308 (N_9308,N_8569,N_8983);
or U9309 (N_9309,N_8794,N_8968);
nor U9310 (N_9310,N_8846,N_8507);
and U9311 (N_9311,N_8520,N_8874);
nand U9312 (N_9312,N_8649,N_8853);
and U9313 (N_9313,N_8932,N_8677);
or U9314 (N_9314,N_8768,N_8869);
nand U9315 (N_9315,N_8551,N_8837);
xor U9316 (N_9316,N_8531,N_8720);
nand U9317 (N_9317,N_8673,N_8750);
and U9318 (N_9318,N_8510,N_8543);
xnor U9319 (N_9319,N_8794,N_8891);
nand U9320 (N_9320,N_8960,N_8708);
xnor U9321 (N_9321,N_8911,N_8714);
nand U9322 (N_9322,N_8920,N_8707);
nand U9323 (N_9323,N_8749,N_8867);
nor U9324 (N_9324,N_8983,N_8840);
nor U9325 (N_9325,N_8695,N_8732);
nor U9326 (N_9326,N_8936,N_8862);
and U9327 (N_9327,N_8825,N_8778);
xnor U9328 (N_9328,N_8952,N_8879);
xor U9329 (N_9329,N_8914,N_8565);
nor U9330 (N_9330,N_8651,N_8514);
xor U9331 (N_9331,N_8607,N_8883);
xor U9332 (N_9332,N_8566,N_8910);
nand U9333 (N_9333,N_8878,N_8568);
and U9334 (N_9334,N_8620,N_8688);
xnor U9335 (N_9335,N_8533,N_8915);
nor U9336 (N_9336,N_8763,N_8978);
or U9337 (N_9337,N_8950,N_8627);
and U9338 (N_9338,N_8867,N_8570);
nor U9339 (N_9339,N_8704,N_8720);
and U9340 (N_9340,N_8688,N_8853);
and U9341 (N_9341,N_8660,N_8915);
and U9342 (N_9342,N_8947,N_8741);
or U9343 (N_9343,N_8575,N_8831);
xor U9344 (N_9344,N_8568,N_8565);
nor U9345 (N_9345,N_8996,N_8843);
nand U9346 (N_9346,N_8774,N_8978);
nor U9347 (N_9347,N_8745,N_8722);
nand U9348 (N_9348,N_8850,N_8601);
nand U9349 (N_9349,N_8541,N_8694);
nand U9350 (N_9350,N_8581,N_8506);
or U9351 (N_9351,N_8857,N_8603);
nor U9352 (N_9352,N_8708,N_8937);
nor U9353 (N_9353,N_8619,N_8986);
nor U9354 (N_9354,N_8711,N_8654);
nand U9355 (N_9355,N_8764,N_8852);
nand U9356 (N_9356,N_8798,N_8878);
nor U9357 (N_9357,N_8699,N_8865);
and U9358 (N_9358,N_8999,N_8955);
nor U9359 (N_9359,N_8890,N_8523);
or U9360 (N_9360,N_8859,N_8962);
nor U9361 (N_9361,N_8608,N_8527);
and U9362 (N_9362,N_8538,N_8571);
and U9363 (N_9363,N_8894,N_8777);
and U9364 (N_9364,N_8957,N_8717);
nand U9365 (N_9365,N_8682,N_8535);
xnor U9366 (N_9366,N_8639,N_8653);
xnor U9367 (N_9367,N_8922,N_8822);
or U9368 (N_9368,N_8661,N_8606);
or U9369 (N_9369,N_8980,N_8905);
nand U9370 (N_9370,N_8741,N_8833);
nand U9371 (N_9371,N_8727,N_8882);
and U9372 (N_9372,N_8851,N_8741);
nor U9373 (N_9373,N_8997,N_8845);
xor U9374 (N_9374,N_8891,N_8593);
xnor U9375 (N_9375,N_8733,N_8745);
xnor U9376 (N_9376,N_8947,N_8786);
or U9377 (N_9377,N_8751,N_8607);
nor U9378 (N_9378,N_8878,N_8804);
and U9379 (N_9379,N_8649,N_8907);
nand U9380 (N_9380,N_8666,N_8514);
and U9381 (N_9381,N_8676,N_8705);
xnor U9382 (N_9382,N_8688,N_8550);
nand U9383 (N_9383,N_8850,N_8691);
nand U9384 (N_9384,N_8591,N_8600);
xnor U9385 (N_9385,N_8847,N_8764);
and U9386 (N_9386,N_8821,N_8657);
xnor U9387 (N_9387,N_8651,N_8833);
nand U9388 (N_9388,N_8960,N_8510);
nand U9389 (N_9389,N_8634,N_8923);
and U9390 (N_9390,N_8548,N_8896);
xnor U9391 (N_9391,N_8751,N_8909);
nor U9392 (N_9392,N_8514,N_8539);
or U9393 (N_9393,N_8694,N_8795);
nand U9394 (N_9394,N_8581,N_8794);
xnor U9395 (N_9395,N_8629,N_8917);
nand U9396 (N_9396,N_8877,N_8507);
nor U9397 (N_9397,N_8780,N_8648);
xor U9398 (N_9398,N_8673,N_8703);
and U9399 (N_9399,N_8845,N_8575);
nor U9400 (N_9400,N_8726,N_8682);
xnor U9401 (N_9401,N_8771,N_8715);
nand U9402 (N_9402,N_8621,N_8556);
nor U9403 (N_9403,N_8963,N_8681);
and U9404 (N_9404,N_8610,N_8577);
xnor U9405 (N_9405,N_8993,N_8842);
or U9406 (N_9406,N_8951,N_8919);
nand U9407 (N_9407,N_8672,N_8767);
or U9408 (N_9408,N_8785,N_8881);
nor U9409 (N_9409,N_8954,N_8596);
or U9410 (N_9410,N_8825,N_8933);
nand U9411 (N_9411,N_8974,N_8853);
and U9412 (N_9412,N_8896,N_8761);
or U9413 (N_9413,N_8967,N_8664);
or U9414 (N_9414,N_8555,N_8993);
and U9415 (N_9415,N_8646,N_8976);
nor U9416 (N_9416,N_8958,N_8782);
nor U9417 (N_9417,N_8619,N_8667);
nor U9418 (N_9418,N_8580,N_8679);
nand U9419 (N_9419,N_8998,N_8665);
xnor U9420 (N_9420,N_8540,N_8987);
nor U9421 (N_9421,N_8914,N_8753);
or U9422 (N_9422,N_8750,N_8934);
xnor U9423 (N_9423,N_8807,N_8515);
nor U9424 (N_9424,N_8682,N_8912);
xor U9425 (N_9425,N_8759,N_8615);
xor U9426 (N_9426,N_8646,N_8555);
nand U9427 (N_9427,N_8814,N_8718);
nor U9428 (N_9428,N_8578,N_8672);
xor U9429 (N_9429,N_8615,N_8664);
nor U9430 (N_9430,N_8796,N_8594);
nand U9431 (N_9431,N_8735,N_8793);
or U9432 (N_9432,N_8819,N_8875);
or U9433 (N_9433,N_8972,N_8648);
or U9434 (N_9434,N_8611,N_8751);
and U9435 (N_9435,N_8845,N_8820);
xnor U9436 (N_9436,N_8550,N_8812);
nand U9437 (N_9437,N_8895,N_8552);
or U9438 (N_9438,N_8691,N_8729);
and U9439 (N_9439,N_8685,N_8711);
nand U9440 (N_9440,N_8740,N_8882);
nor U9441 (N_9441,N_8565,N_8858);
or U9442 (N_9442,N_8657,N_8928);
and U9443 (N_9443,N_8845,N_8943);
or U9444 (N_9444,N_8967,N_8607);
and U9445 (N_9445,N_8988,N_8707);
or U9446 (N_9446,N_8969,N_8949);
nand U9447 (N_9447,N_8708,N_8620);
nand U9448 (N_9448,N_8728,N_8850);
and U9449 (N_9449,N_8686,N_8970);
nor U9450 (N_9450,N_8523,N_8702);
nor U9451 (N_9451,N_8576,N_8991);
and U9452 (N_9452,N_8950,N_8644);
nand U9453 (N_9453,N_8956,N_8857);
nand U9454 (N_9454,N_8549,N_8588);
xnor U9455 (N_9455,N_8545,N_8783);
or U9456 (N_9456,N_8896,N_8656);
and U9457 (N_9457,N_8580,N_8959);
xnor U9458 (N_9458,N_8907,N_8995);
nand U9459 (N_9459,N_8927,N_8574);
nand U9460 (N_9460,N_8843,N_8593);
xor U9461 (N_9461,N_8977,N_8887);
nor U9462 (N_9462,N_8931,N_8596);
or U9463 (N_9463,N_8984,N_8847);
nand U9464 (N_9464,N_8749,N_8956);
xor U9465 (N_9465,N_8732,N_8524);
and U9466 (N_9466,N_8970,N_8818);
nor U9467 (N_9467,N_8870,N_8958);
nor U9468 (N_9468,N_8738,N_8722);
xnor U9469 (N_9469,N_8727,N_8815);
or U9470 (N_9470,N_8653,N_8500);
or U9471 (N_9471,N_8593,N_8544);
and U9472 (N_9472,N_8556,N_8750);
and U9473 (N_9473,N_8770,N_8693);
nand U9474 (N_9474,N_8906,N_8627);
nand U9475 (N_9475,N_8851,N_8646);
and U9476 (N_9476,N_8707,N_8712);
or U9477 (N_9477,N_8828,N_8829);
xor U9478 (N_9478,N_8508,N_8778);
or U9479 (N_9479,N_8932,N_8734);
and U9480 (N_9480,N_8590,N_8609);
and U9481 (N_9481,N_8787,N_8790);
or U9482 (N_9482,N_8812,N_8820);
or U9483 (N_9483,N_8573,N_8938);
and U9484 (N_9484,N_8616,N_8534);
nor U9485 (N_9485,N_8742,N_8821);
xor U9486 (N_9486,N_8514,N_8555);
nor U9487 (N_9487,N_8964,N_8890);
xor U9488 (N_9488,N_8748,N_8639);
xor U9489 (N_9489,N_8795,N_8753);
nor U9490 (N_9490,N_8884,N_8677);
nand U9491 (N_9491,N_8672,N_8982);
nand U9492 (N_9492,N_8665,N_8571);
nor U9493 (N_9493,N_8946,N_8514);
and U9494 (N_9494,N_8840,N_8822);
or U9495 (N_9495,N_8631,N_8680);
nand U9496 (N_9496,N_8913,N_8845);
or U9497 (N_9497,N_8623,N_8877);
nor U9498 (N_9498,N_8800,N_8843);
nand U9499 (N_9499,N_8936,N_8832);
nor U9500 (N_9500,N_9445,N_9274);
xnor U9501 (N_9501,N_9298,N_9493);
xnor U9502 (N_9502,N_9201,N_9376);
and U9503 (N_9503,N_9122,N_9154);
and U9504 (N_9504,N_9343,N_9346);
nand U9505 (N_9505,N_9347,N_9296);
and U9506 (N_9506,N_9246,N_9242);
xnor U9507 (N_9507,N_9489,N_9425);
xnor U9508 (N_9508,N_9208,N_9049);
xnor U9509 (N_9509,N_9216,N_9000);
and U9510 (N_9510,N_9041,N_9476);
nand U9511 (N_9511,N_9318,N_9410);
or U9512 (N_9512,N_9002,N_9282);
or U9513 (N_9513,N_9147,N_9072);
nand U9514 (N_9514,N_9052,N_9170);
and U9515 (N_9515,N_9075,N_9311);
xnor U9516 (N_9516,N_9183,N_9111);
nand U9517 (N_9517,N_9247,N_9300);
nor U9518 (N_9518,N_9426,N_9283);
nand U9519 (N_9519,N_9254,N_9007);
nand U9520 (N_9520,N_9448,N_9320);
or U9521 (N_9521,N_9357,N_9179);
and U9522 (N_9522,N_9088,N_9317);
and U9523 (N_9523,N_9329,N_9397);
xnor U9524 (N_9524,N_9125,N_9023);
xor U9525 (N_9525,N_9387,N_9288);
xor U9526 (N_9526,N_9197,N_9146);
xnor U9527 (N_9527,N_9182,N_9020);
nand U9528 (N_9528,N_9248,N_9130);
or U9529 (N_9529,N_9290,N_9071);
nand U9530 (N_9530,N_9332,N_9095);
xor U9531 (N_9531,N_9386,N_9018);
or U9532 (N_9532,N_9098,N_9084);
or U9533 (N_9533,N_9213,N_9359);
and U9534 (N_9534,N_9207,N_9136);
and U9535 (N_9535,N_9110,N_9285);
nor U9536 (N_9536,N_9228,N_9243);
or U9537 (N_9537,N_9444,N_9077);
and U9538 (N_9538,N_9336,N_9356);
and U9539 (N_9539,N_9087,N_9051);
nor U9540 (N_9540,N_9458,N_9379);
nand U9541 (N_9541,N_9139,N_9280);
nand U9542 (N_9542,N_9423,N_9424);
xor U9543 (N_9543,N_9019,N_9177);
or U9544 (N_9544,N_9085,N_9488);
nand U9545 (N_9545,N_9468,N_9331);
nand U9546 (N_9546,N_9160,N_9099);
nand U9547 (N_9547,N_9017,N_9200);
xnor U9548 (N_9548,N_9047,N_9112);
or U9549 (N_9549,N_9148,N_9039);
nor U9550 (N_9550,N_9005,N_9116);
xor U9551 (N_9551,N_9048,N_9355);
nor U9552 (N_9552,N_9025,N_9297);
nand U9553 (N_9553,N_9181,N_9178);
nand U9554 (N_9554,N_9212,N_9471);
and U9555 (N_9555,N_9313,N_9496);
and U9556 (N_9556,N_9241,N_9202);
nand U9557 (N_9557,N_9255,N_9367);
or U9558 (N_9558,N_9138,N_9481);
nand U9559 (N_9559,N_9253,N_9231);
nor U9560 (N_9560,N_9074,N_9024);
nor U9561 (N_9561,N_9368,N_9454);
or U9562 (N_9562,N_9264,N_9121);
xor U9563 (N_9563,N_9319,N_9028);
and U9564 (N_9564,N_9119,N_9302);
nor U9565 (N_9565,N_9133,N_9321);
xnor U9566 (N_9566,N_9350,N_9413);
nor U9567 (N_9567,N_9187,N_9362);
and U9568 (N_9568,N_9268,N_9330);
nor U9569 (N_9569,N_9045,N_9279);
or U9570 (N_9570,N_9064,N_9295);
nand U9571 (N_9571,N_9272,N_9161);
or U9572 (N_9572,N_9401,N_9115);
nand U9573 (N_9573,N_9262,N_9103);
or U9574 (N_9574,N_9309,N_9046);
or U9575 (N_9575,N_9276,N_9456);
and U9576 (N_9576,N_9173,N_9435);
xor U9577 (N_9577,N_9478,N_9096);
nand U9578 (N_9578,N_9114,N_9155);
nand U9579 (N_9579,N_9428,N_9440);
nor U9580 (N_9580,N_9480,N_9249);
and U9581 (N_9581,N_9037,N_9433);
or U9582 (N_9582,N_9061,N_9301);
nor U9583 (N_9583,N_9180,N_9384);
nand U9584 (N_9584,N_9315,N_9162);
nor U9585 (N_9585,N_9093,N_9135);
nor U9586 (N_9586,N_9391,N_9159);
nand U9587 (N_9587,N_9223,N_9150);
and U9588 (N_9588,N_9271,N_9165);
and U9589 (N_9589,N_9073,N_9040);
and U9590 (N_9590,N_9123,N_9273);
nor U9591 (N_9591,N_9153,N_9059);
xor U9592 (N_9592,N_9070,N_9237);
xnor U9593 (N_9593,N_9167,N_9034);
or U9594 (N_9594,N_9191,N_9469);
or U9595 (N_9595,N_9461,N_9172);
nor U9596 (N_9596,N_9383,N_9326);
or U9597 (N_9597,N_9199,N_9217);
xor U9598 (N_9598,N_9221,N_9451);
or U9599 (N_9599,N_9261,N_9265);
nor U9600 (N_9600,N_9141,N_9432);
xnor U9601 (N_9601,N_9094,N_9239);
xor U9602 (N_9602,N_9081,N_9335);
xnor U9603 (N_9603,N_9224,N_9475);
xor U9604 (N_9604,N_9235,N_9486);
nand U9605 (N_9605,N_9310,N_9342);
xor U9606 (N_9606,N_9405,N_9232);
and U9607 (N_9607,N_9462,N_9079);
nor U9608 (N_9608,N_9464,N_9057);
xnor U9609 (N_9609,N_9403,N_9184);
nand U9610 (N_9610,N_9101,N_9375);
nand U9611 (N_9611,N_9299,N_9055);
xor U9612 (N_9612,N_9487,N_9370);
xnor U9613 (N_9613,N_9108,N_9015);
and U9614 (N_9614,N_9149,N_9473);
or U9615 (N_9615,N_9082,N_9441);
nand U9616 (N_9616,N_9465,N_9490);
and U9617 (N_9617,N_9113,N_9186);
nor U9618 (N_9618,N_9419,N_9080);
or U9619 (N_9619,N_9427,N_9286);
nand U9620 (N_9620,N_9474,N_9304);
and U9621 (N_9621,N_9090,N_9230);
nand U9622 (N_9622,N_9120,N_9291);
or U9623 (N_9623,N_9270,N_9078);
and U9624 (N_9624,N_9126,N_9043);
or U9625 (N_9625,N_9348,N_9013);
xor U9626 (N_9626,N_9158,N_9219);
nand U9627 (N_9627,N_9409,N_9325);
nand U9628 (N_9628,N_9229,N_9227);
nand U9629 (N_9629,N_9267,N_9214);
and U9630 (N_9630,N_9430,N_9118);
nand U9631 (N_9631,N_9014,N_9164);
and U9632 (N_9632,N_9374,N_9281);
nor U9633 (N_9633,N_9363,N_9257);
or U9634 (N_9634,N_9222,N_9065);
xnor U9635 (N_9635,N_9022,N_9289);
xnor U9636 (N_9636,N_9328,N_9463);
nand U9637 (N_9637,N_9422,N_9420);
and U9638 (N_9638,N_9189,N_9127);
nor U9639 (N_9639,N_9009,N_9226);
nor U9640 (N_9640,N_9132,N_9244);
nor U9641 (N_9641,N_9238,N_9069);
xor U9642 (N_9642,N_9196,N_9381);
nand U9643 (N_9643,N_9377,N_9482);
or U9644 (N_9644,N_9408,N_9275);
and U9645 (N_9645,N_9091,N_9131);
or U9646 (N_9646,N_9354,N_9016);
and U9647 (N_9647,N_9142,N_9156);
or U9648 (N_9648,N_9263,N_9305);
and U9649 (N_9649,N_9452,N_9042);
nor U9650 (N_9650,N_9442,N_9412);
nor U9651 (N_9651,N_9012,N_9259);
and U9652 (N_9652,N_9446,N_9307);
and U9653 (N_9653,N_9483,N_9416);
or U9654 (N_9654,N_9027,N_9100);
or U9655 (N_9655,N_9373,N_9011);
and U9656 (N_9656,N_9056,N_9415);
nor U9657 (N_9657,N_9010,N_9092);
or U9658 (N_9658,N_9021,N_9004);
xor U9659 (N_9659,N_9245,N_9492);
xor U9660 (N_9660,N_9431,N_9421);
and U9661 (N_9661,N_9068,N_9215);
or U9662 (N_9662,N_9392,N_9236);
xor U9663 (N_9663,N_9459,N_9322);
and U9664 (N_9664,N_9358,N_9411);
or U9665 (N_9665,N_9001,N_9060);
xor U9666 (N_9666,N_9434,N_9292);
nand U9667 (N_9667,N_9107,N_9390);
or U9668 (N_9668,N_9455,N_9117);
nand U9669 (N_9669,N_9366,N_9352);
nand U9670 (N_9670,N_9175,N_9349);
nor U9671 (N_9671,N_9385,N_9378);
xnor U9672 (N_9672,N_9460,N_9364);
nand U9673 (N_9673,N_9063,N_9449);
nand U9674 (N_9674,N_9157,N_9417);
or U9675 (N_9675,N_9109,N_9256);
or U9676 (N_9676,N_9033,N_9333);
xor U9677 (N_9677,N_9437,N_9031);
or U9678 (N_9678,N_9233,N_9220);
or U9679 (N_9679,N_9171,N_9436);
nor U9680 (N_9680,N_9260,N_9076);
xor U9681 (N_9681,N_9128,N_9407);
nand U9682 (N_9682,N_9185,N_9396);
xor U9683 (N_9683,N_9163,N_9457);
xnor U9684 (N_9684,N_9176,N_9168);
and U9685 (N_9685,N_9404,N_9470);
and U9686 (N_9686,N_9388,N_9209);
nor U9687 (N_9687,N_9479,N_9102);
nor U9688 (N_9688,N_9344,N_9036);
or U9689 (N_9689,N_9303,N_9269);
and U9690 (N_9690,N_9026,N_9193);
or U9691 (N_9691,N_9466,N_9351);
nand U9692 (N_9692,N_9053,N_9395);
xor U9693 (N_9693,N_9205,N_9341);
xor U9694 (N_9694,N_9394,N_9306);
or U9695 (N_9695,N_9365,N_9277);
or U9696 (N_9696,N_9083,N_9323);
nor U9697 (N_9697,N_9287,N_9258);
xnor U9698 (N_9698,N_9204,N_9006);
or U9699 (N_9699,N_9369,N_9485);
nand U9700 (N_9700,N_9278,N_9089);
nand U9701 (N_9701,N_9467,N_9316);
nand U9702 (N_9702,N_9166,N_9003);
or U9703 (N_9703,N_9145,N_9308);
and U9704 (N_9704,N_9495,N_9151);
nor U9705 (N_9705,N_9058,N_9169);
or U9706 (N_9706,N_9406,N_9044);
xor U9707 (N_9707,N_9340,N_9438);
nor U9708 (N_9708,N_9453,N_9327);
xnor U9709 (N_9709,N_9443,N_9345);
and U9710 (N_9710,N_9477,N_9030);
xnor U9711 (N_9711,N_9174,N_9097);
xor U9712 (N_9712,N_9314,N_9491);
nor U9713 (N_9713,N_9414,N_9372);
nand U9714 (N_9714,N_9393,N_9353);
or U9715 (N_9715,N_9266,N_9293);
and U9716 (N_9716,N_9198,N_9211);
xnor U9717 (N_9717,N_9054,N_9137);
nand U9718 (N_9718,N_9339,N_9399);
and U9719 (N_9719,N_9494,N_9140);
nor U9720 (N_9720,N_9206,N_9250);
nand U9721 (N_9721,N_9062,N_9400);
nand U9722 (N_9722,N_9143,N_9499);
or U9723 (N_9723,N_9398,N_9035);
or U9724 (N_9724,N_9134,N_9324);
xnor U9725 (N_9725,N_9360,N_9447);
or U9726 (N_9726,N_9144,N_9402);
nor U9727 (N_9727,N_9029,N_9251);
xor U9728 (N_9728,N_9195,N_9429);
xor U9729 (N_9729,N_9450,N_9067);
and U9730 (N_9730,N_9338,N_9152);
xor U9731 (N_9731,N_9389,N_9050);
nand U9732 (N_9732,N_9190,N_9008);
or U9733 (N_9733,N_9225,N_9371);
nor U9734 (N_9734,N_9192,N_9104);
xor U9735 (N_9735,N_9124,N_9472);
or U9736 (N_9736,N_9086,N_9203);
nand U9737 (N_9737,N_9129,N_9361);
or U9738 (N_9738,N_9380,N_9240);
nand U9739 (N_9739,N_9210,N_9105);
nor U9740 (N_9740,N_9418,N_9194);
nand U9741 (N_9741,N_9382,N_9038);
xnor U9742 (N_9742,N_9066,N_9284);
and U9743 (N_9743,N_9234,N_9484);
xnor U9744 (N_9744,N_9498,N_9252);
nand U9745 (N_9745,N_9032,N_9439);
or U9746 (N_9746,N_9334,N_9497);
nor U9747 (N_9747,N_9294,N_9312);
and U9748 (N_9748,N_9106,N_9188);
nor U9749 (N_9749,N_9218,N_9337);
xnor U9750 (N_9750,N_9291,N_9294);
or U9751 (N_9751,N_9207,N_9361);
xor U9752 (N_9752,N_9222,N_9329);
nand U9753 (N_9753,N_9005,N_9327);
nor U9754 (N_9754,N_9081,N_9273);
and U9755 (N_9755,N_9057,N_9408);
nand U9756 (N_9756,N_9015,N_9093);
xnor U9757 (N_9757,N_9167,N_9151);
or U9758 (N_9758,N_9192,N_9298);
nor U9759 (N_9759,N_9183,N_9172);
or U9760 (N_9760,N_9418,N_9223);
xnor U9761 (N_9761,N_9480,N_9148);
nand U9762 (N_9762,N_9219,N_9097);
nand U9763 (N_9763,N_9005,N_9104);
or U9764 (N_9764,N_9178,N_9156);
nand U9765 (N_9765,N_9237,N_9322);
xor U9766 (N_9766,N_9111,N_9440);
and U9767 (N_9767,N_9458,N_9265);
nand U9768 (N_9768,N_9469,N_9030);
xnor U9769 (N_9769,N_9155,N_9015);
or U9770 (N_9770,N_9213,N_9266);
or U9771 (N_9771,N_9215,N_9219);
or U9772 (N_9772,N_9468,N_9397);
and U9773 (N_9773,N_9315,N_9095);
xnor U9774 (N_9774,N_9021,N_9276);
and U9775 (N_9775,N_9275,N_9284);
xnor U9776 (N_9776,N_9498,N_9283);
nor U9777 (N_9777,N_9365,N_9248);
or U9778 (N_9778,N_9200,N_9379);
nand U9779 (N_9779,N_9283,N_9390);
and U9780 (N_9780,N_9161,N_9409);
and U9781 (N_9781,N_9442,N_9329);
nor U9782 (N_9782,N_9060,N_9295);
and U9783 (N_9783,N_9220,N_9270);
or U9784 (N_9784,N_9182,N_9168);
xor U9785 (N_9785,N_9438,N_9150);
and U9786 (N_9786,N_9119,N_9065);
xor U9787 (N_9787,N_9396,N_9401);
nand U9788 (N_9788,N_9007,N_9487);
xor U9789 (N_9789,N_9161,N_9480);
xor U9790 (N_9790,N_9297,N_9186);
xor U9791 (N_9791,N_9456,N_9322);
nand U9792 (N_9792,N_9129,N_9090);
xnor U9793 (N_9793,N_9328,N_9000);
or U9794 (N_9794,N_9398,N_9356);
nor U9795 (N_9795,N_9277,N_9495);
and U9796 (N_9796,N_9250,N_9349);
or U9797 (N_9797,N_9341,N_9121);
or U9798 (N_9798,N_9006,N_9412);
or U9799 (N_9799,N_9009,N_9280);
nor U9800 (N_9800,N_9041,N_9450);
or U9801 (N_9801,N_9463,N_9382);
or U9802 (N_9802,N_9371,N_9054);
and U9803 (N_9803,N_9080,N_9083);
xor U9804 (N_9804,N_9130,N_9063);
nand U9805 (N_9805,N_9178,N_9152);
and U9806 (N_9806,N_9483,N_9189);
and U9807 (N_9807,N_9499,N_9307);
xor U9808 (N_9808,N_9131,N_9188);
or U9809 (N_9809,N_9135,N_9427);
or U9810 (N_9810,N_9451,N_9241);
nor U9811 (N_9811,N_9178,N_9018);
xnor U9812 (N_9812,N_9437,N_9306);
xnor U9813 (N_9813,N_9334,N_9414);
nand U9814 (N_9814,N_9333,N_9203);
and U9815 (N_9815,N_9295,N_9236);
or U9816 (N_9816,N_9135,N_9315);
nand U9817 (N_9817,N_9038,N_9307);
xor U9818 (N_9818,N_9208,N_9241);
and U9819 (N_9819,N_9098,N_9152);
and U9820 (N_9820,N_9238,N_9234);
and U9821 (N_9821,N_9387,N_9484);
or U9822 (N_9822,N_9239,N_9262);
nor U9823 (N_9823,N_9310,N_9266);
and U9824 (N_9824,N_9490,N_9364);
and U9825 (N_9825,N_9306,N_9484);
nand U9826 (N_9826,N_9396,N_9054);
nand U9827 (N_9827,N_9137,N_9199);
nor U9828 (N_9828,N_9462,N_9215);
and U9829 (N_9829,N_9391,N_9149);
and U9830 (N_9830,N_9143,N_9337);
xnor U9831 (N_9831,N_9122,N_9269);
xnor U9832 (N_9832,N_9324,N_9319);
xnor U9833 (N_9833,N_9149,N_9443);
nor U9834 (N_9834,N_9230,N_9470);
and U9835 (N_9835,N_9155,N_9001);
and U9836 (N_9836,N_9389,N_9198);
xnor U9837 (N_9837,N_9023,N_9308);
xnor U9838 (N_9838,N_9346,N_9113);
xnor U9839 (N_9839,N_9327,N_9115);
and U9840 (N_9840,N_9168,N_9383);
and U9841 (N_9841,N_9153,N_9000);
nand U9842 (N_9842,N_9115,N_9043);
xor U9843 (N_9843,N_9379,N_9226);
xnor U9844 (N_9844,N_9053,N_9067);
or U9845 (N_9845,N_9284,N_9090);
nand U9846 (N_9846,N_9140,N_9110);
and U9847 (N_9847,N_9254,N_9304);
and U9848 (N_9848,N_9055,N_9251);
nor U9849 (N_9849,N_9031,N_9281);
nand U9850 (N_9850,N_9015,N_9235);
or U9851 (N_9851,N_9003,N_9302);
and U9852 (N_9852,N_9498,N_9475);
xor U9853 (N_9853,N_9447,N_9481);
nand U9854 (N_9854,N_9495,N_9183);
or U9855 (N_9855,N_9388,N_9446);
nand U9856 (N_9856,N_9165,N_9460);
or U9857 (N_9857,N_9102,N_9058);
xnor U9858 (N_9858,N_9018,N_9015);
or U9859 (N_9859,N_9152,N_9156);
xnor U9860 (N_9860,N_9413,N_9219);
or U9861 (N_9861,N_9104,N_9259);
or U9862 (N_9862,N_9005,N_9450);
xnor U9863 (N_9863,N_9371,N_9342);
nor U9864 (N_9864,N_9357,N_9457);
nor U9865 (N_9865,N_9419,N_9267);
and U9866 (N_9866,N_9387,N_9109);
and U9867 (N_9867,N_9000,N_9011);
and U9868 (N_9868,N_9482,N_9487);
or U9869 (N_9869,N_9257,N_9240);
nand U9870 (N_9870,N_9204,N_9017);
xnor U9871 (N_9871,N_9116,N_9478);
nand U9872 (N_9872,N_9205,N_9216);
nor U9873 (N_9873,N_9079,N_9400);
xnor U9874 (N_9874,N_9054,N_9289);
nor U9875 (N_9875,N_9202,N_9146);
nor U9876 (N_9876,N_9144,N_9001);
and U9877 (N_9877,N_9425,N_9468);
nor U9878 (N_9878,N_9407,N_9317);
nand U9879 (N_9879,N_9314,N_9174);
nor U9880 (N_9880,N_9427,N_9417);
or U9881 (N_9881,N_9197,N_9099);
xnor U9882 (N_9882,N_9195,N_9382);
nand U9883 (N_9883,N_9271,N_9066);
nor U9884 (N_9884,N_9284,N_9391);
and U9885 (N_9885,N_9332,N_9394);
nand U9886 (N_9886,N_9237,N_9129);
and U9887 (N_9887,N_9467,N_9466);
or U9888 (N_9888,N_9129,N_9083);
or U9889 (N_9889,N_9416,N_9446);
xor U9890 (N_9890,N_9333,N_9498);
xnor U9891 (N_9891,N_9404,N_9323);
nand U9892 (N_9892,N_9362,N_9451);
and U9893 (N_9893,N_9467,N_9109);
xor U9894 (N_9894,N_9098,N_9427);
xor U9895 (N_9895,N_9152,N_9125);
nor U9896 (N_9896,N_9327,N_9368);
nand U9897 (N_9897,N_9199,N_9154);
xor U9898 (N_9898,N_9194,N_9486);
xnor U9899 (N_9899,N_9325,N_9074);
xor U9900 (N_9900,N_9492,N_9303);
or U9901 (N_9901,N_9160,N_9489);
or U9902 (N_9902,N_9041,N_9485);
and U9903 (N_9903,N_9407,N_9434);
or U9904 (N_9904,N_9104,N_9441);
or U9905 (N_9905,N_9392,N_9161);
or U9906 (N_9906,N_9236,N_9131);
nand U9907 (N_9907,N_9121,N_9240);
and U9908 (N_9908,N_9199,N_9338);
or U9909 (N_9909,N_9439,N_9173);
or U9910 (N_9910,N_9388,N_9264);
and U9911 (N_9911,N_9318,N_9045);
xnor U9912 (N_9912,N_9127,N_9172);
xnor U9913 (N_9913,N_9275,N_9070);
xor U9914 (N_9914,N_9362,N_9119);
and U9915 (N_9915,N_9413,N_9018);
xnor U9916 (N_9916,N_9363,N_9336);
nor U9917 (N_9917,N_9458,N_9238);
nand U9918 (N_9918,N_9452,N_9465);
nor U9919 (N_9919,N_9448,N_9197);
or U9920 (N_9920,N_9056,N_9061);
or U9921 (N_9921,N_9282,N_9043);
nor U9922 (N_9922,N_9305,N_9269);
nor U9923 (N_9923,N_9321,N_9418);
or U9924 (N_9924,N_9252,N_9138);
and U9925 (N_9925,N_9352,N_9213);
xnor U9926 (N_9926,N_9093,N_9205);
and U9927 (N_9927,N_9352,N_9117);
and U9928 (N_9928,N_9483,N_9336);
or U9929 (N_9929,N_9196,N_9265);
and U9930 (N_9930,N_9314,N_9480);
xnor U9931 (N_9931,N_9062,N_9486);
and U9932 (N_9932,N_9349,N_9253);
xor U9933 (N_9933,N_9458,N_9086);
nor U9934 (N_9934,N_9439,N_9232);
or U9935 (N_9935,N_9286,N_9084);
nand U9936 (N_9936,N_9479,N_9477);
or U9937 (N_9937,N_9058,N_9124);
or U9938 (N_9938,N_9364,N_9280);
and U9939 (N_9939,N_9296,N_9159);
nor U9940 (N_9940,N_9108,N_9091);
xor U9941 (N_9941,N_9339,N_9458);
xnor U9942 (N_9942,N_9378,N_9040);
and U9943 (N_9943,N_9122,N_9303);
or U9944 (N_9944,N_9148,N_9280);
or U9945 (N_9945,N_9036,N_9471);
nand U9946 (N_9946,N_9063,N_9209);
or U9947 (N_9947,N_9384,N_9028);
nand U9948 (N_9948,N_9009,N_9243);
xor U9949 (N_9949,N_9220,N_9475);
nand U9950 (N_9950,N_9087,N_9119);
or U9951 (N_9951,N_9353,N_9270);
or U9952 (N_9952,N_9281,N_9478);
xnor U9953 (N_9953,N_9347,N_9287);
nor U9954 (N_9954,N_9139,N_9169);
nor U9955 (N_9955,N_9409,N_9358);
nor U9956 (N_9956,N_9128,N_9331);
nand U9957 (N_9957,N_9000,N_9289);
and U9958 (N_9958,N_9259,N_9263);
or U9959 (N_9959,N_9385,N_9442);
nand U9960 (N_9960,N_9497,N_9100);
or U9961 (N_9961,N_9116,N_9437);
or U9962 (N_9962,N_9140,N_9421);
xor U9963 (N_9963,N_9382,N_9316);
nand U9964 (N_9964,N_9060,N_9247);
nand U9965 (N_9965,N_9425,N_9263);
nor U9966 (N_9966,N_9293,N_9287);
and U9967 (N_9967,N_9454,N_9421);
and U9968 (N_9968,N_9358,N_9278);
or U9969 (N_9969,N_9080,N_9269);
nand U9970 (N_9970,N_9441,N_9331);
and U9971 (N_9971,N_9039,N_9180);
or U9972 (N_9972,N_9412,N_9033);
xnor U9973 (N_9973,N_9152,N_9316);
or U9974 (N_9974,N_9106,N_9439);
or U9975 (N_9975,N_9389,N_9210);
or U9976 (N_9976,N_9025,N_9245);
and U9977 (N_9977,N_9131,N_9241);
nand U9978 (N_9978,N_9342,N_9204);
or U9979 (N_9979,N_9298,N_9318);
and U9980 (N_9980,N_9018,N_9025);
or U9981 (N_9981,N_9433,N_9114);
and U9982 (N_9982,N_9456,N_9079);
or U9983 (N_9983,N_9276,N_9041);
and U9984 (N_9984,N_9448,N_9015);
nor U9985 (N_9985,N_9004,N_9496);
nor U9986 (N_9986,N_9482,N_9340);
or U9987 (N_9987,N_9298,N_9459);
and U9988 (N_9988,N_9273,N_9397);
nand U9989 (N_9989,N_9387,N_9430);
nor U9990 (N_9990,N_9081,N_9139);
and U9991 (N_9991,N_9356,N_9388);
nor U9992 (N_9992,N_9148,N_9220);
xnor U9993 (N_9993,N_9495,N_9351);
nand U9994 (N_9994,N_9317,N_9452);
nand U9995 (N_9995,N_9418,N_9334);
nand U9996 (N_9996,N_9337,N_9093);
nor U9997 (N_9997,N_9211,N_9299);
or U9998 (N_9998,N_9204,N_9449);
xor U9999 (N_9999,N_9422,N_9160);
xor U10000 (N_10000,N_9883,N_9723);
nand U10001 (N_10001,N_9540,N_9682);
nand U10002 (N_10002,N_9502,N_9720);
or U10003 (N_10003,N_9640,N_9725);
nand U10004 (N_10004,N_9577,N_9797);
and U10005 (N_10005,N_9510,N_9798);
xor U10006 (N_10006,N_9863,N_9922);
xnor U10007 (N_10007,N_9971,N_9851);
and U10008 (N_10008,N_9748,N_9956);
nand U10009 (N_10009,N_9561,N_9930);
or U10010 (N_10010,N_9519,N_9989);
xnor U10011 (N_10011,N_9882,N_9943);
or U10012 (N_10012,N_9981,N_9909);
and U10013 (N_10013,N_9539,N_9856);
nand U10014 (N_10014,N_9733,N_9941);
xnor U10015 (N_10015,N_9508,N_9694);
nor U10016 (N_10016,N_9554,N_9859);
xor U10017 (N_10017,N_9513,N_9946);
or U10018 (N_10018,N_9902,N_9764);
xor U10019 (N_10019,N_9611,N_9945);
and U10020 (N_10020,N_9904,N_9613);
or U10021 (N_10021,N_9881,N_9954);
nand U10022 (N_10022,N_9993,N_9701);
nor U10023 (N_10023,N_9610,N_9911);
nor U10024 (N_10024,N_9855,N_9949);
nor U10025 (N_10025,N_9889,N_9848);
or U10026 (N_10026,N_9573,N_9631);
and U10027 (N_10027,N_9576,N_9766);
nor U10028 (N_10028,N_9826,N_9567);
xor U10029 (N_10029,N_9521,N_9982);
nand U10030 (N_10030,N_9762,N_9532);
nor U10031 (N_10031,N_9799,N_9660);
nor U10032 (N_10032,N_9979,N_9794);
nor U10033 (N_10033,N_9505,N_9822);
or U10034 (N_10034,N_9808,N_9780);
and U10035 (N_10035,N_9783,N_9589);
nor U10036 (N_10036,N_9538,N_9996);
or U10037 (N_10037,N_9973,N_9663);
nand U10038 (N_10038,N_9927,N_9583);
or U10039 (N_10039,N_9626,N_9813);
or U10040 (N_10040,N_9793,N_9671);
nand U10041 (N_10041,N_9667,N_9807);
nor U10042 (N_10042,N_9568,N_9959);
or U10043 (N_10043,N_9509,N_9637);
or U10044 (N_10044,N_9575,N_9974);
nand U10045 (N_10045,N_9620,N_9650);
nand U10046 (N_10046,N_9885,N_9999);
or U10047 (N_10047,N_9534,N_9920);
nor U10048 (N_10048,N_9767,N_9892);
nor U10049 (N_10049,N_9811,N_9511);
or U10050 (N_10050,N_9714,N_9659);
nor U10051 (N_10051,N_9960,N_9925);
xnor U10052 (N_10052,N_9668,N_9695);
nand U10053 (N_10053,N_9845,N_9501);
and U10054 (N_10054,N_9983,N_9543);
nand U10055 (N_10055,N_9756,N_9947);
or U10056 (N_10056,N_9565,N_9835);
xnor U10057 (N_10057,N_9921,N_9523);
and U10058 (N_10058,N_9522,N_9586);
and U10059 (N_10059,N_9761,N_9884);
or U10060 (N_10060,N_9929,N_9709);
xnor U10061 (N_10061,N_9912,N_9782);
nand U10062 (N_10062,N_9751,N_9990);
or U10063 (N_10063,N_9938,N_9553);
or U10064 (N_10064,N_9646,N_9515);
xnor U10065 (N_10065,N_9525,N_9997);
nand U10066 (N_10066,N_9831,N_9816);
xnor U10067 (N_10067,N_9609,N_9803);
nor U10068 (N_10068,N_9872,N_9625);
nor U10069 (N_10069,N_9757,N_9692);
nand U10070 (N_10070,N_9924,N_9587);
nor U10071 (N_10071,N_9721,N_9559);
nand U10072 (N_10072,N_9791,N_9641);
nor U10073 (N_10073,N_9604,N_9870);
xor U10074 (N_10074,N_9690,N_9893);
xor U10075 (N_10075,N_9994,N_9735);
and U10076 (N_10076,N_9627,N_9548);
or U10077 (N_10077,N_9940,N_9864);
nand U10078 (N_10078,N_9616,N_9693);
xnor U10079 (N_10079,N_9828,N_9744);
xnor U10080 (N_10080,N_9662,N_9913);
or U10081 (N_10081,N_9524,N_9978);
nand U10082 (N_10082,N_9503,N_9857);
nand U10083 (N_10083,N_9526,N_9887);
or U10084 (N_10084,N_9869,N_9873);
or U10085 (N_10085,N_9507,N_9677);
nand U10086 (N_10086,N_9774,N_9699);
nor U10087 (N_10087,N_9908,N_9991);
nor U10088 (N_10088,N_9585,N_9608);
and U10089 (N_10089,N_9739,N_9837);
and U10090 (N_10090,N_9944,N_9528);
xnor U10091 (N_10091,N_9942,N_9633);
xor U10092 (N_10092,N_9648,N_9987);
and U10093 (N_10093,N_9652,N_9895);
and U10094 (N_10094,N_9917,N_9622);
and U10095 (N_10095,N_9854,N_9800);
and U10096 (N_10096,N_9552,N_9918);
and U10097 (N_10097,N_9814,N_9939);
nor U10098 (N_10098,N_9747,N_9796);
and U10099 (N_10099,N_9644,N_9988);
nor U10100 (N_10100,N_9728,N_9995);
nor U10101 (N_10101,N_9719,N_9726);
and U10102 (N_10102,N_9876,N_9969);
nor U10103 (N_10103,N_9787,N_9986);
nand U10104 (N_10104,N_9936,N_9676);
and U10105 (N_10105,N_9951,N_9642);
nor U10106 (N_10106,N_9636,N_9520);
xor U10107 (N_10107,N_9878,N_9843);
nand U10108 (N_10108,N_9562,N_9823);
and U10109 (N_10109,N_9778,N_9672);
xor U10110 (N_10110,N_9957,N_9666);
or U10111 (N_10111,N_9697,N_9915);
and U10112 (N_10112,N_9590,N_9612);
nand U10113 (N_10113,N_9775,N_9619);
nor U10114 (N_10114,N_9817,N_9792);
nand U10115 (N_10115,N_9679,N_9673);
and U10116 (N_10116,N_9500,N_9952);
or U10117 (N_10117,N_9910,N_9829);
and U10118 (N_10118,N_9834,N_9703);
nand U10119 (N_10119,N_9727,N_9595);
xnor U10120 (N_10120,N_9962,N_9614);
nor U10121 (N_10121,N_9606,N_9740);
or U10122 (N_10122,N_9953,N_9842);
and U10123 (N_10123,N_9923,N_9742);
xnor U10124 (N_10124,N_9691,N_9839);
nor U10125 (N_10125,N_9886,N_9897);
xor U10126 (N_10126,N_9985,N_9746);
or U10127 (N_10127,N_9836,N_9722);
nor U10128 (N_10128,N_9686,N_9602);
xnor U10129 (N_10129,N_9972,N_9970);
and U10130 (N_10130,N_9732,N_9653);
xor U10131 (N_10131,N_9853,N_9900);
or U10132 (N_10132,N_9518,N_9651);
nand U10133 (N_10133,N_9765,N_9984);
or U10134 (N_10134,N_9874,N_9901);
xnor U10135 (N_10135,N_9516,N_9621);
or U10136 (N_10136,N_9711,N_9809);
nor U10137 (N_10137,N_9533,N_9632);
xor U10138 (N_10138,N_9950,N_9629);
and U10139 (N_10139,N_9580,N_9541);
nor U10140 (N_10140,N_9934,N_9749);
nor U10141 (N_10141,N_9880,N_9593);
or U10142 (N_10142,N_9907,N_9514);
or U10143 (N_10143,N_9704,N_9750);
nand U10144 (N_10144,N_9932,N_9926);
nand U10145 (N_10145,N_9681,N_9877);
and U10146 (N_10146,N_9708,N_9617);
and U10147 (N_10147,N_9805,N_9731);
nand U10148 (N_10148,N_9958,N_9647);
or U10149 (N_10149,N_9825,N_9919);
xnor U10150 (N_10150,N_9850,N_9776);
nor U10151 (N_10151,N_9928,N_9574);
or U10152 (N_10152,N_9894,N_9675);
nand U10153 (N_10153,N_9866,N_9964);
or U10154 (N_10154,N_9801,N_9753);
nand U10155 (N_10155,N_9896,N_9706);
nand U10156 (N_10156,N_9737,N_9598);
nor U10157 (N_10157,N_9584,N_9862);
xor U10158 (N_10158,N_9578,N_9785);
and U10159 (N_10159,N_9537,N_9821);
or U10160 (N_10160,N_9898,N_9670);
xor U10161 (N_10161,N_9700,N_9569);
xor U10162 (N_10162,N_9899,N_9535);
xor U10163 (N_10163,N_9713,N_9815);
and U10164 (N_10164,N_9931,N_9868);
xnor U10165 (N_10165,N_9555,N_9935);
xor U10166 (N_10166,N_9512,N_9879);
nand U10167 (N_10167,N_9591,N_9819);
or U10168 (N_10168,N_9977,N_9705);
or U10169 (N_10169,N_9802,N_9564);
and U10170 (N_10170,N_9687,N_9968);
nor U10171 (N_10171,N_9556,N_9729);
and U10172 (N_10172,N_9571,N_9818);
and U10173 (N_10173,N_9777,N_9601);
xnor U10174 (N_10174,N_9966,N_9773);
nor U10175 (N_10175,N_9730,N_9891);
xor U10176 (N_10176,N_9804,N_9588);
or U10177 (N_10177,N_9715,N_9716);
xnor U10178 (N_10178,N_9838,N_9654);
or U10179 (N_10179,N_9628,N_9967);
or U10180 (N_10180,N_9531,N_9592);
nor U10181 (N_10181,N_9664,N_9779);
nor U10182 (N_10182,N_9630,N_9661);
nor U10183 (N_10183,N_9560,N_9752);
nand U10184 (N_10184,N_9529,N_9634);
nand U10185 (N_10185,N_9861,N_9674);
nand U10186 (N_10186,N_9658,N_9542);
xnor U10187 (N_10187,N_9841,N_9832);
or U10188 (N_10188,N_9594,N_9965);
nor U10189 (N_10189,N_9955,N_9806);
nor U10190 (N_10190,N_9680,N_9655);
or U10191 (N_10191,N_9784,N_9643);
and U10192 (N_10192,N_9760,N_9645);
xnor U10193 (N_10193,N_9937,N_9558);
and U10194 (N_10194,N_9734,N_9736);
nand U10195 (N_10195,N_9860,N_9656);
xor U10196 (N_10196,N_9768,N_9998);
or U10197 (N_10197,N_9517,N_9506);
nand U10198 (N_10198,N_9827,N_9903);
or U10199 (N_10199,N_9718,N_9772);
nor U10200 (N_10200,N_9605,N_9820);
xnor U10201 (N_10201,N_9890,N_9607);
and U10202 (N_10202,N_9696,N_9738);
xor U10203 (N_10203,N_9812,N_9689);
and U10204 (N_10204,N_9551,N_9688);
xnor U10205 (N_10205,N_9906,N_9635);
xnor U10206 (N_10206,N_9771,N_9840);
nor U10207 (N_10207,N_9530,N_9684);
and U10208 (N_10208,N_9858,N_9702);
and U10209 (N_10209,N_9600,N_9770);
xnor U10210 (N_10210,N_9599,N_9557);
nor U10211 (N_10211,N_9976,N_9685);
xnor U10212 (N_10212,N_9789,N_9638);
xor U10213 (N_10213,N_9741,N_9547);
and U10214 (N_10214,N_9847,N_9724);
or U10215 (N_10215,N_9830,N_9810);
xnor U10216 (N_10216,N_9527,N_9665);
and U10217 (N_10217,N_9623,N_9550);
nor U10218 (N_10218,N_9678,N_9905);
or U10219 (N_10219,N_9743,N_9865);
and U10220 (N_10220,N_9545,N_9849);
or U10221 (N_10221,N_9781,N_9549);
or U10222 (N_10222,N_9790,N_9657);
nor U10223 (N_10223,N_9933,N_9833);
nor U10224 (N_10224,N_9597,N_9871);
xnor U10225 (N_10225,N_9948,N_9624);
nor U10226 (N_10226,N_9759,N_9980);
or U10227 (N_10227,N_9786,N_9754);
nand U10228 (N_10228,N_9572,N_9536);
xnor U10229 (N_10229,N_9563,N_9683);
or U10230 (N_10230,N_9504,N_9992);
or U10231 (N_10231,N_9867,N_9669);
nand U10232 (N_10232,N_9755,N_9846);
nand U10233 (N_10233,N_9875,N_9544);
and U10234 (N_10234,N_9745,N_9707);
or U10235 (N_10235,N_9961,N_9888);
or U10236 (N_10236,N_9582,N_9618);
or U10237 (N_10237,N_9566,N_9710);
and U10238 (N_10238,N_9603,N_9717);
or U10239 (N_10239,N_9763,N_9546);
nand U10240 (N_10240,N_9639,N_9769);
xnor U10241 (N_10241,N_9852,N_9698);
xor U10242 (N_10242,N_9914,N_9579);
nor U10243 (N_10243,N_9844,N_9649);
nand U10244 (N_10244,N_9788,N_9916);
and U10245 (N_10245,N_9570,N_9975);
xor U10246 (N_10246,N_9824,N_9712);
nor U10247 (N_10247,N_9581,N_9795);
and U10248 (N_10248,N_9963,N_9758);
nand U10249 (N_10249,N_9615,N_9596);
or U10250 (N_10250,N_9901,N_9612);
nand U10251 (N_10251,N_9923,N_9690);
nand U10252 (N_10252,N_9765,N_9665);
and U10253 (N_10253,N_9597,N_9762);
nor U10254 (N_10254,N_9802,N_9600);
or U10255 (N_10255,N_9676,N_9729);
nand U10256 (N_10256,N_9658,N_9645);
or U10257 (N_10257,N_9930,N_9939);
nand U10258 (N_10258,N_9599,N_9868);
nor U10259 (N_10259,N_9524,N_9760);
xnor U10260 (N_10260,N_9854,N_9915);
xor U10261 (N_10261,N_9926,N_9817);
nor U10262 (N_10262,N_9940,N_9525);
xnor U10263 (N_10263,N_9780,N_9969);
nor U10264 (N_10264,N_9827,N_9590);
xor U10265 (N_10265,N_9969,N_9632);
xor U10266 (N_10266,N_9735,N_9897);
nor U10267 (N_10267,N_9968,N_9664);
nand U10268 (N_10268,N_9585,N_9629);
xor U10269 (N_10269,N_9753,N_9505);
or U10270 (N_10270,N_9954,N_9773);
or U10271 (N_10271,N_9627,N_9618);
or U10272 (N_10272,N_9957,N_9507);
nand U10273 (N_10273,N_9525,N_9882);
nand U10274 (N_10274,N_9689,N_9904);
nor U10275 (N_10275,N_9503,N_9789);
nor U10276 (N_10276,N_9808,N_9576);
nand U10277 (N_10277,N_9900,N_9524);
nor U10278 (N_10278,N_9583,N_9561);
nor U10279 (N_10279,N_9872,N_9538);
xnor U10280 (N_10280,N_9625,N_9563);
xnor U10281 (N_10281,N_9656,N_9748);
nand U10282 (N_10282,N_9862,N_9516);
and U10283 (N_10283,N_9568,N_9853);
nor U10284 (N_10284,N_9724,N_9969);
nand U10285 (N_10285,N_9638,N_9697);
nand U10286 (N_10286,N_9890,N_9915);
nand U10287 (N_10287,N_9959,N_9851);
and U10288 (N_10288,N_9623,N_9665);
xnor U10289 (N_10289,N_9876,N_9973);
or U10290 (N_10290,N_9959,N_9900);
or U10291 (N_10291,N_9812,N_9825);
xor U10292 (N_10292,N_9585,N_9892);
xor U10293 (N_10293,N_9802,N_9882);
or U10294 (N_10294,N_9772,N_9738);
and U10295 (N_10295,N_9961,N_9799);
nand U10296 (N_10296,N_9634,N_9929);
xor U10297 (N_10297,N_9932,N_9747);
xnor U10298 (N_10298,N_9630,N_9834);
nand U10299 (N_10299,N_9917,N_9977);
or U10300 (N_10300,N_9593,N_9772);
or U10301 (N_10301,N_9810,N_9541);
nor U10302 (N_10302,N_9656,N_9561);
or U10303 (N_10303,N_9581,N_9882);
xnor U10304 (N_10304,N_9750,N_9737);
xnor U10305 (N_10305,N_9602,N_9896);
nand U10306 (N_10306,N_9565,N_9576);
xnor U10307 (N_10307,N_9718,N_9965);
and U10308 (N_10308,N_9984,N_9874);
nor U10309 (N_10309,N_9650,N_9910);
or U10310 (N_10310,N_9677,N_9879);
nand U10311 (N_10311,N_9871,N_9700);
xnor U10312 (N_10312,N_9903,N_9768);
nor U10313 (N_10313,N_9978,N_9620);
xor U10314 (N_10314,N_9947,N_9815);
and U10315 (N_10315,N_9731,N_9860);
nand U10316 (N_10316,N_9594,N_9536);
or U10317 (N_10317,N_9666,N_9517);
and U10318 (N_10318,N_9528,N_9627);
and U10319 (N_10319,N_9566,N_9639);
and U10320 (N_10320,N_9567,N_9763);
xor U10321 (N_10321,N_9757,N_9993);
and U10322 (N_10322,N_9710,N_9999);
or U10323 (N_10323,N_9577,N_9743);
or U10324 (N_10324,N_9739,N_9789);
and U10325 (N_10325,N_9907,N_9597);
nor U10326 (N_10326,N_9717,N_9811);
nor U10327 (N_10327,N_9929,N_9637);
nand U10328 (N_10328,N_9552,N_9762);
nor U10329 (N_10329,N_9547,N_9787);
or U10330 (N_10330,N_9845,N_9822);
xnor U10331 (N_10331,N_9702,N_9756);
xnor U10332 (N_10332,N_9897,N_9586);
nor U10333 (N_10333,N_9844,N_9875);
nor U10334 (N_10334,N_9910,N_9955);
xnor U10335 (N_10335,N_9679,N_9891);
xor U10336 (N_10336,N_9985,N_9842);
nand U10337 (N_10337,N_9999,N_9844);
xnor U10338 (N_10338,N_9627,N_9776);
and U10339 (N_10339,N_9884,N_9734);
or U10340 (N_10340,N_9851,N_9758);
nor U10341 (N_10341,N_9649,N_9633);
and U10342 (N_10342,N_9827,N_9779);
xor U10343 (N_10343,N_9975,N_9838);
nand U10344 (N_10344,N_9789,N_9776);
nand U10345 (N_10345,N_9818,N_9966);
xnor U10346 (N_10346,N_9646,N_9529);
xnor U10347 (N_10347,N_9570,N_9808);
xnor U10348 (N_10348,N_9948,N_9529);
or U10349 (N_10349,N_9583,N_9639);
nor U10350 (N_10350,N_9851,N_9733);
and U10351 (N_10351,N_9778,N_9536);
or U10352 (N_10352,N_9808,N_9560);
nand U10353 (N_10353,N_9998,N_9959);
xnor U10354 (N_10354,N_9922,N_9763);
xor U10355 (N_10355,N_9880,N_9691);
and U10356 (N_10356,N_9688,N_9622);
xor U10357 (N_10357,N_9991,N_9723);
and U10358 (N_10358,N_9731,N_9912);
nand U10359 (N_10359,N_9898,N_9963);
or U10360 (N_10360,N_9835,N_9785);
and U10361 (N_10361,N_9658,N_9844);
nor U10362 (N_10362,N_9858,N_9861);
and U10363 (N_10363,N_9938,N_9960);
xnor U10364 (N_10364,N_9895,N_9637);
or U10365 (N_10365,N_9825,N_9631);
nor U10366 (N_10366,N_9707,N_9850);
nand U10367 (N_10367,N_9560,N_9582);
nand U10368 (N_10368,N_9979,N_9705);
xnor U10369 (N_10369,N_9882,N_9915);
nor U10370 (N_10370,N_9998,N_9824);
nor U10371 (N_10371,N_9902,N_9677);
and U10372 (N_10372,N_9588,N_9910);
or U10373 (N_10373,N_9812,N_9682);
and U10374 (N_10374,N_9788,N_9525);
nor U10375 (N_10375,N_9648,N_9614);
nand U10376 (N_10376,N_9558,N_9882);
nand U10377 (N_10377,N_9612,N_9533);
and U10378 (N_10378,N_9646,N_9649);
nand U10379 (N_10379,N_9572,N_9694);
or U10380 (N_10380,N_9546,N_9797);
and U10381 (N_10381,N_9801,N_9930);
nand U10382 (N_10382,N_9993,N_9833);
or U10383 (N_10383,N_9602,N_9858);
nor U10384 (N_10384,N_9597,N_9751);
nor U10385 (N_10385,N_9835,N_9968);
nor U10386 (N_10386,N_9580,N_9923);
xnor U10387 (N_10387,N_9825,N_9871);
xnor U10388 (N_10388,N_9663,N_9930);
nand U10389 (N_10389,N_9863,N_9703);
nor U10390 (N_10390,N_9861,N_9902);
or U10391 (N_10391,N_9713,N_9832);
nor U10392 (N_10392,N_9994,N_9694);
nor U10393 (N_10393,N_9727,N_9827);
or U10394 (N_10394,N_9772,N_9904);
nand U10395 (N_10395,N_9601,N_9804);
and U10396 (N_10396,N_9541,N_9586);
nand U10397 (N_10397,N_9527,N_9713);
and U10398 (N_10398,N_9712,N_9783);
xor U10399 (N_10399,N_9595,N_9738);
xor U10400 (N_10400,N_9515,N_9726);
xor U10401 (N_10401,N_9934,N_9518);
xor U10402 (N_10402,N_9561,N_9882);
xor U10403 (N_10403,N_9520,N_9879);
or U10404 (N_10404,N_9761,N_9548);
nand U10405 (N_10405,N_9741,N_9577);
and U10406 (N_10406,N_9837,N_9955);
nand U10407 (N_10407,N_9872,N_9575);
and U10408 (N_10408,N_9970,N_9878);
nor U10409 (N_10409,N_9645,N_9753);
and U10410 (N_10410,N_9906,N_9860);
and U10411 (N_10411,N_9667,N_9966);
and U10412 (N_10412,N_9771,N_9942);
xor U10413 (N_10413,N_9779,N_9751);
nand U10414 (N_10414,N_9809,N_9914);
nor U10415 (N_10415,N_9954,N_9843);
nor U10416 (N_10416,N_9952,N_9753);
nor U10417 (N_10417,N_9853,N_9813);
nand U10418 (N_10418,N_9604,N_9643);
and U10419 (N_10419,N_9793,N_9782);
and U10420 (N_10420,N_9655,N_9889);
and U10421 (N_10421,N_9663,N_9940);
nor U10422 (N_10422,N_9536,N_9755);
xnor U10423 (N_10423,N_9863,N_9900);
or U10424 (N_10424,N_9943,N_9743);
xnor U10425 (N_10425,N_9557,N_9500);
xnor U10426 (N_10426,N_9760,N_9620);
nand U10427 (N_10427,N_9745,N_9838);
xor U10428 (N_10428,N_9882,N_9956);
and U10429 (N_10429,N_9802,N_9941);
nor U10430 (N_10430,N_9630,N_9704);
and U10431 (N_10431,N_9519,N_9573);
nor U10432 (N_10432,N_9541,N_9542);
or U10433 (N_10433,N_9860,N_9999);
or U10434 (N_10434,N_9892,N_9600);
nor U10435 (N_10435,N_9916,N_9548);
nor U10436 (N_10436,N_9665,N_9831);
or U10437 (N_10437,N_9572,N_9844);
nor U10438 (N_10438,N_9601,N_9504);
and U10439 (N_10439,N_9822,N_9930);
nor U10440 (N_10440,N_9617,N_9880);
nor U10441 (N_10441,N_9678,N_9692);
nor U10442 (N_10442,N_9760,N_9968);
and U10443 (N_10443,N_9971,N_9716);
or U10444 (N_10444,N_9737,N_9568);
nand U10445 (N_10445,N_9963,N_9685);
and U10446 (N_10446,N_9918,N_9954);
and U10447 (N_10447,N_9960,N_9696);
or U10448 (N_10448,N_9745,N_9725);
nand U10449 (N_10449,N_9921,N_9812);
and U10450 (N_10450,N_9602,N_9642);
or U10451 (N_10451,N_9662,N_9737);
xor U10452 (N_10452,N_9669,N_9887);
nor U10453 (N_10453,N_9670,N_9780);
nor U10454 (N_10454,N_9819,N_9736);
xnor U10455 (N_10455,N_9626,N_9974);
nor U10456 (N_10456,N_9767,N_9752);
nor U10457 (N_10457,N_9936,N_9591);
or U10458 (N_10458,N_9801,N_9595);
or U10459 (N_10459,N_9573,N_9900);
and U10460 (N_10460,N_9812,N_9865);
xnor U10461 (N_10461,N_9527,N_9915);
xor U10462 (N_10462,N_9526,N_9580);
xnor U10463 (N_10463,N_9521,N_9531);
xnor U10464 (N_10464,N_9942,N_9948);
or U10465 (N_10465,N_9890,N_9522);
or U10466 (N_10466,N_9603,N_9797);
and U10467 (N_10467,N_9566,N_9625);
or U10468 (N_10468,N_9920,N_9892);
nor U10469 (N_10469,N_9948,N_9664);
nand U10470 (N_10470,N_9572,N_9745);
and U10471 (N_10471,N_9764,N_9744);
nor U10472 (N_10472,N_9865,N_9883);
and U10473 (N_10473,N_9669,N_9853);
xnor U10474 (N_10474,N_9989,N_9715);
or U10475 (N_10475,N_9535,N_9908);
nor U10476 (N_10476,N_9802,N_9957);
and U10477 (N_10477,N_9646,N_9792);
and U10478 (N_10478,N_9555,N_9602);
and U10479 (N_10479,N_9729,N_9872);
or U10480 (N_10480,N_9582,N_9519);
nor U10481 (N_10481,N_9736,N_9904);
or U10482 (N_10482,N_9505,N_9945);
nor U10483 (N_10483,N_9978,N_9690);
nand U10484 (N_10484,N_9881,N_9586);
nor U10485 (N_10485,N_9990,N_9677);
or U10486 (N_10486,N_9954,N_9889);
xor U10487 (N_10487,N_9550,N_9890);
xnor U10488 (N_10488,N_9611,N_9964);
nand U10489 (N_10489,N_9721,N_9566);
nor U10490 (N_10490,N_9750,N_9513);
nor U10491 (N_10491,N_9561,N_9793);
xor U10492 (N_10492,N_9783,N_9607);
nand U10493 (N_10493,N_9765,N_9546);
nor U10494 (N_10494,N_9876,N_9878);
or U10495 (N_10495,N_9700,N_9925);
nor U10496 (N_10496,N_9567,N_9571);
nor U10497 (N_10497,N_9570,N_9890);
nor U10498 (N_10498,N_9552,N_9554);
nor U10499 (N_10499,N_9835,N_9732);
nor U10500 (N_10500,N_10233,N_10187);
nand U10501 (N_10501,N_10353,N_10319);
xnor U10502 (N_10502,N_10495,N_10481);
and U10503 (N_10503,N_10114,N_10445);
or U10504 (N_10504,N_10119,N_10030);
or U10505 (N_10505,N_10039,N_10407);
nand U10506 (N_10506,N_10386,N_10357);
nor U10507 (N_10507,N_10128,N_10374);
or U10508 (N_10508,N_10431,N_10205);
nand U10509 (N_10509,N_10210,N_10022);
xnor U10510 (N_10510,N_10477,N_10290);
or U10511 (N_10511,N_10420,N_10292);
or U10512 (N_10512,N_10082,N_10235);
nor U10513 (N_10513,N_10466,N_10349);
or U10514 (N_10514,N_10435,N_10281);
xnor U10515 (N_10515,N_10105,N_10230);
nand U10516 (N_10516,N_10024,N_10013);
and U10517 (N_10517,N_10146,N_10427);
and U10518 (N_10518,N_10457,N_10264);
xnor U10519 (N_10519,N_10074,N_10212);
xnor U10520 (N_10520,N_10009,N_10297);
nor U10521 (N_10521,N_10275,N_10261);
and U10522 (N_10522,N_10348,N_10279);
nand U10523 (N_10523,N_10192,N_10117);
nand U10524 (N_10524,N_10143,N_10392);
or U10525 (N_10525,N_10458,N_10299);
and U10526 (N_10526,N_10142,N_10285);
or U10527 (N_10527,N_10454,N_10444);
nor U10528 (N_10528,N_10189,N_10172);
xnor U10529 (N_10529,N_10089,N_10002);
nor U10530 (N_10530,N_10294,N_10482);
nor U10531 (N_10531,N_10472,N_10451);
xnor U10532 (N_10532,N_10116,N_10377);
xnor U10533 (N_10533,N_10220,N_10317);
and U10534 (N_10534,N_10120,N_10470);
or U10535 (N_10535,N_10010,N_10177);
xor U10536 (N_10536,N_10461,N_10456);
or U10537 (N_10537,N_10182,N_10405);
or U10538 (N_10538,N_10314,N_10023);
or U10539 (N_10539,N_10248,N_10197);
and U10540 (N_10540,N_10090,N_10194);
xor U10541 (N_10541,N_10066,N_10442);
nor U10542 (N_10542,N_10065,N_10052);
nor U10543 (N_10543,N_10301,N_10060);
and U10544 (N_10544,N_10343,N_10276);
xnor U10545 (N_10545,N_10153,N_10163);
and U10546 (N_10546,N_10397,N_10487);
xor U10547 (N_10547,N_10211,N_10395);
or U10548 (N_10548,N_10329,N_10325);
and U10549 (N_10549,N_10174,N_10157);
xor U10550 (N_10550,N_10476,N_10139);
nor U10551 (N_10551,N_10446,N_10135);
xor U10552 (N_10552,N_10387,N_10480);
or U10553 (N_10553,N_10436,N_10028);
nand U10554 (N_10554,N_10040,N_10008);
or U10555 (N_10555,N_10308,N_10412);
and U10556 (N_10556,N_10067,N_10450);
nor U10557 (N_10557,N_10096,N_10352);
nand U10558 (N_10558,N_10364,N_10221);
and U10559 (N_10559,N_10134,N_10473);
nor U10560 (N_10560,N_10206,N_10313);
nand U10561 (N_10561,N_10391,N_10488);
nand U10562 (N_10562,N_10147,N_10034);
and U10563 (N_10563,N_10304,N_10263);
nand U10564 (N_10564,N_10136,N_10198);
and U10565 (N_10565,N_10416,N_10241);
and U10566 (N_10566,N_10245,N_10069);
xor U10567 (N_10567,N_10196,N_10402);
and U10568 (N_10568,N_10362,N_10145);
and U10569 (N_10569,N_10358,N_10204);
nor U10570 (N_10570,N_10254,N_10253);
and U10571 (N_10571,N_10166,N_10242);
or U10572 (N_10572,N_10132,N_10266);
nor U10573 (N_10573,N_10422,N_10277);
nand U10574 (N_10574,N_10026,N_10133);
nand U10575 (N_10575,N_10332,N_10497);
or U10576 (N_10576,N_10140,N_10019);
and U10577 (N_10577,N_10462,N_10164);
xnor U10578 (N_10578,N_10268,N_10443);
or U10579 (N_10579,N_10490,N_10366);
xor U10580 (N_10580,N_10186,N_10014);
xnor U10581 (N_10581,N_10403,N_10126);
nand U10582 (N_10582,N_10303,N_10033);
xor U10583 (N_10583,N_10491,N_10367);
and U10584 (N_10584,N_10121,N_10440);
and U10585 (N_10585,N_10141,N_10296);
or U10586 (N_10586,N_10016,N_10193);
nand U10587 (N_10587,N_10478,N_10380);
nand U10588 (N_10588,N_10447,N_10368);
and U10589 (N_10589,N_10410,N_10088);
and U10590 (N_10590,N_10494,N_10102);
or U10591 (N_10591,N_10234,N_10448);
nand U10592 (N_10592,N_10243,N_10224);
and U10593 (N_10593,N_10369,N_10291);
nand U10594 (N_10594,N_10201,N_10180);
xnor U10595 (N_10595,N_10280,N_10104);
nor U10596 (N_10596,N_10094,N_10113);
nor U10597 (N_10597,N_10295,N_10483);
xnor U10598 (N_10598,N_10350,N_10429);
nor U10599 (N_10599,N_10401,N_10095);
or U10600 (N_10600,N_10158,N_10041);
xor U10601 (N_10601,N_10001,N_10346);
or U10602 (N_10602,N_10337,N_10110);
nand U10603 (N_10603,N_10021,N_10236);
and U10604 (N_10604,N_10382,N_10273);
or U10605 (N_10605,N_10389,N_10216);
xnor U10606 (N_10606,N_10306,N_10324);
nor U10607 (N_10607,N_10379,N_10345);
xnor U10608 (N_10608,N_10097,N_10270);
nand U10609 (N_10609,N_10103,N_10231);
nor U10610 (N_10610,N_10137,N_10417);
nor U10611 (N_10611,N_10162,N_10284);
nand U10612 (N_10612,N_10171,N_10426);
nor U10613 (N_10613,N_10093,N_10398);
nand U10614 (N_10614,N_10287,N_10371);
xor U10615 (N_10615,N_10229,N_10131);
nor U10616 (N_10616,N_10181,N_10424);
nand U10617 (N_10617,N_10027,N_10312);
and U10618 (N_10618,N_10214,N_10365);
or U10619 (N_10619,N_10359,N_10286);
nand U10620 (N_10620,N_10053,N_10225);
or U10621 (N_10621,N_10251,N_10475);
and U10622 (N_10622,N_10489,N_10333);
and U10623 (N_10623,N_10161,N_10238);
and U10624 (N_10624,N_10390,N_10288);
xnor U10625 (N_10625,N_10000,N_10079);
nor U10626 (N_10626,N_10252,N_10381);
nor U10627 (N_10627,N_10434,N_10356);
xnor U10628 (N_10628,N_10237,N_10124);
xnor U10629 (N_10629,N_10344,N_10418);
and U10630 (N_10630,N_10107,N_10274);
nand U10631 (N_10631,N_10047,N_10059);
or U10632 (N_10632,N_10415,N_10311);
or U10633 (N_10633,N_10408,N_10072);
nor U10634 (N_10634,N_10265,N_10335);
nor U10635 (N_10635,N_10226,N_10112);
xor U10636 (N_10636,N_10309,N_10191);
or U10637 (N_10637,N_10188,N_10091);
or U10638 (N_10638,N_10115,N_10302);
and U10639 (N_10639,N_10108,N_10207);
nand U10640 (N_10640,N_10051,N_10259);
or U10641 (N_10641,N_10499,N_10320);
nor U10642 (N_10642,N_10098,N_10195);
nand U10643 (N_10643,N_10355,N_10298);
nand U10644 (N_10644,N_10106,N_10068);
nor U10645 (N_10645,N_10151,N_10441);
nand U10646 (N_10646,N_10378,N_10383);
xor U10647 (N_10647,N_10070,N_10471);
and U10648 (N_10648,N_10409,N_10075);
or U10649 (N_10649,N_10239,N_10167);
or U10650 (N_10650,N_10425,N_10496);
nor U10651 (N_10651,N_10086,N_10217);
or U10652 (N_10652,N_10432,N_10032);
nor U10653 (N_10653,N_10076,N_10087);
nor U10654 (N_10654,N_10246,N_10200);
nor U10655 (N_10655,N_10485,N_10006);
or U10656 (N_10656,N_10256,N_10042);
xnor U10657 (N_10657,N_10326,N_10449);
xor U10658 (N_10658,N_10479,N_10049);
xor U10659 (N_10659,N_10351,N_10017);
or U10660 (N_10660,N_10169,N_10249);
nand U10661 (N_10661,N_10227,N_10156);
xnor U10662 (N_10662,N_10213,N_10262);
nand U10663 (N_10663,N_10144,N_10305);
or U10664 (N_10664,N_10050,N_10149);
nor U10665 (N_10665,N_10465,N_10439);
nand U10666 (N_10666,N_10036,N_10111);
and U10667 (N_10667,N_10438,N_10168);
xor U10668 (N_10668,N_10370,N_10150);
xnor U10669 (N_10669,N_10278,N_10469);
xor U10670 (N_10670,N_10179,N_10414);
nor U10671 (N_10671,N_10208,N_10199);
nor U10672 (N_10672,N_10048,N_10393);
or U10673 (N_10673,N_10083,N_10338);
nand U10674 (N_10674,N_10437,N_10073);
nand U10675 (N_10675,N_10260,N_10428);
nand U10676 (N_10676,N_10406,N_10100);
or U10677 (N_10677,N_10218,N_10170);
and U10678 (N_10678,N_10129,N_10413);
nand U10679 (N_10679,N_10453,N_10421);
and U10680 (N_10680,N_10190,N_10498);
or U10681 (N_10681,N_10130,N_10184);
xor U10682 (N_10682,N_10400,N_10258);
xor U10683 (N_10683,N_10148,N_10209);
or U10684 (N_10684,N_10044,N_10080);
and U10685 (N_10685,N_10004,N_10321);
and U10686 (N_10686,N_10484,N_10399);
nor U10687 (N_10687,N_10354,N_10084);
and U10688 (N_10688,N_10007,N_10334);
or U10689 (N_10689,N_10492,N_10430);
xor U10690 (N_10690,N_10029,N_10467);
or U10691 (N_10691,N_10077,N_10394);
nor U10692 (N_10692,N_10085,N_10215);
nand U10693 (N_10693,N_10247,N_10257);
or U10694 (N_10694,N_10056,N_10185);
xor U10695 (N_10695,N_10455,N_10474);
nand U10696 (N_10696,N_10122,N_10384);
nor U10697 (N_10697,N_10336,N_10043);
nand U10698 (N_10698,N_10372,N_10283);
nand U10699 (N_10699,N_10081,N_10183);
nor U10700 (N_10700,N_10018,N_10109);
and U10701 (N_10701,N_10267,N_10493);
xor U10702 (N_10702,N_10176,N_10232);
nor U10703 (N_10703,N_10244,N_10045);
nor U10704 (N_10704,N_10310,N_10057);
and U10705 (N_10705,N_10092,N_10063);
nor U10706 (N_10706,N_10101,N_10361);
nor U10707 (N_10707,N_10300,N_10005);
and U10708 (N_10708,N_10316,N_10322);
nand U10709 (N_10709,N_10376,N_10071);
and U10710 (N_10710,N_10396,N_10078);
xor U10711 (N_10711,N_10038,N_10315);
nand U10712 (N_10712,N_10339,N_10375);
xnor U10713 (N_10713,N_10347,N_10015);
and U10714 (N_10714,N_10293,N_10486);
and U10715 (N_10715,N_10419,N_10271);
xnor U10716 (N_10716,N_10323,N_10464);
nand U10717 (N_10717,N_10055,N_10160);
or U10718 (N_10718,N_10012,N_10341);
and U10719 (N_10719,N_10037,N_10099);
nor U10720 (N_10720,N_10118,N_10219);
xnor U10721 (N_10721,N_10463,N_10318);
nor U10722 (N_10722,N_10031,N_10385);
xor U10723 (N_10723,N_10269,N_10020);
xor U10724 (N_10724,N_10155,N_10203);
nand U10725 (N_10725,N_10154,N_10223);
and U10726 (N_10726,N_10025,N_10046);
or U10727 (N_10727,N_10152,N_10388);
or U10728 (N_10728,N_10222,N_10178);
xor U10729 (N_10729,N_10255,N_10058);
xor U10730 (N_10730,N_10228,N_10202);
or U10731 (N_10731,N_10165,N_10307);
nor U10732 (N_10732,N_10327,N_10289);
nand U10733 (N_10733,N_10411,N_10064);
nand U10734 (N_10734,N_10282,N_10062);
nor U10735 (N_10735,N_10061,N_10360);
and U10736 (N_10736,N_10127,N_10125);
or U10737 (N_10737,N_10423,N_10468);
or U10738 (N_10738,N_10460,N_10250);
or U10739 (N_10739,N_10123,N_10272);
or U10740 (N_10740,N_10404,N_10373);
nor U10741 (N_10741,N_10054,N_10011);
and U10742 (N_10742,N_10240,N_10340);
and U10743 (N_10743,N_10331,N_10159);
and U10744 (N_10744,N_10035,N_10173);
nand U10745 (N_10745,N_10138,N_10175);
xor U10746 (N_10746,N_10433,N_10003);
or U10747 (N_10747,N_10363,N_10328);
xor U10748 (N_10748,N_10342,N_10330);
nor U10749 (N_10749,N_10459,N_10452);
nand U10750 (N_10750,N_10390,N_10353);
and U10751 (N_10751,N_10321,N_10392);
xnor U10752 (N_10752,N_10250,N_10097);
and U10753 (N_10753,N_10428,N_10294);
nor U10754 (N_10754,N_10131,N_10061);
xor U10755 (N_10755,N_10061,N_10202);
and U10756 (N_10756,N_10362,N_10481);
xnor U10757 (N_10757,N_10183,N_10023);
xor U10758 (N_10758,N_10024,N_10438);
and U10759 (N_10759,N_10048,N_10149);
or U10760 (N_10760,N_10168,N_10117);
nand U10761 (N_10761,N_10037,N_10169);
nor U10762 (N_10762,N_10012,N_10322);
xnor U10763 (N_10763,N_10309,N_10458);
and U10764 (N_10764,N_10353,N_10081);
nand U10765 (N_10765,N_10213,N_10119);
nor U10766 (N_10766,N_10397,N_10099);
xnor U10767 (N_10767,N_10021,N_10336);
nor U10768 (N_10768,N_10018,N_10289);
nand U10769 (N_10769,N_10436,N_10495);
and U10770 (N_10770,N_10341,N_10439);
nand U10771 (N_10771,N_10212,N_10243);
and U10772 (N_10772,N_10460,N_10434);
nor U10773 (N_10773,N_10445,N_10292);
or U10774 (N_10774,N_10409,N_10233);
or U10775 (N_10775,N_10296,N_10089);
and U10776 (N_10776,N_10331,N_10002);
and U10777 (N_10777,N_10239,N_10328);
nor U10778 (N_10778,N_10133,N_10038);
xor U10779 (N_10779,N_10456,N_10055);
or U10780 (N_10780,N_10128,N_10002);
or U10781 (N_10781,N_10169,N_10434);
nor U10782 (N_10782,N_10142,N_10173);
and U10783 (N_10783,N_10364,N_10409);
nor U10784 (N_10784,N_10215,N_10251);
nor U10785 (N_10785,N_10116,N_10143);
xor U10786 (N_10786,N_10292,N_10493);
and U10787 (N_10787,N_10062,N_10051);
or U10788 (N_10788,N_10237,N_10405);
nor U10789 (N_10789,N_10475,N_10413);
or U10790 (N_10790,N_10412,N_10330);
or U10791 (N_10791,N_10179,N_10119);
nor U10792 (N_10792,N_10066,N_10228);
nand U10793 (N_10793,N_10331,N_10470);
or U10794 (N_10794,N_10138,N_10020);
xor U10795 (N_10795,N_10139,N_10362);
nor U10796 (N_10796,N_10286,N_10096);
nand U10797 (N_10797,N_10277,N_10116);
or U10798 (N_10798,N_10278,N_10431);
xnor U10799 (N_10799,N_10221,N_10246);
nor U10800 (N_10800,N_10448,N_10421);
xnor U10801 (N_10801,N_10287,N_10466);
or U10802 (N_10802,N_10100,N_10094);
xor U10803 (N_10803,N_10162,N_10174);
nand U10804 (N_10804,N_10392,N_10461);
nand U10805 (N_10805,N_10431,N_10253);
xor U10806 (N_10806,N_10464,N_10059);
nand U10807 (N_10807,N_10170,N_10296);
xor U10808 (N_10808,N_10209,N_10230);
nand U10809 (N_10809,N_10318,N_10142);
xor U10810 (N_10810,N_10216,N_10122);
or U10811 (N_10811,N_10110,N_10129);
or U10812 (N_10812,N_10281,N_10009);
and U10813 (N_10813,N_10191,N_10455);
and U10814 (N_10814,N_10260,N_10107);
xor U10815 (N_10815,N_10184,N_10367);
xnor U10816 (N_10816,N_10228,N_10315);
and U10817 (N_10817,N_10282,N_10472);
and U10818 (N_10818,N_10246,N_10469);
and U10819 (N_10819,N_10093,N_10007);
xnor U10820 (N_10820,N_10344,N_10360);
and U10821 (N_10821,N_10227,N_10068);
nor U10822 (N_10822,N_10268,N_10052);
xor U10823 (N_10823,N_10483,N_10335);
or U10824 (N_10824,N_10336,N_10444);
xor U10825 (N_10825,N_10081,N_10094);
and U10826 (N_10826,N_10353,N_10418);
or U10827 (N_10827,N_10075,N_10079);
nor U10828 (N_10828,N_10111,N_10491);
or U10829 (N_10829,N_10496,N_10034);
xnor U10830 (N_10830,N_10436,N_10226);
xor U10831 (N_10831,N_10193,N_10397);
nor U10832 (N_10832,N_10353,N_10050);
xor U10833 (N_10833,N_10431,N_10372);
nor U10834 (N_10834,N_10325,N_10233);
nand U10835 (N_10835,N_10275,N_10042);
nand U10836 (N_10836,N_10236,N_10096);
xnor U10837 (N_10837,N_10124,N_10037);
nor U10838 (N_10838,N_10315,N_10345);
and U10839 (N_10839,N_10381,N_10191);
nand U10840 (N_10840,N_10126,N_10152);
nor U10841 (N_10841,N_10386,N_10079);
nand U10842 (N_10842,N_10431,N_10468);
nor U10843 (N_10843,N_10328,N_10211);
or U10844 (N_10844,N_10312,N_10285);
nand U10845 (N_10845,N_10418,N_10456);
nand U10846 (N_10846,N_10365,N_10382);
nor U10847 (N_10847,N_10069,N_10118);
and U10848 (N_10848,N_10407,N_10479);
and U10849 (N_10849,N_10269,N_10419);
nand U10850 (N_10850,N_10064,N_10121);
nor U10851 (N_10851,N_10323,N_10005);
xnor U10852 (N_10852,N_10286,N_10497);
xor U10853 (N_10853,N_10131,N_10480);
or U10854 (N_10854,N_10331,N_10284);
xor U10855 (N_10855,N_10288,N_10120);
nor U10856 (N_10856,N_10344,N_10306);
or U10857 (N_10857,N_10329,N_10187);
xor U10858 (N_10858,N_10446,N_10262);
and U10859 (N_10859,N_10242,N_10490);
and U10860 (N_10860,N_10490,N_10305);
xor U10861 (N_10861,N_10021,N_10481);
or U10862 (N_10862,N_10202,N_10309);
or U10863 (N_10863,N_10151,N_10491);
and U10864 (N_10864,N_10480,N_10401);
and U10865 (N_10865,N_10190,N_10395);
nand U10866 (N_10866,N_10226,N_10087);
xnor U10867 (N_10867,N_10433,N_10401);
nand U10868 (N_10868,N_10143,N_10424);
or U10869 (N_10869,N_10096,N_10269);
and U10870 (N_10870,N_10122,N_10203);
or U10871 (N_10871,N_10052,N_10407);
or U10872 (N_10872,N_10354,N_10037);
nor U10873 (N_10873,N_10402,N_10398);
xnor U10874 (N_10874,N_10098,N_10217);
and U10875 (N_10875,N_10473,N_10427);
nor U10876 (N_10876,N_10428,N_10110);
or U10877 (N_10877,N_10174,N_10249);
and U10878 (N_10878,N_10447,N_10323);
xor U10879 (N_10879,N_10272,N_10006);
nand U10880 (N_10880,N_10260,N_10443);
and U10881 (N_10881,N_10485,N_10488);
nand U10882 (N_10882,N_10048,N_10061);
and U10883 (N_10883,N_10301,N_10048);
nand U10884 (N_10884,N_10374,N_10454);
xor U10885 (N_10885,N_10277,N_10103);
or U10886 (N_10886,N_10019,N_10370);
nand U10887 (N_10887,N_10232,N_10250);
nand U10888 (N_10888,N_10364,N_10145);
or U10889 (N_10889,N_10476,N_10421);
nor U10890 (N_10890,N_10429,N_10198);
or U10891 (N_10891,N_10127,N_10038);
xnor U10892 (N_10892,N_10303,N_10485);
and U10893 (N_10893,N_10195,N_10161);
xnor U10894 (N_10894,N_10368,N_10378);
xnor U10895 (N_10895,N_10037,N_10417);
or U10896 (N_10896,N_10232,N_10403);
xnor U10897 (N_10897,N_10276,N_10370);
and U10898 (N_10898,N_10135,N_10444);
nor U10899 (N_10899,N_10480,N_10168);
and U10900 (N_10900,N_10112,N_10203);
xnor U10901 (N_10901,N_10310,N_10263);
or U10902 (N_10902,N_10372,N_10468);
xor U10903 (N_10903,N_10389,N_10306);
and U10904 (N_10904,N_10475,N_10483);
xnor U10905 (N_10905,N_10251,N_10039);
nand U10906 (N_10906,N_10200,N_10177);
and U10907 (N_10907,N_10389,N_10483);
and U10908 (N_10908,N_10309,N_10011);
or U10909 (N_10909,N_10127,N_10305);
nand U10910 (N_10910,N_10089,N_10170);
and U10911 (N_10911,N_10133,N_10282);
xor U10912 (N_10912,N_10146,N_10053);
nand U10913 (N_10913,N_10194,N_10351);
nand U10914 (N_10914,N_10328,N_10209);
and U10915 (N_10915,N_10161,N_10360);
nor U10916 (N_10916,N_10246,N_10078);
nand U10917 (N_10917,N_10319,N_10263);
or U10918 (N_10918,N_10098,N_10281);
or U10919 (N_10919,N_10473,N_10021);
or U10920 (N_10920,N_10388,N_10245);
and U10921 (N_10921,N_10348,N_10463);
or U10922 (N_10922,N_10177,N_10454);
xnor U10923 (N_10923,N_10142,N_10006);
and U10924 (N_10924,N_10454,N_10108);
xor U10925 (N_10925,N_10228,N_10420);
and U10926 (N_10926,N_10246,N_10412);
or U10927 (N_10927,N_10288,N_10256);
nand U10928 (N_10928,N_10363,N_10479);
xnor U10929 (N_10929,N_10386,N_10245);
nor U10930 (N_10930,N_10437,N_10478);
nand U10931 (N_10931,N_10155,N_10074);
nand U10932 (N_10932,N_10005,N_10496);
nand U10933 (N_10933,N_10153,N_10265);
xnor U10934 (N_10934,N_10340,N_10218);
or U10935 (N_10935,N_10072,N_10091);
or U10936 (N_10936,N_10062,N_10107);
nand U10937 (N_10937,N_10442,N_10477);
or U10938 (N_10938,N_10066,N_10467);
xnor U10939 (N_10939,N_10443,N_10447);
or U10940 (N_10940,N_10245,N_10425);
or U10941 (N_10941,N_10254,N_10323);
and U10942 (N_10942,N_10026,N_10207);
or U10943 (N_10943,N_10148,N_10260);
or U10944 (N_10944,N_10402,N_10232);
xnor U10945 (N_10945,N_10428,N_10227);
xnor U10946 (N_10946,N_10476,N_10372);
nand U10947 (N_10947,N_10302,N_10276);
or U10948 (N_10948,N_10421,N_10186);
and U10949 (N_10949,N_10256,N_10339);
or U10950 (N_10950,N_10310,N_10358);
and U10951 (N_10951,N_10346,N_10145);
nor U10952 (N_10952,N_10375,N_10370);
xnor U10953 (N_10953,N_10087,N_10208);
nor U10954 (N_10954,N_10445,N_10362);
nand U10955 (N_10955,N_10035,N_10433);
nor U10956 (N_10956,N_10022,N_10430);
or U10957 (N_10957,N_10036,N_10028);
or U10958 (N_10958,N_10030,N_10481);
and U10959 (N_10959,N_10110,N_10273);
nor U10960 (N_10960,N_10219,N_10019);
nor U10961 (N_10961,N_10459,N_10005);
and U10962 (N_10962,N_10393,N_10114);
xor U10963 (N_10963,N_10473,N_10415);
nand U10964 (N_10964,N_10062,N_10430);
nand U10965 (N_10965,N_10255,N_10061);
nor U10966 (N_10966,N_10263,N_10136);
and U10967 (N_10967,N_10017,N_10297);
nor U10968 (N_10968,N_10247,N_10044);
nor U10969 (N_10969,N_10396,N_10351);
or U10970 (N_10970,N_10016,N_10263);
nor U10971 (N_10971,N_10318,N_10096);
and U10972 (N_10972,N_10227,N_10210);
xnor U10973 (N_10973,N_10275,N_10399);
or U10974 (N_10974,N_10256,N_10143);
and U10975 (N_10975,N_10004,N_10178);
or U10976 (N_10976,N_10201,N_10061);
nand U10977 (N_10977,N_10155,N_10162);
and U10978 (N_10978,N_10162,N_10009);
nand U10979 (N_10979,N_10159,N_10007);
nand U10980 (N_10980,N_10473,N_10141);
xnor U10981 (N_10981,N_10013,N_10283);
xor U10982 (N_10982,N_10166,N_10391);
and U10983 (N_10983,N_10160,N_10104);
and U10984 (N_10984,N_10397,N_10209);
or U10985 (N_10985,N_10106,N_10475);
or U10986 (N_10986,N_10298,N_10085);
or U10987 (N_10987,N_10317,N_10168);
xnor U10988 (N_10988,N_10240,N_10135);
and U10989 (N_10989,N_10332,N_10133);
nor U10990 (N_10990,N_10064,N_10032);
nor U10991 (N_10991,N_10275,N_10153);
nand U10992 (N_10992,N_10464,N_10040);
or U10993 (N_10993,N_10454,N_10099);
and U10994 (N_10994,N_10468,N_10451);
nor U10995 (N_10995,N_10388,N_10355);
nor U10996 (N_10996,N_10384,N_10249);
xnor U10997 (N_10997,N_10384,N_10377);
nor U10998 (N_10998,N_10282,N_10166);
nand U10999 (N_10999,N_10293,N_10346);
or U11000 (N_11000,N_10674,N_10939);
or U11001 (N_11001,N_10745,N_10735);
or U11002 (N_11002,N_10598,N_10794);
or U11003 (N_11003,N_10841,N_10870);
and U11004 (N_11004,N_10512,N_10671);
xor U11005 (N_11005,N_10793,N_10836);
nand U11006 (N_11006,N_10617,N_10531);
and U11007 (N_11007,N_10907,N_10892);
nor U11008 (N_11008,N_10920,N_10867);
or U11009 (N_11009,N_10669,N_10663);
and U11010 (N_11010,N_10860,N_10707);
nor U11011 (N_11011,N_10904,N_10752);
xor U11012 (N_11012,N_10812,N_10866);
nand U11013 (N_11013,N_10642,N_10897);
or U11014 (N_11014,N_10937,N_10846);
nor U11015 (N_11015,N_10758,N_10514);
and U11016 (N_11016,N_10513,N_10574);
nand U11017 (N_11017,N_10965,N_10706);
and U11018 (N_11018,N_10730,N_10894);
and U11019 (N_11019,N_10543,N_10989);
or U11020 (N_11020,N_10868,N_10961);
xor U11021 (N_11021,N_10776,N_10627);
and U11022 (N_11022,N_10905,N_10565);
xor U11023 (N_11023,N_10676,N_10634);
nand U11024 (N_11024,N_10655,N_10819);
or U11025 (N_11025,N_10944,N_10893);
nand U11026 (N_11026,N_10670,N_10788);
xnor U11027 (N_11027,N_10619,N_10733);
and U11028 (N_11028,N_10615,N_10929);
xor U11029 (N_11029,N_10830,N_10908);
nand U11030 (N_11030,N_10532,N_10522);
xnor U11031 (N_11031,N_10861,N_10529);
and U11032 (N_11032,N_10770,N_10833);
nor U11033 (N_11033,N_10999,N_10964);
or U11034 (N_11034,N_10549,N_10504);
nor U11035 (N_11035,N_10986,N_10590);
nor U11036 (N_11036,N_10834,N_10697);
xnor U11037 (N_11037,N_10952,N_10507);
or U11038 (N_11038,N_10879,N_10912);
or U11039 (N_11039,N_10790,N_10963);
xor U11040 (N_11040,N_10643,N_10648);
xor U11041 (N_11041,N_10949,N_10946);
nand U11042 (N_11042,N_10806,N_10816);
or U11043 (N_11043,N_10505,N_10918);
and U11044 (N_11044,N_10661,N_10910);
xor U11045 (N_11045,N_10978,N_10973);
and U11046 (N_11046,N_10888,N_10673);
and U11047 (N_11047,N_10990,N_10659);
xnor U11048 (N_11048,N_10718,N_10589);
and U11049 (N_11049,N_10863,N_10838);
and U11050 (N_11050,N_10564,N_10985);
nor U11051 (N_11051,N_10562,N_10588);
nand U11052 (N_11052,N_10781,N_10962);
or U11053 (N_11053,N_10639,N_10716);
xor U11054 (N_11054,N_10799,N_10556);
and U11055 (N_11055,N_10678,N_10602);
and U11056 (N_11056,N_10778,N_10511);
nand U11057 (N_11057,N_10652,N_10773);
nand U11058 (N_11058,N_10853,N_10815);
and U11059 (N_11059,N_10829,N_10713);
nor U11060 (N_11060,N_10566,N_10597);
xor U11061 (N_11061,N_10624,N_10856);
and U11062 (N_11062,N_10525,N_10613);
nand U11063 (N_11063,N_10572,N_10850);
or U11064 (N_11064,N_10954,N_10967);
xnor U11065 (N_11065,N_10578,N_10821);
and U11066 (N_11066,N_10828,N_10546);
xnor U11067 (N_11067,N_10889,N_10560);
nor U11068 (N_11068,N_10945,N_10646);
or U11069 (N_11069,N_10500,N_10715);
xnor U11070 (N_11070,N_10516,N_10851);
nor U11071 (N_11071,N_10696,N_10877);
or U11072 (N_11072,N_10689,N_10708);
nand U11073 (N_11073,N_10785,N_10909);
and U11074 (N_11074,N_10738,N_10567);
xnor U11075 (N_11075,N_10903,N_10826);
or U11076 (N_11076,N_10784,N_10843);
nor U11077 (N_11077,N_10757,N_10871);
and U11078 (N_11078,N_10876,N_10822);
nor U11079 (N_11079,N_10916,N_10559);
xnor U11080 (N_11080,N_10621,N_10608);
nor U11081 (N_11081,N_10600,N_10641);
and U11082 (N_11082,N_10791,N_10988);
nor U11083 (N_11083,N_10530,N_10596);
and U11084 (N_11084,N_10987,N_10665);
xnor U11085 (N_11085,N_10824,N_10544);
xor U11086 (N_11086,N_10592,N_10796);
or U11087 (N_11087,N_10545,N_10637);
nor U11088 (N_11088,N_10569,N_10691);
nor U11089 (N_11089,N_10755,N_10996);
and U11090 (N_11090,N_10709,N_10979);
nor U11091 (N_11091,N_10900,N_10508);
nor U11092 (N_11092,N_10736,N_10571);
and U11093 (N_11093,N_10629,N_10557);
nand U11094 (N_11094,N_10845,N_10966);
and U11095 (N_11095,N_10664,N_10685);
nor U11096 (N_11096,N_10779,N_10524);
and U11097 (N_11097,N_10695,N_10506);
nand U11098 (N_11098,N_10789,N_10914);
nand U11099 (N_11099,N_10895,N_10743);
and U11100 (N_11100,N_10930,N_10595);
or U11101 (N_11101,N_10694,N_10885);
or U11102 (N_11102,N_10636,N_10977);
nor U11103 (N_11103,N_10787,N_10832);
and U11104 (N_11104,N_10727,N_10968);
nor U11105 (N_11105,N_10734,N_10741);
and U11106 (N_11106,N_10568,N_10911);
nand U11107 (N_11107,N_10917,N_10721);
xnor U11108 (N_11108,N_10679,N_10728);
and U11109 (N_11109,N_10555,N_10874);
nor U11110 (N_11110,N_10609,N_10640);
nand U11111 (N_11111,N_10958,N_10766);
nor U11112 (N_11112,N_10915,N_10724);
nand U11113 (N_11113,N_10971,N_10813);
nor U11114 (N_11114,N_10984,N_10872);
nor U11115 (N_11115,N_10782,N_10519);
nand U11116 (N_11116,N_10924,N_10969);
nand U11117 (N_11117,N_10881,N_10538);
or U11118 (N_11118,N_10825,N_10717);
or U11119 (N_11119,N_10869,N_10528);
or U11120 (N_11120,N_10951,N_10579);
and U11121 (N_11121,N_10680,N_10931);
xor U11122 (N_11122,N_10509,N_10774);
or U11123 (N_11123,N_10786,N_10587);
or U11124 (N_11124,N_10570,N_10804);
xor U11125 (N_11125,N_10623,N_10687);
nor U11126 (N_11126,N_10675,N_10681);
or U11127 (N_11127,N_10810,N_10855);
nor U11128 (N_11128,N_10862,N_10759);
nand U11129 (N_11129,N_10875,N_10701);
nor U11130 (N_11130,N_10501,N_10859);
nor U11131 (N_11131,N_10943,N_10818);
nand U11132 (N_11132,N_10692,N_10731);
or U11133 (N_11133,N_10959,N_10974);
or U11134 (N_11134,N_10960,N_10535);
or U11135 (N_11135,N_10995,N_10657);
xnor U11136 (N_11136,N_10729,N_10823);
nor U11137 (N_11137,N_10814,N_10552);
nand U11138 (N_11138,N_10576,N_10690);
or U11139 (N_11139,N_10645,N_10547);
nand U11140 (N_11140,N_10684,N_10541);
xor U11141 (N_11141,N_10998,N_10882);
xor U11142 (N_11142,N_10980,N_10527);
xor U11143 (N_11143,N_10994,N_10970);
nand U11144 (N_11144,N_10857,N_10662);
and U11145 (N_11145,N_10539,N_10797);
nor U11146 (N_11146,N_10777,N_10982);
nand U11147 (N_11147,N_10714,N_10884);
nor U11148 (N_11148,N_10686,N_10737);
and U11149 (N_11149,N_10933,N_10842);
nand U11150 (N_11150,N_10611,N_10616);
xor U11151 (N_11151,N_10762,N_10769);
nand U11152 (N_11152,N_10754,N_10775);
nand U11153 (N_11153,N_10612,N_10852);
nand U11154 (N_11154,N_10831,N_10873);
nor U11155 (N_11155,N_10534,N_10991);
nor U11156 (N_11156,N_10628,N_10936);
nand U11157 (N_11157,N_10957,N_10660);
xnor U11158 (N_11158,N_10972,N_10503);
nand U11159 (N_11159,N_10551,N_10803);
or U11160 (N_11160,N_10901,N_10618);
and U11161 (N_11161,N_10953,N_10837);
or U11162 (N_11162,N_10536,N_10765);
nor U11163 (N_11163,N_10521,N_10740);
nor U11164 (N_11164,N_10693,N_10800);
xnor U11165 (N_11165,N_10805,N_10599);
nor U11166 (N_11166,N_10750,N_10700);
nor U11167 (N_11167,N_10926,N_10677);
and U11168 (N_11168,N_10561,N_10807);
nor U11169 (N_11169,N_10553,N_10575);
xnor U11170 (N_11170,N_10607,N_10902);
nand U11171 (N_11171,N_10502,N_10703);
xor U11172 (N_11172,N_10667,N_10940);
and U11173 (N_11173,N_10658,N_10771);
nand U11174 (N_11174,N_10583,N_10802);
xor U11175 (N_11175,N_10906,N_10610);
nand U11176 (N_11176,N_10783,N_10809);
nand U11177 (N_11177,N_10848,N_10622);
nor U11178 (N_11178,N_10950,N_10558);
xor U11179 (N_11179,N_10649,N_10742);
nand U11180 (N_11180,N_10927,N_10880);
nor U11181 (N_11181,N_10883,N_10523);
xor U11182 (N_11182,N_10792,N_10919);
xor U11183 (N_11183,N_10651,N_10923);
xnor U11184 (N_11184,N_10760,N_10702);
or U11185 (N_11185,N_10582,N_10753);
nor U11186 (N_11186,N_10698,N_10554);
nand U11187 (N_11187,N_10795,N_10928);
nor U11188 (N_11188,N_10840,N_10533);
xor U11189 (N_11189,N_10748,N_10683);
and U11190 (N_11190,N_10722,N_10710);
or U11191 (N_11191,N_10767,N_10540);
nor U11192 (N_11192,N_10725,N_10938);
nor U11193 (N_11193,N_10934,N_10626);
xor U11194 (N_11194,N_10548,N_10886);
nand U11195 (N_11195,N_10520,N_10847);
xnor U11196 (N_11196,N_10510,N_10711);
and U11197 (N_11197,N_10625,N_10603);
xnor U11198 (N_11198,N_10956,N_10537);
and U11199 (N_11199,N_10633,N_10668);
and U11200 (N_11200,N_10763,N_10947);
nand U11201 (N_11201,N_10817,N_10890);
xnor U11202 (N_11202,N_10732,N_10981);
or U11203 (N_11203,N_10772,N_10808);
or U11204 (N_11204,N_10844,N_10811);
xor U11205 (N_11205,N_10638,N_10997);
and U11206 (N_11206,N_10756,N_10585);
nand U11207 (N_11207,N_10864,N_10712);
xor U11208 (N_11208,N_10898,N_10887);
xor U11209 (N_11209,N_10896,N_10594);
xor U11210 (N_11210,N_10672,N_10891);
and U11211 (N_11211,N_10839,N_10932);
xor U11212 (N_11212,N_10577,N_10726);
nand U11213 (N_11213,N_10542,N_10827);
or U11214 (N_11214,N_10518,N_10699);
xor U11215 (N_11215,N_10780,N_10768);
xor U11216 (N_11216,N_10976,N_10925);
nor U11217 (N_11217,N_10526,N_10644);
or U11218 (N_11218,N_10635,N_10584);
or U11219 (N_11219,N_10922,N_10632);
nand U11220 (N_11220,N_10992,N_10704);
and U11221 (N_11221,N_10746,N_10749);
or U11222 (N_11222,N_10614,N_10656);
nand U11223 (N_11223,N_10620,N_10764);
or U11224 (N_11224,N_10761,N_10515);
xnor U11225 (N_11225,N_10941,N_10688);
xnor U11226 (N_11226,N_10747,N_10604);
nor U11227 (N_11227,N_10650,N_10586);
nand U11228 (N_11228,N_10921,N_10942);
or U11229 (N_11229,N_10563,N_10647);
or U11230 (N_11230,N_10798,N_10719);
xnor U11231 (N_11231,N_10913,N_10751);
and U11232 (N_11232,N_10682,N_10593);
nor U11233 (N_11233,N_10975,N_10865);
and U11234 (N_11234,N_10605,N_10854);
xor U11235 (N_11235,N_10591,N_10580);
or U11236 (N_11236,N_10993,N_10601);
xor U11237 (N_11237,N_10573,N_10858);
nor U11238 (N_11238,N_10630,N_10948);
nand U11239 (N_11239,N_10899,N_10801);
and U11240 (N_11240,N_10935,N_10606);
or U11241 (N_11241,N_10849,N_10955);
nand U11242 (N_11242,N_10653,N_10835);
nor U11243 (N_11243,N_10878,N_10720);
and U11244 (N_11244,N_10723,N_10581);
xnor U11245 (N_11245,N_10820,N_10705);
or U11246 (N_11246,N_10666,N_10744);
and U11247 (N_11247,N_10517,N_10654);
or U11248 (N_11248,N_10983,N_10631);
or U11249 (N_11249,N_10739,N_10550);
and U11250 (N_11250,N_10718,N_10969);
xnor U11251 (N_11251,N_10537,N_10738);
xnor U11252 (N_11252,N_10593,N_10543);
or U11253 (N_11253,N_10705,N_10823);
and U11254 (N_11254,N_10796,N_10854);
xnor U11255 (N_11255,N_10774,N_10896);
and U11256 (N_11256,N_10826,N_10560);
xnor U11257 (N_11257,N_10787,N_10684);
and U11258 (N_11258,N_10921,N_10699);
or U11259 (N_11259,N_10785,N_10662);
or U11260 (N_11260,N_10584,N_10692);
nor U11261 (N_11261,N_10659,N_10678);
nand U11262 (N_11262,N_10678,N_10794);
and U11263 (N_11263,N_10605,N_10996);
nand U11264 (N_11264,N_10603,N_10635);
or U11265 (N_11265,N_10798,N_10868);
or U11266 (N_11266,N_10716,N_10507);
and U11267 (N_11267,N_10622,N_10947);
and U11268 (N_11268,N_10832,N_10911);
nor U11269 (N_11269,N_10969,N_10704);
xnor U11270 (N_11270,N_10977,N_10502);
or U11271 (N_11271,N_10632,N_10608);
or U11272 (N_11272,N_10924,N_10910);
xnor U11273 (N_11273,N_10960,N_10612);
nand U11274 (N_11274,N_10689,N_10700);
and U11275 (N_11275,N_10716,N_10940);
nor U11276 (N_11276,N_10916,N_10843);
nand U11277 (N_11277,N_10556,N_10742);
xnor U11278 (N_11278,N_10546,N_10566);
nor U11279 (N_11279,N_10984,N_10745);
xnor U11280 (N_11280,N_10527,N_10682);
nor U11281 (N_11281,N_10882,N_10969);
and U11282 (N_11282,N_10987,N_10525);
nand U11283 (N_11283,N_10842,N_10967);
nor U11284 (N_11284,N_10727,N_10834);
nand U11285 (N_11285,N_10588,N_10504);
xnor U11286 (N_11286,N_10612,N_10636);
nand U11287 (N_11287,N_10577,N_10773);
or U11288 (N_11288,N_10779,N_10774);
nor U11289 (N_11289,N_10978,N_10627);
xor U11290 (N_11290,N_10925,N_10598);
and U11291 (N_11291,N_10792,N_10766);
nand U11292 (N_11292,N_10833,N_10633);
nor U11293 (N_11293,N_10543,N_10518);
nand U11294 (N_11294,N_10546,N_10940);
nand U11295 (N_11295,N_10647,N_10915);
xor U11296 (N_11296,N_10853,N_10974);
nor U11297 (N_11297,N_10557,N_10861);
and U11298 (N_11298,N_10510,N_10685);
or U11299 (N_11299,N_10704,N_10814);
and U11300 (N_11300,N_10890,N_10848);
or U11301 (N_11301,N_10890,N_10701);
xor U11302 (N_11302,N_10788,N_10577);
and U11303 (N_11303,N_10665,N_10781);
and U11304 (N_11304,N_10730,N_10791);
and U11305 (N_11305,N_10798,N_10510);
and U11306 (N_11306,N_10677,N_10930);
nor U11307 (N_11307,N_10872,N_10889);
xor U11308 (N_11308,N_10687,N_10829);
nand U11309 (N_11309,N_10890,N_10880);
or U11310 (N_11310,N_10534,N_10867);
nand U11311 (N_11311,N_10859,N_10797);
xor U11312 (N_11312,N_10514,N_10604);
and U11313 (N_11313,N_10725,N_10800);
xnor U11314 (N_11314,N_10975,N_10587);
and U11315 (N_11315,N_10912,N_10802);
nand U11316 (N_11316,N_10948,N_10624);
xnor U11317 (N_11317,N_10610,N_10973);
nor U11318 (N_11318,N_10756,N_10707);
and U11319 (N_11319,N_10668,N_10599);
nand U11320 (N_11320,N_10624,N_10521);
nand U11321 (N_11321,N_10962,N_10511);
or U11322 (N_11322,N_10572,N_10947);
and U11323 (N_11323,N_10921,N_10519);
xor U11324 (N_11324,N_10959,N_10737);
nor U11325 (N_11325,N_10946,N_10964);
nor U11326 (N_11326,N_10771,N_10540);
or U11327 (N_11327,N_10619,N_10721);
nor U11328 (N_11328,N_10799,N_10695);
nor U11329 (N_11329,N_10979,N_10590);
xnor U11330 (N_11330,N_10593,N_10634);
nand U11331 (N_11331,N_10703,N_10668);
or U11332 (N_11332,N_10594,N_10773);
nand U11333 (N_11333,N_10832,N_10986);
xnor U11334 (N_11334,N_10714,N_10899);
or U11335 (N_11335,N_10668,N_10827);
and U11336 (N_11336,N_10959,N_10940);
nor U11337 (N_11337,N_10610,N_10895);
nand U11338 (N_11338,N_10600,N_10666);
xor U11339 (N_11339,N_10851,N_10813);
nor U11340 (N_11340,N_10618,N_10816);
and U11341 (N_11341,N_10722,N_10697);
or U11342 (N_11342,N_10986,N_10699);
xnor U11343 (N_11343,N_10910,N_10995);
or U11344 (N_11344,N_10964,N_10640);
nand U11345 (N_11345,N_10835,N_10808);
nand U11346 (N_11346,N_10734,N_10874);
nand U11347 (N_11347,N_10664,N_10973);
or U11348 (N_11348,N_10708,N_10635);
nor U11349 (N_11349,N_10999,N_10980);
nand U11350 (N_11350,N_10682,N_10939);
nand U11351 (N_11351,N_10765,N_10782);
or U11352 (N_11352,N_10785,N_10800);
nand U11353 (N_11353,N_10504,N_10500);
and U11354 (N_11354,N_10911,N_10889);
or U11355 (N_11355,N_10575,N_10809);
nor U11356 (N_11356,N_10580,N_10688);
nor U11357 (N_11357,N_10854,N_10824);
nand U11358 (N_11358,N_10930,N_10648);
nand U11359 (N_11359,N_10627,N_10675);
nor U11360 (N_11360,N_10627,N_10573);
or U11361 (N_11361,N_10551,N_10936);
nor U11362 (N_11362,N_10992,N_10649);
xnor U11363 (N_11363,N_10935,N_10526);
nand U11364 (N_11364,N_10739,N_10648);
and U11365 (N_11365,N_10576,N_10636);
xnor U11366 (N_11366,N_10837,N_10795);
nand U11367 (N_11367,N_10973,N_10629);
nand U11368 (N_11368,N_10503,N_10903);
xor U11369 (N_11369,N_10698,N_10506);
xor U11370 (N_11370,N_10888,N_10999);
nand U11371 (N_11371,N_10793,N_10694);
nor U11372 (N_11372,N_10619,N_10562);
nor U11373 (N_11373,N_10561,N_10519);
nand U11374 (N_11374,N_10501,N_10692);
or U11375 (N_11375,N_10914,N_10533);
or U11376 (N_11376,N_10609,N_10780);
nand U11377 (N_11377,N_10993,N_10815);
and U11378 (N_11378,N_10511,N_10855);
nand U11379 (N_11379,N_10876,N_10879);
nand U11380 (N_11380,N_10720,N_10616);
nor U11381 (N_11381,N_10611,N_10555);
or U11382 (N_11382,N_10658,N_10542);
nor U11383 (N_11383,N_10892,N_10636);
xor U11384 (N_11384,N_10716,N_10926);
nand U11385 (N_11385,N_10649,N_10787);
nor U11386 (N_11386,N_10934,N_10878);
and U11387 (N_11387,N_10562,N_10932);
nand U11388 (N_11388,N_10844,N_10976);
nand U11389 (N_11389,N_10969,N_10782);
nand U11390 (N_11390,N_10637,N_10857);
nand U11391 (N_11391,N_10936,N_10910);
nand U11392 (N_11392,N_10590,N_10719);
and U11393 (N_11393,N_10845,N_10735);
and U11394 (N_11394,N_10956,N_10886);
or U11395 (N_11395,N_10951,N_10828);
and U11396 (N_11396,N_10717,N_10618);
xnor U11397 (N_11397,N_10509,N_10557);
or U11398 (N_11398,N_10763,N_10922);
or U11399 (N_11399,N_10562,N_10960);
and U11400 (N_11400,N_10507,N_10675);
or U11401 (N_11401,N_10946,N_10802);
nand U11402 (N_11402,N_10857,N_10773);
xor U11403 (N_11403,N_10847,N_10904);
nand U11404 (N_11404,N_10962,N_10994);
and U11405 (N_11405,N_10908,N_10618);
and U11406 (N_11406,N_10604,N_10600);
nand U11407 (N_11407,N_10667,N_10566);
nor U11408 (N_11408,N_10627,N_10662);
xnor U11409 (N_11409,N_10640,N_10925);
nor U11410 (N_11410,N_10858,N_10610);
or U11411 (N_11411,N_10954,N_10778);
or U11412 (N_11412,N_10974,N_10824);
and U11413 (N_11413,N_10743,N_10576);
nand U11414 (N_11414,N_10798,N_10708);
nand U11415 (N_11415,N_10615,N_10610);
nor U11416 (N_11416,N_10669,N_10565);
xor U11417 (N_11417,N_10720,N_10785);
or U11418 (N_11418,N_10930,N_10914);
xnor U11419 (N_11419,N_10539,N_10835);
and U11420 (N_11420,N_10797,N_10936);
nand U11421 (N_11421,N_10514,N_10575);
and U11422 (N_11422,N_10500,N_10883);
xnor U11423 (N_11423,N_10789,N_10932);
xor U11424 (N_11424,N_10777,N_10730);
nor U11425 (N_11425,N_10794,N_10926);
xnor U11426 (N_11426,N_10994,N_10990);
nor U11427 (N_11427,N_10916,N_10829);
and U11428 (N_11428,N_10910,N_10697);
nor U11429 (N_11429,N_10568,N_10998);
nand U11430 (N_11430,N_10972,N_10858);
and U11431 (N_11431,N_10944,N_10520);
nand U11432 (N_11432,N_10759,N_10604);
xor U11433 (N_11433,N_10553,N_10540);
and U11434 (N_11434,N_10843,N_10748);
and U11435 (N_11435,N_10863,N_10520);
nor U11436 (N_11436,N_10626,N_10949);
xnor U11437 (N_11437,N_10880,N_10739);
nand U11438 (N_11438,N_10878,N_10573);
nand U11439 (N_11439,N_10700,N_10935);
nor U11440 (N_11440,N_10746,N_10858);
nor U11441 (N_11441,N_10970,N_10706);
xor U11442 (N_11442,N_10619,N_10624);
and U11443 (N_11443,N_10647,N_10541);
nand U11444 (N_11444,N_10910,N_10774);
xnor U11445 (N_11445,N_10504,N_10887);
xor U11446 (N_11446,N_10942,N_10852);
nor U11447 (N_11447,N_10785,N_10742);
nor U11448 (N_11448,N_10676,N_10731);
or U11449 (N_11449,N_10985,N_10720);
nand U11450 (N_11450,N_10524,N_10879);
or U11451 (N_11451,N_10612,N_10787);
and U11452 (N_11452,N_10758,N_10924);
xor U11453 (N_11453,N_10882,N_10849);
or U11454 (N_11454,N_10875,N_10657);
nor U11455 (N_11455,N_10883,N_10514);
and U11456 (N_11456,N_10605,N_10545);
nand U11457 (N_11457,N_10842,N_10683);
or U11458 (N_11458,N_10908,N_10766);
and U11459 (N_11459,N_10799,N_10706);
xnor U11460 (N_11460,N_10783,N_10585);
xnor U11461 (N_11461,N_10814,N_10640);
nor U11462 (N_11462,N_10687,N_10819);
or U11463 (N_11463,N_10769,N_10574);
and U11464 (N_11464,N_10648,N_10757);
xnor U11465 (N_11465,N_10965,N_10733);
xnor U11466 (N_11466,N_10915,N_10928);
nand U11467 (N_11467,N_10658,N_10887);
xnor U11468 (N_11468,N_10736,N_10506);
nand U11469 (N_11469,N_10505,N_10617);
xnor U11470 (N_11470,N_10565,N_10955);
nor U11471 (N_11471,N_10572,N_10670);
nand U11472 (N_11472,N_10996,N_10515);
nor U11473 (N_11473,N_10740,N_10611);
nand U11474 (N_11474,N_10870,N_10932);
nor U11475 (N_11475,N_10997,N_10742);
nand U11476 (N_11476,N_10996,N_10844);
nand U11477 (N_11477,N_10723,N_10689);
nor U11478 (N_11478,N_10774,N_10920);
xnor U11479 (N_11479,N_10569,N_10767);
nand U11480 (N_11480,N_10501,N_10882);
nand U11481 (N_11481,N_10891,N_10508);
and U11482 (N_11482,N_10972,N_10676);
nor U11483 (N_11483,N_10639,N_10918);
nand U11484 (N_11484,N_10649,N_10542);
nor U11485 (N_11485,N_10640,N_10903);
or U11486 (N_11486,N_10938,N_10719);
nor U11487 (N_11487,N_10774,N_10787);
nor U11488 (N_11488,N_10966,N_10515);
nor U11489 (N_11489,N_10625,N_10812);
nor U11490 (N_11490,N_10998,N_10934);
nor U11491 (N_11491,N_10983,N_10946);
and U11492 (N_11492,N_10811,N_10704);
nor U11493 (N_11493,N_10727,N_10612);
xor U11494 (N_11494,N_10573,N_10896);
nand U11495 (N_11495,N_10524,N_10671);
or U11496 (N_11496,N_10723,N_10538);
and U11497 (N_11497,N_10964,N_10988);
and U11498 (N_11498,N_10674,N_10686);
xnor U11499 (N_11499,N_10544,N_10691);
xor U11500 (N_11500,N_11049,N_11028);
nor U11501 (N_11501,N_11042,N_11287);
or U11502 (N_11502,N_11003,N_11172);
or U11503 (N_11503,N_11366,N_11025);
xor U11504 (N_11504,N_11074,N_11324);
nor U11505 (N_11505,N_11082,N_11248);
nand U11506 (N_11506,N_11346,N_11200);
nand U11507 (N_11507,N_11290,N_11458);
nor U11508 (N_11508,N_11405,N_11212);
or U11509 (N_11509,N_11361,N_11024);
nor U11510 (N_11510,N_11055,N_11134);
nand U11511 (N_11511,N_11455,N_11104);
xor U11512 (N_11512,N_11221,N_11018);
and U11513 (N_11513,N_11281,N_11053);
nand U11514 (N_11514,N_11161,N_11297);
and U11515 (N_11515,N_11370,N_11137);
nand U11516 (N_11516,N_11466,N_11288);
or U11517 (N_11517,N_11157,N_11038);
and U11518 (N_11518,N_11249,N_11444);
nand U11519 (N_11519,N_11308,N_11130);
nor U11520 (N_11520,N_11193,N_11262);
nand U11521 (N_11521,N_11479,N_11220);
and U11522 (N_11522,N_11206,N_11277);
nor U11523 (N_11523,N_11012,N_11194);
and U11524 (N_11524,N_11350,N_11171);
and U11525 (N_11525,N_11177,N_11023);
and U11526 (N_11526,N_11340,N_11181);
nor U11527 (N_11527,N_11226,N_11027);
nor U11528 (N_11528,N_11139,N_11227);
nor U11529 (N_11529,N_11187,N_11138);
nand U11530 (N_11530,N_11075,N_11205);
and U11531 (N_11531,N_11261,N_11013);
and U11532 (N_11532,N_11273,N_11257);
nor U11533 (N_11533,N_11339,N_11077);
xor U11534 (N_11534,N_11440,N_11387);
xnor U11535 (N_11535,N_11174,N_11166);
nor U11536 (N_11536,N_11496,N_11404);
xnor U11537 (N_11537,N_11237,N_11017);
nand U11538 (N_11538,N_11449,N_11268);
xnor U11539 (N_11539,N_11219,N_11375);
and U11540 (N_11540,N_11125,N_11253);
nand U11541 (N_11541,N_11167,N_11423);
nor U11542 (N_11542,N_11208,N_11389);
nor U11543 (N_11543,N_11355,N_11446);
or U11544 (N_11544,N_11124,N_11251);
nand U11545 (N_11545,N_11086,N_11477);
nand U11546 (N_11546,N_11425,N_11141);
nor U11547 (N_11547,N_11434,N_11280);
or U11548 (N_11548,N_11397,N_11330);
nor U11549 (N_11549,N_11416,N_11048);
nor U11550 (N_11550,N_11010,N_11345);
nor U11551 (N_11551,N_11060,N_11349);
nand U11552 (N_11552,N_11437,N_11299);
nor U11553 (N_11553,N_11438,N_11307);
or U11554 (N_11554,N_11164,N_11409);
and U11555 (N_11555,N_11005,N_11312);
nor U11556 (N_11556,N_11088,N_11252);
and U11557 (N_11557,N_11402,N_11233);
and U11558 (N_11558,N_11406,N_11238);
or U11559 (N_11559,N_11395,N_11276);
nor U11560 (N_11560,N_11400,N_11169);
or U11561 (N_11561,N_11068,N_11431);
and U11562 (N_11562,N_11443,N_11274);
xnor U11563 (N_11563,N_11015,N_11188);
nand U11564 (N_11564,N_11179,N_11145);
nor U11565 (N_11565,N_11372,N_11032);
and U11566 (N_11566,N_11338,N_11424);
and U11567 (N_11567,N_11064,N_11236);
nand U11568 (N_11568,N_11489,N_11476);
or U11569 (N_11569,N_11398,N_11110);
or U11570 (N_11570,N_11492,N_11057);
and U11571 (N_11571,N_11310,N_11163);
or U11572 (N_11572,N_11359,N_11084);
or U11573 (N_11573,N_11054,N_11180);
xor U11574 (N_11574,N_11436,N_11411);
or U11575 (N_11575,N_11490,N_11391);
xnor U11576 (N_11576,N_11468,N_11302);
xor U11577 (N_11577,N_11083,N_11232);
nor U11578 (N_11578,N_11118,N_11070);
and U11579 (N_11579,N_11327,N_11315);
xor U11580 (N_11580,N_11356,N_11317);
xnor U11581 (N_11581,N_11294,N_11266);
nor U11582 (N_11582,N_11225,N_11422);
xnor U11583 (N_11583,N_11363,N_11323);
nor U11584 (N_11584,N_11195,N_11333);
or U11585 (N_11585,N_11360,N_11269);
nand U11586 (N_11586,N_11108,N_11420);
nand U11587 (N_11587,N_11207,N_11456);
nand U11588 (N_11588,N_11442,N_11170);
nand U11589 (N_11589,N_11494,N_11008);
nand U11590 (N_11590,N_11105,N_11335);
xnor U11591 (N_11591,N_11184,N_11063);
xnor U11592 (N_11592,N_11016,N_11415);
nand U11593 (N_11593,N_11499,N_11247);
nor U11594 (N_11594,N_11351,N_11279);
nor U11595 (N_11595,N_11199,N_11168);
and U11596 (N_11596,N_11058,N_11019);
or U11597 (N_11597,N_11050,N_11198);
nor U11598 (N_11598,N_11433,N_11250);
xnor U11599 (N_11599,N_11450,N_11107);
or U11600 (N_11600,N_11071,N_11471);
or U11601 (N_11601,N_11156,N_11090);
xnor U11602 (N_11602,N_11097,N_11254);
xnor U11603 (N_11603,N_11040,N_11031);
nor U11604 (N_11604,N_11214,N_11210);
xnor U11605 (N_11605,N_11116,N_11044);
and U11606 (N_11606,N_11377,N_11259);
xor U11607 (N_11607,N_11484,N_11240);
nand U11608 (N_11608,N_11011,N_11267);
or U11609 (N_11609,N_11135,N_11401);
nor U11610 (N_11610,N_11213,N_11491);
or U11611 (N_11611,N_11482,N_11224);
xor U11612 (N_11612,N_11403,N_11326);
nor U11613 (N_11613,N_11473,N_11337);
nand U11614 (N_11614,N_11129,N_11147);
xnor U11615 (N_11615,N_11033,N_11182);
and U11616 (N_11616,N_11155,N_11410);
nor U11617 (N_11617,N_11319,N_11460);
or U11618 (N_11618,N_11461,N_11306);
or U11619 (N_11619,N_11223,N_11244);
xor U11620 (N_11620,N_11474,N_11154);
or U11621 (N_11621,N_11119,N_11039);
and U11622 (N_11622,N_11114,N_11497);
nand U11623 (N_11623,N_11041,N_11093);
xnor U11624 (N_11624,N_11457,N_11029);
xnor U11625 (N_11625,N_11352,N_11092);
xnor U11626 (N_11626,N_11439,N_11464);
xnor U11627 (N_11627,N_11385,N_11286);
nand U11628 (N_11628,N_11272,N_11358);
or U11629 (N_11629,N_11045,N_11365);
xor U11630 (N_11630,N_11007,N_11102);
and U11631 (N_11631,N_11301,N_11022);
xnor U11632 (N_11632,N_11472,N_11295);
and U11633 (N_11633,N_11165,N_11435);
nand U11634 (N_11634,N_11133,N_11432);
nand U11635 (N_11635,N_11486,N_11467);
nand U11636 (N_11636,N_11378,N_11412);
or U11637 (N_11637,N_11413,N_11152);
xor U11638 (N_11638,N_11256,N_11140);
nor U11639 (N_11639,N_11127,N_11454);
xnor U11640 (N_11640,N_11201,N_11146);
and U11641 (N_11641,N_11357,N_11209);
xor U11642 (N_11642,N_11382,N_11414);
or U11643 (N_11643,N_11001,N_11160);
and U11644 (N_11644,N_11331,N_11481);
xnor U11645 (N_11645,N_11448,N_11344);
and U11646 (N_11646,N_11478,N_11056);
nor U11647 (N_11647,N_11289,N_11204);
and U11648 (N_11648,N_11293,N_11419);
and U11649 (N_11649,N_11383,N_11441);
xor U11650 (N_11650,N_11392,N_11278);
xnor U11651 (N_11651,N_11354,N_11120);
nor U11652 (N_11652,N_11242,N_11393);
and U11653 (N_11653,N_11325,N_11364);
xnor U11654 (N_11654,N_11483,N_11126);
nor U11655 (N_11655,N_11106,N_11296);
xor U11656 (N_11656,N_11316,N_11283);
and U11657 (N_11657,N_11085,N_11215);
and U11658 (N_11658,N_11390,N_11353);
and U11659 (N_11659,N_11173,N_11043);
nor U11660 (N_11660,N_11131,N_11035);
nor U11661 (N_11661,N_11059,N_11239);
or U11662 (N_11662,N_11004,N_11100);
and U11663 (N_11663,N_11298,N_11094);
nor U11664 (N_11664,N_11109,N_11030);
nand U11665 (N_11665,N_11493,N_11342);
or U11666 (N_11666,N_11121,N_11020);
nand U11667 (N_11667,N_11115,N_11142);
xnor U11668 (N_11668,N_11417,N_11380);
and U11669 (N_11669,N_11159,N_11367);
and U11670 (N_11670,N_11186,N_11381);
xor U11671 (N_11671,N_11037,N_11000);
and U11672 (N_11672,N_11190,N_11488);
nand U11673 (N_11673,N_11255,N_11388);
or U11674 (N_11674,N_11426,N_11246);
or U11675 (N_11675,N_11112,N_11178);
nor U11676 (N_11676,N_11459,N_11128);
nor U11677 (N_11677,N_11322,N_11036);
and U11678 (N_11678,N_11408,N_11101);
xor U11679 (N_11679,N_11051,N_11087);
xnor U11680 (N_11680,N_11061,N_11006);
nand U11681 (N_11681,N_11421,N_11203);
xor U11682 (N_11682,N_11429,N_11123);
and U11683 (N_11683,N_11463,N_11189);
nand U11684 (N_11684,N_11202,N_11111);
xor U11685 (N_11685,N_11122,N_11211);
or U11686 (N_11686,N_11304,N_11487);
nor U11687 (N_11687,N_11270,N_11470);
xor U11688 (N_11688,N_11191,N_11428);
xnor U11689 (N_11689,N_11445,N_11243);
nand U11690 (N_11690,N_11469,N_11291);
and U11691 (N_11691,N_11495,N_11065);
xnor U11692 (N_11692,N_11462,N_11176);
xnor U11693 (N_11693,N_11263,N_11148);
nor U11694 (N_11694,N_11103,N_11334);
or U11695 (N_11695,N_11062,N_11447);
nand U11696 (N_11696,N_11185,N_11218);
and U11697 (N_11697,N_11014,N_11300);
or U11698 (N_11698,N_11052,N_11228);
nor U11699 (N_11699,N_11480,N_11452);
nor U11700 (N_11700,N_11091,N_11197);
xnor U11701 (N_11701,N_11430,N_11321);
nor U11702 (N_11702,N_11332,N_11009);
xor U11703 (N_11703,N_11368,N_11284);
and U11704 (N_11704,N_11089,N_11396);
or U11705 (N_11705,N_11002,N_11231);
nor U11706 (N_11706,N_11230,N_11078);
xnor U11707 (N_11707,N_11079,N_11098);
xor U11708 (N_11708,N_11183,N_11136);
and U11709 (N_11709,N_11026,N_11394);
or U11710 (N_11710,N_11073,N_11271);
and U11711 (N_11711,N_11313,N_11258);
nor U11712 (N_11712,N_11379,N_11407);
and U11713 (N_11713,N_11080,N_11072);
xnor U11714 (N_11714,N_11373,N_11047);
nor U11715 (N_11715,N_11369,N_11453);
and U11716 (N_11716,N_11158,N_11384);
nor U11717 (N_11717,N_11196,N_11343);
or U11718 (N_11718,N_11260,N_11348);
xnor U11719 (N_11719,N_11475,N_11314);
nand U11720 (N_11720,N_11144,N_11099);
nor U11721 (N_11721,N_11418,N_11282);
nand U11722 (N_11722,N_11309,N_11153);
nor U11723 (N_11723,N_11285,N_11498);
xnor U11724 (N_11724,N_11217,N_11485);
or U11725 (N_11725,N_11374,N_11235);
nor U11726 (N_11726,N_11329,N_11150);
or U11727 (N_11727,N_11347,N_11341);
or U11728 (N_11728,N_11096,N_11021);
nor U11729 (N_11729,N_11465,N_11305);
nand U11730 (N_11730,N_11067,N_11371);
and U11731 (N_11731,N_11151,N_11241);
and U11732 (N_11732,N_11376,N_11303);
nor U11733 (N_11733,N_11292,N_11216);
nand U11734 (N_11734,N_11095,N_11275);
or U11735 (N_11735,N_11245,N_11175);
and U11736 (N_11736,N_11222,N_11399);
nor U11737 (N_11737,N_11264,N_11320);
xor U11738 (N_11738,N_11318,N_11149);
nor U11739 (N_11739,N_11081,N_11336);
xor U11740 (N_11740,N_11046,N_11132);
xor U11741 (N_11741,N_11311,N_11069);
nor U11742 (N_11742,N_11117,N_11066);
or U11743 (N_11743,N_11427,N_11386);
and U11744 (N_11744,N_11234,N_11362);
and U11745 (N_11745,N_11143,N_11451);
and U11746 (N_11746,N_11076,N_11113);
nor U11747 (N_11747,N_11328,N_11192);
and U11748 (N_11748,N_11265,N_11162);
nor U11749 (N_11749,N_11229,N_11034);
xor U11750 (N_11750,N_11491,N_11243);
nor U11751 (N_11751,N_11486,N_11372);
and U11752 (N_11752,N_11346,N_11293);
or U11753 (N_11753,N_11426,N_11305);
nor U11754 (N_11754,N_11272,N_11453);
nor U11755 (N_11755,N_11218,N_11289);
nand U11756 (N_11756,N_11279,N_11391);
and U11757 (N_11757,N_11063,N_11171);
nor U11758 (N_11758,N_11202,N_11049);
xor U11759 (N_11759,N_11144,N_11370);
nand U11760 (N_11760,N_11150,N_11465);
xor U11761 (N_11761,N_11146,N_11151);
nor U11762 (N_11762,N_11027,N_11434);
nor U11763 (N_11763,N_11367,N_11435);
or U11764 (N_11764,N_11295,N_11493);
and U11765 (N_11765,N_11473,N_11372);
nand U11766 (N_11766,N_11426,N_11373);
nor U11767 (N_11767,N_11243,N_11482);
or U11768 (N_11768,N_11125,N_11351);
and U11769 (N_11769,N_11487,N_11179);
xnor U11770 (N_11770,N_11099,N_11486);
nor U11771 (N_11771,N_11107,N_11289);
and U11772 (N_11772,N_11248,N_11142);
or U11773 (N_11773,N_11035,N_11350);
nand U11774 (N_11774,N_11177,N_11007);
nor U11775 (N_11775,N_11057,N_11391);
or U11776 (N_11776,N_11311,N_11385);
xnor U11777 (N_11777,N_11161,N_11206);
nand U11778 (N_11778,N_11029,N_11054);
and U11779 (N_11779,N_11026,N_11150);
nand U11780 (N_11780,N_11287,N_11435);
or U11781 (N_11781,N_11437,N_11034);
xor U11782 (N_11782,N_11386,N_11405);
nand U11783 (N_11783,N_11256,N_11492);
nor U11784 (N_11784,N_11036,N_11380);
nand U11785 (N_11785,N_11313,N_11357);
and U11786 (N_11786,N_11004,N_11441);
and U11787 (N_11787,N_11354,N_11316);
nor U11788 (N_11788,N_11230,N_11232);
nor U11789 (N_11789,N_11363,N_11167);
and U11790 (N_11790,N_11102,N_11487);
xnor U11791 (N_11791,N_11195,N_11237);
nor U11792 (N_11792,N_11240,N_11035);
nor U11793 (N_11793,N_11085,N_11471);
xor U11794 (N_11794,N_11260,N_11209);
xnor U11795 (N_11795,N_11201,N_11295);
or U11796 (N_11796,N_11165,N_11163);
xnor U11797 (N_11797,N_11028,N_11347);
nand U11798 (N_11798,N_11360,N_11284);
nor U11799 (N_11799,N_11172,N_11240);
and U11800 (N_11800,N_11241,N_11045);
nor U11801 (N_11801,N_11221,N_11043);
and U11802 (N_11802,N_11074,N_11370);
or U11803 (N_11803,N_11298,N_11338);
xnor U11804 (N_11804,N_11442,N_11450);
or U11805 (N_11805,N_11417,N_11489);
and U11806 (N_11806,N_11321,N_11294);
or U11807 (N_11807,N_11001,N_11173);
or U11808 (N_11808,N_11224,N_11197);
or U11809 (N_11809,N_11332,N_11296);
nor U11810 (N_11810,N_11271,N_11081);
nor U11811 (N_11811,N_11080,N_11298);
xor U11812 (N_11812,N_11254,N_11024);
xnor U11813 (N_11813,N_11086,N_11219);
or U11814 (N_11814,N_11464,N_11322);
and U11815 (N_11815,N_11133,N_11315);
nor U11816 (N_11816,N_11307,N_11064);
and U11817 (N_11817,N_11155,N_11371);
xnor U11818 (N_11818,N_11141,N_11068);
and U11819 (N_11819,N_11064,N_11123);
nand U11820 (N_11820,N_11354,N_11402);
xnor U11821 (N_11821,N_11141,N_11420);
or U11822 (N_11822,N_11190,N_11250);
nand U11823 (N_11823,N_11235,N_11176);
and U11824 (N_11824,N_11163,N_11120);
xor U11825 (N_11825,N_11277,N_11174);
nor U11826 (N_11826,N_11427,N_11371);
or U11827 (N_11827,N_11205,N_11011);
or U11828 (N_11828,N_11268,N_11053);
nor U11829 (N_11829,N_11101,N_11155);
and U11830 (N_11830,N_11245,N_11223);
or U11831 (N_11831,N_11350,N_11076);
or U11832 (N_11832,N_11389,N_11086);
xnor U11833 (N_11833,N_11475,N_11488);
nand U11834 (N_11834,N_11128,N_11243);
xor U11835 (N_11835,N_11300,N_11325);
nand U11836 (N_11836,N_11162,N_11213);
nand U11837 (N_11837,N_11171,N_11352);
nand U11838 (N_11838,N_11277,N_11032);
xnor U11839 (N_11839,N_11463,N_11131);
or U11840 (N_11840,N_11088,N_11267);
xnor U11841 (N_11841,N_11134,N_11159);
nor U11842 (N_11842,N_11285,N_11332);
nand U11843 (N_11843,N_11138,N_11137);
nand U11844 (N_11844,N_11185,N_11378);
and U11845 (N_11845,N_11489,N_11485);
nor U11846 (N_11846,N_11109,N_11406);
nor U11847 (N_11847,N_11024,N_11360);
nand U11848 (N_11848,N_11373,N_11072);
and U11849 (N_11849,N_11237,N_11299);
or U11850 (N_11850,N_11250,N_11460);
nand U11851 (N_11851,N_11159,N_11266);
and U11852 (N_11852,N_11086,N_11124);
and U11853 (N_11853,N_11102,N_11253);
or U11854 (N_11854,N_11136,N_11210);
nor U11855 (N_11855,N_11415,N_11178);
nor U11856 (N_11856,N_11033,N_11116);
and U11857 (N_11857,N_11098,N_11033);
and U11858 (N_11858,N_11415,N_11345);
xor U11859 (N_11859,N_11270,N_11479);
or U11860 (N_11860,N_11328,N_11434);
nor U11861 (N_11861,N_11027,N_11126);
or U11862 (N_11862,N_11014,N_11211);
nand U11863 (N_11863,N_11168,N_11433);
nor U11864 (N_11864,N_11080,N_11031);
xor U11865 (N_11865,N_11216,N_11079);
nand U11866 (N_11866,N_11041,N_11183);
nor U11867 (N_11867,N_11046,N_11375);
nor U11868 (N_11868,N_11291,N_11112);
or U11869 (N_11869,N_11476,N_11376);
or U11870 (N_11870,N_11073,N_11048);
nand U11871 (N_11871,N_11381,N_11492);
or U11872 (N_11872,N_11360,N_11185);
nor U11873 (N_11873,N_11458,N_11461);
and U11874 (N_11874,N_11388,N_11215);
nand U11875 (N_11875,N_11272,N_11196);
nor U11876 (N_11876,N_11490,N_11210);
or U11877 (N_11877,N_11002,N_11153);
nand U11878 (N_11878,N_11283,N_11460);
and U11879 (N_11879,N_11382,N_11422);
xnor U11880 (N_11880,N_11039,N_11010);
nand U11881 (N_11881,N_11344,N_11150);
and U11882 (N_11882,N_11006,N_11144);
xor U11883 (N_11883,N_11194,N_11407);
nand U11884 (N_11884,N_11335,N_11198);
nand U11885 (N_11885,N_11394,N_11411);
and U11886 (N_11886,N_11334,N_11486);
xor U11887 (N_11887,N_11003,N_11037);
xnor U11888 (N_11888,N_11476,N_11102);
nor U11889 (N_11889,N_11140,N_11077);
xor U11890 (N_11890,N_11235,N_11001);
and U11891 (N_11891,N_11265,N_11203);
nand U11892 (N_11892,N_11215,N_11164);
or U11893 (N_11893,N_11133,N_11146);
nor U11894 (N_11894,N_11130,N_11480);
nand U11895 (N_11895,N_11446,N_11458);
or U11896 (N_11896,N_11118,N_11288);
nand U11897 (N_11897,N_11471,N_11178);
and U11898 (N_11898,N_11143,N_11068);
or U11899 (N_11899,N_11269,N_11407);
xor U11900 (N_11900,N_11111,N_11041);
nor U11901 (N_11901,N_11208,N_11117);
xor U11902 (N_11902,N_11224,N_11153);
nor U11903 (N_11903,N_11253,N_11183);
or U11904 (N_11904,N_11290,N_11037);
xnor U11905 (N_11905,N_11400,N_11307);
nor U11906 (N_11906,N_11064,N_11327);
nand U11907 (N_11907,N_11158,N_11400);
or U11908 (N_11908,N_11309,N_11365);
or U11909 (N_11909,N_11106,N_11185);
nor U11910 (N_11910,N_11334,N_11499);
nor U11911 (N_11911,N_11321,N_11316);
and U11912 (N_11912,N_11009,N_11316);
and U11913 (N_11913,N_11247,N_11418);
and U11914 (N_11914,N_11310,N_11075);
nand U11915 (N_11915,N_11411,N_11316);
xor U11916 (N_11916,N_11065,N_11165);
nor U11917 (N_11917,N_11219,N_11015);
nor U11918 (N_11918,N_11165,N_11266);
nor U11919 (N_11919,N_11279,N_11194);
xnor U11920 (N_11920,N_11270,N_11188);
and U11921 (N_11921,N_11003,N_11475);
nor U11922 (N_11922,N_11072,N_11277);
or U11923 (N_11923,N_11017,N_11124);
nor U11924 (N_11924,N_11204,N_11055);
or U11925 (N_11925,N_11249,N_11109);
or U11926 (N_11926,N_11397,N_11030);
nor U11927 (N_11927,N_11235,N_11218);
and U11928 (N_11928,N_11497,N_11269);
and U11929 (N_11929,N_11172,N_11145);
nor U11930 (N_11930,N_11023,N_11211);
nor U11931 (N_11931,N_11010,N_11046);
xnor U11932 (N_11932,N_11180,N_11030);
nor U11933 (N_11933,N_11002,N_11482);
nand U11934 (N_11934,N_11495,N_11370);
nand U11935 (N_11935,N_11314,N_11110);
nor U11936 (N_11936,N_11210,N_11464);
nor U11937 (N_11937,N_11296,N_11269);
nor U11938 (N_11938,N_11056,N_11466);
and U11939 (N_11939,N_11064,N_11317);
or U11940 (N_11940,N_11130,N_11143);
nor U11941 (N_11941,N_11215,N_11160);
nor U11942 (N_11942,N_11435,N_11195);
xor U11943 (N_11943,N_11232,N_11322);
and U11944 (N_11944,N_11067,N_11329);
or U11945 (N_11945,N_11213,N_11060);
nor U11946 (N_11946,N_11253,N_11018);
and U11947 (N_11947,N_11008,N_11483);
or U11948 (N_11948,N_11045,N_11026);
or U11949 (N_11949,N_11077,N_11066);
or U11950 (N_11950,N_11421,N_11488);
and U11951 (N_11951,N_11181,N_11106);
or U11952 (N_11952,N_11335,N_11055);
xor U11953 (N_11953,N_11097,N_11187);
or U11954 (N_11954,N_11289,N_11445);
nand U11955 (N_11955,N_11446,N_11207);
xnor U11956 (N_11956,N_11231,N_11158);
xor U11957 (N_11957,N_11488,N_11193);
xor U11958 (N_11958,N_11491,N_11155);
and U11959 (N_11959,N_11474,N_11390);
or U11960 (N_11960,N_11175,N_11254);
nor U11961 (N_11961,N_11389,N_11378);
nand U11962 (N_11962,N_11293,N_11281);
or U11963 (N_11963,N_11147,N_11433);
or U11964 (N_11964,N_11198,N_11456);
or U11965 (N_11965,N_11017,N_11455);
or U11966 (N_11966,N_11137,N_11135);
or U11967 (N_11967,N_11370,N_11186);
and U11968 (N_11968,N_11237,N_11089);
and U11969 (N_11969,N_11111,N_11052);
nor U11970 (N_11970,N_11059,N_11081);
nand U11971 (N_11971,N_11126,N_11412);
xnor U11972 (N_11972,N_11492,N_11482);
and U11973 (N_11973,N_11364,N_11472);
xnor U11974 (N_11974,N_11436,N_11331);
nand U11975 (N_11975,N_11044,N_11052);
or U11976 (N_11976,N_11119,N_11180);
nor U11977 (N_11977,N_11179,N_11038);
nor U11978 (N_11978,N_11250,N_11296);
or U11979 (N_11979,N_11423,N_11361);
nand U11980 (N_11980,N_11346,N_11451);
xnor U11981 (N_11981,N_11216,N_11427);
and U11982 (N_11982,N_11299,N_11114);
and U11983 (N_11983,N_11020,N_11322);
nor U11984 (N_11984,N_11036,N_11426);
nand U11985 (N_11985,N_11391,N_11293);
xnor U11986 (N_11986,N_11020,N_11283);
nor U11987 (N_11987,N_11033,N_11122);
nand U11988 (N_11988,N_11317,N_11029);
or U11989 (N_11989,N_11249,N_11335);
nand U11990 (N_11990,N_11480,N_11140);
nor U11991 (N_11991,N_11080,N_11313);
nor U11992 (N_11992,N_11410,N_11113);
or U11993 (N_11993,N_11217,N_11182);
nand U11994 (N_11994,N_11485,N_11307);
or U11995 (N_11995,N_11169,N_11477);
or U11996 (N_11996,N_11006,N_11200);
or U11997 (N_11997,N_11437,N_11362);
nor U11998 (N_11998,N_11021,N_11468);
or U11999 (N_11999,N_11005,N_11210);
xor U12000 (N_12000,N_11687,N_11934);
nor U12001 (N_12001,N_11675,N_11800);
xor U12002 (N_12002,N_11691,N_11779);
xnor U12003 (N_12003,N_11791,N_11868);
xor U12004 (N_12004,N_11738,N_11636);
or U12005 (N_12005,N_11917,N_11943);
nand U12006 (N_12006,N_11728,N_11869);
and U12007 (N_12007,N_11511,N_11507);
nand U12008 (N_12008,N_11865,N_11947);
nand U12009 (N_12009,N_11931,N_11935);
xnor U12010 (N_12010,N_11974,N_11645);
nor U12011 (N_12011,N_11912,N_11527);
nor U12012 (N_12012,N_11857,N_11830);
and U12013 (N_12013,N_11977,N_11626);
nand U12014 (N_12014,N_11899,N_11592);
nor U12015 (N_12015,N_11805,N_11590);
or U12016 (N_12016,N_11534,N_11944);
or U12017 (N_12017,N_11674,N_11804);
and U12018 (N_12018,N_11920,N_11818);
and U12019 (N_12019,N_11715,N_11956);
or U12020 (N_12020,N_11753,N_11907);
nor U12021 (N_12021,N_11539,N_11897);
nor U12022 (N_12022,N_11821,N_11562);
xor U12023 (N_12023,N_11593,N_11518);
nand U12024 (N_12024,N_11810,N_11908);
nand U12025 (N_12025,N_11852,N_11996);
xnor U12026 (N_12026,N_11855,N_11789);
nor U12027 (N_12027,N_11754,N_11832);
or U12028 (N_12028,N_11647,N_11723);
and U12029 (N_12029,N_11969,N_11545);
nor U12030 (N_12030,N_11909,N_11929);
nor U12031 (N_12031,N_11811,N_11853);
xnor U12032 (N_12032,N_11762,N_11685);
or U12033 (N_12033,N_11987,N_11550);
nor U12034 (N_12034,N_11758,N_11953);
or U12035 (N_12035,N_11888,N_11631);
xnor U12036 (N_12036,N_11615,N_11793);
xnor U12037 (N_12037,N_11561,N_11981);
xor U12038 (N_12038,N_11538,N_11919);
nor U12039 (N_12039,N_11951,N_11575);
nor U12040 (N_12040,N_11963,N_11748);
and U12041 (N_12041,N_11905,N_11648);
nor U12042 (N_12042,N_11556,N_11960);
nand U12043 (N_12043,N_11672,N_11587);
xor U12044 (N_12044,N_11955,N_11863);
and U12045 (N_12045,N_11773,N_11997);
or U12046 (N_12046,N_11925,N_11620);
or U12047 (N_12047,N_11644,N_11716);
nand U12048 (N_12048,N_11736,N_11559);
and U12049 (N_12049,N_11900,N_11506);
or U12050 (N_12050,N_11973,N_11689);
nand U12051 (N_12051,N_11591,N_11515);
nor U12052 (N_12052,N_11938,N_11928);
nand U12053 (N_12053,N_11597,N_11653);
nor U12054 (N_12054,N_11743,N_11776);
or U12055 (N_12055,N_11967,N_11825);
and U12056 (N_12056,N_11640,N_11734);
nand U12057 (N_12057,N_11598,N_11690);
nand U12058 (N_12058,N_11866,N_11711);
nor U12059 (N_12059,N_11927,N_11623);
and U12060 (N_12060,N_11958,N_11844);
and U12061 (N_12061,N_11815,N_11884);
xnor U12062 (N_12062,N_11764,N_11937);
nor U12063 (N_12063,N_11982,N_11820);
nand U12064 (N_12064,N_11836,N_11721);
nand U12065 (N_12065,N_11979,N_11558);
nor U12066 (N_12066,N_11616,N_11579);
or U12067 (N_12067,N_11998,N_11883);
or U12068 (N_12068,N_11701,N_11509);
xor U12069 (N_12069,N_11601,N_11581);
nand U12070 (N_12070,N_11698,N_11751);
nor U12071 (N_12071,N_11837,N_11708);
or U12072 (N_12072,N_11630,N_11847);
or U12073 (N_12073,N_11795,N_11533);
or U12074 (N_12074,N_11569,N_11911);
nand U12075 (N_12075,N_11681,N_11604);
nor U12076 (N_12076,N_11635,N_11833);
nor U12077 (N_12077,N_11952,N_11964);
and U12078 (N_12078,N_11816,N_11828);
or U12079 (N_12079,N_11642,N_11563);
or U12080 (N_12080,N_11787,N_11633);
nand U12081 (N_12081,N_11877,N_11806);
nand U12082 (N_12082,N_11876,N_11742);
nor U12083 (N_12083,N_11627,N_11880);
xnor U12084 (N_12084,N_11966,N_11885);
or U12085 (N_12085,N_11867,N_11612);
nor U12086 (N_12086,N_11984,N_11763);
xor U12087 (N_12087,N_11817,N_11664);
and U12088 (N_12088,N_11641,N_11582);
nor U12089 (N_12089,N_11812,N_11829);
nor U12090 (N_12090,N_11649,N_11915);
and U12091 (N_12091,N_11896,N_11976);
nand U12092 (N_12092,N_11999,N_11886);
or U12093 (N_12093,N_11891,N_11634);
or U12094 (N_12094,N_11842,N_11946);
and U12095 (N_12095,N_11854,N_11972);
nand U12096 (N_12096,N_11860,N_11991);
or U12097 (N_12097,N_11540,N_11628);
nand U12098 (N_12098,N_11600,N_11898);
and U12099 (N_12099,N_11665,N_11522);
xnor U12100 (N_12100,N_11918,N_11889);
or U12101 (N_12101,N_11676,N_11916);
xor U12102 (N_12102,N_11971,N_11504);
and U12103 (N_12103,N_11894,N_11949);
xnor U12104 (N_12104,N_11731,N_11584);
or U12105 (N_12105,N_11850,N_11528);
and U12106 (N_12106,N_11851,N_11643);
or U12107 (N_12107,N_11835,N_11608);
nand U12108 (N_12108,N_11769,N_11995);
and U12109 (N_12109,N_11679,N_11965);
or U12110 (N_12110,N_11565,N_11605);
or U12111 (N_12111,N_11536,N_11657);
nor U12112 (N_12112,N_11568,N_11726);
xor U12113 (N_12113,N_11710,N_11939);
xor U12114 (N_12114,N_11993,N_11746);
nor U12115 (N_12115,N_11994,N_11864);
or U12116 (N_12116,N_11576,N_11682);
or U12117 (N_12117,N_11555,N_11882);
nor U12118 (N_12118,N_11970,N_11671);
nand U12119 (N_12119,N_11510,N_11872);
nand U12120 (N_12120,N_11503,N_11936);
xnor U12121 (N_12121,N_11759,N_11985);
and U12122 (N_12122,N_11637,N_11992);
nand U12123 (N_12123,N_11923,N_11667);
or U12124 (N_12124,N_11788,N_11525);
nor U12125 (N_12125,N_11839,N_11849);
and U12126 (N_12126,N_11599,N_11914);
nand U12127 (N_12127,N_11890,N_11733);
nand U12128 (N_12128,N_11838,N_11870);
and U12129 (N_12129,N_11501,N_11571);
nor U12130 (N_12130,N_11624,N_11797);
or U12131 (N_12131,N_11941,N_11732);
or U12132 (N_12132,N_11693,N_11529);
nand U12133 (N_12133,N_11695,N_11651);
nand U12134 (N_12134,N_11725,N_11809);
or U12135 (N_12135,N_11703,N_11532);
nand U12136 (N_12136,N_11530,N_11893);
xnor U12137 (N_12137,N_11744,N_11666);
nand U12138 (N_12138,N_11638,N_11989);
nand U12139 (N_12139,N_11574,N_11722);
nor U12140 (N_12140,N_11596,N_11694);
nand U12141 (N_12141,N_11707,N_11735);
xnor U12142 (N_12142,N_11717,N_11547);
nor U12143 (N_12143,N_11611,N_11765);
and U12144 (N_12144,N_11570,N_11901);
xnor U12145 (N_12145,N_11823,N_11546);
or U12146 (N_12146,N_11902,N_11654);
or U12147 (N_12147,N_11807,N_11696);
or U12148 (N_12148,N_11566,N_11803);
nor U12149 (N_12149,N_11517,N_11508);
and U12150 (N_12150,N_11639,N_11606);
xor U12151 (N_12151,N_11777,N_11573);
xor U12152 (N_12152,N_11861,N_11619);
nor U12153 (N_12153,N_11954,N_11712);
xor U12154 (N_12154,N_11609,N_11505);
nand U12155 (N_12155,N_11749,N_11968);
and U12156 (N_12156,N_11756,N_11617);
nand U12157 (N_12157,N_11543,N_11846);
and U12158 (N_12158,N_11680,N_11686);
xnor U12159 (N_12159,N_11551,N_11661);
and U12160 (N_12160,N_11688,N_11845);
and U12161 (N_12161,N_11772,N_11535);
xor U12162 (N_12162,N_11814,N_11990);
and U12163 (N_12163,N_11519,N_11755);
or U12164 (N_12164,N_11771,N_11834);
nor U12165 (N_12165,N_11930,N_11557);
or U12166 (N_12166,N_11502,N_11783);
and U12167 (N_12167,N_11718,N_11841);
and U12168 (N_12168,N_11957,N_11881);
nand U12169 (N_12169,N_11678,N_11782);
and U12170 (N_12170,N_11988,N_11948);
and U12171 (N_12171,N_11613,N_11697);
xor U12172 (N_12172,N_11692,N_11699);
nand U12173 (N_12173,N_11750,N_11516);
xor U12174 (N_12174,N_11719,N_11819);
or U12175 (N_12175,N_11978,N_11942);
or U12176 (N_12176,N_11512,N_11871);
and U12177 (N_12177,N_11781,N_11500);
and U12178 (N_12178,N_11904,N_11760);
nand U12179 (N_12179,N_11727,N_11747);
nor U12180 (N_12180,N_11875,N_11700);
and U12181 (N_12181,N_11632,N_11983);
nor U12182 (N_12182,N_11614,N_11926);
and U12183 (N_12183,N_11745,N_11526);
and U12184 (N_12184,N_11586,N_11521);
nand U12185 (N_12185,N_11858,N_11862);
nand U12186 (N_12186,N_11542,N_11513);
and U12187 (N_12187,N_11741,N_11706);
and U12188 (N_12188,N_11650,N_11794);
or U12189 (N_12189,N_11683,N_11714);
and U12190 (N_12190,N_11702,N_11709);
xnor U12191 (N_12191,N_11652,N_11583);
xor U12192 (N_12192,N_11677,N_11673);
nor U12193 (N_12193,N_11808,N_11713);
and U12194 (N_12194,N_11831,N_11739);
nand U12195 (N_12195,N_11730,N_11729);
xnor U12196 (N_12196,N_11766,N_11924);
nor U12197 (N_12197,N_11541,N_11572);
or U12198 (N_12198,N_11840,N_11775);
and U12199 (N_12199,N_11962,N_11790);
or U12200 (N_12200,N_11553,N_11670);
or U12201 (N_12201,N_11560,N_11906);
or U12202 (N_12202,N_11940,N_11873);
or U12203 (N_12203,N_11813,N_11602);
nor U12204 (N_12204,N_11785,N_11792);
nor U12205 (N_12205,N_11879,N_11887);
or U12206 (N_12206,N_11621,N_11802);
nand U12207 (N_12207,N_11878,N_11520);
nor U12208 (N_12208,N_11577,N_11720);
nor U12209 (N_12209,N_11770,N_11629);
xnor U12210 (N_12210,N_11594,N_11784);
nor U12211 (N_12211,N_11595,N_11655);
xor U12212 (N_12212,N_11778,N_11768);
nor U12213 (N_12213,N_11752,N_11578);
nand U12214 (N_12214,N_11705,N_11827);
xnor U12215 (N_12215,N_11922,N_11589);
and U12216 (N_12216,N_11523,N_11668);
or U12217 (N_12217,N_11903,N_11544);
nand U12218 (N_12218,N_11892,N_11684);
nor U12219 (N_12219,N_11980,N_11514);
nand U12220 (N_12220,N_11859,N_11656);
nand U12221 (N_12221,N_11537,N_11585);
xor U12222 (N_12222,N_11822,N_11824);
or U12223 (N_12223,N_11618,N_11740);
nand U12224 (N_12224,N_11603,N_11625);
nor U12225 (N_12225,N_11801,N_11796);
nand U12226 (N_12226,N_11757,N_11761);
or U12227 (N_12227,N_11856,N_11780);
nor U12228 (N_12228,N_11622,N_11961);
and U12229 (N_12229,N_11895,N_11959);
nand U12230 (N_12230,N_11663,N_11704);
and U12231 (N_12231,N_11986,N_11767);
nor U12232 (N_12232,N_11548,N_11659);
or U12233 (N_12233,N_11932,N_11945);
nor U12234 (N_12234,N_11975,N_11588);
and U12235 (N_12235,N_11564,N_11826);
and U12236 (N_12236,N_11549,N_11843);
or U12237 (N_12237,N_11848,N_11786);
xor U12238 (N_12238,N_11607,N_11921);
nor U12239 (N_12239,N_11524,N_11950);
or U12240 (N_12240,N_11913,N_11646);
or U12241 (N_12241,N_11554,N_11580);
xnor U12242 (N_12242,N_11531,N_11774);
nor U12243 (N_12243,N_11552,N_11910);
nand U12244 (N_12244,N_11610,N_11933);
nor U12245 (N_12245,N_11799,N_11662);
nand U12246 (N_12246,N_11669,N_11724);
or U12247 (N_12247,N_11737,N_11798);
and U12248 (N_12248,N_11874,N_11660);
nor U12249 (N_12249,N_11567,N_11658);
nand U12250 (N_12250,N_11741,N_11648);
or U12251 (N_12251,N_11911,N_11513);
nand U12252 (N_12252,N_11956,N_11758);
xor U12253 (N_12253,N_11998,N_11754);
and U12254 (N_12254,N_11950,N_11500);
xor U12255 (N_12255,N_11939,N_11572);
xor U12256 (N_12256,N_11595,N_11724);
and U12257 (N_12257,N_11961,N_11577);
and U12258 (N_12258,N_11706,N_11530);
nand U12259 (N_12259,N_11774,N_11882);
nor U12260 (N_12260,N_11577,N_11833);
nor U12261 (N_12261,N_11852,N_11946);
and U12262 (N_12262,N_11893,N_11992);
xnor U12263 (N_12263,N_11849,N_11939);
nand U12264 (N_12264,N_11533,N_11789);
and U12265 (N_12265,N_11525,N_11934);
and U12266 (N_12266,N_11989,N_11832);
xor U12267 (N_12267,N_11703,N_11673);
and U12268 (N_12268,N_11822,N_11556);
or U12269 (N_12269,N_11606,N_11817);
and U12270 (N_12270,N_11527,N_11749);
nand U12271 (N_12271,N_11892,N_11634);
nor U12272 (N_12272,N_11821,N_11858);
nor U12273 (N_12273,N_11814,N_11693);
xor U12274 (N_12274,N_11990,N_11936);
xor U12275 (N_12275,N_11579,N_11867);
or U12276 (N_12276,N_11849,N_11606);
or U12277 (N_12277,N_11563,N_11557);
and U12278 (N_12278,N_11984,N_11954);
nand U12279 (N_12279,N_11816,N_11882);
and U12280 (N_12280,N_11541,N_11502);
or U12281 (N_12281,N_11873,N_11926);
and U12282 (N_12282,N_11661,N_11813);
and U12283 (N_12283,N_11670,N_11813);
or U12284 (N_12284,N_11962,N_11508);
nor U12285 (N_12285,N_11743,N_11850);
nand U12286 (N_12286,N_11502,N_11686);
xor U12287 (N_12287,N_11889,N_11733);
nand U12288 (N_12288,N_11800,N_11673);
nor U12289 (N_12289,N_11661,N_11567);
or U12290 (N_12290,N_11629,N_11735);
and U12291 (N_12291,N_11968,N_11831);
and U12292 (N_12292,N_11602,N_11820);
nand U12293 (N_12293,N_11880,N_11989);
xor U12294 (N_12294,N_11515,N_11821);
and U12295 (N_12295,N_11905,N_11946);
and U12296 (N_12296,N_11528,N_11781);
and U12297 (N_12297,N_11545,N_11516);
nand U12298 (N_12298,N_11606,N_11633);
or U12299 (N_12299,N_11891,N_11644);
or U12300 (N_12300,N_11981,N_11802);
and U12301 (N_12301,N_11754,N_11510);
and U12302 (N_12302,N_11689,N_11745);
nor U12303 (N_12303,N_11556,N_11874);
and U12304 (N_12304,N_11577,N_11550);
nor U12305 (N_12305,N_11872,N_11572);
or U12306 (N_12306,N_11560,N_11826);
and U12307 (N_12307,N_11519,N_11658);
and U12308 (N_12308,N_11543,N_11808);
nand U12309 (N_12309,N_11988,N_11892);
or U12310 (N_12310,N_11628,N_11640);
and U12311 (N_12311,N_11612,N_11973);
and U12312 (N_12312,N_11835,N_11580);
xor U12313 (N_12313,N_11955,N_11739);
xor U12314 (N_12314,N_11990,N_11693);
or U12315 (N_12315,N_11666,N_11577);
and U12316 (N_12316,N_11969,N_11550);
nor U12317 (N_12317,N_11962,N_11789);
nand U12318 (N_12318,N_11875,N_11768);
or U12319 (N_12319,N_11664,N_11785);
xnor U12320 (N_12320,N_11642,N_11566);
nor U12321 (N_12321,N_11517,N_11952);
xnor U12322 (N_12322,N_11782,N_11722);
xor U12323 (N_12323,N_11698,N_11569);
nand U12324 (N_12324,N_11638,N_11873);
nand U12325 (N_12325,N_11529,N_11649);
nand U12326 (N_12326,N_11685,N_11599);
or U12327 (N_12327,N_11860,N_11590);
nor U12328 (N_12328,N_11859,N_11914);
and U12329 (N_12329,N_11815,N_11740);
or U12330 (N_12330,N_11611,N_11507);
or U12331 (N_12331,N_11604,N_11816);
or U12332 (N_12332,N_11999,N_11565);
nor U12333 (N_12333,N_11504,N_11555);
and U12334 (N_12334,N_11725,N_11763);
and U12335 (N_12335,N_11778,N_11636);
nor U12336 (N_12336,N_11910,N_11603);
or U12337 (N_12337,N_11536,N_11654);
and U12338 (N_12338,N_11824,N_11978);
and U12339 (N_12339,N_11881,N_11620);
or U12340 (N_12340,N_11833,N_11741);
nor U12341 (N_12341,N_11725,N_11911);
or U12342 (N_12342,N_11714,N_11584);
and U12343 (N_12343,N_11872,N_11983);
nand U12344 (N_12344,N_11590,N_11584);
and U12345 (N_12345,N_11717,N_11926);
and U12346 (N_12346,N_11804,N_11620);
nand U12347 (N_12347,N_11646,N_11533);
xor U12348 (N_12348,N_11919,N_11925);
xnor U12349 (N_12349,N_11585,N_11651);
and U12350 (N_12350,N_11858,N_11514);
or U12351 (N_12351,N_11726,N_11857);
nor U12352 (N_12352,N_11867,N_11762);
nor U12353 (N_12353,N_11840,N_11577);
nor U12354 (N_12354,N_11535,N_11827);
or U12355 (N_12355,N_11938,N_11953);
and U12356 (N_12356,N_11598,N_11651);
or U12357 (N_12357,N_11911,N_11997);
or U12358 (N_12358,N_11653,N_11887);
or U12359 (N_12359,N_11537,N_11688);
and U12360 (N_12360,N_11959,N_11514);
xor U12361 (N_12361,N_11716,N_11936);
and U12362 (N_12362,N_11820,N_11509);
xnor U12363 (N_12363,N_11681,N_11794);
or U12364 (N_12364,N_11749,N_11991);
nor U12365 (N_12365,N_11893,N_11701);
and U12366 (N_12366,N_11636,N_11887);
or U12367 (N_12367,N_11563,N_11544);
nor U12368 (N_12368,N_11563,N_11611);
or U12369 (N_12369,N_11959,N_11875);
xor U12370 (N_12370,N_11760,N_11599);
nor U12371 (N_12371,N_11652,N_11573);
xor U12372 (N_12372,N_11532,N_11625);
nor U12373 (N_12373,N_11807,N_11994);
or U12374 (N_12374,N_11703,N_11818);
nor U12375 (N_12375,N_11944,N_11934);
nand U12376 (N_12376,N_11718,N_11844);
and U12377 (N_12377,N_11798,N_11729);
xnor U12378 (N_12378,N_11811,N_11671);
and U12379 (N_12379,N_11700,N_11575);
nand U12380 (N_12380,N_11996,N_11765);
or U12381 (N_12381,N_11778,N_11764);
nand U12382 (N_12382,N_11923,N_11983);
nand U12383 (N_12383,N_11650,N_11853);
nand U12384 (N_12384,N_11646,N_11600);
xor U12385 (N_12385,N_11589,N_11790);
and U12386 (N_12386,N_11727,N_11604);
nand U12387 (N_12387,N_11617,N_11888);
nor U12388 (N_12388,N_11965,N_11731);
nand U12389 (N_12389,N_11658,N_11657);
and U12390 (N_12390,N_11564,N_11938);
xnor U12391 (N_12391,N_11574,N_11867);
and U12392 (N_12392,N_11775,N_11560);
or U12393 (N_12393,N_11687,N_11675);
nand U12394 (N_12394,N_11918,N_11601);
nor U12395 (N_12395,N_11838,N_11868);
or U12396 (N_12396,N_11560,N_11688);
xnor U12397 (N_12397,N_11853,N_11754);
xnor U12398 (N_12398,N_11917,N_11739);
or U12399 (N_12399,N_11788,N_11838);
xor U12400 (N_12400,N_11845,N_11630);
or U12401 (N_12401,N_11723,N_11561);
and U12402 (N_12402,N_11514,N_11827);
xor U12403 (N_12403,N_11656,N_11645);
or U12404 (N_12404,N_11615,N_11597);
or U12405 (N_12405,N_11506,N_11939);
nor U12406 (N_12406,N_11865,N_11922);
and U12407 (N_12407,N_11863,N_11951);
nor U12408 (N_12408,N_11787,N_11761);
xnor U12409 (N_12409,N_11537,N_11523);
xnor U12410 (N_12410,N_11641,N_11823);
xor U12411 (N_12411,N_11756,N_11947);
xor U12412 (N_12412,N_11607,N_11533);
nand U12413 (N_12413,N_11871,N_11833);
or U12414 (N_12414,N_11793,N_11701);
nor U12415 (N_12415,N_11584,N_11999);
nor U12416 (N_12416,N_11776,N_11979);
xor U12417 (N_12417,N_11925,N_11819);
nand U12418 (N_12418,N_11637,N_11700);
and U12419 (N_12419,N_11999,N_11646);
and U12420 (N_12420,N_11753,N_11652);
nand U12421 (N_12421,N_11508,N_11831);
and U12422 (N_12422,N_11739,N_11918);
nand U12423 (N_12423,N_11843,N_11848);
and U12424 (N_12424,N_11539,N_11584);
nand U12425 (N_12425,N_11505,N_11734);
and U12426 (N_12426,N_11772,N_11987);
xor U12427 (N_12427,N_11746,N_11958);
xor U12428 (N_12428,N_11859,N_11797);
or U12429 (N_12429,N_11601,N_11740);
or U12430 (N_12430,N_11693,N_11854);
nand U12431 (N_12431,N_11960,N_11522);
and U12432 (N_12432,N_11834,N_11600);
nor U12433 (N_12433,N_11554,N_11979);
nor U12434 (N_12434,N_11649,N_11632);
and U12435 (N_12435,N_11622,N_11840);
nand U12436 (N_12436,N_11834,N_11768);
xnor U12437 (N_12437,N_11762,N_11728);
nand U12438 (N_12438,N_11694,N_11844);
nor U12439 (N_12439,N_11647,N_11627);
nand U12440 (N_12440,N_11564,N_11818);
and U12441 (N_12441,N_11862,N_11634);
nor U12442 (N_12442,N_11503,N_11853);
nor U12443 (N_12443,N_11699,N_11903);
nand U12444 (N_12444,N_11868,N_11516);
xor U12445 (N_12445,N_11723,N_11943);
nor U12446 (N_12446,N_11638,N_11624);
nand U12447 (N_12447,N_11883,N_11782);
nand U12448 (N_12448,N_11975,N_11700);
and U12449 (N_12449,N_11599,N_11712);
nand U12450 (N_12450,N_11778,N_11795);
and U12451 (N_12451,N_11865,N_11698);
nor U12452 (N_12452,N_11542,N_11563);
xnor U12453 (N_12453,N_11917,N_11948);
xor U12454 (N_12454,N_11564,N_11700);
or U12455 (N_12455,N_11547,N_11696);
nand U12456 (N_12456,N_11545,N_11554);
or U12457 (N_12457,N_11503,N_11885);
nand U12458 (N_12458,N_11861,N_11532);
or U12459 (N_12459,N_11673,N_11972);
nor U12460 (N_12460,N_11651,N_11707);
or U12461 (N_12461,N_11851,N_11638);
xnor U12462 (N_12462,N_11514,N_11637);
nor U12463 (N_12463,N_11550,N_11575);
or U12464 (N_12464,N_11972,N_11559);
nor U12465 (N_12465,N_11707,N_11939);
nand U12466 (N_12466,N_11666,N_11634);
nor U12467 (N_12467,N_11591,N_11622);
nor U12468 (N_12468,N_11946,N_11845);
nor U12469 (N_12469,N_11900,N_11557);
nor U12470 (N_12470,N_11840,N_11699);
nor U12471 (N_12471,N_11814,N_11978);
xor U12472 (N_12472,N_11729,N_11570);
xor U12473 (N_12473,N_11868,N_11694);
nand U12474 (N_12474,N_11998,N_11542);
and U12475 (N_12475,N_11925,N_11899);
nand U12476 (N_12476,N_11692,N_11916);
and U12477 (N_12477,N_11927,N_11778);
and U12478 (N_12478,N_11721,N_11701);
or U12479 (N_12479,N_11980,N_11910);
and U12480 (N_12480,N_11961,N_11998);
nand U12481 (N_12481,N_11613,N_11736);
nor U12482 (N_12482,N_11767,N_11809);
and U12483 (N_12483,N_11927,N_11677);
xor U12484 (N_12484,N_11973,N_11751);
xor U12485 (N_12485,N_11675,N_11689);
and U12486 (N_12486,N_11709,N_11734);
xor U12487 (N_12487,N_11907,N_11757);
xor U12488 (N_12488,N_11926,N_11628);
xnor U12489 (N_12489,N_11505,N_11759);
nor U12490 (N_12490,N_11917,N_11968);
or U12491 (N_12491,N_11638,N_11589);
and U12492 (N_12492,N_11767,N_11963);
xor U12493 (N_12493,N_11992,N_11685);
or U12494 (N_12494,N_11859,N_11951);
and U12495 (N_12495,N_11702,N_11650);
nor U12496 (N_12496,N_11666,N_11522);
nand U12497 (N_12497,N_11740,N_11823);
or U12498 (N_12498,N_11801,N_11984);
nor U12499 (N_12499,N_11900,N_11614);
and U12500 (N_12500,N_12205,N_12216);
and U12501 (N_12501,N_12400,N_12142);
or U12502 (N_12502,N_12382,N_12024);
and U12503 (N_12503,N_12126,N_12138);
or U12504 (N_12504,N_12094,N_12322);
and U12505 (N_12505,N_12028,N_12344);
and U12506 (N_12506,N_12021,N_12427);
and U12507 (N_12507,N_12303,N_12044);
and U12508 (N_12508,N_12072,N_12281);
nor U12509 (N_12509,N_12485,N_12174);
or U12510 (N_12510,N_12347,N_12495);
nand U12511 (N_12511,N_12135,N_12316);
nand U12512 (N_12512,N_12098,N_12188);
or U12513 (N_12513,N_12484,N_12192);
nor U12514 (N_12514,N_12095,N_12494);
xor U12515 (N_12515,N_12151,N_12114);
or U12516 (N_12516,N_12227,N_12068);
nor U12517 (N_12517,N_12379,N_12388);
xor U12518 (N_12518,N_12050,N_12187);
nor U12519 (N_12519,N_12436,N_12235);
nand U12520 (N_12520,N_12435,N_12224);
nand U12521 (N_12521,N_12118,N_12228);
nor U12522 (N_12522,N_12133,N_12378);
xor U12523 (N_12523,N_12306,N_12023);
nand U12524 (N_12524,N_12444,N_12064);
and U12525 (N_12525,N_12157,N_12487);
nand U12526 (N_12526,N_12014,N_12065);
xnor U12527 (N_12527,N_12083,N_12059);
nand U12528 (N_12528,N_12431,N_12406);
xor U12529 (N_12529,N_12110,N_12343);
nor U12530 (N_12530,N_12348,N_12359);
nand U12531 (N_12531,N_12305,N_12308);
xnor U12532 (N_12532,N_12096,N_12320);
xor U12533 (N_12533,N_12477,N_12450);
or U12534 (N_12534,N_12302,N_12471);
and U12535 (N_12535,N_12200,N_12449);
and U12536 (N_12536,N_12459,N_12461);
nor U12537 (N_12537,N_12319,N_12326);
and U12538 (N_12538,N_12066,N_12409);
and U12539 (N_12539,N_12392,N_12329);
nand U12540 (N_12540,N_12146,N_12060);
nand U12541 (N_12541,N_12411,N_12429);
or U12542 (N_12542,N_12385,N_12036);
nand U12543 (N_12543,N_12264,N_12226);
or U12544 (N_12544,N_12000,N_12152);
or U12545 (N_12545,N_12470,N_12330);
nand U12546 (N_12546,N_12395,N_12207);
or U12547 (N_12547,N_12185,N_12497);
xnor U12548 (N_12548,N_12259,N_12323);
and U12549 (N_12549,N_12015,N_12475);
or U12550 (N_12550,N_12318,N_12310);
nand U12551 (N_12551,N_12209,N_12136);
or U12552 (N_12552,N_12335,N_12258);
or U12553 (N_12553,N_12283,N_12086);
nor U12554 (N_12554,N_12182,N_12147);
or U12555 (N_12555,N_12468,N_12170);
nor U12556 (N_12556,N_12381,N_12440);
xor U12557 (N_12557,N_12054,N_12493);
or U12558 (N_12558,N_12275,N_12332);
or U12559 (N_12559,N_12030,N_12321);
nor U12560 (N_12560,N_12107,N_12001);
and U12561 (N_12561,N_12243,N_12438);
xor U12562 (N_12562,N_12294,N_12109);
nor U12563 (N_12563,N_12043,N_12040);
and U12564 (N_12564,N_12153,N_12102);
xnor U12565 (N_12565,N_12458,N_12353);
nand U12566 (N_12566,N_12422,N_12405);
xnor U12567 (N_12567,N_12082,N_12218);
or U12568 (N_12568,N_12424,N_12012);
xor U12569 (N_12569,N_12402,N_12237);
nand U12570 (N_12570,N_12008,N_12451);
xnor U12571 (N_12571,N_12304,N_12048);
or U12572 (N_12572,N_12181,N_12037);
xor U12573 (N_12573,N_12279,N_12041);
and U12574 (N_12574,N_12499,N_12125);
xor U12575 (N_12575,N_12190,N_12421);
nor U12576 (N_12576,N_12413,N_12467);
nand U12577 (N_12577,N_12139,N_12141);
nand U12578 (N_12578,N_12006,N_12301);
nand U12579 (N_12579,N_12195,N_12180);
or U12580 (N_12580,N_12229,N_12123);
or U12581 (N_12581,N_12293,N_12472);
xor U12582 (N_12582,N_12232,N_12225);
nand U12583 (N_12583,N_12140,N_12375);
and U12584 (N_12584,N_12377,N_12149);
nand U12585 (N_12585,N_12240,N_12105);
xnor U12586 (N_12586,N_12328,N_12437);
nor U12587 (N_12587,N_12013,N_12087);
xor U12588 (N_12588,N_12002,N_12121);
and U12589 (N_12589,N_12313,N_12156);
and U12590 (N_12590,N_12079,N_12277);
nand U12591 (N_12591,N_12069,N_12423);
and U12592 (N_12592,N_12234,N_12291);
and U12593 (N_12593,N_12384,N_12018);
nand U12594 (N_12594,N_12175,N_12492);
xnor U12595 (N_12595,N_12093,N_12331);
or U12596 (N_12596,N_12100,N_12441);
or U12597 (N_12597,N_12389,N_12208);
xnor U12598 (N_12598,N_12434,N_12253);
nand U12599 (N_12599,N_12246,N_12426);
nand U12600 (N_12600,N_12250,N_12496);
nor U12601 (N_12601,N_12158,N_12179);
nor U12602 (N_12602,N_12025,N_12428);
nand U12603 (N_12603,N_12452,N_12124);
nand U12604 (N_12604,N_12113,N_12287);
nand U12605 (N_12605,N_12298,N_12263);
nor U12606 (N_12606,N_12466,N_12349);
nand U12607 (N_12607,N_12486,N_12358);
and U12608 (N_12608,N_12092,N_12333);
nand U12609 (N_12609,N_12202,N_12091);
xor U12610 (N_12610,N_12161,N_12307);
xnor U12611 (N_12611,N_12398,N_12419);
or U12612 (N_12612,N_12111,N_12230);
nor U12613 (N_12613,N_12290,N_12003);
or U12614 (N_12614,N_12249,N_12163);
and U12615 (N_12615,N_12288,N_12233);
or U12616 (N_12616,N_12204,N_12251);
and U12617 (N_12617,N_12296,N_12071);
xnor U12618 (N_12618,N_12193,N_12172);
nand U12619 (N_12619,N_12137,N_12315);
nand U12620 (N_12620,N_12212,N_12324);
nand U12621 (N_12621,N_12143,N_12266);
and U12622 (N_12622,N_12476,N_12401);
or U12623 (N_12623,N_12292,N_12129);
and U12624 (N_12624,N_12289,N_12463);
xnor U12625 (N_12625,N_12254,N_12166);
or U12626 (N_12626,N_12255,N_12311);
or U12627 (N_12627,N_12286,N_12356);
nand U12628 (N_12628,N_12300,N_12346);
nor U12629 (N_12629,N_12155,N_12159);
or U12630 (N_12630,N_12337,N_12352);
nor U12631 (N_12631,N_12242,N_12070);
and U12632 (N_12632,N_12210,N_12061);
or U12633 (N_12633,N_12362,N_12171);
nand U12634 (N_12634,N_12448,N_12122);
or U12635 (N_12635,N_12430,N_12404);
xnor U12636 (N_12636,N_12058,N_12372);
and U12637 (N_12637,N_12414,N_12009);
or U12638 (N_12638,N_12238,N_12005);
xnor U12639 (N_12639,N_12127,N_12017);
or U12640 (N_12640,N_12099,N_12197);
xor U12641 (N_12641,N_12280,N_12269);
or U12642 (N_12642,N_12370,N_12364);
nor U12643 (N_12643,N_12162,N_12177);
xor U12644 (N_12644,N_12183,N_12369);
xor U12645 (N_12645,N_12160,N_12032);
nor U12646 (N_12646,N_12199,N_12261);
and U12647 (N_12647,N_12176,N_12011);
xor U12648 (N_12648,N_12327,N_12273);
nand U12649 (N_12649,N_12101,N_12481);
nand U12650 (N_12650,N_12465,N_12464);
nand U12651 (N_12651,N_12417,N_12154);
nor U12652 (N_12652,N_12407,N_12196);
and U12653 (N_12653,N_12480,N_12057);
nand U12654 (N_12654,N_12265,N_12055);
nand U12655 (N_12655,N_12317,N_12350);
or U12656 (N_12656,N_12173,N_12063);
nand U12657 (N_12657,N_12022,N_12145);
and U12658 (N_12658,N_12272,N_12491);
xnor U12659 (N_12659,N_12164,N_12276);
or U12660 (N_12660,N_12399,N_12239);
nor U12661 (N_12661,N_12046,N_12433);
xor U12662 (N_12662,N_12047,N_12067);
nand U12663 (N_12663,N_12198,N_12189);
nor U12664 (N_12664,N_12144,N_12167);
xnor U12665 (N_12665,N_12020,N_12033);
and U12666 (N_12666,N_12479,N_12203);
nor U12667 (N_12667,N_12034,N_12027);
nand U12668 (N_12668,N_12131,N_12073);
and U12669 (N_12669,N_12412,N_12373);
nor U12670 (N_12670,N_12403,N_12148);
nor U12671 (N_12671,N_12295,N_12045);
xnor U12672 (N_12672,N_12340,N_12446);
or U12673 (N_12673,N_12191,N_12268);
nand U12674 (N_12674,N_12374,N_12488);
xor U12675 (N_12675,N_12038,N_12053);
nor U12676 (N_12676,N_12257,N_12103);
nor U12677 (N_12677,N_12241,N_12049);
nand U12678 (N_12678,N_12090,N_12432);
xnor U12679 (N_12679,N_12278,N_12357);
xnor U12680 (N_12680,N_12483,N_12365);
and U12681 (N_12681,N_12408,N_12222);
or U12682 (N_12682,N_12231,N_12007);
or U12683 (N_12683,N_12325,N_12115);
and U12684 (N_12684,N_12150,N_12097);
nand U12685 (N_12685,N_12425,N_12078);
xor U12686 (N_12686,N_12084,N_12478);
nand U12687 (N_12687,N_12119,N_12267);
nand U12688 (N_12688,N_12285,N_12455);
xnor U12689 (N_12689,N_12474,N_12482);
nor U12690 (N_12690,N_12462,N_12339);
or U12691 (N_12691,N_12355,N_12360);
or U12692 (N_12692,N_12052,N_12415);
nand U12693 (N_12693,N_12074,N_12213);
and U12694 (N_12694,N_12456,N_12080);
and U12695 (N_12695,N_12297,N_12019);
xor U12696 (N_12696,N_12453,N_12442);
nand U12697 (N_12697,N_12390,N_12223);
or U12698 (N_12698,N_12274,N_12178);
and U12699 (N_12699,N_12004,N_12120);
xor U12700 (N_12700,N_12116,N_12186);
nand U12701 (N_12701,N_12108,N_12220);
and U12702 (N_12702,N_12351,N_12056);
nor U12703 (N_12703,N_12393,N_12260);
or U12704 (N_12704,N_12454,N_12397);
nor U12705 (N_12705,N_12312,N_12051);
nand U12706 (N_12706,N_12383,N_12391);
and U12707 (N_12707,N_12029,N_12217);
nand U12708 (N_12708,N_12410,N_12026);
nor U12709 (N_12709,N_12221,N_12284);
nor U12710 (N_12710,N_12387,N_12371);
nor U12711 (N_12711,N_12396,N_12215);
nand U12712 (N_12712,N_12211,N_12081);
nor U12713 (N_12713,N_12016,N_12077);
nand U12714 (N_12714,N_12075,N_12252);
xor U12715 (N_12715,N_12031,N_12342);
and U12716 (N_12716,N_12457,N_12130);
nand U12717 (N_12717,N_12236,N_12117);
or U12718 (N_12718,N_12035,N_12418);
or U12719 (N_12719,N_12194,N_12338);
xor U12720 (N_12720,N_12366,N_12469);
nor U12721 (N_12721,N_12165,N_12394);
xor U12722 (N_12722,N_12345,N_12247);
nand U12723 (N_12723,N_12334,N_12219);
and U12724 (N_12724,N_12244,N_12361);
and U12725 (N_12725,N_12489,N_12245);
nand U12726 (N_12726,N_12104,N_12076);
and U12727 (N_12727,N_12309,N_12443);
or U12728 (N_12728,N_12314,N_12132);
xor U12729 (N_12729,N_12206,N_12184);
nor U12730 (N_12730,N_12439,N_12460);
nor U12731 (N_12731,N_12445,N_12134);
or U12732 (N_12732,N_12128,N_12447);
xor U12733 (N_12733,N_12420,N_12299);
nand U12734 (N_12734,N_12168,N_12112);
and U12735 (N_12735,N_12088,N_12262);
xnor U12736 (N_12736,N_12169,N_12089);
and U12737 (N_12737,N_12380,N_12039);
xor U12738 (N_12738,N_12473,N_12367);
xnor U12739 (N_12739,N_12271,N_12085);
xnor U12740 (N_12740,N_12498,N_12363);
and U12741 (N_12741,N_12062,N_12248);
nor U12742 (N_12742,N_12256,N_12368);
xor U12743 (N_12743,N_12270,N_12376);
xor U12744 (N_12744,N_12354,N_12386);
nand U12745 (N_12745,N_12341,N_12201);
and U12746 (N_12746,N_12282,N_12490);
nor U12747 (N_12747,N_12336,N_12214);
or U12748 (N_12748,N_12416,N_12106);
xnor U12749 (N_12749,N_12010,N_12042);
nor U12750 (N_12750,N_12460,N_12300);
nand U12751 (N_12751,N_12165,N_12103);
or U12752 (N_12752,N_12215,N_12069);
or U12753 (N_12753,N_12420,N_12474);
and U12754 (N_12754,N_12096,N_12019);
xnor U12755 (N_12755,N_12257,N_12396);
nand U12756 (N_12756,N_12068,N_12267);
or U12757 (N_12757,N_12468,N_12068);
and U12758 (N_12758,N_12192,N_12043);
or U12759 (N_12759,N_12134,N_12318);
and U12760 (N_12760,N_12285,N_12148);
or U12761 (N_12761,N_12270,N_12289);
xnor U12762 (N_12762,N_12253,N_12018);
or U12763 (N_12763,N_12059,N_12226);
or U12764 (N_12764,N_12079,N_12254);
and U12765 (N_12765,N_12148,N_12248);
nor U12766 (N_12766,N_12188,N_12024);
nand U12767 (N_12767,N_12154,N_12219);
or U12768 (N_12768,N_12205,N_12041);
xor U12769 (N_12769,N_12080,N_12435);
nand U12770 (N_12770,N_12023,N_12492);
xor U12771 (N_12771,N_12456,N_12207);
nand U12772 (N_12772,N_12244,N_12293);
nor U12773 (N_12773,N_12188,N_12387);
nand U12774 (N_12774,N_12159,N_12400);
and U12775 (N_12775,N_12430,N_12054);
and U12776 (N_12776,N_12238,N_12326);
or U12777 (N_12777,N_12013,N_12304);
and U12778 (N_12778,N_12156,N_12054);
nand U12779 (N_12779,N_12184,N_12385);
or U12780 (N_12780,N_12199,N_12239);
or U12781 (N_12781,N_12024,N_12011);
nor U12782 (N_12782,N_12497,N_12237);
or U12783 (N_12783,N_12360,N_12001);
nand U12784 (N_12784,N_12086,N_12260);
and U12785 (N_12785,N_12102,N_12337);
or U12786 (N_12786,N_12097,N_12170);
nand U12787 (N_12787,N_12484,N_12384);
or U12788 (N_12788,N_12226,N_12148);
xnor U12789 (N_12789,N_12158,N_12355);
and U12790 (N_12790,N_12035,N_12067);
xor U12791 (N_12791,N_12430,N_12086);
and U12792 (N_12792,N_12400,N_12075);
nor U12793 (N_12793,N_12377,N_12276);
nand U12794 (N_12794,N_12319,N_12208);
nand U12795 (N_12795,N_12364,N_12348);
nor U12796 (N_12796,N_12191,N_12183);
and U12797 (N_12797,N_12429,N_12400);
nor U12798 (N_12798,N_12482,N_12064);
and U12799 (N_12799,N_12374,N_12478);
nor U12800 (N_12800,N_12015,N_12063);
nor U12801 (N_12801,N_12489,N_12326);
nand U12802 (N_12802,N_12000,N_12041);
or U12803 (N_12803,N_12116,N_12105);
and U12804 (N_12804,N_12331,N_12298);
xor U12805 (N_12805,N_12327,N_12442);
xnor U12806 (N_12806,N_12006,N_12037);
nor U12807 (N_12807,N_12378,N_12283);
xor U12808 (N_12808,N_12005,N_12090);
and U12809 (N_12809,N_12106,N_12450);
nand U12810 (N_12810,N_12254,N_12308);
nor U12811 (N_12811,N_12293,N_12248);
nor U12812 (N_12812,N_12439,N_12099);
nor U12813 (N_12813,N_12297,N_12102);
nor U12814 (N_12814,N_12143,N_12240);
xor U12815 (N_12815,N_12173,N_12108);
xor U12816 (N_12816,N_12260,N_12085);
nor U12817 (N_12817,N_12283,N_12453);
or U12818 (N_12818,N_12285,N_12119);
xor U12819 (N_12819,N_12259,N_12338);
and U12820 (N_12820,N_12212,N_12277);
or U12821 (N_12821,N_12118,N_12040);
xnor U12822 (N_12822,N_12453,N_12416);
nor U12823 (N_12823,N_12414,N_12487);
nand U12824 (N_12824,N_12013,N_12108);
and U12825 (N_12825,N_12455,N_12064);
xor U12826 (N_12826,N_12027,N_12025);
nor U12827 (N_12827,N_12077,N_12026);
xnor U12828 (N_12828,N_12294,N_12179);
or U12829 (N_12829,N_12198,N_12270);
xnor U12830 (N_12830,N_12258,N_12046);
xnor U12831 (N_12831,N_12009,N_12407);
and U12832 (N_12832,N_12249,N_12143);
or U12833 (N_12833,N_12097,N_12447);
xnor U12834 (N_12834,N_12082,N_12103);
nor U12835 (N_12835,N_12028,N_12267);
nand U12836 (N_12836,N_12132,N_12026);
and U12837 (N_12837,N_12298,N_12386);
nor U12838 (N_12838,N_12039,N_12345);
or U12839 (N_12839,N_12111,N_12457);
and U12840 (N_12840,N_12490,N_12400);
or U12841 (N_12841,N_12203,N_12496);
nand U12842 (N_12842,N_12086,N_12118);
or U12843 (N_12843,N_12159,N_12432);
xor U12844 (N_12844,N_12287,N_12016);
nor U12845 (N_12845,N_12270,N_12310);
nand U12846 (N_12846,N_12370,N_12256);
nand U12847 (N_12847,N_12087,N_12040);
nor U12848 (N_12848,N_12272,N_12027);
xnor U12849 (N_12849,N_12149,N_12210);
xor U12850 (N_12850,N_12264,N_12432);
and U12851 (N_12851,N_12068,N_12136);
and U12852 (N_12852,N_12366,N_12346);
xor U12853 (N_12853,N_12133,N_12238);
xnor U12854 (N_12854,N_12381,N_12030);
xor U12855 (N_12855,N_12228,N_12026);
nor U12856 (N_12856,N_12498,N_12161);
nor U12857 (N_12857,N_12257,N_12044);
nand U12858 (N_12858,N_12032,N_12465);
xnor U12859 (N_12859,N_12428,N_12260);
and U12860 (N_12860,N_12190,N_12315);
and U12861 (N_12861,N_12060,N_12141);
and U12862 (N_12862,N_12064,N_12174);
nor U12863 (N_12863,N_12476,N_12442);
nor U12864 (N_12864,N_12494,N_12155);
nand U12865 (N_12865,N_12142,N_12366);
nand U12866 (N_12866,N_12028,N_12461);
xor U12867 (N_12867,N_12375,N_12095);
nand U12868 (N_12868,N_12276,N_12485);
nand U12869 (N_12869,N_12416,N_12102);
xor U12870 (N_12870,N_12300,N_12101);
nand U12871 (N_12871,N_12108,N_12175);
and U12872 (N_12872,N_12135,N_12091);
xor U12873 (N_12873,N_12368,N_12319);
and U12874 (N_12874,N_12318,N_12450);
xor U12875 (N_12875,N_12368,N_12299);
xor U12876 (N_12876,N_12210,N_12288);
or U12877 (N_12877,N_12384,N_12479);
xnor U12878 (N_12878,N_12112,N_12237);
nand U12879 (N_12879,N_12122,N_12368);
xnor U12880 (N_12880,N_12023,N_12036);
or U12881 (N_12881,N_12031,N_12438);
nor U12882 (N_12882,N_12436,N_12181);
or U12883 (N_12883,N_12088,N_12370);
xor U12884 (N_12884,N_12224,N_12057);
nand U12885 (N_12885,N_12377,N_12134);
xnor U12886 (N_12886,N_12258,N_12495);
and U12887 (N_12887,N_12091,N_12457);
or U12888 (N_12888,N_12363,N_12212);
or U12889 (N_12889,N_12471,N_12224);
xnor U12890 (N_12890,N_12474,N_12247);
or U12891 (N_12891,N_12325,N_12018);
nor U12892 (N_12892,N_12485,N_12478);
xor U12893 (N_12893,N_12476,N_12145);
and U12894 (N_12894,N_12422,N_12484);
or U12895 (N_12895,N_12376,N_12310);
nand U12896 (N_12896,N_12224,N_12013);
or U12897 (N_12897,N_12206,N_12456);
and U12898 (N_12898,N_12430,N_12489);
nand U12899 (N_12899,N_12475,N_12092);
and U12900 (N_12900,N_12216,N_12076);
or U12901 (N_12901,N_12400,N_12185);
xor U12902 (N_12902,N_12391,N_12275);
xnor U12903 (N_12903,N_12007,N_12357);
nand U12904 (N_12904,N_12053,N_12280);
or U12905 (N_12905,N_12170,N_12264);
xor U12906 (N_12906,N_12287,N_12407);
or U12907 (N_12907,N_12016,N_12341);
and U12908 (N_12908,N_12195,N_12445);
or U12909 (N_12909,N_12321,N_12132);
nand U12910 (N_12910,N_12496,N_12497);
xnor U12911 (N_12911,N_12390,N_12210);
and U12912 (N_12912,N_12055,N_12011);
or U12913 (N_12913,N_12439,N_12476);
or U12914 (N_12914,N_12428,N_12218);
nor U12915 (N_12915,N_12316,N_12010);
nand U12916 (N_12916,N_12311,N_12138);
and U12917 (N_12917,N_12007,N_12422);
xnor U12918 (N_12918,N_12046,N_12173);
nor U12919 (N_12919,N_12054,N_12141);
and U12920 (N_12920,N_12433,N_12362);
xnor U12921 (N_12921,N_12031,N_12193);
nand U12922 (N_12922,N_12271,N_12141);
nor U12923 (N_12923,N_12163,N_12126);
nor U12924 (N_12924,N_12010,N_12050);
or U12925 (N_12925,N_12153,N_12031);
nand U12926 (N_12926,N_12236,N_12096);
nor U12927 (N_12927,N_12482,N_12499);
and U12928 (N_12928,N_12362,N_12117);
and U12929 (N_12929,N_12111,N_12119);
or U12930 (N_12930,N_12401,N_12126);
nor U12931 (N_12931,N_12045,N_12173);
nand U12932 (N_12932,N_12238,N_12419);
and U12933 (N_12933,N_12251,N_12148);
xor U12934 (N_12934,N_12120,N_12382);
and U12935 (N_12935,N_12294,N_12306);
nand U12936 (N_12936,N_12121,N_12070);
or U12937 (N_12937,N_12380,N_12253);
or U12938 (N_12938,N_12365,N_12175);
xnor U12939 (N_12939,N_12226,N_12029);
nor U12940 (N_12940,N_12285,N_12208);
or U12941 (N_12941,N_12292,N_12466);
and U12942 (N_12942,N_12454,N_12014);
xor U12943 (N_12943,N_12398,N_12061);
xnor U12944 (N_12944,N_12042,N_12468);
nand U12945 (N_12945,N_12395,N_12181);
or U12946 (N_12946,N_12231,N_12474);
nand U12947 (N_12947,N_12295,N_12215);
or U12948 (N_12948,N_12465,N_12266);
nor U12949 (N_12949,N_12327,N_12007);
or U12950 (N_12950,N_12166,N_12253);
and U12951 (N_12951,N_12015,N_12119);
nor U12952 (N_12952,N_12234,N_12044);
and U12953 (N_12953,N_12453,N_12419);
nor U12954 (N_12954,N_12060,N_12259);
or U12955 (N_12955,N_12259,N_12165);
or U12956 (N_12956,N_12499,N_12172);
and U12957 (N_12957,N_12091,N_12099);
nand U12958 (N_12958,N_12139,N_12063);
or U12959 (N_12959,N_12331,N_12338);
or U12960 (N_12960,N_12394,N_12434);
nor U12961 (N_12961,N_12293,N_12115);
nor U12962 (N_12962,N_12344,N_12286);
nor U12963 (N_12963,N_12130,N_12100);
xnor U12964 (N_12964,N_12164,N_12279);
nor U12965 (N_12965,N_12095,N_12055);
or U12966 (N_12966,N_12456,N_12043);
or U12967 (N_12967,N_12075,N_12004);
and U12968 (N_12968,N_12338,N_12207);
and U12969 (N_12969,N_12474,N_12161);
nor U12970 (N_12970,N_12344,N_12033);
and U12971 (N_12971,N_12311,N_12477);
nand U12972 (N_12972,N_12175,N_12039);
nand U12973 (N_12973,N_12171,N_12386);
or U12974 (N_12974,N_12292,N_12445);
or U12975 (N_12975,N_12470,N_12327);
nand U12976 (N_12976,N_12086,N_12100);
and U12977 (N_12977,N_12093,N_12494);
nand U12978 (N_12978,N_12132,N_12391);
nor U12979 (N_12979,N_12389,N_12279);
and U12980 (N_12980,N_12282,N_12035);
nor U12981 (N_12981,N_12102,N_12477);
nor U12982 (N_12982,N_12484,N_12004);
nand U12983 (N_12983,N_12223,N_12039);
nor U12984 (N_12984,N_12395,N_12150);
or U12985 (N_12985,N_12479,N_12347);
or U12986 (N_12986,N_12435,N_12213);
and U12987 (N_12987,N_12428,N_12122);
nor U12988 (N_12988,N_12051,N_12359);
or U12989 (N_12989,N_12295,N_12420);
or U12990 (N_12990,N_12215,N_12072);
or U12991 (N_12991,N_12211,N_12318);
or U12992 (N_12992,N_12179,N_12037);
xor U12993 (N_12993,N_12232,N_12064);
nor U12994 (N_12994,N_12256,N_12297);
xnor U12995 (N_12995,N_12457,N_12351);
nor U12996 (N_12996,N_12137,N_12355);
xnor U12997 (N_12997,N_12344,N_12457);
xnor U12998 (N_12998,N_12069,N_12297);
nand U12999 (N_12999,N_12173,N_12243);
xnor U13000 (N_13000,N_12979,N_12699);
nor U13001 (N_13001,N_12723,N_12968);
nand U13002 (N_13002,N_12502,N_12836);
and U13003 (N_13003,N_12798,N_12581);
nor U13004 (N_13004,N_12654,N_12986);
or U13005 (N_13005,N_12542,N_12609);
nand U13006 (N_13006,N_12861,N_12557);
nor U13007 (N_13007,N_12693,N_12824);
or U13008 (N_13008,N_12662,N_12500);
nor U13009 (N_13009,N_12527,N_12991);
xnor U13010 (N_13010,N_12620,N_12615);
or U13011 (N_13011,N_12882,N_12994);
or U13012 (N_13012,N_12833,N_12822);
and U13013 (N_13013,N_12807,N_12738);
nor U13014 (N_13014,N_12586,N_12667);
and U13015 (N_13015,N_12672,N_12935);
nand U13016 (N_13016,N_12821,N_12666);
xnor U13017 (N_13017,N_12754,N_12934);
nor U13018 (N_13018,N_12504,N_12990);
nor U13019 (N_13019,N_12685,N_12567);
nor U13020 (N_13020,N_12634,N_12982);
or U13021 (N_13021,N_12701,N_12563);
or U13022 (N_13022,N_12573,N_12903);
nor U13023 (N_13023,N_12963,N_12681);
and U13024 (N_13024,N_12985,N_12704);
and U13025 (N_13025,N_12925,N_12564);
and U13026 (N_13026,N_12971,N_12628);
or U13027 (N_13027,N_12695,N_12651);
or U13028 (N_13028,N_12718,N_12892);
and U13029 (N_13029,N_12605,N_12868);
and U13030 (N_13030,N_12853,N_12977);
or U13031 (N_13031,N_12881,N_12801);
and U13032 (N_13032,N_12682,N_12866);
and U13033 (N_13033,N_12931,N_12817);
nor U13034 (N_13034,N_12538,N_12570);
xnor U13035 (N_13035,N_12629,N_12904);
nor U13036 (N_13036,N_12746,N_12589);
nand U13037 (N_13037,N_12772,N_12552);
or U13038 (N_13038,N_12829,N_12601);
nand U13039 (N_13039,N_12919,N_12785);
xnor U13040 (N_13040,N_12549,N_12956);
nand U13041 (N_13041,N_12593,N_12890);
nand U13042 (N_13042,N_12803,N_12618);
nor U13043 (N_13043,N_12837,N_12722);
and U13044 (N_13044,N_12811,N_12802);
xor U13045 (N_13045,N_12724,N_12870);
xnor U13046 (N_13046,N_12988,N_12550);
xnor U13047 (N_13047,N_12600,N_12747);
xor U13048 (N_13048,N_12731,N_12611);
and U13049 (N_13049,N_12613,N_12729);
and U13050 (N_13050,N_12976,N_12621);
xor U13051 (N_13051,N_12938,N_12595);
and U13052 (N_13052,N_12766,N_12540);
and U13053 (N_13053,N_12865,N_12883);
or U13054 (N_13054,N_12740,N_12920);
or U13055 (N_13055,N_12660,N_12761);
nand U13056 (N_13056,N_12598,N_12503);
and U13057 (N_13057,N_12707,N_12544);
or U13058 (N_13058,N_12716,N_12688);
nor U13059 (N_13059,N_12607,N_12653);
and U13060 (N_13060,N_12973,N_12583);
or U13061 (N_13061,N_12505,N_12838);
or U13062 (N_13062,N_12676,N_12764);
or U13063 (N_13063,N_12794,N_12936);
or U13064 (N_13064,N_12610,N_12584);
nand U13065 (N_13065,N_12683,N_12686);
nand U13066 (N_13066,N_12839,N_12757);
nand U13067 (N_13067,N_12906,N_12874);
and U13068 (N_13068,N_12671,N_12888);
xor U13069 (N_13069,N_12900,N_12663);
xor U13070 (N_13070,N_12594,N_12655);
xnor U13071 (N_13071,N_12674,N_12698);
nor U13072 (N_13072,N_12614,N_12929);
xor U13073 (N_13073,N_12516,N_12733);
or U13074 (N_13074,N_12842,N_12657);
or U13075 (N_13075,N_12548,N_12827);
xor U13076 (N_13076,N_12849,N_12534);
and U13077 (N_13077,N_12518,N_12526);
and U13078 (N_13078,N_12792,N_12898);
or U13079 (N_13079,N_12645,N_12820);
and U13080 (N_13080,N_12575,N_12725);
or U13081 (N_13081,N_12665,N_12913);
or U13082 (N_13082,N_12649,N_12640);
nor U13083 (N_13083,N_12889,N_12560);
xnor U13084 (N_13084,N_12886,N_12891);
nand U13085 (N_13085,N_12744,N_12750);
nand U13086 (N_13086,N_12790,N_12636);
nor U13087 (N_13087,N_12546,N_12514);
nor U13088 (N_13088,N_12727,N_12940);
nor U13089 (N_13089,N_12694,N_12751);
xnor U13090 (N_13090,N_12510,N_12901);
xor U13091 (N_13091,N_12709,N_12561);
and U13092 (N_13092,N_12847,N_12533);
nand U13093 (N_13093,N_12808,N_12714);
xor U13094 (N_13094,N_12644,N_12659);
nand U13095 (N_13095,N_12530,N_12748);
xnor U13096 (N_13096,N_12713,N_12577);
and U13097 (N_13097,N_12582,N_12742);
xnor U13098 (N_13098,N_12781,N_12675);
or U13099 (N_13099,N_12843,N_12623);
xor U13100 (N_13100,N_12871,N_12869);
xnor U13101 (N_13101,N_12953,N_12543);
nand U13102 (N_13102,N_12622,N_12630);
xor U13103 (N_13103,N_12780,N_12765);
and U13104 (N_13104,N_12983,N_12535);
nand U13105 (N_13105,N_12749,N_12728);
nand U13106 (N_13106,N_12778,N_12668);
nand U13107 (N_13107,N_12914,N_12517);
or U13108 (N_13108,N_12545,N_12773);
xnor U13109 (N_13109,N_12720,N_12952);
nor U13110 (N_13110,N_12632,N_12819);
and U13111 (N_13111,N_12721,N_12943);
or U13112 (N_13112,N_12831,N_12834);
nand U13113 (N_13113,N_12887,N_12933);
and U13114 (N_13114,N_12856,N_12715);
or U13115 (N_13115,N_12958,N_12736);
or U13116 (N_13116,N_12854,N_12558);
or U13117 (N_13117,N_12588,N_12812);
or U13118 (N_13118,N_12522,N_12612);
and U13119 (N_13119,N_12814,N_12585);
or U13120 (N_13120,N_12760,N_12692);
xor U13121 (N_13121,N_12680,N_12597);
or U13122 (N_13122,N_12996,N_12762);
nor U13123 (N_13123,N_12712,N_12506);
nand U13124 (N_13124,N_12818,N_12587);
nand U13125 (N_13125,N_12771,N_12711);
nor U13126 (N_13126,N_12578,N_12945);
xnor U13127 (N_13127,N_12603,N_12816);
or U13128 (N_13128,N_12921,N_12826);
nand U13129 (N_13129,N_12909,N_12697);
and U13130 (N_13130,N_12507,N_12590);
nand U13131 (N_13131,N_12551,N_12974);
nand U13132 (N_13132,N_12939,N_12813);
xnor U13133 (N_13133,N_12599,N_12998);
nand U13134 (N_13134,N_12975,N_12775);
nand U13135 (N_13135,N_12702,N_12776);
and U13136 (N_13136,N_12965,N_12860);
nand U13137 (N_13137,N_12689,N_12596);
nand U13138 (N_13138,N_12783,N_12930);
and U13139 (N_13139,N_12574,N_12743);
and U13140 (N_13140,N_12539,N_12878);
or U13141 (N_13141,N_12922,N_12911);
nand U13142 (N_13142,N_12606,N_12896);
and U13143 (N_13143,N_12917,N_12893);
nand U13144 (N_13144,N_12806,N_12602);
and U13145 (N_13145,N_12541,N_12732);
nor U13146 (N_13146,N_12905,N_12559);
xor U13147 (N_13147,N_12608,N_12524);
or U13148 (N_13148,N_12954,N_12823);
nor U13149 (N_13149,N_12670,N_12705);
or U13150 (N_13150,N_12993,N_12850);
nand U13151 (N_13151,N_12815,N_12787);
xnor U13152 (N_13152,N_12571,N_12924);
nand U13153 (N_13153,N_12664,N_12719);
nor U13154 (N_13154,N_12568,N_12942);
and U13155 (N_13155,N_12832,N_12679);
nand U13156 (N_13156,N_12637,N_12992);
nand U13157 (N_13157,N_12912,N_12959);
nand U13158 (N_13158,N_12797,N_12997);
xnor U13159 (N_13159,N_12946,N_12923);
nor U13160 (N_13160,N_12995,N_12638);
and U13161 (N_13161,N_12684,N_12619);
nand U13162 (N_13162,N_12885,N_12528);
nor U13163 (N_13163,N_12768,N_12782);
nor U13164 (N_13164,N_12576,N_12937);
xnor U13165 (N_13165,N_12691,N_12572);
xnor U13166 (N_13166,N_12647,N_12875);
nand U13167 (N_13167,N_12753,N_12512);
xnor U13168 (N_13168,N_12795,N_12627);
or U13169 (N_13169,N_12916,N_12737);
nand U13170 (N_13170,N_12981,N_12678);
nor U13171 (N_13171,N_12767,N_12643);
nor U13172 (N_13172,N_12579,N_12846);
xnor U13173 (N_13173,N_12537,N_12523);
xnor U13174 (N_13174,N_12915,N_12932);
xor U13175 (N_13175,N_12918,N_12774);
or U13176 (N_13176,N_12966,N_12756);
nand U13177 (N_13177,N_12957,N_12509);
nor U13178 (N_13178,N_12970,N_12745);
nand U13179 (N_13179,N_12984,N_12784);
xnor U13180 (N_13180,N_12927,N_12648);
or U13181 (N_13181,N_12501,N_12859);
nand U13182 (N_13182,N_12562,N_12789);
nand U13183 (N_13183,N_12658,N_12592);
xnor U13184 (N_13184,N_12960,N_12763);
xnor U13185 (N_13185,N_12706,N_12964);
and U13186 (N_13186,N_12703,N_12828);
or U13187 (N_13187,N_12641,N_12752);
xor U13188 (N_13188,N_12687,N_12642);
nor U13189 (N_13189,N_12978,N_12639);
or U13190 (N_13190,N_12532,N_12989);
nand U13191 (N_13191,N_12793,N_12565);
nand U13192 (N_13192,N_12730,N_12734);
nand U13193 (N_13193,N_12758,N_12513);
and U13194 (N_13194,N_12877,N_12910);
nand U13195 (N_13195,N_12962,N_12786);
and U13196 (N_13196,N_12536,N_12656);
and U13197 (N_13197,N_12830,N_12791);
nor U13198 (N_13198,N_12616,N_12858);
or U13199 (N_13199,N_12626,N_12961);
xnor U13200 (N_13200,N_12999,N_12520);
nand U13201 (N_13201,N_12947,N_12708);
xor U13202 (N_13202,N_12553,N_12604);
xnor U13203 (N_13203,N_12862,N_12805);
nor U13204 (N_13204,N_12863,N_12873);
nor U13205 (N_13205,N_12969,N_12769);
xnor U13206 (N_13206,N_12710,N_12788);
and U13207 (N_13207,N_12897,N_12726);
or U13208 (N_13208,N_12796,N_12580);
nor U13209 (N_13209,N_12677,N_12741);
or U13210 (N_13210,N_12569,N_12696);
nor U13211 (N_13211,N_12884,N_12944);
nand U13212 (N_13212,N_12739,N_12880);
or U13213 (N_13213,N_12625,N_12799);
and U13214 (N_13214,N_12700,N_12872);
and U13215 (N_13215,N_12972,N_12646);
and U13216 (N_13216,N_12948,N_12717);
xor U13217 (N_13217,N_12661,N_12809);
nor U13218 (N_13218,N_12690,N_12650);
nor U13219 (N_13219,N_12508,N_12907);
and U13220 (N_13220,N_12902,N_12857);
xor U13221 (N_13221,N_12669,N_12556);
nor U13222 (N_13222,N_12851,N_12804);
xnor U13223 (N_13223,N_12735,N_12554);
nand U13224 (N_13224,N_12840,N_12531);
or U13225 (N_13225,N_12908,N_12519);
and U13226 (N_13226,N_12800,N_12779);
nand U13227 (N_13227,N_12899,N_12928);
nand U13228 (N_13228,N_12951,N_12864);
xor U13229 (N_13229,N_12825,N_12926);
nor U13230 (N_13230,N_12624,N_12652);
and U13231 (N_13231,N_12879,N_12950);
or U13232 (N_13232,N_12810,N_12759);
nand U13233 (N_13233,N_12949,N_12835);
and U13234 (N_13234,N_12980,N_12967);
nand U13235 (N_13235,N_12755,N_12955);
nor U13236 (N_13236,N_12515,N_12631);
nor U13237 (N_13237,N_12867,N_12777);
or U13238 (N_13238,N_12617,N_12848);
or U13239 (N_13239,N_12566,N_12841);
xor U13240 (N_13240,N_12525,N_12511);
xnor U13241 (N_13241,N_12633,N_12852);
and U13242 (N_13242,N_12895,N_12941);
or U13243 (N_13243,N_12844,N_12770);
and U13244 (N_13244,N_12635,N_12673);
or U13245 (N_13245,N_12876,N_12591);
or U13246 (N_13246,N_12521,N_12529);
or U13247 (N_13247,N_12894,N_12855);
nor U13248 (N_13248,N_12555,N_12845);
nand U13249 (N_13249,N_12987,N_12547);
xnor U13250 (N_13250,N_12788,N_12601);
nand U13251 (N_13251,N_12664,N_12730);
xor U13252 (N_13252,N_12897,N_12810);
or U13253 (N_13253,N_12534,N_12854);
or U13254 (N_13254,N_12871,N_12794);
and U13255 (N_13255,N_12668,N_12871);
and U13256 (N_13256,N_12946,N_12995);
and U13257 (N_13257,N_12606,N_12548);
or U13258 (N_13258,N_12793,N_12506);
or U13259 (N_13259,N_12526,N_12757);
nor U13260 (N_13260,N_12634,N_12670);
nor U13261 (N_13261,N_12906,N_12640);
or U13262 (N_13262,N_12708,N_12799);
nor U13263 (N_13263,N_12798,N_12695);
nor U13264 (N_13264,N_12761,N_12827);
or U13265 (N_13265,N_12678,N_12927);
or U13266 (N_13266,N_12597,N_12594);
nor U13267 (N_13267,N_12514,N_12859);
and U13268 (N_13268,N_12578,N_12869);
nor U13269 (N_13269,N_12731,N_12732);
or U13270 (N_13270,N_12989,N_12850);
and U13271 (N_13271,N_12730,N_12525);
xnor U13272 (N_13272,N_12613,N_12836);
xor U13273 (N_13273,N_12795,N_12787);
nand U13274 (N_13274,N_12664,N_12905);
xor U13275 (N_13275,N_12615,N_12521);
nor U13276 (N_13276,N_12874,N_12600);
nor U13277 (N_13277,N_12631,N_12534);
nor U13278 (N_13278,N_12884,N_12516);
or U13279 (N_13279,N_12783,N_12910);
nand U13280 (N_13280,N_12942,N_12514);
xnor U13281 (N_13281,N_12881,N_12637);
or U13282 (N_13282,N_12945,N_12576);
nand U13283 (N_13283,N_12822,N_12625);
nand U13284 (N_13284,N_12673,N_12927);
nand U13285 (N_13285,N_12927,N_12844);
and U13286 (N_13286,N_12669,N_12760);
and U13287 (N_13287,N_12522,N_12500);
xor U13288 (N_13288,N_12864,N_12588);
xor U13289 (N_13289,N_12873,N_12794);
nand U13290 (N_13290,N_12916,N_12632);
xnor U13291 (N_13291,N_12785,N_12584);
nand U13292 (N_13292,N_12673,N_12595);
nor U13293 (N_13293,N_12505,N_12557);
or U13294 (N_13294,N_12898,N_12999);
and U13295 (N_13295,N_12560,N_12800);
nor U13296 (N_13296,N_12559,N_12732);
xor U13297 (N_13297,N_12822,N_12619);
xor U13298 (N_13298,N_12502,N_12578);
xor U13299 (N_13299,N_12890,N_12978);
xnor U13300 (N_13300,N_12724,N_12655);
nand U13301 (N_13301,N_12896,N_12777);
xor U13302 (N_13302,N_12741,N_12512);
nor U13303 (N_13303,N_12544,N_12833);
xor U13304 (N_13304,N_12734,N_12938);
nor U13305 (N_13305,N_12754,N_12858);
nor U13306 (N_13306,N_12965,N_12800);
nand U13307 (N_13307,N_12812,N_12679);
nor U13308 (N_13308,N_12881,N_12650);
nand U13309 (N_13309,N_12966,N_12903);
or U13310 (N_13310,N_12795,N_12708);
xnor U13311 (N_13311,N_12640,N_12710);
nor U13312 (N_13312,N_12690,N_12506);
xnor U13313 (N_13313,N_12511,N_12921);
or U13314 (N_13314,N_12507,N_12573);
xor U13315 (N_13315,N_12944,N_12610);
and U13316 (N_13316,N_12816,N_12543);
nor U13317 (N_13317,N_12734,N_12683);
or U13318 (N_13318,N_12796,N_12651);
or U13319 (N_13319,N_12751,N_12606);
and U13320 (N_13320,N_12936,N_12514);
xor U13321 (N_13321,N_12676,N_12919);
xor U13322 (N_13322,N_12913,N_12647);
nor U13323 (N_13323,N_12503,N_12996);
or U13324 (N_13324,N_12812,N_12621);
xnor U13325 (N_13325,N_12867,N_12805);
or U13326 (N_13326,N_12760,N_12681);
or U13327 (N_13327,N_12920,N_12665);
nor U13328 (N_13328,N_12779,N_12661);
xnor U13329 (N_13329,N_12916,N_12927);
nand U13330 (N_13330,N_12835,N_12530);
nand U13331 (N_13331,N_12510,N_12505);
xor U13332 (N_13332,N_12648,N_12705);
nor U13333 (N_13333,N_12818,N_12789);
and U13334 (N_13334,N_12725,N_12707);
and U13335 (N_13335,N_12560,N_12850);
xor U13336 (N_13336,N_12670,N_12566);
and U13337 (N_13337,N_12683,N_12664);
nor U13338 (N_13338,N_12767,N_12615);
nor U13339 (N_13339,N_12504,N_12576);
nand U13340 (N_13340,N_12676,N_12701);
or U13341 (N_13341,N_12692,N_12983);
or U13342 (N_13342,N_12800,N_12863);
nand U13343 (N_13343,N_12859,N_12938);
nor U13344 (N_13344,N_12593,N_12969);
xnor U13345 (N_13345,N_12633,N_12900);
nand U13346 (N_13346,N_12809,N_12791);
xnor U13347 (N_13347,N_12895,N_12716);
nand U13348 (N_13348,N_12893,N_12537);
nor U13349 (N_13349,N_12901,N_12803);
or U13350 (N_13350,N_12924,N_12942);
nor U13351 (N_13351,N_12832,N_12592);
nor U13352 (N_13352,N_12698,N_12892);
or U13353 (N_13353,N_12995,N_12798);
xnor U13354 (N_13354,N_12751,N_12834);
nand U13355 (N_13355,N_12680,N_12614);
nand U13356 (N_13356,N_12925,N_12690);
or U13357 (N_13357,N_12609,N_12601);
and U13358 (N_13358,N_12983,N_12622);
or U13359 (N_13359,N_12923,N_12519);
nor U13360 (N_13360,N_12987,N_12586);
xnor U13361 (N_13361,N_12683,N_12892);
nor U13362 (N_13362,N_12742,N_12903);
or U13363 (N_13363,N_12888,N_12972);
or U13364 (N_13364,N_12527,N_12713);
xor U13365 (N_13365,N_12674,N_12568);
and U13366 (N_13366,N_12924,N_12600);
nand U13367 (N_13367,N_12941,N_12769);
and U13368 (N_13368,N_12582,N_12947);
and U13369 (N_13369,N_12920,N_12867);
nand U13370 (N_13370,N_12846,N_12897);
nand U13371 (N_13371,N_12818,N_12915);
nand U13372 (N_13372,N_12856,N_12501);
nand U13373 (N_13373,N_12582,N_12887);
nand U13374 (N_13374,N_12982,N_12852);
xor U13375 (N_13375,N_12594,N_12675);
nor U13376 (N_13376,N_12610,N_12972);
and U13377 (N_13377,N_12630,N_12543);
and U13378 (N_13378,N_12738,N_12831);
nor U13379 (N_13379,N_12779,N_12915);
or U13380 (N_13380,N_12675,N_12882);
xnor U13381 (N_13381,N_12505,N_12984);
xor U13382 (N_13382,N_12838,N_12541);
nand U13383 (N_13383,N_12561,N_12827);
xor U13384 (N_13384,N_12892,N_12651);
nand U13385 (N_13385,N_12927,N_12764);
nor U13386 (N_13386,N_12831,N_12792);
and U13387 (N_13387,N_12985,N_12935);
xnor U13388 (N_13388,N_12995,N_12654);
nor U13389 (N_13389,N_12548,N_12975);
nor U13390 (N_13390,N_12883,N_12930);
and U13391 (N_13391,N_12974,N_12772);
or U13392 (N_13392,N_12882,N_12884);
and U13393 (N_13393,N_12553,N_12518);
nor U13394 (N_13394,N_12928,N_12581);
or U13395 (N_13395,N_12948,N_12672);
xnor U13396 (N_13396,N_12613,N_12529);
xnor U13397 (N_13397,N_12590,N_12503);
or U13398 (N_13398,N_12958,N_12873);
nand U13399 (N_13399,N_12858,N_12785);
and U13400 (N_13400,N_12661,N_12865);
nand U13401 (N_13401,N_12648,N_12630);
or U13402 (N_13402,N_12990,N_12651);
xnor U13403 (N_13403,N_12659,N_12900);
or U13404 (N_13404,N_12966,N_12595);
or U13405 (N_13405,N_12712,N_12597);
nand U13406 (N_13406,N_12990,N_12552);
and U13407 (N_13407,N_12919,N_12767);
xor U13408 (N_13408,N_12728,N_12515);
nand U13409 (N_13409,N_12671,N_12713);
nand U13410 (N_13410,N_12535,N_12941);
nand U13411 (N_13411,N_12726,N_12665);
nand U13412 (N_13412,N_12897,N_12896);
xor U13413 (N_13413,N_12518,N_12636);
nor U13414 (N_13414,N_12623,N_12664);
or U13415 (N_13415,N_12645,N_12532);
nor U13416 (N_13416,N_12963,N_12977);
xor U13417 (N_13417,N_12619,N_12950);
or U13418 (N_13418,N_12782,N_12853);
or U13419 (N_13419,N_12924,N_12624);
xor U13420 (N_13420,N_12659,N_12768);
nand U13421 (N_13421,N_12634,N_12548);
nand U13422 (N_13422,N_12654,N_12916);
or U13423 (N_13423,N_12533,N_12518);
xnor U13424 (N_13424,N_12877,N_12613);
nor U13425 (N_13425,N_12738,N_12715);
xor U13426 (N_13426,N_12813,N_12758);
nor U13427 (N_13427,N_12764,N_12821);
xnor U13428 (N_13428,N_12598,N_12690);
or U13429 (N_13429,N_12564,N_12704);
and U13430 (N_13430,N_12609,N_12641);
nor U13431 (N_13431,N_12875,N_12926);
nor U13432 (N_13432,N_12841,N_12770);
or U13433 (N_13433,N_12580,N_12616);
nor U13434 (N_13434,N_12910,N_12822);
or U13435 (N_13435,N_12988,N_12581);
xor U13436 (N_13436,N_12903,N_12727);
xnor U13437 (N_13437,N_12948,N_12636);
and U13438 (N_13438,N_12932,N_12618);
nor U13439 (N_13439,N_12991,N_12834);
xor U13440 (N_13440,N_12866,N_12727);
nand U13441 (N_13441,N_12531,N_12872);
xor U13442 (N_13442,N_12920,N_12733);
or U13443 (N_13443,N_12902,N_12880);
or U13444 (N_13444,N_12725,N_12976);
or U13445 (N_13445,N_12597,N_12674);
and U13446 (N_13446,N_12833,N_12889);
and U13447 (N_13447,N_12921,N_12984);
or U13448 (N_13448,N_12869,N_12653);
nor U13449 (N_13449,N_12877,N_12677);
and U13450 (N_13450,N_12986,N_12509);
nor U13451 (N_13451,N_12966,N_12751);
nor U13452 (N_13452,N_12760,N_12945);
xor U13453 (N_13453,N_12776,N_12513);
and U13454 (N_13454,N_12894,N_12530);
or U13455 (N_13455,N_12780,N_12993);
or U13456 (N_13456,N_12988,N_12868);
xnor U13457 (N_13457,N_12523,N_12629);
xnor U13458 (N_13458,N_12661,N_12863);
and U13459 (N_13459,N_12837,N_12542);
or U13460 (N_13460,N_12517,N_12787);
and U13461 (N_13461,N_12808,N_12761);
nand U13462 (N_13462,N_12504,N_12935);
nor U13463 (N_13463,N_12616,N_12573);
xor U13464 (N_13464,N_12686,N_12960);
and U13465 (N_13465,N_12799,N_12973);
xor U13466 (N_13466,N_12698,N_12804);
xor U13467 (N_13467,N_12711,N_12989);
or U13468 (N_13468,N_12705,N_12681);
or U13469 (N_13469,N_12668,N_12959);
nand U13470 (N_13470,N_12638,N_12661);
and U13471 (N_13471,N_12582,N_12553);
nor U13472 (N_13472,N_12722,N_12925);
or U13473 (N_13473,N_12837,N_12761);
or U13474 (N_13474,N_12940,N_12621);
nor U13475 (N_13475,N_12589,N_12983);
nand U13476 (N_13476,N_12676,N_12720);
nor U13477 (N_13477,N_12507,N_12757);
or U13478 (N_13478,N_12806,N_12933);
nand U13479 (N_13479,N_12933,N_12675);
nor U13480 (N_13480,N_12658,N_12806);
nand U13481 (N_13481,N_12988,N_12713);
or U13482 (N_13482,N_12759,N_12738);
and U13483 (N_13483,N_12570,N_12605);
xor U13484 (N_13484,N_12603,N_12557);
xor U13485 (N_13485,N_12536,N_12843);
nor U13486 (N_13486,N_12617,N_12966);
nor U13487 (N_13487,N_12621,N_12713);
nor U13488 (N_13488,N_12693,N_12683);
nand U13489 (N_13489,N_12792,N_12786);
or U13490 (N_13490,N_12872,N_12653);
xnor U13491 (N_13491,N_12590,N_12530);
and U13492 (N_13492,N_12767,N_12698);
or U13493 (N_13493,N_12822,N_12864);
or U13494 (N_13494,N_12961,N_12786);
or U13495 (N_13495,N_12795,N_12605);
xor U13496 (N_13496,N_12661,N_12709);
and U13497 (N_13497,N_12719,N_12780);
and U13498 (N_13498,N_12966,N_12767);
xnor U13499 (N_13499,N_12633,N_12677);
xnor U13500 (N_13500,N_13044,N_13076);
nor U13501 (N_13501,N_13100,N_13167);
xnor U13502 (N_13502,N_13374,N_13348);
xor U13503 (N_13503,N_13036,N_13081);
nor U13504 (N_13504,N_13109,N_13275);
nand U13505 (N_13505,N_13042,N_13116);
nand U13506 (N_13506,N_13331,N_13318);
and U13507 (N_13507,N_13032,N_13266);
xnor U13508 (N_13508,N_13020,N_13435);
nand U13509 (N_13509,N_13096,N_13367);
nor U13510 (N_13510,N_13199,N_13261);
and U13511 (N_13511,N_13077,N_13064);
xor U13512 (N_13512,N_13004,N_13383);
xor U13513 (N_13513,N_13001,N_13097);
nor U13514 (N_13514,N_13115,N_13466);
xnor U13515 (N_13515,N_13169,N_13016);
and U13516 (N_13516,N_13457,N_13163);
nand U13517 (N_13517,N_13024,N_13217);
xnor U13518 (N_13518,N_13089,N_13084);
xnor U13519 (N_13519,N_13280,N_13062);
and U13520 (N_13520,N_13083,N_13472);
xor U13521 (N_13521,N_13209,N_13030);
xnor U13522 (N_13522,N_13498,N_13464);
nor U13523 (N_13523,N_13304,N_13104);
xnor U13524 (N_13524,N_13182,N_13018);
nand U13525 (N_13525,N_13454,N_13067);
nor U13526 (N_13526,N_13279,N_13238);
nor U13527 (N_13527,N_13229,N_13282);
xor U13528 (N_13528,N_13090,N_13372);
nand U13529 (N_13529,N_13392,N_13002);
nor U13530 (N_13530,N_13074,N_13135);
and U13531 (N_13531,N_13215,N_13206);
and U13532 (N_13532,N_13327,N_13223);
and U13533 (N_13533,N_13330,N_13160);
or U13534 (N_13534,N_13311,N_13333);
nor U13535 (N_13535,N_13164,N_13156);
and U13536 (N_13536,N_13134,N_13469);
xnor U13537 (N_13537,N_13099,N_13259);
nor U13538 (N_13538,N_13413,N_13336);
nor U13539 (N_13539,N_13176,N_13225);
and U13540 (N_13540,N_13026,N_13143);
xor U13541 (N_13541,N_13031,N_13071);
or U13542 (N_13542,N_13483,N_13384);
or U13543 (N_13543,N_13029,N_13468);
or U13544 (N_13544,N_13411,N_13147);
and U13545 (N_13545,N_13010,N_13086);
nand U13546 (N_13546,N_13178,N_13356);
and U13547 (N_13547,N_13398,N_13401);
and U13548 (N_13548,N_13495,N_13276);
and U13549 (N_13549,N_13226,N_13270);
or U13550 (N_13550,N_13066,N_13428);
nand U13551 (N_13551,N_13354,N_13375);
xnor U13552 (N_13552,N_13475,N_13341);
and U13553 (N_13553,N_13204,N_13378);
or U13554 (N_13554,N_13052,N_13055);
nor U13555 (N_13555,N_13414,N_13349);
xnor U13556 (N_13556,N_13257,N_13192);
and U13557 (N_13557,N_13335,N_13347);
xor U13558 (N_13558,N_13023,N_13014);
xor U13559 (N_13559,N_13314,N_13344);
nand U13560 (N_13560,N_13301,N_13049);
xnor U13561 (N_13561,N_13012,N_13079);
nor U13562 (N_13562,N_13456,N_13309);
xnor U13563 (N_13563,N_13091,N_13343);
and U13564 (N_13564,N_13442,N_13120);
and U13565 (N_13565,N_13073,N_13465);
xnor U13566 (N_13566,N_13022,N_13037);
and U13567 (N_13567,N_13230,N_13438);
or U13568 (N_13568,N_13153,N_13476);
and U13569 (N_13569,N_13114,N_13441);
and U13570 (N_13570,N_13048,N_13019);
and U13571 (N_13571,N_13264,N_13339);
xnor U13572 (N_13572,N_13286,N_13009);
nor U13573 (N_13573,N_13350,N_13497);
and U13574 (N_13574,N_13158,N_13122);
and U13575 (N_13575,N_13272,N_13306);
and U13576 (N_13576,N_13373,N_13346);
nor U13577 (N_13577,N_13111,N_13034);
and U13578 (N_13578,N_13144,N_13072);
nand U13579 (N_13579,N_13486,N_13364);
nor U13580 (N_13580,N_13103,N_13208);
or U13581 (N_13581,N_13060,N_13434);
or U13582 (N_13582,N_13202,N_13363);
and U13583 (N_13583,N_13105,N_13235);
or U13584 (N_13584,N_13488,N_13271);
nor U13585 (N_13585,N_13345,N_13180);
or U13586 (N_13586,N_13119,N_13239);
or U13587 (N_13587,N_13439,N_13462);
or U13588 (N_13588,N_13210,N_13485);
or U13589 (N_13589,N_13360,N_13050);
nand U13590 (N_13590,N_13278,N_13234);
xor U13591 (N_13591,N_13431,N_13017);
nand U13592 (N_13592,N_13420,N_13289);
or U13593 (N_13593,N_13492,N_13222);
nand U13594 (N_13594,N_13075,N_13008);
nand U13595 (N_13595,N_13013,N_13139);
nor U13596 (N_13596,N_13007,N_13426);
nor U13597 (N_13597,N_13386,N_13455);
nor U13598 (N_13598,N_13387,N_13186);
and U13599 (N_13599,N_13214,N_13342);
xor U13600 (N_13600,N_13452,N_13292);
nor U13601 (N_13601,N_13285,N_13437);
xnor U13602 (N_13602,N_13124,N_13481);
and U13603 (N_13603,N_13394,N_13358);
or U13604 (N_13604,N_13220,N_13027);
xnor U13605 (N_13605,N_13250,N_13005);
and U13606 (N_13606,N_13379,N_13151);
nor U13607 (N_13607,N_13480,N_13338);
nand U13608 (N_13608,N_13258,N_13396);
xnor U13609 (N_13609,N_13415,N_13205);
nand U13610 (N_13610,N_13274,N_13409);
nand U13611 (N_13611,N_13427,N_13425);
xnor U13612 (N_13612,N_13294,N_13011);
nor U13613 (N_13613,N_13376,N_13224);
nor U13614 (N_13614,N_13080,N_13232);
or U13615 (N_13615,N_13319,N_13039);
nand U13616 (N_13616,N_13450,N_13293);
nand U13617 (N_13617,N_13118,N_13328);
or U13618 (N_13618,N_13211,N_13045);
or U13619 (N_13619,N_13252,N_13227);
xnor U13620 (N_13620,N_13106,N_13407);
nor U13621 (N_13621,N_13253,N_13391);
and U13622 (N_13622,N_13221,N_13213);
nor U13623 (N_13623,N_13203,N_13136);
nand U13624 (N_13624,N_13059,N_13410);
or U13625 (N_13625,N_13175,N_13127);
and U13626 (N_13626,N_13057,N_13451);
nand U13627 (N_13627,N_13085,N_13445);
nor U13628 (N_13628,N_13417,N_13150);
xnor U13629 (N_13629,N_13329,N_13402);
nor U13630 (N_13630,N_13051,N_13113);
nor U13631 (N_13631,N_13003,N_13082);
and U13632 (N_13632,N_13322,N_13194);
or U13633 (N_13633,N_13078,N_13006);
nor U13634 (N_13634,N_13473,N_13168);
or U13635 (N_13635,N_13334,N_13133);
nor U13636 (N_13636,N_13423,N_13098);
and U13637 (N_13637,N_13162,N_13303);
nand U13638 (N_13638,N_13095,N_13295);
nand U13639 (N_13639,N_13448,N_13128);
nand U13640 (N_13640,N_13325,N_13200);
or U13641 (N_13641,N_13132,N_13389);
and U13642 (N_13642,N_13240,N_13371);
nand U13643 (N_13643,N_13092,N_13038);
nor U13644 (N_13644,N_13035,N_13043);
nand U13645 (N_13645,N_13377,N_13302);
xnor U13646 (N_13646,N_13471,N_13479);
and U13647 (N_13647,N_13297,N_13185);
and U13648 (N_13648,N_13110,N_13123);
or U13649 (N_13649,N_13467,N_13416);
or U13650 (N_13650,N_13056,N_13284);
nor U13651 (N_13651,N_13197,N_13490);
nand U13652 (N_13652,N_13256,N_13443);
or U13653 (N_13653,N_13310,N_13172);
nand U13654 (N_13654,N_13494,N_13184);
nor U13655 (N_13655,N_13242,N_13419);
nor U13656 (N_13656,N_13424,N_13088);
xnor U13657 (N_13657,N_13193,N_13323);
nor U13658 (N_13658,N_13187,N_13236);
and U13659 (N_13659,N_13130,N_13444);
or U13660 (N_13660,N_13093,N_13228);
nand U13661 (N_13661,N_13421,N_13255);
or U13662 (N_13662,N_13070,N_13207);
nor U13663 (N_13663,N_13245,N_13041);
or U13664 (N_13664,N_13370,N_13154);
or U13665 (N_13665,N_13432,N_13171);
and U13666 (N_13666,N_13247,N_13148);
nor U13667 (N_13667,N_13404,N_13137);
or U13668 (N_13668,N_13068,N_13142);
or U13669 (N_13669,N_13196,N_13246);
and U13670 (N_13670,N_13179,N_13361);
nand U13671 (N_13671,N_13000,N_13254);
nand U13672 (N_13672,N_13216,N_13487);
xor U13673 (N_13673,N_13496,N_13244);
and U13674 (N_13674,N_13155,N_13308);
and U13675 (N_13675,N_13183,N_13291);
nand U13676 (N_13676,N_13381,N_13260);
nand U13677 (N_13677,N_13288,N_13198);
and U13678 (N_13678,N_13368,N_13300);
xor U13679 (N_13679,N_13365,N_13320);
or U13680 (N_13680,N_13273,N_13277);
and U13681 (N_13681,N_13460,N_13237);
xnor U13682 (N_13682,N_13287,N_13219);
and U13683 (N_13683,N_13299,N_13140);
xnor U13684 (N_13684,N_13040,N_13212);
nand U13685 (N_13685,N_13065,N_13298);
xnor U13686 (N_13686,N_13493,N_13249);
nor U13687 (N_13687,N_13382,N_13138);
nor U13688 (N_13688,N_13046,N_13033);
nand U13689 (N_13689,N_13296,N_13403);
nand U13690 (N_13690,N_13269,N_13161);
or U13691 (N_13691,N_13484,N_13129);
and U13692 (N_13692,N_13170,N_13353);
and U13693 (N_13693,N_13145,N_13332);
nor U13694 (N_13694,N_13061,N_13406);
nand U13695 (N_13695,N_13290,N_13218);
nand U13696 (N_13696,N_13313,N_13355);
and U13697 (N_13697,N_13181,N_13251);
or U13698 (N_13698,N_13028,N_13446);
or U13699 (N_13699,N_13305,N_13397);
and U13700 (N_13700,N_13312,N_13380);
and U13701 (N_13701,N_13400,N_13357);
nor U13702 (N_13702,N_13453,N_13021);
or U13703 (N_13703,N_13094,N_13173);
xnor U13704 (N_13704,N_13117,N_13440);
and U13705 (N_13705,N_13316,N_13131);
xor U13706 (N_13706,N_13359,N_13201);
or U13707 (N_13707,N_13054,N_13315);
nor U13708 (N_13708,N_13429,N_13478);
or U13709 (N_13709,N_13188,N_13388);
nand U13710 (N_13710,N_13047,N_13108);
nand U13711 (N_13711,N_13262,N_13195);
or U13712 (N_13712,N_13463,N_13231);
or U13713 (N_13713,N_13321,N_13477);
nand U13714 (N_13714,N_13352,N_13399);
xor U13715 (N_13715,N_13191,N_13102);
or U13716 (N_13716,N_13177,N_13053);
nand U13717 (N_13717,N_13190,N_13449);
or U13718 (N_13718,N_13362,N_13165);
nor U13719 (N_13719,N_13326,N_13015);
nand U13720 (N_13720,N_13491,N_13307);
xor U13721 (N_13721,N_13366,N_13159);
and U13722 (N_13722,N_13243,N_13166);
nor U13723 (N_13723,N_13126,N_13087);
and U13724 (N_13724,N_13470,N_13174);
xor U13725 (N_13725,N_13459,N_13058);
and U13726 (N_13726,N_13149,N_13233);
and U13727 (N_13727,N_13418,N_13241);
and U13728 (N_13728,N_13265,N_13283);
or U13729 (N_13729,N_13121,N_13405);
xor U13730 (N_13730,N_13107,N_13351);
xnor U13731 (N_13731,N_13063,N_13461);
nand U13732 (N_13732,N_13436,N_13430);
nor U13733 (N_13733,N_13141,N_13433);
xor U13734 (N_13734,N_13489,N_13125);
xor U13735 (N_13735,N_13152,N_13324);
or U13736 (N_13736,N_13263,N_13069);
nand U13737 (N_13737,N_13408,N_13395);
and U13738 (N_13738,N_13482,N_13189);
and U13739 (N_13739,N_13157,N_13447);
xnor U13740 (N_13740,N_13369,N_13385);
nand U13741 (N_13741,N_13474,N_13340);
or U13742 (N_13742,N_13499,N_13390);
xnor U13743 (N_13743,N_13146,N_13112);
xor U13744 (N_13744,N_13412,N_13281);
xor U13745 (N_13745,N_13337,N_13025);
or U13746 (N_13746,N_13317,N_13393);
nor U13747 (N_13747,N_13267,N_13101);
nand U13748 (N_13748,N_13268,N_13248);
xnor U13749 (N_13749,N_13422,N_13458);
nand U13750 (N_13750,N_13304,N_13422);
and U13751 (N_13751,N_13492,N_13186);
xnor U13752 (N_13752,N_13482,N_13337);
xnor U13753 (N_13753,N_13048,N_13348);
or U13754 (N_13754,N_13325,N_13017);
xnor U13755 (N_13755,N_13003,N_13341);
nor U13756 (N_13756,N_13375,N_13395);
nor U13757 (N_13757,N_13281,N_13269);
xnor U13758 (N_13758,N_13453,N_13263);
or U13759 (N_13759,N_13329,N_13462);
nand U13760 (N_13760,N_13227,N_13005);
nor U13761 (N_13761,N_13143,N_13260);
nor U13762 (N_13762,N_13365,N_13162);
xnor U13763 (N_13763,N_13359,N_13335);
nor U13764 (N_13764,N_13149,N_13103);
nand U13765 (N_13765,N_13216,N_13058);
nor U13766 (N_13766,N_13027,N_13252);
nor U13767 (N_13767,N_13072,N_13410);
nand U13768 (N_13768,N_13407,N_13217);
xnor U13769 (N_13769,N_13289,N_13495);
xor U13770 (N_13770,N_13289,N_13186);
or U13771 (N_13771,N_13368,N_13288);
xnor U13772 (N_13772,N_13455,N_13399);
or U13773 (N_13773,N_13318,N_13312);
xnor U13774 (N_13774,N_13495,N_13305);
nand U13775 (N_13775,N_13417,N_13405);
nor U13776 (N_13776,N_13295,N_13128);
nand U13777 (N_13777,N_13298,N_13281);
xor U13778 (N_13778,N_13221,N_13055);
and U13779 (N_13779,N_13269,N_13319);
nor U13780 (N_13780,N_13329,N_13178);
or U13781 (N_13781,N_13221,N_13448);
nand U13782 (N_13782,N_13264,N_13269);
xnor U13783 (N_13783,N_13295,N_13371);
nand U13784 (N_13784,N_13169,N_13226);
xor U13785 (N_13785,N_13490,N_13035);
or U13786 (N_13786,N_13402,N_13326);
or U13787 (N_13787,N_13081,N_13082);
xnor U13788 (N_13788,N_13218,N_13274);
nor U13789 (N_13789,N_13110,N_13269);
or U13790 (N_13790,N_13031,N_13337);
or U13791 (N_13791,N_13455,N_13427);
nand U13792 (N_13792,N_13243,N_13104);
nand U13793 (N_13793,N_13352,N_13424);
or U13794 (N_13794,N_13020,N_13143);
nand U13795 (N_13795,N_13399,N_13437);
or U13796 (N_13796,N_13143,N_13067);
xnor U13797 (N_13797,N_13269,N_13365);
xor U13798 (N_13798,N_13037,N_13051);
nor U13799 (N_13799,N_13132,N_13279);
nor U13800 (N_13800,N_13420,N_13170);
nand U13801 (N_13801,N_13290,N_13485);
and U13802 (N_13802,N_13185,N_13415);
or U13803 (N_13803,N_13038,N_13387);
nand U13804 (N_13804,N_13473,N_13326);
and U13805 (N_13805,N_13023,N_13432);
nand U13806 (N_13806,N_13248,N_13036);
nand U13807 (N_13807,N_13052,N_13326);
and U13808 (N_13808,N_13422,N_13329);
nor U13809 (N_13809,N_13315,N_13162);
or U13810 (N_13810,N_13175,N_13341);
xor U13811 (N_13811,N_13150,N_13115);
nand U13812 (N_13812,N_13190,N_13396);
xnor U13813 (N_13813,N_13163,N_13337);
nor U13814 (N_13814,N_13339,N_13257);
nand U13815 (N_13815,N_13058,N_13404);
and U13816 (N_13816,N_13027,N_13412);
xor U13817 (N_13817,N_13147,N_13427);
nand U13818 (N_13818,N_13018,N_13326);
or U13819 (N_13819,N_13040,N_13339);
xnor U13820 (N_13820,N_13186,N_13392);
nor U13821 (N_13821,N_13471,N_13089);
xnor U13822 (N_13822,N_13061,N_13246);
xnor U13823 (N_13823,N_13071,N_13259);
nand U13824 (N_13824,N_13291,N_13436);
nand U13825 (N_13825,N_13476,N_13490);
xor U13826 (N_13826,N_13163,N_13327);
nor U13827 (N_13827,N_13147,N_13408);
nand U13828 (N_13828,N_13187,N_13327);
nand U13829 (N_13829,N_13220,N_13234);
nand U13830 (N_13830,N_13020,N_13182);
or U13831 (N_13831,N_13263,N_13140);
or U13832 (N_13832,N_13120,N_13443);
nand U13833 (N_13833,N_13020,N_13337);
xor U13834 (N_13834,N_13022,N_13318);
nand U13835 (N_13835,N_13118,N_13243);
and U13836 (N_13836,N_13419,N_13480);
and U13837 (N_13837,N_13170,N_13468);
nand U13838 (N_13838,N_13137,N_13370);
nand U13839 (N_13839,N_13314,N_13451);
nor U13840 (N_13840,N_13223,N_13266);
nand U13841 (N_13841,N_13349,N_13023);
nor U13842 (N_13842,N_13047,N_13288);
nor U13843 (N_13843,N_13387,N_13174);
nor U13844 (N_13844,N_13030,N_13043);
xor U13845 (N_13845,N_13272,N_13153);
and U13846 (N_13846,N_13003,N_13456);
nor U13847 (N_13847,N_13281,N_13138);
and U13848 (N_13848,N_13453,N_13159);
nand U13849 (N_13849,N_13005,N_13439);
or U13850 (N_13850,N_13238,N_13409);
or U13851 (N_13851,N_13416,N_13228);
nand U13852 (N_13852,N_13173,N_13379);
and U13853 (N_13853,N_13415,N_13332);
or U13854 (N_13854,N_13459,N_13122);
xnor U13855 (N_13855,N_13343,N_13159);
or U13856 (N_13856,N_13288,N_13314);
nor U13857 (N_13857,N_13393,N_13009);
nor U13858 (N_13858,N_13417,N_13096);
xor U13859 (N_13859,N_13405,N_13425);
nor U13860 (N_13860,N_13042,N_13255);
and U13861 (N_13861,N_13375,N_13436);
and U13862 (N_13862,N_13291,N_13099);
nand U13863 (N_13863,N_13092,N_13185);
xnor U13864 (N_13864,N_13301,N_13210);
or U13865 (N_13865,N_13147,N_13086);
nor U13866 (N_13866,N_13115,N_13315);
xnor U13867 (N_13867,N_13471,N_13328);
and U13868 (N_13868,N_13228,N_13477);
xor U13869 (N_13869,N_13486,N_13303);
or U13870 (N_13870,N_13208,N_13345);
or U13871 (N_13871,N_13055,N_13110);
and U13872 (N_13872,N_13308,N_13175);
and U13873 (N_13873,N_13037,N_13136);
xnor U13874 (N_13874,N_13273,N_13353);
nand U13875 (N_13875,N_13022,N_13198);
or U13876 (N_13876,N_13425,N_13397);
nand U13877 (N_13877,N_13411,N_13337);
and U13878 (N_13878,N_13103,N_13359);
xnor U13879 (N_13879,N_13401,N_13150);
nor U13880 (N_13880,N_13074,N_13232);
and U13881 (N_13881,N_13131,N_13102);
and U13882 (N_13882,N_13449,N_13486);
xor U13883 (N_13883,N_13207,N_13468);
or U13884 (N_13884,N_13474,N_13397);
and U13885 (N_13885,N_13231,N_13222);
xor U13886 (N_13886,N_13022,N_13028);
xor U13887 (N_13887,N_13092,N_13210);
nand U13888 (N_13888,N_13264,N_13196);
nand U13889 (N_13889,N_13459,N_13108);
nand U13890 (N_13890,N_13071,N_13007);
or U13891 (N_13891,N_13275,N_13262);
nand U13892 (N_13892,N_13364,N_13293);
nor U13893 (N_13893,N_13118,N_13482);
and U13894 (N_13894,N_13495,N_13439);
and U13895 (N_13895,N_13477,N_13347);
nand U13896 (N_13896,N_13470,N_13319);
and U13897 (N_13897,N_13215,N_13053);
xor U13898 (N_13898,N_13000,N_13329);
or U13899 (N_13899,N_13348,N_13447);
and U13900 (N_13900,N_13316,N_13407);
and U13901 (N_13901,N_13346,N_13189);
xnor U13902 (N_13902,N_13389,N_13260);
and U13903 (N_13903,N_13421,N_13493);
nand U13904 (N_13904,N_13071,N_13106);
nand U13905 (N_13905,N_13300,N_13320);
xor U13906 (N_13906,N_13074,N_13077);
and U13907 (N_13907,N_13235,N_13107);
or U13908 (N_13908,N_13283,N_13267);
and U13909 (N_13909,N_13089,N_13211);
or U13910 (N_13910,N_13419,N_13307);
nor U13911 (N_13911,N_13112,N_13306);
nand U13912 (N_13912,N_13122,N_13460);
or U13913 (N_13913,N_13314,N_13473);
xor U13914 (N_13914,N_13140,N_13439);
nor U13915 (N_13915,N_13424,N_13356);
or U13916 (N_13916,N_13444,N_13020);
nand U13917 (N_13917,N_13016,N_13448);
nor U13918 (N_13918,N_13482,N_13285);
xnor U13919 (N_13919,N_13260,N_13302);
xor U13920 (N_13920,N_13116,N_13151);
and U13921 (N_13921,N_13342,N_13001);
nor U13922 (N_13922,N_13425,N_13102);
xnor U13923 (N_13923,N_13047,N_13129);
nor U13924 (N_13924,N_13201,N_13409);
nor U13925 (N_13925,N_13083,N_13487);
nor U13926 (N_13926,N_13430,N_13187);
nand U13927 (N_13927,N_13275,N_13406);
or U13928 (N_13928,N_13429,N_13381);
and U13929 (N_13929,N_13130,N_13478);
and U13930 (N_13930,N_13190,N_13180);
or U13931 (N_13931,N_13203,N_13228);
xor U13932 (N_13932,N_13032,N_13271);
or U13933 (N_13933,N_13022,N_13494);
nand U13934 (N_13934,N_13067,N_13073);
xor U13935 (N_13935,N_13000,N_13017);
nand U13936 (N_13936,N_13327,N_13343);
nand U13937 (N_13937,N_13458,N_13061);
or U13938 (N_13938,N_13125,N_13353);
nand U13939 (N_13939,N_13477,N_13216);
nor U13940 (N_13940,N_13359,N_13186);
or U13941 (N_13941,N_13052,N_13285);
or U13942 (N_13942,N_13384,N_13448);
nor U13943 (N_13943,N_13451,N_13267);
nor U13944 (N_13944,N_13175,N_13037);
and U13945 (N_13945,N_13420,N_13325);
xnor U13946 (N_13946,N_13303,N_13200);
or U13947 (N_13947,N_13348,N_13003);
nor U13948 (N_13948,N_13258,N_13002);
or U13949 (N_13949,N_13016,N_13458);
nand U13950 (N_13950,N_13222,N_13319);
nor U13951 (N_13951,N_13195,N_13023);
xnor U13952 (N_13952,N_13138,N_13424);
nor U13953 (N_13953,N_13211,N_13279);
xor U13954 (N_13954,N_13481,N_13159);
nand U13955 (N_13955,N_13437,N_13239);
and U13956 (N_13956,N_13435,N_13299);
nand U13957 (N_13957,N_13451,N_13365);
and U13958 (N_13958,N_13272,N_13427);
and U13959 (N_13959,N_13156,N_13228);
and U13960 (N_13960,N_13118,N_13466);
xor U13961 (N_13961,N_13295,N_13179);
nand U13962 (N_13962,N_13278,N_13112);
nor U13963 (N_13963,N_13154,N_13342);
and U13964 (N_13964,N_13220,N_13377);
or U13965 (N_13965,N_13011,N_13248);
xor U13966 (N_13966,N_13281,N_13146);
and U13967 (N_13967,N_13181,N_13065);
and U13968 (N_13968,N_13397,N_13073);
and U13969 (N_13969,N_13376,N_13214);
nor U13970 (N_13970,N_13490,N_13125);
or U13971 (N_13971,N_13113,N_13056);
xnor U13972 (N_13972,N_13236,N_13265);
nor U13973 (N_13973,N_13164,N_13480);
nor U13974 (N_13974,N_13187,N_13015);
xnor U13975 (N_13975,N_13414,N_13393);
nand U13976 (N_13976,N_13150,N_13078);
nor U13977 (N_13977,N_13096,N_13489);
nor U13978 (N_13978,N_13146,N_13150);
and U13979 (N_13979,N_13387,N_13498);
nand U13980 (N_13980,N_13196,N_13223);
and U13981 (N_13981,N_13450,N_13029);
and U13982 (N_13982,N_13010,N_13464);
nand U13983 (N_13983,N_13377,N_13042);
or U13984 (N_13984,N_13413,N_13166);
and U13985 (N_13985,N_13381,N_13152);
nor U13986 (N_13986,N_13431,N_13050);
xnor U13987 (N_13987,N_13204,N_13408);
or U13988 (N_13988,N_13496,N_13485);
xor U13989 (N_13989,N_13210,N_13299);
nand U13990 (N_13990,N_13236,N_13417);
nor U13991 (N_13991,N_13090,N_13067);
nor U13992 (N_13992,N_13374,N_13235);
and U13993 (N_13993,N_13181,N_13341);
xor U13994 (N_13994,N_13162,N_13469);
xnor U13995 (N_13995,N_13115,N_13269);
or U13996 (N_13996,N_13401,N_13327);
nor U13997 (N_13997,N_13371,N_13030);
nand U13998 (N_13998,N_13394,N_13348);
or U13999 (N_13999,N_13470,N_13152);
or U14000 (N_14000,N_13699,N_13513);
and U14001 (N_14001,N_13773,N_13539);
or U14002 (N_14002,N_13662,N_13534);
xnor U14003 (N_14003,N_13988,N_13587);
and U14004 (N_14004,N_13922,N_13613);
and U14005 (N_14005,N_13728,N_13933);
or U14006 (N_14006,N_13678,N_13734);
nand U14007 (N_14007,N_13574,N_13865);
xnor U14008 (N_14008,N_13564,N_13704);
nand U14009 (N_14009,N_13626,N_13677);
and U14010 (N_14010,N_13900,N_13603);
nor U14011 (N_14011,N_13731,N_13670);
or U14012 (N_14012,N_13596,N_13952);
nor U14013 (N_14013,N_13751,N_13632);
xnor U14014 (N_14014,N_13785,N_13909);
nand U14015 (N_14015,N_13913,N_13762);
xnor U14016 (N_14016,N_13690,N_13759);
xnor U14017 (N_14017,N_13761,N_13580);
or U14018 (N_14018,N_13606,N_13554);
or U14019 (N_14019,N_13683,N_13710);
nor U14020 (N_14020,N_13857,N_13852);
or U14021 (N_14021,N_13671,N_13996);
and U14022 (N_14022,N_13843,N_13904);
xor U14023 (N_14023,N_13879,N_13732);
or U14024 (N_14024,N_13873,N_13923);
or U14025 (N_14025,N_13726,N_13625);
and U14026 (N_14026,N_13541,N_13559);
nand U14027 (N_14027,N_13660,N_13514);
or U14028 (N_14028,N_13977,N_13902);
xor U14029 (N_14029,N_13543,N_13911);
xor U14030 (N_14030,N_13816,N_13803);
xnor U14031 (N_14031,N_13984,N_13552);
nor U14032 (N_14032,N_13818,N_13739);
or U14033 (N_14033,N_13951,N_13948);
nand U14034 (N_14034,N_13727,N_13793);
or U14035 (N_14035,N_13569,N_13832);
nand U14036 (N_14036,N_13730,N_13782);
xor U14037 (N_14037,N_13932,N_13776);
or U14038 (N_14038,N_13939,N_13797);
nor U14039 (N_14039,N_13975,N_13535);
nand U14040 (N_14040,N_13839,N_13525);
or U14041 (N_14041,N_13508,N_13691);
or U14042 (N_14042,N_13860,N_13805);
xnor U14043 (N_14043,N_13877,N_13510);
xor U14044 (N_14044,N_13589,N_13602);
or U14045 (N_14045,N_13848,N_13504);
or U14046 (N_14046,N_13601,N_13550);
nor U14047 (N_14047,N_13791,N_13636);
nor U14048 (N_14048,N_13743,N_13693);
nand U14049 (N_14049,N_13694,N_13612);
nor U14050 (N_14050,N_13910,N_13680);
or U14051 (N_14051,N_13701,N_13876);
xnor U14052 (N_14052,N_13674,N_13740);
xnor U14053 (N_14053,N_13545,N_13868);
or U14054 (N_14054,N_13511,N_13649);
nand U14055 (N_14055,N_13597,N_13944);
nand U14056 (N_14056,N_13755,N_13926);
xnor U14057 (N_14057,N_13611,N_13970);
nand U14058 (N_14058,N_13706,N_13972);
xnor U14059 (N_14059,N_13795,N_13924);
and U14060 (N_14060,N_13617,N_13815);
nor U14061 (N_14061,N_13528,N_13658);
and U14062 (N_14062,N_13682,N_13708);
and U14063 (N_14063,N_13769,N_13647);
xor U14064 (N_14064,N_13886,N_13746);
and U14065 (N_14065,N_13512,N_13960);
nand U14066 (N_14066,N_13973,N_13692);
and U14067 (N_14067,N_13789,N_13982);
nand U14068 (N_14068,N_13507,N_13990);
nand U14069 (N_14069,N_13527,N_13925);
xor U14070 (N_14070,N_13827,N_13506);
or U14071 (N_14071,N_13542,N_13723);
nand U14072 (N_14072,N_13711,N_13563);
nand U14073 (N_14073,N_13936,N_13661);
xnor U14074 (N_14074,N_13778,N_13771);
and U14075 (N_14075,N_13631,N_13872);
nand U14076 (N_14076,N_13808,N_13917);
xnor U14077 (N_14077,N_13942,N_13969);
or U14078 (N_14078,N_13903,N_13515);
nand U14079 (N_14079,N_13830,N_13600);
and U14080 (N_14080,N_13599,N_13666);
or U14081 (N_14081,N_13798,N_13834);
xnor U14082 (N_14082,N_13548,N_13918);
or U14083 (N_14083,N_13919,N_13958);
xor U14084 (N_14084,N_13891,N_13814);
nand U14085 (N_14085,N_13657,N_13572);
or U14086 (N_14086,N_13801,N_13651);
nand U14087 (N_14087,N_13754,N_13573);
or U14088 (N_14088,N_13985,N_13520);
xor U14089 (N_14089,N_13591,N_13757);
nand U14090 (N_14090,N_13595,N_13957);
or U14091 (N_14091,N_13862,N_13709);
nand U14092 (N_14092,N_13800,N_13875);
nor U14093 (N_14093,N_13817,N_13640);
or U14094 (N_14094,N_13863,N_13607);
nor U14095 (N_14095,N_13522,N_13689);
nor U14096 (N_14096,N_13796,N_13654);
nor U14097 (N_14097,N_13532,N_13828);
and U14098 (N_14098,N_13652,N_13979);
and U14099 (N_14099,N_13943,N_13623);
or U14100 (N_14100,N_13745,N_13570);
xnor U14101 (N_14101,N_13887,N_13837);
xor U14102 (N_14102,N_13859,N_13737);
nor U14103 (N_14103,N_13538,N_13581);
or U14104 (N_14104,N_13655,N_13976);
nor U14105 (N_14105,N_13802,N_13838);
and U14106 (N_14106,N_13729,N_13788);
xor U14107 (N_14107,N_13669,N_13653);
nand U14108 (N_14108,N_13850,N_13955);
or U14109 (N_14109,N_13518,N_13790);
nor U14110 (N_14110,N_13588,N_13779);
nand U14111 (N_14111,N_13610,N_13676);
xor U14112 (N_14112,N_13836,N_13864);
or U14113 (N_14113,N_13594,N_13644);
nand U14114 (N_14114,N_13722,N_13811);
nor U14115 (N_14115,N_13561,N_13686);
nand U14116 (N_14116,N_13978,N_13786);
nand U14117 (N_14117,N_13540,N_13920);
or U14118 (N_14118,N_13664,N_13768);
or U14119 (N_14119,N_13861,N_13735);
nand U14120 (N_14120,N_13592,N_13703);
nand U14121 (N_14121,N_13697,N_13738);
and U14122 (N_14122,N_13530,N_13568);
and U14123 (N_14123,N_13974,N_13983);
or U14124 (N_14124,N_13893,N_13713);
and U14125 (N_14125,N_13643,N_13878);
xor U14126 (N_14126,N_13645,N_13914);
and U14127 (N_14127,N_13787,N_13945);
nor U14128 (N_14128,N_13831,N_13899);
nor U14129 (N_14129,N_13823,N_13698);
xor U14130 (N_14130,N_13609,N_13712);
xor U14131 (N_14131,N_13720,N_13915);
nand U14132 (N_14132,N_13668,N_13966);
nor U14133 (N_14133,N_13935,N_13560);
xor U14134 (N_14134,N_13721,N_13533);
nor U14135 (N_14135,N_13883,N_13557);
nand U14136 (N_14136,N_13696,N_13956);
or U14137 (N_14137,N_13847,N_13810);
or U14138 (N_14138,N_13824,N_13665);
xnor U14139 (N_14139,N_13896,N_13517);
nand U14140 (N_14140,N_13963,N_13908);
xnor U14141 (N_14141,N_13889,N_13667);
xor U14142 (N_14142,N_13705,N_13833);
nand U14143 (N_14143,N_13844,N_13566);
nor U14144 (N_14144,N_13871,N_13736);
nor U14145 (N_14145,N_13965,N_13562);
xor U14146 (N_14146,N_13585,N_13584);
nand U14147 (N_14147,N_13916,N_13715);
and U14148 (N_14148,N_13905,N_13894);
or U14149 (N_14149,N_13509,N_13981);
xor U14150 (N_14150,N_13901,N_13890);
or U14151 (N_14151,N_13760,N_13961);
nand U14152 (N_14152,N_13544,N_13546);
nand U14153 (N_14153,N_13885,N_13576);
and U14154 (N_14154,N_13930,N_13880);
nor U14155 (N_14155,N_13579,N_13741);
and U14156 (N_14156,N_13764,N_13502);
and U14157 (N_14157,N_13641,N_13679);
and U14158 (N_14158,N_13639,N_13853);
xor U14159 (N_14159,N_13971,N_13804);
or U14160 (N_14160,N_13964,N_13633);
nor U14161 (N_14161,N_13571,N_13770);
and U14162 (N_14162,N_13551,N_13884);
nor U14163 (N_14163,N_13794,N_13888);
nand U14164 (N_14164,N_13567,N_13642);
and U14165 (N_14165,N_13986,N_13772);
or U14166 (N_14166,N_13650,N_13851);
nor U14167 (N_14167,N_13687,N_13822);
nor U14168 (N_14168,N_13744,N_13912);
nand U14169 (N_14169,N_13558,N_13813);
and U14170 (N_14170,N_13947,N_13583);
and U14171 (N_14171,N_13577,N_13842);
nand U14172 (N_14172,N_13934,N_13637);
and U14173 (N_14173,N_13582,N_13999);
xnor U14174 (N_14174,N_13684,N_13598);
nand U14175 (N_14175,N_13608,N_13941);
xnor U14176 (N_14176,N_13840,N_13898);
or U14177 (N_14177,N_13749,N_13774);
nand U14178 (N_14178,N_13688,N_13892);
xor U14179 (N_14179,N_13987,N_13619);
nor U14180 (N_14180,N_13624,N_13663);
nand U14181 (N_14181,N_13531,N_13807);
xnor U14182 (N_14182,N_13718,N_13565);
xnor U14183 (N_14183,N_13767,N_13881);
or U14184 (N_14184,N_13505,N_13781);
and U14185 (N_14185,N_13656,N_13950);
or U14186 (N_14186,N_13556,N_13784);
or U14187 (N_14187,N_13503,N_13618);
or U14188 (N_14188,N_13766,N_13742);
xnor U14189 (N_14189,N_13959,N_13821);
and U14190 (N_14190,N_13994,N_13590);
xor U14191 (N_14191,N_13681,N_13825);
xnor U14192 (N_14192,N_13792,N_13938);
xor U14193 (N_14193,N_13700,N_13748);
xor U14194 (N_14194,N_13616,N_13858);
xor U14195 (N_14195,N_13995,N_13841);
nor U14196 (N_14196,N_13758,N_13622);
and U14197 (N_14197,N_13869,N_13967);
xor U14198 (N_14198,N_13635,N_13605);
nand U14199 (N_14199,N_13829,N_13929);
xor U14200 (N_14200,N_13968,N_13549);
nor U14201 (N_14201,N_13954,N_13991);
nor U14202 (N_14202,N_13946,N_13646);
or U14203 (N_14203,N_13989,N_13500);
nor U14204 (N_14204,N_13849,N_13707);
nand U14205 (N_14205,N_13940,N_13586);
nor U14206 (N_14206,N_13675,N_13621);
and U14207 (N_14207,N_13702,N_13553);
nand U14208 (N_14208,N_13536,N_13716);
nand U14209 (N_14209,N_13529,N_13928);
or U14210 (N_14210,N_13614,N_13931);
nand U14211 (N_14211,N_13799,N_13882);
nor U14212 (N_14212,N_13783,N_13523);
nand U14213 (N_14213,N_13714,N_13980);
xor U14214 (N_14214,N_13866,N_13906);
nor U14215 (N_14215,N_13685,N_13673);
nor U14216 (N_14216,N_13993,N_13672);
xnor U14217 (N_14217,N_13780,N_13725);
and U14218 (N_14218,N_13519,N_13765);
or U14219 (N_14219,N_13820,N_13845);
nand U14220 (N_14220,N_13921,N_13907);
and U14221 (N_14221,N_13620,N_13547);
nand U14222 (N_14222,N_13937,N_13638);
or U14223 (N_14223,N_13809,N_13719);
or U14224 (N_14224,N_13634,N_13752);
nand U14225 (N_14225,N_13695,N_13927);
and U14226 (N_14226,N_13724,N_13593);
xnor U14227 (N_14227,N_13867,N_13998);
nor U14228 (N_14228,N_13575,N_13775);
nor U14229 (N_14229,N_13854,N_13750);
or U14230 (N_14230,N_13897,N_13870);
nand U14231 (N_14231,N_13953,N_13846);
or U14232 (N_14232,N_13997,N_13615);
or U14233 (N_14233,N_13524,N_13537);
and U14234 (N_14234,N_13501,N_13874);
nor U14235 (N_14235,N_13753,N_13962);
nor U14236 (N_14236,N_13604,N_13763);
xor U14237 (N_14237,N_13578,N_13648);
or U14238 (N_14238,N_13806,N_13992);
and U14239 (N_14239,N_13521,N_13895);
nor U14240 (N_14240,N_13555,N_13628);
and U14241 (N_14241,N_13717,N_13526);
or U14242 (N_14242,N_13630,N_13856);
nor U14243 (N_14243,N_13756,N_13855);
nand U14244 (N_14244,N_13747,N_13819);
nand U14245 (N_14245,N_13627,N_13629);
or U14246 (N_14246,N_13516,N_13949);
and U14247 (N_14247,N_13659,N_13777);
nor U14248 (N_14248,N_13835,N_13826);
or U14249 (N_14249,N_13733,N_13812);
xor U14250 (N_14250,N_13782,N_13688);
xor U14251 (N_14251,N_13773,N_13542);
nor U14252 (N_14252,N_13768,N_13833);
nor U14253 (N_14253,N_13845,N_13988);
nand U14254 (N_14254,N_13655,N_13656);
xnor U14255 (N_14255,N_13548,N_13553);
nor U14256 (N_14256,N_13657,N_13937);
nor U14257 (N_14257,N_13695,N_13539);
or U14258 (N_14258,N_13665,N_13759);
xor U14259 (N_14259,N_13624,N_13636);
xnor U14260 (N_14260,N_13695,N_13769);
xor U14261 (N_14261,N_13846,N_13842);
nor U14262 (N_14262,N_13917,N_13981);
nand U14263 (N_14263,N_13669,N_13841);
nor U14264 (N_14264,N_13683,N_13908);
xor U14265 (N_14265,N_13740,N_13911);
and U14266 (N_14266,N_13670,N_13895);
or U14267 (N_14267,N_13820,N_13824);
nor U14268 (N_14268,N_13776,N_13552);
or U14269 (N_14269,N_13870,N_13786);
and U14270 (N_14270,N_13892,N_13647);
nor U14271 (N_14271,N_13755,N_13748);
nor U14272 (N_14272,N_13928,N_13707);
or U14273 (N_14273,N_13881,N_13989);
nor U14274 (N_14274,N_13776,N_13943);
or U14275 (N_14275,N_13506,N_13861);
and U14276 (N_14276,N_13568,N_13563);
nor U14277 (N_14277,N_13865,N_13890);
nor U14278 (N_14278,N_13563,N_13616);
nand U14279 (N_14279,N_13903,N_13519);
xnor U14280 (N_14280,N_13507,N_13599);
and U14281 (N_14281,N_13797,N_13564);
and U14282 (N_14282,N_13516,N_13751);
nor U14283 (N_14283,N_13672,N_13847);
nand U14284 (N_14284,N_13581,N_13940);
and U14285 (N_14285,N_13584,N_13670);
xnor U14286 (N_14286,N_13696,N_13661);
nor U14287 (N_14287,N_13570,N_13954);
xor U14288 (N_14288,N_13920,N_13677);
nand U14289 (N_14289,N_13643,N_13952);
or U14290 (N_14290,N_13988,N_13637);
nand U14291 (N_14291,N_13582,N_13671);
nand U14292 (N_14292,N_13987,N_13664);
and U14293 (N_14293,N_13669,N_13619);
nand U14294 (N_14294,N_13809,N_13799);
or U14295 (N_14295,N_13694,N_13902);
nand U14296 (N_14296,N_13898,N_13509);
or U14297 (N_14297,N_13501,N_13532);
nor U14298 (N_14298,N_13558,N_13737);
nand U14299 (N_14299,N_13556,N_13835);
nor U14300 (N_14300,N_13586,N_13995);
or U14301 (N_14301,N_13987,N_13830);
xnor U14302 (N_14302,N_13972,N_13618);
xnor U14303 (N_14303,N_13799,N_13600);
nor U14304 (N_14304,N_13970,N_13541);
nor U14305 (N_14305,N_13950,N_13667);
nor U14306 (N_14306,N_13644,N_13597);
and U14307 (N_14307,N_13963,N_13965);
nor U14308 (N_14308,N_13843,N_13933);
nor U14309 (N_14309,N_13617,N_13600);
nor U14310 (N_14310,N_13952,N_13966);
nand U14311 (N_14311,N_13991,N_13773);
xor U14312 (N_14312,N_13570,N_13654);
or U14313 (N_14313,N_13947,N_13620);
or U14314 (N_14314,N_13850,N_13602);
nor U14315 (N_14315,N_13662,N_13940);
nand U14316 (N_14316,N_13782,N_13898);
nand U14317 (N_14317,N_13507,N_13663);
nand U14318 (N_14318,N_13885,N_13785);
nand U14319 (N_14319,N_13587,N_13711);
nor U14320 (N_14320,N_13786,N_13921);
or U14321 (N_14321,N_13533,N_13909);
xnor U14322 (N_14322,N_13957,N_13945);
nor U14323 (N_14323,N_13662,N_13529);
nand U14324 (N_14324,N_13934,N_13658);
and U14325 (N_14325,N_13827,N_13772);
and U14326 (N_14326,N_13906,N_13993);
nand U14327 (N_14327,N_13815,N_13769);
xnor U14328 (N_14328,N_13792,N_13513);
or U14329 (N_14329,N_13524,N_13546);
xor U14330 (N_14330,N_13787,N_13747);
and U14331 (N_14331,N_13908,N_13614);
and U14332 (N_14332,N_13783,N_13713);
xor U14333 (N_14333,N_13901,N_13802);
and U14334 (N_14334,N_13823,N_13522);
and U14335 (N_14335,N_13987,N_13564);
or U14336 (N_14336,N_13661,N_13514);
nor U14337 (N_14337,N_13662,N_13584);
nor U14338 (N_14338,N_13787,N_13659);
nor U14339 (N_14339,N_13973,N_13543);
nor U14340 (N_14340,N_13878,N_13986);
or U14341 (N_14341,N_13567,N_13754);
and U14342 (N_14342,N_13909,N_13985);
or U14343 (N_14343,N_13829,N_13594);
nand U14344 (N_14344,N_13858,N_13694);
nor U14345 (N_14345,N_13925,N_13602);
nor U14346 (N_14346,N_13851,N_13994);
nand U14347 (N_14347,N_13577,N_13975);
or U14348 (N_14348,N_13931,N_13721);
nand U14349 (N_14349,N_13788,N_13807);
nand U14350 (N_14350,N_13674,N_13770);
nand U14351 (N_14351,N_13850,N_13590);
nand U14352 (N_14352,N_13857,N_13589);
nand U14353 (N_14353,N_13770,N_13860);
or U14354 (N_14354,N_13692,N_13739);
and U14355 (N_14355,N_13793,N_13798);
nor U14356 (N_14356,N_13613,N_13641);
nand U14357 (N_14357,N_13561,N_13763);
or U14358 (N_14358,N_13947,N_13910);
or U14359 (N_14359,N_13558,N_13506);
and U14360 (N_14360,N_13621,N_13770);
nor U14361 (N_14361,N_13582,N_13542);
nand U14362 (N_14362,N_13544,N_13849);
nand U14363 (N_14363,N_13644,N_13906);
nor U14364 (N_14364,N_13613,N_13778);
and U14365 (N_14365,N_13917,N_13525);
nor U14366 (N_14366,N_13864,N_13781);
or U14367 (N_14367,N_13736,N_13902);
nand U14368 (N_14368,N_13905,N_13556);
or U14369 (N_14369,N_13787,N_13662);
nor U14370 (N_14370,N_13531,N_13523);
xor U14371 (N_14371,N_13527,N_13988);
nand U14372 (N_14372,N_13814,N_13731);
and U14373 (N_14373,N_13901,N_13634);
or U14374 (N_14374,N_13606,N_13996);
and U14375 (N_14375,N_13863,N_13601);
nand U14376 (N_14376,N_13711,N_13863);
xnor U14377 (N_14377,N_13638,N_13920);
nor U14378 (N_14378,N_13961,N_13817);
nor U14379 (N_14379,N_13768,N_13841);
or U14380 (N_14380,N_13623,N_13885);
xnor U14381 (N_14381,N_13940,N_13816);
and U14382 (N_14382,N_13887,N_13521);
nor U14383 (N_14383,N_13515,N_13530);
and U14384 (N_14384,N_13730,N_13752);
xnor U14385 (N_14385,N_13599,N_13604);
nor U14386 (N_14386,N_13605,N_13766);
xor U14387 (N_14387,N_13978,N_13748);
nand U14388 (N_14388,N_13936,N_13786);
xnor U14389 (N_14389,N_13691,N_13827);
xnor U14390 (N_14390,N_13941,N_13736);
xor U14391 (N_14391,N_13582,N_13688);
xor U14392 (N_14392,N_13822,N_13522);
nand U14393 (N_14393,N_13625,N_13795);
nor U14394 (N_14394,N_13948,N_13688);
nor U14395 (N_14395,N_13913,N_13622);
or U14396 (N_14396,N_13873,N_13580);
nand U14397 (N_14397,N_13961,N_13861);
nand U14398 (N_14398,N_13588,N_13763);
nor U14399 (N_14399,N_13646,N_13694);
and U14400 (N_14400,N_13798,N_13501);
and U14401 (N_14401,N_13589,N_13966);
nor U14402 (N_14402,N_13914,N_13756);
and U14403 (N_14403,N_13977,N_13594);
nor U14404 (N_14404,N_13959,N_13644);
xnor U14405 (N_14405,N_13779,N_13925);
or U14406 (N_14406,N_13563,N_13837);
or U14407 (N_14407,N_13734,N_13928);
nor U14408 (N_14408,N_13704,N_13604);
and U14409 (N_14409,N_13997,N_13632);
nor U14410 (N_14410,N_13892,N_13880);
and U14411 (N_14411,N_13736,N_13732);
nand U14412 (N_14412,N_13931,N_13681);
nor U14413 (N_14413,N_13670,N_13503);
nor U14414 (N_14414,N_13565,N_13599);
nand U14415 (N_14415,N_13676,N_13707);
xor U14416 (N_14416,N_13690,N_13763);
xor U14417 (N_14417,N_13974,N_13867);
or U14418 (N_14418,N_13792,N_13637);
nor U14419 (N_14419,N_13627,N_13967);
or U14420 (N_14420,N_13639,N_13641);
and U14421 (N_14421,N_13907,N_13559);
or U14422 (N_14422,N_13528,N_13992);
and U14423 (N_14423,N_13530,N_13725);
nor U14424 (N_14424,N_13839,N_13732);
xor U14425 (N_14425,N_13951,N_13910);
nor U14426 (N_14426,N_13832,N_13717);
nand U14427 (N_14427,N_13788,N_13600);
nor U14428 (N_14428,N_13790,N_13535);
nor U14429 (N_14429,N_13501,N_13577);
nor U14430 (N_14430,N_13771,N_13874);
or U14431 (N_14431,N_13526,N_13639);
and U14432 (N_14432,N_13660,N_13695);
nand U14433 (N_14433,N_13876,N_13641);
or U14434 (N_14434,N_13713,N_13500);
nand U14435 (N_14435,N_13546,N_13830);
or U14436 (N_14436,N_13656,N_13627);
nand U14437 (N_14437,N_13842,N_13782);
or U14438 (N_14438,N_13898,N_13654);
or U14439 (N_14439,N_13662,N_13657);
or U14440 (N_14440,N_13692,N_13708);
nand U14441 (N_14441,N_13969,N_13710);
nand U14442 (N_14442,N_13659,N_13534);
xnor U14443 (N_14443,N_13960,N_13767);
and U14444 (N_14444,N_13592,N_13902);
nor U14445 (N_14445,N_13685,N_13597);
xor U14446 (N_14446,N_13874,N_13517);
or U14447 (N_14447,N_13879,N_13896);
or U14448 (N_14448,N_13780,N_13783);
or U14449 (N_14449,N_13699,N_13943);
xnor U14450 (N_14450,N_13910,N_13510);
nor U14451 (N_14451,N_13741,N_13659);
and U14452 (N_14452,N_13999,N_13944);
nand U14453 (N_14453,N_13812,N_13829);
xnor U14454 (N_14454,N_13541,N_13694);
nand U14455 (N_14455,N_13907,N_13822);
or U14456 (N_14456,N_13972,N_13838);
nand U14457 (N_14457,N_13664,N_13737);
nor U14458 (N_14458,N_13917,N_13807);
xor U14459 (N_14459,N_13761,N_13988);
or U14460 (N_14460,N_13700,N_13977);
nor U14461 (N_14461,N_13609,N_13953);
and U14462 (N_14462,N_13949,N_13906);
nand U14463 (N_14463,N_13639,N_13633);
and U14464 (N_14464,N_13927,N_13685);
nand U14465 (N_14465,N_13715,N_13562);
nand U14466 (N_14466,N_13590,N_13733);
nand U14467 (N_14467,N_13720,N_13800);
xor U14468 (N_14468,N_13961,N_13801);
nand U14469 (N_14469,N_13972,N_13508);
nor U14470 (N_14470,N_13964,N_13893);
nor U14471 (N_14471,N_13739,N_13979);
or U14472 (N_14472,N_13804,N_13726);
nor U14473 (N_14473,N_13632,N_13604);
nor U14474 (N_14474,N_13810,N_13749);
nand U14475 (N_14475,N_13852,N_13781);
nor U14476 (N_14476,N_13887,N_13650);
xnor U14477 (N_14477,N_13589,N_13707);
and U14478 (N_14478,N_13988,N_13734);
nand U14479 (N_14479,N_13718,N_13739);
nand U14480 (N_14480,N_13887,N_13862);
nand U14481 (N_14481,N_13907,N_13766);
xnor U14482 (N_14482,N_13892,N_13991);
and U14483 (N_14483,N_13768,N_13639);
xnor U14484 (N_14484,N_13692,N_13819);
and U14485 (N_14485,N_13885,N_13686);
xor U14486 (N_14486,N_13564,N_13801);
or U14487 (N_14487,N_13850,N_13605);
and U14488 (N_14488,N_13715,N_13767);
and U14489 (N_14489,N_13775,N_13622);
xor U14490 (N_14490,N_13500,N_13661);
and U14491 (N_14491,N_13658,N_13906);
nor U14492 (N_14492,N_13633,N_13625);
and U14493 (N_14493,N_13656,N_13979);
or U14494 (N_14494,N_13737,N_13914);
and U14495 (N_14495,N_13842,N_13851);
xor U14496 (N_14496,N_13505,N_13773);
xor U14497 (N_14497,N_13710,N_13557);
and U14498 (N_14498,N_13674,N_13568);
nor U14499 (N_14499,N_13649,N_13951);
nor U14500 (N_14500,N_14449,N_14351);
xnor U14501 (N_14501,N_14496,N_14306);
or U14502 (N_14502,N_14477,N_14290);
nor U14503 (N_14503,N_14371,N_14051);
xnor U14504 (N_14504,N_14014,N_14191);
nor U14505 (N_14505,N_14322,N_14105);
or U14506 (N_14506,N_14283,N_14455);
and U14507 (N_14507,N_14197,N_14463);
nor U14508 (N_14508,N_14280,N_14245);
nand U14509 (N_14509,N_14128,N_14244);
nand U14510 (N_14510,N_14001,N_14331);
nor U14511 (N_14511,N_14470,N_14252);
nand U14512 (N_14512,N_14316,N_14321);
nor U14513 (N_14513,N_14412,N_14293);
and U14514 (N_14514,N_14210,N_14088);
nor U14515 (N_14515,N_14203,N_14053);
nor U14516 (N_14516,N_14281,N_14450);
nand U14517 (N_14517,N_14284,N_14246);
and U14518 (N_14518,N_14359,N_14074);
and U14519 (N_14519,N_14374,N_14383);
and U14520 (N_14520,N_14274,N_14048);
nor U14521 (N_14521,N_14260,N_14380);
nor U14522 (N_14522,N_14036,N_14382);
nand U14523 (N_14523,N_14190,N_14399);
nand U14524 (N_14524,N_14462,N_14405);
xnor U14525 (N_14525,N_14234,N_14159);
nor U14526 (N_14526,N_14440,N_14254);
xnor U14527 (N_14527,N_14062,N_14097);
and U14528 (N_14528,N_14023,N_14498);
and U14529 (N_14529,N_14099,N_14481);
xor U14530 (N_14530,N_14150,N_14340);
xor U14531 (N_14531,N_14186,N_14305);
nor U14532 (N_14532,N_14257,N_14390);
xor U14533 (N_14533,N_14117,N_14028);
xnor U14534 (N_14534,N_14221,N_14483);
nand U14535 (N_14535,N_14213,N_14156);
nor U14536 (N_14536,N_14182,N_14204);
and U14537 (N_14537,N_14148,N_14427);
nand U14538 (N_14538,N_14335,N_14010);
nor U14539 (N_14539,N_14441,N_14072);
and U14540 (N_14540,N_14307,N_14250);
nand U14541 (N_14541,N_14485,N_14188);
or U14542 (N_14542,N_14352,N_14233);
xor U14543 (N_14543,N_14466,N_14047);
and U14544 (N_14544,N_14157,N_14172);
and U14545 (N_14545,N_14024,N_14366);
nor U14546 (N_14546,N_14119,N_14478);
nand U14547 (N_14547,N_14318,N_14343);
nand U14548 (N_14548,N_14033,N_14431);
nand U14549 (N_14549,N_14385,N_14253);
and U14550 (N_14550,N_14314,N_14226);
and U14551 (N_14551,N_14402,N_14227);
nor U14552 (N_14552,N_14400,N_14414);
nor U14553 (N_14553,N_14046,N_14039);
nor U14554 (N_14554,N_14453,N_14208);
and U14555 (N_14555,N_14107,N_14392);
or U14556 (N_14556,N_14050,N_14138);
nand U14557 (N_14557,N_14230,N_14472);
and U14558 (N_14558,N_14177,N_14375);
nand U14559 (N_14559,N_14396,N_14214);
nor U14560 (N_14560,N_14241,N_14258);
or U14561 (N_14561,N_14327,N_14304);
nand U14562 (N_14562,N_14184,N_14266);
and U14563 (N_14563,N_14339,N_14419);
xnor U14564 (N_14564,N_14346,N_14476);
xor U14565 (N_14565,N_14464,N_14377);
xor U14566 (N_14566,N_14229,N_14296);
xnor U14567 (N_14567,N_14285,N_14178);
xor U14568 (N_14568,N_14486,N_14139);
nand U14569 (N_14569,N_14168,N_14360);
nor U14570 (N_14570,N_14243,N_14474);
or U14571 (N_14571,N_14131,N_14002);
nor U14572 (N_14572,N_14120,N_14092);
nand U14573 (N_14573,N_14066,N_14320);
nand U14574 (N_14574,N_14457,N_14038);
or U14575 (N_14575,N_14282,N_14323);
or U14576 (N_14576,N_14479,N_14225);
or U14577 (N_14577,N_14052,N_14170);
xor U14578 (N_14578,N_14146,N_14135);
and U14579 (N_14579,N_14403,N_14433);
and U14580 (N_14580,N_14446,N_14432);
nor U14581 (N_14581,N_14019,N_14009);
xnor U14582 (N_14582,N_14421,N_14086);
or U14583 (N_14583,N_14220,N_14013);
nor U14584 (N_14584,N_14059,N_14140);
and U14585 (N_14585,N_14060,N_14337);
xnor U14586 (N_14586,N_14232,N_14174);
nor U14587 (N_14587,N_14347,N_14034);
or U14588 (N_14588,N_14448,N_14078);
xnor U14589 (N_14589,N_14287,N_14492);
nand U14590 (N_14590,N_14218,N_14027);
xnor U14591 (N_14591,N_14365,N_14397);
nand U14592 (N_14592,N_14118,N_14101);
xor U14593 (N_14593,N_14011,N_14087);
xnor U14594 (N_14594,N_14445,N_14085);
nand U14595 (N_14595,N_14319,N_14357);
nor U14596 (N_14596,N_14373,N_14268);
and U14597 (N_14597,N_14249,N_14133);
nand U14598 (N_14598,N_14151,N_14176);
and U14599 (N_14599,N_14354,N_14144);
and U14600 (N_14600,N_14183,N_14363);
xor U14601 (N_14601,N_14114,N_14493);
or U14602 (N_14602,N_14008,N_14137);
nor U14603 (N_14603,N_14317,N_14263);
xnor U14604 (N_14604,N_14018,N_14299);
and U14605 (N_14605,N_14029,N_14003);
nor U14606 (N_14606,N_14211,N_14413);
or U14607 (N_14607,N_14270,N_14216);
or U14608 (N_14608,N_14080,N_14149);
nand U14609 (N_14609,N_14193,N_14124);
or U14610 (N_14610,N_14329,N_14169);
nor U14611 (N_14611,N_14298,N_14006);
nor U14612 (N_14612,N_14103,N_14369);
and U14613 (N_14613,N_14364,N_14461);
xor U14614 (N_14614,N_14411,N_14235);
or U14615 (N_14615,N_14044,N_14143);
nand U14616 (N_14616,N_14104,N_14109);
nand U14617 (N_14617,N_14292,N_14026);
and U14618 (N_14618,N_14388,N_14022);
nand U14619 (N_14619,N_14196,N_14325);
xnor U14620 (N_14620,N_14279,N_14082);
nor U14621 (N_14621,N_14090,N_14404);
or U14622 (N_14622,N_14112,N_14110);
nor U14623 (N_14623,N_14259,N_14032);
xnor U14624 (N_14624,N_14091,N_14145);
and U14625 (N_14625,N_14152,N_14198);
xnor U14626 (N_14626,N_14180,N_14142);
nor U14627 (N_14627,N_14348,N_14163);
and U14628 (N_14628,N_14065,N_14125);
nand U14629 (N_14629,N_14452,N_14158);
or U14630 (N_14630,N_14093,N_14269);
and U14631 (N_14631,N_14242,N_14236);
nand U14632 (N_14632,N_14239,N_14495);
xor U14633 (N_14633,N_14195,N_14378);
nand U14634 (N_14634,N_14376,N_14206);
nor U14635 (N_14635,N_14302,N_14491);
or U14636 (N_14636,N_14294,N_14056);
nand U14637 (N_14637,N_14115,N_14326);
or U14638 (N_14638,N_14437,N_14007);
nand U14639 (N_14639,N_14015,N_14394);
nand U14640 (N_14640,N_14454,N_14031);
nor U14641 (N_14641,N_14154,N_14408);
xnor U14642 (N_14642,N_14418,N_14079);
or U14643 (N_14643,N_14291,N_14488);
nor U14644 (N_14644,N_14460,N_14422);
nor U14645 (N_14645,N_14286,N_14406);
xnor U14646 (N_14646,N_14219,N_14123);
and U14647 (N_14647,N_14428,N_14181);
nor U14648 (N_14648,N_14289,N_14012);
and U14649 (N_14649,N_14054,N_14271);
or U14650 (N_14650,N_14370,N_14116);
nand U14651 (N_14651,N_14071,N_14121);
or U14652 (N_14652,N_14349,N_14132);
nand U14653 (N_14653,N_14467,N_14353);
nand U14654 (N_14654,N_14179,N_14468);
nand U14655 (N_14655,N_14267,N_14251);
nor U14656 (N_14656,N_14338,N_14275);
nor U14657 (N_14657,N_14362,N_14041);
and U14658 (N_14658,N_14155,N_14173);
nand U14659 (N_14659,N_14122,N_14113);
xnor U14660 (N_14660,N_14458,N_14215);
xor U14661 (N_14661,N_14407,N_14222);
nand U14662 (N_14662,N_14200,N_14309);
or U14663 (N_14663,N_14401,N_14265);
nand U14664 (N_14664,N_14209,N_14487);
and U14665 (N_14665,N_14212,N_14224);
nand U14666 (N_14666,N_14134,N_14482);
xor U14667 (N_14667,N_14175,N_14311);
nor U14668 (N_14668,N_14308,N_14136);
and U14669 (N_14669,N_14389,N_14000);
and U14670 (N_14670,N_14095,N_14430);
xor U14671 (N_14671,N_14126,N_14160);
xor U14672 (N_14672,N_14055,N_14435);
or U14673 (N_14673,N_14465,N_14185);
and U14674 (N_14674,N_14336,N_14301);
xnor U14675 (N_14675,N_14342,N_14303);
and U14676 (N_14676,N_14202,N_14420);
nor U14677 (N_14677,N_14297,N_14442);
nand U14678 (N_14678,N_14164,N_14076);
and U14679 (N_14679,N_14255,N_14187);
nor U14680 (N_14680,N_14248,N_14165);
nand U14681 (N_14681,N_14058,N_14497);
nand U14682 (N_14682,N_14207,N_14004);
or U14683 (N_14683,N_14333,N_14129);
nor U14684 (N_14684,N_14240,N_14276);
and U14685 (N_14685,N_14324,N_14199);
or U14686 (N_14686,N_14094,N_14189);
nand U14687 (N_14687,N_14436,N_14415);
xor U14688 (N_14688,N_14070,N_14098);
nor U14689 (N_14689,N_14330,N_14489);
nor U14690 (N_14690,N_14037,N_14409);
xnor U14691 (N_14691,N_14456,N_14127);
nor U14692 (N_14692,N_14475,N_14391);
nor U14693 (N_14693,N_14130,N_14426);
or U14694 (N_14694,N_14423,N_14021);
nor U14695 (N_14695,N_14379,N_14217);
xnor U14696 (N_14696,N_14057,N_14102);
nor U14697 (N_14697,N_14345,N_14061);
or U14698 (N_14698,N_14025,N_14494);
or U14699 (N_14699,N_14273,N_14484);
and U14700 (N_14700,N_14451,N_14344);
nor U14701 (N_14701,N_14171,N_14328);
nand U14702 (N_14702,N_14398,N_14434);
or U14703 (N_14703,N_14111,N_14334);
and U14704 (N_14704,N_14288,N_14231);
nand U14705 (N_14705,N_14035,N_14238);
nand U14706 (N_14706,N_14499,N_14106);
nand U14707 (N_14707,N_14017,N_14381);
xor U14708 (N_14708,N_14417,N_14272);
nand U14709 (N_14709,N_14443,N_14100);
and U14710 (N_14710,N_14332,N_14147);
nand U14711 (N_14711,N_14069,N_14192);
nor U14712 (N_14712,N_14312,N_14077);
nand U14713 (N_14713,N_14262,N_14194);
nand U14714 (N_14714,N_14490,N_14313);
or U14715 (N_14715,N_14020,N_14416);
or U14716 (N_14716,N_14030,N_14084);
or U14717 (N_14717,N_14310,N_14438);
xnor U14718 (N_14718,N_14469,N_14108);
or U14719 (N_14719,N_14410,N_14201);
and U14720 (N_14720,N_14205,N_14393);
nor U14721 (N_14721,N_14247,N_14045);
xor U14722 (N_14722,N_14261,N_14368);
and U14723 (N_14723,N_14264,N_14425);
or U14724 (N_14724,N_14166,N_14439);
xor U14725 (N_14725,N_14075,N_14063);
and U14726 (N_14726,N_14081,N_14223);
and U14727 (N_14727,N_14384,N_14444);
xnor U14728 (N_14728,N_14042,N_14395);
and U14729 (N_14729,N_14043,N_14162);
xor U14730 (N_14730,N_14355,N_14040);
xor U14731 (N_14731,N_14424,N_14228);
or U14732 (N_14732,N_14064,N_14277);
and U14733 (N_14733,N_14480,N_14167);
nor U14734 (N_14734,N_14473,N_14089);
nor U14735 (N_14735,N_14386,N_14459);
xor U14736 (N_14736,N_14372,N_14367);
nand U14737 (N_14737,N_14278,N_14005);
nand U14738 (N_14738,N_14153,N_14083);
xor U14739 (N_14739,N_14016,N_14096);
nor U14740 (N_14740,N_14161,N_14361);
or U14741 (N_14741,N_14049,N_14350);
xor U14742 (N_14742,N_14141,N_14067);
or U14743 (N_14743,N_14429,N_14447);
and U14744 (N_14744,N_14315,N_14387);
nand U14745 (N_14745,N_14300,N_14356);
and U14746 (N_14746,N_14073,N_14256);
or U14747 (N_14747,N_14068,N_14237);
nor U14748 (N_14748,N_14341,N_14358);
or U14749 (N_14749,N_14471,N_14295);
nor U14750 (N_14750,N_14349,N_14098);
nor U14751 (N_14751,N_14315,N_14105);
nor U14752 (N_14752,N_14092,N_14040);
xnor U14753 (N_14753,N_14200,N_14488);
nor U14754 (N_14754,N_14392,N_14108);
or U14755 (N_14755,N_14304,N_14180);
or U14756 (N_14756,N_14241,N_14056);
and U14757 (N_14757,N_14159,N_14333);
and U14758 (N_14758,N_14236,N_14371);
or U14759 (N_14759,N_14212,N_14343);
and U14760 (N_14760,N_14493,N_14430);
xor U14761 (N_14761,N_14009,N_14223);
nor U14762 (N_14762,N_14482,N_14198);
nor U14763 (N_14763,N_14020,N_14485);
xnor U14764 (N_14764,N_14111,N_14214);
xnor U14765 (N_14765,N_14456,N_14046);
and U14766 (N_14766,N_14276,N_14027);
xnor U14767 (N_14767,N_14463,N_14151);
nor U14768 (N_14768,N_14081,N_14341);
or U14769 (N_14769,N_14028,N_14085);
xnor U14770 (N_14770,N_14239,N_14312);
nor U14771 (N_14771,N_14048,N_14324);
and U14772 (N_14772,N_14201,N_14267);
xor U14773 (N_14773,N_14258,N_14493);
and U14774 (N_14774,N_14409,N_14329);
and U14775 (N_14775,N_14244,N_14099);
or U14776 (N_14776,N_14057,N_14086);
or U14777 (N_14777,N_14444,N_14419);
nor U14778 (N_14778,N_14167,N_14105);
and U14779 (N_14779,N_14172,N_14135);
and U14780 (N_14780,N_14181,N_14026);
xor U14781 (N_14781,N_14237,N_14079);
xor U14782 (N_14782,N_14467,N_14375);
nor U14783 (N_14783,N_14493,N_14259);
nand U14784 (N_14784,N_14458,N_14294);
nand U14785 (N_14785,N_14433,N_14119);
nor U14786 (N_14786,N_14232,N_14303);
and U14787 (N_14787,N_14293,N_14024);
nor U14788 (N_14788,N_14383,N_14236);
and U14789 (N_14789,N_14351,N_14424);
and U14790 (N_14790,N_14272,N_14222);
or U14791 (N_14791,N_14254,N_14326);
nand U14792 (N_14792,N_14153,N_14377);
nand U14793 (N_14793,N_14394,N_14115);
or U14794 (N_14794,N_14163,N_14131);
and U14795 (N_14795,N_14096,N_14480);
or U14796 (N_14796,N_14338,N_14457);
and U14797 (N_14797,N_14351,N_14378);
and U14798 (N_14798,N_14222,N_14332);
nand U14799 (N_14799,N_14121,N_14264);
nand U14800 (N_14800,N_14338,N_14447);
and U14801 (N_14801,N_14272,N_14331);
or U14802 (N_14802,N_14128,N_14034);
xor U14803 (N_14803,N_14060,N_14405);
xor U14804 (N_14804,N_14323,N_14347);
nand U14805 (N_14805,N_14199,N_14047);
xor U14806 (N_14806,N_14473,N_14342);
or U14807 (N_14807,N_14095,N_14388);
nand U14808 (N_14808,N_14445,N_14342);
or U14809 (N_14809,N_14499,N_14100);
xor U14810 (N_14810,N_14339,N_14065);
nor U14811 (N_14811,N_14273,N_14337);
and U14812 (N_14812,N_14153,N_14104);
and U14813 (N_14813,N_14034,N_14055);
and U14814 (N_14814,N_14499,N_14406);
xnor U14815 (N_14815,N_14016,N_14030);
nor U14816 (N_14816,N_14104,N_14273);
xnor U14817 (N_14817,N_14471,N_14288);
nand U14818 (N_14818,N_14493,N_14418);
and U14819 (N_14819,N_14098,N_14460);
nand U14820 (N_14820,N_14076,N_14408);
and U14821 (N_14821,N_14311,N_14438);
nand U14822 (N_14822,N_14313,N_14262);
xor U14823 (N_14823,N_14150,N_14172);
or U14824 (N_14824,N_14102,N_14279);
nand U14825 (N_14825,N_14065,N_14241);
or U14826 (N_14826,N_14480,N_14422);
nand U14827 (N_14827,N_14471,N_14083);
and U14828 (N_14828,N_14246,N_14146);
nor U14829 (N_14829,N_14378,N_14340);
and U14830 (N_14830,N_14392,N_14400);
or U14831 (N_14831,N_14487,N_14227);
nand U14832 (N_14832,N_14189,N_14055);
nor U14833 (N_14833,N_14223,N_14436);
nand U14834 (N_14834,N_14185,N_14166);
and U14835 (N_14835,N_14387,N_14346);
and U14836 (N_14836,N_14473,N_14196);
and U14837 (N_14837,N_14481,N_14207);
and U14838 (N_14838,N_14320,N_14016);
nand U14839 (N_14839,N_14410,N_14061);
and U14840 (N_14840,N_14046,N_14047);
nand U14841 (N_14841,N_14442,N_14370);
and U14842 (N_14842,N_14012,N_14251);
and U14843 (N_14843,N_14353,N_14419);
and U14844 (N_14844,N_14368,N_14497);
and U14845 (N_14845,N_14484,N_14232);
and U14846 (N_14846,N_14077,N_14005);
or U14847 (N_14847,N_14028,N_14475);
or U14848 (N_14848,N_14114,N_14483);
nand U14849 (N_14849,N_14135,N_14119);
xor U14850 (N_14850,N_14470,N_14172);
or U14851 (N_14851,N_14158,N_14090);
and U14852 (N_14852,N_14024,N_14446);
or U14853 (N_14853,N_14350,N_14498);
or U14854 (N_14854,N_14010,N_14328);
and U14855 (N_14855,N_14046,N_14408);
nor U14856 (N_14856,N_14248,N_14333);
nor U14857 (N_14857,N_14274,N_14062);
xor U14858 (N_14858,N_14080,N_14079);
nor U14859 (N_14859,N_14199,N_14025);
nand U14860 (N_14860,N_14184,N_14210);
or U14861 (N_14861,N_14261,N_14354);
nor U14862 (N_14862,N_14192,N_14055);
nand U14863 (N_14863,N_14327,N_14020);
and U14864 (N_14864,N_14166,N_14058);
and U14865 (N_14865,N_14122,N_14202);
xnor U14866 (N_14866,N_14324,N_14030);
nor U14867 (N_14867,N_14186,N_14104);
and U14868 (N_14868,N_14158,N_14343);
or U14869 (N_14869,N_14185,N_14257);
nor U14870 (N_14870,N_14160,N_14371);
or U14871 (N_14871,N_14047,N_14138);
and U14872 (N_14872,N_14465,N_14333);
nor U14873 (N_14873,N_14337,N_14277);
or U14874 (N_14874,N_14013,N_14355);
xnor U14875 (N_14875,N_14125,N_14451);
and U14876 (N_14876,N_14008,N_14025);
and U14877 (N_14877,N_14025,N_14463);
xnor U14878 (N_14878,N_14324,N_14353);
nand U14879 (N_14879,N_14196,N_14464);
and U14880 (N_14880,N_14032,N_14471);
nand U14881 (N_14881,N_14243,N_14334);
nand U14882 (N_14882,N_14432,N_14276);
nand U14883 (N_14883,N_14299,N_14303);
xor U14884 (N_14884,N_14397,N_14415);
or U14885 (N_14885,N_14277,N_14117);
nor U14886 (N_14886,N_14265,N_14445);
and U14887 (N_14887,N_14116,N_14462);
nand U14888 (N_14888,N_14354,N_14271);
nand U14889 (N_14889,N_14475,N_14379);
or U14890 (N_14890,N_14244,N_14211);
nand U14891 (N_14891,N_14206,N_14061);
or U14892 (N_14892,N_14411,N_14129);
nor U14893 (N_14893,N_14316,N_14291);
nor U14894 (N_14894,N_14347,N_14313);
or U14895 (N_14895,N_14210,N_14351);
nor U14896 (N_14896,N_14199,N_14293);
and U14897 (N_14897,N_14168,N_14047);
nand U14898 (N_14898,N_14010,N_14413);
nor U14899 (N_14899,N_14111,N_14459);
nand U14900 (N_14900,N_14274,N_14260);
xnor U14901 (N_14901,N_14019,N_14059);
xnor U14902 (N_14902,N_14261,N_14039);
nor U14903 (N_14903,N_14029,N_14115);
or U14904 (N_14904,N_14164,N_14157);
xnor U14905 (N_14905,N_14340,N_14064);
nand U14906 (N_14906,N_14399,N_14104);
xor U14907 (N_14907,N_14316,N_14295);
xnor U14908 (N_14908,N_14303,N_14062);
or U14909 (N_14909,N_14007,N_14360);
nor U14910 (N_14910,N_14209,N_14315);
nand U14911 (N_14911,N_14060,N_14324);
nor U14912 (N_14912,N_14462,N_14188);
or U14913 (N_14913,N_14249,N_14358);
or U14914 (N_14914,N_14414,N_14191);
xnor U14915 (N_14915,N_14186,N_14065);
and U14916 (N_14916,N_14207,N_14451);
nand U14917 (N_14917,N_14067,N_14241);
xor U14918 (N_14918,N_14113,N_14332);
and U14919 (N_14919,N_14057,N_14404);
xor U14920 (N_14920,N_14035,N_14223);
nor U14921 (N_14921,N_14246,N_14305);
nand U14922 (N_14922,N_14445,N_14090);
or U14923 (N_14923,N_14085,N_14025);
nor U14924 (N_14924,N_14043,N_14102);
nand U14925 (N_14925,N_14180,N_14027);
or U14926 (N_14926,N_14431,N_14022);
xnor U14927 (N_14927,N_14302,N_14325);
nand U14928 (N_14928,N_14086,N_14477);
and U14929 (N_14929,N_14378,N_14274);
xnor U14930 (N_14930,N_14159,N_14162);
and U14931 (N_14931,N_14025,N_14010);
or U14932 (N_14932,N_14282,N_14371);
nand U14933 (N_14933,N_14329,N_14156);
nand U14934 (N_14934,N_14038,N_14441);
xor U14935 (N_14935,N_14449,N_14446);
nand U14936 (N_14936,N_14146,N_14400);
nand U14937 (N_14937,N_14220,N_14477);
and U14938 (N_14938,N_14130,N_14371);
nor U14939 (N_14939,N_14016,N_14060);
nand U14940 (N_14940,N_14127,N_14176);
or U14941 (N_14941,N_14477,N_14361);
nand U14942 (N_14942,N_14093,N_14366);
nor U14943 (N_14943,N_14168,N_14329);
xnor U14944 (N_14944,N_14215,N_14280);
nor U14945 (N_14945,N_14239,N_14030);
xor U14946 (N_14946,N_14177,N_14230);
nor U14947 (N_14947,N_14320,N_14252);
nor U14948 (N_14948,N_14284,N_14074);
and U14949 (N_14949,N_14255,N_14275);
nand U14950 (N_14950,N_14083,N_14277);
xnor U14951 (N_14951,N_14050,N_14057);
or U14952 (N_14952,N_14444,N_14129);
nor U14953 (N_14953,N_14496,N_14380);
and U14954 (N_14954,N_14456,N_14339);
xor U14955 (N_14955,N_14275,N_14237);
and U14956 (N_14956,N_14178,N_14365);
or U14957 (N_14957,N_14429,N_14317);
nor U14958 (N_14958,N_14291,N_14498);
and U14959 (N_14959,N_14184,N_14444);
nor U14960 (N_14960,N_14403,N_14055);
nand U14961 (N_14961,N_14446,N_14196);
xnor U14962 (N_14962,N_14137,N_14219);
or U14963 (N_14963,N_14154,N_14217);
nand U14964 (N_14964,N_14295,N_14149);
nor U14965 (N_14965,N_14311,N_14006);
xnor U14966 (N_14966,N_14120,N_14311);
xor U14967 (N_14967,N_14148,N_14484);
and U14968 (N_14968,N_14064,N_14190);
and U14969 (N_14969,N_14034,N_14271);
xnor U14970 (N_14970,N_14188,N_14302);
or U14971 (N_14971,N_14165,N_14202);
xnor U14972 (N_14972,N_14054,N_14078);
nand U14973 (N_14973,N_14242,N_14033);
nand U14974 (N_14974,N_14191,N_14274);
nand U14975 (N_14975,N_14239,N_14259);
nand U14976 (N_14976,N_14103,N_14243);
and U14977 (N_14977,N_14155,N_14484);
xor U14978 (N_14978,N_14246,N_14136);
and U14979 (N_14979,N_14102,N_14014);
nand U14980 (N_14980,N_14417,N_14409);
nand U14981 (N_14981,N_14040,N_14108);
nor U14982 (N_14982,N_14060,N_14226);
and U14983 (N_14983,N_14189,N_14386);
nand U14984 (N_14984,N_14308,N_14199);
nand U14985 (N_14985,N_14458,N_14452);
nor U14986 (N_14986,N_14113,N_14198);
xor U14987 (N_14987,N_14236,N_14142);
or U14988 (N_14988,N_14429,N_14102);
or U14989 (N_14989,N_14002,N_14154);
xnor U14990 (N_14990,N_14278,N_14279);
nor U14991 (N_14991,N_14365,N_14271);
and U14992 (N_14992,N_14453,N_14469);
or U14993 (N_14993,N_14121,N_14154);
nor U14994 (N_14994,N_14316,N_14402);
xnor U14995 (N_14995,N_14441,N_14483);
or U14996 (N_14996,N_14310,N_14344);
and U14997 (N_14997,N_14411,N_14383);
and U14998 (N_14998,N_14088,N_14421);
and U14999 (N_14999,N_14218,N_14494);
nand UO_0 (O_0,N_14982,N_14718);
xnor UO_1 (O_1,N_14734,N_14891);
nand UO_2 (O_2,N_14987,N_14903);
xnor UO_3 (O_3,N_14793,N_14604);
nand UO_4 (O_4,N_14904,N_14876);
or UO_5 (O_5,N_14881,N_14935);
nand UO_6 (O_6,N_14698,N_14675);
xnor UO_7 (O_7,N_14629,N_14530);
and UO_8 (O_8,N_14852,N_14589);
nand UO_9 (O_9,N_14840,N_14551);
nand UO_10 (O_10,N_14562,N_14528);
xor UO_11 (O_11,N_14612,N_14785);
nor UO_12 (O_12,N_14522,N_14520);
and UO_13 (O_13,N_14864,N_14556);
or UO_14 (O_14,N_14662,N_14906);
nor UO_15 (O_15,N_14776,N_14536);
nand UO_16 (O_16,N_14704,N_14567);
xor UO_17 (O_17,N_14569,N_14839);
and UO_18 (O_18,N_14884,N_14598);
nand UO_19 (O_19,N_14766,N_14751);
and UO_20 (O_20,N_14601,N_14654);
nor UO_21 (O_21,N_14949,N_14981);
and UO_22 (O_22,N_14989,N_14773);
nand UO_23 (O_23,N_14771,N_14874);
nand UO_24 (O_24,N_14679,N_14533);
xor UO_25 (O_25,N_14924,N_14827);
nand UO_26 (O_26,N_14653,N_14646);
nand UO_27 (O_27,N_14507,N_14568);
nor UO_28 (O_28,N_14972,N_14710);
xor UO_29 (O_29,N_14740,N_14505);
and UO_30 (O_30,N_14560,N_14756);
xor UO_31 (O_31,N_14965,N_14558);
xor UO_32 (O_32,N_14790,N_14846);
or UO_33 (O_33,N_14579,N_14597);
xnor UO_34 (O_34,N_14584,N_14768);
nand UO_35 (O_35,N_14594,N_14655);
or UO_36 (O_36,N_14978,N_14842);
nor UO_37 (O_37,N_14592,N_14697);
nand UO_38 (O_38,N_14921,N_14755);
nand UO_39 (O_39,N_14923,N_14915);
or UO_40 (O_40,N_14749,N_14600);
xor UO_41 (O_41,N_14943,N_14788);
xnor UO_42 (O_42,N_14540,N_14649);
and UO_43 (O_43,N_14825,N_14815);
nor UO_44 (O_44,N_14831,N_14832);
or UO_45 (O_45,N_14913,N_14549);
nand UO_46 (O_46,N_14779,N_14931);
or UO_47 (O_47,N_14626,N_14919);
or UO_48 (O_48,N_14585,N_14714);
xor UO_49 (O_49,N_14819,N_14859);
or UO_50 (O_50,N_14786,N_14680);
nand UO_51 (O_51,N_14880,N_14747);
and UO_52 (O_52,N_14835,N_14983);
nor UO_53 (O_53,N_14848,N_14553);
nor UO_54 (O_54,N_14609,N_14555);
xor UO_55 (O_55,N_14878,N_14684);
nor UO_56 (O_56,N_14810,N_14761);
xnor UO_57 (O_57,N_14503,N_14844);
or UO_58 (O_58,N_14741,N_14535);
or UO_59 (O_59,N_14525,N_14527);
xor UO_60 (O_60,N_14754,N_14713);
or UO_61 (O_61,N_14944,N_14501);
nand UO_62 (O_62,N_14865,N_14582);
or UO_63 (O_63,N_14886,N_14664);
xor UO_64 (O_64,N_14709,N_14705);
and UO_65 (O_65,N_14621,N_14985);
and UO_66 (O_66,N_14937,N_14509);
and UO_67 (O_67,N_14628,N_14619);
or UO_68 (O_68,N_14733,N_14753);
and UO_69 (O_69,N_14606,N_14860);
xor UO_70 (O_70,N_14663,N_14712);
and UO_71 (O_71,N_14564,N_14991);
and UO_72 (O_72,N_14523,N_14632);
or UO_73 (O_73,N_14538,N_14678);
xor UO_74 (O_74,N_14807,N_14820);
xor UO_75 (O_75,N_14932,N_14506);
and UO_76 (O_76,N_14951,N_14833);
or UO_77 (O_77,N_14732,N_14566);
xor UO_78 (O_78,N_14830,N_14805);
nand UO_79 (O_79,N_14554,N_14877);
or UO_80 (O_80,N_14961,N_14813);
nor UO_81 (O_81,N_14973,N_14959);
xnor UO_82 (O_82,N_14681,N_14752);
nand UO_83 (O_83,N_14542,N_14795);
nand UO_84 (O_84,N_14611,N_14623);
nor UO_85 (O_85,N_14745,N_14939);
and UO_86 (O_86,N_14797,N_14563);
nand UO_87 (O_87,N_14581,N_14834);
and UO_88 (O_88,N_14724,N_14738);
nor UO_89 (O_89,N_14955,N_14706);
or UO_90 (O_90,N_14764,N_14984);
xor UO_91 (O_91,N_14822,N_14950);
and UO_92 (O_92,N_14742,N_14690);
or UO_93 (O_93,N_14896,N_14658);
nor UO_94 (O_94,N_14513,N_14873);
nand UO_95 (O_95,N_14858,N_14963);
and UO_96 (O_96,N_14673,N_14999);
nor UO_97 (O_97,N_14739,N_14909);
and UO_98 (O_98,N_14784,N_14707);
and UO_99 (O_99,N_14573,N_14547);
nor UO_100 (O_100,N_14660,N_14758);
nand UO_101 (O_101,N_14996,N_14731);
nand UO_102 (O_102,N_14635,N_14767);
nand UO_103 (O_103,N_14726,N_14613);
nor UO_104 (O_104,N_14941,N_14644);
nand UO_105 (O_105,N_14798,N_14716);
nor UO_106 (O_106,N_14537,N_14637);
and UO_107 (O_107,N_14970,N_14721);
and UO_108 (O_108,N_14723,N_14574);
or UO_109 (O_109,N_14605,N_14759);
nand UO_110 (O_110,N_14922,N_14521);
nand UO_111 (O_111,N_14901,N_14998);
and UO_112 (O_112,N_14997,N_14518);
nor UO_113 (O_113,N_14648,N_14593);
nand UO_114 (O_114,N_14847,N_14888);
and UO_115 (O_115,N_14502,N_14791);
xnor UO_116 (O_116,N_14603,N_14920);
or UO_117 (O_117,N_14953,N_14727);
nor UO_118 (O_118,N_14954,N_14770);
nor UO_119 (O_119,N_14661,N_14866);
xnor UO_120 (O_120,N_14682,N_14557);
nand UO_121 (O_121,N_14657,N_14514);
xnor UO_122 (O_122,N_14602,N_14689);
nand UO_123 (O_123,N_14668,N_14722);
nand UO_124 (O_124,N_14836,N_14801);
nand UO_125 (O_125,N_14652,N_14552);
nand UO_126 (O_126,N_14572,N_14889);
nor UO_127 (O_127,N_14647,N_14804);
nand UO_128 (O_128,N_14890,N_14599);
or UO_129 (O_129,N_14700,N_14960);
nand UO_130 (O_130,N_14559,N_14760);
nand UO_131 (O_131,N_14728,N_14578);
and UO_132 (O_132,N_14976,N_14942);
nor UO_133 (O_133,N_14843,N_14677);
xor UO_134 (O_134,N_14957,N_14672);
nand UO_135 (O_135,N_14945,N_14691);
nand UO_136 (O_136,N_14643,N_14841);
xnor UO_137 (O_137,N_14783,N_14868);
and UO_138 (O_138,N_14683,N_14782);
nor UO_139 (O_139,N_14781,N_14817);
nor UO_140 (O_140,N_14516,N_14777);
nor UO_141 (O_141,N_14787,N_14634);
xor UO_142 (O_142,N_14561,N_14853);
xor UO_143 (O_143,N_14814,N_14746);
and UO_144 (O_144,N_14715,N_14762);
nor UO_145 (O_145,N_14640,N_14616);
or UO_146 (O_146,N_14799,N_14774);
or UO_147 (O_147,N_14818,N_14656);
and UO_148 (O_148,N_14702,N_14674);
nand UO_149 (O_149,N_14630,N_14809);
nand UO_150 (O_150,N_14837,N_14615);
and UO_151 (O_151,N_14899,N_14948);
and UO_152 (O_152,N_14975,N_14927);
xnor UO_153 (O_153,N_14703,N_14812);
and UO_154 (O_154,N_14631,N_14570);
xnor UO_155 (O_155,N_14838,N_14974);
nand UO_156 (O_156,N_14962,N_14544);
or UO_157 (O_157,N_14821,N_14515);
nor UO_158 (O_158,N_14775,N_14968);
or UO_159 (O_159,N_14645,N_14519);
xor UO_160 (O_160,N_14571,N_14531);
nand UO_161 (O_161,N_14686,N_14665);
or UO_162 (O_162,N_14845,N_14875);
or UO_163 (O_163,N_14946,N_14808);
xor UO_164 (O_164,N_14938,N_14666);
xnor UO_165 (O_165,N_14826,N_14918);
and UO_166 (O_166,N_14622,N_14641);
xor UO_167 (O_167,N_14737,N_14977);
or UO_168 (O_168,N_14511,N_14928);
xnor UO_169 (O_169,N_14806,N_14895);
nand UO_170 (O_170,N_14929,N_14794);
and UO_171 (O_171,N_14869,N_14796);
and UO_172 (O_172,N_14883,N_14917);
and UO_173 (O_173,N_14851,N_14550);
nand UO_174 (O_174,N_14517,N_14699);
or UO_175 (O_175,N_14988,N_14912);
and UO_176 (O_176,N_14855,N_14701);
nand UO_177 (O_177,N_14894,N_14930);
nor UO_178 (O_178,N_14575,N_14638);
nand UO_179 (O_179,N_14828,N_14729);
nand UO_180 (O_180,N_14992,N_14980);
nand UO_181 (O_181,N_14879,N_14580);
xnor UO_182 (O_182,N_14867,N_14688);
and UO_183 (O_183,N_14757,N_14824);
nor UO_184 (O_184,N_14743,N_14636);
or UO_185 (O_185,N_14548,N_14720);
nand UO_186 (O_186,N_14914,N_14565);
and UO_187 (O_187,N_14995,N_14882);
xnor UO_188 (O_188,N_14769,N_14934);
nand UO_189 (O_189,N_14711,N_14504);
and UO_190 (O_190,N_14532,N_14862);
and UO_191 (O_191,N_14971,N_14614);
nor UO_192 (O_192,N_14811,N_14633);
nor UO_193 (O_193,N_14534,N_14687);
and UO_194 (O_194,N_14861,N_14926);
or UO_195 (O_195,N_14789,N_14803);
xnor UO_196 (O_196,N_14854,N_14541);
nor UO_197 (O_197,N_14908,N_14586);
and UO_198 (O_198,N_14545,N_14670);
nand UO_199 (O_199,N_14748,N_14671);
and UO_200 (O_200,N_14529,N_14897);
nand UO_201 (O_201,N_14667,N_14856);
and UO_202 (O_202,N_14650,N_14870);
and UO_203 (O_203,N_14676,N_14588);
xor UO_204 (O_204,N_14508,N_14823);
nor UO_205 (O_205,N_14816,N_14624);
nor UO_206 (O_206,N_14956,N_14872);
nand UO_207 (O_207,N_14990,N_14587);
nand UO_208 (O_208,N_14947,N_14893);
or UO_209 (O_209,N_14608,N_14750);
nor UO_210 (O_210,N_14898,N_14863);
or UO_211 (O_211,N_14902,N_14730);
nor UO_212 (O_212,N_14925,N_14576);
nor UO_213 (O_213,N_14979,N_14543);
and UO_214 (O_214,N_14850,N_14696);
nand UO_215 (O_215,N_14911,N_14964);
nand UO_216 (O_216,N_14717,N_14546);
and UO_217 (O_217,N_14892,N_14857);
nor UO_218 (O_218,N_14642,N_14607);
or UO_219 (O_219,N_14763,N_14617);
and UO_220 (O_220,N_14887,N_14933);
or UO_221 (O_221,N_14591,N_14910);
nand UO_222 (O_222,N_14958,N_14765);
xnor UO_223 (O_223,N_14871,N_14772);
nand UO_224 (O_224,N_14595,N_14627);
and UO_225 (O_225,N_14526,N_14610);
and UO_226 (O_226,N_14802,N_14651);
and UO_227 (O_227,N_14695,N_14618);
and UO_228 (O_228,N_14524,N_14669);
xor UO_229 (O_229,N_14500,N_14800);
xor UO_230 (O_230,N_14639,N_14916);
nand UO_231 (O_231,N_14829,N_14778);
nand UO_232 (O_232,N_14969,N_14659);
xor UO_233 (O_233,N_14539,N_14967);
or UO_234 (O_234,N_14692,N_14966);
nor UO_235 (O_235,N_14885,N_14719);
and UO_236 (O_236,N_14735,N_14590);
and UO_237 (O_237,N_14725,N_14993);
and UO_238 (O_238,N_14849,N_14986);
and UO_239 (O_239,N_14792,N_14744);
nand UO_240 (O_240,N_14596,N_14936);
and UO_241 (O_241,N_14693,N_14994);
nand UO_242 (O_242,N_14952,N_14940);
xnor UO_243 (O_243,N_14900,N_14708);
xor UO_244 (O_244,N_14694,N_14907);
nor UO_245 (O_245,N_14583,N_14625);
nand UO_246 (O_246,N_14620,N_14510);
or UO_247 (O_247,N_14512,N_14780);
or UO_248 (O_248,N_14577,N_14736);
or UO_249 (O_249,N_14905,N_14685);
xnor UO_250 (O_250,N_14958,N_14862);
or UO_251 (O_251,N_14532,N_14871);
nor UO_252 (O_252,N_14798,N_14719);
or UO_253 (O_253,N_14618,N_14944);
nand UO_254 (O_254,N_14841,N_14528);
and UO_255 (O_255,N_14722,N_14923);
xor UO_256 (O_256,N_14670,N_14897);
nand UO_257 (O_257,N_14661,N_14645);
and UO_258 (O_258,N_14718,N_14751);
and UO_259 (O_259,N_14831,N_14788);
nor UO_260 (O_260,N_14877,N_14637);
nand UO_261 (O_261,N_14752,N_14664);
xor UO_262 (O_262,N_14580,N_14853);
and UO_263 (O_263,N_14742,N_14835);
xor UO_264 (O_264,N_14573,N_14649);
nor UO_265 (O_265,N_14529,N_14502);
xnor UO_266 (O_266,N_14920,N_14522);
nor UO_267 (O_267,N_14627,N_14809);
nand UO_268 (O_268,N_14793,N_14651);
nor UO_269 (O_269,N_14596,N_14632);
and UO_270 (O_270,N_14759,N_14617);
nand UO_271 (O_271,N_14598,N_14665);
and UO_272 (O_272,N_14843,N_14895);
nor UO_273 (O_273,N_14756,N_14510);
nand UO_274 (O_274,N_14625,N_14676);
xor UO_275 (O_275,N_14700,N_14906);
or UO_276 (O_276,N_14566,N_14579);
nand UO_277 (O_277,N_14839,N_14958);
or UO_278 (O_278,N_14720,N_14618);
nor UO_279 (O_279,N_14907,N_14859);
and UO_280 (O_280,N_14596,N_14548);
nand UO_281 (O_281,N_14551,N_14980);
nor UO_282 (O_282,N_14686,N_14991);
and UO_283 (O_283,N_14883,N_14704);
nand UO_284 (O_284,N_14946,N_14924);
and UO_285 (O_285,N_14959,N_14550);
xor UO_286 (O_286,N_14635,N_14510);
or UO_287 (O_287,N_14615,N_14860);
xor UO_288 (O_288,N_14720,N_14732);
nand UO_289 (O_289,N_14661,N_14829);
and UO_290 (O_290,N_14807,N_14956);
nand UO_291 (O_291,N_14849,N_14578);
and UO_292 (O_292,N_14968,N_14896);
nand UO_293 (O_293,N_14800,N_14649);
nor UO_294 (O_294,N_14865,N_14679);
and UO_295 (O_295,N_14605,N_14536);
or UO_296 (O_296,N_14510,N_14546);
nand UO_297 (O_297,N_14836,N_14827);
nand UO_298 (O_298,N_14940,N_14845);
xnor UO_299 (O_299,N_14619,N_14577);
nor UO_300 (O_300,N_14730,N_14573);
nand UO_301 (O_301,N_14695,N_14986);
nand UO_302 (O_302,N_14773,N_14934);
or UO_303 (O_303,N_14845,N_14678);
nor UO_304 (O_304,N_14682,N_14694);
and UO_305 (O_305,N_14827,N_14720);
nand UO_306 (O_306,N_14931,N_14676);
or UO_307 (O_307,N_14833,N_14855);
nand UO_308 (O_308,N_14828,N_14704);
nor UO_309 (O_309,N_14998,N_14972);
or UO_310 (O_310,N_14925,N_14642);
and UO_311 (O_311,N_14753,N_14831);
and UO_312 (O_312,N_14798,N_14975);
or UO_313 (O_313,N_14634,N_14555);
or UO_314 (O_314,N_14620,N_14570);
and UO_315 (O_315,N_14806,N_14840);
xnor UO_316 (O_316,N_14504,N_14522);
xnor UO_317 (O_317,N_14579,N_14525);
xor UO_318 (O_318,N_14836,N_14849);
nor UO_319 (O_319,N_14706,N_14832);
or UO_320 (O_320,N_14962,N_14923);
xnor UO_321 (O_321,N_14503,N_14671);
or UO_322 (O_322,N_14983,N_14656);
nor UO_323 (O_323,N_14691,N_14814);
and UO_324 (O_324,N_14716,N_14563);
nor UO_325 (O_325,N_14840,N_14653);
nand UO_326 (O_326,N_14881,N_14947);
and UO_327 (O_327,N_14791,N_14727);
xor UO_328 (O_328,N_14836,N_14806);
xor UO_329 (O_329,N_14849,N_14553);
and UO_330 (O_330,N_14812,N_14942);
and UO_331 (O_331,N_14565,N_14838);
and UO_332 (O_332,N_14713,N_14970);
xnor UO_333 (O_333,N_14771,N_14529);
xnor UO_334 (O_334,N_14694,N_14997);
xor UO_335 (O_335,N_14893,N_14912);
nand UO_336 (O_336,N_14690,N_14532);
and UO_337 (O_337,N_14666,N_14543);
nand UO_338 (O_338,N_14653,N_14663);
nor UO_339 (O_339,N_14760,N_14673);
nand UO_340 (O_340,N_14722,N_14799);
xor UO_341 (O_341,N_14870,N_14964);
nor UO_342 (O_342,N_14582,N_14563);
nand UO_343 (O_343,N_14695,N_14780);
nand UO_344 (O_344,N_14767,N_14892);
or UO_345 (O_345,N_14847,N_14513);
or UO_346 (O_346,N_14908,N_14511);
or UO_347 (O_347,N_14858,N_14709);
nand UO_348 (O_348,N_14875,N_14626);
or UO_349 (O_349,N_14611,N_14628);
nand UO_350 (O_350,N_14842,N_14662);
and UO_351 (O_351,N_14548,N_14610);
or UO_352 (O_352,N_14560,N_14955);
and UO_353 (O_353,N_14732,N_14661);
or UO_354 (O_354,N_14568,N_14530);
nor UO_355 (O_355,N_14804,N_14632);
xnor UO_356 (O_356,N_14755,N_14682);
or UO_357 (O_357,N_14965,N_14542);
nand UO_358 (O_358,N_14595,N_14763);
nand UO_359 (O_359,N_14850,N_14553);
or UO_360 (O_360,N_14897,N_14802);
or UO_361 (O_361,N_14695,N_14932);
nand UO_362 (O_362,N_14552,N_14730);
xor UO_363 (O_363,N_14778,N_14970);
nand UO_364 (O_364,N_14913,N_14536);
and UO_365 (O_365,N_14809,N_14988);
nand UO_366 (O_366,N_14567,N_14916);
or UO_367 (O_367,N_14795,N_14778);
or UO_368 (O_368,N_14668,N_14515);
and UO_369 (O_369,N_14537,N_14554);
and UO_370 (O_370,N_14768,N_14675);
and UO_371 (O_371,N_14588,N_14820);
nor UO_372 (O_372,N_14681,N_14590);
or UO_373 (O_373,N_14949,N_14741);
or UO_374 (O_374,N_14605,N_14651);
nand UO_375 (O_375,N_14720,N_14680);
xnor UO_376 (O_376,N_14885,N_14634);
or UO_377 (O_377,N_14927,N_14614);
nand UO_378 (O_378,N_14851,N_14841);
and UO_379 (O_379,N_14775,N_14515);
xnor UO_380 (O_380,N_14834,N_14895);
nor UO_381 (O_381,N_14881,N_14954);
xor UO_382 (O_382,N_14900,N_14573);
nand UO_383 (O_383,N_14539,N_14986);
nor UO_384 (O_384,N_14650,N_14887);
or UO_385 (O_385,N_14516,N_14941);
nor UO_386 (O_386,N_14968,N_14751);
nor UO_387 (O_387,N_14904,N_14924);
nand UO_388 (O_388,N_14893,N_14916);
nor UO_389 (O_389,N_14552,N_14997);
or UO_390 (O_390,N_14630,N_14658);
and UO_391 (O_391,N_14609,N_14697);
xnor UO_392 (O_392,N_14852,N_14955);
xor UO_393 (O_393,N_14640,N_14854);
and UO_394 (O_394,N_14825,N_14864);
xor UO_395 (O_395,N_14875,N_14771);
or UO_396 (O_396,N_14546,N_14692);
or UO_397 (O_397,N_14963,N_14628);
nand UO_398 (O_398,N_14689,N_14849);
nand UO_399 (O_399,N_14973,N_14649);
xor UO_400 (O_400,N_14773,N_14771);
and UO_401 (O_401,N_14701,N_14851);
and UO_402 (O_402,N_14670,N_14892);
nor UO_403 (O_403,N_14815,N_14645);
and UO_404 (O_404,N_14973,N_14900);
xnor UO_405 (O_405,N_14817,N_14974);
or UO_406 (O_406,N_14754,N_14691);
nor UO_407 (O_407,N_14672,N_14648);
xor UO_408 (O_408,N_14795,N_14929);
xor UO_409 (O_409,N_14742,N_14960);
nor UO_410 (O_410,N_14873,N_14960);
nor UO_411 (O_411,N_14745,N_14905);
xor UO_412 (O_412,N_14941,N_14710);
xor UO_413 (O_413,N_14744,N_14962);
xnor UO_414 (O_414,N_14725,N_14985);
xnor UO_415 (O_415,N_14532,N_14652);
and UO_416 (O_416,N_14958,N_14568);
nand UO_417 (O_417,N_14977,N_14836);
xor UO_418 (O_418,N_14993,N_14904);
nor UO_419 (O_419,N_14936,N_14676);
nor UO_420 (O_420,N_14838,N_14819);
or UO_421 (O_421,N_14598,N_14960);
xnor UO_422 (O_422,N_14869,N_14893);
nor UO_423 (O_423,N_14779,N_14739);
and UO_424 (O_424,N_14720,N_14803);
nor UO_425 (O_425,N_14602,N_14548);
xnor UO_426 (O_426,N_14656,N_14904);
or UO_427 (O_427,N_14543,N_14980);
nand UO_428 (O_428,N_14544,N_14629);
nand UO_429 (O_429,N_14823,N_14872);
and UO_430 (O_430,N_14668,N_14921);
and UO_431 (O_431,N_14810,N_14956);
nor UO_432 (O_432,N_14744,N_14674);
nand UO_433 (O_433,N_14974,N_14675);
nand UO_434 (O_434,N_14902,N_14657);
or UO_435 (O_435,N_14789,N_14775);
nand UO_436 (O_436,N_14879,N_14778);
nand UO_437 (O_437,N_14515,N_14901);
nor UO_438 (O_438,N_14591,N_14695);
nand UO_439 (O_439,N_14764,N_14802);
nor UO_440 (O_440,N_14894,N_14709);
or UO_441 (O_441,N_14849,N_14550);
nor UO_442 (O_442,N_14755,N_14721);
xor UO_443 (O_443,N_14590,N_14956);
nand UO_444 (O_444,N_14559,N_14803);
and UO_445 (O_445,N_14762,N_14904);
or UO_446 (O_446,N_14959,N_14896);
nand UO_447 (O_447,N_14982,N_14742);
nor UO_448 (O_448,N_14886,N_14722);
or UO_449 (O_449,N_14718,N_14846);
or UO_450 (O_450,N_14899,N_14570);
or UO_451 (O_451,N_14578,N_14793);
nand UO_452 (O_452,N_14678,N_14868);
xnor UO_453 (O_453,N_14753,N_14920);
or UO_454 (O_454,N_14716,N_14839);
and UO_455 (O_455,N_14822,N_14527);
or UO_456 (O_456,N_14533,N_14802);
nand UO_457 (O_457,N_14603,N_14870);
xnor UO_458 (O_458,N_14591,N_14511);
and UO_459 (O_459,N_14629,N_14810);
or UO_460 (O_460,N_14923,N_14536);
nand UO_461 (O_461,N_14734,N_14652);
or UO_462 (O_462,N_14847,N_14896);
nor UO_463 (O_463,N_14561,N_14589);
nand UO_464 (O_464,N_14909,N_14854);
nor UO_465 (O_465,N_14569,N_14576);
or UO_466 (O_466,N_14673,N_14834);
or UO_467 (O_467,N_14876,N_14997);
xnor UO_468 (O_468,N_14923,N_14702);
xor UO_469 (O_469,N_14910,N_14593);
or UO_470 (O_470,N_14885,N_14615);
or UO_471 (O_471,N_14765,N_14725);
nor UO_472 (O_472,N_14895,N_14771);
xnor UO_473 (O_473,N_14998,N_14988);
nand UO_474 (O_474,N_14711,N_14833);
xor UO_475 (O_475,N_14891,N_14568);
and UO_476 (O_476,N_14963,N_14759);
nand UO_477 (O_477,N_14541,N_14921);
xnor UO_478 (O_478,N_14822,N_14786);
and UO_479 (O_479,N_14930,N_14755);
nor UO_480 (O_480,N_14568,N_14964);
xnor UO_481 (O_481,N_14753,N_14679);
xor UO_482 (O_482,N_14698,N_14708);
nand UO_483 (O_483,N_14520,N_14665);
or UO_484 (O_484,N_14885,N_14824);
and UO_485 (O_485,N_14783,N_14765);
nand UO_486 (O_486,N_14576,N_14894);
nand UO_487 (O_487,N_14678,N_14776);
nor UO_488 (O_488,N_14850,N_14710);
nor UO_489 (O_489,N_14726,N_14828);
or UO_490 (O_490,N_14863,N_14929);
xnor UO_491 (O_491,N_14519,N_14830);
nand UO_492 (O_492,N_14742,N_14702);
and UO_493 (O_493,N_14768,N_14869);
and UO_494 (O_494,N_14984,N_14904);
nand UO_495 (O_495,N_14655,N_14700);
xnor UO_496 (O_496,N_14609,N_14940);
nand UO_497 (O_497,N_14690,N_14882);
nor UO_498 (O_498,N_14939,N_14710);
nand UO_499 (O_499,N_14799,N_14635);
xnor UO_500 (O_500,N_14794,N_14988);
nor UO_501 (O_501,N_14828,N_14936);
nor UO_502 (O_502,N_14562,N_14755);
nand UO_503 (O_503,N_14954,N_14537);
nand UO_504 (O_504,N_14716,N_14588);
nand UO_505 (O_505,N_14773,N_14827);
and UO_506 (O_506,N_14969,N_14533);
and UO_507 (O_507,N_14724,N_14924);
or UO_508 (O_508,N_14837,N_14907);
and UO_509 (O_509,N_14988,N_14927);
nand UO_510 (O_510,N_14851,N_14644);
or UO_511 (O_511,N_14711,N_14631);
xnor UO_512 (O_512,N_14690,N_14634);
nor UO_513 (O_513,N_14797,N_14584);
and UO_514 (O_514,N_14688,N_14947);
or UO_515 (O_515,N_14980,N_14797);
nand UO_516 (O_516,N_14814,N_14686);
and UO_517 (O_517,N_14622,N_14577);
or UO_518 (O_518,N_14770,N_14554);
nand UO_519 (O_519,N_14879,N_14745);
nand UO_520 (O_520,N_14642,N_14748);
or UO_521 (O_521,N_14595,N_14728);
xnor UO_522 (O_522,N_14567,N_14775);
and UO_523 (O_523,N_14765,N_14892);
nor UO_524 (O_524,N_14752,N_14639);
nor UO_525 (O_525,N_14512,N_14824);
nor UO_526 (O_526,N_14893,N_14662);
and UO_527 (O_527,N_14762,N_14582);
or UO_528 (O_528,N_14665,N_14587);
or UO_529 (O_529,N_14547,N_14997);
nor UO_530 (O_530,N_14538,N_14785);
xnor UO_531 (O_531,N_14856,N_14833);
and UO_532 (O_532,N_14930,N_14949);
and UO_533 (O_533,N_14725,N_14830);
or UO_534 (O_534,N_14934,N_14618);
nand UO_535 (O_535,N_14600,N_14906);
nand UO_536 (O_536,N_14641,N_14740);
nand UO_537 (O_537,N_14522,N_14975);
nor UO_538 (O_538,N_14845,N_14880);
xnor UO_539 (O_539,N_14866,N_14939);
or UO_540 (O_540,N_14664,N_14773);
or UO_541 (O_541,N_14659,N_14786);
and UO_542 (O_542,N_14910,N_14523);
and UO_543 (O_543,N_14622,N_14914);
and UO_544 (O_544,N_14904,N_14502);
or UO_545 (O_545,N_14725,N_14809);
and UO_546 (O_546,N_14521,N_14576);
nor UO_547 (O_547,N_14534,N_14966);
xor UO_548 (O_548,N_14544,N_14970);
nor UO_549 (O_549,N_14519,N_14594);
nand UO_550 (O_550,N_14843,N_14944);
nor UO_551 (O_551,N_14832,N_14973);
nand UO_552 (O_552,N_14863,N_14956);
nor UO_553 (O_553,N_14753,N_14636);
and UO_554 (O_554,N_14788,N_14555);
nand UO_555 (O_555,N_14678,N_14755);
xor UO_556 (O_556,N_14765,N_14966);
xnor UO_557 (O_557,N_14697,N_14718);
nand UO_558 (O_558,N_14683,N_14746);
nand UO_559 (O_559,N_14960,N_14782);
xor UO_560 (O_560,N_14577,N_14541);
nand UO_561 (O_561,N_14757,N_14550);
and UO_562 (O_562,N_14570,N_14893);
and UO_563 (O_563,N_14939,N_14884);
or UO_564 (O_564,N_14954,N_14601);
xnor UO_565 (O_565,N_14819,N_14679);
or UO_566 (O_566,N_14866,N_14519);
nand UO_567 (O_567,N_14696,N_14668);
nand UO_568 (O_568,N_14558,N_14682);
nand UO_569 (O_569,N_14727,N_14744);
xnor UO_570 (O_570,N_14699,N_14848);
xnor UO_571 (O_571,N_14928,N_14684);
or UO_572 (O_572,N_14572,N_14535);
nand UO_573 (O_573,N_14667,N_14805);
xnor UO_574 (O_574,N_14713,N_14952);
xnor UO_575 (O_575,N_14989,N_14547);
nor UO_576 (O_576,N_14615,N_14896);
nand UO_577 (O_577,N_14718,N_14814);
and UO_578 (O_578,N_14938,N_14590);
xnor UO_579 (O_579,N_14655,N_14783);
xnor UO_580 (O_580,N_14993,N_14894);
nand UO_581 (O_581,N_14508,N_14521);
nor UO_582 (O_582,N_14643,N_14979);
nand UO_583 (O_583,N_14950,N_14997);
nand UO_584 (O_584,N_14876,N_14639);
or UO_585 (O_585,N_14812,N_14682);
xnor UO_586 (O_586,N_14596,N_14851);
xor UO_587 (O_587,N_14914,N_14739);
or UO_588 (O_588,N_14964,N_14743);
xnor UO_589 (O_589,N_14936,N_14765);
and UO_590 (O_590,N_14773,N_14943);
or UO_591 (O_591,N_14812,N_14954);
nand UO_592 (O_592,N_14962,N_14976);
xor UO_593 (O_593,N_14676,N_14688);
xnor UO_594 (O_594,N_14910,N_14559);
nor UO_595 (O_595,N_14788,N_14739);
or UO_596 (O_596,N_14563,N_14956);
and UO_597 (O_597,N_14846,N_14705);
xor UO_598 (O_598,N_14684,N_14979);
nand UO_599 (O_599,N_14934,N_14812);
nor UO_600 (O_600,N_14685,N_14885);
nand UO_601 (O_601,N_14668,N_14692);
nor UO_602 (O_602,N_14880,N_14821);
nand UO_603 (O_603,N_14651,N_14997);
or UO_604 (O_604,N_14689,N_14898);
and UO_605 (O_605,N_14989,N_14895);
or UO_606 (O_606,N_14884,N_14590);
and UO_607 (O_607,N_14718,N_14845);
or UO_608 (O_608,N_14702,N_14966);
nand UO_609 (O_609,N_14870,N_14817);
nor UO_610 (O_610,N_14893,N_14741);
or UO_611 (O_611,N_14519,N_14574);
xor UO_612 (O_612,N_14560,N_14642);
nor UO_613 (O_613,N_14799,N_14537);
nand UO_614 (O_614,N_14836,N_14769);
nor UO_615 (O_615,N_14898,N_14780);
nor UO_616 (O_616,N_14723,N_14682);
and UO_617 (O_617,N_14747,N_14623);
nand UO_618 (O_618,N_14831,N_14922);
or UO_619 (O_619,N_14989,N_14697);
and UO_620 (O_620,N_14653,N_14770);
xor UO_621 (O_621,N_14515,N_14503);
nand UO_622 (O_622,N_14844,N_14903);
nor UO_623 (O_623,N_14602,N_14518);
or UO_624 (O_624,N_14652,N_14581);
or UO_625 (O_625,N_14764,N_14677);
and UO_626 (O_626,N_14795,N_14639);
xor UO_627 (O_627,N_14717,N_14817);
or UO_628 (O_628,N_14707,N_14884);
xnor UO_629 (O_629,N_14774,N_14856);
and UO_630 (O_630,N_14824,N_14693);
nand UO_631 (O_631,N_14782,N_14784);
xnor UO_632 (O_632,N_14718,N_14736);
nor UO_633 (O_633,N_14514,N_14944);
and UO_634 (O_634,N_14990,N_14602);
nand UO_635 (O_635,N_14595,N_14758);
xnor UO_636 (O_636,N_14604,N_14806);
nand UO_637 (O_637,N_14764,N_14566);
or UO_638 (O_638,N_14961,N_14907);
nor UO_639 (O_639,N_14690,N_14545);
xnor UO_640 (O_640,N_14528,N_14963);
and UO_641 (O_641,N_14588,N_14571);
nor UO_642 (O_642,N_14515,N_14915);
nor UO_643 (O_643,N_14673,N_14531);
and UO_644 (O_644,N_14651,N_14885);
nand UO_645 (O_645,N_14588,N_14856);
xnor UO_646 (O_646,N_14920,N_14988);
nand UO_647 (O_647,N_14893,N_14813);
and UO_648 (O_648,N_14883,N_14738);
and UO_649 (O_649,N_14586,N_14698);
and UO_650 (O_650,N_14530,N_14752);
nand UO_651 (O_651,N_14597,N_14940);
xor UO_652 (O_652,N_14734,N_14541);
and UO_653 (O_653,N_14665,N_14987);
or UO_654 (O_654,N_14977,N_14848);
nor UO_655 (O_655,N_14750,N_14891);
and UO_656 (O_656,N_14608,N_14912);
and UO_657 (O_657,N_14723,N_14605);
xor UO_658 (O_658,N_14873,N_14640);
nor UO_659 (O_659,N_14914,N_14510);
and UO_660 (O_660,N_14711,N_14748);
xor UO_661 (O_661,N_14621,N_14796);
nor UO_662 (O_662,N_14709,N_14913);
nor UO_663 (O_663,N_14752,N_14869);
nor UO_664 (O_664,N_14655,N_14880);
xor UO_665 (O_665,N_14547,N_14572);
or UO_666 (O_666,N_14513,N_14789);
xor UO_667 (O_667,N_14605,N_14642);
nor UO_668 (O_668,N_14845,N_14827);
and UO_669 (O_669,N_14791,N_14749);
or UO_670 (O_670,N_14840,N_14950);
nand UO_671 (O_671,N_14608,N_14867);
and UO_672 (O_672,N_14510,N_14601);
nand UO_673 (O_673,N_14985,N_14829);
or UO_674 (O_674,N_14997,N_14931);
nand UO_675 (O_675,N_14659,N_14778);
nand UO_676 (O_676,N_14867,N_14928);
and UO_677 (O_677,N_14724,N_14650);
and UO_678 (O_678,N_14866,N_14632);
nand UO_679 (O_679,N_14861,N_14955);
nand UO_680 (O_680,N_14624,N_14608);
and UO_681 (O_681,N_14732,N_14592);
or UO_682 (O_682,N_14857,N_14745);
xor UO_683 (O_683,N_14928,N_14650);
nand UO_684 (O_684,N_14563,N_14927);
or UO_685 (O_685,N_14628,N_14847);
and UO_686 (O_686,N_14523,N_14500);
nor UO_687 (O_687,N_14902,N_14971);
nand UO_688 (O_688,N_14592,N_14789);
xor UO_689 (O_689,N_14562,N_14974);
nand UO_690 (O_690,N_14752,N_14862);
xnor UO_691 (O_691,N_14744,N_14683);
and UO_692 (O_692,N_14801,N_14637);
xnor UO_693 (O_693,N_14637,N_14566);
xor UO_694 (O_694,N_14723,N_14706);
nand UO_695 (O_695,N_14709,N_14692);
nor UO_696 (O_696,N_14737,N_14664);
nand UO_697 (O_697,N_14948,N_14547);
and UO_698 (O_698,N_14577,N_14652);
and UO_699 (O_699,N_14616,N_14668);
xor UO_700 (O_700,N_14600,N_14992);
nor UO_701 (O_701,N_14691,N_14937);
xor UO_702 (O_702,N_14687,N_14800);
and UO_703 (O_703,N_14848,N_14992);
xor UO_704 (O_704,N_14611,N_14753);
or UO_705 (O_705,N_14845,N_14858);
or UO_706 (O_706,N_14586,N_14795);
and UO_707 (O_707,N_14572,N_14954);
nand UO_708 (O_708,N_14578,N_14571);
and UO_709 (O_709,N_14921,N_14768);
or UO_710 (O_710,N_14646,N_14688);
xnor UO_711 (O_711,N_14725,N_14640);
nor UO_712 (O_712,N_14770,N_14546);
or UO_713 (O_713,N_14743,N_14969);
or UO_714 (O_714,N_14699,N_14647);
nand UO_715 (O_715,N_14800,N_14907);
nor UO_716 (O_716,N_14777,N_14917);
nand UO_717 (O_717,N_14691,N_14706);
nor UO_718 (O_718,N_14715,N_14883);
and UO_719 (O_719,N_14875,N_14944);
and UO_720 (O_720,N_14852,N_14646);
xnor UO_721 (O_721,N_14804,N_14675);
xor UO_722 (O_722,N_14929,N_14770);
and UO_723 (O_723,N_14733,N_14746);
nand UO_724 (O_724,N_14537,N_14944);
or UO_725 (O_725,N_14867,N_14864);
xnor UO_726 (O_726,N_14638,N_14801);
xnor UO_727 (O_727,N_14506,N_14617);
nand UO_728 (O_728,N_14854,N_14704);
nor UO_729 (O_729,N_14625,N_14998);
nor UO_730 (O_730,N_14979,N_14965);
nor UO_731 (O_731,N_14871,N_14765);
nor UO_732 (O_732,N_14953,N_14544);
nand UO_733 (O_733,N_14755,N_14821);
and UO_734 (O_734,N_14556,N_14597);
nand UO_735 (O_735,N_14598,N_14855);
and UO_736 (O_736,N_14770,N_14797);
nor UO_737 (O_737,N_14743,N_14778);
nor UO_738 (O_738,N_14939,N_14834);
and UO_739 (O_739,N_14990,N_14852);
nor UO_740 (O_740,N_14540,N_14830);
nand UO_741 (O_741,N_14965,N_14880);
nand UO_742 (O_742,N_14912,N_14817);
and UO_743 (O_743,N_14863,N_14786);
xor UO_744 (O_744,N_14874,N_14861);
nor UO_745 (O_745,N_14989,N_14529);
nand UO_746 (O_746,N_14553,N_14851);
nor UO_747 (O_747,N_14625,N_14565);
and UO_748 (O_748,N_14805,N_14679);
or UO_749 (O_749,N_14598,N_14883);
or UO_750 (O_750,N_14854,N_14901);
nor UO_751 (O_751,N_14829,N_14825);
and UO_752 (O_752,N_14783,N_14820);
or UO_753 (O_753,N_14946,N_14820);
xor UO_754 (O_754,N_14978,N_14761);
xor UO_755 (O_755,N_14620,N_14648);
or UO_756 (O_756,N_14517,N_14693);
or UO_757 (O_757,N_14940,N_14678);
xnor UO_758 (O_758,N_14676,N_14528);
nand UO_759 (O_759,N_14912,N_14735);
xor UO_760 (O_760,N_14969,N_14959);
and UO_761 (O_761,N_14911,N_14739);
and UO_762 (O_762,N_14998,N_14795);
xor UO_763 (O_763,N_14735,N_14785);
nand UO_764 (O_764,N_14997,N_14864);
xor UO_765 (O_765,N_14549,N_14994);
or UO_766 (O_766,N_14818,N_14624);
or UO_767 (O_767,N_14610,N_14607);
nand UO_768 (O_768,N_14794,N_14986);
nand UO_769 (O_769,N_14614,N_14605);
nor UO_770 (O_770,N_14931,N_14516);
xnor UO_771 (O_771,N_14996,N_14840);
nand UO_772 (O_772,N_14561,N_14580);
or UO_773 (O_773,N_14569,N_14552);
xor UO_774 (O_774,N_14812,N_14849);
xnor UO_775 (O_775,N_14783,N_14888);
xor UO_776 (O_776,N_14890,N_14541);
nor UO_777 (O_777,N_14690,N_14792);
nand UO_778 (O_778,N_14824,N_14988);
nor UO_779 (O_779,N_14752,N_14886);
nand UO_780 (O_780,N_14873,N_14504);
or UO_781 (O_781,N_14793,N_14687);
and UO_782 (O_782,N_14704,N_14766);
xnor UO_783 (O_783,N_14890,N_14747);
nor UO_784 (O_784,N_14537,N_14628);
nor UO_785 (O_785,N_14884,N_14929);
nor UO_786 (O_786,N_14511,N_14806);
or UO_787 (O_787,N_14994,N_14910);
xor UO_788 (O_788,N_14748,N_14638);
xor UO_789 (O_789,N_14699,N_14582);
xor UO_790 (O_790,N_14886,N_14718);
xor UO_791 (O_791,N_14570,N_14728);
nor UO_792 (O_792,N_14597,N_14732);
or UO_793 (O_793,N_14862,N_14511);
or UO_794 (O_794,N_14656,N_14785);
nand UO_795 (O_795,N_14712,N_14659);
and UO_796 (O_796,N_14653,N_14661);
and UO_797 (O_797,N_14755,N_14578);
and UO_798 (O_798,N_14908,N_14954);
xor UO_799 (O_799,N_14570,N_14729);
or UO_800 (O_800,N_14772,N_14666);
or UO_801 (O_801,N_14832,N_14612);
nand UO_802 (O_802,N_14729,N_14900);
xor UO_803 (O_803,N_14999,N_14959);
and UO_804 (O_804,N_14731,N_14527);
and UO_805 (O_805,N_14503,N_14550);
and UO_806 (O_806,N_14927,N_14684);
or UO_807 (O_807,N_14854,N_14590);
and UO_808 (O_808,N_14978,N_14896);
or UO_809 (O_809,N_14612,N_14509);
nand UO_810 (O_810,N_14909,N_14503);
xor UO_811 (O_811,N_14632,N_14803);
nor UO_812 (O_812,N_14808,N_14516);
or UO_813 (O_813,N_14780,N_14952);
or UO_814 (O_814,N_14991,N_14568);
xnor UO_815 (O_815,N_14858,N_14944);
nand UO_816 (O_816,N_14633,N_14942);
xor UO_817 (O_817,N_14755,N_14862);
nor UO_818 (O_818,N_14743,N_14838);
nor UO_819 (O_819,N_14561,N_14730);
nor UO_820 (O_820,N_14687,N_14594);
nand UO_821 (O_821,N_14857,N_14582);
or UO_822 (O_822,N_14993,N_14803);
xnor UO_823 (O_823,N_14851,N_14689);
nor UO_824 (O_824,N_14712,N_14548);
and UO_825 (O_825,N_14962,N_14748);
xor UO_826 (O_826,N_14978,N_14721);
xor UO_827 (O_827,N_14857,N_14547);
xor UO_828 (O_828,N_14878,N_14746);
and UO_829 (O_829,N_14506,N_14853);
nor UO_830 (O_830,N_14545,N_14525);
xor UO_831 (O_831,N_14739,N_14866);
xor UO_832 (O_832,N_14779,N_14927);
nand UO_833 (O_833,N_14778,N_14690);
or UO_834 (O_834,N_14971,N_14802);
nor UO_835 (O_835,N_14881,N_14840);
or UO_836 (O_836,N_14559,N_14885);
xor UO_837 (O_837,N_14844,N_14886);
nor UO_838 (O_838,N_14804,N_14659);
xnor UO_839 (O_839,N_14764,N_14646);
or UO_840 (O_840,N_14981,N_14730);
and UO_841 (O_841,N_14735,N_14978);
nand UO_842 (O_842,N_14609,N_14704);
nor UO_843 (O_843,N_14528,N_14911);
nand UO_844 (O_844,N_14659,N_14706);
nand UO_845 (O_845,N_14577,N_14988);
or UO_846 (O_846,N_14863,N_14800);
and UO_847 (O_847,N_14901,N_14570);
nand UO_848 (O_848,N_14520,N_14702);
nor UO_849 (O_849,N_14936,N_14859);
or UO_850 (O_850,N_14619,N_14665);
xor UO_851 (O_851,N_14718,N_14896);
or UO_852 (O_852,N_14968,N_14881);
nor UO_853 (O_853,N_14566,N_14956);
or UO_854 (O_854,N_14501,N_14807);
nand UO_855 (O_855,N_14734,N_14581);
nand UO_856 (O_856,N_14527,N_14753);
or UO_857 (O_857,N_14885,N_14544);
xnor UO_858 (O_858,N_14773,N_14624);
nand UO_859 (O_859,N_14555,N_14989);
nor UO_860 (O_860,N_14612,N_14574);
xor UO_861 (O_861,N_14508,N_14681);
xnor UO_862 (O_862,N_14657,N_14585);
xor UO_863 (O_863,N_14753,N_14592);
and UO_864 (O_864,N_14618,N_14611);
and UO_865 (O_865,N_14578,N_14739);
nor UO_866 (O_866,N_14816,N_14518);
or UO_867 (O_867,N_14632,N_14604);
nand UO_868 (O_868,N_14529,N_14648);
xor UO_869 (O_869,N_14723,N_14527);
and UO_870 (O_870,N_14861,N_14792);
or UO_871 (O_871,N_14892,N_14648);
nand UO_872 (O_872,N_14731,N_14828);
or UO_873 (O_873,N_14776,N_14582);
and UO_874 (O_874,N_14761,N_14725);
and UO_875 (O_875,N_14552,N_14506);
xnor UO_876 (O_876,N_14517,N_14592);
nor UO_877 (O_877,N_14602,N_14555);
nor UO_878 (O_878,N_14702,N_14917);
and UO_879 (O_879,N_14833,N_14510);
nand UO_880 (O_880,N_14533,N_14890);
xnor UO_881 (O_881,N_14666,N_14631);
and UO_882 (O_882,N_14952,N_14933);
nand UO_883 (O_883,N_14784,N_14885);
xor UO_884 (O_884,N_14602,N_14523);
or UO_885 (O_885,N_14866,N_14738);
or UO_886 (O_886,N_14880,N_14721);
nand UO_887 (O_887,N_14642,N_14879);
and UO_888 (O_888,N_14997,N_14605);
or UO_889 (O_889,N_14640,N_14968);
xor UO_890 (O_890,N_14874,N_14967);
nand UO_891 (O_891,N_14897,N_14796);
xor UO_892 (O_892,N_14580,N_14704);
xnor UO_893 (O_893,N_14985,N_14699);
nand UO_894 (O_894,N_14518,N_14800);
and UO_895 (O_895,N_14532,N_14968);
or UO_896 (O_896,N_14653,N_14815);
nand UO_897 (O_897,N_14546,N_14907);
and UO_898 (O_898,N_14715,N_14737);
xor UO_899 (O_899,N_14665,N_14692);
or UO_900 (O_900,N_14707,N_14764);
nand UO_901 (O_901,N_14949,N_14746);
or UO_902 (O_902,N_14547,N_14623);
xnor UO_903 (O_903,N_14812,N_14732);
and UO_904 (O_904,N_14828,N_14718);
and UO_905 (O_905,N_14592,N_14809);
and UO_906 (O_906,N_14605,N_14978);
nor UO_907 (O_907,N_14769,N_14729);
nor UO_908 (O_908,N_14615,N_14985);
and UO_909 (O_909,N_14987,N_14674);
nand UO_910 (O_910,N_14941,N_14942);
nand UO_911 (O_911,N_14688,N_14605);
nand UO_912 (O_912,N_14619,N_14630);
nor UO_913 (O_913,N_14728,N_14614);
or UO_914 (O_914,N_14865,N_14758);
nor UO_915 (O_915,N_14897,N_14815);
and UO_916 (O_916,N_14837,N_14703);
or UO_917 (O_917,N_14553,N_14830);
xor UO_918 (O_918,N_14804,N_14504);
or UO_919 (O_919,N_14783,N_14588);
xnor UO_920 (O_920,N_14970,N_14744);
or UO_921 (O_921,N_14744,N_14614);
nand UO_922 (O_922,N_14767,N_14692);
and UO_923 (O_923,N_14576,N_14909);
nor UO_924 (O_924,N_14939,N_14854);
xor UO_925 (O_925,N_14970,N_14859);
nand UO_926 (O_926,N_14610,N_14810);
and UO_927 (O_927,N_14956,N_14984);
nand UO_928 (O_928,N_14725,N_14531);
xor UO_929 (O_929,N_14834,N_14564);
or UO_930 (O_930,N_14539,N_14639);
nor UO_931 (O_931,N_14805,N_14946);
nor UO_932 (O_932,N_14814,N_14689);
nor UO_933 (O_933,N_14945,N_14717);
nor UO_934 (O_934,N_14521,N_14976);
nor UO_935 (O_935,N_14569,N_14895);
nand UO_936 (O_936,N_14635,N_14577);
nand UO_937 (O_937,N_14878,N_14685);
nand UO_938 (O_938,N_14604,N_14571);
and UO_939 (O_939,N_14525,N_14846);
nor UO_940 (O_940,N_14682,N_14849);
nor UO_941 (O_941,N_14883,N_14718);
or UO_942 (O_942,N_14686,N_14545);
nor UO_943 (O_943,N_14939,N_14837);
and UO_944 (O_944,N_14743,N_14649);
xnor UO_945 (O_945,N_14770,N_14705);
xnor UO_946 (O_946,N_14921,N_14908);
nand UO_947 (O_947,N_14551,N_14693);
and UO_948 (O_948,N_14981,N_14618);
xor UO_949 (O_949,N_14972,N_14932);
nor UO_950 (O_950,N_14968,N_14550);
nor UO_951 (O_951,N_14769,N_14964);
or UO_952 (O_952,N_14899,N_14585);
xnor UO_953 (O_953,N_14822,N_14757);
nand UO_954 (O_954,N_14707,N_14877);
nand UO_955 (O_955,N_14777,N_14900);
or UO_956 (O_956,N_14558,N_14881);
xnor UO_957 (O_957,N_14885,N_14748);
or UO_958 (O_958,N_14674,N_14995);
and UO_959 (O_959,N_14730,N_14570);
xor UO_960 (O_960,N_14915,N_14652);
nand UO_961 (O_961,N_14557,N_14989);
xor UO_962 (O_962,N_14746,N_14739);
or UO_963 (O_963,N_14816,N_14978);
nand UO_964 (O_964,N_14995,N_14990);
xor UO_965 (O_965,N_14604,N_14865);
xor UO_966 (O_966,N_14673,N_14915);
and UO_967 (O_967,N_14556,N_14944);
xor UO_968 (O_968,N_14998,N_14516);
and UO_969 (O_969,N_14515,N_14847);
xnor UO_970 (O_970,N_14782,N_14977);
and UO_971 (O_971,N_14598,N_14932);
nand UO_972 (O_972,N_14853,N_14666);
xor UO_973 (O_973,N_14597,N_14588);
nor UO_974 (O_974,N_14728,N_14529);
nor UO_975 (O_975,N_14543,N_14746);
or UO_976 (O_976,N_14677,N_14980);
xor UO_977 (O_977,N_14759,N_14804);
and UO_978 (O_978,N_14959,N_14592);
and UO_979 (O_979,N_14855,N_14970);
and UO_980 (O_980,N_14881,N_14742);
nor UO_981 (O_981,N_14570,N_14681);
and UO_982 (O_982,N_14555,N_14600);
or UO_983 (O_983,N_14906,N_14805);
and UO_984 (O_984,N_14662,N_14509);
and UO_985 (O_985,N_14600,N_14890);
or UO_986 (O_986,N_14885,N_14510);
xnor UO_987 (O_987,N_14801,N_14735);
nor UO_988 (O_988,N_14797,N_14762);
and UO_989 (O_989,N_14914,N_14549);
or UO_990 (O_990,N_14573,N_14877);
xnor UO_991 (O_991,N_14644,N_14911);
and UO_992 (O_992,N_14881,N_14778);
xnor UO_993 (O_993,N_14790,N_14653);
nor UO_994 (O_994,N_14552,N_14819);
nor UO_995 (O_995,N_14833,N_14939);
xor UO_996 (O_996,N_14619,N_14617);
or UO_997 (O_997,N_14796,N_14531);
and UO_998 (O_998,N_14759,N_14732);
nand UO_999 (O_999,N_14770,N_14809);
or UO_1000 (O_1000,N_14838,N_14632);
and UO_1001 (O_1001,N_14866,N_14877);
nand UO_1002 (O_1002,N_14985,N_14750);
and UO_1003 (O_1003,N_14709,N_14706);
nor UO_1004 (O_1004,N_14646,N_14605);
nor UO_1005 (O_1005,N_14598,N_14573);
and UO_1006 (O_1006,N_14956,N_14557);
or UO_1007 (O_1007,N_14743,N_14594);
and UO_1008 (O_1008,N_14624,N_14950);
and UO_1009 (O_1009,N_14781,N_14752);
and UO_1010 (O_1010,N_14789,N_14654);
xor UO_1011 (O_1011,N_14577,N_14884);
nand UO_1012 (O_1012,N_14587,N_14623);
nor UO_1013 (O_1013,N_14773,N_14657);
nand UO_1014 (O_1014,N_14997,N_14779);
nor UO_1015 (O_1015,N_14521,N_14728);
nor UO_1016 (O_1016,N_14535,N_14932);
and UO_1017 (O_1017,N_14679,N_14609);
xnor UO_1018 (O_1018,N_14659,N_14714);
nand UO_1019 (O_1019,N_14960,N_14589);
nor UO_1020 (O_1020,N_14739,N_14732);
nand UO_1021 (O_1021,N_14947,N_14956);
and UO_1022 (O_1022,N_14710,N_14852);
nand UO_1023 (O_1023,N_14611,N_14663);
and UO_1024 (O_1024,N_14500,N_14874);
nand UO_1025 (O_1025,N_14579,N_14515);
xor UO_1026 (O_1026,N_14699,N_14874);
nand UO_1027 (O_1027,N_14800,N_14643);
nand UO_1028 (O_1028,N_14855,N_14820);
or UO_1029 (O_1029,N_14693,N_14563);
or UO_1030 (O_1030,N_14518,N_14724);
or UO_1031 (O_1031,N_14973,N_14537);
and UO_1032 (O_1032,N_14533,N_14636);
and UO_1033 (O_1033,N_14583,N_14626);
or UO_1034 (O_1034,N_14698,N_14863);
xor UO_1035 (O_1035,N_14816,N_14869);
or UO_1036 (O_1036,N_14943,N_14500);
and UO_1037 (O_1037,N_14872,N_14580);
nor UO_1038 (O_1038,N_14917,N_14634);
nand UO_1039 (O_1039,N_14687,N_14846);
and UO_1040 (O_1040,N_14722,N_14837);
nor UO_1041 (O_1041,N_14728,N_14539);
nor UO_1042 (O_1042,N_14947,N_14990);
or UO_1043 (O_1043,N_14897,N_14993);
nor UO_1044 (O_1044,N_14683,N_14688);
and UO_1045 (O_1045,N_14504,N_14950);
and UO_1046 (O_1046,N_14990,N_14770);
nand UO_1047 (O_1047,N_14906,N_14556);
xnor UO_1048 (O_1048,N_14538,N_14504);
nor UO_1049 (O_1049,N_14806,N_14886);
and UO_1050 (O_1050,N_14803,N_14807);
nor UO_1051 (O_1051,N_14646,N_14920);
nor UO_1052 (O_1052,N_14553,N_14595);
nor UO_1053 (O_1053,N_14956,N_14848);
nand UO_1054 (O_1054,N_14764,N_14547);
or UO_1055 (O_1055,N_14603,N_14724);
nor UO_1056 (O_1056,N_14608,N_14524);
or UO_1057 (O_1057,N_14518,N_14810);
and UO_1058 (O_1058,N_14804,N_14746);
and UO_1059 (O_1059,N_14581,N_14551);
nand UO_1060 (O_1060,N_14772,N_14918);
and UO_1061 (O_1061,N_14928,N_14795);
xor UO_1062 (O_1062,N_14517,N_14556);
and UO_1063 (O_1063,N_14535,N_14882);
or UO_1064 (O_1064,N_14822,N_14613);
nand UO_1065 (O_1065,N_14869,N_14712);
nor UO_1066 (O_1066,N_14666,N_14822);
xor UO_1067 (O_1067,N_14712,N_14791);
or UO_1068 (O_1068,N_14900,N_14953);
and UO_1069 (O_1069,N_14921,N_14850);
nand UO_1070 (O_1070,N_14877,N_14701);
and UO_1071 (O_1071,N_14924,N_14721);
xor UO_1072 (O_1072,N_14599,N_14507);
and UO_1073 (O_1073,N_14949,N_14512);
nand UO_1074 (O_1074,N_14940,N_14741);
nor UO_1075 (O_1075,N_14741,N_14618);
xor UO_1076 (O_1076,N_14534,N_14905);
nand UO_1077 (O_1077,N_14964,N_14742);
nor UO_1078 (O_1078,N_14634,N_14812);
nor UO_1079 (O_1079,N_14688,N_14642);
xor UO_1080 (O_1080,N_14842,N_14632);
or UO_1081 (O_1081,N_14668,N_14789);
nand UO_1082 (O_1082,N_14755,N_14780);
or UO_1083 (O_1083,N_14629,N_14927);
and UO_1084 (O_1084,N_14944,N_14833);
xor UO_1085 (O_1085,N_14667,N_14970);
xor UO_1086 (O_1086,N_14639,N_14698);
nand UO_1087 (O_1087,N_14666,N_14820);
or UO_1088 (O_1088,N_14626,N_14690);
xor UO_1089 (O_1089,N_14880,N_14838);
or UO_1090 (O_1090,N_14806,N_14533);
and UO_1091 (O_1091,N_14635,N_14949);
xnor UO_1092 (O_1092,N_14547,N_14944);
xnor UO_1093 (O_1093,N_14615,N_14634);
or UO_1094 (O_1094,N_14839,N_14844);
xnor UO_1095 (O_1095,N_14989,N_14565);
or UO_1096 (O_1096,N_14640,N_14531);
xor UO_1097 (O_1097,N_14711,N_14500);
or UO_1098 (O_1098,N_14786,N_14867);
nand UO_1099 (O_1099,N_14980,N_14637);
or UO_1100 (O_1100,N_14804,N_14699);
xor UO_1101 (O_1101,N_14854,N_14889);
nand UO_1102 (O_1102,N_14661,N_14714);
nand UO_1103 (O_1103,N_14964,N_14628);
xnor UO_1104 (O_1104,N_14650,N_14640);
and UO_1105 (O_1105,N_14504,N_14648);
nand UO_1106 (O_1106,N_14993,N_14824);
nand UO_1107 (O_1107,N_14763,N_14638);
xnor UO_1108 (O_1108,N_14652,N_14712);
nor UO_1109 (O_1109,N_14929,N_14971);
xnor UO_1110 (O_1110,N_14702,N_14822);
nand UO_1111 (O_1111,N_14682,N_14516);
or UO_1112 (O_1112,N_14938,N_14778);
xor UO_1113 (O_1113,N_14526,N_14736);
and UO_1114 (O_1114,N_14612,N_14997);
nor UO_1115 (O_1115,N_14864,N_14992);
or UO_1116 (O_1116,N_14592,N_14548);
or UO_1117 (O_1117,N_14573,N_14956);
xor UO_1118 (O_1118,N_14988,N_14510);
and UO_1119 (O_1119,N_14644,N_14814);
or UO_1120 (O_1120,N_14774,N_14638);
or UO_1121 (O_1121,N_14771,N_14979);
xor UO_1122 (O_1122,N_14558,N_14855);
and UO_1123 (O_1123,N_14505,N_14733);
nor UO_1124 (O_1124,N_14942,N_14792);
nor UO_1125 (O_1125,N_14590,N_14625);
nor UO_1126 (O_1126,N_14818,N_14598);
nor UO_1127 (O_1127,N_14709,N_14829);
nor UO_1128 (O_1128,N_14630,N_14546);
xor UO_1129 (O_1129,N_14637,N_14900);
and UO_1130 (O_1130,N_14828,N_14649);
and UO_1131 (O_1131,N_14780,N_14557);
xnor UO_1132 (O_1132,N_14991,N_14776);
or UO_1133 (O_1133,N_14511,N_14969);
xnor UO_1134 (O_1134,N_14685,N_14536);
or UO_1135 (O_1135,N_14648,N_14972);
nand UO_1136 (O_1136,N_14599,N_14596);
xnor UO_1137 (O_1137,N_14542,N_14559);
nor UO_1138 (O_1138,N_14938,N_14574);
nor UO_1139 (O_1139,N_14916,N_14817);
nor UO_1140 (O_1140,N_14983,N_14595);
nand UO_1141 (O_1141,N_14650,N_14973);
nand UO_1142 (O_1142,N_14596,N_14827);
nor UO_1143 (O_1143,N_14553,N_14662);
nor UO_1144 (O_1144,N_14599,N_14623);
and UO_1145 (O_1145,N_14619,N_14720);
nand UO_1146 (O_1146,N_14513,N_14962);
or UO_1147 (O_1147,N_14719,N_14675);
xnor UO_1148 (O_1148,N_14987,N_14983);
xnor UO_1149 (O_1149,N_14958,N_14638);
nor UO_1150 (O_1150,N_14787,N_14613);
nor UO_1151 (O_1151,N_14928,N_14870);
or UO_1152 (O_1152,N_14959,N_14789);
xor UO_1153 (O_1153,N_14609,N_14948);
or UO_1154 (O_1154,N_14726,N_14765);
nor UO_1155 (O_1155,N_14866,N_14529);
or UO_1156 (O_1156,N_14623,N_14963);
or UO_1157 (O_1157,N_14845,N_14684);
xor UO_1158 (O_1158,N_14558,N_14790);
xor UO_1159 (O_1159,N_14571,N_14980);
or UO_1160 (O_1160,N_14731,N_14563);
nand UO_1161 (O_1161,N_14700,N_14511);
or UO_1162 (O_1162,N_14909,N_14930);
or UO_1163 (O_1163,N_14888,N_14673);
nand UO_1164 (O_1164,N_14605,N_14789);
or UO_1165 (O_1165,N_14543,N_14816);
or UO_1166 (O_1166,N_14899,N_14862);
nand UO_1167 (O_1167,N_14693,N_14593);
or UO_1168 (O_1168,N_14543,N_14512);
nand UO_1169 (O_1169,N_14832,N_14740);
and UO_1170 (O_1170,N_14996,N_14725);
nor UO_1171 (O_1171,N_14853,N_14866);
xor UO_1172 (O_1172,N_14631,N_14572);
nand UO_1173 (O_1173,N_14509,N_14903);
and UO_1174 (O_1174,N_14569,N_14704);
xor UO_1175 (O_1175,N_14521,N_14593);
and UO_1176 (O_1176,N_14999,N_14846);
xnor UO_1177 (O_1177,N_14831,N_14907);
nor UO_1178 (O_1178,N_14606,N_14903);
nand UO_1179 (O_1179,N_14958,N_14580);
or UO_1180 (O_1180,N_14634,N_14880);
nor UO_1181 (O_1181,N_14824,N_14960);
and UO_1182 (O_1182,N_14864,N_14573);
or UO_1183 (O_1183,N_14659,N_14989);
nand UO_1184 (O_1184,N_14557,N_14584);
xnor UO_1185 (O_1185,N_14559,N_14646);
and UO_1186 (O_1186,N_14998,N_14818);
and UO_1187 (O_1187,N_14663,N_14735);
or UO_1188 (O_1188,N_14541,N_14790);
xnor UO_1189 (O_1189,N_14739,N_14838);
nor UO_1190 (O_1190,N_14960,N_14987);
nand UO_1191 (O_1191,N_14522,N_14627);
and UO_1192 (O_1192,N_14925,N_14577);
xnor UO_1193 (O_1193,N_14749,N_14640);
nor UO_1194 (O_1194,N_14755,N_14684);
nand UO_1195 (O_1195,N_14893,N_14633);
and UO_1196 (O_1196,N_14518,N_14988);
or UO_1197 (O_1197,N_14662,N_14554);
and UO_1198 (O_1198,N_14943,N_14853);
or UO_1199 (O_1199,N_14806,N_14816);
and UO_1200 (O_1200,N_14588,N_14503);
and UO_1201 (O_1201,N_14742,N_14790);
nand UO_1202 (O_1202,N_14910,N_14594);
xnor UO_1203 (O_1203,N_14682,N_14673);
nor UO_1204 (O_1204,N_14585,N_14518);
xor UO_1205 (O_1205,N_14656,N_14982);
or UO_1206 (O_1206,N_14782,N_14866);
xor UO_1207 (O_1207,N_14534,N_14790);
nand UO_1208 (O_1208,N_14937,N_14731);
nor UO_1209 (O_1209,N_14900,N_14706);
and UO_1210 (O_1210,N_14752,N_14797);
nor UO_1211 (O_1211,N_14735,N_14778);
xor UO_1212 (O_1212,N_14761,N_14977);
xnor UO_1213 (O_1213,N_14603,N_14542);
nand UO_1214 (O_1214,N_14745,N_14724);
or UO_1215 (O_1215,N_14714,N_14750);
or UO_1216 (O_1216,N_14501,N_14684);
nand UO_1217 (O_1217,N_14827,N_14657);
nand UO_1218 (O_1218,N_14978,N_14825);
and UO_1219 (O_1219,N_14947,N_14579);
or UO_1220 (O_1220,N_14822,N_14874);
xor UO_1221 (O_1221,N_14632,N_14881);
nand UO_1222 (O_1222,N_14782,N_14827);
nor UO_1223 (O_1223,N_14553,N_14895);
or UO_1224 (O_1224,N_14764,N_14560);
xnor UO_1225 (O_1225,N_14601,N_14864);
xnor UO_1226 (O_1226,N_14523,N_14614);
nor UO_1227 (O_1227,N_14668,N_14953);
or UO_1228 (O_1228,N_14963,N_14632);
xnor UO_1229 (O_1229,N_14943,N_14640);
xnor UO_1230 (O_1230,N_14703,N_14810);
or UO_1231 (O_1231,N_14657,N_14975);
and UO_1232 (O_1232,N_14796,N_14538);
nor UO_1233 (O_1233,N_14522,N_14819);
nor UO_1234 (O_1234,N_14881,N_14683);
xor UO_1235 (O_1235,N_14553,N_14706);
and UO_1236 (O_1236,N_14861,N_14990);
xnor UO_1237 (O_1237,N_14558,N_14828);
or UO_1238 (O_1238,N_14589,N_14895);
and UO_1239 (O_1239,N_14657,N_14837);
nand UO_1240 (O_1240,N_14922,N_14599);
nand UO_1241 (O_1241,N_14684,N_14692);
and UO_1242 (O_1242,N_14663,N_14629);
and UO_1243 (O_1243,N_14679,N_14958);
nand UO_1244 (O_1244,N_14653,N_14911);
nand UO_1245 (O_1245,N_14729,N_14789);
nor UO_1246 (O_1246,N_14682,N_14689);
nor UO_1247 (O_1247,N_14664,N_14862);
nor UO_1248 (O_1248,N_14613,N_14987);
nor UO_1249 (O_1249,N_14957,N_14614);
nand UO_1250 (O_1250,N_14772,N_14869);
xnor UO_1251 (O_1251,N_14677,N_14850);
nand UO_1252 (O_1252,N_14897,N_14951);
nand UO_1253 (O_1253,N_14562,N_14714);
and UO_1254 (O_1254,N_14924,N_14916);
or UO_1255 (O_1255,N_14835,N_14833);
or UO_1256 (O_1256,N_14574,N_14536);
or UO_1257 (O_1257,N_14671,N_14553);
nor UO_1258 (O_1258,N_14557,N_14969);
nor UO_1259 (O_1259,N_14636,N_14723);
nand UO_1260 (O_1260,N_14841,N_14569);
or UO_1261 (O_1261,N_14750,N_14779);
nor UO_1262 (O_1262,N_14994,N_14937);
nor UO_1263 (O_1263,N_14612,N_14526);
nand UO_1264 (O_1264,N_14561,N_14902);
xnor UO_1265 (O_1265,N_14876,N_14940);
xnor UO_1266 (O_1266,N_14766,N_14850);
nor UO_1267 (O_1267,N_14658,N_14634);
nor UO_1268 (O_1268,N_14659,N_14775);
and UO_1269 (O_1269,N_14666,N_14993);
nor UO_1270 (O_1270,N_14699,N_14868);
and UO_1271 (O_1271,N_14781,N_14597);
or UO_1272 (O_1272,N_14899,N_14668);
nor UO_1273 (O_1273,N_14584,N_14848);
nand UO_1274 (O_1274,N_14670,N_14962);
nand UO_1275 (O_1275,N_14595,N_14517);
and UO_1276 (O_1276,N_14872,N_14585);
or UO_1277 (O_1277,N_14527,N_14599);
and UO_1278 (O_1278,N_14912,N_14646);
or UO_1279 (O_1279,N_14755,N_14765);
xnor UO_1280 (O_1280,N_14616,N_14851);
and UO_1281 (O_1281,N_14571,N_14860);
or UO_1282 (O_1282,N_14948,N_14835);
or UO_1283 (O_1283,N_14829,N_14895);
nor UO_1284 (O_1284,N_14747,N_14962);
or UO_1285 (O_1285,N_14776,N_14789);
or UO_1286 (O_1286,N_14644,N_14845);
and UO_1287 (O_1287,N_14621,N_14815);
and UO_1288 (O_1288,N_14516,N_14523);
xnor UO_1289 (O_1289,N_14632,N_14718);
xnor UO_1290 (O_1290,N_14709,N_14983);
nand UO_1291 (O_1291,N_14906,N_14809);
nor UO_1292 (O_1292,N_14501,N_14703);
or UO_1293 (O_1293,N_14501,N_14610);
nand UO_1294 (O_1294,N_14837,N_14782);
nand UO_1295 (O_1295,N_14790,N_14816);
xor UO_1296 (O_1296,N_14950,N_14944);
nand UO_1297 (O_1297,N_14751,N_14752);
nor UO_1298 (O_1298,N_14804,N_14818);
and UO_1299 (O_1299,N_14658,N_14821);
nor UO_1300 (O_1300,N_14942,N_14890);
and UO_1301 (O_1301,N_14948,N_14953);
and UO_1302 (O_1302,N_14883,N_14758);
and UO_1303 (O_1303,N_14965,N_14814);
nor UO_1304 (O_1304,N_14690,N_14623);
xor UO_1305 (O_1305,N_14852,N_14566);
or UO_1306 (O_1306,N_14506,N_14639);
nor UO_1307 (O_1307,N_14749,N_14967);
nor UO_1308 (O_1308,N_14892,N_14943);
xor UO_1309 (O_1309,N_14688,N_14622);
nand UO_1310 (O_1310,N_14727,N_14576);
and UO_1311 (O_1311,N_14844,N_14709);
xnor UO_1312 (O_1312,N_14615,N_14560);
or UO_1313 (O_1313,N_14892,N_14911);
nand UO_1314 (O_1314,N_14508,N_14502);
nand UO_1315 (O_1315,N_14985,N_14862);
and UO_1316 (O_1316,N_14907,N_14749);
or UO_1317 (O_1317,N_14922,N_14934);
nor UO_1318 (O_1318,N_14945,N_14535);
nor UO_1319 (O_1319,N_14862,N_14841);
nor UO_1320 (O_1320,N_14544,N_14525);
and UO_1321 (O_1321,N_14820,N_14708);
xor UO_1322 (O_1322,N_14752,N_14576);
nor UO_1323 (O_1323,N_14951,N_14644);
or UO_1324 (O_1324,N_14545,N_14602);
or UO_1325 (O_1325,N_14870,N_14648);
nand UO_1326 (O_1326,N_14513,N_14610);
nand UO_1327 (O_1327,N_14796,N_14972);
xnor UO_1328 (O_1328,N_14585,N_14773);
or UO_1329 (O_1329,N_14776,N_14843);
or UO_1330 (O_1330,N_14710,N_14994);
or UO_1331 (O_1331,N_14675,N_14547);
nand UO_1332 (O_1332,N_14550,N_14759);
and UO_1333 (O_1333,N_14753,N_14728);
nand UO_1334 (O_1334,N_14518,N_14655);
nor UO_1335 (O_1335,N_14872,N_14927);
xnor UO_1336 (O_1336,N_14634,N_14752);
nand UO_1337 (O_1337,N_14574,N_14766);
or UO_1338 (O_1338,N_14722,N_14965);
nand UO_1339 (O_1339,N_14911,N_14584);
and UO_1340 (O_1340,N_14557,N_14886);
or UO_1341 (O_1341,N_14968,N_14598);
nor UO_1342 (O_1342,N_14937,N_14892);
nor UO_1343 (O_1343,N_14675,N_14729);
or UO_1344 (O_1344,N_14781,N_14589);
and UO_1345 (O_1345,N_14689,N_14874);
and UO_1346 (O_1346,N_14544,N_14901);
nand UO_1347 (O_1347,N_14929,N_14933);
and UO_1348 (O_1348,N_14935,N_14878);
xnor UO_1349 (O_1349,N_14599,N_14880);
and UO_1350 (O_1350,N_14680,N_14713);
xnor UO_1351 (O_1351,N_14946,N_14666);
xor UO_1352 (O_1352,N_14653,N_14755);
and UO_1353 (O_1353,N_14595,N_14593);
or UO_1354 (O_1354,N_14541,N_14740);
and UO_1355 (O_1355,N_14976,N_14849);
or UO_1356 (O_1356,N_14758,N_14564);
and UO_1357 (O_1357,N_14908,N_14651);
nor UO_1358 (O_1358,N_14521,N_14729);
xnor UO_1359 (O_1359,N_14533,N_14531);
or UO_1360 (O_1360,N_14994,N_14541);
xor UO_1361 (O_1361,N_14903,N_14567);
nor UO_1362 (O_1362,N_14691,N_14537);
and UO_1363 (O_1363,N_14538,N_14547);
xnor UO_1364 (O_1364,N_14942,N_14823);
and UO_1365 (O_1365,N_14606,N_14560);
or UO_1366 (O_1366,N_14828,N_14518);
nand UO_1367 (O_1367,N_14904,N_14648);
and UO_1368 (O_1368,N_14583,N_14853);
nand UO_1369 (O_1369,N_14733,N_14555);
xnor UO_1370 (O_1370,N_14610,N_14534);
nand UO_1371 (O_1371,N_14606,N_14865);
nand UO_1372 (O_1372,N_14626,N_14903);
or UO_1373 (O_1373,N_14625,N_14558);
and UO_1374 (O_1374,N_14796,N_14623);
nand UO_1375 (O_1375,N_14727,N_14834);
nand UO_1376 (O_1376,N_14557,N_14691);
and UO_1377 (O_1377,N_14925,N_14972);
xor UO_1378 (O_1378,N_14935,N_14964);
nor UO_1379 (O_1379,N_14929,N_14587);
nand UO_1380 (O_1380,N_14849,N_14512);
nand UO_1381 (O_1381,N_14991,N_14783);
or UO_1382 (O_1382,N_14968,N_14656);
nand UO_1383 (O_1383,N_14739,N_14523);
xor UO_1384 (O_1384,N_14799,N_14930);
nand UO_1385 (O_1385,N_14893,N_14836);
nand UO_1386 (O_1386,N_14553,N_14751);
xor UO_1387 (O_1387,N_14698,N_14802);
xnor UO_1388 (O_1388,N_14937,N_14725);
nand UO_1389 (O_1389,N_14964,N_14631);
or UO_1390 (O_1390,N_14807,N_14941);
and UO_1391 (O_1391,N_14902,N_14866);
xor UO_1392 (O_1392,N_14626,N_14758);
nor UO_1393 (O_1393,N_14914,N_14888);
nand UO_1394 (O_1394,N_14546,N_14713);
nor UO_1395 (O_1395,N_14955,N_14992);
nor UO_1396 (O_1396,N_14746,N_14585);
nand UO_1397 (O_1397,N_14915,N_14651);
xnor UO_1398 (O_1398,N_14899,N_14867);
nor UO_1399 (O_1399,N_14888,N_14591);
or UO_1400 (O_1400,N_14897,N_14906);
xor UO_1401 (O_1401,N_14515,N_14722);
xnor UO_1402 (O_1402,N_14565,N_14643);
xor UO_1403 (O_1403,N_14620,N_14780);
or UO_1404 (O_1404,N_14685,N_14858);
nand UO_1405 (O_1405,N_14778,N_14722);
and UO_1406 (O_1406,N_14669,N_14835);
nor UO_1407 (O_1407,N_14939,N_14696);
and UO_1408 (O_1408,N_14587,N_14863);
or UO_1409 (O_1409,N_14587,N_14858);
or UO_1410 (O_1410,N_14960,N_14711);
or UO_1411 (O_1411,N_14656,N_14712);
nand UO_1412 (O_1412,N_14715,N_14924);
nand UO_1413 (O_1413,N_14831,N_14513);
xor UO_1414 (O_1414,N_14623,N_14758);
or UO_1415 (O_1415,N_14684,N_14602);
and UO_1416 (O_1416,N_14628,N_14693);
and UO_1417 (O_1417,N_14762,N_14896);
nand UO_1418 (O_1418,N_14828,N_14797);
xor UO_1419 (O_1419,N_14766,N_14891);
nor UO_1420 (O_1420,N_14744,N_14971);
nor UO_1421 (O_1421,N_14979,N_14846);
nor UO_1422 (O_1422,N_14901,N_14809);
nor UO_1423 (O_1423,N_14785,N_14690);
xnor UO_1424 (O_1424,N_14706,N_14593);
nor UO_1425 (O_1425,N_14613,N_14753);
or UO_1426 (O_1426,N_14955,N_14939);
nand UO_1427 (O_1427,N_14892,N_14590);
or UO_1428 (O_1428,N_14843,N_14513);
nor UO_1429 (O_1429,N_14715,N_14820);
nand UO_1430 (O_1430,N_14891,N_14832);
and UO_1431 (O_1431,N_14746,N_14587);
nand UO_1432 (O_1432,N_14733,N_14761);
xnor UO_1433 (O_1433,N_14663,N_14708);
nand UO_1434 (O_1434,N_14539,N_14700);
and UO_1435 (O_1435,N_14843,N_14771);
or UO_1436 (O_1436,N_14893,N_14677);
and UO_1437 (O_1437,N_14939,N_14902);
and UO_1438 (O_1438,N_14678,N_14674);
or UO_1439 (O_1439,N_14952,N_14559);
xnor UO_1440 (O_1440,N_14534,N_14531);
nor UO_1441 (O_1441,N_14725,N_14974);
xor UO_1442 (O_1442,N_14746,N_14935);
xor UO_1443 (O_1443,N_14743,N_14684);
and UO_1444 (O_1444,N_14974,N_14723);
or UO_1445 (O_1445,N_14751,N_14914);
xnor UO_1446 (O_1446,N_14677,N_14605);
or UO_1447 (O_1447,N_14577,N_14798);
xnor UO_1448 (O_1448,N_14991,N_14913);
and UO_1449 (O_1449,N_14695,N_14516);
or UO_1450 (O_1450,N_14732,N_14708);
xnor UO_1451 (O_1451,N_14842,N_14937);
or UO_1452 (O_1452,N_14808,N_14835);
and UO_1453 (O_1453,N_14780,N_14765);
and UO_1454 (O_1454,N_14795,N_14800);
and UO_1455 (O_1455,N_14767,N_14816);
nor UO_1456 (O_1456,N_14718,N_14901);
xor UO_1457 (O_1457,N_14618,N_14505);
xnor UO_1458 (O_1458,N_14971,N_14881);
and UO_1459 (O_1459,N_14894,N_14619);
or UO_1460 (O_1460,N_14689,N_14951);
and UO_1461 (O_1461,N_14988,N_14953);
or UO_1462 (O_1462,N_14710,N_14986);
or UO_1463 (O_1463,N_14900,N_14685);
or UO_1464 (O_1464,N_14516,N_14883);
xor UO_1465 (O_1465,N_14829,N_14599);
and UO_1466 (O_1466,N_14537,N_14788);
nand UO_1467 (O_1467,N_14878,N_14507);
and UO_1468 (O_1468,N_14683,N_14575);
nor UO_1469 (O_1469,N_14825,N_14796);
or UO_1470 (O_1470,N_14652,N_14502);
and UO_1471 (O_1471,N_14600,N_14796);
or UO_1472 (O_1472,N_14854,N_14652);
or UO_1473 (O_1473,N_14812,N_14968);
or UO_1474 (O_1474,N_14906,N_14960);
nor UO_1475 (O_1475,N_14509,N_14828);
or UO_1476 (O_1476,N_14584,N_14649);
nor UO_1477 (O_1477,N_14816,N_14775);
nor UO_1478 (O_1478,N_14635,N_14961);
nor UO_1479 (O_1479,N_14988,N_14539);
or UO_1480 (O_1480,N_14859,N_14628);
or UO_1481 (O_1481,N_14605,N_14521);
and UO_1482 (O_1482,N_14934,N_14745);
nor UO_1483 (O_1483,N_14828,N_14977);
nor UO_1484 (O_1484,N_14728,N_14505);
nor UO_1485 (O_1485,N_14908,N_14732);
nor UO_1486 (O_1486,N_14693,N_14815);
xor UO_1487 (O_1487,N_14871,N_14965);
nand UO_1488 (O_1488,N_14576,N_14605);
xor UO_1489 (O_1489,N_14864,N_14543);
xnor UO_1490 (O_1490,N_14884,N_14738);
nor UO_1491 (O_1491,N_14633,N_14540);
or UO_1492 (O_1492,N_14609,N_14582);
nand UO_1493 (O_1493,N_14560,N_14869);
xnor UO_1494 (O_1494,N_14741,N_14863);
nor UO_1495 (O_1495,N_14839,N_14911);
nand UO_1496 (O_1496,N_14818,N_14879);
nor UO_1497 (O_1497,N_14578,N_14674);
nand UO_1498 (O_1498,N_14779,N_14534);
nand UO_1499 (O_1499,N_14839,N_14624);
xnor UO_1500 (O_1500,N_14970,N_14882);
xnor UO_1501 (O_1501,N_14886,N_14579);
or UO_1502 (O_1502,N_14834,N_14742);
nand UO_1503 (O_1503,N_14630,N_14748);
and UO_1504 (O_1504,N_14718,N_14794);
nor UO_1505 (O_1505,N_14984,N_14682);
and UO_1506 (O_1506,N_14907,N_14919);
xor UO_1507 (O_1507,N_14911,N_14997);
nand UO_1508 (O_1508,N_14672,N_14947);
and UO_1509 (O_1509,N_14847,N_14786);
xnor UO_1510 (O_1510,N_14647,N_14823);
nor UO_1511 (O_1511,N_14963,N_14742);
or UO_1512 (O_1512,N_14814,N_14779);
or UO_1513 (O_1513,N_14577,N_14793);
or UO_1514 (O_1514,N_14633,N_14732);
and UO_1515 (O_1515,N_14519,N_14506);
xnor UO_1516 (O_1516,N_14612,N_14531);
and UO_1517 (O_1517,N_14558,N_14690);
or UO_1518 (O_1518,N_14753,N_14973);
or UO_1519 (O_1519,N_14519,N_14600);
xor UO_1520 (O_1520,N_14854,N_14518);
and UO_1521 (O_1521,N_14860,N_14599);
nand UO_1522 (O_1522,N_14880,N_14830);
xnor UO_1523 (O_1523,N_14982,N_14644);
nand UO_1524 (O_1524,N_14665,N_14927);
or UO_1525 (O_1525,N_14700,N_14887);
nand UO_1526 (O_1526,N_14641,N_14823);
nand UO_1527 (O_1527,N_14704,N_14689);
or UO_1528 (O_1528,N_14671,N_14839);
or UO_1529 (O_1529,N_14961,N_14999);
nor UO_1530 (O_1530,N_14613,N_14821);
and UO_1531 (O_1531,N_14790,N_14860);
nand UO_1532 (O_1532,N_14808,N_14926);
nor UO_1533 (O_1533,N_14888,N_14796);
nor UO_1534 (O_1534,N_14525,N_14697);
nor UO_1535 (O_1535,N_14899,N_14526);
or UO_1536 (O_1536,N_14890,N_14548);
nor UO_1537 (O_1537,N_14845,N_14807);
and UO_1538 (O_1538,N_14833,N_14921);
and UO_1539 (O_1539,N_14564,N_14784);
nor UO_1540 (O_1540,N_14589,N_14750);
nor UO_1541 (O_1541,N_14933,N_14543);
xnor UO_1542 (O_1542,N_14732,N_14914);
and UO_1543 (O_1543,N_14843,N_14943);
and UO_1544 (O_1544,N_14998,N_14641);
nand UO_1545 (O_1545,N_14639,N_14764);
and UO_1546 (O_1546,N_14617,N_14841);
xnor UO_1547 (O_1547,N_14951,N_14931);
xor UO_1548 (O_1548,N_14821,N_14688);
or UO_1549 (O_1549,N_14823,N_14653);
xnor UO_1550 (O_1550,N_14539,N_14521);
or UO_1551 (O_1551,N_14556,N_14550);
xnor UO_1552 (O_1552,N_14961,N_14884);
xor UO_1553 (O_1553,N_14889,N_14829);
xor UO_1554 (O_1554,N_14890,N_14881);
or UO_1555 (O_1555,N_14602,N_14994);
xor UO_1556 (O_1556,N_14894,N_14618);
or UO_1557 (O_1557,N_14534,N_14862);
xor UO_1558 (O_1558,N_14812,N_14890);
xnor UO_1559 (O_1559,N_14823,N_14500);
and UO_1560 (O_1560,N_14695,N_14829);
xor UO_1561 (O_1561,N_14788,N_14559);
nor UO_1562 (O_1562,N_14905,N_14635);
xor UO_1563 (O_1563,N_14916,N_14613);
or UO_1564 (O_1564,N_14563,N_14860);
nor UO_1565 (O_1565,N_14965,N_14695);
nor UO_1566 (O_1566,N_14913,N_14599);
nor UO_1567 (O_1567,N_14581,N_14542);
xnor UO_1568 (O_1568,N_14590,N_14516);
nand UO_1569 (O_1569,N_14917,N_14794);
nand UO_1570 (O_1570,N_14696,N_14543);
nand UO_1571 (O_1571,N_14845,N_14893);
nor UO_1572 (O_1572,N_14900,N_14888);
or UO_1573 (O_1573,N_14544,N_14658);
nand UO_1574 (O_1574,N_14717,N_14955);
nand UO_1575 (O_1575,N_14835,N_14507);
nor UO_1576 (O_1576,N_14796,N_14854);
xor UO_1577 (O_1577,N_14898,N_14799);
and UO_1578 (O_1578,N_14514,N_14734);
nor UO_1579 (O_1579,N_14922,N_14781);
xnor UO_1580 (O_1580,N_14606,N_14911);
and UO_1581 (O_1581,N_14863,N_14614);
nand UO_1582 (O_1582,N_14900,N_14809);
or UO_1583 (O_1583,N_14869,N_14983);
and UO_1584 (O_1584,N_14900,N_14855);
xor UO_1585 (O_1585,N_14619,N_14985);
nor UO_1586 (O_1586,N_14696,N_14583);
xnor UO_1587 (O_1587,N_14787,N_14692);
xnor UO_1588 (O_1588,N_14681,N_14692);
or UO_1589 (O_1589,N_14953,N_14780);
or UO_1590 (O_1590,N_14808,N_14809);
xnor UO_1591 (O_1591,N_14754,N_14598);
xnor UO_1592 (O_1592,N_14633,N_14858);
or UO_1593 (O_1593,N_14512,N_14698);
and UO_1594 (O_1594,N_14681,N_14854);
nand UO_1595 (O_1595,N_14684,N_14669);
and UO_1596 (O_1596,N_14986,N_14996);
or UO_1597 (O_1597,N_14956,N_14985);
xnor UO_1598 (O_1598,N_14995,N_14709);
nand UO_1599 (O_1599,N_14703,N_14915);
nor UO_1600 (O_1600,N_14957,N_14564);
and UO_1601 (O_1601,N_14953,N_14975);
and UO_1602 (O_1602,N_14981,N_14607);
and UO_1603 (O_1603,N_14824,N_14955);
xnor UO_1604 (O_1604,N_14883,N_14915);
xnor UO_1605 (O_1605,N_14830,N_14973);
or UO_1606 (O_1606,N_14892,N_14673);
and UO_1607 (O_1607,N_14945,N_14955);
nor UO_1608 (O_1608,N_14776,N_14640);
and UO_1609 (O_1609,N_14831,N_14658);
xnor UO_1610 (O_1610,N_14511,N_14856);
or UO_1611 (O_1611,N_14844,N_14915);
xnor UO_1612 (O_1612,N_14700,N_14640);
or UO_1613 (O_1613,N_14962,N_14887);
xor UO_1614 (O_1614,N_14863,N_14886);
nor UO_1615 (O_1615,N_14635,N_14541);
nor UO_1616 (O_1616,N_14560,N_14677);
nand UO_1617 (O_1617,N_14858,N_14705);
nor UO_1618 (O_1618,N_14835,N_14856);
nor UO_1619 (O_1619,N_14811,N_14917);
nor UO_1620 (O_1620,N_14735,N_14669);
or UO_1621 (O_1621,N_14839,N_14840);
nor UO_1622 (O_1622,N_14541,N_14505);
and UO_1623 (O_1623,N_14518,N_14755);
or UO_1624 (O_1624,N_14769,N_14888);
and UO_1625 (O_1625,N_14943,N_14847);
xor UO_1626 (O_1626,N_14700,N_14882);
nor UO_1627 (O_1627,N_14567,N_14570);
or UO_1628 (O_1628,N_14522,N_14615);
xnor UO_1629 (O_1629,N_14935,N_14868);
nor UO_1630 (O_1630,N_14505,N_14669);
nand UO_1631 (O_1631,N_14868,N_14747);
nor UO_1632 (O_1632,N_14832,N_14716);
nand UO_1633 (O_1633,N_14883,N_14523);
nor UO_1634 (O_1634,N_14704,N_14813);
and UO_1635 (O_1635,N_14950,N_14948);
nand UO_1636 (O_1636,N_14900,N_14776);
nand UO_1637 (O_1637,N_14733,N_14707);
nand UO_1638 (O_1638,N_14674,N_14682);
xor UO_1639 (O_1639,N_14562,N_14905);
nand UO_1640 (O_1640,N_14978,N_14664);
or UO_1641 (O_1641,N_14786,N_14984);
and UO_1642 (O_1642,N_14641,N_14981);
and UO_1643 (O_1643,N_14508,N_14820);
nand UO_1644 (O_1644,N_14967,N_14668);
or UO_1645 (O_1645,N_14823,N_14915);
or UO_1646 (O_1646,N_14512,N_14662);
nor UO_1647 (O_1647,N_14783,N_14764);
or UO_1648 (O_1648,N_14506,N_14720);
xor UO_1649 (O_1649,N_14898,N_14741);
and UO_1650 (O_1650,N_14549,N_14762);
nor UO_1651 (O_1651,N_14651,N_14575);
xnor UO_1652 (O_1652,N_14576,N_14823);
and UO_1653 (O_1653,N_14990,N_14764);
nor UO_1654 (O_1654,N_14586,N_14988);
nand UO_1655 (O_1655,N_14967,N_14565);
nor UO_1656 (O_1656,N_14686,N_14947);
and UO_1657 (O_1657,N_14677,N_14883);
nand UO_1658 (O_1658,N_14912,N_14673);
nand UO_1659 (O_1659,N_14984,N_14554);
or UO_1660 (O_1660,N_14635,N_14857);
nand UO_1661 (O_1661,N_14991,N_14584);
xnor UO_1662 (O_1662,N_14772,N_14936);
nand UO_1663 (O_1663,N_14545,N_14834);
nand UO_1664 (O_1664,N_14798,N_14732);
or UO_1665 (O_1665,N_14555,N_14696);
and UO_1666 (O_1666,N_14857,N_14893);
nor UO_1667 (O_1667,N_14936,N_14548);
and UO_1668 (O_1668,N_14835,N_14892);
or UO_1669 (O_1669,N_14992,N_14706);
xnor UO_1670 (O_1670,N_14726,N_14699);
nand UO_1671 (O_1671,N_14987,N_14697);
nor UO_1672 (O_1672,N_14660,N_14743);
nor UO_1673 (O_1673,N_14590,N_14648);
xnor UO_1674 (O_1674,N_14979,N_14541);
nor UO_1675 (O_1675,N_14742,N_14842);
nand UO_1676 (O_1676,N_14962,N_14892);
xor UO_1677 (O_1677,N_14626,N_14554);
nand UO_1678 (O_1678,N_14995,N_14642);
or UO_1679 (O_1679,N_14911,N_14616);
xnor UO_1680 (O_1680,N_14911,N_14764);
nand UO_1681 (O_1681,N_14639,N_14737);
nand UO_1682 (O_1682,N_14917,N_14887);
and UO_1683 (O_1683,N_14858,N_14764);
xnor UO_1684 (O_1684,N_14837,N_14511);
nand UO_1685 (O_1685,N_14504,N_14855);
nand UO_1686 (O_1686,N_14793,N_14933);
xnor UO_1687 (O_1687,N_14882,N_14918);
and UO_1688 (O_1688,N_14726,N_14819);
nor UO_1689 (O_1689,N_14531,N_14607);
nor UO_1690 (O_1690,N_14603,N_14648);
xor UO_1691 (O_1691,N_14965,N_14732);
and UO_1692 (O_1692,N_14620,N_14781);
xor UO_1693 (O_1693,N_14832,N_14713);
xnor UO_1694 (O_1694,N_14995,N_14835);
or UO_1695 (O_1695,N_14951,N_14706);
xnor UO_1696 (O_1696,N_14590,N_14809);
or UO_1697 (O_1697,N_14728,N_14645);
xor UO_1698 (O_1698,N_14562,N_14718);
or UO_1699 (O_1699,N_14688,N_14698);
nor UO_1700 (O_1700,N_14868,N_14567);
and UO_1701 (O_1701,N_14759,N_14897);
and UO_1702 (O_1702,N_14680,N_14789);
xor UO_1703 (O_1703,N_14860,N_14828);
xor UO_1704 (O_1704,N_14987,N_14675);
or UO_1705 (O_1705,N_14780,N_14581);
or UO_1706 (O_1706,N_14667,N_14931);
nor UO_1707 (O_1707,N_14750,N_14868);
nor UO_1708 (O_1708,N_14752,N_14896);
nand UO_1709 (O_1709,N_14879,N_14605);
or UO_1710 (O_1710,N_14892,N_14856);
or UO_1711 (O_1711,N_14753,N_14542);
xor UO_1712 (O_1712,N_14761,N_14996);
and UO_1713 (O_1713,N_14779,N_14937);
xor UO_1714 (O_1714,N_14698,N_14552);
nor UO_1715 (O_1715,N_14806,N_14575);
nand UO_1716 (O_1716,N_14882,N_14583);
and UO_1717 (O_1717,N_14967,N_14868);
nor UO_1718 (O_1718,N_14857,N_14830);
nor UO_1719 (O_1719,N_14754,N_14749);
or UO_1720 (O_1720,N_14635,N_14657);
nor UO_1721 (O_1721,N_14966,N_14530);
xnor UO_1722 (O_1722,N_14864,N_14961);
nand UO_1723 (O_1723,N_14643,N_14991);
nand UO_1724 (O_1724,N_14997,N_14894);
nor UO_1725 (O_1725,N_14644,N_14811);
nor UO_1726 (O_1726,N_14936,N_14551);
or UO_1727 (O_1727,N_14839,N_14873);
and UO_1728 (O_1728,N_14506,N_14833);
xor UO_1729 (O_1729,N_14729,N_14643);
xor UO_1730 (O_1730,N_14995,N_14939);
or UO_1731 (O_1731,N_14753,N_14641);
xnor UO_1732 (O_1732,N_14604,N_14894);
or UO_1733 (O_1733,N_14949,N_14630);
and UO_1734 (O_1734,N_14585,N_14770);
or UO_1735 (O_1735,N_14587,N_14932);
or UO_1736 (O_1736,N_14878,N_14672);
xnor UO_1737 (O_1737,N_14623,N_14786);
nand UO_1738 (O_1738,N_14969,N_14902);
nor UO_1739 (O_1739,N_14559,N_14686);
or UO_1740 (O_1740,N_14971,N_14688);
nor UO_1741 (O_1741,N_14647,N_14872);
or UO_1742 (O_1742,N_14801,N_14945);
and UO_1743 (O_1743,N_14904,N_14712);
nor UO_1744 (O_1744,N_14900,N_14954);
nor UO_1745 (O_1745,N_14937,N_14764);
xnor UO_1746 (O_1746,N_14686,N_14896);
or UO_1747 (O_1747,N_14603,N_14755);
xnor UO_1748 (O_1748,N_14588,N_14762);
nor UO_1749 (O_1749,N_14622,N_14944);
or UO_1750 (O_1750,N_14684,N_14773);
and UO_1751 (O_1751,N_14898,N_14633);
nand UO_1752 (O_1752,N_14739,N_14908);
and UO_1753 (O_1753,N_14983,N_14730);
and UO_1754 (O_1754,N_14813,N_14756);
nand UO_1755 (O_1755,N_14840,N_14678);
or UO_1756 (O_1756,N_14599,N_14992);
nand UO_1757 (O_1757,N_14826,N_14794);
or UO_1758 (O_1758,N_14719,N_14934);
nand UO_1759 (O_1759,N_14506,N_14875);
and UO_1760 (O_1760,N_14501,N_14749);
nor UO_1761 (O_1761,N_14616,N_14633);
or UO_1762 (O_1762,N_14711,N_14549);
and UO_1763 (O_1763,N_14877,N_14592);
nand UO_1764 (O_1764,N_14783,N_14848);
nor UO_1765 (O_1765,N_14622,N_14737);
nor UO_1766 (O_1766,N_14957,N_14974);
or UO_1767 (O_1767,N_14588,N_14798);
nand UO_1768 (O_1768,N_14894,N_14773);
or UO_1769 (O_1769,N_14726,N_14997);
nand UO_1770 (O_1770,N_14983,N_14796);
xnor UO_1771 (O_1771,N_14889,N_14516);
nand UO_1772 (O_1772,N_14579,N_14602);
nor UO_1773 (O_1773,N_14844,N_14679);
nor UO_1774 (O_1774,N_14608,N_14873);
nand UO_1775 (O_1775,N_14768,N_14977);
nand UO_1776 (O_1776,N_14784,N_14923);
or UO_1777 (O_1777,N_14566,N_14797);
nand UO_1778 (O_1778,N_14746,N_14959);
xnor UO_1779 (O_1779,N_14578,N_14601);
nand UO_1780 (O_1780,N_14884,N_14767);
and UO_1781 (O_1781,N_14878,N_14850);
xnor UO_1782 (O_1782,N_14819,N_14752);
and UO_1783 (O_1783,N_14624,N_14675);
nand UO_1784 (O_1784,N_14846,N_14981);
and UO_1785 (O_1785,N_14701,N_14630);
xor UO_1786 (O_1786,N_14921,N_14505);
nand UO_1787 (O_1787,N_14587,N_14546);
and UO_1788 (O_1788,N_14704,N_14712);
or UO_1789 (O_1789,N_14684,N_14573);
or UO_1790 (O_1790,N_14830,N_14535);
nor UO_1791 (O_1791,N_14843,N_14669);
and UO_1792 (O_1792,N_14711,N_14618);
nand UO_1793 (O_1793,N_14804,N_14775);
nand UO_1794 (O_1794,N_14573,N_14699);
nand UO_1795 (O_1795,N_14794,N_14588);
and UO_1796 (O_1796,N_14635,N_14549);
xor UO_1797 (O_1797,N_14755,N_14939);
nand UO_1798 (O_1798,N_14678,N_14783);
nand UO_1799 (O_1799,N_14912,N_14505);
nand UO_1800 (O_1800,N_14774,N_14893);
and UO_1801 (O_1801,N_14918,N_14815);
and UO_1802 (O_1802,N_14884,N_14970);
nand UO_1803 (O_1803,N_14646,N_14987);
and UO_1804 (O_1804,N_14911,N_14978);
or UO_1805 (O_1805,N_14532,N_14898);
nand UO_1806 (O_1806,N_14662,N_14542);
xnor UO_1807 (O_1807,N_14679,N_14890);
or UO_1808 (O_1808,N_14541,N_14935);
and UO_1809 (O_1809,N_14737,N_14884);
or UO_1810 (O_1810,N_14644,N_14756);
xnor UO_1811 (O_1811,N_14744,N_14980);
xor UO_1812 (O_1812,N_14711,N_14770);
nand UO_1813 (O_1813,N_14955,N_14957);
nand UO_1814 (O_1814,N_14608,N_14742);
xor UO_1815 (O_1815,N_14589,N_14665);
nand UO_1816 (O_1816,N_14947,N_14797);
xor UO_1817 (O_1817,N_14728,N_14947);
xnor UO_1818 (O_1818,N_14524,N_14895);
nand UO_1819 (O_1819,N_14902,N_14941);
xnor UO_1820 (O_1820,N_14808,N_14918);
nand UO_1821 (O_1821,N_14540,N_14775);
nand UO_1822 (O_1822,N_14830,N_14682);
nor UO_1823 (O_1823,N_14923,N_14952);
xor UO_1824 (O_1824,N_14909,N_14586);
and UO_1825 (O_1825,N_14578,N_14629);
nand UO_1826 (O_1826,N_14972,N_14621);
nor UO_1827 (O_1827,N_14786,N_14517);
or UO_1828 (O_1828,N_14850,N_14661);
nand UO_1829 (O_1829,N_14596,N_14698);
nor UO_1830 (O_1830,N_14951,N_14622);
nand UO_1831 (O_1831,N_14881,N_14505);
xnor UO_1832 (O_1832,N_14582,N_14721);
nor UO_1833 (O_1833,N_14548,N_14521);
or UO_1834 (O_1834,N_14662,N_14873);
nand UO_1835 (O_1835,N_14961,N_14752);
nor UO_1836 (O_1836,N_14855,N_14860);
xor UO_1837 (O_1837,N_14796,N_14709);
and UO_1838 (O_1838,N_14941,N_14812);
nand UO_1839 (O_1839,N_14940,N_14942);
nor UO_1840 (O_1840,N_14938,N_14955);
xnor UO_1841 (O_1841,N_14843,N_14632);
or UO_1842 (O_1842,N_14906,N_14533);
and UO_1843 (O_1843,N_14763,N_14575);
nor UO_1844 (O_1844,N_14991,N_14769);
or UO_1845 (O_1845,N_14829,N_14827);
xor UO_1846 (O_1846,N_14861,N_14584);
and UO_1847 (O_1847,N_14521,N_14620);
or UO_1848 (O_1848,N_14914,N_14794);
xnor UO_1849 (O_1849,N_14697,N_14985);
nor UO_1850 (O_1850,N_14711,N_14854);
xor UO_1851 (O_1851,N_14582,N_14825);
xnor UO_1852 (O_1852,N_14663,N_14722);
xor UO_1853 (O_1853,N_14980,N_14813);
xor UO_1854 (O_1854,N_14761,N_14976);
nand UO_1855 (O_1855,N_14989,N_14748);
or UO_1856 (O_1856,N_14702,N_14566);
and UO_1857 (O_1857,N_14502,N_14672);
nor UO_1858 (O_1858,N_14992,N_14867);
and UO_1859 (O_1859,N_14721,N_14969);
or UO_1860 (O_1860,N_14700,N_14972);
and UO_1861 (O_1861,N_14700,N_14791);
nor UO_1862 (O_1862,N_14910,N_14830);
or UO_1863 (O_1863,N_14922,N_14850);
xnor UO_1864 (O_1864,N_14834,N_14882);
nor UO_1865 (O_1865,N_14983,N_14687);
and UO_1866 (O_1866,N_14523,N_14598);
or UO_1867 (O_1867,N_14902,N_14539);
xnor UO_1868 (O_1868,N_14600,N_14576);
and UO_1869 (O_1869,N_14861,N_14734);
nor UO_1870 (O_1870,N_14597,N_14514);
and UO_1871 (O_1871,N_14984,N_14885);
and UO_1872 (O_1872,N_14850,N_14906);
nand UO_1873 (O_1873,N_14622,N_14523);
nor UO_1874 (O_1874,N_14693,N_14764);
and UO_1875 (O_1875,N_14762,N_14524);
and UO_1876 (O_1876,N_14758,N_14841);
nor UO_1877 (O_1877,N_14944,N_14948);
xnor UO_1878 (O_1878,N_14857,N_14707);
nor UO_1879 (O_1879,N_14898,N_14993);
xor UO_1880 (O_1880,N_14828,N_14685);
and UO_1881 (O_1881,N_14935,N_14720);
and UO_1882 (O_1882,N_14841,N_14669);
or UO_1883 (O_1883,N_14504,N_14540);
nor UO_1884 (O_1884,N_14669,N_14978);
xor UO_1885 (O_1885,N_14508,N_14839);
nand UO_1886 (O_1886,N_14880,N_14909);
nand UO_1887 (O_1887,N_14930,N_14629);
nand UO_1888 (O_1888,N_14743,N_14784);
or UO_1889 (O_1889,N_14949,N_14923);
xor UO_1890 (O_1890,N_14710,N_14862);
and UO_1891 (O_1891,N_14921,N_14552);
nor UO_1892 (O_1892,N_14501,N_14698);
nand UO_1893 (O_1893,N_14926,N_14678);
and UO_1894 (O_1894,N_14841,N_14892);
and UO_1895 (O_1895,N_14958,N_14913);
nor UO_1896 (O_1896,N_14855,N_14963);
and UO_1897 (O_1897,N_14586,N_14604);
nand UO_1898 (O_1898,N_14928,N_14781);
or UO_1899 (O_1899,N_14918,N_14720);
and UO_1900 (O_1900,N_14613,N_14857);
and UO_1901 (O_1901,N_14819,N_14922);
nor UO_1902 (O_1902,N_14856,N_14811);
nand UO_1903 (O_1903,N_14853,N_14900);
nor UO_1904 (O_1904,N_14840,N_14680);
xor UO_1905 (O_1905,N_14719,N_14858);
nor UO_1906 (O_1906,N_14929,N_14817);
nand UO_1907 (O_1907,N_14920,N_14883);
and UO_1908 (O_1908,N_14646,N_14508);
nand UO_1909 (O_1909,N_14755,N_14910);
nand UO_1910 (O_1910,N_14925,N_14674);
and UO_1911 (O_1911,N_14536,N_14813);
xor UO_1912 (O_1912,N_14806,N_14931);
nand UO_1913 (O_1913,N_14828,N_14806);
or UO_1914 (O_1914,N_14823,N_14945);
nor UO_1915 (O_1915,N_14720,N_14850);
and UO_1916 (O_1916,N_14643,N_14876);
nor UO_1917 (O_1917,N_14860,N_14621);
xnor UO_1918 (O_1918,N_14837,N_14927);
and UO_1919 (O_1919,N_14691,N_14670);
xnor UO_1920 (O_1920,N_14863,N_14595);
and UO_1921 (O_1921,N_14527,N_14647);
or UO_1922 (O_1922,N_14851,N_14708);
and UO_1923 (O_1923,N_14514,N_14706);
and UO_1924 (O_1924,N_14911,N_14703);
and UO_1925 (O_1925,N_14859,N_14610);
nor UO_1926 (O_1926,N_14775,N_14857);
and UO_1927 (O_1927,N_14902,N_14653);
or UO_1928 (O_1928,N_14806,N_14510);
and UO_1929 (O_1929,N_14515,N_14672);
nand UO_1930 (O_1930,N_14879,N_14710);
and UO_1931 (O_1931,N_14512,N_14912);
and UO_1932 (O_1932,N_14906,N_14502);
nand UO_1933 (O_1933,N_14531,N_14856);
nand UO_1934 (O_1934,N_14860,N_14560);
or UO_1935 (O_1935,N_14576,N_14697);
nor UO_1936 (O_1936,N_14895,N_14541);
xor UO_1937 (O_1937,N_14815,N_14872);
and UO_1938 (O_1938,N_14735,N_14998);
nand UO_1939 (O_1939,N_14580,N_14707);
xnor UO_1940 (O_1940,N_14559,N_14977);
nor UO_1941 (O_1941,N_14724,N_14566);
nor UO_1942 (O_1942,N_14749,N_14756);
nand UO_1943 (O_1943,N_14539,N_14973);
or UO_1944 (O_1944,N_14870,N_14744);
and UO_1945 (O_1945,N_14879,N_14722);
or UO_1946 (O_1946,N_14918,N_14593);
nand UO_1947 (O_1947,N_14989,N_14931);
or UO_1948 (O_1948,N_14768,N_14721);
and UO_1949 (O_1949,N_14890,N_14500);
xor UO_1950 (O_1950,N_14591,N_14978);
xor UO_1951 (O_1951,N_14509,N_14820);
and UO_1952 (O_1952,N_14747,N_14825);
and UO_1953 (O_1953,N_14698,N_14616);
nand UO_1954 (O_1954,N_14809,N_14538);
or UO_1955 (O_1955,N_14901,N_14802);
or UO_1956 (O_1956,N_14528,N_14589);
and UO_1957 (O_1957,N_14637,N_14777);
or UO_1958 (O_1958,N_14666,N_14894);
and UO_1959 (O_1959,N_14519,N_14572);
nor UO_1960 (O_1960,N_14812,N_14896);
nor UO_1961 (O_1961,N_14679,N_14884);
or UO_1962 (O_1962,N_14632,N_14913);
xnor UO_1963 (O_1963,N_14951,N_14905);
nor UO_1964 (O_1964,N_14615,N_14681);
and UO_1965 (O_1965,N_14631,N_14902);
xnor UO_1966 (O_1966,N_14809,N_14695);
nor UO_1967 (O_1967,N_14500,N_14756);
or UO_1968 (O_1968,N_14913,N_14818);
nor UO_1969 (O_1969,N_14666,N_14757);
nand UO_1970 (O_1970,N_14516,N_14945);
xor UO_1971 (O_1971,N_14815,N_14712);
or UO_1972 (O_1972,N_14875,N_14742);
and UO_1973 (O_1973,N_14627,N_14643);
nand UO_1974 (O_1974,N_14559,N_14929);
xor UO_1975 (O_1975,N_14788,N_14918);
xnor UO_1976 (O_1976,N_14780,N_14626);
nor UO_1977 (O_1977,N_14935,N_14778);
xor UO_1978 (O_1978,N_14609,N_14685);
nor UO_1979 (O_1979,N_14805,N_14564);
xor UO_1980 (O_1980,N_14904,N_14901);
xor UO_1981 (O_1981,N_14817,N_14639);
or UO_1982 (O_1982,N_14586,N_14779);
nand UO_1983 (O_1983,N_14839,N_14777);
nor UO_1984 (O_1984,N_14669,N_14885);
or UO_1985 (O_1985,N_14733,N_14803);
or UO_1986 (O_1986,N_14652,N_14947);
nand UO_1987 (O_1987,N_14733,N_14934);
or UO_1988 (O_1988,N_14948,N_14707);
xor UO_1989 (O_1989,N_14724,N_14970);
xnor UO_1990 (O_1990,N_14847,N_14607);
or UO_1991 (O_1991,N_14547,N_14791);
or UO_1992 (O_1992,N_14686,N_14594);
or UO_1993 (O_1993,N_14906,N_14702);
nand UO_1994 (O_1994,N_14728,N_14886);
and UO_1995 (O_1995,N_14957,N_14933);
nand UO_1996 (O_1996,N_14842,N_14715);
nor UO_1997 (O_1997,N_14754,N_14980);
nor UO_1998 (O_1998,N_14671,N_14997);
and UO_1999 (O_1999,N_14763,N_14736);
endmodule