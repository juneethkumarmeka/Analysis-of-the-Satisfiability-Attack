module basic_3000_30000_3500_60_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1590,In_1080);
and U1 (N_1,In_1267,In_2411);
nor U2 (N_2,In_526,In_1359);
and U3 (N_3,In_17,In_2612);
nor U4 (N_4,In_2243,In_947);
nand U5 (N_5,In_2174,In_1989);
xor U6 (N_6,In_710,In_1765);
and U7 (N_7,In_298,In_1429);
xnor U8 (N_8,In_136,In_2169);
nand U9 (N_9,In_696,In_1568);
nor U10 (N_10,In_1304,In_330);
and U11 (N_11,In_771,In_2880);
and U12 (N_12,In_2781,In_731);
xnor U13 (N_13,In_2493,In_2358);
xor U14 (N_14,In_217,In_921);
nand U15 (N_15,In_169,In_2038);
or U16 (N_16,In_1792,In_2412);
nand U17 (N_17,In_2527,In_549);
nand U18 (N_18,In_98,In_2101);
and U19 (N_19,In_1443,In_334);
and U20 (N_20,In_943,In_901);
xor U21 (N_21,In_1068,In_1285);
or U22 (N_22,In_2553,In_903);
nand U23 (N_23,In_2333,In_2481);
or U24 (N_24,In_855,In_1456);
and U25 (N_25,In_232,In_1261);
xor U26 (N_26,In_2018,In_2548);
or U27 (N_27,In_1274,In_654);
or U28 (N_28,In_97,In_284);
nor U29 (N_29,In_2277,In_867);
or U30 (N_30,In_186,In_1944);
and U31 (N_31,In_2012,In_2646);
nor U32 (N_32,In_2338,In_2124);
or U33 (N_33,In_2276,In_2099);
xnor U34 (N_34,In_1420,In_1868);
or U35 (N_35,In_1287,In_2424);
nand U36 (N_36,In_2793,In_1754);
or U37 (N_37,In_777,In_474);
or U38 (N_38,In_285,In_322);
xor U39 (N_39,In_1288,In_1560);
or U40 (N_40,In_1182,In_1796);
or U41 (N_41,In_627,In_2474);
nor U42 (N_42,In_519,In_2000);
xor U43 (N_43,In_114,In_2479);
nor U44 (N_44,In_2418,In_1004);
nand U45 (N_45,In_1519,In_2465);
or U46 (N_46,In_1451,In_2986);
nand U47 (N_47,In_58,In_2787);
nor U48 (N_48,In_1262,In_2208);
and U49 (N_49,In_2354,In_1840);
xnor U50 (N_50,In_1242,In_119);
nor U51 (N_51,In_806,In_818);
nor U52 (N_52,In_2566,In_1457);
and U53 (N_53,In_1079,In_52);
xor U54 (N_54,In_1331,In_2789);
nand U55 (N_55,In_2336,In_1425);
or U56 (N_56,In_1394,In_1890);
or U57 (N_57,In_329,In_828);
and U58 (N_58,In_96,In_888);
xnor U59 (N_59,In_2438,In_1014);
nand U60 (N_60,In_651,In_1380);
nor U61 (N_61,In_2247,In_335);
nand U62 (N_62,In_2503,In_385);
nor U63 (N_63,In_869,In_2011);
or U64 (N_64,In_2298,In_184);
nor U65 (N_65,In_1298,In_1887);
and U66 (N_66,In_2,In_2305);
nand U67 (N_67,In_410,In_1454);
nor U68 (N_68,In_69,In_2102);
nor U69 (N_69,In_1027,In_573);
nor U70 (N_70,In_1585,In_827);
nand U71 (N_71,In_1985,In_922);
nand U72 (N_72,In_1689,In_1111);
or U73 (N_73,In_387,In_2818);
nor U74 (N_74,In_791,In_1591);
and U75 (N_75,In_2840,In_2025);
xnor U76 (N_76,In_1662,In_1812);
xnor U77 (N_77,In_2579,In_727);
nand U78 (N_78,In_1637,In_1431);
nor U79 (N_79,In_583,In_2398);
or U80 (N_80,In_1946,In_113);
nand U81 (N_81,In_733,In_1151);
nor U82 (N_82,In_1815,In_1373);
or U83 (N_83,In_1473,In_2218);
and U84 (N_84,In_2065,In_879);
nand U85 (N_85,In_1776,In_2064);
or U86 (N_86,In_2052,In_2036);
nor U87 (N_87,In_1609,In_2334);
nor U88 (N_88,In_311,In_674);
or U89 (N_89,In_1066,In_214);
and U90 (N_90,In_688,In_1413);
nand U91 (N_91,In_1337,In_253);
or U92 (N_92,In_1836,In_2794);
nor U93 (N_93,In_820,In_2642);
xnor U94 (N_94,In_912,In_368);
and U95 (N_95,In_2130,In_2197);
nor U96 (N_96,In_1048,In_460);
and U97 (N_97,In_1118,In_178);
nor U98 (N_98,In_2563,In_786);
xor U99 (N_99,In_625,In_540);
nor U100 (N_100,In_2976,In_2999);
or U101 (N_101,In_163,In_487);
or U102 (N_102,In_1500,In_2687);
or U103 (N_103,In_2615,In_269);
xnor U104 (N_104,In_2453,In_109);
nand U105 (N_105,In_751,In_1641);
nand U106 (N_106,In_937,In_1286);
nor U107 (N_107,In_1977,In_1283);
nor U108 (N_108,In_15,In_575);
or U109 (N_109,In_824,In_224);
or U110 (N_110,In_860,In_1496);
nand U111 (N_111,In_913,In_100);
or U112 (N_112,In_476,In_1844);
nor U113 (N_113,In_250,In_395);
xor U114 (N_114,In_963,In_459);
nand U115 (N_115,In_292,In_2511);
nand U116 (N_116,In_356,In_1924);
or U117 (N_117,In_1067,In_837);
or U118 (N_118,In_11,In_2447);
xnor U119 (N_119,In_2349,In_1691);
xnor U120 (N_120,In_453,In_1702);
and U121 (N_121,In_2824,In_2826);
or U122 (N_122,In_2114,In_2881);
nand U123 (N_123,In_1408,In_1990);
or U124 (N_124,In_1667,In_1056);
and U125 (N_125,In_2600,In_2945);
nand U126 (N_126,In_461,In_1140);
and U127 (N_127,In_929,In_2559);
xnor U128 (N_128,In_2293,In_1356);
nand U129 (N_129,In_71,In_588);
xor U130 (N_130,In_1579,In_2737);
nand U131 (N_131,In_2365,In_2386);
nor U132 (N_132,In_1153,In_1130);
xor U133 (N_133,In_2369,In_634);
or U134 (N_134,In_1584,In_545);
and U135 (N_135,In_1763,In_2636);
nand U136 (N_136,In_48,In_1043);
xnor U137 (N_137,In_344,In_1777);
nor U138 (N_138,In_889,In_2068);
and U139 (N_139,In_1994,In_2594);
nor U140 (N_140,In_2931,In_631);
xor U141 (N_141,In_1921,In_1101);
and U142 (N_142,In_760,In_2673);
nand U143 (N_143,In_386,In_744);
xor U144 (N_144,In_278,In_600);
nor U145 (N_145,In_673,In_2454);
nand U146 (N_146,In_1205,In_1538);
and U147 (N_147,In_884,In_146);
and U148 (N_148,In_1319,In_655);
or U149 (N_149,In_231,In_2359);
xnor U150 (N_150,In_2170,In_166);
or U151 (N_151,In_633,In_1406);
or U152 (N_152,In_962,In_944);
and U153 (N_153,In_2764,In_1248);
xnor U154 (N_154,In_1338,In_353);
and U155 (N_155,In_2192,In_2225);
nand U156 (N_156,In_2287,In_2165);
or U157 (N_157,In_2928,In_440);
nor U158 (N_158,In_985,In_939);
and U159 (N_159,In_2907,In_1599);
or U160 (N_160,In_572,In_2806);
xnor U161 (N_161,In_1279,In_2808);
and U162 (N_162,In_1476,In_1759);
or U163 (N_163,In_1612,In_1097);
xnor U164 (N_164,In_925,In_340);
or U165 (N_165,In_1929,In_565);
or U166 (N_166,In_2699,In_582);
or U167 (N_167,In_1016,In_1530);
or U168 (N_168,In_2867,In_1789);
nor U169 (N_169,In_832,In_1136);
nor U170 (N_170,In_1647,In_28);
and U171 (N_171,In_435,In_2959);
and U172 (N_172,In_2416,In_2206);
xnor U173 (N_173,In_2519,In_2091);
and U174 (N_174,In_672,In_1635);
nor U175 (N_175,In_1155,In_2708);
xor U176 (N_176,In_216,In_2421);
nor U177 (N_177,In_2207,In_1104);
xor U178 (N_178,In_2877,In_2326);
nor U179 (N_179,In_892,In_2097);
nor U180 (N_180,In_1170,In_2657);
nor U181 (N_181,In_314,In_1212);
xor U182 (N_182,In_1758,In_2357);
xor U183 (N_183,In_968,In_1349);
or U184 (N_184,In_2490,In_2163);
xor U185 (N_185,In_1088,In_2450);
xor U186 (N_186,In_648,In_341);
or U187 (N_187,In_2397,In_2990);
or U188 (N_188,In_2087,In_873);
nand U189 (N_189,In_1955,In_2848);
and U190 (N_190,In_1762,In_2337);
or U191 (N_191,In_684,In_1709);
and U192 (N_192,In_1638,In_2596);
nor U193 (N_193,In_374,In_1226);
or U194 (N_194,In_809,In_172);
nand U195 (N_195,In_319,In_2142);
nor U196 (N_196,In_2683,In_2984);
xor U197 (N_197,In_381,In_1015);
xor U198 (N_198,In_569,In_2953);
nand U199 (N_199,In_1387,In_2680);
and U200 (N_200,In_1588,In_220);
nand U201 (N_201,In_112,In_1653);
and U202 (N_202,In_2392,In_518);
or U203 (N_203,In_2092,In_2057);
and U204 (N_204,In_2827,In_405);
xnor U205 (N_205,In_1362,In_2788);
and U206 (N_206,In_51,In_323);
and U207 (N_207,In_2987,In_636);
nand U208 (N_208,In_55,In_427);
xnor U209 (N_209,In_1664,In_83);
and U210 (N_210,In_1911,In_612);
and U211 (N_211,In_1305,In_2573);
xnor U212 (N_212,In_605,In_693);
nand U213 (N_213,In_1766,In_854);
xor U214 (N_214,In_1509,In_1845);
nor U215 (N_215,In_21,In_899);
xor U216 (N_216,In_739,In_2194);
nor U217 (N_217,In_520,In_1031);
nor U218 (N_218,In_1650,In_1505);
xnor U219 (N_219,In_975,In_2946);
nand U220 (N_220,In_1736,In_1983);
and U221 (N_221,In_1366,In_2965);
or U222 (N_222,In_1649,In_522);
and U223 (N_223,In_376,In_1448);
nand U224 (N_224,In_2510,In_1619);
nand U225 (N_225,In_1536,In_1995);
or U226 (N_226,In_1761,In_2263);
nand U227 (N_227,In_1094,In_2484);
or U228 (N_228,In_2284,In_874);
nor U229 (N_229,In_2430,In_1106);
and U230 (N_230,In_1144,In_2962);
nor U231 (N_231,In_2295,In_2060);
nand U232 (N_232,In_1225,In_2921);
nand U233 (N_233,In_1369,In_1190);
or U234 (N_234,In_825,In_2279);
nor U235 (N_235,In_2204,In_1992);
xnor U236 (N_236,In_1199,In_2633);
nand U237 (N_237,In_2653,In_2157);
nor U238 (N_238,In_665,In_312);
nor U239 (N_239,In_1823,In_441);
or U240 (N_240,In_2384,In_1901);
or U241 (N_241,In_2193,In_1438);
nor U242 (N_242,In_2339,In_442);
and U243 (N_243,In_974,In_2368);
or U244 (N_244,In_581,In_1577);
nand U245 (N_245,In_1827,In_1959);
nor U246 (N_246,In_713,In_1250);
nor U247 (N_247,In_76,In_2509);
xor U248 (N_248,In_1316,In_2260);
and U249 (N_249,In_2380,In_558);
or U250 (N_250,In_641,In_388);
nand U251 (N_251,In_143,In_140);
nand U252 (N_252,In_2982,In_1208);
nor U253 (N_253,In_1102,In_446);
nor U254 (N_254,In_1883,In_2108);
and U255 (N_255,In_2672,In_2906);
or U256 (N_256,In_1308,In_130);
xor U257 (N_257,In_199,In_2677);
or U258 (N_258,In_270,In_1863);
xor U259 (N_259,In_1401,In_1038);
and U260 (N_260,In_683,In_895);
and U261 (N_261,In_1487,In_2311);
xnor U262 (N_262,In_1085,In_2448);
and U263 (N_263,In_1397,In_1069);
or U264 (N_264,In_258,In_858);
and U265 (N_265,In_2032,In_1514);
and U266 (N_266,In_1341,In_1533);
nor U267 (N_267,In_1978,In_2608);
xnor U268 (N_268,In_1042,In_1324);
and U269 (N_269,In_1122,In_756);
or U270 (N_270,In_2776,In_304);
xor U271 (N_271,In_72,In_1192);
xnor U272 (N_272,In_1698,In_1628);
nor U273 (N_273,In_121,In_1028);
xnor U274 (N_274,In_243,In_370);
nor U275 (N_275,In_2783,In_1180);
xnor U276 (N_276,In_2151,In_406);
nand U277 (N_277,In_2584,In_916);
nor U278 (N_278,In_1292,In_1618);
and U279 (N_279,In_205,In_2229);
or U280 (N_280,In_307,In_1668);
or U281 (N_281,In_2756,In_622);
nand U282 (N_282,In_2909,In_138);
nand U283 (N_283,In_1893,In_2146);
nor U284 (N_284,In_372,In_1488);
nor U285 (N_285,In_265,In_462);
or U286 (N_286,In_394,In_1091);
nor U287 (N_287,In_779,In_2991);
nand U288 (N_288,In_1961,In_2113);
or U289 (N_289,In_475,In_2892);
or U290 (N_290,In_2139,In_559);
xnor U291 (N_291,In_2128,In_2992);
or U292 (N_292,In_1917,In_923);
or U293 (N_293,In_2037,In_1976);
and U294 (N_294,In_1484,In_1072);
nand U295 (N_295,In_1553,In_288);
and U296 (N_296,In_2937,In_1318);
and U297 (N_297,In_2237,In_2977);
nor U298 (N_298,In_1718,In_2288);
and U299 (N_299,In_339,In_1074);
and U300 (N_300,In_983,In_1158);
or U301 (N_301,In_430,In_591);
and U302 (N_302,In_1073,In_1439);
and U303 (N_303,In_1971,In_93);
nand U304 (N_304,In_272,In_663);
xnor U305 (N_305,In_525,In_2785);
nor U306 (N_306,In_2310,In_2825);
nor U307 (N_307,In_347,In_2010);
nand U308 (N_308,In_528,In_2645);
nand U309 (N_309,In_2950,In_2849);
nor U310 (N_310,In_1389,In_1149);
nand U311 (N_311,In_197,In_2890);
or U312 (N_312,In_2956,In_2722);
or U313 (N_313,In_3,In_1113);
nand U314 (N_314,In_592,In_675);
and U315 (N_315,In_2771,In_1051);
xor U316 (N_316,In_1972,In_1573);
nand U317 (N_317,In_1184,In_2241);
nand U318 (N_318,In_2410,In_1851);
and U319 (N_319,In_653,In_1813);
and U320 (N_320,In_2779,In_1854);
and U321 (N_321,In_141,In_1321);
xnor U322 (N_322,In_2993,In_1974);
xor U323 (N_323,In_1541,In_2539);
nand U324 (N_324,In_1903,In_2674);
nor U325 (N_325,In_116,In_2486);
and U326 (N_326,In_1265,In_987);
nand U327 (N_327,In_457,In_2115);
xnor U328 (N_328,In_1703,In_2148);
or U329 (N_329,In_389,In_752);
xnor U330 (N_330,In_1633,In_808);
nor U331 (N_331,In_439,In_2127);
or U332 (N_332,In_1034,In_1760);
nand U333 (N_333,In_772,In_2058);
nand U334 (N_334,In_1816,In_1201);
nor U335 (N_335,In_1059,In_2132);
xnor U336 (N_336,In_1352,In_2883);
and U337 (N_337,In_1630,In_1862);
or U338 (N_338,In_2094,In_871);
and U339 (N_339,In_7,In_2071);
nand U340 (N_340,In_2641,In_2195);
or U341 (N_341,In_1567,In_1729);
xor U342 (N_342,In_1159,In_1108);
xor U343 (N_343,In_746,In_2464);
and U344 (N_344,In_1295,In_630);
and U345 (N_345,In_1041,In_1753);
xnor U346 (N_346,In_2855,In_1866);
or U347 (N_347,In_1023,In_1865);
nand U348 (N_348,In_924,In_382);
xor U349 (N_349,In_705,In_180);
and U350 (N_350,In_539,In_431);
xor U351 (N_351,In_246,In_1859);
nand U352 (N_352,In_2317,In_2552);
nand U353 (N_353,In_2595,In_813);
nor U354 (N_354,In_2210,In_1071);
and U355 (N_355,In_416,In_807);
or U356 (N_356,In_2433,In_2891);
or U357 (N_357,In_1648,In_2766);
nand U358 (N_358,In_1154,In_1679);
and U359 (N_359,In_2182,In_1646);
and U360 (N_360,In_346,In_1234);
xor U361 (N_361,In_1026,In_82);
nand U362 (N_362,In_1755,In_1824);
nor U363 (N_363,In_213,In_979);
and U364 (N_364,In_1000,In_730);
xnor U365 (N_365,In_498,In_81);
nand U366 (N_366,In_715,In_1639);
nor U367 (N_367,In_695,In_2575);
xnor U368 (N_368,In_666,In_2226);
nand U369 (N_369,In_1671,In_2168);
or U370 (N_370,In_2924,In_1938);
or U371 (N_371,In_2420,In_2003);
or U372 (N_372,In_876,In_2807);
nor U373 (N_373,In_129,In_1606);
nor U374 (N_374,In_1818,In_1915);
and U375 (N_375,In_2487,In_1907);
or U376 (N_376,In_719,In_907);
and U377 (N_377,In_229,In_2744);
and U378 (N_378,In_1344,In_2428);
or U379 (N_379,In_1968,In_1426);
nor U380 (N_380,In_1396,In_2658);
xnor U381 (N_381,In_2352,In_1046);
and U382 (N_382,In_2385,In_2030);
or U383 (N_383,In_2665,In_2162);
or U384 (N_384,In_1299,In_183);
and U385 (N_385,In_1945,In_606);
nor U386 (N_386,In_1368,In_1681);
xor U387 (N_387,In_1166,In_646);
nand U388 (N_388,In_2831,In_2692);
nand U389 (N_389,In_302,In_601);
nand U390 (N_390,In_609,In_1284);
or U391 (N_391,In_2245,In_2864);
nor U392 (N_392,In_2703,In_2666);
xor U393 (N_393,In_687,In_1586);
xnor U394 (N_394,In_2440,In_221);
xnor U395 (N_395,In_557,In_1807);
xnor U396 (N_396,In_2521,In_1377);
nand U397 (N_397,In_1922,In_2014);
xor U398 (N_398,In_1297,In_2171);
nand U399 (N_399,In_101,In_532);
and U400 (N_400,In_2270,In_1788);
and U401 (N_401,In_2083,In_2620);
nor U402 (N_402,In_2696,In_996);
or U403 (N_403,In_762,In_1427);
xor U404 (N_404,In_768,In_2353);
nand U405 (N_405,In_403,In_1084);
nor U406 (N_406,In_1460,In_2639);
nor U407 (N_407,In_308,In_1418);
and U408 (N_408,In_433,In_2179);
nand U409 (N_409,In_1914,In_639);
xnor U410 (N_410,In_511,In_2517);
and U411 (N_411,In_1405,In_2387);
xnor U412 (N_412,In_2007,In_1269);
nor U413 (N_413,In_2852,In_2340);
xor U414 (N_414,In_2273,In_1918);
nand U415 (N_415,In_1733,In_967);
xnor U416 (N_416,In_780,In_978);
and U417 (N_417,In_742,In_484);
nand U418 (N_418,In_738,In_623);
or U419 (N_419,In_92,In_1219);
and U420 (N_420,In_2372,In_2224);
nor U421 (N_421,In_620,In_1659);
and U422 (N_422,In_1958,In_1882);
and U423 (N_423,In_126,In_1957);
nor U424 (N_424,In_1187,In_348);
nand U425 (N_425,In_383,In_1675);
and U426 (N_426,In_1544,In_2186);
and U427 (N_427,In_1402,In_906);
nand U428 (N_428,In_2901,In_908);
or U429 (N_429,In_2155,In_2315);
and U430 (N_430,In_86,In_1064);
and U431 (N_431,In_852,In_2478);
or U432 (N_432,In_1363,In_276);
nand U433 (N_433,In_2500,In_2899);
xor U434 (N_434,In_1683,In_2327);
nor U435 (N_435,In_2572,In_470);
xnor U436 (N_436,In_1876,In_2451);
nand U437 (N_437,In_375,In_198);
nor U438 (N_438,In_2655,In_2160);
and U439 (N_439,In_479,In_574);
xor U440 (N_440,In_2396,In_2467);
nand U441 (N_441,In_2274,In_320);
or U442 (N_442,In_645,In_1390);
xnor U443 (N_443,In_2832,In_1078);
xor U444 (N_444,In_1748,In_286);
xnor U445 (N_445,In_282,In_1853);
nor U446 (N_446,In_2107,In_2271);
nor U447 (N_447,In_2916,In_707);
or U448 (N_448,In_753,In_426);
nand U449 (N_449,In_1486,In_2253);
nand U450 (N_450,In_1723,In_652);
nand U451 (N_451,In_154,In_993);
nor U452 (N_452,In_1361,In_1183);
xor U453 (N_453,In_1229,In_2971);
nand U454 (N_454,In_1843,In_2323);
xnor U455 (N_455,In_2862,In_26);
and U456 (N_456,In_1569,In_2203);
nor U457 (N_457,In_2388,In_1083);
nand U458 (N_458,In_1194,In_162);
xor U459 (N_459,In_2498,In_1143);
nand U460 (N_460,In_2020,In_1047);
nand U461 (N_461,In_2502,In_1019);
and U462 (N_462,In_1602,In_524);
and U463 (N_463,In_318,In_2117);
nor U464 (N_464,In_2111,In_782);
or U465 (N_465,In_2660,In_1861);
xnor U466 (N_466,In_1332,In_1597);
xor U467 (N_467,In_399,In_1365);
nand U468 (N_468,In_1172,In_25);
nor U469 (N_469,In_351,In_1139);
nand U470 (N_470,In_2935,In_610);
xnor U471 (N_471,In_160,In_1940);
nor U472 (N_472,In_404,In_2709);
xor U473 (N_473,In_2164,In_640);
nand U474 (N_474,In_2382,In_1741);
nand U475 (N_475,In_1003,In_567);
and U476 (N_476,In_826,In_1065);
nor U477 (N_477,In_1708,In_1704);
and U478 (N_478,In_1554,In_2452);
nor U479 (N_479,In_56,In_632);
or U480 (N_480,In_1701,In_2325);
and U481 (N_481,In_716,In_89);
and U482 (N_482,In_1355,In_393);
or U483 (N_483,In_2266,In_1690);
and U484 (N_484,In_1670,In_697);
or U485 (N_485,In_900,In_1204);
and U486 (N_486,In_1601,In_992);
nor U487 (N_487,In_210,In_2347);
nand U488 (N_488,In_2792,In_2180);
xnor U489 (N_489,In_1873,In_438);
and U490 (N_490,In_1773,In_2044);
or U491 (N_491,In_1858,In_1545);
nand U492 (N_492,In_1459,In_483);
nor U493 (N_493,In_1570,In_2540);
xnor U494 (N_494,In_1479,In_1846);
nor U495 (N_495,In_1221,In_2516);
and U496 (N_496,In_554,In_233);
and U497 (N_497,In_1339,In_1012);
nand U498 (N_498,In_2096,In_817);
or U499 (N_499,In_1749,In_291);
xor U500 (N_500,In_2045,N_417);
nand U501 (N_501,N_202,In_757);
or U502 (N_502,In_2542,In_1987);
nand U503 (N_503,In_2462,In_571);
or U504 (N_504,In_2930,In_1195);
xnor U505 (N_505,In_1657,In_495);
nor U506 (N_506,In_1507,In_2069);
nor U507 (N_507,In_2616,In_321);
nand U508 (N_508,In_244,N_121);
nand U509 (N_509,In_2659,In_481);
nand U510 (N_510,In_796,In_2681);
nand U511 (N_511,In_2834,In_1969);
and U512 (N_512,In_1598,N_151);
xor U513 (N_513,In_2120,In_1804);
and U514 (N_514,In_2413,In_1605);
or U515 (N_515,In_1781,In_2408);
nand U516 (N_516,In_1138,N_28);
and U517 (N_517,In_909,In_1849);
and U518 (N_518,N_282,In_1481);
or U519 (N_519,In_2118,In_1616);
nor U520 (N_520,In_2029,In_2219);
and U521 (N_521,In_464,In_513);
nor U522 (N_522,In_794,N_47);
or U523 (N_523,In_986,N_158);
xor U524 (N_524,In_1993,In_2654);
nor U525 (N_525,In_2131,In_537);
nand U526 (N_526,In_1548,In_473);
nor U527 (N_527,In_373,N_248);
or U528 (N_528,In_2800,In_170);
nand U529 (N_529,N_79,In_2013);
xor U530 (N_530,In_354,N_147);
nand U531 (N_531,In_2076,N_16);
or U532 (N_532,In_2422,In_125);
nor U533 (N_533,In_1611,In_2280);
and U534 (N_534,N_252,In_2439);
nand U535 (N_535,In_2407,In_2585);
and U536 (N_536,N_13,In_502);
nand U537 (N_537,In_1927,In_1163);
and U538 (N_538,In_2866,In_788);
and U539 (N_539,In_658,In_190);
xnor U540 (N_540,In_930,N_281);
nand U541 (N_541,N_344,In_2080);
nand U542 (N_542,In_830,In_997);
or U543 (N_543,In_2985,In_2414);
or U544 (N_544,In_1469,In_2803);
and U545 (N_545,In_767,In_1740);
nand U546 (N_546,In_1705,In_970);
xor U547 (N_547,In_2499,In_68);
xnor U548 (N_548,In_2066,In_2850);
nand U549 (N_549,N_438,In_488);
or U550 (N_550,In_134,In_2640);
nand U551 (N_551,In_2488,In_2587);
or U552 (N_552,In_413,In_1587);
or U553 (N_553,N_349,In_1923);
and U554 (N_554,N_89,In_425);
xnor U555 (N_555,In_75,N_45);
nand U556 (N_556,In_1926,In_2939);
nand U557 (N_557,In_1385,In_2141);
nor U558 (N_558,N_378,In_2150);
nor U559 (N_559,In_1629,N_362);
nor U560 (N_560,In_2294,In_1835);
xor U561 (N_561,In_2248,In_2627);
and U562 (N_562,In_2602,In_268);
nand U563 (N_563,In_2258,In_1092);
or U564 (N_564,N_97,In_2341);
and U565 (N_565,In_749,In_2300);
nand U566 (N_566,In_1948,In_1864);
nor U567 (N_567,N_80,N_387);
xor U568 (N_568,In_946,N_214);
and U569 (N_569,In_2605,In_1164);
nor U570 (N_570,In_2469,N_432);
and U571 (N_571,In_2839,In_2236);
nor U572 (N_572,In_1450,In_1778);
nor U573 (N_573,In_299,In_1712);
nor U574 (N_574,In_102,In_325);
nand U575 (N_575,In_724,In_1191);
nand U576 (N_576,In_882,In_1565);
or U577 (N_577,In_1784,In_2161);
or U578 (N_578,In_1888,In_1045);
and U579 (N_579,N_470,In_2547);
and U580 (N_580,In_562,N_472);
or U581 (N_581,In_1271,In_2167);
and U582 (N_582,In_338,In_1855);
nor U583 (N_583,N_419,In_1526);
or U584 (N_584,In_336,N_167);
nor U585 (N_585,N_446,N_133);
nor U586 (N_586,N_452,In_1124);
xor U587 (N_587,In_2567,In_2482);
nand U588 (N_588,In_1523,In_2137);
xnor U589 (N_589,In_455,N_361);
or U590 (N_590,N_306,In_1435);
xor U591 (N_591,In_1902,In_2628);
nand U592 (N_592,N_40,N_160);
xnor U593 (N_593,In_834,In_1135);
and U594 (N_594,In_548,In_2177);
nor U595 (N_595,In_2817,N_294);
nand U596 (N_596,In_2028,In_174);
xnor U597 (N_597,In_2925,In_1198);
xnor U598 (N_598,In_1826,In_2695);
nor U599 (N_599,In_822,N_261);
or U600 (N_600,In_2304,N_291);
or U601 (N_601,In_773,In_2773);
nor U602 (N_602,In_1800,N_142);
nand U603 (N_603,In_982,N_418);
nor U604 (N_604,N_2,In_42);
and U605 (N_605,In_2942,In_1510);
and U606 (N_606,In_2468,In_2172);
nor U607 (N_607,N_174,In_966);
xor U608 (N_608,In_555,In_401);
or U609 (N_609,In_1774,In_1549);
xnor U610 (N_610,In_364,N_444);
nand U611 (N_611,In_2205,N_139);
and U612 (N_612,N_257,In_2235);
nor U613 (N_613,In_245,In_776);
and U614 (N_614,In_1055,In_2606);
nor U615 (N_615,N_435,In_589);
and U616 (N_616,N_104,In_1906);
xnor U617 (N_617,In_1658,In_2973);
nor U618 (N_618,In_1525,In_2719);
and U619 (N_619,In_2023,In_507);
or U620 (N_620,N_118,N_222);
nand U621 (N_621,In_1428,In_1475);
nor U622 (N_622,N_269,In_1447);
and U623 (N_623,In_2431,In_2811);
nor U624 (N_624,In_1407,In_408);
or U625 (N_625,N_190,In_61);
nor U626 (N_626,In_816,N_279);
nor U627 (N_627,N_57,N_474);
xnor U628 (N_628,N_347,In_2745);
nand U629 (N_629,In_2888,N_92);
and U630 (N_630,In_1176,N_199);
or U631 (N_631,In_2798,In_1512);
nor U632 (N_632,In_2212,In_423);
and U633 (N_633,In_1706,In_712);
xor U634 (N_634,In_277,In_1809);
nor U635 (N_635,In_1539,In_541);
and U636 (N_636,In_24,In_1098);
and U637 (N_637,In_783,In_1445);
nand U638 (N_638,N_210,N_488);
nor U639 (N_639,In_2061,In_227);
xor U640 (N_640,N_408,N_385);
nand U641 (N_641,In_397,In_2185);
and U642 (N_642,N_30,In_54);
or U643 (N_643,N_178,In_2742);
or U644 (N_644,N_366,In_685);
xnor U645 (N_645,In_2835,In_2401);
nand U646 (N_646,In_1325,In_1013);
nand U647 (N_647,In_2138,In_1884);
or U648 (N_648,In_2736,In_2047);
or U649 (N_649,In_706,In_1449);
xnor U650 (N_650,In_1384,In_1309);
nand U651 (N_651,In_2870,In_660);
or U652 (N_652,In_2508,In_972);
nand U653 (N_653,In_412,In_561);
or U654 (N_654,In_736,N_401);
and U655 (N_655,In_2455,In_2590);
nor U656 (N_656,In_1966,In_1687);
nor U657 (N_657,N_264,N_274);
and U658 (N_658,N_336,In_841);
xor U659 (N_659,In_2570,In_90);
and U660 (N_660,In_57,In_2955);
nor U661 (N_661,In_1581,In_1677);
and U662 (N_662,In_449,N_410);
nand U663 (N_663,In_2988,In_1320);
nor U664 (N_664,In_1037,In_862);
or U665 (N_665,N_235,In_447);
nand U666 (N_666,N_414,In_2213);
nand U667 (N_667,In_1471,N_430);
xor U668 (N_668,N_128,In_1623);
and U669 (N_669,In_833,In_94);
or U670 (N_670,N_186,In_2958);
nor U671 (N_671,In_1468,In_1086);
or U672 (N_672,N_215,N_364);
or U673 (N_673,In_2480,In_2176);
nor U674 (N_674,N_426,In_1382);
and U675 (N_675,N_475,In_2927);
nor U676 (N_676,In_875,In_1007);
nor U677 (N_677,In_2292,In_2932);
and U678 (N_678,In_2733,In_1988);
xnor U679 (N_679,N_496,In_1147);
or U680 (N_680,N_255,N_478);
xnor U681 (N_681,In_1424,N_67);
or U682 (N_682,In_2373,In_764);
or U683 (N_683,N_152,In_192);
xnor U684 (N_684,In_2321,In_2529);
and U685 (N_685,In_714,In_1970);
or U686 (N_686,In_2809,In_2694);
or U687 (N_687,N_224,In_456);
nand U688 (N_688,In_815,In_2147);
nand U689 (N_689,N_131,In_2393);
or U690 (N_690,In_1107,N_403);
nor U691 (N_691,In_1409,In_1515);
xor U692 (N_692,In_1772,In_2442);
or U693 (N_693,In_2759,N_10);
nand U694 (N_694,In_521,In_2129);
or U695 (N_695,N_90,In_236);
nand U696 (N_696,In_263,In_306);
nor U697 (N_697,N_0,In_2119);
nor U698 (N_698,In_576,N_148);
xor U699 (N_699,In_2889,In_1213);
or U700 (N_700,In_2701,In_781);
xnor U701 (N_701,N_53,In_2555);
or U702 (N_702,N_168,In_342);
or U703 (N_703,In_196,In_938);
or U704 (N_704,N_290,In_547);
and U705 (N_705,In_1561,In_2048);
nand U706 (N_706,In_711,In_2026);
or U707 (N_707,In_1370,In_802);
and U708 (N_708,In_1672,In_1464);
and U709 (N_709,N_352,In_1595);
nor U710 (N_710,In_785,In_2721);
and U711 (N_711,In_139,In_2233);
or U712 (N_712,In_2140,N_113);
or U713 (N_713,In_702,In_1644);
or U714 (N_714,N_115,In_1886);
or U715 (N_715,N_337,In_611);
nor U716 (N_716,In_251,In_1152);
nor U717 (N_717,N_331,In_703);
nor U718 (N_718,In_1137,In_932);
and U719 (N_719,In_990,N_319);
nor U720 (N_720,In_1388,N_320);
or U721 (N_721,In_85,In_1757);
nor U722 (N_722,In_1764,In_480);
nor U723 (N_723,In_2922,In_2629);
nand U724 (N_724,In_2782,N_342);
and U725 (N_725,In_1133,In_1105);
or U726 (N_726,In_861,In_2319);
and U727 (N_727,In_1642,N_179);
nor U728 (N_728,N_494,In_1880);
nor U729 (N_729,In_1119,In_2868);
nor U730 (N_730,In_1033,In_700);
nand U731 (N_731,N_35,In_2485);
nor U732 (N_732,In_1110,In_1898);
and U733 (N_733,In_2109,In_1819);
or U734 (N_734,In_2718,In_2996);
xor U735 (N_735,N_101,N_476);
xnor U736 (N_736,In_2441,In_1684);
and U737 (N_737,In_436,In_1063);
and U738 (N_738,In_2784,In_1255);
xnor U739 (N_739,N_383,In_2704);
nand U740 (N_740,In_2483,In_857);
nor U741 (N_741,In_2191,In_998);
nand U742 (N_742,In_2860,In_2894);
xor U743 (N_743,In_2152,N_273);
nor U744 (N_744,In_2753,N_216);
nor U745 (N_745,N_50,In_1030);
nand U746 (N_746,In_2897,N_449);
or U747 (N_747,In_2477,In_1342);
and U748 (N_748,In_1714,In_2873);
nor U749 (N_749,In_2915,In_563);
or U750 (N_750,In_1960,In_1724);
nor U751 (N_751,In_132,In_1127);
nor U752 (N_752,In_1148,In_1259);
and U753 (N_753,N_99,In_2126);
and U754 (N_754,In_1527,In_1235);
nor U755 (N_755,In_177,In_988);
or U756 (N_756,N_180,In_1371);
nand U757 (N_757,In_2583,In_2972);
xnor U758 (N_758,In_2379,In_2123);
xnor U759 (N_759,In_690,In_2790);
xnor U760 (N_760,In_247,In_989);
nor U761 (N_761,In_1099,N_379);
nand U762 (N_762,In_2227,In_1266);
and U763 (N_763,N_398,N_125);
or U764 (N_764,In_1001,In_2898);
nand U765 (N_765,In_161,In_2648);
or U766 (N_766,In_2974,In_1949);
or U767 (N_767,N_358,In_2153);
and U768 (N_768,N_194,In_1302);
or U769 (N_769,In_1433,In_949);
and U770 (N_770,In_218,N_272);
or U771 (N_771,In_279,In_2732);
or U772 (N_772,In_99,In_896);
nor U773 (N_773,In_91,In_814);
or U774 (N_774,In_1270,In_2638);
and U775 (N_775,In_2275,In_2621);
and U776 (N_776,In_2727,In_2513);
nand U777 (N_777,In_1141,In_1392);
or U778 (N_778,In_1395,In_398);
xnor U779 (N_779,In_617,In_797);
or U780 (N_780,In_2272,In_1348);
nand U781 (N_781,In_2613,N_498);
xor U782 (N_782,In_2749,N_463);
and U783 (N_783,In_43,In_885);
and U784 (N_784,N_11,In_1608);
or U785 (N_785,In_2940,In_1211);
and U786 (N_786,In_10,In_1202);
xnor U787 (N_787,In_2328,In_2093);
nor U788 (N_788,In_597,In_118);
nor U789 (N_789,In_407,In_2656);
and U790 (N_790,In_1767,In_8);
or U791 (N_791,In_1751,N_441);
or U792 (N_792,In_1333,In_2884);
and U793 (N_793,In_2778,In_1743);
xnor U794 (N_794,N_250,In_1592);
nand U795 (N_795,In_1223,In_800);
or U796 (N_796,In_2090,In_503);
and U797 (N_797,In_845,In_2961);
or U798 (N_798,In_2330,In_1963);
and U799 (N_799,N_3,N_22);
and U800 (N_800,In_1947,N_293);
or U801 (N_801,In_911,In_1323);
and U802 (N_802,In_2728,In_774);
or U803 (N_803,N_395,N_12);
nor U804 (N_804,In_1008,In_1942);
nor U805 (N_805,In_1984,N_150);
or U806 (N_806,In_1794,In_1953);
and U807 (N_807,In_2926,N_374);
or U808 (N_808,N_334,N_469);
nor U809 (N_809,N_271,In_2306);
and U810 (N_810,In_241,N_52);
and U811 (N_811,In_2432,In_2593);
xnor U812 (N_812,In_2805,In_1593);
or U813 (N_813,In_1442,N_58);
xor U814 (N_814,In_1497,In_726);
or U815 (N_815,In_747,In_2079);
or U816 (N_816,In_980,In_84);
nor U817 (N_817,N_345,In_508);
or U818 (N_818,In_358,In_2214);
and U819 (N_819,In_485,In_941);
nor U820 (N_820,In_1498,In_1490);
or U821 (N_821,In_1378,N_9);
nor U822 (N_822,In_1281,In_1177);
nand U823 (N_823,In_1694,N_493);
nand U824 (N_824,In_2743,In_1173);
xor U825 (N_825,In_390,In_1317);
nor U826 (N_826,In_1022,In_267);
nor U827 (N_827,In_257,In_1002);
xnor U828 (N_828,In_516,In_1054);
and U829 (N_829,In_1673,In_1666);
nor U830 (N_830,In_2216,In_1747);
nand U831 (N_831,In_1480,N_303);
nand U832 (N_832,In_1735,In_1872);
xor U833 (N_833,In_969,In_745);
nand U834 (N_834,In_1156,In_1557);
or U835 (N_835,In_2067,In_1126);
xor U836 (N_836,In_1374,N_330);
or U837 (N_837,In_1057,N_377);
nand U838 (N_838,In_2089,In_2324);
xnor U839 (N_839,In_1303,In_2562);
or U840 (N_840,In_1935,In_315);
nand U841 (N_841,In_662,In_458);
xor U842 (N_842,In_1090,In_1412);
nand U843 (N_843,N_481,N_46);
nor U844 (N_844,In_150,In_2632);
nand U845 (N_845,In_956,In_1478);
nor U846 (N_846,N_132,In_2016);
nand U847 (N_847,In_699,In_844);
or U848 (N_848,In_2663,N_297);
or U849 (N_849,N_317,In_850);
nor U850 (N_850,In_2531,In_202);
nand U851 (N_851,In_737,In_1932);
and U852 (N_852,In_1228,N_88);
xor U853 (N_853,N_249,N_36);
or U854 (N_854,In_748,In_2390);
xnor U855 (N_855,In_1474,In_2975);
or U856 (N_856,In_151,In_2853);
and U857 (N_857,In_2537,In_1808);
xor U858 (N_858,In_463,In_357);
and U859 (N_859,In_2712,In_619);
and U860 (N_860,In_2599,In_2551);
or U861 (N_861,In_78,In_621);
or U862 (N_862,In_2550,In_775);
xnor U863 (N_863,In_836,In_1967);
nor U864 (N_864,In_343,In_2603);
nand U865 (N_865,N_308,In_1263);
nand U866 (N_866,In_1786,In_1502);
and U867 (N_867,In_1301,In_155);
xnor U868 (N_868,In_1787,In_2980);
xnor U869 (N_869,In_371,In_647);
xor U870 (N_870,N_55,In_2098);
and U871 (N_871,In_2230,In_2842);
nor U872 (N_872,In_510,In_1411);
nor U873 (N_873,In_2181,In_1169);
and U874 (N_874,N_166,N_87);
xnor U875 (N_875,N_238,In_496);
xor U876 (N_876,In_570,In_1050);
nand U877 (N_877,In_740,In_1874);
nand U878 (N_878,In_1699,In_1185);
and U879 (N_879,In_847,In_2816);
or U880 (N_880,In_2845,In_1710);
and U881 (N_881,In_2664,In_1115);
xor U882 (N_882,In_40,In_1437);
nand U883 (N_883,In_1215,In_1603);
and U884 (N_884,N_84,In_2887);
or U885 (N_885,In_30,N_464);
nand U886 (N_886,N_208,In_2082);
and U887 (N_887,In_2815,In_2088);
nand U888 (N_888,In_1555,In_2458);
nand U889 (N_889,N_312,In_1719);
nor U890 (N_890,In_1006,In_877);
and U891 (N_891,In_2741,N_176);
nor U892 (N_892,In_36,In_1869);
and U893 (N_893,In_2923,In_1803);
and U894 (N_894,In_147,N_465);
or U895 (N_895,In_2581,In_2662);
and U896 (N_896,In_1383,N_371);
or U897 (N_897,N_23,In_692);
and U898 (N_898,In_1233,N_233);
nor U899 (N_899,In_2814,In_465);
and U900 (N_900,N_143,In_878);
nand U901 (N_901,In_1351,In_14);
nor U902 (N_902,In_686,In_2688);
nor U903 (N_903,In_964,In_914);
and U904 (N_904,N_314,N_268);
nand U905 (N_905,N_433,In_1607);
nand U906 (N_906,N_318,In_500);
or U907 (N_907,In_1660,N_239);
xor U908 (N_908,In_1347,In_1707);
xnor U909 (N_909,In_789,N_263);
nor U910 (N_910,In_859,In_2943);
or U911 (N_911,In_1227,In_2370);
nor U912 (N_912,N_284,In_981);
or U913 (N_913,In_153,In_2564);
nor U914 (N_914,In_856,In_1540);
xor U915 (N_915,In_1956,In_2775);
nor U916 (N_916,N_453,In_16);
xnor U917 (N_917,In_1217,N_431);
nand U918 (N_918,In_2437,N_247);
or U919 (N_919,N_254,In_1165);
or U920 (N_920,In_2202,In_2989);
nor U921 (N_921,In_2456,In_2734);
nand U922 (N_922,N_165,N_86);
nand U923 (N_923,In_2598,In_2403);
xor U924 (N_924,In_2024,In_2144);
or U925 (N_925,N_412,In_2588);
xor U926 (N_926,In_1838,N_388);
nand U927 (N_927,In_919,In_2329);
and U928 (N_928,In_2557,In_959);
nor U929 (N_929,In_2843,In_2578);
and U930 (N_930,N_230,In_2434);
nand U931 (N_931,In_863,In_1326);
nand U932 (N_932,In_2078,In_536);
and U933 (N_933,In_428,In_2470);
nand U934 (N_934,In_1962,In_1529);
or U935 (N_935,In_420,In_961);
or U936 (N_936,In_2647,In_2549);
nand U937 (N_937,In_33,In_977);
xnor U938 (N_938,N_295,N_187);
nand U939 (N_939,In_1952,In_2256);
xnor U940 (N_940,N_348,In_2059);
nand U941 (N_941,In_870,In_872);
or U942 (N_942,In_2409,In_189);
or U943 (N_943,N_153,In_2738);
xnor U944 (N_944,N_287,In_2399);
nor U945 (N_945,In_1483,In_2283);
xnor U946 (N_946,In_2211,N_209);
nor U947 (N_947,In_195,In_2905);
or U948 (N_948,In_2571,In_523);
nor U949 (N_949,In_709,In_158);
nand U950 (N_950,In_848,In_2426);
nand U951 (N_951,N_161,In_1768);
or U952 (N_952,N_471,In_1645);
xor U953 (N_953,In_1249,In_1082);
xor U954 (N_954,In_957,In_534);
nor U955 (N_955,In_1693,In_778);
nand U956 (N_956,In_853,In_819);
or U957 (N_957,In_2404,In_1727);
and U958 (N_958,In_2833,In_1626);
and U959 (N_959,In_77,N_114);
nand U960 (N_960,N_311,In_530);
xnor U961 (N_961,In_527,In_2307);
nand U962 (N_962,In_1375,In_1214);
xor U963 (N_963,N_439,In_1446);
xnor U964 (N_964,In_1093,In_482);
nor U965 (N_965,In_1582,In_2021);
xor U966 (N_966,In_2903,In_2039);
or U967 (N_967,N_69,In_1264);
xor U968 (N_968,In_1458,N_20);
nand U969 (N_969,N_212,In_2820);
and U970 (N_970,In_866,N_145);
nand U971 (N_971,In_790,In_363);
and U972 (N_972,N_220,In_313);
nor U973 (N_973,N_499,In_303);
and U974 (N_974,In_2345,In_248);
or U975 (N_975,N_275,N_299);
nor U976 (N_976,In_843,In_424);
nor U977 (N_977,In_1181,In_2027);
and U978 (N_978,In_927,In_1912);
and U979 (N_979,In_194,In_2910);
and U980 (N_980,In_1745,N_105);
xnor U981 (N_981,In_2105,In_2200);
xor U982 (N_982,In_531,In_1580);
and U983 (N_983,In_2591,In_1661);
or U984 (N_984,In_584,In_256);
and U985 (N_985,In_2072,In_1240);
and U986 (N_986,In_1495,In_2331);
xnor U987 (N_987,N_265,In_1620);
xor U988 (N_988,In_1025,In_2528);
and U989 (N_989,In_187,In_2017);
and U990 (N_990,N_427,In_1837);
nor U991 (N_991,In_179,In_1276);
xnor U992 (N_992,N_428,In_493);
xnor U993 (N_993,In_1174,In_324);
xnor U994 (N_994,In_219,In_761);
nor U995 (N_995,In_333,N_226);
and U996 (N_996,In_1795,In_1186);
and U997 (N_997,In_454,N_71);
or U998 (N_998,In_936,N_137);
nand U999 (N_999,In_1241,In_1919);
nand U1000 (N_1000,In_20,In_2046);
xor U1001 (N_1001,In_41,N_102);
nand U1002 (N_1002,In_2250,N_770);
nor U1003 (N_1003,In_955,In_2242);
nand U1004 (N_1004,In_2313,In_1996);
nor U1005 (N_1005,In_2356,N_302);
nand U1006 (N_1006,In_242,In_103);
and U1007 (N_1007,In_477,In_59);
nor U1008 (N_1008,In_47,In_1291);
nor U1009 (N_1009,N_519,In_234);
or U1010 (N_1010,N_738,N_637);
and U1011 (N_1011,In_1998,In_467);
nand U1012 (N_1012,In_928,N_981);
nand U1013 (N_1013,In_305,In_65);
nand U1014 (N_1014,In_1831,N_886);
or U1015 (N_1015,In_1360,In_1273);
nor U1016 (N_1016,N_877,In_203);
xnor U1017 (N_1017,In_108,In_1910);
and U1018 (N_1018,In_1403,N_696);
nor U1019 (N_1019,In_191,N_33);
or U1020 (N_1020,In_2084,N_75);
nand U1021 (N_1021,In_2652,N_579);
or U1022 (N_1022,In_823,In_50);
xnor U1023 (N_1023,N_896,In_1132);
nand U1024 (N_1024,In_1537,In_1518);
and U1025 (N_1025,In_2702,In_2670);
and U1026 (N_1026,N_63,N_182);
nand U1027 (N_1027,In_1343,N_994);
nor U1028 (N_1028,N_556,In_396);
or U1029 (N_1029,In_1289,N_384);
nand U1030 (N_1030,In_1930,In_2522);
and U1031 (N_1031,In_628,N_929);
nand U1032 (N_1032,In_793,In_260);
xnor U1033 (N_1033,In_1870,In_734);
and U1034 (N_1034,In_131,In_331);
and U1035 (N_1035,In_2019,N_778);
nor U1036 (N_1036,N_109,In_2760);
nand U1037 (N_1037,N_506,In_1049);
nand U1038 (N_1038,N_669,In_851);
xor U1039 (N_1039,N_389,In_225);
nor U1040 (N_1040,N_577,N_926);
and U1041 (N_1041,In_1997,N_631);
nor U1042 (N_1042,N_706,N_390);
or U1043 (N_1043,In_1522,In_2847);
nand U1044 (N_1044,In_275,N_138);
and U1045 (N_1045,In_2005,In_1485);
nand U1046 (N_1046,N_951,N_876);
or U1047 (N_1047,In_505,N_566);
nor U1048 (N_1048,N_309,N_136);
nor U1049 (N_1049,In_2051,In_237);
nor U1050 (N_1050,In_2312,N_856);
and U1051 (N_1051,N_867,In_2624);
nor U1052 (N_1052,In_228,N_826);
and U1053 (N_1053,In_1688,N_783);
or U1054 (N_1054,In_2472,In_698);
and U1055 (N_1055,In_1076,In_626);
xor U1056 (N_1056,N_155,In_2104);
xor U1057 (N_1057,N_993,N_141);
or U1058 (N_1058,In_1622,N_454);
xnor U1059 (N_1059,In_1501,In_2534);
and U1060 (N_1060,In_497,In_23);
nand U1061 (N_1061,In_1860,N_760);
or U1062 (N_1062,In_1531,In_283);
nor U1063 (N_1063,In_670,In_886);
xor U1064 (N_1064,In_2457,In_917);
xnor U1065 (N_1065,N_847,In_432);
nor U1066 (N_1066,In_204,In_1559);
and U1067 (N_1067,In_1613,In_1193);
and U1068 (N_1068,In_173,In_1532);
nand U1069 (N_1069,In_2362,N_741);
or U1070 (N_1070,N_402,N_304);
nor U1071 (N_1071,N_947,N_690);
or U1072 (N_1072,N_528,N_500);
nand U1073 (N_1073,In_1018,In_1462);
nand U1074 (N_1074,N_177,N_667);
and U1075 (N_1075,N_779,N_467);
nand U1076 (N_1076,In_2320,N_436);
nor U1077 (N_1077,N_686,N_743);
or U1078 (N_1078,In_369,N_718);
nand U1079 (N_1079,In_411,In_2846);
and U1080 (N_1080,N_861,In_2445);
or U1081 (N_1081,N_405,In_2998);
nor U1082 (N_1082,In_2857,N_193);
nand U1083 (N_1083,In_1416,In_1715);
nand U1084 (N_1084,N_582,N_484);
nand U1085 (N_1085,In_902,N_323);
xor U1086 (N_1086,In_2690,N_731);
and U1087 (N_1087,N_697,In_230);
nor U1088 (N_1088,In_2158,N_935);
or U1089 (N_1089,In_649,In_1131);
or U1090 (N_1090,In_1146,In_883);
and U1091 (N_1091,N_440,In_2644);
or U1092 (N_1092,In_128,N_195);
or U1093 (N_1093,In_255,N_727);
nand U1094 (N_1094,In_167,N_333);
nand U1095 (N_1095,In_360,In_1197);
nand U1096 (N_1096,N_285,In_1793);
or U1097 (N_1097,N_883,N_791);
and U1098 (N_1098,In_1472,In_1077);
nor U1099 (N_1099,N_38,In_2649);
nand U1100 (N_1100,N_231,In_2343);
or U1101 (N_1101,In_1430,In_1722);
xnor U1102 (N_1102,N_539,N_585);
nand U1103 (N_1103,N_283,In_2056);
nor U1104 (N_1104,N_32,N_700);
or U1105 (N_1105,In_556,N_624);
or U1106 (N_1106,In_2761,N_234);
xor U1107 (N_1107,In_578,In_1780);
xor U1108 (N_1108,In_1504,In_211);
nor U1109 (N_1109,In_466,In_729);
or U1110 (N_1110,In_529,In_1891);
or U1111 (N_1111,In_2693,In_1224);
or U1112 (N_1112,N_66,In_2002);
and U1113 (N_1113,N_326,In_2769);
and U1114 (N_1114,In_1121,In_1188);
xnor U1115 (N_1115,N_945,N_798);
xnor U1116 (N_1116,N_713,N_678);
and U1117 (N_1117,In_1506,In_2332);
xor U1118 (N_1118,N_999,In_2427);
and U1119 (N_1119,N_854,In_607);
xor U1120 (N_1120,N_359,In_238);
xor U1121 (N_1121,In_469,In_2222);
nor U1122 (N_1122,N_31,N_429);
xor U1123 (N_1123,In_942,In_758);
xnor U1124 (N_1124,In_2122,In_2893);
nand U1125 (N_1125,N_692,N_267);
nand U1126 (N_1126,In_2705,N_110);
or U1127 (N_1127,In_677,In_2851);
and U1128 (N_1128,N_916,N_985);
nand U1129 (N_1129,In_1852,N_660);
xnor U1130 (N_1130,N_938,In_2791);
or U1131 (N_1131,In_2514,In_1491);
and U1132 (N_1132,In_326,N_838);
nor U1133 (N_1133,In_2837,N_974);
xnor U1134 (N_1134,In_2908,In_2110);
or U1135 (N_1135,In_515,N_758);
xor U1136 (N_1136,N_748,In_2254);
nor U1137 (N_1137,In_2869,In_2515);
xor U1138 (N_1138,In_2473,N_533);
nand U1139 (N_1139,In_1278,In_1928);
nand U1140 (N_1140,In_1563,In_2981);
nor U1141 (N_1141,In_437,In_1934);
xnor U1142 (N_1142,In_1398,N_460);
and U1143 (N_1143,In_2936,In_1625);
nor U1144 (N_1144,N_550,In_2774);
or U1145 (N_1145,N_485,In_2267);
and U1146 (N_1146,In_1280,In_1889);
and U1147 (N_1147,In_1404,N_807);
nand U1148 (N_1148,In_599,N_200);
and U1149 (N_1149,In_2812,In_754);
or U1150 (N_1150,N_122,In_1621);
or U1151 (N_1151,In_0,N_975);
xnor U1152 (N_1152,N_885,N_534);
and U1153 (N_1153,In_421,In_1452);
or U1154 (N_1154,N_561,In_2874);
or U1155 (N_1155,N_386,In_1799);
nand U1156 (N_1156,In_831,In_1716);
and U1157 (N_1157,N_832,In_868);
or U1158 (N_1158,In_2617,N_107);
and U1159 (N_1159,In_1811,N_661);
nand U1160 (N_1160,In_1440,N_749);
or U1161 (N_1161,N_662,In_934);
or U1162 (N_1162,N_657,N_732);
xor U1163 (N_1163,In_543,In_2342);
or U1164 (N_1164,N_913,In_865);
or U1165 (N_1165,N_653,In_2074);
nand U1166 (N_1166,In_1461,In_1805);
nand U1167 (N_1167,In_2747,In_2765);
xor U1168 (N_1168,N_703,In_1770);
nand U1169 (N_1169,N_707,N_942);
nand U1170 (N_1170,N_651,N_455);
and U1171 (N_1171,N_251,In_2752);
or U1172 (N_1172,N_559,In_750);
nand U1173 (N_1173,In_2262,N_943);
nand U1174 (N_1174,N_369,N_170);
or U1175 (N_1175,In_2746,N_140);
xnor U1176 (N_1176,N_375,In_2100);
and U1177 (N_1177,N_466,N_923);
or U1178 (N_1178,In_2706,In_1179);
nor U1179 (N_1179,N_747,In_722);
or U1180 (N_1180,N_381,N_18);
or U1181 (N_1181,N_537,In_1624);
xnor U1182 (N_1182,In_2377,N_524);
or U1183 (N_1183,In_2166,In_1771);
and U1184 (N_1184,N_822,In_842);
and U1185 (N_1185,In_1627,In_182);
nand U1186 (N_1186,In_720,In_32);
and U1187 (N_1187,N_702,In_2489);
nand U1188 (N_1188,In_478,In_765);
and U1189 (N_1189,In_2879,In_1614);
and U1190 (N_1190,N_356,In_6);
nand U1191 (N_1191,N_684,In_2423);
xnor U1192 (N_1192,N_831,In_1508);
or U1193 (N_1193,N_613,In_2651);
and U1194 (N_1194,In_2301,In_262);
or U1195 (N_1195,In_1678,In_2240);
xor U1196 (N_1196,In_2856,N_357);
xnor U1197 (N_1197,N_560,In_1817);
nand U1198 (N_1198,In_2876,N_457);
nor U1199 (N_1199,N_545,In_1336);
nand U1200 (N_1200,N_672,N_882);
nor U1201 (N_1201,N_450,N_363);
and U1202 (N_1202,In_2406,N_189);
or U1203 (N_1203,In_723,In_2697);
or U1204 (N_1204,In_638,In_615);
nand U1205 (N_1205,In_656,N_73);
and U1206 (N_1206,In_2556,N_391);
nor U1207 (N_1207,In_624,N_941);
and U1208 (N_1208,In_838,In_2201);
and U1209 (N_1209,In_1,In_2611);
nor U1210 (N_1210,In_2405,In_795);
nor U1211 (N_1211,N_688,In_1089);
and U1212 (N_1212,In_2520,In_1434);
nand U1213 (N_1213,In_35,N_756);
or U1214 (N_1214,N_871,In_1245);
or U1215 (N_1215,N_979,N_786);
xor U1216 (N_1216,In_350,N_610);
xor U1217 (N_1217,In_743,In_659);
xnor U1218 (N_1218,In_1354,In_1878);
and U1219 (N_1219,In_1275,In_1600);
and U1220 (N_1220,In_1419,In_2863);
nand U1221 (N_1221,In_300,N_574);
nand U1222 (N_1222,In_948,In_249);
xor U1223 (N_1223,N_256,N_752);
or U1224 (N_1224,In_2360,In_1243);
xnor U1225 (N_1225,In_616,In_1021);
nor U1226 (N_1226,N_768,In_361);
and U1227 (N_1227,In_2711,In_1254);
xor U1228 (N_1228,N_666,N_716);
or U1229 (N_1229,N_812,N_744);
and U1230 (N_1230,In_2554,N_677);
xnor U1231 (N_1231,N_644,In_2389);
and U1232 (N_1232,In_1973,In_950);
and U1233 (N_1233,In_1441,In_721);
nor U1234 (N_1234,In_2675,In_2106);
or U1235 (N_1235,In_1410,In_2255);
nor U1236 (N_1236,In_414,In_2249);
xor U1237 (N_1237,N_399,In_2967);
or U1238 (N_1238,N_77,In_95);
nor U1239 (N_1239,In_1791,In_1520);
or U1240 (N_1240,N_784,In_2221);
or U1241 (N_1241,N_396,In_2823);
and U1242 (N_1242,In_1036,In_952);
or U1243 (N_1243,In_769,N_448);
or U1244 (N_1244,N_370,In_1892);
or U1245 (N_1245,In_2698,N_350);
nor U1246 (N_1246,N_298,In_2103);
nand U1247 (N_1247,In_2371,In_1367);
xnor U1248 (N_1248,N_803,N_793);
nand U1249 (N_1249,In_2316,N_810);
xor U1250 (N_1250,N_964,In_419);
nand U1251 (N_1251,N_596,In_1571);
nor U1252 (N_1252,In_2008,In_898);
xnor U1253 (N_1253,In_891,In_566);
nor U1254 (N_1254,N_206,N_632);
nor U1255 (N_1255,N_825,In_2070);
or U1256 (N_1256,In_1790,In_2968);
nor U1257 (N_1257,N_787,In_2361);
nand U1258 (N_1258,In_1636,In_9);
or U1259 (N_1259,In_2795,In_2476);
nor U1260 (N_1260,N_984,In_1654);
and U1261 (N_1261,N_602,N_987);
nor U1262 (N_1262,In_821,N_904);
and U1263 (N_1263,In_679,N_56);
nor U1264 (N_1264,N_996,In_1943);
or U1265 (N_1265,In_2391,In_2582);
or U1266 (N_1266,In_535,In_2523);
or U1267 (N_1267,In_45,In_2268);
or U1268 (N_1268,N_715,In_2715);
or U1269 (N_1269,In_18,In_142);
xor U1270 (N_1270,In_603,In_1676);
or U1271 (N_1271,In_1696,N_674);
nor U1272 (N_1272,In_1253,In_2189);
xor U1273 (N_1273,In_2947,In_1294);
xnor U1274 (N_1274,N_917,In_2730);
xor U1275 (N_1275,N_988,N_725);
xnor U1276 (N_1276,In_2637,In_1822);
nor U1277 (N_1277,N_864,N_982);
or U1278 (N_1278,In_2896,In_805);
nor U1279 (N_1279,In_2173,N_865);
and U1280 (N_1280,In_2053,N_108);
xor U1281 (N_1281,In_1313,In_1350);
nor U1282 (N_1282,N_641,N_37);
nand U1283 (N_1283,In_80,In_499);
and U1284 (N_1284,In_2346,In_784);
and U1285 (N_1285,In_984,N_289);
or U1286 (N_1286,In_34,N_719);
xnor U1287 (N_1287,In_694,N_796);
or U1288 (N_1288,In_2770,In_1830);
and U1289 (N_1289,N_699,N_734);
and U1290 (N_1290,N_164,In_1257);
nor U1291 (N_1291,N_849,N_971);
and U1292 (N_1292,N_483,In_200);
nor U1293 (N_1293,In_2190,In_2054);
and U1294 (N_1294,N_920,In_2133);
nand U1295 (N_1295,N_751,N_874);
or U1296 (N_1296,In_1894,N_586);
or U1297 (N_1297,In_209,N_4);
nor U1298 (N_1298,N_81,In_637);
xnor U1299 (N_1299,N_530,N_609);
or U1300 (N_1300,In_377,In_37);
or U1301 (N_1301,N_244,In_2259);
and U1302 (N_1302,N_407,N_729);
and U1303 (N_1303,In_2929,In_1421);
nor U1304 (N_1304,In_1455,In_1231);
xor U1305 (N_1305,N_423,In_1775);
nor U1306 (N_1306,N_451,In_1828);
nor U1307 (N_1307,In_2278,N_486);
nand U1308 (N_1308,N_733,In_1499);
and U1309 (N_1309,In_1307,In_31);
or U1310 (N_1310,N_372,In_586);
nand U1311 (N_1311,In_2215,N_619);
xnor U1312 (N_1312,N_636,In_2322);
nor U1313 (N_1313,N_592,In_1329);
or U1314 (N_1314,In_2882,N_606);
nand U1315 (N_1315,In_400,In_1128);
and U1316 (N_1316,N_958,In_2917);
xnor U1317 (N_1317,In_310,In_1246);
nor U1318 (N_1318,In_2757,In_2758);
and U1319 (N_1319,In_417,N_924);
and U1320 (N_1320,In_2495,In_171);
xor U1321 (N_1321,In_812,In_560);
or U1322 (N_1322,In_1937,In_1052);
and U1323 (N_1323,N_270,N_895);
xor U1324 (N_1324,In_1643,In_2444);
xor U1325 (N_1325,In_2209,In_1335);
xnor U1326 (N_1326,N_884,N_927);
or U1327 (N_1327,N_621,In_897);
and U1328 (N_1328,In_2378,N_670);
nor U1329 (N_1329,In_2460,N_722);
xor U1330 (N_1330,N_135,In_650);
xnor U1331 (N_1331,N_956,N_62);
nor U1332 (N_1332,N_338,N_616);
nor U1333 (N_1333,In_940,In_1856);
and U1334 (N_1334,N_603,In_2735);
nor U1335 (N_1335,In_1686,In_492);
nor U1336 (N_1336,In_46,N_156);
and U1337 (N_1337,N_184,In_2610);
xnor U1338 (N_1338,N_936,N_420);
nand U1339 (N_1339,N_880,In_418);
and U1340 (N_1340,N_966,In_840);
or U1341 (N_1341,N_197,In_409);
and U1342 (N_1342,N_780,In_1070);
and U1343 (N_1343,In_1189,In_1087);
or U1344 (N_1344,In_995,In_1574);
nor U1345 (N_1345,N_968,N_322);
nor U1346 (N_1346,In_145,In_2836);
and U1347 (N_1347,In_2086,In_2801);
and U1348 (N_1348,In_1268,In_2900);
nand U1349 (N_1349,N_790,N_836);
xor U1350 (N_1350,In_240,In_544);
or U1351 (N_1351,In_999,In_1564);
and U1352 (N_1352,N_888,In_2904);
or U1353 (N_1353,In_2885,N_578);
or U1354 (N_1354,N_663,In_2364);
nand U1355 (N_1355,In_2919,In_846);
and U1356 (N_1356,In_735,In_1296);
or U1357 (N_1357,N_960,In_935);
or U1358 (N_1358,In_2296,N_277);
nor U1359 (N_1359,N_413,In_2754);
nor U1360 (N_1360,N_461,In_1897);
xor U1361 (N_1361,In_2966,In_2383);
nor U1362 (N_1362,In_1832,N_305);
nor U1363 (N_1363,In_2802,In_799);
or U1364 (N_1364,N_425,N_593);
or U1365 (N_1365,In_259,N_415);
and U1366 (N_1366,In_1939,In_2886);
nor U1367 (N_1367,In_2748,In_1558);
or U1368 (N_1368,In_62,In_2724);
and U1369 (N_1369,In_2143,In_1040);
nand U1370 (N_1370,In_309,In_5);
nor U1371 (N_1371,N_902,In_2819);
nand U1372 (N_1372,N_54,In_2350);
nor U1373 (N_1373,In_301,In_1682);
xor U1374 (N_1374,N_497,N_818);
nor U1375 (N_1375,N_26,In_2912);
or U1376 (N_1376,In_669,In_704);
and U1377 (N_1377,N_570,In_2303);
and U1378 (N_1378,In_239,N_907);
xnor U1379 (N_1379,N_529,N_698);
or U1380 (N_1380,N_563,In_2055);
nand U1381 (N_1381,In_546,In_1806);
and U1382 (N_1382,N_116,N_739);
xnor U1383 (N_1383,N_146,In_164);
nand U1384 (N_1384,In_2544,N_552);
nand U1385 (N_1385,In_120,In_2435);
nand U1386 (N_1386,N_491,In_1477);
nand U1387 (N_1387,In_2592,In_2042);
or U1388 (N_1388,N_568,In_1493);
nand U1389 (N_1389,In_2031,N_321);
or U1390 (N_1390,In_598,In_2859);
or U1391 (N_1391,In_70,In_1979);
nand U1392 (N_1392,In_1327,In_366);
or U1393 (N_1393,N_517,In_1857);
nand U1394 (N_1394,N_60,N_591);
nand U1395 (N_1395,In_2895,In_2308);
xor U1396 (N_1396,N_767,N_24);
and U1397 (N_1397,N_397,In_585);
nor U1398 (N_1398,In_105,In_1282);
xnor U1399 (N_1399,In_643,In_918);
and U1400 (N_1400,In_1640,N_213);
nor U1401 (N_1401,In_2344,In_2739);
or U1402 (N_1402,N_259,In_676);
nor U1403 (N_1403,In_289,In_2786);
or U1404 (N_1404,In_839,N_655);
nand U1405 (N_1405,In_2723,In_235);
and U1406 (N_1406,N_100,N_633);
and U1407 (N_1407,N_355,In_2918);
and U1408 (N_1408,In_1632,N_149);
nor U1409 (N_1409,In_1821,N_682);
nand U1410 (N_1410,In_1528,In_1109);
and U1411 (N_1411,N_325,In_359);
nand U1412 (N_1412,N_788,In_953);
and U1413 (N_1413,N_307,In_1422);
and U1414 (N_1414,N_512,In_1999);
xor U1415 (N_1415,N_799,N_324);
nor U1416 (N_1416,In_1695,In_2121);
xnor U1417 (N_1417,In_1905,N_514);
or U1418 (N_1418,N_456,N_774);
and U1419 (N_1419,In_1467,N_952);
or U1420 (N_1420,N_573,In_2717);
xor U1421 (N_1421,In_1908,In_2355);
nor U1422 (N_1422,N_15,In_1310);
or U1423 (N_1423,In_328,N_808);
or U1424 (N_1424,In_849,N_736);
and U1425 (N_1425,N_94,N_409);
nand U1426 (N_1426,N_532,In_550);
nand U1427 (N_1427,N_462,In_1244);
xor U1428 (N_1428,N_117,N_64);
and U1429 (N_1429,In_1725,N_236);
xnor U1430 (N_1430,In_514,In_355);
or U1431 (N_1431,In_2063,N_376);
nor U1432 (N_1432,In_1965,In_1340);
nand U1433 (N_1433,N_781,N_694);
nand U1434 (N_1434,In_2395,In_608);
xor U1435 (N_1435,In_741,In_1732);
and U1436 (N_1436,In_445,In_2033);
and U1437 (N_1437,In_2631,In_1322);
xnor U1438 (N_1438,N_919,In_2799);
or U1439 (N_1439,In_176,N_754);
and U1440 (N_1440,In_392,N_998);
or U1441 (N_1441,In_208,In_1986);
and U1442 (N_1442,In_104,N_106);
nor U1443 (N_1443,In_811,N_642);
nor U1444 (N_1444,In_1256,In_1936);
or U1445 (N_1445,In_644,In_2006);
or U1446 (N_1446,N_933,In_19);
and U1447 (N_1447,In_2034,In_951);
and U1448 (N_1448,In_2145,In_2865);
and U1449 (N_1449,In_2618,In_415);
or U1450 (N_1450,In_2979,N_851);
xnor U1451 (N_1451,N_819,In_1516);
xor U1452 (N_1452,In_2135,In_2234);
nand U1453 (N_1453,N_163,In_1300);
and U1454 (N_1454,In_1386,In_452);
nand U1455 (N_1455,In_613,N_296);
nand U1456 (N_1456,In_1717,N_74);
xor U1457 (N_1457,In_596,N_159);
or U1458 (N_1458,In_2244,In_1583);
xor U1459 (N_1459,N_535,In_2156);
nand U1460 (N_1460,In_110,In_1991);
and U1461 (N_1461,N_693,N_315);
nor U1462 (N_1462,In_835,In_1663);
nor U1463 (N_1463,N_468,In_1311);
xnor U1464 (N_1464,In_1913,N_590);
xnor U1465 (N_1465,In_2545,N_188);
xnor U1466 (N_1466,In_66,N_341);
nor U1467 (N_1467,In_337,In_2400);
nand U1468 (N_1468,In_1312,N_416);
or U1469 (N_1469,In_1178,In_1353);
or U1470 (N_1470,In_165,N_675);
nor U1471 (N_1471,N_201,N_630);
nor U1472 (N_1472,In_1125,In_2264);
or U1473 (N_1473,N_879,In_2286);
xnor U1474 (N_1474,N_542,In_261);
or U1475 (N_1475,In_2750,In_29);
and U1476 (N_1476,N_848,N_720);
and U1477 (N_1477,In_2957,In_2081);
nor U1478 (N_1478,N_584,In_2780);
xor U1479 (N_1479,N_761,N_652);
nor U1480 (N_1480,In_2040,In_954);
nand U1481 (N_1481,N_583,N_811);
or U1482 (N_1482,In_2538,In_1801);
xor U1483 (N_1483,In_657,N_804);
and U1484 (N_1484,In_2949,N_658);
xnor U1485 (N_1485,In_2417,In_2689);
nor U1486 (N_1486,N_340,In_2475);
and U1487 (N_1487,In_2116,In_2536);
or U1488 (N_1488,In_642,N_853);
or U1489 (N_1489,N_894,In_1933);
or U1490 (N_1490,N_858,In_1652);
nor U1491 (N_1491,In_1511,In_1950);
nor U1492 (N_1492,In_2822,N_480);
xor U1493 (N_1493,In_1572,In_1482);
and U1494 (N_1494,N_766,In_1035);
nor U1495 (N_1495,In_64,In_264);
and U1496 (N_1496,N_989,N_912);
nand U1497 (N_1497,N_957,In_63);
xnor U1498 (N_1498,N_42,N_243);
and U1499 (N_1499,N_620,In_2561);
or U1500 (N_1500,In_391,N_313);
nand U1501 (N_1501,In_661,N_1381);
or U1502 (N_1502,N_68,N_557);
xor U1503 (N_1503,N_878,In_384);
or U1504 (N_1504,In_1655,N_1322);
or U1505 (N_1505,N_759,N_599);
and U1506 (N_1506,N_1350,N_855);
or U1507 (N_1507,N_701,N_422);
nor U1508 (N_1508,N_129,In_1756);
or U1509 (N_1509,In_2533,N_824);
nor U1510 (N_1510,In_2601,In_2532);
nor U1511 (N_1511,N_1207,In_1237);
nand U1512 (N_1512,N_1129,N_1254);
nand U1513 (N_1513,N_991,N_614);
nor U1514 (N_1514,N_977,In_755);
or U1515 (N_1515,N_1005,N_223);
nor U1516 (N_1516,N_510,In_1941);
or U1517 (N_1517,N_6,N_800);
nand U1518 (N_1518,In_352,In_1517);
and U1519 (N_1519,N_1013,N_1190);
nor U1520 (N_1520,N_588,N_327);
nor U1521 (N_1521,N_558,N_627);
xor U1522 (N_1522,In_1489,N_1116);
or U1523 (N_1523,In_1400,N_1267);
nor U1524 (N_1524,In_2871,N_329);
or U1525 (N_1525,In_2740,N_595);
nand U1526 (N_1526,In_2314,N_1353);
nand U1527 (N_1527,N_622,In_614);
nand U1528 (N_1528,N_1138,N_1201);
nor U1529 (N_1529,N_640,N_1217);
and U1530 (N_1530,N_1428,N_43);
xor U1531 (N_1531,In_2077,N_120);
xnor U1532 (N_1532,In_1314,In_1345);
and U1533 (N_1533,N_477,N_1124);
or U1534 (N_1534,N_555,In_1216);
xnor U1535 (N_1535,N_1194,N_25);
nand U1536 (N_1536,N_1315,N_1367);
nand U1537 (N_1537,N_664,N_1492);
nand U1538 (N_1538,In_1415,N_1310);
nor U1539 (N_1539,In_1547,N_571);
xnor U1540 (N_1540,N_709,In_732);
or U1541 (N_1541,In_2466,In_1011);
or U1542 (N_1542,N_538,In_1739);
nand U1543 (N_1543,In_1521,N_615);
xnor U1544 (N_1544,N_1480,In_1150);
nor U1545 (N_1545,In_2726,In_422);
and U1546 (N_1546,N_1317,In_1782);
and U1547 (N_1547,In_1391,N_1227);
or U1548 (N_1548,In_1981,In_2049);
xnor U1549 (N_1549,N_1282,In_2461);
xnor U1550 (N_1550,In_2541,N_903);
or U1551 (N_1551,In_2518,N_1109);
or U1552 (N_1552,In_2463,In_193);
nand U1553 (N_1553,N_253,N_1074);
or U1554 (N_1554,In_115,N_507);
or U1555 (N_1555,In_281,In_1982);
and U1556 (N_1556,N_354,In_39);
xor U1557 (N_1557,N_1351,In_691);
xnor U1558 (N_1558,In_2691,N_1467);
nor U1559 (N_1559,In_2729,In_1009);
nor U1560 (N_1560,In_629,N_1061);
and U1561 (N_1561,In_960,N_1081);
xnor U1562 (N_1562,N_278,N_406);
nand U1563 (N_1563,In_2471,In_274);
xor U1564 (N_1564,N_1120,N_1417);
and U1565 (N_1565,In_1552,In_2035);
nor U1566 (N_1566,N_1283,In_137);
or U1567 (N_1567,N_1141,N_260);
or U1568 (N_1568,N_949,In_1881);
xnor U1569 (N_1569,N_954,In_864);
or U1570 (N_1570,In_894,N_1030);
nor U1571 (N_1571,N_1152,In_2661);
nand U1572 (N_1572,N_735,N_946);
nand U1573 (N_1573,N_495,N_1098);
nand U1574 (N_1574,In_1720,In_2269);
nand U1575 (N_1575,In_2136,N_1281);
nor U1576 (N_1576,In_671,N_351);
nor U1577 (N_1577,N_650,N_1246);
nor U1578 (N_1578,In_1820,In_2607);
and U1579 (N_1579,N_1214,N_14);
nor U1580 (N_1580,In_2459,In_2714);
or U1581 (N_1581,N_1135,In_67);
xnor U1582 (N_1582,N_34,In_2952);
or U1583 (N_1583,N_598,N_513);
nor U1584 (N_1584,N_889,N_1003);
and U1585 (N_1585,N_1232,In_123);
nand U1586 (N_1586,In_1239,N_509);
or U1587 (N_1587,In_379,N_567);
or U1588 (N_1588,N_41,N_915);
nor U1589 (N_1589,In_4,N_990);
nor U1590 (N_1590,In_2650,N_820);
and U1591 (N_1591,In_1542,N_1452);
xnor U1592 (N_1592,In_226,N_421);
and U1593 (N_1593,In_1711,N_207);
nor U1594 (N_1594,N_1481,N_1365);
or U1595 (N_1595,N_373,N_1076);
or U1596 (N_1596,In_2838,N_911);
or U1597 (N_1597,In_1543,In_2015);
or U1598 (N_1598,In_1465,In_1900);
and U1599 (N_1599,N_300,N_515);
or U1600 (N_1600,In_1925,N_857);
nor U1601 (N_1601,N_1017,N_1431);
nand U1602 (N_1602,N_1369,N_1142);
nand U1603 (N_1603,N_1108,In_2073);
xor U1604 (N_1604,In_517,N_875);
xnor U1605 (N_1605,N_1421,N_1089);
nand U1606 (N_1606,N_976,N_198);
and U1607 (N_1607,In_188,In_1444);
and U1608 (N_1608,N_1088,In_2810);
and U1609 (N_1609,In_1875,N_1086);
nor U1610 (N_1610,In_1162,In_2496);
or U1611 (N_1611,In_1258,N_1231);
xor U1612 (N_1612,N_773,In_2198);
and U1613 (N_1613,In_1129,N_1011);
or U1614 (N_1614,In_88,N_1334);
and U1615 (N_1615,N_1101,N_1024);
nor U1616 (N_1616,N_932,N_643);
nand U1617 (N_1617,N_394,N_1338);
and U1618 (N_1618,In_2994,N_1050);
nor U1619 (N_1619,N_1128,N_837);
nand U1620 (N_1620,In_2777,In_1631);
and U1621 (N_1621,N_648,N_1489);
or U1622 (N_1622,In_910,N_1060);
and U1623 (N_1623,N_1434,N_1200);
xnor U1624 (N_1624,In_1020,N_1271);
nor U1625 (N_1625,N_1257,N_901);
and U1626 (N_1626,N_676,N_1162);
xor U1627 (N_1627,In_1596,N_124);
nand U1628 (N_1628,In_973,In_2576);
or U1629 (N_1629,In_2804,N_44);
nor U1630 (N_1630,In_1196,In_1842);
or U1631 (N_1631,In_1576,In_1238);
or U1632 (N_1632,N_1158,N_1497);
or U1633 (N_1633,In_881,N_1176);
nand U1634 (N_1634,N_1027,N_1057);
nand U1635 (N_1635,N_872,N_228);
nand U1636 (N_1636,N_1019,N_575);
nor U1637 (N_1637,N_1187,In_280);
nor U1638 (N_1638,N_504,N_508);
or U1639 (N_1639,N_1078,In_590);
xnor U1640 (N_1640,N_1029,In_1615);
nor U1641 (N_1641,N_459,N_1382);
xnor U1642 (N_1642,N_1203,N_1117);
or U1643 (N_1643,N_782,In_1251);
or U1644 (N_1644,In_2685,N_601);
nand U1645 (N_1645,In_106,In_2772);
and U1646 (N_1646,N_1000,N_1325);
nand U1647 (N_1647,N_939,N_554);
xor U1648 (N_1648,N_1303,N_1033);
or U1649 (N_1649,N_541,N_520);
xnor U1650 (N_1650,N_1179,In_689);
xor U1651 (N_1651,In_2948,In_2184);
nand U1652 (N_1652,N_27,N_828);
and U1653 (N_1653,N_191,In_568);
nand U1654 (N_1654,In_2050,N_1055);
xor U1655 (N_1655,In_1005,N_1296);
or U1656 (N_1656,N_1211,In_1463);
nand U1657 (N_1657,In_1453,N_1276);
nand U1658 (N_1658,N_587,N_1484);
or U1659 (N_1659,In_1737,N_157);
and U1660 (N_1660,N_1132,In_2546);
xnor U1661 (N_1661,In_290,N_1172);
xnor U1662 (N_1662,N_1251,N_1002);
or U1663 (N_1663,In_2565,In_1209);
and U1664 (N_1664,N_1197,In_1713);
or U1665 (N_1665,N_1306,N_240);
nand U1666 (N_1666,N_785,In_2829);
and U1667 (N_1667,N_130,N_1261);
nor U1668 (N_1668,N_772,N_1105);
and U1669 (N_1669,In_2875,In_708);
nand U1670 (N_1670,N_1499,N_687);
nor U1671 (N_1671,N_95,N_1279);
nor U1672 (N_1672,In_491,N_1453);
or U1673 (N_1673,In_509,In_1293);
nor U1674 (N_1674,N_1448,In_53);
xnor U1675 (N_1675,N_607,In_2914);
and U1676 (N_1676,In_254,In_2676);
nor U1677 (N_1677,N_1240,In_681);
nand U1678 (N_1678,N_597,N_1479);
xor U1679 (N_1679,In_2686,N_1161);
xor U1680 (N_1680,N_970,N_411);
xnor U1681 (N_1681,N_1359,N_1034);
and U1682 (N_1682,In_564,In_1306);
and U1683 (N_1683,N_1102,In_2821);
xnor U1684 (N_1684,In_2861,In_2796);
and U1685 (N_1685,N_1372,In_2963);
nor U1686 (N_1686,N_656,N_1163);
nor U1687 (N_1687,N_721,N_492);
xor U1688 (N_1688,N_1385,N_301);
nor U1689 (N_1689,In_1364,In_345);
and U1690 (N_1690,N_1407,N_1239);
or U1691 (N_1691,N_91,In_1566);
and U1692 (N_1692,In_327,In_1044);
and U1693 (N_1693,N_679,N_1149);
or U1694 (N_1694,In_2911,N_526);
nor U1695 (N_1695,In_2281,In_111);
xor U1696 (N_1696,In_365,N_777);
nand U1697 (N_1697,N_1447,In_595);
and U1698 (N_1698,N_955,N_1400);
nand U1699 (N_1699,N_205,N_1420);
nor U1700 (N_1700,N_1191,In_2004);
xnor U1701 (N_1701,N_866,N_685);
nor U1702 (N_1702,N_1223,In_1750);
xnor U1703 (N_1703,N_806,N_1196);
xor U1704 (N_1704,N_887,N_1286);
nor U1705 (N_1705,N_869,N_1326);
nor U1706 (N_1706,In_1896,N_905);
xor U1707 (N_1707,In_2265,N_1474);
nor U1708 (N_1708,N_1256,N_1064);
nand U1709 (N_1709,In_2348,N_1386);
xnor U1710 (N_1710,In_1358,In_2751);
and U1711 (N_1711,N_1424,N_997);
xor U1712 (N_1712,In_770,In_2041);
nor U1713 (N_1713,In_1575,In_444);
nor U1714 (N_1714,N_1415,In_725);
or U1715 (N_1715,N_1263,In_1206);
nand U1716 (N_1716,N_551,In_1203);
xnor U1717 (N_1717,N_1169,In_2299);
nand U1718 (N_1718,N_841,N_1457);
nand U1719 (N_1719,N_1210,N_1174);
xnor U1720 (N_1720,N_1487,N_183);
xor U1721 (N_1721,N_1371,N_922);
xnor U1722 (N_1722,N_1260,In_2920);
nand U1723 (N_1723,In_1414,In_1779);
nor U1724 (N_1724,In_2504,In_450);
nand U1725 (N_1725,N_1291,N_639);
and U1726 (N_1726,N_1370,N_78);
xnor U1727 (N_1727,N_1314,N_925);
or U1728 (N_1728,N_1340,N_1311);
nor U1729 (N_1729,N_1028,N_76);
nor U1730 (N_1730,N_1418,In_1120);
nand U1731 (N_1731,N_1486,N_1236);
nand U1732 (N_1732,N_1139,In_2604);
or U1733 (N_1733,N_262,N_730);
and U1734 (N_1734,In_1423,N_776);
and U1735 (N_1735,In_577,In_2710);
and U1736 (N_1736,In_580,In_2668);
nand U1737 (N_1737,In_2619,N_1097);
xnor U1738 (N_1738,N_1171,N_1083);
xor U1739 (N_1739,In_157,N_1166);
xor U1740 (N_1740,In_1556,N_1301);
xor U1741 (N_1741,In_2960,N_85);
nor U1742 (N_1742,N_1490,N_1319);
xnor U1743 (N_1743,In_472,N_834);
nor U1744 (N_1744,N_1344,N_1307);
and U1745 (N_1745,In_2232,N_1045);
nand U1746 (N_1746,N_1373,N_1237);
nor U1747 (N_1747,In_2366,In_2767);
nor U1748 (N_1748,In_2095,N_1248);
xor U1749 (N_1749,N_948,N_647);
xor U1750 (N_1750,In_668,N_611);
or U1751 (N_1751,N_978,In_156);
nand U1752 (N_1752,In_2574,N_445);
or U1753 (N_1753,N_225,In_1871);
xnor U1754 (N_1754,In_2679,In_1834);
nor U1755 (N_1755,In_122,N_646);
nor U1756 (N_1756,In_1810,N_1006);
or U1757 (N_1757,In_587,N_544);
nand U1758 (N_1758,In_2501,N_346);
nand U1759 (N_1759,N_1241,N_245);
nand U1760 (N_1760,In_2512,N_1004);
or U1761 (N_1761,N_1391,N_1459);
and U1762 (N_1762,In_1885,N_892);
xor U1763 (N_1763,N_119,N_1249);
and U1764 (N_1764,In_759,N_961);
or U1765 (N_1765,In_1134,N_1008);
nor U1766 (N_1766,In_1697,N_809);
xnor U1767 (N_1767,N_1022,N_1477);
nand U1768 (N_1768,N_1001,N_1295);
or U1769 (N_1769,In_1674,N_852);
xnor U1770 (N_1770,N_1184,In_1470);
nand U1771 (N_1771,N_1329,N_1094);
xor U1772 (N_1772,N_1041,N_1327);
and U1773 (N_1773,In_667,N_1360);
or U1774 (N_1774,In_933,In_1847);
or U1775 (N_1775,N_1037,In_2944);
xnor U1776 (N_1776,N_1247,In_2394);
or U1777 (N_1777,N_967,N_645);
nand U1778 (N_1778,In_2112,In_1075);
xnor U1779 (N_1779,In_594,N_940);
nor U1780 (N_1780,N_745,In_2085);
nand U1781 (N_1781,N_1189,N_203);
nor U1782 (N_1782,N_490,N_400);
and U1783 (N_1783,N_1328,N_1432);
and U1784 (N_1784,In_215,N_950);
and U1785 (N_1785,N_1183,In_2872);
nand U1786 (N_1786,In_2425,N_1273);
or U1787 (N_1787,In_223,In_1916);
and U1788 (N_1788,In_2375,In_1534);
and U1789 (N_1789,N_266,In_2995);
xnor U1790 (N_1790,In_2125,In_27);
and U1791 (N_1791,In_1017,In_2149);
or U1792 (N_1792,N_531,In_2282);
xnor U1793 (N_1793,N_1445,N_1304);
or U1794 (N_1794,N_1253,In_2828);
nor U1795 (N_1795,In_2285,N_1460);
nand U1796 (N_1796,N_1488,In_1656);
and U1797 (N_1797,N_805,N_1018);
and U1798 (N_1798,N_959,N_1048);
and U1799 (N_1799,N_1090,In_2491);
xor U1800 (N_1800,N_380,In_2402);
and U1801 (N_1801,N_1361,N_1438);
nor U1802 (N_1802,In_1692,N_292);
xnor U1803 (N_1803,N_1178,In_2768);
or U1804 (N_1804,In_1247,In_2290);
xnor U1805 (N_1805,N_1093,N_181);
or U1806 (N_1806,N_218,In_471);
nor U1807 (N_1807,In_1432,N_604);
xor U1808 (N_1808,In_965,N_1377);
nor U1809 (N_1809,In_763,In_144);
nand U1810 (N_1810,In_316,N_908);
and U1811 (N_1811,In_79,N_1387);
or U1812 (N_1812,N_937,In_1103);
nand U1813 (N_1813,N_1485,N_1035);
nor U1814 (N_1814,N_689,N_980);
and U1815 (N_1815,N_458,N_1228);
nor U1816 (N_1816,N_1072,N_1458);
xnor U1817 (N_1817,In_915,N_525);
nor U1818 (N_1818,N_310,N_1259);
xor U1819 (N_1819,N_1243,N_612);
or U1820 (N_1820,N_65,In_2630);
nor U1821 (N_1821,In_798,In_2878);
nand U1822 (N_1822,N_724,In_1746);
nand U1823 (N_1823,In_958,N_775);
nor U1824 (N_1824,N_173,In_512);
xor U1825 (N_1825,N_714,In_1503);
or U1826 (N_1826,In_2609,N_1274);
xor U1827 (N_1827,In_1372,In_1062);
or U1828 (N_1828,In_717,N_1275);
nor U1829 (N_1829,N_629,In_1895);
nor U1830 (N_1830,In_1114,N_1091);
nor U1831 (N_1831,In_2978,N_757);
xor U1832 (N_1832,In_293,N_1235);
or U1833 (N_1833,N_1396,N_1233);
nand U1834 (N_1834,N_96,N_1087);
xnor U1835 (N_1835,In_1879,In_1802);
xnor U1836 (N_1836,N_815,N_1137);
and U1837 (N_1837,N_523,N_723);
and U1838 (N_1838,In_926,N_1204);
nor U1839 (N_1839,N_649,N_840);
nand U1840 (N_1840,N_1242,N_1390);
or U1841 (N_1841,N_258,N_1364);
nand U1842 (N_1842,In_2964,In_551);
or U1843 (N_1843,N_740,In_2577);
nor U1844 (N_1844,N_61,N_1066);
or U1845 (N_1845,N_21,N_335);
and U1846 (N_1846,N_1280,N_1422);
and U1847 (N_1847,N_1079,In_2187);
xnor U1848 (N_1848,In_1116,N_1368);
and U1849 (N_1849,In_1376,In_1145);
and U1850 (N_1850,In_317,N_873);
nand U1851 (N_1851,N_1054,N_712);
xor U1852 (N_1852,N_1252,N_1449);
nor U1853 (N_1853,N_1442,In_367);
and U1854 (N_1854,N_765,In_1466);
xor U1855 (N_1855,In_2682,In_1785);
and U1856 (N_1856,N_1414,In_494);
xnor U1857 (N_1857,N_870,N_842);
and U1858 (N_1858,In_1058,N_1348);
and U1859 (N_1859,In_2188,N_1229);
xnor U1860 (N_1860,N_1318,N_126);
xor U1861 (N_1861,N_1012,N_434);
xor U1862 (N_1862,N_930,In_2297);
nor U1863 (N_1863,In_1328,N_1297);
xor U1864 (N_1864,N_746,N_1482);
nor U1865 (N_1865,N_1416,In_1175);
nand U1866 (N_1866,In_74,In_2217);
or U1867 (N_1867,N_1443,In_1330);
or U1868 (N_1868,In_893,N_845);
and U1869 (N_1869,In_2854,N_863);
nor U1870 (N_1870,In_680,N_962);
or U1871 (N_1871,In_2335,N_1164);
or U1872 (N_1872,N_368,N_1224);
or U1873 (N_1873,N_1192,N_764);
nor U1874 (N_1874,In_2954,In_1232);
and U1875 (N_1875,N_769,N_1264);
nor U1876 (N_1876,N_1168,N_898);
nand U1877 (N_1877,N_1230,In_2231);
nand U1878 (N_1878,N_382,In_2635);
and U1879 (N_1879,N_339,N_1126);
xor U1880 (N_1880,In_678,N_442);
nand U1881 (N_1881,In_538,N_1413);
nor U1882 (N_1882,In_402,In_2238);
or U1883 (N_1883,N_482,N_1268);
or U1884 (N_1884,N_1209,N_1071);
and U1885 (N_1885,N_899,N_1068);
nand U1886 (N_1886,N_654,N_443);
and U1887 (N_1887,N_1333,N_594);
xnor U1888 (N_1888,In_829,In_1290);
and U1889 (N_1889,N_5,In_1357);
nor U1890 (N_1890,In_2560,In_618);
xnor U1891 (N_1891,N_1148,N_797);
or U1892 (N_1892,In_2535,In_2731);
and U1893 (N_1893,In_542,In_1731);
and U1894 (N_1894,In_468,In_1346);
nor U1895 (N_1895,In_2526,N_728);
nor U1896 (N_1896,In_2075,In_448);
and U1897 (N_1897,In_2022,N_1419);
and U1898 (N_1898,N_1380,N_1265);
and U1899 (N_1899,N_794,N_1342);
nand U1900 (N_1900,N_1435,In_2969);
nor U1901 (N_1901,In_2597,N_1);
xnor U1902 (N_1902,In_803,N_1155);
nand U1903 (N_1903,N_316,In_2199);
nand U1904 (N_1904,N_789,In_297);
nor U1905 (N_1905,N_1177,N_1346);
or U1906 (N_1906,In_2246,In_2351);
nor U1907 (N_1907,In_206,N_830);
or U1908 (N_1908,N_1337,In_107);
nand U1909 (N_1909,In_533,In_2001);
xnor U1910 (N_1910,N_1285,N_726);
and U1911 (N_1911,In_1222,N_1498);
nor U1912 (N_1912,In_792,N_1007);
and U1913 (N_1913,In_2558,In_971);
xnor U1914 (N_1914,N_813,N_1389);
and U1915 (N_1915,N_1115,N_928);
or U1916 (N_1916,In_1029,N_1495);
nor U1917 (N_1917,In_1742,In_1393);
nand U1918 (N_1918,In_664,N_1404);
or U1919 (N_1919,N_1299,In_804);
nor U1920 (N_1920,N_1429,In_1546);
or U1921 (N_1921,N_823,In_1524);
nor U1922 (N_1922,N_1216,N_1053);
and U1923 (N_1923,N_1305,In_2858);
nor U1924 (N_1924,N_540,N_1100);
nand U1925 (N_1925,N_829,In_1877);
nor U1926 (N_1926,N_673,N_742);
nor U1927 (N_1927,In_945,In_1100);
or U1928 (N_1928,N_521,N_1451);
and U1929 (N_1929,N_237,In_451);
nor U1930 (N_1930,N_1069,N_360);
nor U1931 (N_1931,In_273,N_103);
nor U1932 (N_1932,N_111,In_1417);
or U1933 (N_1933,N_221,In_1379);
or U1934 (N_1934,N_1044,N_70);
nor U1935 (N_1935,In_490,In_1604);
nand U1936 (N_1936,N_232,N_1106);
nand U1937 (N_1937,N_1426,N_1312);
or U1938 (N_1938,N_1051,N_1021);
xnor U1939 (N_1939,In_635,N_992);
xnor U1940 (N_1940,In_931,N_48);
nand U1941 (N_1941,N_1343,N_1406);
and U1942 (N_1942,In_295,In_1277);
nand U1943 (N_1943,N_518,In_2707);
nor U1944 (N_1944,N_1475,N_1110);
nand U1945 (N_1945,N_522,N_328);
nand U1946 (N_1946,In_2844,N_1255);
and U1947 (N_1947,N_172,In_1096);
and U1948 (N_1948,N_1375,N_1425);
xor U1949 (N_1949,N_49,In_766);
nand U1950 (N_1950,N_217,In_1399);
nor U1951 (N_1951,N_447,N_659);
and U1952 (N_1952,In_2589,N_1095);
or U1953 (N_1953,In_880,In_1829);
xor U1954 (N_1954,N_1104,In_1252);
and U1955 (N_1955,In_552,N_1272);
xnor U1956 (N_1956,N_1026,N_1378);
xor U1957 (N_1957,N_1345,N_835);
nand U1958 (N_1958,In_1798,In_1617);
nor U1959 (N_1959,In_2302,N_1402);
or U1960 (N_1960,N_1388,N_1473);
xor U1961 (N_1961,N_1058,N_29);
and U1962 (N_1962,In_1744,N_705);
nand U1963 (N_1963,In_1610,In_2009);
nor U1964 (N_1964,N_1323,N_1309);
and U1965 (N_1965,N_1040,N_1131);
nor U1966 (N_1966,N_1193,N_1153);
or U1967 (N_1967,In_2363,N_562);
and U1968 (N_1968,In_149,N_1096);
nand U1969 (N_1969,In_2376,In_2902);
nor U1970 (N_1970,In_2220,N_1185);
nand U1971 (N_1971,In_2154,N_1494);
xor U1972 (N_1972,N_1221,In_2568);
xnor U1973 (N_1973,N_1080,N_51);
or U1974 (N_1974,In_1220,In_920);
xnor U1975 (N_1975,In_1931,In_1060);
xnor U1976 (N_1976,In_506,N_546);
nand U1977 (N_1977,In_2625,In_1850);
xor U1978 (N_1978,N_1316,In_2580);
nor U1979 (N_1979,In_2797,N_134);
nor U1980 (N_1980,N_1165,N_1266);
nand U1981 (N_1981,In_378,N_755);
xnor U1982 (N_1982,N_1463,N_1444);
and U1983 (N_1983,In_1160,N_665);
and U1984 (N_1984,In_2062,N_1175);
nand U1985 (N_1985,In_1024,In_13);
nor U1986 (N_1986,N_802,In_49);
and U1987 (N_1987,N_995,N_1277);
nor U1988 (N_1988,N_1202,N_392);
nor U1989 (N_1989,N_404,N_1288);
nand U1990 (N_1990,In_2933,In_2841);
nand U1991 (N_1991,N_1441,N_1151);
and U1992 (N_1992,In_2713,N_839);
or U1993 (N_1993,N_548,In_207);
and U1994 (N_1994,In_501,N_1140);
nor U1995 (N_1995,In_994,In_1783);
xnor U1996 (N_1996,N_881,N_1399);
nand U1997 (N_1997,N_1195,N_353);
xor U1998 (N_1998,N_1123,N_1349);
nor U1999 (N_1999,N_1466,N_1393);
nand U2000 (N_2000,N_1742,N_1455);
or U2001 (N_2001,N_1712,N_1036);
nand U2002 (N_2002,N_1976,N_931);
nand U2003 (N_2003,In_2700,N_1213);
xor U2004 (N_2004,N_1691,N_1689);
nor U2005 (N_2005,N_1493,In_1685);
or U2006 (N_2006,N_625,N_668);
xnor U2007 (N_2007,N_1837,N_1752);
or U2008 (N_2008,N_1219,N_1956);
nor U2009 (N_2009,N_1144,N_1578);
nor U2010 (N_2010,N_1154,N_1205);
nor U2011 (N_2011,In_2725,In_1207);
nand U2012 (N_2012,N_1146,In_1236);
xnor U2013 (N_2013,In_434,N_1979);
nor U2014 (N_2014,N_1244,N_1864);
xor U2015 (N_2015,N_1825,N_1791);
nor U2016 (N_2016,In_2623,N_1496);
nor U2017 (N_2017,N_1454,N_1808);
or U2018 (N_2018,N_1067,N_1650);
nor U2019 (N_2019,N_1563,N_704);
and U2020 (N_2020,N_1743,N_1682);
and U2021 (N_2021,N_1354,N_1596);
or U2022 (N_2022,N_1626,N_1932);
nor U2023 (N_2023,N_1796,N_833);
or U2024 (N_2024,N_1575,N_1939);
and U2025 (N_2025,N_1977,N_1822);
nor U2026 (N_2026,N_1292,N_1947);
nor U2027 (N_2027,N_1332,In_1669);
xnor U2028 (N_2028,N_671,N_1619);
or U2029 (N_2029,N_367,N_1500);
nor U2030 (N_2030,N_1554,In_1218);
or U2031 (N_2031,In_486,N_711);
nor U2032 (N_2032,N_1504,N_1476);
xnor U2033 (N_2033,N_1700,N_944);
or U2034 (N_2034,In_1315,N_1685);
xor U2035 (N_2035,N_1545,N_1828);
or U2036 (N_2036,N_1468,N_1208);
nand U2037 (N_2037,N_1586,N_762);
xnor U2038 (N_2038,In_1492,N_817);
or U2039 (N_2039,In_1825,In_2586);
and U2040 (N_2040,N_1641,N_1841);
nor U2041 (N_2041,N_1509,N_241);
nor U2042 (N_2042,N_1865,N_1948);
nand U2043 (N_2043,N_1324,N_1678);
nor U2044 (N_2044,N_1234,In_2043);
xnor U2045 (N_2045,N_1411,N_1651);
nand U2046 (N_2046,In_1721,N_1802);
nor U2047 (N_2047,N_1082,In_2257);
nand U2048 (N_2048,N_1625,N_343);
nor U2049 (N_2049,N_1680,In_2228);
or U2050 (N_2050,In_2196,N_1518);
nand U2051 (N_2051,N_1649,N_1972);
and U2052 (N_2052,N_1262,N_1674);
and U2053 (N_2053,N_1536,N_1880);
xnor U2054 (N_2054,N_1795,N_1958);
nand U2055 (N_2055,N_1892,N_1788);
xnor U2056 (N_2056,N_8,N_1456);
xor U2057 (N_2057,N_1412,N_1998);
nor U2058 (N_2058,N_1919,N_1996);
nor U2059 (N_2059,N_1830,In_159);
nor U2060 (N_2060,N_986,N_1289);
nor U2061 (N_2061,N_1553,N_827);
xor U2062 (N_2062,N_1949,N_1647);
nand U2063 (N_2063,N_1258,N_1754);
nand U2064 (N_2064,N_1639,N_1125);
and U2065 (N_2065,N_1245,N_1917);
xor U2066 (N_2066,N_1065,N_1898);
and U2067 (N_2067,In_1728,N_1521);
nand U2068 (N_2068,N_1888,N_1820);
or U2069 (N_2069,N_1122,N_934);
or U2070 (N_2070,N_1912,In_252);
and U2071 (N_2071,N_1963,N_1737);
xor U2072 (N_2072,In_2626,N_1711);
or U2073 (N_2073,N_963,N_1510);
or U2074 (N_2074,N_1534,N_1582);
or U2075 (N_2075,N_1198,N_1075);
nand U2076 (N_2076,In_701,N_1654);
xor U2077 (N_2077,N_1629,N_1661);
or U2078 (N_2078,N_1695,In_1550);
or U2079 (N_2079,N_1780,N_1910);
xor U2080 (N_2080,N_1982,N_1968);
nor U2081 (N_2081,In_1123,In_1010);
or U2082 (N_2082,N_850,N_1751);
and U2083 (N_2083,N_1890,In_38);
nor U2084 (N_2084,N_1199,N_1612);
xor U2085 (N_2085,N_1928,N_1590);
nor U2086 (N_2086,N_1895,N_1779);
or U2087 (N_2087,N_1562,N_1733);
or U2088 (N_2088,N_1893,N_1512);
nand U2089 (N_2089,N_1570,N_144);
nor U2090 (N_2090,N_1226,N_1686);
nand U2091 (N_2091,N_1907,N_1580);
xor U2092 (N_2092,N_1507,In_201);
and U2093 (N_2093,N_1719,N_1464);
or U2094 (N_2094,In_2159,N_503);
nand U2095 (N_2095,N_1611,N_1409);
or U2096 (N_2096,N_1084,N_1505);
or U2097 (N_2097,N_1847,In_1171);
nor U2098 (N_2098,N_1430,N_1293);
xnor U2099 (N_2099,N_1757,N_1748);
nand U2100 (N_2100,N_1843,In_2934);
xor U2101 (N_2101,N_680,N_83);
xnor U2102 (N_2102,N_1698,N_1585);
nand U2103 (N_2103,N_516,N_623);
and U2104 (N_2104,In_1839,N_1506);
and U2105 (N_2105,In_2291,N_1839);
xor U2106 (N_2106,N_1491,N_1556);
and U2107 (N_2107,In_44,N_1595);
or U2108 (N_2108,In_1230,N_1362);
or U2109 (N_2109,N_1728,N_1765);
nor U2110 (N_2110,N_1914,N_1167);
and U2111 (N_2111,In_332,In_1980);
or U2112 (N_2112,N_605,N_1924);
and U2113 (N_2113,N_1107,N_1114);
nand U2114 (N_2114,N_953,N_1659);
or U2115 (N_2115,In_1909,N_816);
and U2116 (N_2116,N_1668,N_1112);
or U2117 (N_2117,In_2813,N_1683);
xor U2118 (N_2118,N_1127,N_1778);
nor U2119 (N_2119,N_1587,N_1222);
or U2120 (N_2120,N_1789,N_1383);
or U2121 (N_2121,In_1867,In_2134);
and U2122 (N_2122,N_1602,N_1809);
nor U2123 (N_2123,In_2494,N_1744);
nand U2124 (N_2124,N_1635,In_2178);
and U2125 (N_2125,N_1618,N_969);
or U2126 (N_2126,N_1771,N_681);
nor U2127 (N_2127,N_1799,N_1501);
or U2128 (N_2128,N_1538,N_1878);
nor U2129 (N_2129,N_918,N_1971);
or U2130 (N_2130,N_1571,N_1056);
xor U2131 (N_2131,In_2913,N_1284);
xnor U2132 (N_2132,N_1885,N_1750);
and U2133 (N_2133,N_39,N_1186);
or U2134 (N_2134,In_1168,N_1806);
nor U2135 (N_2135,N_1594,N_1836);
xor U2136 (N_2136,In_504,N_1657);
and U2137 (N_2137,N_1792,N_1039);
xnor U2138 (N_2138,N_1298,N_1860);
nand U2139 (N_2139,N_600,N_634);
nor U2140 (N_2140,N_1760,N_1631);
nand U2141 (N_2141,N_1656,N_1930);
and U2142 (N_2142,N_1833,N_1092);
xnor U2143 (N_2143,N_1063,In_349);
or U2144 (N_2144,N_1693,N_750);
nor U2145 (N_2145,N_489,N_1180);
xnor U2146 (N_2146,N_1598,N_1016);
nand U2147 (N_2147,N_1755,In_2524);
nand U2148 (N_2148,N_1940,N_1552);
nand U2149 (N_2149,N_1920,N_1964);
xor U2150 (N_2150,N_1876,N_1692);
nand U2151 (N_2151,N_1601,N_1990);
nand U2152 (N_2152,N_1250,N_1136);
or U2153 (N_2153,N_196,In_1964);
and U2154 (N_2154,N_1727,N_1574);
and U2155 (N_2155,In_1112,N_890);
and U2156 (N_2156,In_294,N_973);
and U2157 (N_2157,N_1954,In_2374);
nor U2158 (N_2158,In_2667,N_1915);
or U2159 (N_2159,In_1157,N_1352);
nand U2160 (N_2160,In_1436,N_1664);
or U2161 (N_2161,N_1992,N_1665);
nand U2162 (N_2162,N_1845,N_1931);
or U2163 (N_2163,N_1675,N_717);
or U2164 (N_2164,N_1800,In_890);
nor U2165 (N_2165,N_569,N_1522);
xnor U2166 (N_2166,In_212,N_1519);
nor U2167 (N_2167,N_1950,N_1623);
xor U2168 (N_2168,N_914,N_1608);
nand U2169 (N_2169,N_814,N_1777);
or U2170 (N_2170,N_227,N_897);
and U2171 (N_2171,N_1900,N_1085);
nor U2172 (N_2172,In_1535,N_1886);
xnor U2173 (N_2173,N_1716,N_1863);
nand U2174 (N_2174,In_2449,N_1824);
or U2175 (N_2175,N_1991,N_626);
xnor U2176 (N_2176,N_1831,N_1206);
nand U2177 (N_2177,N_1902,N_1745);
nand U2178 (N_2178,N_868,N_1614);
nor U2179 (N_2179,N_1812,In_2309);
xnor U2180 (N_2180,N_1569,In_602);
nor U2181 (N_2181,N_1541,N_710);
and U2182 (N_2182,N_1667,In_2525);
nand U2183 (N_2183,In_168,N_1640);
or U2184 (N_2184,N_1730,N_1861);
and U2185 (N_2185,N_1896,N_1014);
and U2186 (N_2186,N_1133,In_2289);
xor U2187 (N_2187,N_1916,In_2543);
and U2188 (N_2188,N_1989,N_1038);
and U2189 (N_2189,N_843,N_204);
nand U2190 (N_2190,N_1546,N_801);
nand U2191 (N_2191,N_1798,N_1523);
and U2192 (N_2192,N_1713,N_1515);
nor U2193 (N_2193,N_1440,N_1150);
and U2194 (N_2194,N_1883,N_1856);
nor U2195 (N_2195,N_1903,N_1827);
nor U2196 (N_2196,N_1540,N_1547);
xor U2197 (N_2197,N_1600,N_1870);
nor U2198 (N_2198,N_1846,N_1899);
xnor U2199 (N_2199,In_2367,N_860);
or U2200 (N_2200,N_1694,N_565);
nand U2201 (N_2201,N_1995,N_1557);
nor U2202 (N_2202,N_98,N_1768);
or U2203 (N_2203,N_795,N_1627);
and U2204 (N_2204,N_424,In_2970);
and U2205 (N_2205,N_1398,In_1161);
nand U2206 (N_2206,N_1118,N_1810);
nor U2207 (N_2207,In_2941,N_276);
nor U2208 (N_2208,N_1520,In_1381);
nor U2209 (N_2209,In_185,In_991);
and U2210 (N_2210,N_1981,N_1103);
nor U2211 (N_2211,N_1994,N_1469);
nand U2212 (N_2212,In_296,N_1551);
xnor U2213 (N_2213,N_1023,N_1834);
or U2214 (N_2214,In_593,In_1032);
nor U2215 (N_2215,N_1046,N_1781);
nor U2216 (N_2216,N_1607,N_1478);
nor U2217 (N_2217,N_1558,N_1565);
nand U2218 (N_2218,N_1729,N_1508);
nand U2219 (N_2219,N_1739,N_1873);
nor U2220 (N_2220,N_1672,N_1049);
xor U2221 (N_2221,N_1734,N_1592);
nand U2222 (N_2222,N_1572,In_287);
or U2223 (N_2223,N_82,N_1539);
nand U2224 (N_2224,N_1042,N_1736);
nor U2225 (N_2225,N_219,N_1816);
xor U2226 (N_2226,N_1529,N_1662);
xor U2227 (N_2227,N_1278,N_859);
nand U2228 (N_2228,N_1134,In_1665);
nor U2229 (N_2229,In_1904,N_1462);
or U2230 (N_2230,In_1726,In_1848);
xor U2231 (N_2231,N_1671,N_1531);
nand U2232 (N_2232,N_1819,N_1938);
nand U2233 (N_2233,N_1741,N_1908);
nand U2234 (N_2234,In_73,In_1738);
or U2235 (N_2235,N_1967,N_1767);
or U2236 (N_2236,N_1723,N_1461);
nor U2237 (N_2237,N_1677,N_1697);
and U2238 (N_2238,N_1269,N_1960);
or U2239 (N_2239,N_1805,N_1363);
nand U2240 (N_2240,N_1159,N_1997);
xnor U2241 (N_2241,N_1502,N_1170);
or U2242 (N_2242,N_910,N_175);
or U2243 (N_2243,N_1395,N_1379);
and U2244 (N_2244,N_1591,N_1111);
or U2245 (N_2245,N_1944,N_1704);
or U2246 (N_2246,In_2622,N_1740);
and U2247 (N_2247,N_1483,N_17);
nand U2248 (N_2248,N_844,In_266);
or U2249 (N_2249,N_1528,In_1551);
nand U2250 (N_2250,N_1408,N_1218);
or U2251 (N_2251,N_1270,In_117);
nand U2252 (N_2252,N_1423,In_1578);
nor U2253 (N_2253,N_1842,N_1517);
nand U2254 (N_2254,In_1167,N_1709);
nand U2255 (N_2255,N_1904,N_1313);
and U2256 (N_2256,N_1855,In_2223);
nor U2257 (N_2257,N_792,N_1643);
xnor U2258 (N_2258,In_1920,In_787);
and U2259 (N_2259,N_983,N_242);
nor U2260 (N_2260,N_1676,N_162);
nand U2261 (N_2261,N_628,N_1714);
or U2262 (N_2262,N_1999,N_753);
nand U2263 (N_2263,N_1579,N_1644);
nor U2264 (N_2264,N_1433,N_618);
or U2265 (N_2265,In_2239,N_1926);
nand U2266 (N_2266,N_683,N_1181);
and U2267 (N_2267,N_1220,N_1813);
nor U2268 (N_2268,N_1762,In_579);
nand U2269 (N_2269,N_1130,N_479);
nor U2270 (N_2270,N_1962,N_332);
and U2271 (N_2271,N_246,N_1630);
nand U2272 (N_2272,N_1725,N_1772);
nand U2273 (N_2273,In_2569,N_1559);
and U2274 (N_2274,N_1758,N_1437);
or U2275 (N_2275,N_1212,In_2755);
or U2276 (N_2276,N_1394,N_1610);
and U2277 (N_2277,N_1616,N_1160);
nor U2278 (N_2278,In_87,N_1875);
or U2279 (N_2279,N_1537,N_1869);
nor U2280 (N_2280,N_1622,N_900);
nand U2281 (N_2281,N_1696,In_2497);
and U2282 (N_2282,In_2997,N_1636);
or U2283 (N_2283,N_1854,N_1868);
nand U2284 (N_2284,N_1986,N_1606);
and U2285 (N_2285,In_2446,N_1776);
xor U2286 (N_2286,In_443,N_1059);
nor U2287 (N_2287,In_1814,N_1867);
nand U2288 (N_2288,N_502,N_1550);
nor U2289 (N_2289,N_771,In_1594);
nand U2290 (N_2290,N_1533,In_1260);
xnor U2291 (N_2291,N_1188,N_1628);
and U2292 (N_2292,N_1603,N_1043);
or U2293 (N_2293,N_1584,N_1405);
and U2294 (N_2294,In_2671,N_1403);
nand U2295 (N_2295,N_1859,N_1561);
nand U2296 (N_2296,N_1439,In_1975);
or U2297 (N_2297,In_1589,N_1020);
nand U2298 (N_2298,N_1753,N_1573);
nand U2299 (N_2299,N_1514,N_638);
nand U2300 (N_2300,N_1366,N_1634);
xnor U2301 (N_2301,N_1790,In_1734);
nor U2302 (N_2302,N_1710,N_1113);
xnor U2303 (N_2303,N_1897,In_2830);
xnor U2304 (N_2304,N_1588,In_1210);
and U2305 (N_2305,In_1797,N_1025);
xnor U2306 (N_2306,N_1866,N_1663);
nor U2307 (N_2307,In_2763,In_2419);
xnor U2308 (N_2308,N_1735,N_1673);
nand U2309 (N_2309,N_1985,N_1544);
nor U2310 (N_2310,N_1156,In_801);
xnor U2311 (N_2311,N_393,In_2505);
and U2312 (N_2312,N_1599,N_1613);
nand U2313 (N_2313,In_2381,N_1761);
and U2314 (N_2314,N_1701,N_1681);
or U2315 (N_2315,N_543,N_1721);
or U2316 (N_2316,N_1465,In_148);
xnor U2317 (N_2317,N_1576,In_728);
or U2318 (N_2318,N_1182,N_1984);
nand U2319 (N_2319,N_1913,N_505);
xnor U2320 (N_2320,N_691,In_2252);
xnor U2321 (N_2321,N_123,N_1308);
xor U2322 (N_2322,N_1376,N_112);
or U2323 (N_2323,N_1620,In_976);
nand U2324 (N_2324,N_1705,N_1959);
nor U2325 (N_2325,In_1081,N_1666);
nor U2326 (N_2326,N_1637,N_1764);
xor U2327 (N_2327,N_1881,N_1450);
nor U2328 (N_2328,In_271,N_1794);
nor U2329 (N_2329,N_1589,N_1974);
nor U2330 (N_2330,N_286,In_887);
nor U2331 (N_2331,N_1031,N_127);
and U2332 (N_2332,N_1560,In_2443);
and U2333 (N_2333,N_59,N_1225);
nor U2334 (N_2334,N_1535,N_553);
and U2335 (N_2335,N_1357,N_1922);
and U2336 (N_2336,N_1943,N_229);
and U2337 (N_2337,N_821,In_1841);
and U2338 (N_2338,In_1494,N_1401);
nor U2339 (N_2339,In_682,N_1929);
or U2340 (N_2340,N_1786,In_2720);
nand U2341 (N_2341,N_1966,N_1879);
nor U2342 (N_2342,N_1969,N_1320);
or U2343 (N_2343,N_1909,N_1850);
xnor U2344 (N_2344,In_2938,N_549);
and U2345 (N_2345,In_1053,N_1838);
xnor U2346 (N_2346,N_1718,N_1987);
nor U2347 (N_2347,N_1503,N_1852);
or U2348 (N_2348,N_1858,N_1993);
nand U2349 (N_2349,N_1609,In_904);
xor U2350 (N_2350,In_718,N_1787);
nand U2351 (N_2351,In_1951,In_2175);
nand U2352 (N_2352,N_1801,N_1119);
or U2353 (N_2353,N_1906,N_1935);
and U2354 (N_2354,N_1471,N_1951);
nand U2355 (N_2355,N_1525,In_380);
nor U2356 (N_2356,N_1032,N_1374);
nor U2357 (N_2357,N_1526,N_589);
and U2358 (N_2358,N_1882,In_2506);
and U2359 (N_2359,N_511,In_2634);
xor U2360 (N_2360,N_1294,N_1961);
or U2361 (N_2361,N_1957,In_1730);
nand U2362 (N_2362,In_175,N_1568);
or U2363 (N_2363,N_1911,N_1872);
and U2364 (N_2364,N_192,N_1918);
and U2365 (N_2365,N_1707,In_2429);
xnor U2366 (N_2366,In_1634,N_1604);
and U2367 (N_2367,N_1832,N_288);
nor U2368 (N_2368,N_1980,N_1720);
nand U2369 (N_2369,N_547,In_124);
or U2370 (N_2370,N_1669,N_1953);
or U2371 (N_2371,N_1699,N_1516);
xnor U2372 (N_2372,N_1384,N_1901);
xnor U2373 (N_2373,N_1410,N_1703);
nor U2374 (N_2374,N_1642,N_1143);
or U2375 (N_2375,N_862,N_1321);
or U2376 (N_2376,N_1077,N_1874);
or U2377 (N_2377,N_1891,In_12);
xnor U2378 (N_2378,N_1746,N_1527);
xnor U2379 (N_2379,In_152,N_1670);
nand U2380 (N_2380,N_72,N_617);
and U2381 (N_2381,N_708,N_1062);
and U2382 (N_2382,In_1680,N_1652);
nand U2383 (N_2383,N_906,N_1923);
or U2384 (N_2384,N_909,N_1238);
nand U2385 (N_2385,N_1624,N_1446);
nor U2386 (N_2386,N_1392,In_1142);
nand U2387 (N_2387,N_1355,In_2678);
nand U2388 (N_2388,In_604,In_1899);
xnor U2389 (N_2389,N_1427,In_222);
nand U2390 (N_2390,N_1638,In_1039);
or U2391 (N_2391,N_965,N_1356);
and U2392 (N_2392,N_1593,N_1287);
or U2393 (N_2393,In_2261,In_1095);
nor U2394 (N_2394,N_921,N_1532);
nor U2395 (N_2395,In_2492,In_429);
or U2396 (N_2396,N_487,N_1717);
xnor U2397 (N_2397,N_1010,N_1581);
and U2398 (N_2398,N_1555,N_1782);
xnor U2399 (N_2399,In_2507,N_1988);
nand U2400 (N_2400,In_553,N_1783);
nand U2401 (N_2401,N_1769,N_1804);
and U2402 (N_2402,N_1679,N_7);
xnor U2403 (N_2403,N_1814,N_1542);
nand U2404 (N_2404,N_1965,N_1763);
or U2405 (N_2405,N_1687,N_1853);
or U2406 (N_2406,In_2318,N_1633);
or U2407 (N_2407,In_2183,N_1121);
xnor U2408 (N_2408,N_1936,N_1347);
and U2409 (N_2409,N_1894,N_1621);
or U2410 (N_2410,N_1811,N_1341);
nor U2411 (N_2411,N_1770,N_1818);
nand U2412 (N_2412,N_1331,N_635);
or U2413 (N_2413,N_763,N_185);
nor U2414 (N_2414,N_1945,In_135);
or U2415 (N_2415,N_1793,N_608);
or U2416 (N_2416,N_1070,N_1871);
xnor U2417 (N_2417,In_2669,N_1823);
or U2418 (N_2418,N_1844,In_1651);
or U2419 (N_2419,N_893,In_362);
xnor U2420 (N_2420,N_1983,In_1117);
nand U2421 (N_2421,In_1513,N_1513);
nor U2422 (N_2422,N_1862,N_1955);
xnor U2423 (N_2423,In_181,In_1954);
and U2424 (N_2424,N_501,N_1690);
nand U2425 (N_2425,N_1583,N_695);
xor U2426 (N_2426,N_1889,N_581);
nor U2427 (N_2427,N_1548,N_1829);
nor U2428 (N_2428,N_1978,In_2684);
xor U2429 (N_2429,N_1884,N_211);
nor U2430 (N_2430,N_1336,N_1702);
or U2431 (N_2431,N_1759,N_1927);
nand U2432 (N_2432,N_1731,N_1684);
nand U2433 (N_2433,N_1877,In_2716);
nand U2434 (N_2434,In_2415,In_2643);
nand U2435 (N_2435,N_1339,In_1200);
nor U2436 (N_2436,N_1925,In_1752);
xor U2437 (N_2437,N_1658,N_737);
and U2438 (N_2438,N_1784,In_2251);
and U2439 (N_2439,N_572,In_2614);
or U2440 (N_2440,N_1732,N_576);
xor U2441 (N_2441,In_22,N_1848);
nand U2442 (N_2442,N_1826,N_1887);
or U2443 (N_2443,N_1747,N_1803);
nand U2444 (N_2444,N_1145,N_1300);
nor U2445 (N_2445,In_2436,N_1302);
nor U2446 (N_2446,N_1335,In_2951);
nand U2447 (N_2447,In_60,N_536);
or U2448 (N_2448,N_1605,N_1566);
nor U2449 (N_2449,In_1700,N_1738);
or U2450 (N_2450,N_1397,N_527);
nand U2451 (N_2451,N_1933,N_1946);
nand U2452 (N_2452,N_1597,N_154);
and U2453 (N_2453,N_1358,N_171);
and U2454 (N_2454,N_1785,N_1436);
or U2455 (N_2455,N_580,N_437);
or U2456 (N_2456,N_1632,N_1934);
xnor U2457 (N_2457,In_2762,N_1815);
or U2458 (N_2458,N_1942,In_127);
nand U2459 (N_2459,N_169,In_905);
or U2460 (N_2460,N_1009,N_1724);
and U2461 (N_2461,N_1708,N_1715);
nand U2462 (N_2462,N_1564,N_280);
nand U2463 (N_2463,In_133,N_1821);
or U2464 (N_2464,N_1645,N_972);
or U2465 (N_2465,N_1937,N_1726);
and U2466 (N_2466,N_93,N_1617);
and U2467 (N_2467,N_1756,N_1722);
nand U2468 (N_2468,N_1849,In_2983);
or U2469 (N_2469,N_1660,In_1334);
xnor U2470 (N_2470,N_1290,N_1524);
and U2471 (N_2471,N_365,N_1648);
or U2472 (N_2472,In_2530,N_1807);
or U2473 (N_2473,N_1851,N_1973);
and U2474 (N_2474,N_1905,In_1562);
nand U2475 (N_2475,In_1769,N_1797);
nor U2476 (N_2476,N_1615,N_1775);
xor U2477 (N_2477,N_1015,N_1157);
nor U2478 (N_2478,N_1646,N_1173);
or U2479 (N_2479,N_1706,N_1549);
or U2480 (N_2480,N_1470,N_891);
nor U2481 (N_2481,N_1099,N_1543);
nor U2482 (N_2482,N_1511,N_1817);
and U2483 (N_2483,N_846,N_1073);
nor U2484 (N_2484,N_1921,N_564);
and U2485 (N_2485,N_1472,N_1655);
nand U2486 (N_2486,In_1061,N_1215);
or U2487 (N_2487,N_473,N_1749);
nor U2488 (N_2488,N_1774,N_1577);
nor U2489 (N_2489,N_1857,N_1147);
nor U2490 (N_2490,N_1840,N_1975);
nand U2491 (N_2491,N_1941,N_1835);
nor U2492 (N_2492,N_1766,N_1653);
nand U2493 (N_2493,N_1047,In_489);
nand U2494 (N_2494,N_1330,N_1970);
or U2495 (N_2495,N_1567,N_1530);
or U2496 (N_2496,In_810,N_19);
nand U2497 (N_2497,N_1052,In_1272);
nor U2498 (N_2498,N_1688,N_1952);
nand U2499 (N_2499,In_1833,N_1773);
nor U2500 (N_2500,N_2048,N_2269);
nor U2501 (N_2501,N_2240,N_2257);
or U2502 (N_2502,N_2029,N_2049);
nor U2503 (N_2503,N_2180,N_2274);
nand U2504 (N_2504,N_2174,N_2143);
and U2505 (N_2505,N_2043,N_2056);
and U2506 (N_2506,N_2051,N_2114);
and U2507 (N_2507,N_2386,N_2271);
or U2508 (N_2508,N_2395,N_2241);
nand U2509 (N_2509,N_2231,N_2286);
and U2510 (N_2510,N_2443,N_2107);
nand U2511 (N_2511,N_2467,N_2189);
nor U2512 (N_2512,N_2208,N_2102);
and U2513 (N_2513,N_2431,N_2360);
and U2514 (N_2514,N_2116,N_2289);
xor U2515 (N_2515,N_2325,N_2130);
nand U2516 (N_2516,N_2454,N_2217);
and U2517 (N_2517,N_2017,N_2003);
xnor U2518 (N_2518,N_2005,N_2149);
xnor U2519 (N_2519,N_2178,N_2158);
nand U2520 (N_2520,N_2153,N_2299);
nor U2521 (N_2521,N_2383,N_2479);
nor U2522 (N_2522,N_2193,N_2280);
nand U2523 (N_2523,N_2027,N_2119);
nand U2524 (N_2524,N_2080,N_2447);
nor U2525 (N_2525,N_2076,N_2261);
xnor U2526 (N_2526,N_2159,N_2310);
nor U2527 (N_2527,N_2334,N_2046);
nand U2528 (N_2528,N_2109,N_2446);
nor U2529 (N_2529,N_2074,N_2175);
nor U2530 (N_2530,N_2246,N_2353);
and U2531 (N_2531,N_2319,N_2282);
nand U2532 (N_2532,N_2172,N_2326);
nand U2533 (N_2533,N_2087,N_2458);
nand U2534 (N_2534,N_2224,N_2053);
nand U2535 (N_2535,N_2018,N_2419);
nor U2536 (N_2536,N_2373,N_2062);
or U2537 (N_2537,N_2389,N_2044);
nor U2538 (N_2538,N_2335,N_2132);
nand U2539 (N_2539,N_2392,N_2259);
nor U2540 (N_2540,N_2409,N_2004);
and U2541 (N_2541,N_2456,N_2230);
and U2542 (N_2542,N_2434,N_2337);
xnor U2543 (N_2543,N_2380,N_2264);
nor U2544 (N_2544,N_2059,N_2416);
or U2545 (N_2545,N_2463,N_2105);
nor U2546 (N_2546,N_2472,N_2369);
xnor U2547 (N_2547,N_2055,N_2313);
and U2548 (N_2548,N_2081,N_2393);
or U2549 (N_2549,N_2290,N_2164);
and U2550 (N_2550,N_2331,N_2417);
nand U2551 (N_2551,N_2001,N_2405);
nand U2552 (N_2552,N_2077,N_2427);
and U2553 (N_2553,N_2491,N_2414);
nor U2554 (N_2554,N_2209,N_2041);
and U2555 (N_2555,N_2420,N_2365);
nor U2556 (N_2556,N_2212,N_2268);
nor U2557 (N_2557,N_2254,N_2407);
and U2558 (N_2558,N_2194,N_2247);
and U2559 (N_2559,N_2453,N_2021);
and U2560 (N_2560,N_2204,N_2113);
xnor U2561 (N_2561,N_2430,N_2371);
nand U2562 (N_2562,N_2484,N_2078);
or U2563 (N_2563,N_2281,N_2002);
nor U2564 (N_2564,N_2296,N_2378);
xor U2565 (N_2565,N_2134,N_2066);
and U2566 (N_2566,N_2201,N_2276);
xnor U2567 (N_2567,N_2010,N_2375);
or U2568 (N_2568,N_2390,N_2303);
and U2569 (N_2569,N_2352,N_2112);
and U2570 (N_2570,N_2169,N_2070);
and U2571 (N_2571,N_2318,N_2258);
nor U2572 (N_2572,N_2450,N_2161);
nor U2573 (N_2573,N_2069,N_2232);
nor U2574 (N_2574,N_2357,N_2412);
nand U2575 (N_2575,N_2248,N_2227);
nand U2576 (N_2576,N_2031,N_2411);
nor U2577 (N_2577,N_2439,N_2157);
and U2578 (N_2578,N_2354,N_2493);
or U2579 (N_2579,N_2129,N_2034);
or U2580 (N_2580,N_2368,N_2497);
or U2581 (N_2581,N_2477,N_2014);
nor U2582 (N_2582,N_2495,N_2327);
and U2583 (N_2583,N_2460,N_2347);
nand U2584 (N_2584,N_2328,N_2060);
and U2585 (N_2585,N_2302,N_2263);
xor U2586 (N_2586,N_2402,N_2103);
or U2587 (N_2587,N_2061,N_2473);
nor U2588 (N_2588,N_2344,N_2391);
nand U2589 (N_2589,N_2421,N_2401);
xor U2590 (N_2590,N_2128,N_2397);
and U2591 (N_2591,N_2323,N_2451);
and U2592 (N_2592,N_2410,N_2287);
nor U2593 (N_2593,N_2297,N_2091);
or U2594 (N_2594,N_2432,N_2184);
nor U2595 (N_2595,N_2213,N_2220);
and U2596 (N_2596,N_2016,N_2028);
xor U2597 (N_2597,N_2396,N_2173);
and U2598 (N_2598,N_2162,N_2433);
nand U2599 (N_2599,N_2403,N_2082);
nor U2600 (N_2600,N_2415,N_2118);
nor U2601 (N_2601,N_2144,N_2047);
and U2602 (N_2602,N_2171,N_2320);
or U2603 (N_2603,N_2340,N_2481);
and U2604 (N_2604,N_2349,N_2355);
or U2605 (N_2605,N_2022,N_2131);
nand U2606 (N_2606,N_2448,N_2306);
nor U2607 (N_2607,N_2475,N_2272);
or U2608 (N_2608,N_2015,N_2309);
or U2609 (N_2609,N_2007,N_2223);
xor U2610 (N_2610,N_2499,N_2202);
nor U2611 (N_2611,N_2457,N_2452);
and U2612 (N_2612,N_2459,N_2238);
nor U2613 (N_2613,N_2152,N_2185);
nand U2614 (N_2614,N_2404,N_2345);
nor U2615 (N_2615,N_2426,N_2425);
xnor U2616 (N_2616,N_2093,N_2068);
xor U2617 (N_2617,N_2214,N_2123);
nor U2618 (N_2618,N_2233,N_2110);
nand U2619 (N_2619,N_2301,N_2229);
nor U2620 (N_2620,N_2079,N_2145);
or U2621 (N_2621,N_2435,N_2058);
and U2622 (N_2622,N_2200,N_2064);
xnor U2623 (N_2623,N_2124,N_2215);
or U2624 (N_2624,N_2364,N_2097);
or U2625 (N_2625,N_2418,N_2026);
nor U2626 (N_2626,N_2199,N_2490);
xnor U2627 (N_2627,N_2099,N_2298);
nand U2628 (N_2628,N_2422,N_2492);
xor U2629 (N_2629,N_2137,N_2198);
nand U2630 (N_2630,N_2476,N_2210);
and U2631 (N_2631,N_2317,N_2341);
xor U2632 (N_2632,N_2376,N_2275);
nor U2633 (N_2633,N_2192,N_2032);
nand U2634 (N_2634,N_2339,N_2382);
and U2635 (N_2635,N_2139,N_2398);
and U2636 (N_2636,N_2019,N_2350);
nor U2637 (N_2637,N_2075,N_2181);
nor U2638 (N_2638,N_2088,N_2030);
xor U2639 (N_2639,N_2024,N_2000);
nor U2640 (N_2640,N_2251,N_2179);
nand U2641 (N_2641,N_2195,N_2045);
or U2642 (N_2642,N_2218,N_2265);
and U2643 (N_2643,N_2065,N_2293);
xnor U2644 (N_2644,N_2182,N_2284);
xor U2645 (N_2645,N_2141,N_2150);
nand U2646 (N_2646,N_2073,N_2226);
xnor U2647 (N_2647,N_2020,N_2106);
nor U2648 (N_2648,N_2166,N_2489);
xor U2649 (N_2649,N_2314,N_2108);
xnor U2650 (N_2650,N_2142,N_2387);
nand U2651 (N_2651,N_2351,N_2071);
nor U2652 (N_2652,N_2362,N_2140);
xnor U2653 (N_2653,N_2285,N_2363);
nand U2654 (N_2654,N_2009,N_2312);
nor U2655 (N_2655,N_2190,N_2292);
nor U2656 (N_2656,N_2243,N_2307);
nand U2657 (N_2657,N_2321,N_2168);
and U2658 (N_2658,N_2260,N_2085);
nor U2659 (N_2659,N_2438,N_2205);
xnor U2660 (N_2660,N_2316,N_2191);
nand U2661 (N_2661,N_2187,N_2366);
and U2662 (N_2662,N_2277,N_2167);
nand U2663 (N_2663,N_2278,N_2372);
nor U2664 (N_2664,N_2428,N_2295);
and U2665 (N_2665,N_2008,N_2449);
nor U2666 (N_2666,N_2120,N_2235);
xor U2667 (N_2667,N_2206,N_2133);
and U2668 (N_2668,N_2092,N_2104);
xor U2669 (N_2669,N_2012,N_2474);
or U2670 (N_2670,N_2083,N_2222);
nand U2671 (N_2671,N_2154,N_2203);
nor U2672 (N_2672,N_2267,N_2468);
xor U2673 (N_2673,N_2057,N_2388);
nand U2674 (N_2674,N_2244,N_2135);
xnor U2675 (N_2675,N_2332,N_2115);
nor U2676 (N_2676,N_2485,N_2394);
or U2677 (N_2677,N_2160,N_2121);
nand U2678 (N_2678,N_2408,N_2186);
nand U2679 (N_2679,N_2177,N_2288);
nand U2680 (N_2680,N_2228,N_2465);
and U2681 (N_2681,N_2336,N_2305);
or U2682 (N_2682,N_2219,N_2245);
nand U2683 (N_2683,N_2283,N_2252);
and U2684 (N_2684,N_2111,N_2338);
and U2685 (N_2685,N_2216,N_2399);
nor U2686 (N_2686,N_2126,N_2471);
or U2687 (N_2687,N_2165,N_2480);
or U2688 (N_2688,N_2013,N_2063);
nor U2689 (N_2689,N_2455,N_2170);
or U2690 (N_2690,N_2122,N_2176);
nor U2691 (N_2691,N_2052,N_2033);
nor U2692 (N_2692,N_2308,N_2072);
and U2693 (N_2693,N_2279,N_2006);
xnor U2694 (N_2694,N_2155,N_2211);
or U2695 (N_2695,N_2042,N_2342);
or U2696 (N_2696,N_2196,N_2400);
nor U2697 (N_2697,N_2098,N_2406);
or U2698 (N_2698,N_2300,N_2482);
nor U2699 (N_2699,N_2011,N_2094);
nor U2700 (N_2700,N_2225,N_2035);
nand U2701 (N_2701,N_2151,N_2429);
and U2702 (N_2702,N_2040,N_2067);
and U2703 (N_2703,N_2294,N_2377);
xnor U2704 (N_2704,N_2125,N_2221);
or U2705 (N_2705,N_2037,N_2462);
and U2706 (N_2706,N_2498,N_2148);
nand U2707 (N_2707,N_2236,N_2095);
and U2708 (N_2708,N_2117,N_2343);
and U2709 (N_2709,N_2466,N_2358);
or U2710 (N_2710,N_2483,N_2273);
and U2711 (N_2711,N_2054,N_2470);
and U2712 (N_2712,N_2253,N_2050);
nor U2713 (N_2713,N_2437,N_2234);
xor U2714 (N_2714,N_2038,N_2478);
and U2715 (N_2715,N_2440,N_2488);
xnor U2716 (N_2716,N_2262,N_2138);
nor U2717 (N_2717,N_2348,N_2100);
nand U2718 (N_2718,N_2239,N_2423);
or U2719 (N_2719,N_2197,N_2090);
or U2720 (N_2720,N_2370,N_2384);
nand U2721 (N_2721,N_2356,N_2207);
nor U2722 (N_2722,N_2445,N_2464);
nor U2723 (N_2723,N_2023,N_2333);
nand U2724 (N_2724,N_2315,N_2266);
and U2725 (N_2725,N_2101,N_2096);
xnor U2726 (N_2726,N_2361,N_2469);
nand U2727 (N_2727,N_2329,N_2461);
nor U2728 (N_2728,N_2330,N_2270);
nand U2729 (N_2729,N_2436,N_2494);
nand U2730 (N_2730,N_2324,N_2486);
nand U2731 (N_2731,N_2163,N_2322);
xnor U2732 (N_2732,N_2441,N_2255);
and U2733 (N_2733,N_2359,N_2442);
and U2734 (N_2734,N_2136,N_2025);
or U2735 (N_2735,N_2424,N_2311);
nand U2736 (N_2736,N_2367,N_2146);
nor U2737 (N_2737,N_2291,N_2086);
nor U2738 (N_2738,N_2256,N_2250);
or U2739 (N_2739,N_2381,N_2496);
or U2740 (N_2740,N_2188,N_2036);
nand U2741 (N_2741,N_2413,N_2084);
nand U2742 (N_2742,N_2249,N_2242);
and U2743 (N_2743,N_2379,N_2487);
or U2744 (N_2744,N_2127,N_2089);
and U2745 (N_2745,N_2374,N_2183);
xnor U2746 (N_2746,N_2385,N_2346);
and U2747 (N_2747,N_2156,N_2039);
and U2748 (N_2748,N_2304,N_2237);
nor U2749 (N_2749,N_2444,N_2147);
nor U2750 (N_2750,N_2254,N_2314);
nand U2751 (N_2751,N_2363,N_2320);
and U2752 (N_2752,N_2481,N_2080);
or U2753 (N_2753,N_2448,N_2220);
nand U2754 (N_2754,N_2078,N_2310);
nor U2755 (N_2755,N_2316,N_2461);
nor U2756 (N_2756,N_2121,N_2003);
and U2757 (N_2757,N_2110,N_2374);
xor U2758 (N_2758,N_2363,N_2220);
or U2759 (N_2759,N_2293,N_2465);
nand U2760 (N_2760,N_2179,N_2123);
nand U2761 (N_2761,N_2208,N_2004);
nand U2762 (N_2762,N_2106,N_2339);
nand U2763 (N_2763,N_2429,N_2218);
nand U2764 (N_2764,N_2196,N_2447);
or U2765 (N_2765,N_2397,N_2166);
xnor U2766 (N_2766,N_2209,N_2231);
nor U2767 (N_2767,N_2248,N_2262);
and U2768 (N_2768,N_2337,N_2313);
nor U2769 (N_2769,N_2245,N_2302);
nor U2770 (N_2770,N_2221,N_2190);
or U2771 (N_2771,N_2292,N_2231);
xor U2772 (N_2772,N_2100,N_2137);
nor U2773 (N_2773,N_2031,N_2180);
and U2774 (N_2774,N_2334,N_2087);
nor U2775 (N_2775,N_2326,N_2164);
and U2776 (N_2776,N_2160,N_2439);
or U2777 (N_2777,N_2410,N_2094);
nor U2778 (N_2778,N_2210,N_2423);
or U2779 (N_2779,N_2235,N_2133);
nand U2780 (N_2780,N_2448,N_2076);
nor U2781 (N_2781,N_2335,N_2432);
nor U2782 (N_2782,N_2045,N_2105);
and U2783 (N_2783,N_2112,N_2204);
xnor U2784 (N_2784,N_2041,N_2096);
nor U2785 (N_2785,N_2103,N_2213);
xor U2786 (N_2786,N_2418,N_2262);
or U2787 (N_2787,N_2420,N_2147);
nand U2788 (N_2788,N_2044,N_2442);
nand U2789 (N_2789,N_2132,N_2480);
xnor U2790 (N_2790,N_2383,N_2332);
xor U2791 (N_2791,N_2043,N_2422);
and U2792 (N_2792,N_2408,N_2314);
and U2793 (N_2793,N_2230,N_2209);
and U2794 (N_2794,N_2421,N_2434);
and U2795 (N_2795,N_2050,N_2149);
nor U2796 (N_2796,N_2188,N_2322);
xor U2797 (N_2797,N_2245,N_2049);
and U2798 (N_2798,N_2245,N_2318);
or U2799 (N_2799,N_2128,N_2186);
nand U2800 (N_2800,N_2087,N_2144);
and U2801 (N_2801,N_2094,N_2359);
nor U2802 (N_2802,N_2294,N_2215);
nor U2803 (N_2803,N_2079,N_2199);
or U2804 (N_2804,N_2251,N_2102);
nor U2805 (N_2805,N_2259,N_2493);
and U2806 (N_2806,N_2370,N_2294);
or U2807 (N_2807,N_2440,N_2304);
xor U2808 (N_2808,N_2355,N_2441);
or U2809 (N_2809,N_2301,N_2481);
nand U2810 (N_2810,N_2188,N_2487);
xnor U2811 (N_2811,N_2318,N_2177);
xor U2812 (N_2812,N_2162,N_2439);
or U2813 (N_2813,N_2079,N_2102);
and U2814 (N_2814,N_2362,N_2424);
nand U2815 (N_2815,N_2199,N_2045);
or U2816 (N_2816,N_2350,N_2025);
and U2817 (N_2817,N_2079,N_2379);
xor U2818 (N_2818,N_2416,N_2431);
and U2819 (N_2819,N_2497,N_2419);
nor U2820 (N_2820,N_2054,N_2368);
nor U2821 (N_2821,N_2456,N_2321);
nor U2822 (N_2822,N_2297,N_2070);
nor U2823 (N_2823,N_2414,N_2228);
and U2824 (N_2824,N_2450,N_2499);
or U2825 (N_2825,N_2245,N_2084);
xor U2826 (N_2826,N_2450,N_2318);
nor U2827 (N_2827,N_2096,N_2418);
and U2828 (N_2828,N_2296,N_2313);
and U2829 (N_2829,N_2394,N_2413);
nor U2830 (N_2830,N_2281,N_2042);
or U2831 (N_2831,N_2330,N_2006);
or U2832 (N_2832,N_2321,N_2043);
or U2833 (N_2833,N_2151,N_2330);
or U2834 (N_2834,N_2119,N_2023);
nand U2835 (N_2835,N_2168,N_2467);
nand U2836 (N_2836,N_2243,N_2395);
and U2837 (N_2837,N_2236,N_2385);
xor U2838 (N_2838,N_2011,N_2271);
nand U2839 (N_2839,N_2481,N_2430);
nor U2840 (N_2840,N_2073,N_2452);
or U2841 (N_2841,N_2198,N_2227);
or U2842 (N_2842,N_2157,N_2035);
nor U2843 (N_2843,N_2130,N_2180);
nor U2844 (N_2844,N_2037,N_2478);
nor U2845 (N_2845,N_2467,N_2159);
nand U2846 (N_2846,N_2093,N_2235);
xnor U2847 (N_2847,N_2145,N_2191);
xor U2848 (N_2848,N_2203,N_2426);
nand U2849 (N_2849,N_2374,N_2179);
xnor U2850 (N_2850,N_2274,N_2423);
and U2851 (N_2851,N_2431,N_2035);
xor U2852 (N_2852,N_2329,N_2125);
or U2853 (N_2853,N_2161,N_2084);
or U2854 (N_2854,N_2276,N_2010);
xor U2855 (N_2855,N_2077,N_2093);
nand U2856 (N_2856,N_2228,N_2257);
and U2857 (N_2857,N_2309,N_2203);
nor U2858 (N_2858,N_2415,N_2327);
nor U2859 (N_2859,N_2151,N_2186);
nand U2860 (N_2860,N_2436,N_2185);
nand U2861 (N_2861,N_2379,N_2070);
nand U2862 (N_2862,N_2460,N_2011);
nor U2863 (N_2863,N_2024,N_2475);
nand U2864 (N_2864,N_2297,N_2499);
or U2865 (N_2865,N_2407,N_2245);
nor U2866 (N_2866,N_2372,N_2145);
nand U2867 (N_2867,N_2477,N_2175);
xor U2868 (N_2868,N_2206,N_2338);
nor U2869 (N_2869,N_2332,N_2438);
xnor U2870 (N_2870,N_2292,N_2242);
nand U2871 (N_2871,N_2365,N_2256);
nand U2872 (N_2872,N_2253,N_2178);
or U2873 (N_2873,N_2117,N_2288);
or U2874 (N_2874,N_2239,N_2014);
nor U2875 (N_2875,N_2216,N_2454);
xnor U2876 (N_2876,N_2072,N_2497);
and U2877 (N_2877,N_2099,N_2316);
xnor U2878 (N_2878,N_2341,N_2151);
xor U2879 (N_2879,N_2419,N_2397);
nor U2880 (N_2880,N_2150,N_2081);
xor U2881 (N_2881,N_2464,N_2259);
or U2882 (N_2882,N_2248,N_2049);
xor U2883 (N_2883,N_2308,N_2232);
xor U2884 (N_2884,N_2069,N_2363);
or U2885 (N_2885,N_2490,N_2312);
nand U2886 (N_2886,N_2299,N_2207);
or U2887 (N_2887,N_2411,N_2268);
nand U2888 (N_2888,N_2101,N_2286);
xor U2889 (N_2889,N_2260,N_2061);
and U2890 (N_2890,N_2215,N_2323);
xor U2891 (N_2891,N_2278,N_2265);
nand U2892 (N_2892,N_2226,N_2216);
nor U2893 (N_2893,N_2415,N_2412);
or U2894 (N_2894,N_2086,N_2295);
nand U2895 (N_2895,N_2061,N_2187);
nor U2896 (N_2896,N_2110,N_2416);
xnor U2897 (N_2897,N_2288,N_2448);
nand U2898 (N_2898,N_2433,N_2333);
or U2899 (N_2899,N_2166,N_2035);
xnor U2900 (N_2900,N_2342,N_2333);
xor U2901 (N_2901,N_2034,N_2006);
nand U2902 (N_2902,N_2039,N_2302);
xor U2903 (N_2903,N_2343,N_2036);
xnor U2904 (N_2904,N_2248,N_2428);
nor U2905 (N_2905,N_2214,N_2185);
or U2906 (N_2906,N_2311,N_2131);
or U2907 (N_2907,N_2015,N_2342);
xnor U2908 (N_2908,N_2413,N_2026);
and U2909 (N_2909,N_2454,N_2358);
nor U2910 (N_2910,N_2023,N_2007);
nand U2911 (N_2911,N_2431,N_2174);
or U2912 (N_2912,N_2301,N_2432);
or U2913 (N_2913,N_2456,N_2329);
or U2914 (N_2914,N_2122,N_2267);
nand U2915 (N_2915,N_2180,N_2476);
nor U2916 (N_2916,N_2141,N_2201);
nor U2917 (N_2917,N_2186,N_2099);
nor U2918 (N_2918,N_2366,N_2254);
xor U2919 (N_2919,N_2079,N_2089);
and U2920 (N_2920,N_2421,N_2348);
xor U2921 (N_2921,N_2024,N_2172);
nand U2922 (N_2922,N_2189,N_2314);
xnor U2923 (N_2923,N_2048,N_2333);
and U2924 (N_2924,N_2057,N_2341);
or U2925 (N_2925,N_2196,N_2261);
and U2926 (N_2926,N_2061,N_2108);
xnor U2927 (N_2927,N_2464,N_2307);
xor U2928 (N_2928,N_2463,N_2213);
or U2929 (N_2929,N_2221,N_2222);
xnor U2930 (N_2930,N_2439,N_2292);
and U2931 (N_2931,N_2181,N_2171);
or U2932 (N_2932,N_2399,N_2439);
and U2933 (N_2933,N_2054,N_2327);
nor U2934 (N_2934,N_2350,N_2129);
nor U2935 (N_2935,N_2417,N_2202);
and U2936 (N_2936,N_2181,N_2439);
or U2937 (N_2937,N_2315,N_2139);
and U2938 (N_2938,N_2296,N_2125);
nor U2939 (N_2939,N_2100,N_2426);
or U2940 (N_2940,N_2237,N_2042);
or U2941 (N_2941,N_2397,N_2201);
or U2942 (N_2942,N_2163,N_2111);
and U2943 (N_2943,N_2090,N_2394);
or U2944 (N_2944,N_2246,N_2390);
nand U2945 (N_2945,N_2478,N_2335);
and U2946 (N_2946,N_2057,N_2324);
or U2947 (N_2947,N_2132,N_2292);
or U2948 (N_2948,N_2200,N_2016);
nor U2949 (N_2949,N_2407,N_2472);
nand U2950 (N_2950,N_2088,N_2335);
nor U2951 (N_2951,N_2168,N_2226);
nand U2952 (N_2952,N_2150,N_2191);
xor U2953 (N_2953,N_2288,N_2091);
xor U2954 (N_2954,N_2468,N_2248);
nor U2955 (N_2955,N_2164,N_2067);
or U2956 (N_2956,N_2416,N_2290);
and U2957 (N_2957,N_2173,N_2314);
nor U2958 (N_2958,N_2150,N_2303);
nand U2959 (N_2959,N_2474,N_2390);
nor U2960 (N_2960,N_2124,N_2041);
nor U2961 (N_2961,N_2227,N_2066);
nand U2962 (N_2962,N_2321,N_2151);
nand U2963 (N_2963,N_2089,N_2031);
nand U2964 (N_2964,N_2427,N_2404);
or U2965 (N_2965,N_2338,N_2186);
and U2966 (N_2966,N_2489,N_2247);
xor U2967 (N_2967,N_2131,N_2492);
xnor U2968 (N_2968,N_2277,N_2266);
nor U2969 (N_2969,N_2106,N_2018);
and U2970 (N_2970,N_2350,N_2234);
or U2971 (N_2971,N_2452,N_2470);
xor U2972 (N_2972,N_2138,N_2113);
and U2973 (N_2973,N_2241,N_2139);
nand U2974 (N_2974,N_2442,N_2357);
nor U2975 (N_2975,N_2268,N_2277);
nor U2976 (N_2976,N_2217,N_2245);
nand U2977 (N_2977,N_2366,N_2227);
xor U2978 (N_2978,N_2076,N_2424);
or U2979 (N_2979,N_2303,N_2075);
nor U2980 (N_2980,N_2260,N_2399);
xor U2981 (N_2981,N_2442,N_2274);
or U2982 (N_2982,N_2418,N_2008);
nor U2983 (N_2983,N_2457,N_2232);
nor U2984 (N_2984,N_2415,N_2265);
nor U2985 (N_2985,N_2341,N_2326);
xor U2986 (N_2986,N_2238,N_2338);
or U2987 (N_2987,N_2425,N_2313);
nor U2988 (N_2988,N_2053,N_2126);
nor U2989 (N_2989,N_2422,N_2270);
nand U2990 (N_2990,N_2266,N_2481);
nand U2991 (N_2991,N_2162,N_2142);
nor U2992 (N_2992,N_2257,N_2256);
xor U2993 (N_2993,N_2338,N_2283);
nand U2994 (N_2994,N_2083,N_2133);
xnor U2995 (N_2995,N_2383,N_2409);
nor U2996 (N_2996,N_2430,N_2373);
nand U2997 (N_2997,N_2290,N_2371);
nor U2998 (N_2998,N_2486,N_2414);
and U2999 (N_2999,N_2022,N_2252);
or U3000 (N_3000,N_2647,N_2967);
xnor U3001 (N_3001,N_2636,N_2630);
nand U3002 (N_3002,N_2528,N_2873);
and U3003 (N_3003,N_2853,N_2608);
or U3004 (N_3004,N_2567,N_2592);
nor U3005 (N_3005,N_2750,N_2622);
xor U3006 (N_3006,N_2736,N_2947);
nand U3007 (N_3007,N_2661,N_2614);
xnor U3008 (N_3008,N_2638,N_2707);
or U3009 (N_3009,N_2639,N_2844);
and U3010 (N_3010,N_2949,N_2932);
nor U3011 (N_3011,N_2723,N_2913);
or U3012 (N_3012,N_2655,N_2749);
nor U3013 (N_3013,N_2910,N_2602);
or U3014 (N_3014,N_2806,N_2951);
and U3015 (N_3015,N_2888,N_2535);
xnor U3016 (N_3016,N_2775,N_2727);
or U3017 (N_3017,N_2869,N_2817);
nor U3018 (N_3018,N_2526,N_2722);
or U3019 (N_3019,N_2942,N_2937);
nor U3020 (N_3020,N_2955,N_2768);
or U3021 (N_3021,N_2551,N_2934);
nand U3022 (N_3022,N_2856,N_2771);
nand U3023 (N_3023,N_2677,N_2863);
nor U3024 (N_3024,N_2599,N_2816);
nor U3025 (N_3025,N_2812,N_2555);
nand U3026 (N_3026,N_2995,N_2593);
xnor U3027 (N_3027,N_2524,N_2579);
and U3028 (N_3028,N_2890,N_2763);
nor U3029 (N_3029,N_2719,N_2505);
and U3030 (N_3030,N_2893,N_2559);
and U3031 (N_3031,N_2785,N_2633);
xor U3032 (N_3032,N_2927,N_2804);
or U3033 (N_3033,N_2635,N_2987);
or U3034 (N_3034,N_2936,N_2918);
xor U3035 (N_3035,N_2646,N_2714);
or U3036 (N_3036,N_2504,N_2781);
nand U3037 (N_3037,N_2566,N_2859);
nand U3038 (N_3038,N_2813,N_2626);
xnor U3039 (N_3039,N_2867,N_2653);
xnor U3040 (N_3040,N_2693,N_2849);
nand U3041 (N_3041,N_2583,N_2997);
or U3042 (N_3042,N_2931,N_2684);
or U3043 (N_3043,N_2857,N_2687);
xnor U3044 (N_3044,N_2905,N_2974);
nand U3045 (N_3045,N_2836,N_2916);
nor U3046 (N_3046,N_2810,N_2782);
xor U3047 (N_3047,N_2939,N_2897);
and U3048 (N_3048,N_2858,N_2521);
nor U3049 (N_3049,N_2909,N_2900);
and U3050 (N_3050,N_2685,N_2514);
nand U3051 (N_3051,N_2770,N_2944);
or U3052 (N_3052,N_2801,N_2848);
or U3053 (N_3053,N_2582,N_2531);
xor U3054 (N_3054,N_2837,N_2780);
nand U3055 (N_3055,N_2713,N_2985);
nor U3056 (N_3056,N_2720,N_2898);
and U3057 (N_3057,N_2965,N_2778);
nand U3058 (N_3058,N_2652,N_2969);
or U3059 (N_3059,N_2598,N_2620);
or U3060 (N_3060,N_2532,N_2701);
nor U3061 (N_3061,N_2676,N_2520);
or U3062 (N_3062,N_2922,N_2980);
and U3063 (N_3063,N_2843,N_2797);
or U3064 (N_3064,N_2966,N_2889);
nand U3065 (N_3065,N_2891,N_2503);
nor U3066 (N_3066,N_2549,N_2870);
xnor U3067 (N_3067,N_2590,N_2809);
and U3068 (N_3068,N_2610,N_2774);
nand U3069 (N_3069,N_2794,N_2989);
and U3070 (N_3070,N_2656,N_2654);
nor U3071 (N_3071,N_2699,N_2712);
nor U3072 (N_3072,N_2850,N_2698);
and U3073 (N_3073,N_2577,N_2605);
xor U3074 (N_3074,N_2865,N_2525);
and U3075 (N_3075,N_2904,N_2546);
xor U3076 (N_3076,N_2686,N_2740);
xor U3077 (N_3077,N_2758,N_2747);
xor U3078 (N_3078,N_2772,N_2507);
xor U3079 (N_3079,N_2615,N_2923);
nand U3080 (N_3080,N_2788,N_2991);
and U3081 (N_3081,N_2711,N_2820);
nand U3082 (N_3082,N_2764,N_2935);
nand U3083 (N_3083,N_2954,N_2612);
nor U3084 (N_3084,N_2883,N_2641);
and U3085 (N_3085,N_2721,N_2545);
and U3086 (N_3086,N_2829,N_2956);
or U3087 (N_3087,N_2501,N_2790);
xor U3088 (N_3088,N_2570,N_2755);
xnor U3089 (N_3089,N_2650,N_2887);
or U3090 (N_3090,N_2841,N_2563);
or U3091 (N_3091,N_2730,N_2851);
nor U3092 (N_3092,N_2729,N_2990);
and U3093 (N_3093,N_2793,N_2564);
nor U3094 (N_3094,N_2901,N_2648);
and U3095 (N_3095,N_2695,N_2678);
nor U3096 (N_3096,N_2600,N_2732);
nand U3097 (N_3097,N_2899,N_2971);
nand U3098 (N_3098,N_2575,N_2968);
nand U3099 (N_3099,N_2613,N_2716);
nand U3100 (N_3100,N_2784,N_2536);
nand U3101 (N_3101,N_2674,N_2673);
nor U3102 (N_3102,N_2643,N_2538);
and U3103 (N_3103,N_2999,N_2717);
nor U3104 (N_3104,N_2511,N_2627);
nor U3105 (N_3105,N_2534,N_2731);
nand U3106 (N_3106,N_2562,N_2880);
nor U3107 (N_3107,N_2948,N_2765);
and U3108 (N_3108,N_2573,N_2862);
xnor U3109 (N_3109,N_2961,N_2920);
and U3110 (N_3110,N_2928,N_2798);
xnor U3111 (N_3111,N_2941,N_2726);
nor U3112 (N_3112,N_2751,N_2914);
nor U3113 (N_3113,N_2973,N_2854);
nor U3114 (N_3114,N_2527,N_2984);
xor U3115 (N_3115,N_2586,N_2940);
and U3116 (N_3116,N_2666,N_2894);
xor U3117 (N_3117,N_2537,N_2581);
or U3118 (N_3118,N_2609,N_2960);
or U3119 (N_3119,N_2933,N_2675);
or U3120 (N_3120,N_2539,N_2815);
and U3121 (N_3121,N_2972,N_2706);
and U3122 (N_3122,N_2547,N_2607);
nor U3123 (N_3123,N_2983,N_2710);
xor U3124 (N_3124,N_2540,N_2616);
nand U3125 (N_3125,N_2629,N_2659);
xnor U3126 (N_3126,N_2981,N_2557);
and U3127 (N_3127,N_2625,N_2632);
nor U3128 (N_3128,N_2805,N_2508);
nor U3129 (N_3129,N_2776,N_2550);
nor U3130 (N_3130,N_2752,N_2822);
and U3131 (N_3131,N_2779,N_2753);
nand U3132 (N_3132,N_2825,N_2881);
and U3133 (N_3133,N_2572,N_2522);
xnor U3134 (N_3134,N_2634,N_2548);
nand U3135 (N_3135,N_2876,N_2975);
or U3136 (N_3136,N_2672,N_2819);
or U3137 (N_3137,N_2544,N_2606);
xor U3138 (N_3138,N_2631,N_2560);
nor U3139 (N_3139,N_2943,N_2530);
and U3140 (N_3140,N_2908,N_2715);
xnor U3141 (N_3141,N_2733,N_2574);
and U3142 (N_3142,N_2906,N_2515);
nor U3143 (N_3143,N_2831,N_2748);
and U3144 (N_3144,N_2946,N_2868);
or U3145 (N_3145,N_2957,N_2872);
and U3146 (N_3146,N_2847,N_2818);
and U3147 (N_3147,N_2604,N_2619);
and U3148 (N_3148,N_2926,N_2651);
and U3149 (N_3149,N_2879,N_2533);
xnor U3150 (N_3150,N_2742,N_2724);
nand U3151 (N_3151,N_2644,N_2689);
nor U3152 (N_3152,N_2786,N_2864);
nand U3153 (N_3153,N_2512,N_2777);
nand U3154 (N_3154,N_2958,N_2688);
xor U3155 (N_3155,N_2554,N_2866);
nand U3156 (N_3156,N_2696,N_2628);
nor U3157 (N_3157,N_2697,N_2725);
nand U3158 (N_3158,N_2911,N_2561);
nor U3159 (N_3159,N_2553,N_2704);
xor U3160 (N_3160,N_2840,N_2787);
nor U3161 (N_3161,N_2657,N_2878);
and U3162 (N_3162,N_2513,N_2611);
and U3163 (N_3163,N_2875,N_2976);
or U3164 (N_3164,N_2921,N_2962);
xor U3165 (N_3165,N_2552,N_2664);
xor U3166 (N_3166,N_2744,N_2993);
or U3167 (N_3167,N_2930,N_2811);
and U3168 (N_3168,N_2800,N_2737);
xnor U3169 (N_3169,N_2500,N_2978);
xnor U3170 (N_3170,N_2681,N_2986);
xnor U3171 (N_3171,N_2588,N_2692);
and U3172 (N_3172,N_2743,N_2649);
xor U3173 (N_3173,N_2658,N_2877);
or U3174 (N_3174,N_2585,N_2821);
xnor U3175 (N_3175,N_2739,N_2846);
nand U3176 (N_3176,N_2506,N_2591);
nor U3177 (N_3177,N_2871,N_2708);
nand U3178 (N_3178,N_2669,N_2959);
xor U3179 (N_3179,N_2754,N_2834);
nand U3180 (N_3180,N_2694,N_2827);
xor U3181 (N_3181,N_2766,N_2642);
xor U3182 (N_3182,N_2667,N_2728);
nor U3183 (N_3183,N_2556,N_2663);
and U3184 (N_3184,N_2569,N_2830);
xnor U3185 (N_3185,N_2919,N_2882);
nor U3186 (N_3186,N_2580,N_2759);
or U3187 (N_3187,N_2529,N_2587);
nand U3188 (N_3188,N_2568,N_2795);
nor U3189 (N_3189,N_2640,N_2799);
and U3190 (N_3190,N_2892,N_2839);
nand U3191 (N_3191,N_2623,N_2571);
nor U3192 (N_3192,N_2601,N_2789);
xnor U3193 (N_3193,N_2769,N_2895);
nand U3194 (N_3194,N_2746,N_2907);
and U3195 (N_3195,N_2828,N_2679);
nor U3196 (N_3196,N_2807,N_2925);
nor U3197 (N_3197,N_2584,N_2802);
or U3198 (N_3198,N_2665,N_2705);
or U3199 (N_3199,N_2796,N_2523);
nand U3200 (N_3200,N_2808,N_2924);
nor U3201 (N_3201,N_2950,N_2860);
xnor U3202 (N_3202,N_2690,N_2668);
nor U3203 (N_3203,N_2516,N_2833);
nand U3204 (N_3204,N_2745,N_2576);
nor U3205 (N_3205,N_2541,N_2783);
nor U3206 (N_3206,N_2502,N_2542);
and U3207 (N_3207,N_2845,N_2578);
xor U3208 (N_3208,N_2979,N_2671);
nor U3209 (N_3209,N_2660,N_2594);
nand U3210 (N_3210,N_2886,N_2756);
xor U3211 (N_3211,N_2682,N_2734);
nor U3212 (N_3212,N_2992,N_2518);
nor U3213 (N_3213,N_2741,N_2703);
xor U3214 (N_3214,N_2597,N_2824);
nand U3215 (N_3215,N_2510,N_2953);
nor U3216 (N_3216,N_2803,N_2996);
or U3217 (N_3217,N_2823,N_2977);
nand U3218 (N_3218,N_2683,N_2761);
and U3219 (N_3219,N_2994,N_2709);
nand U3220 (N_3220,N_2637,N_2963);
and U3221 (N_3221,N_2964,N_2838);
and U3222 (N_3222,N_2791,N_2517);
and U3223 (N_3223,N_2998,N_2814);
nor U3224 (N_3224,N_2903,N_2670);
nand U3225 (N_3225,N_2595,N_2915);
nor U3226 (N_3226,N_2874,N_2662);
or U3227 (N_3227,N_2762,N_2896);
nor U3228 (N_3228,N_2912,N_2735);
nor U3229 (N_3229,N_2760,N_2589);
nor U3230 (N_3230,N_2603,N_2596);
or U3231 (N_3231,N_2982,N_2970);
nor U3232 (N_3232,N_2884,N_2509);
nor U3233 (N_3233,N_2618,N_2757);
nor U3234 (N_3234,N_2773,N_2543);
nor U3235 (N_3235,N_2861,N_2938);
nand U3236 (N_3236,N_2702,N_2621);
nand U3237 (N_3237,N_2988,N_2700);
nand U3238 (N_3238,N_2691,N_2945);
nor U3239 (N_3239,N_2855,N_2832);
nand U3240 (N_3240,N_2718,N_2738);
or U3241 (N_3241,N_2519,N_2792);
xor U3242 (N_3242,N_2680,N_2835);
nor U3243 (N_3243,N_2826,N_2902);
and U3244 (N_3244,N_2565,N_2645);
nand U3245 (N_3245,N_2558,N_2917);
nor U3246 (N_3246,N_2852,N_2624);
or U3247 (N_3247,N_2767,N_2929);
or U3248 (N_3248,N_2842,N_2617);
and U3249 (N_3249,N_2885,N_2952);
and U3250 (N_3250,N_2973,N_2808);
nor U3251 (N_3251,N_2561,N_2883);
and U3252 (N_3252,N_2818,N_2548);
or U3253 (N_3253,N_2969,N_2857);
xnor U3254 (N_3254,N_2971,N_2880);
or U3255 (N_3255,N_2725,N_2934);
nand U3256 (N_3256,N_2658,N_2908);
and U3257 (N_3257,N_2603,N_2999);
xnor U3258 (N_3258,N_2750,N_2857);
nor U3259 (N_3259,N_2695,N_2791);
nand U3260 (N_3260,N_2608,N_2950);
xnor U3261 (N_3261,N_2957,N_2793);
nand U3262 (N_3262,N_2538,N_2617);
nand U3263 (N_3263,N_2740,N_2729);
and U3264 (N_3264,N_2962,N_2775);
nor U3265 (N_3265,N_2825,N_2529);
nor U3266 (N_3266,N_2862,N_2605);
and U3267 (N_3267,N_2639,N_2942);
and U3268 (N_3268,N_2510,N_2773);
and U3269 (N_3269,N_2983,N_2898);
nor U3270 (N_3270,N_2786,N_2905);
or U3271 (N_3271,N_2952,N_2534);
nand U3272 (N_3272,N_2614,N_2755);
nor U3273 (N_3273,N_2916,N_2576);
nor U3274 (N_3274,N_2952,N_2964);
nand U3275 (N_3275,N_2503,N_2589);
nor U3276 (N_3276,N_2946,N_2890);
or U3277 (N_3277,N_2813,N_2955);
or U3278 (N_3278,N_2677,N_2983);
and U3279 (N_3279,N_2874,N_2716);
xnor U3280 (N_3280,N_2719,N_2993);
or U3281 (N_3281,N_2948,N_2764);
and U3282 (N_3282,N_2697,N_2729);
or U3283 (N_3283,N_2531,N_2538);
nor U3284 (N_3284,N_2593,N_2765);
nor U3285 (N_3285,N_2743,N_2877);
or U3286 (N_3286,N_2749,N_2614);
or U3287 (N_3287,N_2854,N_2752);
nor U3288 (N_3288,N_2656,N_2760);
xor U3289 (N_3289,N_2715,N_2628);
nor U3290 (N_3290,N_2509,N_2807);
and U3291 (N_3291,N_2819,N_2994);
nor U3292 (N_3292,N_2664,N_2642);
nand U3293 (N_3293,N_2797,N_2689);
and U3294 (N_3294,N_2788,N_2838);
nor U3295 (N_3295,N_2677,N_2521);
nor U3296 (N_3296,N_2891,N_2589);
or U3297 (N_3297,N_2920,N_2849);
xor U3298 (N_3298,N_2579,N_2822);
nor U3299 (N_3299,N_2732,N_2656);
and U3300 (N_3300,N_2798,N_2819);
nor U3301 (N_3301,N_2585,N_2865);
nand U3302 (N_3302,N_2909,N_2823);
xnor U3303 (N_3303,N_2849,N_2814);
nor U3304 (N_3304,N_2964,N_2953);
nand U3305 (N_3305,N_2899,N_2644);
and U3306 (N_3306,N_2640,N_2838);
nand U3307 (N_3307,N_2603,N_2554);
nand U3308 (N_3308,N_2818,N_2892);
nand U3309 (N_3309,N_2579,N_2936);
nand U3310 (N_3310,N_2737,N_2870);
and U3311 (N_3311,N_2831,N_2755);
nand U3312 (N_3312,N_2528,N_2771);
nor U3313 (N_3313,N_2640,N_2982);
xor U3314 (N_3314,N_2899,N_2882);
and U3315 (N_3315,N_2736,N_2968);
or U3316 (N_3316,N_2686,N_2671);
or U3317 (N_3317,N_2880,N_2678);
or U3318 (N_3318,N_2684,N_2923);
nand U3319 (N_3319,N_2507,N_2646);
nand U3320 (N_3320,N_2587,N_2570);
nand U3321 (N_3321,N_2984,N_2797);
nor U3322 (N_3322,N_2788,N_2721);
or U3323 (N_3323,N_2731,N_2559);
xnor U3324 (N_3324,N_2807,N_2557);
or U3325 (N_3325,N_2792,N_2622);
or U3326 (N_3326,N_2854,N_2858);
nor U3327 (N_3327,N_2565,N_2843);
xor U3328 (N_3328,N_2682,N_2748);
nand U3329 (N_3329,N_2711,N_2732);
nor U3330 (N_3330,N_2562,N_2728);
and U3331 (N_3331,N_2918,N_2566);
and U3332 (N_3332,N_2662,N_2579);
or U3333 (N_3333,N_2749,N_2914);
xnor U3334 (N_3334,N_2929,N_2728);
or U3335 (N_3335,N_2881,N_2982);
and U3336 (N_3336,N_2961,N_2824);
and U3337 (N_3337,N_2643,N_2562);
xnor U3338 (N_3338,N_2744,N_2506);
xnor U3339 (N_3339,N_2920,N_2535);
or U3340 (N_3340,N_2948,N_2711);
nor U3341 (N_3341,N_2517,N_2799);
nor U3342 (N_3342,N_2563,N_2827);
nand U3343 (N_3343,N_2903,N_2883);
or U3344 (N_3344,N_2818,N_2596);
and U3345 (N_3345,N_2918,N_2891);
xnor U3346 (N_3346,N_2852,N_2973);
xnor U3347 (N_3347,N_2735,N_2725);
nand U3348 (N_3348,N_2880,N_2900);
nor U3349 (N_3349,N_2629,N_2671);
nand U3350 (N_3350,N_2976,N_2591);
nand U3351 (N_3351,N_2774,N_2606);
or U3352 (N_3352,N_2798,N_2616);
nor U3353 (N_3353,N_2772,N_2920);
nor U3354 (N_3354,N_2906,N_2798);
and U3355 (N_3355,N_2793,N_2613);
or U3356 (N_3356,N_2986,N_2946);
and U3357 (N_3357,N_2704,N_2601);
or U3358 (N_3358,N_2755,N_2886);
or U3359 (N_3359,N_2746,N_2902);
nor U3360 (N_3360,N_2512,N_2894);
xnor U3361 (N_3361,N_2805,N_2930);
or U3362 (N_3362,N_2624,N_2887);
nor U3363 (N_3363,N_2850,N_2970);
or U3364 (N_3364,N_2790,N_2613);
nand U3365 (N_3365,N_2891,N_2701);
nand U3366 (N_3366,N_2867,N_2755);
and U3367 (N_3367,N_2545,N_2603);
nor U3368 (N_3368,N_2648,N_2873);
xor U3369 (N_3369,N_2673,N_2854);
or U3370 (N_3370,N_2989,N_2637);
or U3371 (N_3371,N_2729,N_2826);
nor U3372 (N_3372,N_2880,N_2508);
xnor U3373 (N_3373,N_2683,N_2919);
or U3374 (N_3374,N_2874,N_2864);
nand U3375 (N_3375,N_2871,N_2792);
xnor U3376 (N_3376,N_2636,N_2957);
or U3377 (N_3377,N_2755,N_2980);
or U3378 (N_3378,N_2799,N_2591);
nor U3379 (N_3379,N_2716,N_2777);
xor U3380 (N_3380,N_2933,N_2618);
nor U3381 (N_3381,N_2614,N_2919);
and U3382 (N_3382,N_2659,N_2570);
xor U3383 (N_3383,N_2854,N_2543);
nor U3384 (N_3384,N_2729,N_2584);
xnor U3385 (N_3385,N_2846,N_2997);
nand U3386 (N_3386,N_2768,N_2988);
nand U3387 (N_3387,N_2574,N_2515);
and U3388 (N_3388,N_2893,N_2909);
nor U3389 (N_3389,N_2564,N_2969);
nor U3390 (N_3390,N_2878,N_2949);
nand U3391 (N_3391,N_2626,N_2791);
or U3392 (N_3392,N_2784,N_2968);
nor U3393 (N_3393,N_2713,N_2677);
nor U3394 (N_3394,N_2873,N_2590);
or U3395 (N_3395,N_2579,N_2829);
or U3396 (N_3396,N_2656,N_2720);
nand U3397 (N_3397,N_2577,N_2632);
xnor U3398 (N_3398,N_2711,N_2527);
nor U3399 (N_3399,N_2876,N_2756);
and U3400 (N_3400,N_2846,N_2683);
xor U3401 (N_3401,N_2569,N_2782);
nand U3402 (N_3402,N_2676,N_2851);
xor U3403 (N_3403,N_2723,N_2542);
xor U3404 (N_3404,N_2923,N_2599);
nand U3405 (N_3405,N_2946,N_2981);
or U3406 (N_3406,N_2767,N_2643);
or U3407 (N_3407,N_2771,N_2596);
nor U3408 (N_3408,N_2871,N_2910);
xor U3409 (N_3409,N_2649,N_2733);
xnor U3410 (N_3410,N_2633,N_2922);
and U3411 (N_3411,N_2522,N_2580);
xor U3412 (N_3412,N_2816,N_2956);
nand U3413 (N_3413,N_2553,N_2807);
nand U3414 (N_3414,N_2885,N_2630);
or U3415 (N_3415,N_2578,N_2791);
or U3416 (N_3416,N_2752,N_2797);
or U3417 (N_3417,N_2782,N_2797);
and U3418 (N_3418,N_2788,N_2500);
and U3419 (N_3419,N_2612,N_2832);
xnor U3420 (N_3420,N_2761,N_2865);
and U3421 (N_3421,N_2937,N_2731);
xor U3422 (N_3422,N_2728,N_2776);
and U3423 (N_3423,N_2717,N_2586);
xor U3424 (N_3424,N_2518,N_2794);
and U3425 (N_3425,N_2745,N_2660);
nor U3426 (N_3426,N_2973,N_2788);
nand U3427 (N_3427,N_2953,N_2569);
nor U3428 (N_3428,N_2580,N_2838);
xnor U3429 (N_3429,N_2789,N_2827);
nor U3430 (N_3430,N_2950,N_2789);
or U3431 (N_3431,N_2983,N_2784);
nor U3432 (N_3432,N_2986,N_2753);
nand U3433 (N_3433,N_2792,N_2655);
or U3434 (N_3434,N_2697,N_2632);
nand U3435 (N_3435,N_2652,N_2755);
xor U3436 (N_3436,N_2705,N_2633);
or U3437 (N_3437,N_2682,N_2576);
xnor U3438 (N_3438,N_2893,N_2892);
or U3439 (N_3439,N_2702,N_2568);
nor U3440 (N_3440,N_2533,N_2891);
and U3441 (N_3441,N_2690,N_2731);
nand U3442 (N_3442,N_2597,N_2634);
or U3443 (N_3443,N_2653,N_2663);
xor U3444 (N_3444,N_2927,N_2558);
nand U3445 (N_3445,N_2747,N_2589);
and U3446 (N_3446,N_2768,N_2803);
or U3447 (N_3447,N_2783,N_2649);
nor U3448 (N_3448,N_2865,N_2874);
and U3449 (N_3449,N_2780,N_2590);
xor U3450 (N_3450,N_2620,N_2953);
nor U3451 (N_3451,N_2587,N_2989);
xnor U3452 (N_3452,N_2808,N_2615);
nand U3453 (N_3453,N_2610,N_2575);
nand U3454 (N_3454,N_2536,N_2631);
xor U3455 (N_3455,N_2903,N_2860);
xor U3456 (N_3456,N_2962,N_2920);
xnor U3457 (N_3457,N_2668,N_2703);
nand U3458 (N_3458,N_2584,N_2597);
nand U3459 (N_3459,N_2695,N_2709);
and U3460 (N_3460,N_2627,N_2795);
nand U3461 (N_3461,N_2980,N_2649);
and U3462 (N_3462,N_2591,N_2755);
xnor U3463 (N_3463,N_2986,N_2912);
or U3464 (N_3464,N_2879,N_2545);
xnor U3465 (N_3465,N_2609,N_2510);
or U3466 (N_3466,N_2788,N_2649);
nand U3467 (N_3467,N_2542,N_2642);
nand U3468 (N_3468,N_2663,N_2922);
nand U3469 (N_3469,N_2652,N_2597);
nand U3470 (N_3470,N_2776,N_2789);
xnor U3471 (N_3471,N_2537,N_2885);
nor U3472 (N_3472,N_2883,N_2857);
xor U3473 (N_3473,N_2715,N_2708);
and U3474 (N_3474,N_2847,N_2789);
and U3475 (N_3475,N_2642,N_2909);
xnor U3476 (N_3476,N_2935,N_2771);
and U3477 (N_3477,N_2747,N_2708);
nand U3478 (N_3478,N_2623,N_2638);
or U3479 (N_3479,N_2621,N_2794);
or U3480 (N_3480,N_2647,N_2842);
nand U3481 (N_3481,N_2921,N_2873);
nand U3482 (N_3482,N_2861,N_2541);
and U3483 (N_3483,N_2543,N_2756);
and U3484 (N_3484,N_2824,N_2748);
and U3485 (N_3485,N_2870,N_2585);
nand U3486 (N_3486,N_2530,N_2665);
nor U3487 (N_3487,N_2602,N_2874);
and U3488 (N_3488,N_2752,N_2883);
nor U3489 (N_3489,N_2951,N_2727);
xnor U3490 (N_3490,N_2963,N_2898);
nor U3491 (N_3491,N_2930,N_2822);
or U3492 (N_3492,N_2596,N_2665);
xnor U3493 (N_3493,N_2502,N_2653);
or U3494 (N_3494,N_2650,N_2604);
nor U3495 (N_3495,N_2608,N_2626);
nor U3496 (N_3496,N_2924,N_2583);
xnor U3497 (N_3497,N_2913,N_2989);
or U3498 (N_3498,N_2714,N_2657);
xnor U3499 (N_3499,N_2521,N_2939);
nor U3500 (N_3500,N_3399,N_3300);
and U3501 (N_3501,N_3303,N_3231);
xnor U3502 (N_3502,N_3316,N_3113);
or U3503 (N_3503,N_3497,N_3205);
nor U3504 (N_3504,N_3382,N_3446);
xor U3505 (N_3505,N_3293,N_3371);
xor U3506 (N_3506,N_3027,N_3030);
nor U3507 (N_3507,N_3328,N_3122);
nor U3508 (N_3508,N_3039,N_3199);
and U3509 (N_3509,N_3173,N_3290);
nor U3510 (N_3510,N_3387,N_3332);
xor U3511 (N_3511,N_3344,N_3133);
nand U3512 (N_3512,N_3313,N_3451);
nand U3513 (N_3513,N_3288,N_3402);
xnor U3514 (N_3514,N_3032,N_3120);
xor U3515 (N_3515,N_3262,N_3241);
nor U3516 (N_3516,N_3442,N_3363);
xnor U3517 (N_3517,N_3105,N_3216);
nor U3518 (N_3518,N_3406,N_3237);
or U3519 (N_3519,N_3349,N_3396);
and U3520 (N_3520,N_3153,N_3114);
and U3521 (N_3521,N_3395,N_3071);
nand U3522 (N_3522,N_3226,N_3289);
nand U3523 (N_3523,N_3412,N_3211);
or U3524 (N_3524,N_3162,N_3061);
and U3525 (N_3525,N_3111,N_3339);
xor U3526 (N_3526,N_3381,N_3421);
xnor U3527 (N_3527,N_3002,N_3471);
xnor U3528 (N_3528,N_3491,N_3207);
nor U3529 (N_3529,N_3408,N_3334);
nand U3530 (N_3530,N_3012,N_3273);
xor U3531 (N_3531,N_3452,N_3213);
nor U3532 (N_3532,N_3178,N_3464);
xor U3533 (N_3533,N_3304,N_3040);
nand U3534 (N_3534,N_3478,N_3070);
or U3535 (N_3535,N_3065,N_3468);
and U3536 (N_3536,N_3416,N_3020);
or U3537 (N_3537,N_3377,N_3081);
nor U3538 (N_3538,N_3414,N_3209);
or U3539 (N_3539,N_3054,N_3128);
nor U3540 (N_3540,N_3482,N_3248);
nand U3541 (N_3541,N_3068,N_3346);
nand U3542 (N_3542,N_3260,N_3082);
nor U3543 (N_3543,N_3141,N_3287);
or U3544 (N_3544,N_3087,N_3426);
nor U3545 (N_3545,N_3234,N_3411);
or U3546 (N_3546,N_3256,N_3484);
xor U3547 (N_3547,N_3341,N_3161);
nand U3548 (N_3548,N_3024,N_3158);
nor U3549 (N_3549,N_3218,N_3157);
nand U3550 (N_3550,N_3429,N_3324);
and U3551 (N_3551,N_3135,N_3221);
nor U3552 (N_3552,N_3163,N_3492);
xnor U3553 (N_3553,N_3035,N_3000);
or U3554 (N_3554,N_3046,N_3127);
and U3555 (N_3555,N_3370,N_3448);
nor U3556 (N_3556,N_3169,N_3499);
or U3557 (N_3557,N_3297,N_3208);
or U3558 (N_3558,N_3494,N_3319);
or U3559 (N_3559,N_3280,N_3115);
or U3560 (N_3560,N_3415,N_3188);
and U3561 (N_3561,N_3258,N_3025);
nand U3562 (N_3562,N_3080,N_3291);
nand U3563 (N_3563,N_3224,N_3362);
or U3564 (N_3564,N_3233,N_3239);
xnor U3565 (N_3565,N_3299,N_3050);
or U3566 (N_3566,N_3393,N_3250);
nand U3567 (N_3567,N_3252,N_3434);
nand U3568 (N_3568,N_3329,N_3198);
or U3569 (N_3569,N_3347,N_3197);
xor U3570 (N_3570,N_3182,N_3456);
or U3571 (N_3571,N_3463,N_3166);
nand U3572 (N_3572,N_3298,N_3243);
xor U3573 (N_3573,N_3172,N_3441);
and U3574 (N_3574,N_3194,N_3193);
nand U3575 (N_3575,N_3259,N_3453);
nand U3576 (N_3576,N_3074,N_3123);
or U3577 (N_3577,N_3493,N_3321);
xor U3578 (N_3578,N_3345,N_3326);
nand U3579 (N_3579,N_3450,N_3380);
and U3580 (N_3580,N_3026,N_3325);
nand U3581 (N_3581,N_3044,N_3296);
and U3582 (N_3582,N_3496,N_3033);
and U3583 (N_3583,N_3160,N_3394);
nor U3584 (N_3584,N_3306,N_3190);
nand U3585 (N_3585,N_3047,N_3097);
or U3586 (N_3586,N_3433,N_3227);
nor U3587 (N_3587,N_3112,N_3184);
xor U3588 (N_3588,N_3352,N_3419);
or U3589 (N_3589,N_3094,N_3018);
and U3590 (N_3590,N_3417,N_3389);
nand U3591 (N_3591,N_3171,N_3454);
or U3592 (N_3592,N_3486,N_3053);
nor U3593 (N_3593,N_3440,N_3311);
or U3594 (N_3594,N_3320,N_3420);
nand U3595 (N_3595,N_3257,N_3058);
nand U3596 (N_3596,N_3125,N_3129);
and U3597 (N_3597,N_3401,N_3375);
nor U3598 (N_3598,N_3130,N_3409);
nand U3599 (N_3599,N_3055,N_3202);
and U3600 (N_3600,N_3118,N_3254);
or U3601 (N_3601,N_3430,N_3479);
nand U3602 (N_3602,N_3147,N_3146);
and U3603 (N_3603,N_3388,N_3108);
or U3604 (N_3604,N_3268,N_3364);
or U3605 (N_3605,N_3351,N_3003);
xor U3606 (N_3606,N_3144,N_3398);
xor U3607 (N_3607,N_3170,N_3210);
and U3608 (N_3608,N_3480,N_3487);
and U3609 (N_3609,N_3117,N_3283);
xor U3610 (N_3610,N_3469,N_3315);
nand U3611 (N_3611,N_3110,N_3309);
nand U3612 (N_3612,N_3088,N_3271);
nor U3613 (N_3613,N_3266,N_3028);
or U3614 (N_3614,N_3472,N_3225);
or U3615 (N_3615,N_3159,N_3383);
and U3616 (N_3616,N_3090,N_3278);
nand U3617 (N_3617,N_3140,N_3067);
xor U3618 (N_3618,N_3041,N_3009);
nor U3619 (N_3619,N_3253,N_3124);
nor U3620 (N_3620,N_3089,N_3425);
or U3621 (N_3621,N_3302,N_3010);
nor U3622 (N_3622,N_3473,N_3338);
or U3623 (N_3623,N_3154,N_3066);
xnor U3624 (N_3624,N_3078,N_3455);
nor U3625 (N_3625,N_3063,N_3336);
nor U3626 (N_3626,N_3385,N_3116);
xnor U3627 (N_3627,N_3145,N_3051);
and U3628 (N_3628,N_3143,N_3481);
xnor U3629 (N_3629,N_3354,N_3312);
or U3630 (N_3630,N_3413,N_3107);
nand U3631 (N_3631,N_3263,N_3092);
and U3632 (N_3632,N_3474,N_3337);
and U3633 (N_3633,N_3236,N_3077);
nor U3634 (N_3634,N_3437,N_3436);
and U3635 (N_3635,N_3151,N_3174);
nand U3636 (N_3636,N_3431,N_3242);
nor U3637 (N_3637,N_3137,N_3164);
nand U3638 (N_3638,N_3103,N_3037);
xor U3639 (N_3639,N_3305,N_3477);
xnor U3640 (N_3640,N_3121,N_3060);
nor U3641 (N_3641,N_3269,N_3084);
and U3642 (N_3642,N_3232,N_3353);
nor U3643 (N_3643,N_3367,N_3428);
xnor U3644 (N_3644,N_3438,N_3176);
and U3645 (N_3645,N_3222,N_3148);
and U3646 (N_3646,N_3284,N_3294);
and U3647 (N_3647,N_3203,N_3049);
or U3648 (N_3648,N_3310,N_3057);
nand U3649 (N_3649,N_3457,N_3014);
nand U3650 (N_3650,N_3004,N_3156);
or U3651 (N_3651,N_3475,N_3376);
xnor U3652 (N_3652,N_3189,N_3272);
nand U3653 (N_3653,N_3458,N_3056);
nand U3654 (N_3654,N_3368,N_3228);
and U3655 (N_3655,N_3072,N_3181);
nand U3656 (N_3656,N_3245,N_3318);
or U3657 (N_3657,N_3330,N_3490);
xnor U3658 (N_3658,N_3183,N_3333);
or U3659 (N_3659,N_3007,N_3085);
nand U3660 (N_3660,N_3031,N_3251);
and U3661 (N_3661,N_3192,N_3186);
and U3662 (N_3662,N_3264,N_3403);
or U3663 (N_3663,N_3465,N_3132);
or U3664 (N_3664,N_3292,N_3285);
and U3665 (N_3665,N_3261,N_3134);
xor U3666 (N_3666,N_3323,N_3276);
and U3667 (N_3667,N_3390,N_3043);
or U3668 (N_3668,N_3099,N_3369);
nor U3669 (N_3669,N_3255,N_3142);
nor U3670 (N_3670,N_3348,N_3204);
and U3671 (N_3671,N_3314,N_3498);
or U3672 (N_3672,N_3042,N_3340);
xor U3673 (N_3673,N_3350,N_3214);
or U3674 (N_3674,N_3019,N_3317);
nor U3675 (N_3675,N_3435,N_3422);
and U3676 (N_3676,N_3286,N_3126);
or U3677 (N_3677,N_3373,N_3235);
and U3678 (N_3678,N_3476,N_3104);
nor U3679 (N_3679,N_3036,N_3360);
or U3680 (N_3680,N_3136,N_3444);
and U3681 (N_3681,N_3073,N_3076);
xnor U3682 (N_3682,N_3384,N_3201);
nand U3683 (N_3683,N_3219,N_3101);
nand U3684 (N_3684,N_3005,N_3083);
nor U3685 (N_3685,N_3270,N_3462);
nand U3686 (N_3686,N_3048,N_3374);
and U3687 (N_3687,N_3343,N_3206);
and U3688 (N_3688,N_3021,N_3460);
and U3689 (N_3689,N_3307,N_3366);
or U3690 (N_3690,N_3196,N_3249);
nor U3691 (N_3691,N_3372,N_3013);
nand U3692 (N_3692,N_3277,N_3139);
and U3693 (N_3693,N_3275,N_3185);
nand U3694 (N_3694,N_3495,N_3467);
nor U3695 (N_3695,N_3075,N_3017);
nor U3696 (N_3696,N_3295,N_3223);
xor U3697 (N_3697,N_3001,N_3424);
nor U3698 (N_3698,N_3327,N_3488);
and U3699 (N_3699,N_3358,N_3230);
nor U3700 (N_3700,N_3449,N_3404);
or U3701 (N_3701,N_3086,N_3008);
nand U3702 (N_3702,N_3100,N_3215);
nand U3703 (N_3703,N_3432,N_3445);
nor U3704 (N_3704,N_3168,N_3357);
and U3705 (N_3705,N_3093,N_3443);
nand U3706 (N_3706,N_3418,N_3155);
or U3707 (N_3707,N_3267,N_3091);
xor U3708 (N_3708,N_3180,N_3483);
or U3709 (N_3709,N_3392,N_3405);
nand U3710 (N_3710,N_3059,N_3301);
and U3711 (N_3711,N_3423,N_3011);
xor U3712 (N_3712,N_3187,N_3029);
nor U3713 (N_3713,N_3331,N_3152);
and U3714 (N_3714,N_3064,N_3379);
nand U3715 (N_3715,N_3427,N_3265);
nor U3716 (N_3716,N_3220,N_3023);
and U3717 (N_3717,N_3274,N_3335);
xnor U3718 (N_3718,N_3397,N_3052);
and U3719 (N_3719,N_3038,N_3281);
nor U3720 (N_3720,N_3282,N_3109);
nor U3721 (N_3721,N_3119,N_3470);
and U3722 (N_3722,N_3240,N_3167);
xor U3723 (N_3723,N_3138,N_3102);
or U3724 (N_3724,N_3355,N_3342);
xor U3725 (N_3725,N_3175,N_3062);
and U3726 (N_3726,N_3177,N_3361);
and U3727 (N_3727,N_3485,N_3096);
nand U3728 (N_3728,N_3247,N_3200);
xnor U3729 (N_3729,N_3212,N_3022);
and U3730 (N_3730,N_3391,N_3439);
xnor U3731 (N_3731,N_3034,N_3165);
xor U3732 (N_3732,N_3131,N_3238);
nand U3733 (N_3733,N_3191,N_3106);
xor U3734 (N_3734,N_3095,N_3217);
nor U3735 (N_3735,N_3466,N_3461);
nand U3736 (N_3736,N_3308,N_3015);
nor U3737 (N_3737,N_3378,N_3149);
nand U3738 (N_3738,N_3098,N_3150);
nor U3739 (N_3739,N_3244,N_3006);
nor U3740 (N_3740,N_3386,N_3359);
and U3741 (N_3741,N_3322,N_3016);
nand U3742 (N_3742,N_3356,N_3195);
nor U3743 (N_3743,N_3365,N_3229);
xor U3744 (N_3744,N_3410,N_3179);
and U3745 (N_3745,N_3079,N_3400);
nand U3746 (N_3746,N_3279,N_3489);
xnor U3747 (N_3747,N_3459,N_3407);
and U3748 (N_3748,N_3447,N_3069);
or U3749 (N_3749,N_3246,N_3045);
xnor U3750 (N_3750,N_3095,N_3252);
nand U3751 (N_3751,N_3261,N_3310);
nor U3752 (N_3752,N_3364,N_3405);
or U3753 (N_3753,N_3197,N_3468);
or U3754 (N_3754,N_3498,N_3136);
xnor U3755 (N_3755,N_3491,N_3466);
xnor U3756 (N_3756,N_3450,N_3051);
or U3757 (N_3757,N_3203,N_3105);
nor U3758 (N_3758,N_3311,N_3325);
xor U3759 (N_3759,N_3437,N_3478);
nor U3760 (N_3760,N_3316,N_3163);
or U3761 (N_3761,N_3196,N_3004);
nand U3762 (N_3762,N_3355,N_3222);
xor U3763 (N_3763,N_3015,N_3356);
and U3764 (N_3764,N_3052,N_3214);
nor U3765 (N_3765,N_3329,N_3457);
or U3766 (N_3766,N_3471,N_3165);
nor U3767 (N_3767,N_3130,N_3255);
or U3768 (N_3768,N_3041,N_3394);
xor U3769 (N_3769,N_3081,N_3211);
nor U3770 (N_3770,N_3288,N_3298);
nor U3771 (N_3771,N_3198,N_3462);
xnor U3772 (N_3772,N_3156,N_3208);
or U3773 (N_3773,N_3460,N_3277);
xnor U3774 (N_3774,N_3013,N_3335);
or U3775 (N_3775,N_3347,N_3132);
xnor U3776 (N_3776,N_3308,N_3072);
and U3777 (N_3777,N_3485,N_3029);
and U3778 (N_3778,N_3060,N_3449);
and U3779 (N_3779,N_3112,N_3228);
or U3780 (N_3780,N_3322,N_3353);
or U3781 (N_3781,N_3390,N_3471);
or U3782 (N_3782,N_3287,N_3008);
xor U3783 (N_3783,N_3051,N_3304);
and U3784 (N_3784,N_3215,N_3467);
nor U3785 (N_3785,N_3152,N_3020);
nand U3786 (N_3786,N_3277,N_3474);
nand U3787 (N_3787,N_3375,N_3216);
nor U3788 (N_3788,N_3134,N_3346);
and U3789 (N_3789,N_3158,N_3464);
or U3790 (N_3790,N_3163,N_3268);
nor U3791 (N_3791,N_3475,N_3344);
nor U3792 (N_3792,N_3079,N_3044);
nor U3793 (N_3793,N_3262,N_3042);
or U3794 (N_3794,N_3110,N_3224);
xnor U3795 (N_3795,N_3480,N_3144);
xor U3796 (N_3796,N_3226,N_3322);
xnor U3797 (N_3797,N_3304,N_3387);
xnor U3798 (N_3798,N_3068,N_3427);
xor U3799 (N_3799,N_3459,N_3124);
xor U3800 (N_3800,N_3165,N_3263);
or U3801 (N_3801,N_3223,N_3320);
nand U3802 (N_3802,N_3236,N_3395);
nand U3803 (N_3803,N_3432,N_3301);
or U3804 (N_3804,N_3384,N_3252);
or U3805 (N_3805,N_3277,N_3242);
nand U3806 (N_3806,N_3442,N_3307);
xnor U3807 (N_3807,N_3119,N_3008);
xnor U3808 (N_3808,N_3154,N_3136);
or U3809 (N_3809,N_3070,N_3182);
nor U3810 (N_3810,N_3483,N_3090);
or U3811 (N_3811,N_3436,N_3413);
or U3812 (N_3812,N_3072,N_3229);
and U3813 (N_3813,N_3042,N_3330);
or U3814 (N_3814,N_3060,N_3481);
xor U3815 (N_3815,N_3058,N_3267);
xor U3816 (N_3816,N_3196,N_3088);
or U3817 (N_3817,N_3261,N_3027);
or U3818 (N_3818,N_3154,N_3134);
nor U3819 (N_3819,N_3253,N_3132);
and U3820 (N_3820,N_3455,N_3423);
or U3821 (N_3821,N_3346,N_3138);
nand U3822 (N_3822,N_3176,N_3392);
nor U3823 (N_3823,N_3096,N_3079);
xor U3824 (N_3824,N_3134,N_3130);
xor U3825 (N_3825,N_3416,N_3208);
or U3826 (N_3826,N_3390,N_3234);
or U3827 (N_3827,N_3242,N_3149);
nor U3828 (N_3828,N_3142,N_3204);
nor U3829 (N_3829,N_3322,N_3192);
nor U3830 (N_3830,N_3052,N_3251);
and U3831 (N_3831,N_3015,N_3313);
nand U3832 (N_3832,N_3319,N_3384);
and U3833 (N_3833,N_3303,N_3306);
or U3834 (N_3834,N_3250,N_3408);
or U3835 (N_3835,N_3040,N_3078);
nor U3836 (N_3836,N_3337,N_3387);
nor U3837 (N_3837,N_3187,N_3150);
and U3838 (N_3838,N_3169,N_3417);
nor U3839 (N_3839,N_3403,N_3140);
nor U3840 (N_3840,N_3476,N_3303);
and U3841 (N_3841,N_3264,N_3372);
or U3842 (N_3842,N_3169,N_3211);
nand U3843 (N_3843,N_3412,N_3092);
or U3844 (N_3844,N_3284,N_3495);
and U3845 (N_3845,N_3129,N_3021);
or U3846 (N_3846,N_3312,N_3096);
and U3847 (N_3847,N_3397,N_3246);
xor U3848 (N_3848,N_3271,N_3073);
xor U3849 (N_3849,N_3202,N_3028);
or U3850 (N_3850,N_3248,N_3050);
nand U3851 (N_3851,N_3490,N_3289);
or U3852 (N_3852,N_3150,N_3463);
nor U3853 (N_3853,N_3000,N_3103);
xnor U3854 (N_3854,N_3015,N_3282);
nand U3855 (N_3855,N_3432,N_3205);
xnor U3856 (N_3856,N_3277,N_3294);
or U3857 (N_3857,N_3075,N_3348);
nor U3858 (N_3858,N_3014,N_3271);
nor U3859 (N_3859,N_3488,N_3491);
xnor U3860 (N_3860,N_3430,N_3076);
nand U3861 (N_3861,N_3221,N_3469);
nand U3862 (N_3862,N_3470,N_3058);
xor U3863 (N_3863,N_3102,N_3048);
or U3864 (N_3864,N_3109,N_3443);
nor U3865 (N_3865,N_3073,N_3119);
or U3866 (N_3866,N_3058,N_3178);
xor U3867 (N_3867,N_3439,N_3216);
and U3868 (N_3868,N_3395,N_3169);
or U3869 (N_3869,N_3440,N_3290);
or U3870 (N_3870,N_3400,N_3366);
xor U3871 (N_3871,N_3363,N_3228);
and U3872 (N_3872,N_3191,N_3214);
xor U3873 (N_3873,N_3091,N_3405);
and U3874 (N_3874,N_3247,N_3497);
xnor U3875 (N_3875,N_3394,N_3335);
nand U3876 (N_3876,N_3163,N_3051);
or U3877 (N_3877,N_3036,N_3176);
xnor U3878 (N_3878,N_3364,N_3382);
and U3879 (N_3879,N_3009,N_3429);
or U3880 (N_3880,N_3326,N_3251);
and U3881 (N_3881,N_3383,N_3218);
nor U3882 (N_3882,N_3376,N_3287);
nor U3883 (N_3883,N_3026,N_3159);
and U3884 (N_3884,N_3003,N_3368);
xor U3885 (N_3885,N_3254,N_3162);
nand U3886 (N_3886,N_3383,N_3037);
or U3887 (N_3887,N_3064,N_3390);
or U3888 (N_3888,N_3221,N_3400);
and U3889 (N_3889,N_3204,N_3154);
xnor U3890 (N_3890,N_3046,N_3240);
xor U3891 (N_3891,N_3094,N_3110);
nor U3892 (N_3892,N_3186,N_3073);
nor U3893 (N_3893,N_3166,N_3407);
nor U3894 (N_3894,N_3041,N_3374);
and U3895 (N_3895,N_3228,N_3026);
or U3896 (N_3896,N_3484,N_3027);
nand U3897 (N_3897,N_3336,N_3402);
xor U3898 (N_3898,N_3236,N_3338);
nor U3899 (N_3899,N_3384,N_3101);
and U3900 (N_3900,N_3496,N_3136);
or U3901 (N_3901,N_3465,N_3142);
or U3902 (N_3902,N_3045,N_3362);
or U3903 (N_3903,N_3481,N_3474);
nor U3904 (N_3904,N_3208,N_3226);
and U3905 (N_3905,N_3405,N_3084);
xnor U3906 (N_3906,N_3033,N_3082);
or U3907 (N_3907,N_3084,N_3362);
nor U3908 (N_3908,N_3239,N_3444);
xor U3909 (N_3909,N_3445,N_3051);
or U3910 (N_3910,N_3482,N_3253);
xor U3911 (N_3911,N_3123,N_3028);
nor U3912 (N_3912,N_3160,N_3199);
xnor U3913 (N_3913,N_3285,N_3471);
nand U3914 (N_3914,N_3116,N_3439);
xor U3915 (N_3915,N_3110,N_3276);
nand U3916 (N_3916,N_3480,N_3130);
and U3917 (N_3917,N_3442,N_3132);
and U3918 (N_3918,N_3404,N_3386);
nor U3919 (N_3919,N_3129,N_3457);
nand U3920 (N_3920,N_3065,N_3383);
xnor U3921 (N_3921,N_3224,N_3161);
or U3922 (N_3922,N_3477,N_3448);
xor U3923 (N_3923,N_3337,N_3197);
nand U3924 (N_3924,N_3130,N_3290);
nor U3925 (N_3925,N_3013,N_3420);
and U3926 (N_3926,N_3174,N_3048);
nor U3927 (N_3927,N_3380,N_3170);
nor U3928 (N_3928,N_3039,N_3386);
nor U3929 (N_3929,N_3241,N_3211);
xnor U3930 (N_3930,N_3210,N_3238);
xor U3931 (N_3931,N_3146,N_3021);
or U3932 (N_3932,N_3177,N_3107);
and U3933 (N_3933,N_3483,N_3114);
xnor U3934 (N_3934,N_3044,N_3105);
xor U3935 (N_3935,N_3336,N_3451);
and U3936 (N_3936,N_3196,N_3320);
nor U3937 (N_3937,N_3205,N_3076);
nand U3938 (N_3938,N_3058,N_3372);
and U3939 (N_3939,N_3474,N_3031);
and U3940 (N_3940,N_3040,N_3476);
nor U3941 (N_3941,N_3149,N_3125);
and U3942 (N_3942,N_3073,N_3328);
xor U3943 (N_3943,N_3022,N_3452);
and U3944 (N_3944,N_3215,N_3131);
xnor U3945 (N_3945,N_3231,N_3058);
nor U3946 (N_3946,N_3494,N_3129);
or U3947 (N_3947,N_3441,N_3105);
nor U3948 (N_3948,N_3270,N_3199);
xor U3949 (N_3949,N_3482,N_3139);
or U3950 (N_3950,N_3015,N_3009);
xor U3951 (N_3951,N_3208,N_3388);
or U3952 (N_3952,N_3441,N_3391);
nor U3953 (N_3953,N_3457,N_3025);
nor U3954 (N_3954,N_3457,N_3323);
or U3955 (N_3955,N_3327,N_3138);
and U3956 (N_3956,N_3433,N_3212);
and U3957 (N_3957,N_3015,N_3031);
nor U3958 (N_3958,N_3305,N_3365);
xnor U3959 (N_3959,N_3084,N_3495);
or U3960 (N_3960,N_3066,N_3394);
xnor U3961 (N_3961,N_3446,N_3434);
nand U3962 (N_3962,N_3193,N_3484);
xor U3963 (N_3963,N_3432,N_3012);
or U3964 (N_3964,N_3286,N_3005);
nor U3965 (N_3965,N_3452,N_3167);
and U3966 (N_3966,N_3373,N_3329);
or U3967 (N_3967,N_3203,N_3345);
xor U3968 (N_3968,N_3352,N_3109);
and U3969 (N_3969,N_3490,N_3029);
nand U3970 (N_3970,N_3443,N_3199);
xnor U3971 (N_3971,N_3386,N_3329);
nand U3972 (N_3972,N_3182,N_3033);
xor U3973 (N_3973,N_3016,N_3160);
nand U3974 (N_3974,N_3326,N_3245);
or U3975 (N_3975,N_3164,N_3295);
xnor U3976 (N_3976,N_3237,N_3021);
or U3977 (N_3977,N_3227,N_3267);
nor U3978 (N_3978,N_3122,N_3295);
or U3979 (N_3979,N_3125,N_3188);
nand U3980 (N_3980,N_3030,N_3226);
and U3981 (N_3981,N_3047,N_3245);
nor U3982 (N_3982,N_3076,N_3285);
or U3983 (N_3983,N_3456,N_3331);
and U3984 (N_3984,N_3289,N_3181);
nor U3985 (N_3985,N_3059,N_3121);
or U3986 (N_3986,N_3327,N_3055);
or U3987 (N_3987,N_3086,N_3430);
nand U3988 (N_3988,N_3418,N_3229);
or U3989 (N_3989,N_3012,N_3254);
or U3990 (N_3990,N_3366,N_3358);
or U3991 (N_3991,N_3173,N_3005);
nor U3992 (N_3992,N_3148,N_3237);
nor U3993 (N_3993,N_3413,N_3382);
xnor U3994 (N_3994,N_3331,N_3375);
nor U3995 (N_3995,N_3340,N_3344);
nand U3996 (N_3996,N_3161,N_3144);
nor U3997 (N_3997,N_3018,N_3377);
xnor U3998 (N_3998,N_3192,N_3055);
nand U3999 (N_3999,N_3399,N_3184);
or U4000 (N_4000,N_3726,N_3755);
and U4001 (N_4001,N_3993,N_3778);
xor U4002 (N_4002,N_3945,N_3767);
or U4003 (N_4003,N_3903,N_3527);
nor U4004 (N_4004,N_3813,N_3799);
nor U4005 (N_4005,N_3992,N_3591);
and U4006 (N_4006,N_3761,N_3782);
xor U4007 (N_4007,N_3800,N_3821);
or U4008 (N_4008,N_3777,N_3578);
and U4009 (N_4009,N_3811,N_3564);
nand U4010 (N_4010,N_3636,N_3968);
nor U4011 (N_4011,N_3889,N_3931);
xnor U4012 (N_4012,N_3960,N_3852);
xnor U4013 (N_4013,N_3505,N_3856);
or U4014 (N_4014,N_3633,N_3624);
nand U4015 (N_4015,N_3626,N_3601);
or U4016 (N_4016,N_3594,N_3603);
or U4017 (N_4017,N_3619,N_3693);
or U4018 (N_4018,N_3970,N_3609);
xor U4019 (N_4019,N_3611,N_3516);
xor U4020 (N_4020,N_3635,N_3628);
nor U4021 (N_4021,N_3994,N_3886);
xor U4022 (N_4022,N_3969,N_3823);
or U4023 (N_4023,N_3597,N_3937);
or U4024 (N_4024,N_3834,N_3908);
nand U4025 (N_4025,N_3882,N_3736);
and U4026 (N_4026,N_3739,N_3890);
or U4027 (N_4027,N_3538,N_3654);
nor U4028 (N_4028,N_3612,N_3793);
and U4029 (N_4029,N_3589,N_3868);
or U4030 (N_4030,N_3754,N_3731);
and U4031 (N_4031,N_3928,N_3871);
nor U4032 (N_4032,N_3748,N_3849);
or U4033 (N_4033,N_3763,N_3837);
xor U4034 (N_4034,N_3744,N_3796);
or U4035 (N_4035,N_3789,N_3511);
nand U4036 (N_4036,N_3634,N_3714);
or U4037 (N_4037,N_3791,N_3965);
nand U4038 (N_4038,N_3874,N_3632);
nor U4039 (N_4039,N_3547,N_3536);
or U4040 (N_4040,N_3529,N_3776);
nand U4041 (N_4041,N_3764,N_3661);
xnor U4042 (N_4042,N_3618,N_3853);
xor U4043 (N_4043,N_3845,N_3814);
nand U4044 (N_4044,N_3762,N_3985);
nor U4045 (N_4045,N_3947,N_3738);
nand U4046 (N_4046,N_3501,N_3899);
or U4047 (N_4047,N_3808,N_3592);
xnor U4048 (N_4048,N_3866,N_3510);
nand U4049 (N_4049,N_3953,N_3673);
and U4050 (N_4050,N_3923,N_3952);
and U4051 (N_4051,N_3785,N_3700);
and U4052 (N_4052,N_3690,N_3996);
nor U4053 (N_4053,N_3920,N_3936);
and U4054 (N_4054,N_3876,N_3548);
nor U4055 (N_4055,N_3758,N_3540);
xor U4056 (N_4056,N_3695,N_3881);
and U4057 (N_4057,N_3686,N_3981);
and U4058 (N_4058,N_3584,N_3598);
or U4059 (N_4059,N_3961,N_3602);
xor U4060 (N_4060,N_3827,N_3894);
nor U4061 (N_4061,N_3751,N_3949);
xnor U4062 (N_4062,N_3655,N_3519);
nand U4063 (N_4063,N_3508,N_3709);
nor U4064 (N_4064,N_3573,N_3708);
nor U4065 (N_4065,N_3722,N_3566);
nor U4066 (N_4066,N_3787,N_3581);
or U4067 (N_4067,N_3614,N_3604);
and U4068 (N_4068,N_3507,N_3696);
nor U4069 (N_4069,N_3770,N_3746);
nand U4070 (N_4070,N_3599,N_3942);
or U4071 (N_4071,N_3660,N_3650);
or U4072 (N_4072,N_3699,N_3870);
or U4073 (N_4073,N_3518,N_3735);
and U4074 (N_4074,N_3546,N_3561);
xnor U4075 (N_4075,N_3750,N_3804);
and U4076 (N_4076,N_3898,N_3846);
xor U4077 (N_4077,N_3532,N_3840);
nor U4078 (N_4078,N_3930,N_3590);
or U4079 (N_4079,N_3905,N_3829);
nand U4080 (N_4080,N_3506,N_3932);
or U4081 (N_4081,N_3806,N_3753);
xor U4082 (N_4082,N_3613,N_3712);
xnor U4083 (N_4083,N_3583,N_3891);
xnor U4084 (N_4084,N_3523,N_3911);
nor U4085 (N_4085,N_3522,N_3774);
nor U4086 (N_4086,N_3810,N_3623);
nor U4087 (N_4087,N_3986,N_3784);
and U4088 (N_4088,N_3772,N_3860);
xnor U4089 (N_4089,N_3976,N_3902);
nor U4090 (N_4090,N_3545,N_3617);
and U4091 (N_4091,N_3641,N_3557);
xnor U4092 (N_4092,N_3901,N_3677);
nand U4093 (N_4093,N_3848,N_3504);
nor U4094 (N_4094,N_3863,N_3983);
xor U4095 (N_4095,N_3728,N_3732);
or U4096 (N_4096,N_3987,N_3704);
or U4097 (N_4097,N_3734,N_3600);
nand U4098 (N_4098,N_3576,N_3858);
or U4099 (N_4099,N_3727,N_3502);
xor U4100 (N_4100,N_3649,N_3857);
nand U4101 (N_4101,N_3662,N_3659);
and U4102 (N_4102,N_3512,N_3574);
or U4103 (N_4103,N_3797,N_3570);
nand U4104 (N_4104,N_3543,N_3539);
xor U4105 (N_4105,N_3577,N_3657);
or U4106 (N_4106,N_3990,N_3526);
nand U4107 (N_4107,N_3999,N_3706);
and U4108 (N_4108,N_3842,N_3742);
xor U4109 (N_4109,N_3653,N_3652);
nand U4110 (N_4110,N_3517,N_3851);
and U4111 (N_4111,N_3670,N_3995);
or U4112 (N_4112,N_3955,N_3984);
nand U4113 (N_4113,N_3847,N_3817);
and U4114 (N_4114,N_3957,N_3528);
nand U4115 (N_4115,N_3752,N_3741);
and U4116 (N_4116,N_3631,N_3725);
nor U4117 (N_4117,N_3646,N_3718);
and U4118 (N_4118,N_3552,N_3689);
xor U4119 (N_4119,N_3688,N_3922);
nor U4120 (N_4120,N_3558,N_3974);
and U4121 (N_4121,N_3503,N_3958);
nand U4122 (N_4122,N_3831,N_3771);
nand U4123 (N_4123,N_3861,N_3684);
nand U4124 (N_4124,N_3525,N_3766);
nor U4125 (N_4125,N_3559,N_3954);
nor U4126 (N_4126,N_3925,N_3675);
or U4127 (N_4127,N_3674,N_3768);
or U4128 (N_4128,N_3884,N_3524);
nand U4129 (N_4129,N_3521,N_3575);
and U4130 (N_4130,N_3988,N_3586);
and U4131 (N_4131,N_3658,N_3667);
nor U4132 (N_4132,N_3998,N_3531);
xnor U4133 (N_4133,N_3694,N_3825);
and U4134 (N_4134,N_3605,N_3865);
or U4135 (N_4135,N_3835,N_3883);
or U4136 (N_4136,N_3941,N_3839);
nor U4137 (N_4137,N_3702,N_3900);
nand U4138 (N_4138,N_3569,N_3643);
nor U4139 (N_4139,N_3500,N_3756);
nand U4140 (N_4140,N_3801,N_3701);
xnor U4141 (N_4141,N_3982,N_3541);
or U4142 (N_4142,N_3980,N_3724);
nand U4143 (N_4143,N_3879,N_3710);
nand U4144 (N_4144,N_3671,N_3807);
nor U4145 (N_4145,N_3897,N_3888);
nand U4146 (N_4146,N_3838,N_3779);
xnor U4147 (N_4147,N_3615,N_3780);
nand U4148 (N_4148,N_3647,N_3940);
or U4149 (N_4149,N_3924,N_3571);
xor U4150 (N_4150,N_3743,N_3535);
nor U4151 (N_4151,N_3560,N_3864);
nor U4152 (N_4152,N_3610,N_3629);
xor U4153 (N_4153,N_3580,N_3794);
xnor U4154 (N_4154,N_3959,N_3929);
nand U4155 (N_4155,N_3622,N_3562);
or U4156 (N_4156,N_3593,N_3991);
xnor U4157 (N_4157,N_3668,N_3515);
and U4158 (N_4158,N_3703,N_3565);
or U4159 (N_4159,N_3676,N_3509);
nand U4160 (N_4160,N_3933,N_3773);
nand U4161 (N_4161,N_3841,N_3788);
xnor U4162 (N_4162,N_3651,N_3585);
and U4163 (N_4163,N_3715,N_3830);
nor U4164 (N_4164,N_3733,N_3663);
xor U4165 (N_4165,N_3783,N_3859);
or U4166 (N_4166,N_3645,N_3910);
nand U4167 (N_4167,N_3926,N_3716);
xor U4168 (N_4168,N_3582,N_3587);
and U4169 (N_4169,N_3698,N_3775);
and U4170 (N_4170,N_3588,N_3943);
xor U4171 (N_4171,N_3648,N_3549);
nor U4172 (N_4172,N_3912,N_3963);
nor U4173 (N_4173,N_3909,N_3914);
or U4174 (N_4174,N_3544,N_3664);
nor U4175 (N_4175,N_3944,N_3869);
nand U4176 (N_4176,N_3572,N_3828);
and U4177 (N_4177,N_3730,N_3880);
xnor U4178 (N_4178,N_3621,N_3826);
nand U4179 (N_4179,N_3514,N_3805);
xnor U4180 (N_4180,N_3967,N_3973);
nor U4181 (N_4181,N_3935,N_3620);
nand U4182 (N_4182,N_3537,N_3567);
or U4183 (N_4183,N_3946,N_3760);
xor U4184 (N_4184,N_3534,N_3956);
nand U4185 (N_4185,N_3917,N_3563);
xnor U4186 (N_4186,N_3697,N_3885);
or U4187 (N_4187,N_3906,N_3681);
nor U4188 (N_4188,N_3872,N_3579);
and U4189 (N_4189,N_3607,N_3542);
and U4190 (N_4190,N_3627,N_3938);
and U4191 (N_4191,N_3637,N_3692);
and U4192 (N_4192,N_3873,N_3729);
xnor U4193 (N_4193,N_3989,N_3792);
or U4194 (N_4194,N_3669,N_3568);
nor U4195 (N_4195,N_3844,N_3533);
nor U4196 (N_4196,N_3639,N_3972);
and U4197 (N_4197,N_3875,N_3878);
xnor U4198 (N_4198,N_3737,N_3820);
nor U4199 (N_4199,N_3862,N_3608);
xnor U4200 (N_4200,N_3962,N_3950);
nor U4201 (N_4201,N_3665,N_3616);
nand U4202 (N_4202,N_3822,N_3964);
or U4203 (N_4203,N_3893,N_3530);
nand U4204 (N_4204,N_3555,N_3915);
or U4205 (N_4205,N_3802,N_3790);
nand U4206 (N_4206,N_3855,N_3606);
xor U4207 (N_4207,N_3556,N_3713);
and U4208 (N_4208,N_3812,N_3843);
and U4209 (N_4209,N_3749,N_3682);
nor U4210 (N_4210,N_3877,N_3680);
or U4211 (N_4211,N_3717,N_3769);
nor U4212 (N_4212,N_3679,N_3683);
nand U4213 (N_4213,N_3971,N_3720);
or U4214 (N_4214,N_3978,N_3833);
or U4215 (N_4215,N_3818,N_3721);
and U4216 (N_4216,N_3951,N_3997);
xor U4217 (N_4217,N_3832,N_3815);
and U4218 (N_4218,N_3656,N_3892);
or U4219 (N_4219,N_3740,N_3747);
nand U4220 (N_4220,N_3719,N_3850);
or U4221 (N_4221,N_3757,N_3975);
nor U4222 (N_4222,N_3644,N_3795);
nor U4223 (N_4223,N_3685,N_3687);
nand U4224 (N_4224,N_3921,N_3711);
xor U4225 (N_4225,N_3819,N_3895);
xnor U4226 (N_4226,N_3979,N_3642);
nor U4227 (N_4227,N_3678,N_3550);
or U4228 (N_4228,N_3809,N_3836);
xnor U4229 (N_4229,N_3916,N_3596);
xor U4230 (N_4230,N_3939,N_3707);
nand U4231 (N_4231,N_3904,N_3553);
or U4232 (N_4232,N_3907,N_3765);
xnor U4233 (N_4233,N_3625,N_3927);
and U4234 (N_4234,N_3919,N_3640);
xnor U4235 (N_4235,N_3630,N_3723);
nor U4236 (N_4236,N_3513,N_3666);
and U4237 (N_4237,N_3896,N_3781);
or U4238 (N_4238,N_3918,N_3816);
nor U4239 (N_4239,N_3913,N_3824);
xor U4240 (N_4240,N_3691,N_3977);
nor U4241 (N_4241,N_3887,N_3867);
nor U4242 (N_4242,N_3854,N_3554);
and U4243 (N_4243,N_3638,N_3798);
and U4244 (N_4244,N_3786,N_3745);
and U4245 (N_4245,N_3551,N_3520);
or U4246 (N_4246,N_3759,N_3966);
xor U4247 (N_4247,N_3803,N_3705);
nand U4248 (N_4248,N_3672,N_3948);
nor U4249 (N_4249,N_3934,N_3595);
nor U4250 (N_4250,N_3613,N_3959);
and U4251 (N_4251,N_3881,N_3698);
xor U4252 (N_4252,N_3924,N_3949);
nand U4253 (N_4253,N_3541,N_3815);
nand U4254 (N_4254,N_3564,N_3616);
nand U4255 (N_4255,N_3871,N_3783);
nor U4256 (N_4256,N_3863,N_3832);
and U4257 (N_4257,N_3671,N_3992);
nand U4258 (N_4258,N_3979,N_3981);
xor U4259 (N_4259,N_3996,N_3556);
or U4260 (N_4260,N_3971,N_3598);
nor U4261 (N_4261,N_3893,N_3655);
nand U4262 (N_4262,N_3728,N_3787);
nor U4263 (N_4263,N_3798,N_3743);
nor U4264 (N_4264,N_3987,N_3656);
xor U4265 (N_4265,N_3943,N_3647);
nand U4266 (N_4266,N_3645,N_3827);
xor U4267 (N_4267,N_3565,N_3588);
and U4268 (N_4268,N_3762,N_3502);
and U4269 (N_4269,N_3981,N_3915);
and U4270 (N_4270,N_3920,N_3629);
or U4271 (N_4271,N_3549,N_3972);
xnor U4272 (N_4272,N_3968,N_3751);
and U4273 (N_4273,N_3859,N_3549);
or U4274 (N_4274,N_3670,N_3807);
nand U4275 (N_4275,N_3797,N_3603);
nor U4276 (N_4276,N_3622,N_3944);
and U4277 (N_4277,N_3838,N_3515);
and U4278 (N_4278,N_3932,N_3768);
or U4279 (N_4279,N_3542,N_3563);
or U4280 (N_4280,N_3942,N_3580);
xnor U4281 (N_4281,N_3983,N_3954);
or U4282 (N_4282,N_3500,N_3512);
nor U4283 (N_4283,N_3905,N_3655);
xor U4284 (N_4284,N_3504,N_3596);
and U4285 (N_4285,N_3848,N_3655);
or U4286 (N_4286,N_3583,N_3728);
nor U4287 (N_4287,N_3775,N_3735);
and U4288 (N_4288,N_3727,N_3513);
xor U4289 (N_4289,N_3888,N_3864);
and U4290 (N_4290,N_3794,N_3771);
nor U4291 (N_4291,N_3805,N_3880);
and U4292 (N_4292,N_3648,N_3650);
nand U4293 (N_4293,N_3774,N_3770);
nand U4294 (N_4294,N_3899,N_3946);
xnor U4295 (N_4295,N_3621,N_3568);
or U4296 (N_4296,N_3599,N_3529);
nor U4297 (N_4297,N_3643,N_3660);
and U4298 (N_4298,N_3991,N_3837);
or U4299 (N_4299,N_3800,N_3580);
and U4300 (N_4300,N_3904,N_3513);
nand U4301 (N_4301,N_3814,N_3716);
and U4302 (N_4302,N_3860,N_3846);
xnor U4303 (N_4303,N_3699,N_3740);
or U4304 (N_4304,N_3697,N_3635);
nand U4305 (N_4305,N_3522,N_3919);
or U4306 (N_4306,N_3856,N_3537);
nand U4307 (N_4307,N_3916,N_3728);
nor U4308 (N_4308,N_3899,N_3522);
nand U4309 (N_4309,N_3582,N_3667);
and U4310 (N_4310,N_3708,N_3624);
xnor U4311 (N_4311,N_3726,N_3501);
xor U4312 (N_4312,N_3908,N_3999);
and U4313 (N_4313,N_3782,N_3885);
nor U4314 (N_4314,N_3510,N_3958);
and U4315 (N_4315,N_3744,N_3605);
and U4316 (N_4316,N_3644,N_3725);
or U4317 (N_4317,N_3868,N_3732);
xnor U4318 (N_4318,N_3510,N_3651);
or U4319 (N_4319,N_3647,N_3945);
xnor U4320 (N_4320,N_3620,N_3786);
xnor U4321 (N_4321,N_3763,N_3879);
and U4322 (N_4322,N_3671,N_3618);
and U4323 (N_4323,N_3963,N_3733);
and U4324 (N_4324,N_3565,N_3882);
nor U4325 (N_4325,N_3727,N_3948);
and U4326 (N_4326,N_3502,N_3676);
nand U4327 (N_4327,N_3863,N_3719);
nand U4328 (N_4328,N_3792,N_3674);
and U4329 (N_4329,N_3534,N_3743);
or U4330 (N_4330,N_3514,N_3679);
nor U4331 (N_4331,N_3665,N_3931);
nand U4332 (N_4332,N_3726,N_3867);
or U4333 (N_4333,N_3668,N_3650);
nor U4334 (N_4334,N_3661,N_3713);
nor U4335 (N_4335,N_3814,N_3509);
nor U4336 (N_4336,N_3698,N_3659);
nor U4337 (N_4337,N_3599,N_3548);
and U4338 (N_4338,N_3801,N_3714);
xor U4339 (N_4339,N_3906,N_3803);
and U4340 (N_4340,N_3983,N_3979);
nor U4341 (N_4341,N_3739,N_3545);
or U4342 (N_4342,N_3697,N_3937);
or U4343 (N_4343,N_3677,N_3614);
xor U4344 (N_4344,N_3977,N_3827);
xnor U4345 (N_4345,N_3824,N_3975);
or U4346 (N_4346,N_3671,N_3878);
and U4347 (N_4347,N_3671,N_3804);
nor U4348 (N_4348,N_3964,N_3848);
nor U4349 (N_4349,N_3842,N_3533);
and U4350 (N_4350,N_3802,N_3590);
and U4351 (N_4351,N_3839,N_3939);
xor U4352 (N_4352,N_3573,N_3543);
nor U4353 (N_4353,N_3742,N_3642);
nor U4354 (N_4354,N_3740,N_3535);
nor U4355 (N_4355,N_3534,N_3708);
xnor U4356 (N_4356,N_3568,N_3901);
nor U4357 (N_4357,N_3641,N_3573);
and U4358 (N_4358,N_3918,N_3819);
xor U4359 (N_4359,N_3904,N_3644);
xnor U4360 (N_4360,N_3731,N_3728);
nor U4361 (N_4361,N_3664,N_3774);
xor U4362 (N_4362,N_3640,N_3699);
and U4363 (N_4363,N_3938,N_3818);
and U4364 (N_4364,N_3746,N_3661);
xor U4365 (N_4365,N_3890,N_3729);
nand U4366 (N_4366,N_3510,N_3518);
or U4367 (N_4367,N_3900,N_3804);
xor U4368 (N_4368,N_3502,N_3685);
and U4369 (N_4369,N_3618,N_3862);
nor U4370 (N_4370,N_3952,N_3815);
or U4371 (N_4371,N_3606,N_3618);
and U4372 (N_4372,N_3893,N_3952);
and U4373 (N_4373,N_3619,N_3617);
and U4374 (N_4374,N_3540,N_3738);
and U4375 (N_4375,N_3549,N_3698);
or U4376 (N_4376,N_3791,N_3730);
xor U4377 (N_4377,N_3966,N_3850);
nand U4378 (N_4378,N_3831,N_3954);
or U4379 (N_4379,N_3577,N_3555);
nand U4380 (N_4380,N_3655,N_3739);
and U4381 (N_4381,N_3804,N_3566);
nand U4382 (N_4382,N_3843,N_3826);
nand U4383 (N_4383,N_3559,N_3612);
or U4384 (N_4384,N_3629,N_3700);
nor U4385 (N_4385,N_3847,N_3918);
and U4386 (N_4386,N_3538,N_3793);
nand U4387 (N_4387,N_3782,N_3774);
and U4388 (N_4388,N_3679,N_3605);
nor U4389 (N_4389,N_3651,N_3675);
or U4390 (N_4390,N_3626,N_3522);
nor U4391 (N_4391,N_3818,N_3569);
and U4392 (N_4392,N_3543,N_3949);
and U4393 (N_4393,N_3952,N_3651);
nor U4394 (N_4394,N_3610,N_3622);
or U4395 (N_4395,N_3926,N_3830);
nand U4396 (N_4396,N_3684,N_3763);
nor U4397 (N_4397,N_3510,N_3639);
or U4398 (N_4398,N_3920,N_3915);
or U4399 (N_4399,N_3947,N_3856);
nor U4400 (N_4400,N_3588,N_3689);
or U4401 (N_4401,N_3811,N_3735);
and U4402 (N_4402,N_3700,N_3918);
xnor U4403 (N_4403,N_3925,N_3614);
and U4404 (N_4404,N_3643,N_3809);
nor U4405 (N_4405,N_3850,N_3818);
nor U4406 (N_4406,N_3504,N_3872);
or U4407 (N_4407,N_3742,N_3741);
or U4408 (N_4408,N_3845,N_3552);
nor U4409 (N_4409,N_3889,N_3673);
nand U4410 (N_4410,N_3939,N_3937);
and U4411 (N_4411,N_3991,N_3794);
and U4412 (N_4412,N_3892,N_3764);
nor U4413 (N_4413,N_3717,N_3526);
or U4414 (N_4414,N_3850,N_3993);
nand U4415 (N_4415,N_3674,N_3555);
xor U4416 (N_4416,N_3583,N_3917);
and U4417 (N_4417,N_3563,N_3947);
nand U4418 (N_4418,N_3591,N_3707);
and U4419 (N_4419,N_3905,N_3624);
and U4420 (N_4420,N_3852,N_3594);
and U4421 (N_4421,N_3995,N_3529);
or U4422 (N_4422,N_3642,N_3592);
or U4423 (N_4423,N_3869,N_3817);
xnor U4424 (N_4424,N_3876,N_3957);
or U4425 (N_4425,N_3881,N_3612);
xor U4426 (N_4426,N_3780,N_3922);
xnor U4427 (N_4427,N_3886,N_3879);
and U4428 (N_4428,N_3873,N_3552);
or U4429 (N_4429,N_3556,N_3730);
and U4430 (N_4430,N_3671,N_3547);
nand U4431 (N_4431,N_3771,N_3884);
and U4432 (N_4432,N_3961,N_3503);
xor U4433 (N_4433,N_3773,N_3682);
or U4434 (N_4434,N_3880,N_3773);
xnor U4435 (N_4435,N_3580,N_3549);
nand U4436 (N_4436,N_3720,N_3600);
xor U4437 (N_4437,N_3767,N_3527);
or U4438 (N_4438,N_3674,N_3691);
nand U4439 (N_4439,N_3914,N_3630);
and U4440 (N_4440,N_3810,N_3833);
or U4441 (N_4441,N_3606,N_3531);
xor U4442 (N_4442,N_3799,N_3883);
nor U4443 (N_4443,N_3789,N_3918);
or U4444 (N_4444,N_3647,N_3790);
or U4445 (N_4445,N_3788,N_3898);
nand U4446 (N_4446,N_3956,N_3698);
nor U4447 (N_4447,N_3888,N_3941);
xor U4448 (N_4448,N_3810,N_3533);
nand U4449 (N_4449,N_3694,N_3837);
nor U4450 (N_4450,N_3970,N_3742);
nand U4451 (N_4451,N_3587,N_3639);
nor U4452 (N_4452,N_3889,N_3948);
nor U4453 (N_4453,N_3659,N_3758);
or U4454 (N_4454,N_3929,N_3817);
nor U4455 (N_4455,N_3834,N_3563);
and U4456 (N_4456,N_3854,N_3890);
nor U4457 (N_4457,N_3609,N_3742);
nor U4458 (N_4458,N_3945,N_3547);
and U4459 (N_4459,N_3984,N_3736);
xor U4460 (N_4460,N_3805,N_3693);
xor U4461 (N_4461,N_3914,N_3527);
xnor U4462 (N_4462,N_3754,N_3900);
and U4463 (N_4463,N_3621,N_3795);
nor U4464 (N_4464,N_3811,N_3593);
or U4465 (N_4465,N_3627,N_3698);
nand U4466 (N_4466,N_3675,N_3760);
xor U4467 (N_4467,N_3783,N_3751);
nand U4468 (N_4468,N_3939,N_3789);
nand U4469 (N_4469,N_3835,N_3542);
nand U4470 (N_4470,N_3785,N_3550);
and U4471 (N_4471,N_3972,N_3648);
or U4472 (N_4472,N_3995,N_3705);
xor U4473 (N_4473,N_3605,N_3909);
nor U4474 (N_4474,N_3789,N_3629);
or U4475 (N_4475,N_3538,N_3823);
nor U4476 (N_4476,N_3528,N_3985);
xor U4477 (N_4477,N_3803,N_3675);
nor U4478 (N_4478,N_3604,N_3751);
xnor U4479 (N_4479,N_3596,N_3581);
nand U4480 (N_4480,N_3858,N_3579);
or U4481 (N_4481,N_3705,N_3898);
nand U4482 (N_4482,N_3596,N_3740);
or U4483 (N_4483,N_3600,N_3634);
nor U4484 (N_4484,N_3911,N_3711);
nor U4485 (N_4485,N_3988,N_3547);
nand U4486 (N_4486,N_3909,N_3675);
or U4487 (N_4487,N_3532,N_3736);
and U4488 (N_4488,N_3960,N_3963);
nand U4489 (N_4489,N_3997,N_3750);
or U4490 (N_4490,N_3693,N_3691);
nor U4491 (N_4491,N_3622,N_3641);
nor U4492 (N_4492,N_3598,N_3627);
nand U4493 (N_4493,N_3680,N_3540);
or U4494 (N_4494,N_3619,N_3815);
or U4495 (N_4495,N_3902,N_3545);
nor U4496 (N_4496,N_3580,N_3736);
and U4497 (N_4497,N_3579,N_3732);
nand U4498 (N_4498,N_3717,N_3706);
nand U4499 (N_4499,N_3997,N_3715);
nand U4500 (N_4500,N_4091,N_4305);
nor U4501 (N_4501,N_4063,N_4335);
and U4502 (N_4502,N_4077,N_4172);
xor U4503 (N_4503,N_4245,N_4273);
xnor U4504 (N_4504,N_4035,N_4226);
nand U4505 (N_4505,N_4036,N_4376);
or U4506 (N_4506,N_4332,N_4361);
or U4507 (N_4507,N_4186,N_4067);
nand U4508 (N_4508,N_4040,N_4331);
xor U4509 (N_4509,N_4086,N_4194);
nor U4510 (N_4510,N_4400,N_4025);
xor U4511 (N_4511,N_4125,N_4060);
xor U4512 (N_4512,N_4492,N_4249);
xor U4513 (N_4513,N_4047,N_4113);
or U4514 (N_4514,N_4201,N_4151);
nor U4515 (N_4515,N_4355,N_4014);
or U4516 (N_4516,N_4246,N_4394);
and U4517 (N_4517,N_4437,N_4193);
nand U4518 (N_4518,N_4037,N_4208);
nand U4519 (N_4519,N_4428,N_4433);
nand U4520 (N_4520,N_4384,N_4257);
or U4521 (N_4521,N_4385,N_4300);
nor U4522 (N_4522,N_4184,N_4110);
nand U4523 (N_4523,N_4468,N_4476);
xor U4524 (N_4524,N_4012,N_4311);
nand U4525 (N_4525,N_4043,N_4371);
nand U4526 (N_4526,N_4416,N_4262);
or U4527 (N_4527,N_4239,N_4165);
or U4528 (N_4528,N_4176,N_4189);
nor U4529 (N_4529,N_4150,N_4408);
nand U4530 (N_4530,N_4350,N_4209);
xnor U4531 (N_4531,N_4268,N_4310);
nand U4532 (N_4532,N_4248,N_4377);
nand U4533 (N_4533,N_4022,N_4164);
xnor U4534 (N_4534,N_4061,N_4382);
xnor U4535 (N_4535,N_4316,N_4052);
nor U4536 (N_4536,N_4017,N_4308);
xor U4537 (N_4537,N_4159,N_4409);
or U4538 (N_4538,N_4447,N_4432);
nor U4539 (N_4539,N_4030,N_4028);
or U4540 (N_4540,N_4267,N_4140);
or U4541 (N_4541,N_4190,N_4281);
xnor U4542 (N_4542,N_4462,N_4117);
nor U4543 (N_4543,N_4352,N_4356);
nor U4544 (N_4544,N_4469,N_4059);
xnor U4545 (N_4545,N_4290,N_4001);
xor U4546 (N_4546,N_4450,N_4082);
xor U4547 (N_4547,N_4284,N_4103);
xor U4548 (N_4548,N_4449,N_4474);
and U4549 (N_4549,N_4288,N_4473);
or U4550 (N_4550,N_4235,N_4013);
nand U4551 (N_4551,N_4326,N_4074);
nor U4552 (N_4552,N_4481,N_4057);
or U4553 (N_4553,N_4141,N_4445);
xor U4554 (N_4554,N_4265,N_4405);
and U4555 (N_4555,N_4031,N_4497);
and U4556 (N_4556,N_4324,N_4272);
and U4557 (N_4557,N_4049,N_4493);
and U4558 (N_4558,N_4083,N_4198);
and U4559 (N_4559,N_4155,N_4419);
nor U4560 (N_4560,N_4005,N_4329);
and U4561 (N_4561,N_4283,N_4487);
nor U4562 (N_4562,N_4375,N_4348);
and U4563 (N_4563,N_4475,N_4102);
and U4564 (N_4564,N_4156,N_4451);
xor U4565 (N_4565,N_4282,N_4051);
xor U4566 (N_4566,N_4360,N_4423);
xor U4567 (N_4567,N_4130,N_4232);
or U4568 (N_4568,N_4230,N_4336);
nand U4569 (N_4569,N_4259,N_4009);
nand U4570 (N_4570,N_4349,N_4264);
and U4571 (N_4571,N_4179,N_4483);
nor U4572 (N_4572,N_4167,N_4390);
and U4573 (N_4573,N_4065,N_4459);
and U4574 (N_4574,N_4171,N_4307);
nand U4575 (N_4575,N_4149,N_4136);
or U4576 (N_4576,N_4023,N_4453);
xor U4577 (N_4577,N_4489,N_4106);
nor U4578 (N_4578,N_4027,N_4018);
and U4579 (N_4579,N_4442,N_4285);
xor U4580 (N_4580,N_4147,N_4068);
xor U4581 (N_4581,N_4032,N_4217);
nor U4582 (N_4582,N_4048,N_4266);
nand U4583 (N_4583,N_4046,N_4019);
xnor U4584 (N_4584,N_4465,N_4378);
and U4585 (N_4585,N_4407,N_4173);
xor U4586 (N_4586,N_4343,N_4302);
and U4587 (N_4587,N_4139,N_4325);
and U4588 (N_4588,N_4162,N_4116);
nor U4589 (N_4589,N_4389,N_4322);
nor U4590 (N_4590,N_4295,N_4353);
nand U4591 (N_4591,N_4367,N_4188);
or U4592 (N_4592,N_4304,N_4112);
xnor U4593 (N_4593,N_4138,N_4271);
nor U4594 (N_4594,N_4470,N_4085);
or U4595 (N_4595,N_4318,N_4101);
xnor U4596 (N_4596,N_4128,N_4328);
xnor U4597 (N_4597,N_4344,N_4134);
and U4598 (N_4598,N_4253,N_4126);
and U4599 (N_4599,N_4274,N_4477);
or U4600 (N_4600,N_4054,N_4413);
or U4601 (N_4601,N_4105,N_4440);
xnor U4602 (N_4602,N_4157,N_4498);
nand U4603 (N_4603,N_4119,N_4338);
xnor U4604 (N_4604,N_4296,N_4278);
and U4605 (N_4605,N_4287,N_4058);
or U4606 (N_4606,N_4072,N_4491);
nand U4607 (N_4607,N_4369,N_4455);
nor U4608 (N_4608,N_4174,N_4404);
and U4609 (N_4609,N_4132,N_4270);
or U4610 (N_4610,N_4301,N_4321);
and U4611 (N_4611,N_4096,N_4414);
nor U4612 (N_4612,N_4251,N_4045);
nor U4613 (N_4613,N_4438,N_4216);
xor U4614 (N_4614,N_4050,N_4062);
or U4615 (N_4615,N_4412,N_4280);
nand U4616 (N_4616,N_4279,N_4206);
or U4617 (N_4617,N_4364,N_4418);
or U4618 (N_4618,N_4241,N_4368);
or U4619 (N_4619,N_4247,N_4426);
nor U4620 (N_4620,N_4381,N_4143);
xor U4621 (N_4621,N_4000,N_4224);
nor U4622 (N_4622,N_4160,N_4185);
xnor U4623 (N_4623,N_4238,N_4029);
or U4624 (N_4624,N_4439,N_4341);
xor U4625 (N_4625,N_4098,N_4292);
nor U4626 (N_4626,N_4212,N_4457);
nor U4627 (N_4627,N_4215,N_4395);
nand U4628 (N_4628,N_4242,N_4410);
nor U4629 (N_4629,N_4118,N_4231);
xor U4630 (N_4630,N_4435,N_4214);
nand U4631 (N_4631,N_4056,N_4456);
nand U4632 (N_4632,N_4181,N_4454);
or U4633 (N_4633,N_4354,N_4084);
nand U4634 (N_4634,N_4261,N_4298);
or U4635 (N_4635,N_4195,N_4007);
and U4636 (N_4636,N_4494,N_4145);
nand U4637 (N_4637,N_4297,N_4041);
and U4638 (N_4638,N_4004,N_4166);
or U4639 (N_4639,N_4221,N_4120);
nor U4640 (N_4640,N_4396,N_4357);
nand U4641 (N_4641,N_4109,N_4299);
xnor U4642 (N_4642,N_4406,N_4011);
or U4643 (N_4643,N_4129,N_4383);
nand U4644 (N_4644,N_4127,N_4071);
and U4645 (N_4645,N_4220,N_4202);
nor U4646 (N_4646,N_4170,N_4327);
and U4647 (N_4647,N_4076,N_4399);
nand U4648 (N_4648,N_4227,N_4183);
xnor U4649 (N_4649,N_4393,N_4380);
nand U4650 (N_4650,N_4003,N_4291);
xnor U4651 (N_4651,N_4340,N_4496);
and U4652 (N_4652,N_4342,N_4225);
and U4653 (N_4653,N_4484,N_4234);
or U4654 (N_4654,N_4169,N_4191);
or U4655 (N_4655,N_4320,N_4345);
or U4656 (N_4656,N_4448,N_4482);
and U4657 (N_4657,N_4233,N_4275);
xnor U4658 (N_4658,N_4252,N_4055);
xor U4659 (N_4659,N_4124,N_4314);
nand U4660 (N_4660,N_4333,N_4488);
nand U4661 (N_4661,N_4420,N_4269);
nand U4662 (N_4662,N_4016,N_4089);
nand U4663 (N_4663,N_4010,N_4163);
nand U4664 (N_4664,N_4108,N_4152);
nor U4665 (N_4665,N_4460,N_4315);
nand U4666 (N_4666,N_4236,N_4339);
nor U4667 (N_4667,N_4372,N_4200);
nand U4668 (N_4668,N_4480,N_4008);
or U4669 (N_4669,N_4417,N_4095);
xnor U4670 (N_4670,N_4244,N_4452);
nor U4671 (N_4671,N_4490,N_4218);
xor U4672 (N_4672,N_4064,N_4180);
xnor U4673 (N_4673,N_4122,N_4430);
and U4674 (N_4674,N_4207,N_4254);
xor U4675 (N_4675,N_4197,N_4351);
xor U4676 (N_4676,N_4079,N_4359);
nor U4677 (N_4677,N_4222,N_4002);
nor U4678 (N_4678,N_4177,N_4427);
xor U4679 (N_4679,N_4346,N_4114);
xor U4680 (N_4680,N_4024,N_4075);
nand U4681 (N_4681,N_4429,N_4153);
nor U4682 (N_4682,N_4317,N_4443);
or U4683 (N_4683,N_4038,N_4158);
and U4684 (N_4684,N_4495,N_4020);
and U4685 (N_4685,N_4458,N_4323);
nand U4686 (N_4686,N_4363,N_4373);
or U4687 (N_4687,N_4306,N_4366);
nand U4688 (N_4688,N_4277,N_4203);
nor U4689 (N_4689,N_4276,N_4379);
nor U4690 (N_4690,N_4478,N_4263);
nor U4691 (N_4691,N_4078,N_4178);
xor U4692 (N_4692,N_4100,N_4256);
nor U4693 (N_4693,N_4303,N_4391);
nand U4694 (N_4694,N_4388,N_4196);
nand U4695 (N_4695,N_4199,N_4467);
xor U4696 (N_4696,N_4499,N_4090);
or U4697 (N_4697,N_4133,N_4365);
xor U4698 (N_4698,N_4088,N_4415);
nand U4699 (N_4699,N_4260,N_4210);
or U4700 (N_4700,N_4081,N_4204);
nor U4701 (N_4701,N_4123,N_4104);
xnor U4702 (N_4702,N_4431,N_4289);
xor U4703 (N_4703,N_4485,N_4182);
nand U4704 (N_4704,N_4099,N_4312);
or U4705 (N_4705,N_4034,N_4015);
xor U4706 (N_4706,N_4347,N_4161);
xnor U4707 (N_4707,N_4142,N_4080);
xor U4708 (N_4708,N_4131,N_4403);
nand U4709 (N_4709,N_4334,N_4187);
or U4710 (N_4710,N_4211,N_4472);
or U4711 (N_4711,N_4309,N_4137);
nand U4712 (N_4712,N_4436,N_4111);
nor U4713 (N_4713,N_4471,N_4397);
and U4714 (N_4714,N_4069,N_4337);
xnor U4715 (N_4715,N_4370,N_4286);
and U4716 (N_4716,N_4107,N_4093);
nand U4717 (N_4717,N_4402,N_4135);
xnor U4718 (N_4718,N_4479,N_4087);
nor U4719 (N_4719,N_4044,N_4464);
and U4720 (N_4720,N_4401,N_4148);
xnor U4721 (N_4721,N_4255,N_4319);
and U4722 (N_4722,N_4066,N_4121);
or U4723 (N_4723,N_4042,N_4374);
nor U4724 (N_4724,N_4258,N_4228);
nor U4725 (N_4725,N_4229,N_4421);
nor U4726 (N_4726,N_4094,N_4073);
and U4727 (N_4727,N_4205,N_4033);
or U4728 (N_4728,N_4039,N_4387);
and U4729 (N_4729,N_4293,N_4237);
or U4730 (N_4730,N_4154,N_4219);
nor U4731 (N_4731,N_4386,N_4243);
xor U4732 (N_4732,N_4398,N_4146);
xor U4733 (N_4733,N_4021,N_4358);
or U4734 (N_4734,N_4250,N_4330);
nand U4735 (N_4735,N_4313,N_4006);
nand U4736 (N_4736,N_4392,N_4240);
or U4737 (N_4737,N_4223,N_4441);
xnor U4738 (N_4738,N_4026,N_4444);
or U4739 (N_4739,N_4466,N_4053);
xor U4740 (N_4740,N_4144,N_4362);
or U4741 (N_4741,N_4463,N_4168);
and U4742 (N_4742,N_4092,N_4486);
nand U4743 (N_4743,N_4097,N_4213);
or U4744 (N_4744,N_4425,N_4192);
or U4745 (N_4745,N_4070,N_4115);
nand U4746 (N_4746,N_4422,N_4461);
xnor U4747 (N_4747,N_4294,N_4446);
xnor U4748 (N_4748,N_4175,N_4411);
or U4749 (N_4749,N_4434,N_4424);
nor U4750 (N_4750,N_4312,N_4157);
nor U4751 (N_4751,N_4078,N_4046);
xnor U4752 (N_4752,N_4393,N_4333);
xor U4753 (N_4753,N_4202,N_4493);
nor U4754 (N_4754,N_4018,N_4331);
and U4755 (N_4755,N_4347,N_4278);
nor U4756 (N_4756,N_4052,N_4416);
and U4757 (N_4757,N_4421,N_4182);
xor U4758 (N_4758,N_4187,N_4228);
or U4759 (N_4759,N_4243,N_4300);
and U4760 (N_4760,N_4479,N_4074);
nand U4761 (N_4761,N_4117,N_4141);
nand U4762 (N_4762,N_4129,N_4304);
nor U4763 (N_4763,N_4437,N_4240);
and U4764 (N_4764,N_4438,N_4331);
and U4765 (N_4765,N_4113,N_4032);
nand U4766 (N_4766,N_4366,N_4072);
xnor U4767 (N_4767,N_4050,N_4396);
nor U4768 (N_4768,N_4333,N_4014);
or U4769 (N_4769,N_4042,N_4262);
and U4770 (N_4770,N_4120,N_4070);
nor U4771 (N_4771,N_4219,N_4165);
and U4772 (N_4772,N_4246,N_4164);
nand U4773 (N_4773,N_4192,N_4242);
and U4774 (N_4774,N_4410,N_4399);
nor U4775 (N_4775,N_4455,N_4492);
nand U4776 (N_4776,N_4432,N_4337);
xor U4777 (N_4777,N_4060,N_4040);
nor U4778 (N_4778,N_4159,N_4126);
xor U4779 (N_4779,N_4430,N_4121);
or U4780 (N_4780,N_4405,N_4125);
xnor U4781 (N_4781,N_4120,N_4415);
and U4782 (N_4782,N_4088,N_4148);
xor U4783 (N_4783,N_4397,N_4282);
nor U4784 (N_4784,N_4187,N_4410);
and U4785 (N_4785,N_4411,N_4278);
xor U4786 (N_4786,N_4192,N_4299);
nand U4787 (N_4787,N_4484,N_4388);
nand U4788 (N_4788,N_4117,N_4318);
nor U4789 (N_4789,N_4078,N_4081);
nor U4790 (N_4790,N_4146,N_4085);
xnor U4791 (N_4791,N_4090,N_4410);
nand U4792 (N_4792,N_4495,N_4367);
nor U4793 (N_4793,N_4016,N_4400);
xor U4794 (N_4794,N_4317,N_4062);
and U4795 (N_4795,N_4457,N_4210);
nor U4796 (N_4796,N_4302,N_4201);
xor U4797 (N_4797,N_4388,N_4498);
nand U4798 (N_4798,N_4449,N_4125);
or U4799 (N_4799,N_4048,N_4151);
and U4800 (N_4800,N_4053,N_4400);
nand U4801 (N_4801,N_4412,N_4346);
nand U4802 (N_4802,N_4461,N_4328);
and U4803 (N_4803,N_4051,N_4274);
or U4804 (N_4804,N_4420,N_4241);
or U4805 (N_4805,N_4288,N_4150);
xor U4806 (N_4806,N_4071,N_4129);
nor U4807 (N_4807,N_4366,N_4040);
or U4808 (N_4808,N_4316,N_4381);
nand U4809 (N_4809,N_4271,N_4088);
or U4810 (N_4810,N_4006,N_4039);
xnor U4811 (N_4811,N_4249,N_4337);
or U4812 (N_4812,N_4305,N_4124);
and U4813 (N_4813,N_4101,N_4019);
xor U4814 (N_4814,N_4287,N_4089);
nand U4815 (N_4815,N_4049,N_4130);
nor U4816 (N_4816,N_4020,N_4393);
xor U4817 (N_4817,N_4272,N_4091);
xnor U4818 (N_4818,N_4051,N_4496);
nand U4819 (N_4819,N_4251,N_4261);
xnor U4820 (N_4820,N_4459,N_4247);
nand U4821 (N_4821,N_4174,N_4402);
and U4822 (N_4822,N_4324,N_4200);
nor U4823 (N_4823,N_4437,N_4211);
or U4824 (N_4824,N_4203,N_4036);
xor U4825 (N_4825,N_4068,N_4369);
nand U4826 (N_4826,N_4032,N_4414);
and U4827 (N_4827,N_4489,N_4323);
or U4828 (N_4828,N_4201,N_4313);
nand U4829 (N_4829,N_4409,N_4115);
nand U4830 (N_4830,N_4039,N_4392);
xnor U4831 (N_4831,N_4080,N_4049);
and U4832 (N_4832,N_4325,N_4406);
and U4833 (N_4833,N_4197,N_4138);
nand U4834 (N_4834,N_4442,N_4492);
nand U4835 (N_4835,N_4402,N_4088);
nand U4836 (N_4836,N_4441,N_4180);
and U4837 (N_4837,N_4481,N_4458);
nor U4838 (N_4838,N_4099,N_4085);
xor U4839 (N_4839,N_4112,N_4276);
nand U4840 (N_4840,N_4231,N_4283);
or U4841 (N_4841,N_4399,N_4329);
and U4842 (N_4842,N_4015,N_4092);
xnor U4843 (N_4843,N_4207,N_4108);
or U4844 (N_4844,N_4070,N_4127);
nand U4845 (N_4845,N_4468,N_4021);
nor U4846 (N_4846,N_4309,N_4108);
or U4847 (N_4847,N_4375,N_4229);
or U4848 (N_4848,N_4338,N_4118);
or U4849 (N_4849,N_4105,N_4289);
xnor U4850 (N_4850,N_4227,N_4343);
xor U4851 (N_4851,N_4199,N_4103);
nand U4852 (N_4852,N_4196,N_4010);
or U4853 (N_4853,N_4050,N_4013);
nor U4854 (N_4854,N_4205,N_4258);
and U4855 (N_4855,N_4102,N_4009);
and U4856 (N_4856,N_4435,N_4293);
nor U4857 (N_4857,N_4474,N_4265);
nand U4858 (N_4858,N_4095,N_4243);
and U4859 (N_4859,N_4305,N_4076);
xnor U4860 (N_4860,N_4113,N_4281);
and U4861 (N_4861,N_4390,N_4189);
and U4862 (N_4862,N_4108,N_4296);
xor U4863 (N_4863,N_4387,N_4214);
or U4864 (N_4864,N_4129,N_4140);
or U4865 (N_4865,N_4017,N_4428);
nor U4866 (N_4866,N_4312,N_4365);
xnor U4867 (N_4867,N_4373,N_4456);
or U4868 (N_4868,N_4150,N_4446);
xor U4869 (N_4869,N_4140,N_4245);
or U4870 (N_4870,N_4299,N_4226);
and U4871 (N_4871,N_4010,N_4152);
nand U4872 (N_4872,N_4415,N_4383);
and U4873 (N_4873,N_4490,N_4092);
or U4874 (N_4874,N_4280,N_4124);
nor U4875 (N_4875,N_4132,N_4450);
xor U4876 (N_4876,N_4042,N_4267);
or U4877 (N_4877,N_4243,N_4337);
nor U4878 (N_4878,N_4357,N_4352);
nand U4879 (N_4879,N_4088,N_4346);
or U4880 (N_4880,N_4096,N_4262);
nor U4881 (N_4881,N_4287,N_4377);
xnor U4882 (N_4882,N_4348,N_4225);
xnor U4883 (N_4883,N_4416,N_4343);
or U4884 (N_4884,N_4201,N_4175);
xor U4885 (N_4885,N_4164,N_4103);
or U4886 (N_4886,N_4250,N_4392);
and U4887 (N_4887,N_4493,N_4325);
nor U4888 (N_4888,N_4123,N_4327);
or U4889 (N_4889,N_4208,N_4337);
xor U4890 (N_4890,N_4301,N_4152);
xor U4891 (N_4891,N_4398,N_4205);
nor U4892 (N_4892,N_4230,N_4481);
or U4893 (N_4893,N_4481,N_4180);
xor U4894 (N_4894,N_4233,N_4025);
nand U4895 (N_4895,N_4066,N_4360);
xnor U4896 (N_4896,N_4438,N_4319);
or U4897 (N_4897,N_4262,N_4112);
nand U4898 (N_4898,N_4141,N_4030);
nor U4899 (N_4899,N_4004,N_4469);
and U4900 (N_4900,N_4339,N_4239);
nand U4901 (N_4901,N_4167,N_4415);
or U4902 (N_4902,N_4301,N_4367);
nor U4903 (N_4903,N_4488,N_4224);
nor U4904 (N_4904,N_4472,N_4196);
xnor U4905 (N_4905,N_4085,N_4290);
xor U4906 (N_4906,N_4219,N_4228);
nor U4907 (N_4907,N_4280,N_4331);
or U4908 (N_4908,N_4034,N_4499);
nor U4909 (N_4909,N_4109,N_4203);
and U4910 (N_4910,N_4374,N_4437);
nand U4911 (N_4911,N_4251,N_4068);
or U4912 (N_4912,N_4220,N_4169);
nor U4913 (N_4913,N_4301,N_4194);
nand U4914 (N_4914,N_4113,N_4176);
xor U4915 (N_4915,N_4231,N_4171);
xnor U4916 (N_4916,N_4046,N_4466);
nor U4917 (N_4917,N_4484,N_4495);
nand U4918 (N_4918,N_4185,N_4360);
xnor U4919 (N_4919,N_4078,N_4228);
or U4920 (N_4920,N_4041,N_4069);
and U4921 (N_4921,N_4063,N_4243);
or U4922 (N_4922,N_4462,N_4060);
or U4923 (N_4923,N_4055,N_4209);
or U4924 (N_4924,N_4453,N_4239);
and U4925 (N_4925,N_4105,N_4388);
and U4926 (N_4926,N_4420,N_4135);
nor U4927 (N_4927,N_4217,N_4010);
nor U4928 (N_4928,N_4209,N_4409);
nand U4929 (N_4929,N_4102,N_4035);
nand U4930 (N_4930,N_4334,N_4425);
and U4931 (N_4931,N_4228,N_4411);
and U4932 (N_4932,N_4458,N_4421);
nor U4933 (N_4933,N_4211,N_4353);
nand U4934 (N_4934,N_4396,N_4295);
and U4935 (N_4935,N_4161,N_4322);
and U4936 (N_4936,N_4489,N_4192);
xnor U4937 (N_4937,N_4298,N_4204);
xnor U4938 (N_4938,N_4248,N_4002);
xnor U4939 (N_4939,N_4023,N_4298);
nand U4940 (N_4940,N_4045,N_4491);
and U4941 (N_4941,N_4463,N_4331);
xnor U4942 (N_4942,N_4200,N_4444);
nand U4943 (N_4943,N_4025,N_4029);
or U4944 (N_4944,N_4225,N_4194);
and U4945 (N_4945,N_4080,N_4010);
and U4946 (N_4946,N_4417,N_4381);
nand U4947 (N_4947,N_4496,N_4110);
or U4948 (N_4948,N_4303,N_4360);
nand U4949 (N_4949,N_4179,N_4005);
and U4950 (N_4950,N_4318,N_4023);
or U4951 (N_4951,N_4062,N_4217);
nand U4952 (N_4952,N_4383,N_4476);
nand U4953 (N_4953,N_4279,N_4281);
nor U4954 (N_4954,N_4004,N_4106);
nand U4955 (N_4955,N_4175,N_4113);
xor U4956 (N_4956,N_4215,N_4368);
and U4957 (N_4957,N_4080,N_4361);
nor U4958 (N_4958,N_4108,N_4097);
and U4959 (N_4959,N_4446,N_4469);
xnor U4960 (N_4960,N_4295,N_4490);
xor U4961 (N_4961,N_4447,N_4129);
and U4962 (N_4962,N_4139,N_4157);
or U4963 (N_4963,N_4147,N_4367);
and U4964 (N_4964,N_4085,N_4276);
nand U4965 (N_4965,N_4465,N_4143);
xnor U4966 (N_4966,N_4188,N_4461);
and U4967 (N_4967,N_4237,N_4344);
nor U4968 (N_4968,N_4438,N_4167);
nor U4969 (N_4969,N_4005,N_4452);
or U4970 (N_4970,N_4132,N_4312);
nor U4971 (N_4971,N_4181,N_4484);
xnor U4972 (N_4972,N_4164,N_4293);
nand U4973 (N_4973,N_4219,N_4351);
nand U4974 (N_4974,N_4482,N_4014);
or U4975 (N_4975,N_4294,N_4471);
nand U4976 (N_4976,N_4173,N_4204);
xnor U4977 (N_4977,N_4491,N_4437);
or U4978 (N_4978,N_4365,N_4045);
and U4979 (N_4979,N_4145,N_4314);
xor U4980 (N_4980,N_4152,N_4046);
nor U4981 (N_4981,N_4076,N_4450);
or U4982 (N_4982,N_4185,N_4188);
and U4983 (N_4983,N_4114,N_4478);
and U4984 (N_4984,N_4145,N_4052);
nor U4985 (N_4985,N_4492,N_4283);
nand U4986 (N_4986,N_4133,N_4173);
or U4987 (N_4987,N_4109,N_4295);
and U4988 (N_4988,N_4007,N_4352);
xnor U4989 (N_4989,N_4463,N_4088);
nor U4990 (N_4990,N_4217,N_4350);
nand U4991 (N_4991,N_4373,N_4157);
nand U4992 (N_4992,N_4409,N_4065);
and U4993 (N_4993,N_4124,N_4165);
and U4994 (N_4994,N_4051,N_4482);
and U4995 (N_4995,N_4300,N_4158);
nand U4996 (N_4996,N_4169,N_4321);
and U4997 (N_4997,N_4080,N_4286);
nor U4998 (N_4998,N_4440,N_4056);
nand U4999 (N_4999,N_4410,N_4317);
nor U5000 (N_5000,N_4710,N_4917);
nor U5001 (N_5001,N_4930,N_4530);
xnor U5002 (N_5002,N_4866,N_4638);
xnor U5003 (N_5003,N_4782,N_4983);
nand U5004 (N_5004,N_4566,N_4745);
nor U5005 (N_5005,N_4807,N_4615);
and U5006 (N_5006,N_4741,N_4814);
or U5007 (N_5007,N_4786,N_4996);
nand U5008 (N_5008,N_4771,N_4751);
nor U5009 (N_5009,N_4598,N_4711);
xor U5010 (N_5010,N_4992,N_4521);
xor U5011 (N_5011,N_4676,N_4664);
or U5012 (N_5012,N_4952,N_4997);
and U5013 (N_5013,N_4858,N_4876);
or U5014 (N_5014,N_4599,N_4731);
nor U5015 (N_5015,N_4763,N_4922);
or U5016 (N_5016,N_4575,N_4647);
nor U5017 (N_5017,N_4901,N_4853);
and U5018 (N_5018,N_4720,N_4685);
or U5019 (N_5019,N_4523,N_4601);
and U5020 (N_5020,N_4822,N_4879);
and U5021 (N_5021,N_4804,N_4981);
xor U5022 (N_5022,N_4847,N_4666);
nor U5023 (N_5023,N_4977,N_4948);
or U5024 (N_5024,N_4932,N_4975);
xor U5025 (N_5025,N_4660,N_4768);
nand U5026 (N_5026,N_4640,N_4818);
xor U5027 (N_5027,N_4584,N_4979);
xnor U5028 (N_5028,N_4592,N_4773);
xnor U5029 (N_5029,N_4928,N_4648);
nand U5030 (N_5030,N_4891,N_4792);
nor U5031 (N_5031,N_4689,N_4848);
and U5032 (N_5032,N_4626,N_4667);
and U5033 (N_5033,N_4500,N_4759);
nor U5034 (N_5034,N_4984,N_4968);
and U5035 (N_5035,N_4620,N_4945);
nor U5036 (N_5036,N_4650,N_4836);
nand U5037 (N_5037,N_4699,N_4549);
nand U5038 (N_5038,N_4908,N_4903);
nor U5039 (N_5039,N_4933,N_4535);
or U5040 (N_5040,N_4779,N_4559);
xnor U5041 (N_5041,N_4865,N_4834);
nand U5042 (N_5042,N_4766,N_4752);
and U5043 (N_5043,N_4639,N_4576);
nand U5044 (N_5044,N_4713,N_4817);
or U5045 (N_5045,N_4927,N_4955);
or U5046 (N_5046,N_4800,N_4950);
nor U5047 (N_5047,N_4596,N_4693);
and U5048 (N_5048,N_4655,N_4862);
nor U5049 (N_5049,N_4803,N_4514);
and U5050 (N_5050,N_4509,N_4993);
nand U5051 (N_5051,N_4816,N_4556);
or U5052 (N_5052,N_4548,N_4663);
or U5053 (N_5053,N_4574,N_4597);
or U5054 (N_5054,N_4854,N_4668);
and U5055 (N_5055,N_4569,N_4623);
xnor U5056 (N_5056,N_4838,N_4571);
and U5057 (N_5057,N_4538,N_4856);
nand U5058 (N_5058,N_4806,N_4906);
nor U5059 (N_5059,N_4555,N_4701);
xnor U5060 (N_5060,N_4839,N_4939);
or U5061 (N_5061,N_4990,N_4941);
and U5062 (N_5062,N_4832,N_4929);
xor U5063 (N_5063,N_4855,N_4815);
or U5064 (N_5064,N_4805,N_4557);
nand U5065 (N_5065,N_4777,N_4962);
and U5066 (N_5066,N_4624,N_4653);
and U5067 (N_5067,N_4649,N_4830);
nor U5068 (N_5068,N_4687,N_4723);
nand U5069 (N_5069,N_4565,N_4508);
nand U5070 (N_5070,N_4696,N_4673);
nand U5071 (N_5071,N_4905,N_4622);
xor U5072 (N_5072,N_4821,N_4618);
xor U5073 (N_5073,N_4645,N_4616);
xor U5074 (N_5074,N_4560,N_4543);
nor U5075 (N_5075,N_4705,N_4988);
or U5076 (N_5076,N_4845,N_4788);
xor U5077 (N_5077,N_4775,N_4769);
nand U5078 (N_5078,N_4878,N_4896);
or U5079 (N_5079,N_4913,N_4679);
xor U5080 (N_5080,N_4884,N_4613);
nand U5081 (N_5081,N_4674,N_4706);
nand U5082 (N_5082,N_4875,N_4860);
nand U5083 (N_5083,N_4629,N_4880);
nand U5084 (N_5084,N_4600,N_4553);
nor U5085 (N_5085,N_4558,N_4784);
nand U5086 (N_5086,N_4778,N_4973);
nor U5087 (N_5087,N_4582,N_4909);
nor U5088 (N_5088,N_4892,N_4749);
xnor U5089 (N_5089,N_4820,N_4529);
or U5090 (N_5090,N_4697,N_4946);
nor U5091 (N_5091,N_4810,N_4522);
nor U5092 (N_5092,N_4965,N_4811);
and U5093 (N_5093,N_4942,N_4641);
nand U5094 (N_5094,N_4943,N_4722);
xor U5095 (N_5095,N_4897,N_4552);
and U5096 (N_5096,N_4874,N_4665);
nand U5097 (N_5097,N_4873,N_4895);
nand U5098 (N_5098,N_4868,N_4935);
nand U5099 (N_5099,N_4900,N_4716);
nand U5100 (N_5100,N_4672,N_4694);
xnor U5101 (N_5101,N_4812,N_4835);
xor U5102 (N_5102,N_4586,N_4502);
and U5103 (N_5103,N_4888,N_4528);
and U5104 (N_5104,N_4846,N_4633);
nand U5105 (N_5105,N_4525,N_4515);
nor U5106 (N_5106,N_4670,N_4877);
nand U5107 (N_5107,N_4541,N_4849);
and U5108 (N_5108,N_4739,N_4572);
or U5109 (N_5109,N_4585,N_4999);
or U5110 (N_5110,N_4724,N_4774);
or U5111 (N_5111,N_4958,N_4504);
and U5112 (N_5112,N_4591,N_4910);
nand U5113 (N_5113,N_4954,N_4579);
and U5114 (N_5114,N_4748,N_4813);
or U5115 (N_5115,N_4707,N_4651);
and U5116 (N_5116,N_4914,N_4911);
and U5117 (N_5117,N_4513,N_4989);
nand U5118 (N_5118,N_4947,N_4700);
or U5119 (N_5119,N_4551,N_4826);
nand U5120 (N_5120,N_4869,N_4680);
nand U5121 (N_5121,N_4730,N_4704);
nand U5122 (N_5122,N_4683,N_4899);
or U5123 (N_5123,N_4539,N_4787);
or U5124 (N_5124,N_4533,N_4671);
and U5125 (N_5125,N_4505,N_4503);
xnor U5126 (N_5126,N_4636,N_4631);
or U5127 (N_5127,N_4758,N_4669);
and U5128 (N_5128,N_4681,N_4634);
nor U5129 (N_5129,N_4755,N_4844);
nand U5130 (N_5130,N_4644,N_4790);
nand U5131 (N_5131,N_4921,N_4767);
nand U5132 (N_5132,N_4986,N_4841);
nand U5133 (N_5133,N_4702,N_4991);
xor U5134 (N_5134,N_4791,N_4957);
xnor U5135 (N_5135,N_4537,N_4761);
nand U5136 (N_5136,N_4516,N_4536);
nand U5137 (N_5137,N_4887,N_4898);
xnor U5138 (N_5138,N_4708,N_4995);
or U5139 (N_5139,N_4610,N_4840);
or U5140 (N_5140,N_4594,N_4978);
nor U5141 (N_5141,N_4765,N_4859);
nand U5142 (N_5142,N_4886,N_4916);
xor U5143 (N_5143,N_4940,N_4587);
xor U5144 (N_5144,N_4870,N_4926);
xnor U5145 (N_5145,N_4581,N_4678);
xor U5146 (N_5146,N_4643,N_4562);
nor U5147 (N_5147,N_4617,N_4867);
or U5148 (N_5148,N_4686,N_4726);
xnor U5149 (N_5149,N_4823,N_4715);
xnor U5150 (N_5150,N_4744,N_4628);
and U5151 (N_5151,N_4692,N_4570);
or U5152 (N_5152,N_4656,N_4621);
nand U5153 (N_5153,N_4825,N_4843);
nand U5154 (N_5154,N_4980,N_4554);
nor U5155 (N_5155,N_4563,N_4662);
nor U5156 (N_5156,N_4785,N_4902);
or U5157 (N_5157,N_4519,N_4593);
xnor U5158 (N_5158,N_4881,N_4695);
xnor U5159 (N_5159,N_4719,N_4518);
nand U5160 (N_5160,N_4799,N_4918);
nand U5161 (N_5161,N_4863,N_4831);
xor U5162 (N_5162,N_4937,N_4544);
or U5163 (N_5163,N_4520,N_4770);
nor U5164 (N_5164,N_4737,N_4583);
nor U5165 (N_5165,N_4534,N_4953);
xnor U5166 (N_5166,N_4608,N_4746);
nor U5167 (N_5167,N_4998,N_4925);
nand U5168 (N_5168,N_4951,N_4819);
xor U5169 (N_5169,N_4959,N_4506);
nor U5170 (N_5170,N_4754,N_4550);
xor U5171 (N_5171,N_4691,N_4760);
and U5172 (N_5172,N_4732,N_4736);
and U5173 (N_5173,N_4966,N_4837);
xor U5174 (N_5174,N_4646,N_4976);
and U5175 (N_5175,N_4772,N_4642);
xor U5176 (N_5176,N_4956,N_4904);
or U5177 (N_5177,N_4923,N_4637);
nand U5178 (N_5178,N_4627,N_4580);
and U5179 (N_5179,N_4728,N_4611);
nor U5180 (N_5180,N_4657,N_4603);
xor U5181 (N_5181,N_4578,N_4824);
or U5182 (N_5182,N_4764,N_4564);
nand U5183 (N_5183,N_4793,N_4507);
nand U5184 (N_5184,N_4501,N_4964);
xor U5185 (N_5185,N_4912,N_4781);
xnor U5186 (N_5186,N_4721,N_4568);
or U5187 (N_5187,N_4717,N_4531);
and U5188 (N_5188,N_4776,N_4654);
nand U5189 (N_5189,N_4851,N_4725);
or U5190 (N_5190,N_4658,N_4738);
or U5191 (N_5191,N_4742,N_4794);
and U5192 (N_5192,N_4974,N_4567);
nand U5193 (N_5193,N_4606,N_4795);
or U5194 (N_5194,N_4698,N_4783);
or U5195 (N_5195,N_4652,N_4734);
nand U5196 (N_5196,N_4612,N_4740);
and U5197 (N_5197,N_4987,N_4588);
nand U5198 (N_5198,N_4526,N_4789);
or U5199 (N_5199,N_4960,N_4907);
or U5200 (N_5200,N_4915,N_4938);
nand U5201 (N_5201,N_4632,N_4970);
or U5202 (N_5202,N_4750,N_4972);
and U5203 (N_5203,N_4540,N_4690);
nor U5204 (N_5204,N_4573,N_4971);
and U5205 (N_5205,N_4602,N_4524);
xor U5206 (N_5206,N_4797,N_4532);
nor U5207 (N_5207,N_4614,N_4625);
nor U5208 (N_5208,N_4510,N_4590);
xor U5209 (N_5209,N_4883,N_4545);
or U5210 (N_5210,N_4967,N_4934);
and U5211 (N_5211,N_4688,N_4920);
xnor U5212 (N_5212,N_4684,N_4857);
nand U5213 (N_5213,N_4893,N_4703);
nor U5214 (N_5214,N_4630,N_4931);
xor U5215 (N_5215,N_4595,N_4889);
and U5216 (N_5216,N_4809,N_4852);
nand U5217 (N_5217,N_4802,N_4577);
or U5218 (N_5218,N_4963,N_4561);
and U5219 (N_5219,N_4885,N_4735);
nand U5220 (N_5220,N_4808,N_4517);
xor U5221 (N_5221,N_4677,N_4547);
nand U5222 (N_5222,N_4936,N_4605);
nand U5223 (N_5223,N_4753,N_4882);
or U5224 (N_5224,N_4827,N_4944);
nand U5225 (N_5225,N_4682,N_4712);
nand U5226 (N_5226,N_4894,N_4546);
xor U5227 (N_5227,N_4890,N_4661);
nor U5228 (N_5228,N_4756,N_4511);
nor U5229 (N_5229,N_4780,N_4961);
or U5230 (N_5230,N_4919,N_4607);
and U5231 (N_5231,N_4861,N_4743);
or U5232 (N_5232,N_4985,N_4757);
and U5233 (N_5233,N_4709,N_4762);
or U5234 (N_5234,N_4589,N_4512);
xor U5235 (N_5235,N_4924,N_4714);
nor U5236 (N_5236,N_4798,N_4619);
nor U5237 (N_5237,N_4982,N_4542);
or U5238 (N_5238,N_4949,N_4969);
and U5239 (N_5239,N_4872,N_4527);
and U5240 (N_5240,N_4635,N_4828);
and U5241 (N_5241,N_4609,N_4733);
nor U5242 (N_5242,N_4604,N_4718);
and U5243 (N_5243,N_4871,N_4994);
nand U5244 (N_5244,N_4842,N_4796);
or U5245 (N_5245,N_4850,N_4833);
xnor U5246 (N_5246,N_4801,N_4829);
nand U5247 (N_5247,N_4659,N_4747);
or U5248 (N_5248,N_4727,N_4729);
nor U5249 (N_5249,N_4675,N_4864);
and U5250 (N_5250,N_4580,N_4534);
and U5251 (N_5251,N_4617,N_4925);
or U5252 (N_5252,N_4925,N_4961);
and U5253 (N_5253,N_4677,N_4582);
nor U5254 (N_5254,N_4900,N_4595);
xor U5255 (N_5255,N_4831,N_4918);
and U5256 (N_5256,N_4865,N_4789);
xor U5257 (N_5257,N_4905,N_4790);
xnor U5258 (N_5258,N_4924,N_4585);
and U5259 (N_5259,N_4859,N_4658);
nor U5260 (N_5260,N_4712,N_4664);
xor U5261 (N_5261,N_4997,N_4845);
and U5262 (N_5262,N_4521,N_4865);
or U5263 (N_5263,N_4689,N_4969);
and U5264 (N_5264,N_4710,N_4655);
nand U5265 (N_5265,N_4716,N_4948);
and U5266 (N_5266,N_4714,N_4944);
nor U5267 (N_5267,N_4914,N_4730);
nor U5268 (N_5268,N_4710,N_4848);
nor U5269 (N_5269,N_4760,N_4949);
nor U5270 (N_5270,N_4811,N_4906);
xor U5271 (N_5271,N_4804,N_4843);
nor U5272 (N_5272,N_4668,N_4603);
xnor U5273 (N_5273,N_4808,N_4724);
nand U5274 (N_5274,N_4812,N_4846);
nand U5275 (N_5275,N_4634,N_4809);
nand U5276 (N_5276,N_4614,N_4988);
nand U5277 (N_5277,N_4800,N_4761);
and U5278 (N_5278,N_4609,N_4805);
xor U5279 (N_5279,N_4973,N_4529);
nor U5280 (N_5280,N_4820,N_4553);
xnor U5281 (N_5281,N_4639,N_4769);
nand U5282 (N_5282,N_4904,N_4639);
nand U5283 (N_5283,N_4572,N_4664);
or U5284 (N_5284,N_4651,N_4910);
or U5285 (N_5285,N_4837,N_4500);
xor U5286 (N_5286,N_4986,N_4669);
and U5287 (N_5287,N_4876,N_4753);
or U5288 (N_5288,N_4814,N_4504);
or U5289 (N_5289,N_4874,N_4832);
xor U5290 (N_5290,N_4828,N_4781);
xnor U5291 (N_5291,N_4537,N_4559);
nor U5292 (N_5292,N_4838,N_4863);
nand U5293 (N_5293,N_4836,N_4519);
or U5294 (N_5294,N_4598,N_4597);
and U5295 (N_5295,N_4652,N_4531);
nand U5296 (N_5296,N_4690,N_4849);
and U5297 (N_5297,N_4728,N_4953);
nand U5298 (N_5298,N_4893,N_4620);
and U5299 (N_5299,N_4658,N_4632);
xnor U5300 (N_5300,N_4934,N_4555);
or U5301 (N_5301,N_4909,N_4942);
or U5302 (N_5302,N_4966,N_4940);
xnor U5303 (N_5303,N_4505,N_4636);
or U5304 (N_5304,N_4942,N_4669);
nor U5305 (N_5305,N_4903,N_4501);
nor U5306 (N_5306,N_4666,N_4838);
xnor U5307 (N_5307,N_4618,N_4550);
xnor U5308 (N_5308,N_4919,N_4800);
and U5309 (N_5309,N_4557,N_4623);
nand U5310 (N_5310,N_4749,N_4980);
nor U5311 (N_5311,N_4805,N_4615);
nand U5312 (N_5312,N_4560,N_4737);
nand U5313 (N_5313,N_4765,N_4739);
xnor U5314 (N_5314,N_4883,N_4560);
xnor U5315 (N_5315,N_4795,N_4567);
nor U5316 (N_5316,N_4999,N_4574);
xnor U5317 (N_5317,N_4717,N_4629);
xor U5318 (N_5318,N_4957,N_4524);
nor U5319 (N_5319,N_4750,N_4619);
and U5320 (N_5320,N_4905,N_4828);
or U5321 (N_5321,N_4865,N_4997);
nand U5322 (N_5322,N_4794,N_4810);
xor U5323 (N_5323,N_4567,N_4662);
nand U5324 (N_5324,N_4661,N_4518);
or U5325 (N_5325,N_4563,N_4589);
nand U5326 (N_5326,N_4619,N_4739);
xnor U5327 (N_5327,N_4660,N_4504);
nor U5328 (N_5328,N_4856,N_4940);
xnor U5329 (N_5329,N_4522,N_4830);
nor U5330 (N_5330,N_4568,N_4817);
nand U5331 (N_5331,N_4831,N_4694);
xnor U5332 (N_5332,N_4954,N_4816);
and U5333 (N_5333,N_4932,N_4759);
xnor U5334 (N_5334,N_4635,N_4830);
nand U5335 (N_5335,N_4678,N_4536);
xnor U5336 (N_5336,N_4716,N_4586);
or U5337 (N_5337,N_4723,N_4729);
nor U5338 (N_5338,N_4554,N_4887);
and U5339 (N_5339,N_4866,N_4722);
or U5340 (N_5340,N_4516,N_4700);
and U5341 (N_5341,N_4779,N_4666);
nor U5342 (N_5342,N_4915,N_4881);
or U5343 (N_5343,N_4816,N_4723);
nor U5344 (N_5344,N_4835,N_4950);
nand U5345 (N_5345,N_4609,N_4512);
xor U5346 (N_5346,N_4801,N_4622);
nor U5347 (N_5347,N_4518,N_4881);
nor U5348 (N_5348,N_4534,N_4653);
xor U5349 (N_5349,N_4771,N_4984);
nor U5350 (N_5350,N_4557,N_4925);
and U5351 (N_5351,N_4960,N_4779);
xor U5352 (N_5352,N_4846,N_4667);
xor U5353 (N_5353,N_4755,N_4731);
xor U5354 (N_5354,N_4853,N_4844);
or U5355 (N_5355,N_4520,N_4901);
and U5356 (N_5356,N_4569,N_4651);
or U5357 (N_5357,N_4800,N_4638);
nand U5358 (N_5358,N_4549,N_4964);
or U5359 (N_5359,N_4651,N_4600);
and U5360 (N_5360,N_4768,N_4713);
nor U5361 (N_5361,N_4686,N_4799);
or U5362 (N_5362,N_4737,N_4880);
nor U5363 (N_5363,N_4502,N_4588);
nor U5364 (N_5364,N_4616,N_4577);
nor U5365 (N_5365,N_4793,N_4770);
or U5366 (N_5366,N_4853,N_4510);
nand U5367 (N_5367,N_4547,N_4801);
nor U5368 (N_5368,N_4931,N_4629);
nor U5369 (N_5369,N_4524,N_4605);
or U5370 (N_5370,N_4824,N_4675);
xnor U5371 (N_5371,N_4678,N_4731);
xor U5372 (N_5372,N_4515,N_4922);
nor U5373 (N_5373,N_4970,N_4565);
or U5374 (N_5374,N_4824,N_4944);
xor U5375 (N_5375,N_4787,N_4788);
or U5376 (N_5376,N_4679,N_4637);
nor U5377 (N_5377,N_4670,N_4564);
nor U5378 (N_5378,N_4944,N_4847);
and U5379 (N_5379,N_4650,N_4914);
nand U5380 (N_5380,N_4580,N_4866);
and U5381 (N_5381,N_4809,N_4739);
and U5382 (N_5382,N_4791,N_4866);
nand U5383 (N_5383,N_4917,N_4851);
nand U5384 (N_5384,N_4807,N_4644);
or U5385 (N_5385,N_4858,N_4638);
xor U5386 (N_5386,N_4906,N_4762);
xnor U5387 (N_5387,N_4721,N_4973);
nand U5388 (N_5388,N_4633,N_4863);
xor U5389 (N_5389,N_4976,N_4874);
xnor U5390 (N_5390,N_4986,N_4714);
xnor U5391 (N_5391,N_4693,N_4919);
nand U5392 (N_5392,N_4745,N_4820);
xor U5393 (N_5393,N_4810,N_4574);
nand U5394 (N_5394,N_4786,N_4775);
and U5395 (N_5395,N_4611,N_4634);
nand U5396 (N_5396,N_4799,N_4557);
xor U5397 (N_5397,N_4773,N_4885);
nor U5398 (N_5398,N_4988,N_4554);
xor U5399 (N_5399,N_4517,N_4880);
and U5400 (N_5400,N_4765,N_4587);
xnor U5401 (N_5401,N_4594,N_4512);
and U5402 (N_5402,N_4965,N_4555);
xnor U5403 (N_5403,N_4514,N_4659);
or U5404 (N_5404,N_4502,N_4988);
and U5405 (N_5405,N_4932,N_4831);
or U5406 (N_5406,N_4774,N_4909);
or U5407 (N_5407,N_4834,N_4816);
or U5408 (N_5408,N_4794,N_4741);
and U5409 (N_5409,N_4713,N_4910);
or U5410 (N_5410,N_4514,N_4737);
and U5411 (N_5411,N_4599,N_4726);
nor U5412 (N_5412,N_4738,N_4578);
xor U5413 (N_5413,N_4510,N_4635);
xor U5414 (N_5414,N_4580,N_4814);
nor U5415 (N_5415,N_4639,N_4795);
or U5416 (N_5416,N_4716,N_4877);
nor U5417 (N_5417,N_4917,N_4918);
nor U5418 (N_5418,N_4514,N_4931);
or U5419 (N_5419,N_4548,N_4510);
nor U5420 (N_5420,N_4536,N_4722);
and U5421 (N_5421,N_4645,N_4620);
or U5422 (N_5422,N_4719,N_4859);
nor U5423 (N_5423,N_4806,N_4776);
and U5424 (N_5424,N_4750,N_4561);
nor U5425 (N_5425,N_4971,N_4744);
nand U5426 (N_5426,N_4784,N_4516);
nor U5427 (N_5427,N_4729,N_4900);
xor U5428 (N_5428,N_4611,N_4738);
nand U5429 (N_5429,N_4754,N_4831);
nand U5430 (N_5430,N_4769,N_4618);
and U5431 (N_5431,N_4852,N_4859);
or U5432 (N_5432,N_4690,N_4796);
xor U5433 (N_5433,N_4572,N_4545);
or U5434 (N_5434,N_4863,N_4696);
xor U5435 (N_5435,N_4519,N_4755);
or U5436 (N_5436,N_4794,N_4912);
nor U5437 (N_5437,N_4931,N_4880);
and U5438 (N_5438,N_4902,N_4737);
and U5439 (N_5439,N_4535,N_4931);
or U5440 (N_5440,N_4702,N_4718);
nor U5441 (N_5441,N_4837,N_4667);
xor U5442 (N_5442,N_4643,N_4678);
nor U5443 (N_5443,N_4963,N_4637);
nor U5444 (N_5444,N_4501,N_4883);
nor U5445 (N_5445,N_4869,N_4988);
nor U5446 (N_5446,N_4896,N_4521);
nor U5447 (N_5447,N_4631,N_4649);
or U5448 (N_5448,N_4513,N_4549);
nor U5449 (N_5449,N_4884,N_4654);
or U5450 (N_5450,N_4647,N_4697);
or U5451 (N_5451,N_4555,N_4647);
nor U5452 (N_5452,N_4897,N_4648);
nor U5453 (N_5453,N_4603,N_4539);
or U5454 (N_5454,N_4838,N_4937);
nor U5455 (N_5455,N_4961,N_4860);
xnor U5456 (N_5456,N_4718,N_4757);
or U5457 (N_5457,N_4779,N_4809);
and U5458 (N_5458,N_4751,N_4970);
nand U5459 (N_5459,N_4653,N_4646);
nand U5460 (N_5460,N_4627,N_4624);
xor U5461 (N_5461,N_4529,N_4751);
nand U5462 (N_5462,N_4892,N_4970);
nor U5463 (N_5463,N_4912,N_4828);
or U5464 (N_5464,N_4957,N_4781);
nand U5465 (N_5465,N_4997,N_4807);
nand U5466 (N_5466,N_4585,N_4580);
xor U5467 (N_5467,N_4514,N_4982);
xor U5468 (N_5468,N_4599,N_4623);
nand U5469 (N_5469,N_4792,N_4884);
xor U5470 (N_5470,N_4876,N_4863);
nor U5471 (N_5471,N_4864,N_4603);
xor U5472 (N_5472,N_4743,N_4763);
or U5473 (N_5473,N_4744,N_4841);
or U5474 (N_5474,N_4529,N_4593);
nand U5475 (N_5475,N_4608,N_4753);
and U5476 (N_5476,N_4665,N_4574);
or U5477 (N_5477,N_4762,N_4543);
xnor U5478 (N_5478,N_4983,N_4520);
xnor U5479 (N_5479,N_4514,N_4562);
nor U5480 (N_5480,N_4996,N_4986);
xor U5481 (N_5481,N_4747,N_4752);
nand U5482 (N_5482,N_4510,N_4604);
nor U5483 (N_5483,N_4811,N_4870);
or U5484 (N_5484,N_4695,N_4831);
nand U5485 (N_5485,N_4729,N_4771);
and U5486 (N_5486,N_4570,N_4791);
nor U5487 (N_5487,N_4660,N_4630);
or U5488 (N_5488,N_4801,N_4845);
nor U5489 (N_5489,N_4993,N_4724);
nand U5490 (N_5490,N_4826,N_4713);
nand U5491 (N_5491,N_4731,N_4630);
nand U5492 (N_5492,N_4859,N_4830);
xor U5493 (N_5493,N_4543,N_4595);
nor U5494 (N_5494,N_4520,N_4603);
and U5495 (N_5495,N_4734,N_4950);
or U5496 (N_5496,N_4883,N_4807);
or U5497 (N_5497,N_4920,N_4916);
nor U5498 (N_5498,N_4858,N_4513);
or U5499 (N_5499,N_4781,N_4962);
or U5500 (N_5500,N_5318,N_5329);
or U5501 (N_5501,N_5001,N_5358);
nor U5502 (N_5502,N_5095,N_5474);
xnor U5503 (N_5503,N_5301,N_5108);
nand U5504 (N_5504,N_5186,N_5090);
xnor U5505 (N_5505,N_5400,N_5141);
xor U5506 (N_5506,N_5423,N_5128);
nand U5507 (N_5507,N_5196,N_5346);
nor U5508 (N_5508,N_5344,N_5359);
nor U5509 (N_5509,N_5305,N_5435);
xnor U5510 (N_5510,N_5410,N_5322);
or U5511 (N_5511,N_5323,N_5429);
nand U5512 (N_5512,N_5324,N_5038);
and U5513 (N_5513,N_5198,N_5216);
and U5514 (N_5514,N_5149,N_5334);
or U5515 (N_5515,N_5181,N_5194);
xor U5516 (N_5516,N_5471,N_5051);
nand U5517 (N_5517,N_5476,N_5013);
xnor U5518 (N_5518,N_5024,N_5176);
xor U5519 (N_5519,N_5117,N_5310);
or U5520 (N_5520,N_5279,N_5231);
nor U5521 (N_5521,N_5342,N_5010);
nand U5522 (N_5522,N_5477,N_5293);
or U5523 (N_5523,N_5247,N_5481);
and U5524 (N_5524,N_5367,N_5268);
nand U5525 (N_5525,N_5163,N_5138);
nand U5526 (N_5526,N_5100,N_5101);
xnor U5527 (N_5527,N_5497,N_5331);
xnor U5528 (N_5528,N_5345,N_5419);
and U5529 (N_5529,N_5294,N_5364);
and U5530 (N_5530,N_5219,N_5304);
nor U5531 (N_5531,N_5298,N_5485);
nand U5532 (N_5532,N_5234,N_5459);
or U5533 (N_5533,N_5143,N_5058);
nand U5534 (N_5534,N_5228,N_5411);
and U5535 (N_5535,N_5495,N_5416);
nand U5536 (N_5536,N_5157,N_5387);
and U5537 (N_5537,N_5059,N_5484);
xnor U5538 (N_5538,N_5487,N_5320);
nand U5539 (N_5539,N_5252,N_5492);
nand U5540 (N_5540,N_5458,N_5269);
nor U5541 (N_5541,N_5085,N_5054);
xor U5542 (N_5542,N_5473,N_5260);
or U5543 (N_5543,N_5285,N_5086);
and U5544 (N_5544,N_5472,N_5250);
nand U5545 (N_5545,N_5319,N_5347);
nor U5546 (N_5546,N_5061,N_5034);
and U5547 (N_5547,N_5026,N_5464);
nor U5548 (N_5548,N_5210,N_5389);
and U5549 (N_5549,N_5076,N_5047);
or U5550 (N_5550,N_5112,N_5192);
nand U5551 (N_5551,N_5457,N_5207);
and U5552 (N_5552,N_5378,N_5437);
nand U5553 (N_5553,N_5191,N_5494);
nor U5554 (N_5554,N_5355,N_5483);
nor U5555 (N_5555,N_5035,N_5016);
xor U5556 (N_5556,N_5152,N_5146);
xor U5557 (N_5557,N_5221,N_5154);
xnor U5558 (N_5558,N_5450,N_5273);
or U5559 (N_5559,N_5053,N_5111);
and U5560 (N_5560,N_5130,N_5027);
nand U5561 (N_5561,N_5466,N_5372);
nand U5562 (N_5562,N_5271,N_5362);
nand U5563 (N_5563,N_5140,N_5482);
or U5564 (N_5564,N_5277,N_5068);
and U5565 (N_5565,N_5498,N_5158);
xor U5566 (N_5566,N_5036,N_5037);
nand U5567 (N_5567,N_5244,N_5114);
or U5568 (N_5568,N_5230,N_5178);
or U5569 (N_5569,N_5469,N_5204);
nand U5570 (N_5570,N_5105,N_5166);
or U5571 (N_5571,N_5428,N_5071);
nor U5572 (N_5572,N_5360,N_5241);
or U5573 (N_5573,N_5262,N_5041);
and U5574 (N_5574,N_5297,N_5002);
nor U5575 (N_5575,N_5239,N_5353);
and U5576 (N_5576,N_5099,N_5020);
or U5577 (N_5577,N_5448,N_5087);
and U5578 (N_5578,N_5119,N_5357);
and U5579 (N_5579,N_5052,N_5170);
or U5580 (N_5580,N_5415,N_5371);
nand U5581 (N_5581,N_5017,N_5098);
and U5582 (N_5582,N_5366,N_5296);
xor U5583 (N_5583,N_5102,N_5172);
nor U5584 (N_5584,N_5151,N_5461);
xnor U5585 (N_5585,N_5491,N_5070);
nand U5586 (N_5586,N_5409,N_5067);
nor U5587 (N_5587,N_5229,N_5451);
and U5588 (N_5588,N_5201,N_5454);
or U5589 (N_5589,N_5093,N_5225);
and U5590 (N_5590,N_5384,N_5218);
or U5591 (N_5591,N_5327,N_5083);
xor U5592 (N_5592,N_5200,N_5365);
nand U5593 (N_5593,N_5049,N_5385);
nand U5594 (N_5594,N_5177,N_5044);
and U5595 (N_5595,N_5233,N_5014);
or U5596 (N_5596,N_5243,N_5350);
xnor U5597 (N_5597,N_5179,N_5309);
and U5598 (N_5598,N_5321,N_5394);
nand U5599 (N_5599,N_5422,N_5197);
nor U5600 (N_5600,N_5110,N_5470);
nand U5601 (N_5601,N_5300,N_5183);
nor U5602 (N_5602,N_5169,N_5092);
or U5603 (N_5603,N_5155,N_5008);
xor U5604 (N_5604,N_5258,N_5121);
or U5605 (N_5605,N_5281,N_5325);
or U5606 (N_5606,N_5316,N_5440);
nand U5607 (N_5607,N_5261,N_5145);
or U5608 (N_5608,N_5425,N_5465);
or U5609 (N_5609,N_5137,N_5391);
and U5610 (N_5610,N_5289,N_5238);
and U5611 (N_5611,N_5264,N_5308);
xnor U5612 (N_5612,N_5460,N_5147);
or U5613 (N_5613,N_5493,N_5392);
nand U5614 (N_5614,N_5403,N_5224);
or U5615 (N_5615,N_5453,N_5025);
nand U5616 (N_5616,N_5265,N_5184);
nand U5617 (N_5617,N_5259,N_5430);
and U5618 (N_5618,N_5286,N_5267);
nor U5619 (N_5619,N_5215,N_5232);
xor U5620 (N_5620,N_5307,N_5404);
nand U5621 (N_5621,N_5337,N_5222);
and U5622 (N_5622,N_5480,N_5284);
nor U5623 (N_5623,N_5467,N_5116);
nor U5624 (N_5624,N_5018,N_5131);
xnor U5625 (N_5625,N_5383,N_5205);
nand U5626 (N_5626,N_5190,N_5187);
and U5627 (N_5627,N_5275,N_5432);
xor U5628 (N_5628,N_5490,N_5213);
and U5629 (N_5629,N_5336,N_5062);
nand U5630 (N_5630,N_5007,N_5381);
xnor U5631 (N_5631,N_5040,N_5153);
nor U5632 (N_5632,N_5174,N_5256);
or U5633 (N_5633,N_5439,N_5188);
and U5634 (N_5634,N_5019,N_5468);
or U5635 (N_5635,N_5332,N_5314);
and U5636 (N_5636,N_5374,N_5072);
or U5637 (N_5637,N_5398,N_5287);
nor U5638 (N_5638,N_5081,N_5349);
and U5639 (N_5639,N_5000,N_5343);
and U5640 (N_5640,N_5414,N_5074);
or U5641 (N_5641,N_5015,N_5499);
nor U5642 (N_5642,N_5106,N_5050);
and U5643 (N_5643,N_5164,N_5436);
xor U5644 (N_5644,N_5148,N_5280);
nand U5645 (N_5645,N_5063,N_5254);
nor U5646 (N_5646,N_5202,N_5444);
nor U5647 (N_5647,N_5441,N_5122);
nand U5648 (N_5648,N_5126,N_5255);
xor U5649 (N_5649,N_5447,N_5139);
and U5650 (N_5650,N_5113,N_5235);
and U5651 (N_5651,N_5212,N_5171);
or U5652 (N_5652,N_5055,N_5412);
and U5653 (N_5653,N_5132,N_5033);
and U5654 (N_5654,N_5159,N_5368);
nor U5655 (N_5655,N_5393,N_5452);
nand U5656 (N_5656,N_5402,N_5245);
nand U5657 (N_5657,N_5042,N_5333);
nor U5658 (N_5658,N_5237,N_5388);
nand U5659 (N_5659,N_5283,N_5405);
xnor U5660 (N_5660,N_5421,N_5115);
and U5661 (N_5661,N_5442,N_5125);
xnor U5662 (N_5662,N_5278,N_5475);
xor U5663 (N_5663,N_5312,N_5227);
nor U5664 (N_5664,N_5124,N_5397);
nor U5665 (N_5665,N_5065,N_5375);
nand U5666 (N_5666,N_5352,N_5189);
nand U5667 (N_5667,N_5206,N_5377);
nand U5668 (N_5668,N_5299,N_5236);
nor U5669 (N_5669,N_5379,N_5288);
nand U5670 (N_5670,N_5031,N_5407);
or U5671 (N_5671,N_5274,N_5136);
or U5672 (N_5672,N_5445,N_5315);
xnor U5673 (N_5673,N_5091,N_5496);
or U5674 (N_5674,N_5479,N_5162);
nor U5675 (N_5675,N_5069,N_5079);
or U5676 (N_5676,N_5246,N_5376);
xnor U5677 (N_5677,N_5438,N_5075);
and U5678 (N_5678,N_5348,N_5144);
xor U5679 (N_5679,N_5182,N_5449);
xor U5680 (N_5680,N_5317,N_5168);
or U5681 (N_5681,N_5340,N_5313);
and U5682 (N_5682,N_5380,N_5003);
and U5683 (N_5683,N_5276,N_5488);
xor U5684 (N_5684,N_5096,N_5351);
xor U5685 (N_5685,N_5330,N_5030);
xnor U5686 (N_5686,N_5328,N_5272);
nor U5687 (N_5687,N_5386,N_5226);
or U5688 (N_5688,N_5150,N_5193);
and U5689 (N_5689,N_5434,N_5057);
nor U5690 (N_5690,N_5489,N_5303);
xnor U5691 (N_5691,N_5046,N_5180);
nand U5692 (N_5692,N_5039,N_5291);
and U5693 (N_5693,N_5433,N_5413);
xor U5694 (N_5694,N_5064,N_5311);
xor U5695 (N_5695,N_5089,N_5104);
or U5696 (N_5696,N_5107,N_5290);
and U5697 (N_5697,N_5199,N_5292);
xor U5698 (N_5698,N_5456,N_5142);
nor U5699 (N_5699,N_5045,N_5011);
and U5700 (N_5700,N_5338,N_5354);
xor U5701 (N_5701,N_5257,N_5208);
xor U5702 (N_5702,N_5424,N_5134);
xnor U5703 (N_5703,N_5161,N_5195);
or U5704 (N_5704,N_5478,N_5363);
and U5705 (N_5705,N_5427,N_5373);
nor U5706 (N_5706,N_5418,N_5399);
xnor U5707 (N_5707,N_5080,N_5006);
nand U5708 (N_5708,N_5094,N_5266);
xor U5709 (N_5709,N_5078,N_5023);
nor U5710 (N_5710,N_5302,N_5443);
and U5711 (N_5711,N_5408,N_5251);
nor U5712 (N_5712,N_5211,N_5248);
xnor U5713 (N_5713,N_5431,N_5361);
nor U5714 (N_5714,N_5048,N_5009);
xnor U5715 (N_5715,N_5133,N_5295);
nand U5716 (N_5716,N_5109,N_5446);
nand U5717 (N_5717,N_5217,N_5462);
and U5718 (N_5718,N_5056,N_5043);
xor U5719 (N_5719,N_5463,N_5214);
xor U5720 (N_5720,N_5396,N_5077);
xnor U5721 (N_5721,N_5209,N_5253);
or U5722 (N_5722,N_5066,N_5082);
nor U5723 (N_5723,N_5084,N_5203);
and U5724 (N_5724,N_5012,N_5406);
nand U5725 (N_5725,N_5401,N_5135);
and U5726 (N_5726,N_5240,N_5326);
and U5727 (N_5727,N_5088,N_5029);
xnor U5728 (N_5728,N_5120,N_5185);
nor U5729 (N_5729,N_5073,N_5223);
nor U5730 (N_5730,N_5426,N_5242);
and U5731 (N_5731,N_5060,N_5021);
or U5732 (N_5732,N_5028,N_5165);
xnor U5733 (N_5733,N_5335,N_5123);
nor U5734 (N_5734,N_5167,N_5118);
xnor U5735 (N_5735,N_5341,N_5420);
and U5736 (N_5736,N_5220,N_5249);
xor U5737 (N_5737,N_5455,N_5382);
nor U5738 (N_5738,N_5097,N_5173);
and U5739 (N_5739,N_5486,N_5004);
nor U5740 (N_5740,N_5175,N_5417);
and U5741 (N_5741,N_5156,N_5129);
nand U5742 (N_5742,N_5370,N_5103);
xnor U5743 (N_5743,N_5270,N_5127);
or U5744 (N_5744,N_5005,N_5263);
and U5745 (N_5745,N_5356,N_5022);
nand U5746 (N_5746,N_5395,N_5306);
nand U5747 (N_5747,N_5339,N_5160);
nand U5748 (N_5748,N_5282,N_5032);
or U5749 (N_5749,N_5369,N_5390);
or U5750 (N_5750,N_5022,N_5280);
or U5751 (N_5751,N_5328,N_5018);
nand U5752 (N_5752,N_5411,N_5045);
nand U5753 (N_5753,N_5322,N_5345);
nor U5754 (N_5754,N_5044,N_5224);
or U5755 (N_5755,N_5116,N_5027);
xnor U5756 (N_5756,N_5261,N_5378);
xor U5757 (N_5757,N_5275,N_5499);
nor U5758 (N_5758,N_5309,N_5015);
nand U5759 (N_5759,N_5285,N_5462);
or U5760 (N_5760,N_5151,N_5268);
nor U5761 (N_5761,N_5200,N_5266);
nor U5762 (N_5762,N_5020,N_5291);
and U5763 (N_5763,N_5381,N_5259);
or U5764 (N_5764,N_5448,N_5034);
nand U5765 (N_5765,N_5179,N_5463);
or U5766 (N_5766,N_5082,N_5052);
nand U5767 (N_5767,N_5276,N_5056);
xnor U5768 (N_5768,N_5469,N_5392);
and U5769 (N_5769,N_5477,N_5058);
and U5770 (N_5770,N_5034,N_5081);
nor U5771 (N_5771,N_5062,N_5210);
or U5772 (N_5772,N_5219,N_5073);
nand U5773 (N_5773,N_5048,N_5371);
xnor U5774 (N_5774,N_5266,N_5299);
xnor U5775 (N_5775,N_5213,N_5246);
and U5776 (N_5776,N_5100,N_5256);
nor U5777 (N_5777,N_5084,N_5224);
or U5778 (N_5778,N_5134,N_5195);
nor U5779 (N_5779,N_5165,N_5046);
nor U5780 (N_5780,N_5032,N_5378);
nor U5781 (N_5781,N_5347,N_5218);
and U5782 (N_5782,N_5428,N_5310);
nor U5783 (N_5783,N_5109,N_5200);
xnor U5784 (N_5784,N_5443,N_5366);
xor U5785 (N_5785,N_5148,N_5045);
nor U5786 (N_5786,N_5410,N_5300);
nor U5787 (N_5787,N_5211,N_5408);
nor U5788 (N_5788,N_5122,N_5464);
nand U5789 (N_5789,N_5009,N_5107);
or U5790 (N_5790,N_5412,N_5292);
or U5791 (N_5791,N_5353,N_5210);
nor U5792 (N_5792,N_5349,N_5418);
and U5793 (N_5793,N_5266,N_5171);
or U5794 (N_5794,N_5008,N_5018);
nand U5795 (N_5795,N_5068,N_5480);
or U5796 (N_5796,N_5494,N_5416);
and U5797 (N_5797,N_5015,N_5360);
and U5798 (N_5798,N_5169,N_5413);
nand U5799 (N_5799,N_5282,N_5457);
nor U5800 (N_5800,N_5179,N_5491);
nor U5801 (N_5801,N_5441,N_5245);
nor U5802 (N_5802,N_5431,N_5237);
nor U5803 (N_5803,N_5386,N_5348);
or U5804 (N_5804,N_5312,N_5147);
or U5805 (N_5805,N_5230,N_5383);
xnor U5806 (N_5806,N_5373,N_5269);
xor U5807 (N_5807,N_5438,N_5092);
xor U5808 (N_5808,N_5115,N_5034);
or U5809 (N_5809,N_5070,N_5003);
and U5810 (N_5810,N_5394,N_5492);
and U5811 (N_5811,N_5006,N_5460);
xnor U5812 (N_5812,N_5329,N_5403);
or U5813 (N_5813,N_5270,N_5455);
nand U5814 (N_5814,N_5045,N_5214);
xor U5815 (N_5815,N_5119,N_5138);
nand U5816 (N_5816,N_5157,N_5329);
nand U5817 (N_5817,N_5475,N_5352);
nor U5818 (N_5818,N_5165,N_5111);
xnor U5819 (N_5819,N_5027,N_5457);
or U5820 (N_5820,N_5477,N_5014);
nor U5821 (N_5821,N_5478,N_5154);
nand U5822 (N_5822,N_5470,N_5261);
nand U5823 (N_5823,N_5069,N_5373);
nor U5824 (N_5824,N_5272,N_5348);
nand U5825 (N_5825,N_5316,N_5254);
nand U5826 (N_5826,N_5341,N_5223);
or U5827 (N_5827,N_5452,N_5013);
nand U5828 (N_5828,N_5499,N_5130);
xnor U5829 (N_5829,N_5226,N_5456);
or U5830 (N_5830,N_5143,N_5481);
xor U5831 (N_5831,N_5279,N_5392);
nand U5832 (N_5832,N_5159,N_5093);
nor U5833 (N_5833,N_5058,N_5353);
nand U5834 (N_5834,N_5072,N_5377);
nand U5835 (N_5835,N_5298,N_5141);
or U5836 (N_5836,N_5373,N_5027);
and U5837 (N_5837,N_5158,N_5169);
nand U5838 (N_5838,N_5313,N_5461);
or U5839 (N_5839,N_5264,N_5206);
nand U5840 (N_5840,N_5444,N_5273);
or U5841 (N_5841,N_5483,N_5271);
nor U5842 (N_5842,N_5095,N_5357);
or U5843 (N_5843,N_5034,N_5177);
nand U5844 (N_5844,N_5340,N_5118);
or U5845 (N_5845,N_5189,N_5019);
nor U5846 (N_5846,N_5151,N_5221);
and U5847 (N_5847,N_5133,N_5411);
nand U5848 (N_5848,N_5179,N_5213);
or U5849 (N_5849,N_5219,N_5228);
nand U5850 (N_5850,N_5279,N_5165);
or U5851 (N_5851,N_5127,N_5323);
nor U5852 (N_5852,N_5327,N_5168);
nand U5853 (N_5853,N_5037,N_5195);
and U5854 (N_5854,N_5021,N_5123);
xnor U5855 (N_5855,N_5336,N_5446);
or U5856 (N_5856,N_5464,N_5462);
and U5857 (N_5857,N_5042,N_5270);
or U5858 (N_5858,N_5201,N_5191);
or U5859 (N_5859,N_5062,N_5129);
xor U5860 (N_5860,N_5107,N_5209);
and U5861 (N_5861,N_5403,N_5005);
nor U5862 (N_5862,N_5086,N_5118);
or U5863 (N_5863,N_5167,N_5274);
xor U5864 (N_5864,N_5058,N_5398);
nor U5865 (N_5865,N_5225,N_5198);
xor U5866 (N_5866,N_5127,N_5420);
xnor U5867 (N_5867,N_5462,N_5475);
and U5868 (N_5868,N_5144,N_5487);
nand U5869 (N_5869,N_5012,N_5352);
nand U5870 (N_5870,N_5111,N_5064);
xnor U5871 (N_5871,N_5379,N_5069);
or U5872 (N_5872,N_5415,N_5423);
nand U5873 (N_5873,N_5061,N_5420);
nor U5874 (N_5874,N_5434,N_5225);
or U5875 (N_5875,N_5300,N_5145);
xnor U5876 (N_5876,N_5056,N_5117);
and U5877 (N_5877,N_5029,N_5177);
xor U5878 (N_5878,N_5219,N_5176);
xnor U5879 (N_5879,N_5346,N_5084);
xor U5880 (N_5880,N_5262,N_5187);
xnor U5881 (N_5881,N_5416,N_5442);
or U5882 (N_5882,N_5369,N_5231);
xnor U5883 (N_5883,N_5403,N_5239);
and U5884 (N_5884,N_5003,N_5390);
or U5885 (N_5885,N_5032,N_5125);
xnor U5886 (N_5886,N_5469,N_5497);
nand U5887 (N_5887,N_5436,N_5029);
and U5888 (N_5888,N_5495,N_5246);
or U5889 (N_5889,N_5391,N_5181);
or U5890 (N_5890,N_5080,N_5040);
nor U5891 (N_5891,N_5291,N_5224);
or U5892 (N_5892,N_5267,N_5006);
nand U5893 (N_5893,N_5486,N_5288);
nor U5894 (N_5894,N_5199,N_5202);
nor U5895 (N_5895,N_5056,N_5159);
and U5896 (N_5896,N_5355,N_5024);
and U5897 (N_5897,N_5059,N_5459);
and U5898 (N_5898,N_5331,N_5465);
xor U5899 (N_5899,N_5320,N_5400);
nor U5900 (N_5900,N_5271,N_5377);
and U5901 (N_5901,N_5433,N_5087);
nor U5902 (N_5902,N_5343,N_5227);
or U5903 (N_5903,N_5296,N_5093);
or U5904 (N_5904,N_5272,N_5259);
nor U5905 (N_5905,N_5034,N_5168);
or U5906 (N_5906,N_5059,N_5417);
xor U5907 (N_5907,N_5223,N_5428);
xnor U5908 (N_5908,N_5336,N_5049);
and U5909 (N_5909,N_5386,N_5097);
or U5910 (N_5910,N_5215,N_5043);
xor U5911 (N_5911,N_5339,N_5064);
nor U5912 (N_5912,N_5397,N_5009);
or U5913 (N_5913,N_5487,N_5449);
xor U5914 (N_5914,N_5130,N_5361);
and U5915 (N_5915,N_5036,N_5484);
or U5916 (N_5916,N_5402,N_5237);
nand U5917 (N_5917,N_5300,N_5330);
nand U5918 (N_5918,N_5210,N_5366);
and U5919 (N_5919,N_5154,N_5355);
nor U5920 (N_5920,N_5019,N_5161);
or U5921 (N_5921,N_5448,N_5352);
nand U5922 (N_5922,N_5318,N_5036);
and U5923 (N_5923,N_5338,N_5399);
nor U5924 (N_5924,N_5120,N_5380);
xnor U5925 (N_5925,N_5456,N_5293);
xnor U5926 (N_5926,N_5147,N_5065);
nand U5927 (N_5927,N_5054,N_5159);
nand U5928 (N_5928,N_5011,N_5112);
xnor U5929 (N_5929,N_5134,N_5451);
or U5930 (N_5930,N_5209,N_5290);
or U5931 (N_5931,N_5317,N_5447);
xor U5932 (N_5932,N_5256,N_5110);
xor U5933 (N_5933,N_5359,N_5355);
xor U5934 (N_5934,N_5393,N_5160);
xnor U5935 (N_5935,N_5169,N_5017);
or U5936 (N_5936,N_5102,N_5262);
or U5937 (N_5937,N_5250,N_5029);
nand U5938 (N_5938,N_5018,N_5191);
or U5939 (N_5939,N_5428,N_5080);
and U5940 (N_5940,N_5059,N_5106);
nand U5941 (N_5941,N_5183,N_5000);
or U5942 (N_5942,N_5400,N_5107);
nor U5943 (N_5943,N_5044,N_5293);
nor U5944 (N_5944,N_5080,N_5201);
xnor U5945 (N_5945,N_5441,N_5430);
or U5946 (N_5946,N_5182,N_5330);
xnor U5947 (N_5947,N_5430,N_5074);
nor U5948 (N_5948,N_5421,N_5300);
xnor U5949 (N_5949,N_5383,N_5197);
nand U5950 (N_5950,N_5336,N_5063);
and U5951 (N_5951,N_5445,N_5125);
or U5952 (N_5952,N_5269,N_5023);
and U5953 (N_5953,N_5398,N_5069);
or U5954 (N_5954,N_5216,N_5156);
nand U5955 (N_5955,N_5167,N_5223);
nor U5956 (N_5956,N_5325,N_5499);
nor U5957 (N_5957,N_5087,N_5005);
or U5958 (N_5958,N_5201,N_5341);
xnor U5959 (N_5959,N_5164,N_5439);
and U5960 (N_5960,N_5389,N_5264);
and U5961 (N_5961,N_5143,N_5360);
nor U5962 (N_5962,N_5122,N_5092);
and U5963 (N_5963,N_5196,N_5354);
and U5964 (N_5964,N_5487,N_5475);
and U5965 (N_5965,N_5420,N_5462);
and U5966 (N_5966,N_5046,N_5096);
nand U5967 (N_5967,N_5159,N_5334);
or U5968 (N_5968,N_5327,N_5258);
or U5969 (N_5969,N_5233,N_5108);
or U5970 (N_5970,N_5465,N_5052);
or U5971 (N_5971,N_5237,N_5494);
nor U5972 (N_5972,N_5364,N_5300);
nand U5973 (N_5973,N_5434,N_5142);
and U5974 (N_5974,N_5195,N_5326);
nand U5975 (N_5975,N_5304,N_5399);
xor U5976 (N_5976,N_5463,N_5291);
nor U5977 (N_5977,N_5332,N_5031);
nor U5978 (N_5978,N_5378,N_5198);
xor U5979 (N_5979,N_5406,N_5051);
xor U5980 (N_5980,N_5178,N_5135);
nand U5981 (N_5981,N_5004,N_5200);
nand U5982 (N_5982,N_5224,N_5120);
and U5983 (N_5983,N_5034,N_5295);
nand U5984 (N_5984,N_5351,N_5225);
nand U5985 (N_5985,N_5008,N_5225);
xor U5986 (N_5986,N_5311,N_5357);
nor U5987 (N_5987,N_5019,N_5094);
nand U5988 (N_5988,N_5323,N_5241);
or U5989 (N_5989,N_5145,N_5125);
nor U5990 (N_5990,N_5219,N_5243);
nand U5991 (N_5991,N_5480,N_5223);
and U5992 (N_5992,N_5304,N_5130);
or U5993 (N_5993,N_5443,N_5435);
xnor U5994 (N_5994,N_5483,N_5408);
nor U5995 (N_5995,N_5379,N_5167);
and U5996 (N_5996,N_5382,N_5200);
and U5997 (N_5997,N_5024,N_5059);
nand U5998 (N_5998,N_5287,N_5442);
and U5999 (N_5999,N_5232,N_5463);
nand U6000 (N_6000,N_5867,N_5937);
or U6001 (N_6001,N_5744,N_5992);
or U6002 (N_6002,N_5637,N_5971);
xnor U6003 (N_6003,N_5845,N_5524);
xor U6004 (N_6004,N_5757,N_5903);
and U6005 (N_6005,N_5751,N_5513);
or U6006 (N_6006,N_5802,N_5516);
nor U6007 (N_6007,N_5856,N_5866);
or U6008 (N_6008,N_5558,N_5548);
and U6009 (N_6009,N_5763,N_5719);
xnor U6010 (N_6010,N_5964,N_5860);
nand U6011 (N_6011,N_5805,N_5822);
nor U6012 (N_6012,N_5922,N_5855);
nand U6013 (N_6013,N_5512,N_5790);
nor U6014 (N_6014,N_5827,N_5576);
and U6015 (N_6015,N_5655,N_5733);
nand U6016 (N_6016,N_5673,N_5557);
nand U6017 (N_6017,N_5969,N_5975);
nand U6018 (N_6018,N_5534,N_5962);
or U6019 (N_6019,N_5646,N_5839);
xor U6020 (N_6020,N_5919,N_5675);
nor U6021 (N_6021,N_5585,N_5741);
and U6022 (N_6022,N_5792,N_5888);
nor U6023 (N_6023,N_5837,N_5911);
xnor U6024 (N_6024,N_5989,N_5955);
nand U6025 (N_6025,N_5899,N_5731);
xnor U6026 (N_6026,N_5796,N_5862);
xor U6027 (N_6027,N_5959,N_5926);
nand U6028 (N_6028,N_5671,N_5957);
xor U6029 (N_6029,N_5565,N_5521);
nor U6030 (N_6030,N_5659,N_5536);
and U6031 (N_6031,N_5775,N_5873);
nand U6032 (N_6032,N_5658,N_5972);
nor U6033 (N_6033,N_5892,N_5639);
xor U6034 (N_6034,N_5567,N_5766);
or U6035 (N_6035,N_5603,N_5774);
xor U6036 (N_6036,N_5853,N_5600);
and U6037 (N_6037,N_5615,N_5875);
nand U6038 (N_6038,N_5586,N_5609);
xor U6039 (N_6039,N_5829,N_5927);
nand U6040 (N_6040,N_5864,N_5891);
or U6041 (N_6041,N_5677,N_5712);
xnor U6042 (N_6042,N_5840,N_5706);
and U6043 (N_6043,N_5782,N_5676);
nand U6044 (N_6044,N_5778,N_5771);
and U6045 (N_6045,N_5504,N_5532);
or U6046 (N_6046,N_5691,N_5824);
nor U6047 (N_6047,N_5571,N_5589);
nand U6048 (N_6048,N_5803,N_5939);
nand U6049 (N_6049,N_5551,N_5643);
and U6050 (N_6050,N_5921,N_5721);
xor U6051 (N_6051,N_5880,N_5747);
xor U6052 (N_6052,N_5756,N_5727);
and U6053 (N_6053,N_5941,N_5627);
xnor U6054 (N_6054,N_5714,N_5813);
xnor U6055 (N_6055,N_5895,N_5750);
xor U6056 (N_6056,N_5893,N_5647);
or U6057 (N_6057,N_5711,N_5811);
and U6058 (N_6058,N_5987,N_5527);
and U6059 (N_6059,N_5525,N_5529);
and U6060 (N_6060,N_5681,N_5680);
nor U6061 (N_6061,N_5518,N_5799);
and U6062 (N_6062,N_5610,N_5550);
xnor U6063 (N_6063,N_5695,N_5631);
or U6064 (N_6064,N_5979,N_5848);
and U6065 (N_6065,N_5765,N_5668);
xnor U6066 (N_6066,N_5966,N_5601);
or U6067 (N_6067,N_5844,N_5906);
or U6068 (N_6068,N_5735,N_5816);
nand U6069 (N_6069,N_5530,N_5509);
or U6070 (N_6070,N_5692,N_5519);
xnor U6071 (N_6071,N_5849,N_5732);
or U6072 (N_6072,N_5670,N_5683);
or U6073 (N_6073,N_5907,N_5889);
nor U6074 (N_6074,N_5687,N_5597);
nor U6075 (N_6075,N_5770,N_5996);
nor U6076 (N_6076,N_5815,N_5549);
or U6077 (N_6077,N_5638,N_5632);
nor U6078 (N_6078,N_5842,N_5555);
or U6079 (N_6079,N_5994,N_5515);
nor U6080 (N_6080,N_5923,N_5838);
or U6081 (N_6081,N_5868,N_5858);
nor U6082 (N_6082,N_5630,N_5985);
or U6083 (N_6083,N_5833,N_5517);
xnor U6084 (N_6084,N_5781,N_5577);
nand U6085 (N_6085,N_5700,N_5915);
nand U6086 (N_6086,N_5871,N_5737);
nand U6087 (N_6087,N_5722,N_5968);
xor U6088 (N_6088,N_5898,N_5602);
and U6089 (N_6089,N_5552,N_5584);
nand U6090 (N_6090,N_5993,N_5894);
nand U6091 (N_6091,N_5566,N_5901);
or U6092 (N_6092,N_5946,N_5505);
nor U6093 (N_6093,N_5934,N_5544);
and U6094 (N_6094,N_5931,N_5999);
or U6095 (N_6095,N_5531,N_5890);
nand U6096 (N_6096,N_5980,N_5575);
or U6097 (N_6097,N_5773,N_5779);
nand U6098 (N_6098,N_5510,N_5794);
xor U6099 (N_6099,N_5896,N_5948);
xnor U6100 (N_6100,N_5641,N_5562);
or U6101 (N_6101,N_5990,N_5686);
nor U6102 (N_6102,N_5720,N_5857);
nand U6103 (N_6103,N_5998,N_5672);
nand U6104 (N_6104,N_5876,N_5715);
or U6105 (N_6105,N_5607,N_5960);
nand U6106 (N_6106,N_5910,N_5900);
nor U6107 (N_6107,N_5591,N_5956);
nor U6108 (N_6108,N_5523,N_5682);
and U6109 (N_6109,N_5596,N_5707);
or U6110 (N_6110,N_5593,N_5769);
nor U6111 (N_6111,N_5924,N_5705);
xor U6112 (N_6112,N_5717,N_5913);
and U6113 (N_6113,N_5791,N_5991);
or U6114 (N_6114,N_5788,N_5661);
nor U6115 (N_6115,N_5984,N_5718);
nor U6116 (N_6116,N_5635,N_5541);
or U6117 (N_6117,N_5592,N_5743);
nor U6118 (N_6118,N_5808,N_5928);
nand U6119 (N_6119,N_5854,N_5877);
nand U6120 (N_6120,N_5863,N_5563);
nor U6121 (N_6121,N_5542,N_5800);
xor U6122 (N_6122,N_5954,N_5869);
and U6123 (N_6123,N_5986,N_5826);
nor U6124 (N_6124,N_5657,N_5623);
nor U6125 (N_6125,N_5634,N_5832);
nand U6126 (N_6126,N_5724,N_5768);
nor U6127 (N_6127,N_5745,N_5932);
nor U6128 (N_6128,N_5553,N_5581);
or U6129 (N_6129,N_5787,N_5614);
and U6130 (N_6130,N_5943,N_5570);
or U6131 (N_6131,N_5502,N_5633);
and U6132 (N_6132,N_5636,N_5983);
xnor U6133 (N_6133,N_5936,N_5704);
nor U6134 (N_6134,N_5974,N_5713);
and U6135 (N_6135,N_5755,N_5678);
nor U6136 (N_6136,N_5949,N_5716);
or U6137 (N_6137,N_5749,N_5604);
and U6138 (N_6138,N_5746,N_5859);
nor U6139 (N_6139,N_5538,N_5789);
and U6140 (N_6140,N_5835,N_5754);
and U6141 (N_6141,N_5807,N_5709);
or U6142 (N_6142,N_5825,N_5688);
xnor U6143 (N_6143,N_5540,N_5830);
or U6144 (N_6144,N_5560,N_5736);
xor U6145 (N_6145,N_5967,N_5865);
xnor U6146 (N_6146,N_5660,N_5605);
and U6147 (N_6147,N_5621,N_5649);
nand U6148 (N_6148,N_5995,N_5801);
and U6149 (N_6149,N_5651,N_5951);
and U6150 (N_6150,N_5693,N_5702);
nand U6151 (N_6151,N_5982,N_5694);
nor U6152 (N_6152,N_5606,N_5664);
nor U6153 (N_6153,N_5819,N_5624);
nor U6154 (N_6154,N_5760,N_5587);
nor U6155 (N_6155,N_5574,N_5797);
nand U6156 (N_6156,N_5942,N_5742);
xnor U6157 (N_6157,N_5918,N_5929);
or U6158 (N_6158,N_5973,N_5613);
xor U6159 (N_6159,N_5696,N_5500);
nand U6160 (N_6160,N_5508,N_5618);
or U6161 (N_6161,N_5823,N_5626);
and U6162 (N_6162,N_5905,N_5945);
nand U6163 (N_6163,N_5579,N_5662);
and U6164 (N_6164,N_5764,N_5580);
nand U6165 (N_6165,N_5761,N_5885);
xor U6166 (N_6166,N_5667,N_5583);
nor U6167 (N_6167,N_5897,N_5697);
or U6168 (N_6168,N_5762,N_5846);
and U6169 (N_6169,N_5887,N_5752);
xnor U6170 (N_6170,N_5970,N_5511);
or U6171 (N_6171,N_5793,N_5902);
xor U6172 (N_6172,N_5507,N_5818);
or U6173 (N_6173,N_5648,N_5656);
or U6174 (N_6174,N_5546,N_5977);
nor U6175 (N_6175,N_5674,N_5514);
xor U6176 (N_6176,N_5723,N_5817);
xnor U6177 (N_6177,N_5625,N_5599);
or U6178 (N_6178,N_5573,N_5917);
and U6179 (N_6179,N_5690,N_5841);
or U6180 (N_6180,N_5652,N_5726);
nor U6181 (N_6181,N_5556,N_5872);
nand U6182 (N_6182,N_5528,N_5699);
nand U6183 (N_6183,N_5804,N_5644);
nand U6184 (N_6184,N_5947,N_5666);
nor U6185 (N_6185,N_5559,N_5608);
nand U6186 (N_6186,N_5665,N_5965);
nand U6187 (N_6187,N_5976,N_5629);
xor U6188 (N_6188,N_5506,N_5914);
and U6189 (N_6189,N_5795,N_5776);
nand U6190 (N_6190,N_5698,N_5730);
and U6191 (N_6191,N_5847,N_5535);
nand U6192 (N_6192,N_5874,N_5952);
nand U6193 (N_6193,N_5912,N_5501);
nand U6194 (N_6194,N_5963,N_5537);
xor U6195 (N_6195,N_5820,N_5834);
xor U6196 (N_6196,N_5785,N_5748);
nand U6197 (N_6197,N_5828,N_5539);
nor U6198 (N_6198,N_5653,N_5916);
nor U6199 (N_6199,N_5685,N_5753);
or U6200 (N_6200,N_5958,N_5777);
or U6201 (N_6201,N_5852,N_5758);
xor U6202 (N_6202,N_5981,N_5772);
nor U6203 (N_6203,N_5988,N_5739);
nand U6204 (N_6204,N_5798,N_5886);
nor U6205 (N_6205,N_5598,N_5564);
and U6206 (N_6206,N_5590,N_5547);
xor U6207 (N_6207,N_5595,N_5622);
nand U6208 (N_6208,N_5561,N_5831);
nor U6209 (N_6209,N_5679,N_5843);
and U6210 (N_6210,N_5908,N_5810);
nor U6211 (N_6211,N_5882,N_5878);
or U6212 (N_6212,N_5620,N_5526);
or U6213 (N_6213,N_5640,N_5767);
nand U6214 (N_6214,N_5786,N_5814);
xor U6215 (N_6215,N_5684,N_5821);
nand U6216 (N_6216,N_5850,N_5909);
nor U6217 (N_6217,N_5953,N_5728);
xnor U6218 (N_6218,N_5628,N_5520);
nor U6219 (N_6219,N_5870,N_5543);
nand U6220 (N_6220,N_5884,N_5612);
or U6221 (N_6221,N_5545,N_5806);
nand U6222 (N_6222,N_5925,N_5594);
nand U6223 (N_6223,N_5784,N_5780);
or U6224 (N_6224,N_5689,N_5950);
nand U6225 (N_6225,N_5809,N_5812);
nand U6226 (N_6226,N_5582,N_5616);
xnor U6227 (N_6227,N_5533,N_5663);
and U6228 (N_6228,N_5734,N_5940);
xnor U6229 (N_6229,N_5642,N_5978);
xnor U6230 (N_6230,N_5881,N_5725);
or U6231 (N_6231,N_5703,N_5904);
nor U6232 (N_6232,N_5935,N_5961);
xor U6233 (N_6233,N_5569,N_5669);
nor U6234 (N_6234,N_5883,N_5572);
and U6235 (N_6235,N_5554,N_5997);
and U6236 (N_6236,N_5836,N_5933);
nand U6237 (N_6237,N_5861,N_5619);
nand U6238 (N_6238,N_5654,N_5944);
and U6239 (N_6239,N_5729,N_5503);
nand U6240 (N_6240,N_5920,N_5851);
or U6241 (N_6241,N_5930,N_5740);
xnor U6242 (N_6242,N_5645,N_5701);
and U6243 (N_6243,N_5938,N_5650);
nor U6244 (N_6244,N_5879,N_5588);
xnor U6245 (N_6245,N_5708,N_5578);
nor U6246 (N_6246,N_5710,N_5759);
nand U6247 (N_6247,N_5611,N_5783);
and U6248 (N_6248,N_5738,N_5568);
and U6249 (N_6249,N_5617,N_5522);
xnor U6250 (N_6250,N_5910,N_5926);
nand U6251 (N_6251,N_5826,N_5937);
and U6252 (N_6252,N_5587,N_5659);
or U6253 (N_6253,N_5940,N_5976);
or U6254 (N_6254,N_5781,N_5826);
xor U6255 (N_6255,N_5838,N_5509);
nand U6256 (N_6256,N_5704,N_5529);
or U6257 (N_6257,N_5837,N_5680);
or U6258 (N_6258,N_5948,N_5701);
nand U6259 (N_6259,N_5698,N_5651);
nand U6260 (N_6260,N_5843,N_5762);
or U6261 (N_6261,N_5778,N_5701);
or U6262 (N_6262,N_5974,N_5986);
or U6263 (N_6263,N_5875,N_5693);
xnor U6264 (N_6264,N_5629,N_5818);
and U6265 (N_6265,N_5617,N_5586);
xnor U6266 (N_6266,N_5656,N_5741);
or U6267 (N_6267,N_5982,N_5726);
and U6268 (N_6268,N_5570,N_5981);
xnor U6269 (N_6269,N_5540,N_5922);
xnor U6270 (N_6270,N_5991,N_5744);
or U6271 (N_6271,N_5982,N_5640);
nor U6272 (N_6272,N_5803,N_5633);
or U6273 (N_6273,N_5710,N_5653);
nor U6274 (N_6274,N_5838,N_5890);
nor U6275 (N_6275,N_5522,N_5570);
and U6276 (N_6276,N_5784,N_5838);
xor U6277 (N_6277,N_5557,N_5610);
and U6278 (N_6278,N_5943,N_5987);
or U6279 (N_6279,N_5866,N_5962);
nand U6280 (N_6280,N_5866,N_5524);
xor U6281 (N_6281,N_5859,N_5773);
nor U6282 (N_6282,N_5890,N_5981);
nor U6283 (N_6283,N_5745,N_5737);
nand U6284 (N_6284,N_5677,N_5652);
xor U6285 (N_6285,N_5756,N_5662);
nand U6286 (N_6286,N_5701,N_5921);
and U6287 (N_6287,N_5850,N_5873);
or U6288 (N_6288,N_5646,N_5854);
nor U6289 (N_6289,N_5632,N_5553);
nor U6290 (N_6290,N_5969,N_5684);
nor U6291 (N_6291,N_5573,N_5878);
and U6292 (N_6292,N_5930,N_5938);
nor U6293 (N_6293,N_5704,N_5944);
or U6294 (N_6294,N_5758,N_5793);
or U6295 (N_6295,N_5985,N_5661);
and U6296 (N_6296,N_5890,N_5863);
xor U6297 (N_6297,N_5742,N_5931);
nor U6298 (N_6298,N_5546,N_5846);
and U6299 (N_6299,N_5832,N_5542);
nor U6300 (N_6300,N_5654,N_5723);
xor U6301 (N_6301,N_5630,N_5619);
xor U6302 (N_6302,N_5536,N_5770);
or U6303 (N_6303,N_5843,N_5800);
nand U6304 (N_6304,N_5877,N_5883);
nor U6305 (N_6305,N_5511,N_5570);
xnor U6306 (N_6306,N_5971,N_5722);
nand U6307 (N_6307,N_5859,N_5843);
and U6308 (N_6308,N_5819,N_5595);
and U6309 (N_6309,N_5558,N_5609);
nand U6310 (N_6310,N_5873,N_5652);
nor U6311 (N_6311,N_5946,N_5807);
and U6312 (N_6312,N_5683,N_5696);
nor U6313 (N_6313,N_5619,N_5656);
or U6314 (N_6314,N_5662,N_5929);
xnor U6315 (N_6315,N_5507,N_5730);
or U6316 (N_6316,N_5685,N_5693);
and U6317 (N_6317,N_5778,N_5848);
xnor U6318 (N_6318,N_5718,N_5578);
nand U6319 (N_6319,N_5561,N_5690);
nor U6320 (N_6320,N_5895,N_5530);
nand U6321 (N_6321,N_5696,N_5547);
nor U6322 (N_6322,N_5902,N_5923);
and U6323 (N_6323,N_5789,N_5682);
nand U6324 (N_6324,N_5523,N_5969);
and U6325 (N_6325,N_5805,N_5578);
xnor U6326 (N_6326,N_5816,N_5534);
nand U6327 (N_6327,N_5775,N_5645);
xor U6328 (N_6328,N_5772,N_5901);
or U6329 (N_6329,N_5715,N_5569);
or U6330 (N_6330,N_5678,N_5821);
and U6331 (N_6331,N_5916,N_5727);
nand U6332 (N_6332,N_5881,N_5763);
and U6333 (N_6333,N_5616,N_5963);
nor U6334 (N_6334,N_5574,N_5832);
nor U6335 (N_6335,N_5666,N_5786);
xor U6336 (N_6336,N_5596,N_5675);
xor U6337 (N_6337,N_5788,N_5543);
nand U6338 (N_6338,N_5631,N_5956);
and U6339 (N_6339,N_5598,N_5993);
nor U6340 (N_6340,N_5622,N_5827);
and U6341 (N_6341,N_5615,N_5572);
xnor U6342 (N_6342,N_5808,N_5832);
xnor U6343 (N_6343,N_5889,N_5572);
and U6344 (N_6344,N_5866,N_5697);
nand U6345 (N_6345,N_5961,N_5627);
and U6346 (N_6346,N_5918,N_5614);
and U6347 (N_6347,N_5917,N_5861);
xnor U6348 (N_6348,N_5663,N_5742);
and U6349 (N_6349,N_5808,N_5727);
nand U6350 (N_6350,N_5892,N_5891);
nand U6351 (N_6351,N_5841,N_5663);
or U6352 (N_6352,N_5540,N_5940);
or U6353 (N_6353,N_5902,N_5782);
and U6354 (N_6354,N_5924,N_5811);
xnor U6355 (N_6355,N_5501,N_5794);
nand U6356 (N_6356,N_5801,N_5603);
and U6357 (N_6357,N_5724,N_5997);
nand U6358 (N_6358,N_5562,N_5912);
nand U6359 (N_6359,N_5642,N_5847);
and U6360 (N_6360,N_5559,N_5545);
xnor U6361 (N_6361,N_5841,N_5676);
xor U6362 (N_6362,N_5962,N_5829);
xor U6363 (N_6363,N_5794,N_5948);
xnor U6364 (N_6364,N_5824,N_5855);
and U6365 (N_6365,N_5973,N_5520);
nand U6366 (N_6366,N_5784,N_5921);
nor U6367 (N_6367,N_5759,N_5994);
and U6368 (N_6368,N_5712,N_5500);
xor U6369 (N_6369,N_5921,N_5990);
and U6370 (N_6370,N_5538,N_5720);
xor U6371 (N_6371,N_5912,N_5638);
and U6372 (N_6372,N_5602,N_5861);
nand U6373 (N_6373,N_5949,N_5612);
or U6374 (N_6374,N_5768,N_5729);
nand U6375 (N_6375,N_5669,N_5928);
or U6376 (N_6376,N_5749,N_5550);
and U6377 (N_6377,N_5774,N_5793);
xor U6378 (N_6378,N_5965,N_5896);
or U6379 (N_6379,N_5932,N_5749);
or U6380 (N_6380,N_5887,N_5757);
and U6381 (N_6381,N_5599,N_5584);
xor U6382 (N_6382,N_5884,N_5770);
nor U6383 (N_6383,N_5711,N_5740);
nor U6384 (N_6384,N_5756,N_5989);
nor U6385 (N_6385,N_5536,N_5502);
and U6386 (N_6386,N_5855,N_5893);
and U6387 (N_6387,N_5514,N_5664);
or U6388 (N_6388,N_5598,N_5526);
or U6389 (N_6389,N_5576,N_5769);
and U6390 (N_6390,N_5841,N_5797);
or U6391 (N_6391,N_5908,N_5711);
and U6392 (N_6392,N_5641,N_5977);
nor U6393 (N_6393,N_5921,N_5798);
or U6394 (N_6394,N_5670,N_5812);
xnor U6395 (N_6395,N_5944,N_5909);
nand U6396 (N_6396,N_5962,N_5815);
xor U6397 (N_6397,N_5628,N_5874);
or U6398 (N_6398,N_5541,N_5554);
and U6399 (N_6399,N_5595,N_5873);
and U6400 (N_6400,N_5983,N_5800);
and U6401 (N_6401,N_5994,N_5849);
xnor U6402 (N_6402,N_5920,N_5563);
xnor U6403 (N_6403,N_5979,N_5971);
nor U6404 (N_6404,N_5536,N_5814);
or U6405 (N_6405,N_5527,N_5900);
or U6406 (N_6406,N_5880,N_5662);
nand U6407 (N_6407,N_5700,N_5753);
nand U6408 (N_6408,N_5649,N_5502);
nor U6409 (N_6409,N_5793,N_5969);
xnor U6410 (N_6410,N_5757,N_5906);
or U6411 (N_6411,N_5889,N_5542);
nor U6412 (N_6412,N_5991,N_5885);
and U6413 (N_6413,N_5584,N_5756);
xnor U6414 (N_6414,N_5651,N_5772);
xnor U6415 (N_6415,N_5614,N_5555);
or U6416 (N_6416,N_5727,N_5819);
or U6417 (N_6417,N_5922,N_5909);
xor U6418 (N_6418,N_5701,N_5803);
or U6419 (N_6419,N_5860,N_5565);
xnor U6420 (N_6420,N_5611,N_5759);
nand U6421 (N_6421,N_5713,N_5928);
nand U6422 (N_6422,N_5840,N_5627);
and U6423 (N_6423,N_5548,N_5837);
xnor U6424 (N_6424,N_5969,N_5867);
xnor U6425 (N_6425,N_5803,N_5540);
nand U6426 (N_6426,N_5524,N_5827);
xor U6427 (N_6427,N_5677,N_5701);
nand U6428 (N_6428,N_5650,N_5721);
and U6429 (N_6429,N_5535,N_5860);
nand U6430 (N_6430,N_5829,N_5902);
xnor U6431 (N_6431,N_5944,N_5531);
xnor U6432 (N_6432,N_5761,N_5617);
or U6433 (N_6433,N_5512,N_5903);
nand U6434 (N_6434,N_5699,N_5552);
and U6435 (N_6435,N_5980,N_5692);
nor U6436 (N_6436,N_5583,N_5610);
and U6437 (N_6437,N_5856,N_5505);
nand U6438 (N_6438,N_5880,N_5572);
or U6439 (N_6439,N_5818,N_5592);
nand U6440 (N_6440,N_5532,N_5811);
and U6441 (N_6441,N_5656,N_5633);
xor U6442 (N_6442,N_5758,N_5790);
nand U6443 (N_6443,N_5664,N_5599);
xnor U6444 (N_6444,N_5964,N_5945);
and U6445 (N_6445,N_5679,N_5736);
and U6446 (N_6446,N_5730,N_5807);
or U6447 (N_6447,N_5663,N_5677);
nor U6448 (N_6448,N_5706,N_5738);
or U6449 (N_6449,N_5756,N_5665);
and U6450 (N_6450,N_5520,N_5855);
and U6451 (N_6451,N_5711,N_5923);
nor U6452 (N_6452,N_5804,N_5623);
xnor U6453 (N_6453,N_5914,N_5899);
nor U6454 (N_6454,N_5635,N_5880);
nor U6455 (N_6455,N_5618,N_5526);
xor U6456 (N_6456,N_5823,N_5593);
or U6457 (N_6457,N_5502,N_5660);
or U6458 (N_6458,N_5950,N_5970);
nand U6459 (N_6459,N_5539,N_5582);
xor U6460 (N_6460,N_5864,N_5680);
nor U6461 (N_6461,N_5881,N_5699);
nor U6462 (N_6462,N_5980,N_5950);
xnor U6463 (N_6463,N_5795,N_5880);
and U6464 (N_6464,N_5903,N_5866);
nand U6465 (N_6465,N_5507,N_5803);
nor U6466 (N_6466,N_5935,N_5504);
nand U6467 (N_6467,N_5826,N_5960);
and U6468 (N_6468,N_5786,N_5844);
nand U6469 (N_6469,N_5506,N_5626);
nor U6470 (N_6470,N_5670,N_5813);
nor U6471 (N_6471,N_5604,N_5879);
or U6472 (N_6472,N_5506,N_5502);
xor U6473 (N_6473,N_5904,N_5930);
nand U6474 (N_6474,N_5850,N_5705);
nand U6475 (N_6475,N_5516,N_5800);
or U6476 (N_6476,N_5837,N_5725);
xnor U6477 (N_6477,N_5601,N_5578);
and U6478 (N_6478,N_5773,N_5832);
nor U6479 (N_6479,N_5605,N_5811);
nor U6480 (N_6480,N_5577,N_5537);
xor U6481 (N_6481,N_5823,N_5841);
and U6482 (N_6482,N_5555,N_5525);
xor U6483 (N_6483,N_5907,N_5534);
nand U6484 (N_6484,N_5807,N_5647);
and U6485 (N_6485,N_5943,N_5679);
nand U6486 (N_6486,N_5638,N_5665);
nand U6487 (N_6487,N_5864,N_5747);
or U6488 (N_6488,N_5766,N_5912);
nand U6489 (N_6489,N_5675,N_5767);
and U6490 (N_6490,N_5969,N_5723);
and U6491 (N_6491,N_5983,N_5869);
and U6492 (N_6492,N_5811,N_5853);
and U6493 (N_6493,N_5720,N_5543);
and U6494 (N_6494,N_5520,N_5763);
nor U6495 (N_6495,N_5625,N_5519);
nor U6496 (N_6496,N_5581,N_5621);
nand U6497 (N_6497,N_5651,N_5974);
nor U6498 (N_6498,N_5860,N_5931);
and U6499 (N_6499,N_5863,N_5901);
nor U6500 (N_6500,N_6253,N_6245);
and U6501 (N_6501,N_6268,N_6175);
nor U6502 (N_6502,N_6183,N_6275);
nor U6503 (N_6503,N_6481,N_6076);
nand U6504 (N_6504,N_6453,N_6218);
or U6505 (N_6505,N_6290,N_6226);
or U6506 (N_6506,N_6238,N_6373);
nand U6507 (N_6507,N_6011,N_6360);
and U6508 (N_6508,N_6330,N_6000);
or U6509 (N_6509,N_6427,N_6446);
xor U6510 (N_6510,N_6292,N_6270);
or U6511 (N_6511,N_6083,N_6331);
nand U6512 (N_6512,N_6364,N_6149);
or U6513 (N_6513,N_6469,N_6036);
xnor U6514 (N_6514,N_6310,N_6302);
xor U6515 (N_6515,N_6298,N_6382);
nand U6516 (N_6516,N_6420,N_6172);
and U6517 (N_6517,N_6283,N_6239);
nor U6518 (N_6518,N_6317,N_6230);
or U6519 (N_6519,N_6378,N_6143);
nand U6520 (N_6520,N_6102,N_6067);
nor U6521 (N_6521,N_6034,N_6107);
xnor U6522 (N_6522,N_6424,N_6208);
xor U6523 (N_6523,N_6072,N_6397);
or U6524 (N_6524,N_6012,N_6115);
and U6525 (N_6525,N_6286,N_6403);
nand U6526 (N_6526,N_6256,N_6486);
nand U6527 (N_6527,N_6308,N_6181);
or U6528 (N_6528,N_6164,N_6435);
nor U6529 (N_6529,N_6356,N_6161);
nor U6530 (N_6530,N_6361,N_6179);
nand U6531 (N_6531,N_6147,N_6399);
and U6532 (N_6532,N_6199,N_6065);
nand U6533 (N_6533,N_6440,N_6140);
nor U6534 (N_6534,N_6018,N_6359);
or U6535 (N_6535,N_6213,N_6341);
or U6536 (N_6536,N_6030,N_6125);
and U6537 (N_6537,N_6422,N_6372);
nor U6538 (N_6538,N_6200,N_6212);
nand U6539 (N_6539,N_6152,N_6362);
and U6540 (N_6540,N_6309,N_6484);
and U6541 (N_6541,N_6233,N_6137);
xor U6542 (N_6542,N_6479,N_6185);
xor U6543 (N_6543,N_6131,N_6097);
or U6544 (N_6544,N_6421,N_6186);
or U6545 (N_6545,N_6354,N_6414);
nand U6546 (N_6546,N_6498,N_6074);
xor U6547 (N_6547,N_6258,N_6351);
nand U6548 (N_6548,N_6120,N_6350);
nand U6549 (N_6549,N_6098,N_6263);
and U6550 (N_6550,N_6130,N_6059);
or U6551 (N_6551,N_6023,N_6005);
and U6552 (N_6552,N_6156,N_6346);
nor U6553 (N_6553,N_6325,N_6105);
and U6554 (N_6554,N_6339,N_6116);
and U6555 (N_6555,N_6473,N_6291);
xor U6556 (N_6556,N_6410,N_6202);
and U6557 (N_6557,N_6347,N_6269);
or U6558 (N_6558,N_6138,N_6142);
nand U6559 (N_6559,N_6345,N_6439);
nor U6560 (N_6560,N_6264,N_6419);
or U6561 (N_6561,N_6189,N_6044);
and U6562 (N_6562,N_6017,N_6318);
xnor U6563 (N_6563,N_6322,N_6461);
xor U6564 (N_6564,N_6307,N_6383);
nand U6565 (N_6565,N_6124,N_6004);
nand U6566 (N_6566,N_6216,N_6048);
and U6567 (N_6567,N_6211,N_6122);
nor U6568 (N_6568,N_6338,N_6288);
xnor U6569 (N_6569,N_6340,N_6171);
and U6570 (N_6570,N_6118,N_6089);
xnor U6571 (N_6571,N_6304,N_6398);
xnor U6572 (N_6572,N_6491,N_6153);
xor U6573 (N_6573,N_6159,N_6321);
nor U6574 (N_6574,N_6280,N_6032);
or U6575 (N_6575,N_6085,N_6386);
or U6576 (N_6576,N_6002,N_6445);
and U6577 (N_6577,N_6454,N_6141);
xnor U6578 (N_6578,N_6470,N_6409);
or U6579 (N_6579,N_6111,N_6126);
or U6580 (N_6580,N_6042,N_6073);
nand U6581 (N_6581,N_6038,N_6394);
or U6582 (N_6582,N_6084,N_6029);
and U6583 (N_6583,N_6196,N_6492);
xnor U6584 (N_6584,N_6001,N_6224);
nor U6585 (N_6585,N_6274,N_6187);
xnor U6586 (N_6586,N_6231,N_6066);
and U6587 (N_6587,N_6136,N_6430);
xnor U6588 (N_6588,N_6015,N_6062);
nor U6589 (N_6589,N_6476,N_6203);
nand U6590 (N_6590,N_6236,N_6475);
or U6591 (N_6591,N_6123,N_6401);
and U6592 (N_6592,N_6374,N_6194);
nand U6593 (N_6593,N_6027,N_6020);
or U6594 (N_6594,N_6094,N_6244);
xnor U6595 (N_6595,N_6154,N_6367);
nor U6596 (N_6596,N_6273,N_6285);
nand U6597 (N_6597,N_6313,N_6379);
nand U6598 (N_6598,N_6092,N_6369);
and U6599 (N_6599,N_6495,N_6058);
or U6600 (N_6600,N_6319,N_6037);
xnor U6601 (N_6601,N_6197,N_6174);
nand U6602 (N_6602,N_6163,N_6462);
xor U6603 (N_6603,N_6054,N_6243);
nand U6604 (N_6604,N_6443,N_6260);
xor U6605 (N_6605,N_6297,N_6234);
xor U6606 (N_6606,N_6281,N_6381);
nor U6607 (N_6607,N_6368,N_6068);
nor U6608 (N_6608,N_6348,N_6150);
xnor U6609 (N_6609,N_6184,N_6235);
xor U6610 (N_6610,N_6496,N_6464);
or U6611 (N_6611,N_6384,N_6485);
or U6612 (N_6612,N_6342,N_6293);
and U6613 (N_6613,N_6240,N_6219);
nor U6614 (N_6614,N_6389,N_6405);
and U6615 (N_6615,N_6371,N_6315);
nor U6616 (N_6616,N_6333,N_6447);
and U6617 (N_6617,N_6468,N_6434);
xor U6618 (N_6618,N_6177,N_6472);
nor U6619 (N_6619,N_6220,N_6099);
nor U6620 (N_6620,N_6432,N_6489);
or U6621 (N_6621,N_6474,N_6046);
or U6622 (N_6622,N_6225,N_6214);
nor U6623 (N_6623,N_6003,N_6249);
and U6624 (N_6624,N_6449,N_6078);
nor U6625 (N_6625,N_6349,N_6459);
nor U6626 (N_6626,N_6114,N_6113);
xnor U6627 (N_6627,N_6408,N_6128);
nand U6628 (N_6628,N_6336,N_6391);
and U6629 (N_6629,N_6229,N_6277);
xor U6630 (N_6630,N_6148,N_6494);
and U6631 (N_6631,N_6395,N_6357);
nand U6632 (N_6632,N_6320,N_6262);
or U6633 (N_6633,N_6077,N_6019);
and U6634 (N_6634,N_6190,N_6259);
and U6635 (N_6635,N_6396,N_6413);
and U6636 (N_6636,N_6488,N_6400);
or U6637 (N_6637,N_6303,N_6039);
nor U6638 (N_6638,N_6222,N_6178);
nand U6639 (N_6639,N_6271,N_6326);
or U6640 (N_6640,N_6100,N_6112);
nor U6641 (N_6641,N_6021,N_6402);
nand U6642 (N_6642,N_6035,N_6248);
and U6643 (N_6643,N_6109,N_6287);
nor U6644 (N_6644,N_6306,N_6477);
nor U6645 (N_6645,N_6314,N_6296);
or U6646 (N_6646,N_6117,N_6119);
nand U6647 (N_6647,N_6478,N_6146);
nand U6648 (N_6648,N_6192,N_6441);
and U6649 (N_6649,N_6370,N_6110);
nand U6650 (N_6650,N_6053,N_6327);
xnor U6651 (N_6651,N_6416,N_6375);
nor U6652 (N_6652,N_6180,N_6157);
xnor U6653 (N_6653,N_6407,N_6438);
and U6654 (N_6654,N_6193,N_6201);
or U6655 (N_6655,N_6366,N_6063);
and U6656 (N_6656,N_6376,N_6428);
or U6657 (N_6657,N_6237,N_6444);
nor U6658 (N_6658,N_6466,N_6047);
and U6659 (N_6659,N_6052,N_6377);
xnor U6660 (N_6660,N_6168,N_6355);
xor U6661 (N_6661,N_6301,N_6344);
nand U6662 (N_6662,N_6010,N_6431);
nand U6663 (N_6663,N_6448,N_6075);
xor U6664 (N_6664,N_6311,N_6064);
nand U6665 (N_6665,N_6133,N_6255);
nor U6666 (N_6666,N_6204,N_6079);
xnor U6667 (N_6667,N_6300,N_6108);
nand U6668 (N_6668,N_6289,N_6095);
nand U6669 (N_6669,N_6254,N_6247);
nand U6670 (N_6670,N_6134,N_6467);
nor U6671 (N_6671,N_6106,N_6265);
or U6672 (N_6672,N_6206,N_6006);
xor U6673 (N_6673,N_6104,N_6436);
nor U6674 (N_6674,N_6393,N_6312);
nand U6675 (N_6675,N_6267,N_6250);
nor U6676 (N_6676,N_6080,N_6127);
nor U6677 (N_6677,N_6025,N_6071);
nor U6678 (N_6678,N_6167,N_6279);
and U6679 (N_6679,N_6182,N_6090);
nor U6680 (N_6680,N_6013,N_6057);
nand U6681 (N_6681,N_6417,N_6014);
nor U6682 (N_6682,N_6166,N_6324);
or U6683 (N_6683,N_6404,N_6337);
nor U6684 (N_6684,N_6009,N_6016);
nor U6685 (N_6685,N_6132,N_6056);
or U6686 (N_6686,N_6028,N_6335);
xnor U6687 (N_6687,N_6284,N_6261);
nand U6688 (N_6688,N_6195,N_6144);
xor U6689 (N_6689,N_6352,N_6455);
or U6690 (N_6690,N_6087,N_6343);
nand U6691 (N_6691,N_6429,N_6433);
nand U6692 (N_6692,N_6103,N_6165);
nor U6693 (N_6693,N_6101,N_6129);
or U6694 (N_6694,N_6483,N_6460);
nand U6695 (N_6695,N_6257,N_6385);
nand U6696 (N_6696,N_6232,N_6049);
and U6697 (N_6697,N_6266,N_6278);
nand U6698 (N_6698,N_6471,N_6463);
nand U6699 (N_6699,N_6033,N_6198);
xor U6700 (N_6700,N_6051,N_6365);
xnor U6701 (N_6701,N_6145,N_6155);
nand U6702 (N_6702,N_6437,N_6412);
xnor U6703 (N_6703,N_6299,N_6031);
or U6704 (N_6704,N_6426,N_6205);
nor U6705 (N_6705,N_6227,N_6041);
xnor U6706 (N_6706,N_6423,N_6380);
or U6707 (N_6707,N_6295,N_6209);
nand U6708 (N_6708,N_6328,N_6242);
or U6709 (N_6709,N_6294,N_6387);
nor U6710 (N_6710,N_6353,N_6252);
or U6711 (N_6711,N_6050,N_6411);
nor U6712 (N_6712,N_6026,N_6043);
nor U6713 (N_6713,N_6221,N_6045);
nor U6714 (N_6714,N_6480,N_6139);
and U6715 (N_6715,N_6061,N_6497);
xor U6716 (N_6716,N_6188,N_6228);
or U6717 (N_6717,N_6363,N_6091);
xor U6718 (N_6718,N_6173,N_6316);
nor U6719 (N_6719,N_6329,N_6215);
nand U6720 (N_6720,N_6246,N_6388);
nor U6721 (N_6721,N_6450,N_6418);
or U6722 (N_6722,N_6358,N_6169);
nor U6723 (N_6723,N_6055,N_6207);
nor U6724 (N_6724,N_6465,N_6332);
and U6725 (N_6725,N_6191,N_6490);
nor U6726 (N_6726,N_6499,N_6088);
or U6727 (N_6727,N_6070,N_6007);
and U6728 (N_6728,N_6176,N_6415);
nand U6729 (N_6729,N_6323,N_6334);
nor U6730 (N_6730,N_6482,N_6272);
nor U6731 (N_6731,N_6458,N_6008);
and U6732 (N_6732,N_6086,N_6082);
or U6733 (N_6733,N_6457,N_6069);
nand U6734 (N_6734,N_6210,N_6060);
nor U6735 (N_6735,N_6024,N_6241);
or U6736 (N_6736,N_6392,N_6040);
nand U6737 (N_6737,N_6162,N_6487);
and U6738 (N_6738,N_6282,N_6456);
nand U6739 (N_6739,N_6158,N_6390);
and U6740 (N_6740,N_6425,N_6135);
xor U6741 (N_6741,N_6217,N_6160);
nand U6742 (N_6742,N_6096,N_6452);
nor U6743 (N_6743,N_6121,N_6170);
nor U6744 (N_6744,N_6406,N_6251);
or U6745 (N_6745,N_6276,N_6022);
nor U6746 (N_6746,N_6223,N_6093);
xor U6747 (N_6747,N_6151,N_6451);
or U6748 (N_6748,N_6305,N_6493);
xnor U6749 (N_6749,N_6081,N_6442);
or U6750 (N_6750,N_6384,N_6183);
and U6751 (N_6751,N_6248,N_6397);
xnor U6752 (N_6752,N_6187,N_6284);
xnor U6753 (N_6753,N_6179,N_6187);
nor U6754 (N_6754,N_6457,N_6002);
nand U6755 (N_6755,N_6033,N_6359);
xor U6756 (N_6756,N_6041,N_6146);
xor U6757 (N_6757,N_6360,N_6192);
and U6758 (N_6758,N_6314,N_6128);
nand U6759 (N_6759,N_6215,N_6290);
and U6760 (N_6760,N_6080,N_6277);
or U6761 (N_6761,N_6219,N_6408);
nor U6762 (N_6762,N_6416,N_6302);
nor U6763 (N_6763,N_6104,N_6256);
or U6764 (N_6764,N_6368,N_6410);
xor U6765 (N_6765,N_6031,N_6124);
or U6766 (N_6766,N_6350,N_6392);
or U6767 (N_6767,N_6319,N_6385);
or U6768 (N_6768,N_6146,N_6246);
xor U6769 (N_6769,N_6166,N_6351);
and U6770 (N_6770,N_6034,N_6484);
and U6771 (N_6771,N_6144,N_6051);
or U6772 (N_6772,N_6309,N_6210);
xnor U6773 (N_6773,N_6048,N_6494);
nand U6774 (N_6774,N_6130,N_6241);
and U6775 (N_6775,N_6289,N_6475);
xnor U6776 (N_6776,N_6110,N_6228);
nand U6777 (N_6777,N_6342,N_6143);
nand U6778 (N_6778,N_6407,N_6131);
nand U6779 (N_6779,N_6487,N_6128);
nand U6780 (N_6780,N_6322,N_6444);
xnor U6781 (N_6781,N_6480,N_6482);
or U6782 (N_6782,N_6474,N_6333);
xor U6783 (N_6783,N_6111,N_6235);
or U6784 (N_6784,N_6173,N_6351);
nand U6785 (N_6785,N_6051,N_6012);
or U6786 (N_6786,N_6383,N_6157);
nor U6787 (N_6787,N_6490,N_6295);
nand U6788 (N_6788,N_6271,N_6391);
nor U6789 (N_6789,N_6435,N_6242);
nor U6790 (N_6790,N_6076,N_6061);
xor U6791 (N_6791,N_6400,N_6077);
xor U6792 (N_6792,N_6093,N_6107);
nand U6793 (N_6793,N_6368,N_6446);
nand U6794 (N_6794,N_6359,N_6338);
nand U6795 (N_6795,N_6120,N_6441);
xor U6796 (N_6796,N_6367,N_6349);
nand U6797 (N_6797,N_6471,N_6427);
xor U6798 (N_6798,N_6376,N_6155);
nand U6799 (N_6799,N_6324,N_6041);
nand U6800 (N_6800,N_6107,N_6428);
xor U6801 (N_6801,N_6418,N_6227);
nor U6802 (N_6802,N_6137,N_6170);
or U6803 (N_6803,N_6251,N_6398);
xnor U6804 (N_6804,N_6358,N_6326);
and U6805 (N_6805,N_6203,N_6445);
xnor U6806 (N_6806,N_6323,N_6202);
or U6807 (N_6807,N_6370,N_6249);
or U6808 (N_6808,N_6192,N_6034);
nor U6809 (N_6809,N_6123,N_6117);
nand U6810 (N_6810,N_6098,N_6075);
nor U6811 (N_6811,N_6002,N_6178);
xor U6812 (N_6812,N_6177,N_6455);
and U6813 (N_6813,N_6416,N_6075);
and U6814 (N_6814,N_6438,N_6022);
xnor U6815 (N_6815,N_6374,N_6466);
or U6816 (N_6816,N_6191,N_6437);
and U6817 (N_6817,N_6471,N_6155);
and U6818 (N_6818,N_6038,N_6039);
or U6819 (N_6819,N_6027,N_6043);
and U6820 (N_6820,N_6428,N_6315);
nand U6821 (N_6821,N_6046,N_6470);
nand U6822 (N_6822,N_6441,N_6407);
and U6823 (N_6823,N_6129,N_6293);
or U6824 (N_6824,N_6224,N_6327);
or U6825 (N_6825,N_6408,N_6150);
and U6826 (N_6826,N_6057,N_6320);
and U6827 (N_6827,N_6335,N_6133);
nor U6828 (N_6828,N_6041,N_6143);
nor U6829 (N_6829,N_6226,N_6054);
nor U6830 (N_6830,N_6429,N_6042);
xnor U6831 (N_6831,N_6003,N_6045);
and U6832 (N_6832,N_6322,N_6053);
or U6833 (N_6833,N_6008,N_6186);
and U6834 (N_6834,N_6468,N_6287);
nor U6835 (N_6835,N_6380,N_6206);
nor U6836 (N_6836,N_6430,N_6351);
xor U6837 (N_6837,N_6463,N_6316);
and U6838 (N_6838,N_6388,N_6229);
and U6839 (N_6839,N_6047,N_6390);
nor U6840 (N_6840,N_6414,N_6244);
nand U6841 (N_6841,N_6483,N_6398);
xnor U6842 (N_6842,N_6323,N_6395);
or U6843 (N_6843,N_6081,N_6288);
xor U6844 (N_6844,N_6063,N_6336);
nor U6845 (N_6845,N_6133,N_6441);
or U6846 (N_6846,N_6357,N_6214);
nand U6847 (N_6847,N_6103,N_6482);
or U6848 (N_6848,N_6116,N_6245);
and U6849 (N_6849,N_6469,N_6250);
xor U6850 (N_6850,N_6052,N_6104);
xnor U6851 (N_6851,N_6192,N_6359);
xor U6852 (N_6852,N_6421,N_6405);
xnor U6853 (N_6853,N_6010,N_6381);
nand U6854 (N_6854,N_6183,N_6295);
nor U6855 (N_6855,N_6348,N_6178);
nand U6856 (N_6856,N_6063,N_6188);
or U6857 (N_6857,N_6044,N_6338);
and U6858 (N_6858,N_6477,N_6179);
nor U6859 (N_6859,N_6261,N_6227);
nand U6860 (N_6860,N_6089,N_6152);
and U6861 (N_6861,N_6266,N_6261);
or U6862 (N_6862,N_6087,N_6434);
nor U6863 (N_6863,N_6048,N_6188);
xnor U6864 (N_6864,N_6158,N_6456);
xnor U6865 (N_6865,N_6395,N_6440);
nand U6866 (N_6866,N_6074,N_6043);
xnor U6867 (N_6867,N_6177,N_6237);
nand U6868 (N_6868,N_6012,N_6064);
and U6869 (N_6869,N_6179,N_6341);
nor U6870 (N_6870,N_6371,N_6222);
or U6871 (N_6871,N_6470,N_6197);
xor U6872 (N_6872,N_6149,N_6429);
nand U6873 (N_6873,N_6286,N_6006);
nand U6874 (N_6874,N_6168,N_6396);
and U6875 (N_6875,N_6366,N_6124);
or U6876 (N_6876,N_6082,N_6065);
nand U6877 (N_6877,N_6204,N_6152);
xor U6878 (N_6878,N_6345,N_6466);
xnor U6879 (N_6879,N_6082,N_6457);
and U6880 (N_6880,N_6453,N_6290);
and U6881 (N_6881,N_6049,N_6240);
xnor U6882 (N_6882,N_6090,N_6112);
nand U6883 (N_6883,N_6323,N_6234);
nor U6884 (N_6884,N_6398,N_6141);
xor U6885 (N_6885,N_6351,N_6114);
xnor U6886 (N_6886,N_6295,N_6235);
and U6887 (N_6887,N_6368,N_6085);
xnor U6888 (N_6888,N_6416,N_6257);
xor U6889 (N_6889,N_6098,N_6488);
nand U6890 (N_6890,N_6159,N_6496);
or U6891 (N_6891,N_6125,N_6023);
xor U6892 (N_6892,N_6066,N_6466);
nand U6893 (N_6893,N_6466,N_6289);
nor U6894 (N_6894,N_6035,N_6434);
nand U6895 (N_6895,N_6474,N_6028);
or U6896 (N_6896,N_6136,N_6127);
and U6897 (N_6897,N_6407,N_6463);
and U6898 (N_6898,N_6387,N_6031);
nor U6899 (N_6899,N_6245,N_6129);
nand U6900 (N_6900,N_6269,N_6452);
or U6901 (N_6901,N_6136,N_6194);
xnor U6902 (N_6902,N_6320,N_6021);
nor U6903 (N_6903,N_6000,N_6393);
nand U6904 (N_6904,N_6133,N_6487);
nor U6905 (N_6905,N_6021,N_6195);
or U6906 (N_6906,N_6263,N_6231);
nand U6907 (N_6907,N_6228,N_6002);
and U6908 (N_6908,N_6358,N_6247);
nor U6909 (N_6909,N_6184,N_6031);
nor U6910 (N_6910,N_6046,N_6112);
and U6911 (N_6911,N_6060,N_6221);
nor U6912 (N_6912,N_6123,N_6210);
nand U6913 (N_6913,N_6069,N_6212);
xor U6914 (N_6914,N_6410,N_6304);
or U6915 (N_6915,N_6471,N_6469);
nor U6916 (N_6916,N_6173,N_6379);
xnor U6917 (N_6917,N_6202,N_6092);
nor U6918 (N_6918,N_6408,N_6098);
nor U6919 (N_6919,N_6450,N_6291);
and U6920 (N_6920,N_6092,N_6124);
or U6921 (N_6921,N_6004,N_6404);
nor U6922 (N_6922,N_6297,N_6332);
or U6923 (N_6923,N_6005,N_6317);
nor U6924 (N_6924,N_6312,N_6297);
nand U6925 (N_6925,N_6002,N_6233);
nor U6926 (N_6926,N_6291,N_6337);
or U6927 (N_6927,N_6190,N_6282);
nand U6928 (N_6928,N_6132,N_6384);
xor U6929 (N_6929,N_6371,N_6312);
or U6930 (N_6930,N_6004,N_6200);
nand U6931 (N_6931,N_6144,N_6450);
nand U6932 (N_6932,N_6363,N_6011);
nand U6933 (N_6933,N_6240,N_6469);
nor U6934 (N_6934,N_6080,N_6332);
or U6935 (N_6935,N_6238,N_6008);
xnor U6936 (N_6936,N_6331,N_6418);
and U6937 (N_6937,N_6113,N_6237);
nand U6938 (N_6938,N_6058,N_6271);
nor U6939 (N_6939,N_6450,N_6269);
nor U6940 (N_6940,N_6329,N_6076);
xor U6941 (N_6941,N_6240,N_6388);
or U6942 (N_6942,N_6412,N_6290);
xor U6943 (N_6943,N_6477,N_6332);
or U6944 (N_6944,N_6081,N_6299);
or U6945 (N_6945,N_6499,N_6270);
nand U6946 (N_6946,N_6121,N_6423);
nor U6947 (N_6947,N_6424,N_6080);
and U6948 (N_6948,N_6400,N_6463);
nand U6949 (N_6949,N_6490,N_6391);
nand U6950 (N_6950,N_6079,N_6052);
xor U6951 (N_6951,N_6169,N_6137);
nand U6952 (N_6952,N_6115,N_6258);
xnor U6953 (N_6953,N_6015,N_6467);
nand U6954 (N_6954,N_6229,N_6427);
nand U6955 (N_6955,N_6051,N_6004);
or U6956 (N_6956,N_6378,N_6485);
nand U6957 (N_6957,N_6244,N_6044);
xor U6958 (N_6958,N_6344,N_6390);
nand U6959 (N_6959,N_6208,N_6320);
and U6960 (N_6960,N_6499,N_6434);
nor U6961 (N_6961,N_6467,N_6023);
or U6962 (N_6962,N_6243,N_6006);
nand U6963 (N_6963,N_6000,N_6097);
nor U6964 (N_6964,N_6325,N_6287);
or U6965 (N_6965,N_6374,N_6338);
or U6966 (N_6966,N_6420,N_6394);
nand U6967 (N_6967,N_6006,N_6161);
and U6968 (N_6968,N_6317,N_6362);
nand U6969 (N_6969,N_6381,N_6342);
nand U6970 (N_6970,N_6489,N_6097);
nand U6971 (N_6971,N_6378,N_6276);
or U6972 (N_6972,N_6236,N_6370);
and U6973 (N_6973,N_6101,N_6112);
nor U6974 (N_6974,N_6123,N_6245);
nor U6975 (N_6975,N_6390,N_6196);
xnor U6976 (N_6976,N_6077,N_6348);
and U6977 (N_6977,N_6401,N_6249);
xnor U6978 (N_6978,N_6380,N_6403);
or U6979 (N_6979,N_6422,N_6394);
or U6980 (N_6980,N_6064,N_6226);
xor U6981 (N_6981,N_6375,N_6020);
or U6982 (N_6982,N_6370,N_6268);
nor U6983 (N_6983,N_6081,N_6349);
and U6984 (N_6984,N_6398,N_6154);
xnor U6985 (N_6985,N_6343,N_6067);
xnor U6986 (N_6986,N_6474,N_6478);
and U6987 (N_6987,N_6202,N_6137);
and U6988 (N_6988,N_6344,N_6239);
nor U6989 (N_6989,N_6474,N_6020);
nor U6990 (N_6990,N_6303,N_6144);
nor U6991 (N_6991,N_6354,N_6140);
and U6992 (N_6992,N_6092,N_6399);
xnor U6993 (N_6993,N_6116,N_6386);
nor U6994 (N_6994,N_6383,N_6488);
and U6995 (N_6995,N_6130,N_6370);
nand U6996 (N_6996,N_6368,N_6326);
nand U6997 (N_6997,N_6126,N_6173);
nand U6998 (N_6998,N_6085,N_6252);
and U6999 (N_6999,N_6312,N_6091);
xor U7000 (N_7000,N_6800,N_6504);
nor U7001 (N_7001,N_6868,N_6772);
nand U7002 (N_7002,N_6955,N_6838);
and U7003 (N_7003,N_6848,N_6825);
or U7004 (N_7004,N_6974,N_6887);
xnor U7005 (N_7005,N_6514,N_6875);
or U7006 (N_7006,N_6643,N_6761);
and U7007 (N_7007,N_6522,N_6689);
nor U7008 (N_7008,N_6746,N_6702);
nor U7009 (N_7009,N_6804,N_6932);
nand U7010 (N_7010,N_6742,N_6529);
nand U7011 (N_7011,N_6707,N_6612);
nand U7012 (N_7012,N_6677,N_6560);
nor U7013 (N_7013,N_6777,N_6510);
nor U7014 (N_7014,N_6970,N_6715);
xnor U7015 (N_7015,N_6518,N_6999);
nor U7016 (N_7016,N_6841,N_6939);
or U7017 (N_7017,N_6566,N_6549);
and U7018 (N_7018,N_6571,N_6704);
nand U7019 (N_7019,N_6541,N_6521);
xor U7020 (N_7020,N_6894,N_6613);
xnor U7021 (N_7021,N_6703,N_6821);
nand U7022 (N_7022,N_6796,N_6556);
xnor U7023 (N_7023,N_6992,N_6898);
and U7024 (N_7024,N_6771,N_6899);
nand U7025 (N_7025,N_6879,N_6506);
nor U7026 (N_7026,N_6544,N_6591);
xor U7027 (N_7027,N_6980,N_6997);
xnor U7028 (N_7028,N_6690,N_6706);
nand U7029 (N_7029,N_6512,N_6819);
xor U7030 (N_7030,N_6513,N_6602);
and U7031 (N_7031,N_6749,N_6667);
or U7032 (N_7032,N_6880,N_6908);
and U7033 (N_7033,N_6760,N_6826);
or U7034 (N_7034,N_6824,N_6553);
or U7035 (N_7035,N_6960,N_6629);
nor U7036 (N_7036,N_6882,N_6842);
and U7037 (N_7037,N_6928,N_6990);
or U7038 (N_7038,N_6876,N_6666);
xnor U7039 (N_7039,N_6705,N_6779);
and U7040 (N_7040,N_6565,N_6682);
nor U7041 (N_7041,N_6614,N_6993);
xor U7042 (N_7042,N_6603,N_6878);
or U7043 (N_7043,N_6935,N_6822);
xnor U7044 (N_7044,N_6859,N_6937);
nand U7045 (N_7045,N_6710,N_6924);
and U7046 (N_7046,N_6891,N_6526);
and U7047 (N_7047,N_6670,N_6871);
nor U7048 (N_7048,N_6776,N_6775);
or U7049 (N_7049,N_6797,N_6743);
and U7050 (N_7050,N_6933,N_6839);
and U7051 (N_7051,N_6609,N_6605);
xnor U7052 (N_7052,N_6792,N_6511);
nor U7053 (N_7053,N_6691,N_6794);
and U7054 (N_7054,N_6906,N_6961);
nor U7055 (N_7055,N_6720,N_6641);
and U7056 (N_7056,N_6920,N_6642);
and U7057 (N_7057,N_6583,N_6663);
and U7058 (N_7058,N_6767,N_6930);
or U7059 (N_7059,N_6550,N_6534);
and U7060 (N_7060,N_6595,N_6696);
xor U7061 (N_7061,N_6719,N_6991);
nor U7062 (N_7062,N_6814,N_6538);
xnor U7063 (N_7063,N_6721,N_6558);
and U7064 (N_7064,N_6590,N_6766);
nand U7065 (N_7065,N_6733,N_6533);
nand U7066 (N_7066,N_6620,N_6668);
nand U7067 (N_7067,N_6658,N_6604);
nand U7068 (N_7068,N_6503,N_6922);
or U7069 (N_7069,N_6919,N_6686);
nand U7070 (N_7070,N_6574,N_6734);
and U7071 (N_7071,N_6874,N_6805);
nor U7072 (N_7072,N_6896,N_6537);
nand U7073 (N_7073,N_6627,N_6981);
or U7074 (N_7074,N_6827,N_6921);
nand U7075 (N_7075,N_6768,N_6585);
xnor U7076 (N_7076,N_6884,N_6692);
or U7077 (N_7077,N_6925,N_6855);
nand U7078 (N_7078,N_6659,N_6647);
xor U7079 (N_7079,N_6946,N_6632);
and U7080 (N_7080,N_6845,N_6802);
or U7081 (N_7081,N_6987,N_6649);
nor U7082 (N_7082,N_6867,N_6672);
or U7083 (N_7083,N_6739,N_6547);
and U7084 (N_7084,N_6854,N_6587);
xor U7085 (N_7085,N_6909,N_6638);
and U7086 (N_7086,N_6982,N_6971);
nand U7087 (N_7087,N_6509,N_6661);
nand U7088 (N_7088,N_6563,N_6861);
and U7089 (N_7089,N_6718,N_6616);
nand U7090 (N_7090,N_6712,N_6866);
or U7091 (N_7091,N_6724,N_6778);
xnor U7092 (N_7092,N_6834,N_6634);
nor U7093 (N_7093,N_6709,N_6688);
xor U7094 (N_7094,N_6747,N_6823);
nand U7095 (N_7095,N_6601,N_6850);
nor U7096 (N_7096,N_6902,N_6770);
and U7097 (N_7097,N_6944,N_6731);
or U7098 (N_7098,N_6599,N_6941);
nand U7099 (N_7099,N_6586,N_6735);
nand U7100 (N_7100,N_6551,N_6651);
nand U7101 (N_7101,N_6745,N_6964);
and U7102 (N_7102,N_6846,N_6631);
nor U7103 (N_7103,N_6764,N_6699);
nand U7104 (N_7104,N_6817,N_6502);
nor U7105 (N_7105,N_6790,N_6759);
nand U7106 (N_7106,N_6505,N_6674);
xor U7107 (N_7107,N_6519,N_6640);
and U7108 (N_7108,N_6732,N_6931);
xnor U7109 (N_7109,N_6539,N_6729);
or U7110 (N_7110,N_6679,N_6969);
and U7111 (N_7111,N_6542,N_6957);
and U7112 (N_7112,N_6972,N_6918);
nor U7113 (N_7113,N_6532,N_6807);
nand U7114 (N_7114,N_6516,N_6664);
xnor U7115 (N_7115,N_6758,N_6998);
nor U7116 (N_7116,N_6669,N_6515);
nor U7117 (N_7117,N_6607,N_6988);
or U7118 (N_7118,N_6953,N_6520);
or U7119 (N_7119,N_6624,N_6569);
nand U7120 (N_7120,N_6892,N_6913);
xnor U7121 (N_7121,N_6722,N_6837);
nand U7122 (N_7122,N_6831,N_6635);
xor U7123 (N_7123,N_6877,N_6592);
and U7124 (N_7124,N_6996,N_6942);
xor U7125 (N_7125,N_6811,N_6917);
xor U7126 (N_7126,N_6619,N_6596);
or U7127 (N_7127,N_6934,N_6816);
xnor U7128 (N_7128,N_6594,N_6572);
nand U7129 (N_7129,N_6508,N_6750);
xnor U7130 (N_7130,N_6687,N_6528);
or U7131 (N_7131,N_6870,N_6994);
nand U7132 (N_7132,N_6795,N_6812);
and U7133 (N_7133,N_6582,N_6769);
and U7134 (N_7134,N_6501,N_6678);
nand U7135 (N_7135,N_6989,N_6828);
nand U7136 (N_7136,N_6523,N_6864);
nand U7137 (N_7137,N_6956,N_6852);
nor U7138 (N_7138,N_6727,N_6912);
and U7139 (N_7139,N_6858,N_6853);
nand U7140 (N_7140,N_6580,N_6618);
and U7141 (N_7141,N_6781,N_6684);
nand U7142 (N_7142,N_6540,N_6694);
or U7143 (N_7143,N_6889,N_6801);
nor U7144 (N_7144,N_6786,N_6843);
and U7145 (N_7145,N_6923,N_6665);
and U7146 (N_7146,N_6915,N_6726);
xor U7147 (N_7147,N_6847,N_6813);
and U7148 (N_7148,N_6656,N_6683);
xnor U7149 (N_7149,N_6895,N_6789);
nor U7150 (N_7150,N_6728,N_6713);
nand U7151 (N_7151,N_6886,N_6662);
xnor U7152 (N_7152,N_6507,N_6693);
or U7153 (N_7153,N_6737,N_6545);
and U7154 (N_7154,N_6636,N_6783);
nand U7155 (N_7155,N_6985,N_6589);
xor U7156 (N_7156,N_6830,N_6741);
nor U7157 (N_7157,N_6646,N_6714);
xor U7158 (N_7158,N_6657,N_6762);
nor U7159 (N_7159,N_6633,N_6655);
xnor U7160 (N_7160,N_6840,N_6654);
nor U7161 (N_7161,N_6782,N_6927);
or U7162 (N_7162,N_6597,N_6881);
or U7163 (N_7163,N_6623,N_6835);
and U7164 (N_7164,N_6873,N_6500);
and U7165 (N_7165,N_6530,N_6757);
or U7166 (N_7166,N_6904,N_6685);
nor U7167 (N_7167,N_6803,N_6897);
nand U7168 (N_7168,N_6948,N_6975);
xor U7169 (N_7169,N_6773,N_6753);
or U7170 (N_7170,N_6621,N_6697);
nand U7171 (N_7171,N_6744,N_6905);
or U7172 (N_7172,N_6650,N_6730);
nand U7173 (N_7173,N_6865,N_6951);
xnor U7174 (N_7174,N_6611,N_6617);
xnor U7175 (N_7175,N_6829,N_6979);
nand U7176 (N_7176,N_6708,N_6644);
xor U7177 (N_7177,N_6630,N_6626);
and U7178 (N_7178,N_6711,N_6968);
nand U7179 (N_7179,N_6901,N_6725);
nand U7180 (N_7180,N_6639,N_6959);
nor U7181 (N_7181,N_6995,N_6962);
nand U7182 (N_7182,N_6748,N_6863);
or U7183 (N_7183,N_6588,N_6564);
xnor U7184 (N_7184,N_6977,N_6653);
xor U7185 (N_7185,N_6950,N_6716);
and U7186 (N_7186,N_6562,N_6652);
or U7187 (N_7187,N_6754,N_6756);
and U7188 (N_7188,N_6645,N_6567);
and U7189 (N_7189,N_6548,N_6736);
nor U7190 (N_7190,N_6557,N_6543);
and U7191 (N_7191,N_6945,N_6799);
nand U7192 (N_7192,N_6610,N_6675);
nor U7193 (N_7193,N_6555,N_6806);
and U7194 (N_7194,N_6872,N_6517);
nand U7195 (N_7195,N_6860,N_6755);
nand U7196 (N_7196,N_6976,N_6568);
xnor U7197 (N_7197,N_6573,N_6947);
or U7198 (N_7198,N_6926,N_6676);
or U7199 (N_7199,N_6849,N_6949);
or U7200 (N_7200,N_6888,N_6967);
xnor U7201 (N_7201,N_6785,N_6680);
and U7202 (N_7202,N_6784,N_6681);
nand U7203 (N_7203,N_6723,N_6857);
or U7204 (N_7204,N_6907,N_6883);
or U7205 (N_7205,N_6938,N_6965);
and U7206 (N_7206,N_6780,N_6851);
or U7207 (N_7207,N_6910,N_6608);
nor U7208 (N_7208,N_6885,N_6700);
nor U7209 (N_7209,N_6963,N_6600);
or U7210 (N_7210,N_6527,N_6916);
or U7211 (N_7211,N_6820,N_6862);
and U7212 (N_7212,N_6535,N_6524);
nor U7213 (N_7213,N_6958,N_6581);
or U7214 (N_7214,N_6536,N_6628);
nand U7215 (N_7215,N_6798,N_6598);
nor U7216 (N_7216,N_6673,N_6808);
nor U7217 (N_7217,N_6584,N_6815);
nor U7218 (N_7218,N_6738,N_6940);
nand U7219 (N_7219,N_6793,N_6765);
xor U7220 (N_7220,N_6525,N_6983);
and U7221 (N_7221,N_6625,N_6952);
nor U7222 (N_7222,N_6648,N_6869);
or U7223 (N_7223,N_6978,N_6763);
and U7224 (N_7224,N_6809,N_6622);
or U7225 (N_7225,N_6914,N_6890);
nand U7226 (N_7226,N_6740,N_6774);
xnor U7227 (N_7227,N_6787,N_6671);
xor U7228 (N_7228,N_6936,N_6943);
xnor U7229 (N_7229,N_6579,N_6751);
nor U7230 (N_7230,N_6911,N_6752);
or U7231 (N_7231,N_6554,N_6833);
and U7232 (N_7232,N_6570,N_6984);
nor U7233 (N_7233,N_6593,N_6903);
and U7234 (N_7234,N_6698,N_6576);
nor U7235 (N_7235,N_6552,N_6531);
and U7236 (N_7236,N_6701,N_6695);
xor U7237 (N_7237,N_6788,N_6810);
or U7238 (N_7238,N_6836,N_6637);
nor U7239 (N_7239,N_6546,N_6832);
nand U7240 (N_7240,N_6954,N_6818);
or U7241 (N_7241,N_6559,N_6717);
nand U7242 (N_7242,N_6856,N_6660);
xnor U7243 (N_7243,N_6893,N_6561);
nand U7244 (N_7244,N_6966,N_6577);
and U7245 (N_7245,N_6606,N_6575);
nand U7246 (N_7246,N_6578,N_6615);
or U7247 (N_7247,N_6929,N_6791);
nand U7248 (N_7248,N_6900,N_6986);
and U7249 (N_7249,N_6973,N_6844);
and U7250 (N_7250,N_6732,N_6646);
xor U7251 (N_7251,N_6790,N_6882);
nand U7252 (N_7252,N_6956,N_6729);
xnor U7253 (N_7253,N_6520,N_6531);
or U7254 (N_7254,N_6706,N_6810);
and U7255 (N_7255,N_6752,N_6764);
xor U7256 (N_7256,N_6748,N_6604);
nor U7257 (N_7257,N_6684,N_6915);
and U7258 (N_7258,N_6967,N_6927);
and U7259 (N_7259,N_6589,N_6808);
nor U7260 (N_7260,N_6575,N_6964);
and U7261 (N_7261,N_6611,N_6797);
nor U7262 (N_7262,N_6757,N_6536);
nand U7263 (N_7263,N_6651,N_6785);
or U7264 (N_7264,N_6753,N_6594);
nand U7265 (N_7265,N_6786,N_6542);
and U7266 (N_7266,N_6740,N_6859);
or U7267 (N_7267,N_6875,N_6661);
xnor U7268 (N_7268,N_6962,N_6979);
nor U7269 (N_7269,N_6562,N_6929);
nor U7270 (N_7270,N_6535,N_6537);
xnor U7271 (N_7271,N_6972,N_6832);
and U7272 (N_7272,N_6721,N_6529);
nor U7273 (N_7273,N_6611,N_6862);
nand U7274 (N_7274,N_6992,N_6873);
nand U7275 (N_7275,N_6991,N_6593);
nor U7276 (N_7276,N_6562,N_6761);
and U7277 (N_7277,N_6719,N_6681);
nor U7278 (N_7278,N_6901,N_6748);
or U7279 (N_7279,N_6686,N_6878);
nand U7280 (N_7280,N_6762,N_6614);
and U7281 (N_7281,N_6872,N_6515);
or U7282 (N_7282,N_6704,N_6930);
xnor U7283 (N_7283,N_6920,N_6702);
and U7284 (N_7284,N_6976,N_6780);
or U7285 (N_7285,N_6516,N_6707);
and U7286 (N_7286,N_6857,N_6606);
and U7287 (N_7287,N_6702,N_6875);
xnor U7288 (N_7288,N_6609,N_6941);
or U7289 (N_7289,N_6972,N_6584);
xor U7290 (N_7290,N_6905,N_6593);
xor U7291 (N_7291,N_6963,N_6791);
nor U7292 (N_7292,N_6927,N_6744);
xor U7293 (N_7293,N_6862,N_6587);
nand U7294 (N_7294,N_6611,N_6874);
and U7295 (N_7295,N_6720,N_6610);
nor U7296 (N_7296,N_6525,N_6795);
nand U7297 (N_7297,N_6843,N_6864);
or U7298 (N_7298,N_6551,N_6590);
nand U7299 (N_7299,N_6671,N_6829);
or U7300 (N_7300,N_6825,N_6559);
nor U7301 (N_7301,N_6535,N_6646);
xnor U7302 (N_7302,N_6551,N_6531);
and U7303 (N_7303,N_6915,N_6811);
nand U7304 (N_7304,N_6682,N_6703);
nor U7305 (N_7305,N_6588,N_6692);
nor U7306 (N_7306,N_6762,N_6649);
xnor U7307 (N_7307,N_6687,N_6928);
nand U7308 (N_7308,N_6733,N_6898);
or U7309 (N_7309,N_6721,N_6613);
nor U7310 (N_7310,N_6532,N_6846);
or U7311 (N_7311,N_6608,N_6900);
and U7312 (N_7312,N_6628,N_6799);
or U7313 (N_7313,N_6594,N_6720);
or U7314 (N_7314,N_6583,N_6762);
and U7315 (N_7315,N_6922,N_6919);
nand U7316 (N_7316,N_6611,N_6579);
or U7317 (N_7317,N_6576,N_6988);
nand U7318 (N_7318,N_6944,N_6834);
nand U7319 (N_7319,N_6681,N_6607);
nor U7320 (N_7320,N_6737,N_6889);
nor U7321 (N_7321,N_6896,N_6608);
and U7322 (N_7322,N_6604,N_6866);
nor U7323 (N_7323,N_6682,N_6537);
nand U7324 (N_7324,N_6530,N_6559);
and U7325 (N_7325,N_6757,N_6904);
or U7326 (N_7326,N_6929,N_6504);
nor U7327 (N_7327,N_6843,N_6675);
and U7328 (N_7328,N_6776,N_6693);
nor U7329 (N_7329,N_6755,N_6568);
nor U7330 (N_7330,N_6752,N_6653);
xnor U7331 (N_7331,N_6900,N_6993);
and U7332 (N_7332,N_6670,N_6516);
nand U7333 (N_7333,N_6533,N_6898);
nor U7334 (N_7334,N_6948,N_6751);
xnor U7335 (N_7335,N_6657,N_6514);
nand U7336 (N_7336,N_6957,N_6776);
xnor U7337 (N_7337,N_6502,N_6805);
or U7338 (N_7338,N_6763,N_6510);
nand U7339 (N_7339,N_6853,N_6852);
nand U7340 (N_7340,N_6865,N_6734);
and U7341 (N_7341,N_6793,N_6615);
nor U7342 (N_7342,N_6651,N_6655);
and U7343 (N_7343,N_6516,N_6919);
or U7344 (N_7344,N_6515,N_6581);
or U7345 (N_7345,N_6867,N_6518);
xor U7346 (N_7346,N_6875,N_6792);
nor U7347 (N_7347,N_6672,N_6878);
nand U7348 (N_7348,N_6923,N_6833);
nand U7349 (N_7349,N_6561,N_6897);
or U7350 (N_7350,N_6976,N_6575);
nand U7351 (N_7351,N_6726,N_6667);
xor U7352 (N_7352,N_6581,N_6833);
nor U7353 (N_7353,N_6674,N_6504);
nor U7354 (N_7354,N_6586,N_6801);
and U7355 (N_7355,N_6962,N_6672);
or U7356 (N_7356,N_6837,N_6965);
nand U7357 (N_7357,N_6791,N_6905);
nand U7358 (N_7358,N_6838,N_6992);
or U7359 (N_7359,N_6703,N_6909);
nor U7360 (N_7360,N_6704,N_6936);
and U7361 (N_7361,N_6847,N_6749);
or U7362 (N_7362,N_6593,N_6706);
nor U7363 (N_7363,N_6547,N_6582);
and U7364 (N_7364,N_6921,N_6772);
nor U7365 (N_7365,N_6775,N_6931);
nor U7366 (N_7366,N_6737,N_6664);
or U7367 (N_7367,N_6786,N_6868);
xor U7368 (N_7368,N_6648,N_6782);
nor U7369 (N_7369,N_6979,N_6970);
xor U7370 (N_7370,N_6673,N_6774);
or U7371 (N_7371,N_6563,N_6604);
xnor U7372 (N_7372,N_6522,N_6695);
xnor U7373 (N_7373,N_6661,N_6550);
or U7374 (N_7374,N_6740,N_6772);
xor U7375 (N_7375,N_6778,N_6803);
xnor U7376 (N_7376,N_6680,N_6537);
and U7377 (N_7377,N_6652,N_6603);
nor U7378 (N_7378,N_6591,N_6530);
xor U7379 (N_7379,N_6778,N_6577);
nand U7380 (N_7380,N_6904,N_6599);
or U7381 (N_7381,N_6950,N_6914);
and U7382 (N_7382,N_6608,N_6556);
or U7383 (N_7383,N_6586,N_6610);
or U7384 (N_7384,N_6935,N_6650);
or U7385 (N_7385,N_6948,N_6972);
nor U7386 (N_7386,N_6547,N_6644);
or U7387 (N_7387,N_6706,N_6633);
nand U7388 (N_7388,N_6832,N_6919);
nand U7389 (N_7389,N_6994,N_6929);
xor U7390 (N_7390,N_6843,N_6729);
xnor U7391 (N_7391,N_6533,N_6770);
nand U7392 (N_7392,N_6803,N_6786);
and U7393 (N_7393,N_6758,N_6971);
nand U7394 (N_7394,N_6897,N_6973);
nor U7395 (N_7395,N_6671,N_6934);
or U7396 (N_7396,N_6714,N_6702);
or U7397 (N_7397,N_6867,N_6763);
xnor U7398 (N_7398,N_6767,N_6682);
nand U7399 (N_7399,N_6747,N_6842);
nor U7400 (N_7400,N_6659,N_6945);
nor U7401 (N_7401,N_6797,N_6766);
nor U7402 (N_7402,N_6698,N_6506);
or U7403 (N_7403,N_6940,N_6505);
xnor U7404 (N_7404,N_6517,N_6971);
or U7405 (N_7405,N_6988,N_6577);
xnor U7406 (N_7406,N_6953,N_6675);
xor U7407 (N_7407,N_6956,N_6515);
nand U7408 (N_7408,N_6830,N_6767);
or U7409 (N_7409,N_6887,N_6747);
and U7410 (N_7410,N_6965,N_6984);
and U7411 (N_7411,N_6860,N_6601);
or U7412 (N_7412,N_6769,N_6804);
nand U7413 (N_7413,N_6677,N_6921);
nand U7414 (N_7414,N_6604,N_6993);
or U7415 (N_7415,N_6843,N_6962);
nor U7416 (N_7416,N_6856,N_6879);
xnor U7417 (N_7417,N_6743,N_6836);
xor U7418 (N_7418,N_6926,N_6520);
nand U7419 (N_7419,N_6978,N_6807);
nand U7420 (N_7420,N_6971,N_6654);
or U7421 (N_7421,N_6636,N_6505);
and U7422 (N_7422,N_6565,N_6535);
and U7423 (N_7423,N_6619,N_6661);
nor U7424 (N_7424,N_6734,N_6559);
nor U7425 (N_7425,N_6524,N_6544);
nand U7426 (N_7426,N_6840,N_6526);
and U7427 (N_7427,N_6911,N_6742);
xor U7428 (N_7428,N_6629,N_6641);
xnor U7429 (N_7429,N_6906,N_6502);
nand U7430 (N_7430,N_6681,N_6708);
xnor U7431 (N_7431,N_6638,N_6563);
and U7432 (N_7432,N_6550,N_6532);
nor U7433 (N_7433,N_6675,N_6592);
or U7434 (N_7434,N_6522,N_6952);
nor U7435 (N_7435,N_6990,N_6850);
xnor U7436 (N_7436,N_6987,N_6582);
or U7437 (N_7437,N_6856,N_6591);
nor U7438 (N_7438,N_6908,N_6514);
and U7439 (N_7439,N_6702,N_6926);
and U7440 (N_7440,N_6880,N_6763);
nand U7441 (N_7441,N_6851,N_6739);
nor U7442 (N_7442,N_6907,N_6716);
nand U7443 (N_7443,N_6615,N_6819);
nor U7444 (N_7444,N_6721,N_6846);
and U7445 (N_7445,N_6911,N_6626);
and U7446 (N_7446,N_6532,N_6879);
and U7447 (N_7447,N_6879,N_6554);
and U7448 (N_7448,N_6655,N_6739);
and U7449 (N_7449,N_6925,N_6828);
or U7450 (N_7450,N_6968,N_6962);
nand U7451 (N_7451,N_6543,N_6565);
nand U7452 (N_7452,N_6868,N_6572);
or U7453 (N_7453,N_6782,N_6739);
xnor U7454 (N_7454,N_6756,N_6658);
or U7455 (N_7455,N_6665,N_6914);
or U7456 (N_7456,N_6674,N_6586);
nand U7457 (N_7457,N_6685,N_6671);
nand U7458 (N_7458,N_6541,N_6911);
and U7459 (N_7459,N_6959,N_6773);
nor U7460 (N_7460,N_6929,N_6891);
or U7461 (N_7461,N_6642,N_6944);
and U7462 (N_7462,N_6544,N_6581);
and U7463 (N_7463,N_6969,N_6899);
xnor U7464 (N_7464,N_6909,N_6962);
and U7465 (N_7465,N_6852,N_6829);
or U7466 (N_7466,N_6912,N_6921);
and U7467 (N_7467,N_6582,N_6847);
xor U7468 (N_7468,N_6906,N_6981);
nor U7469 (N_7469,N_6995,N_6987);
nand U7470 (N_7470,N_6626,N_6643);
nor U7471 (N_7471,N_6661,N_6834);
or U7472 (N_7472,N_6648,N_6849);
nor U7473 (N_7473,N_6813,N_6874);
or U7474 (N_7474,N_6947,N_6669);
nand U7475 (N_7475,N_6912,N_6549);
nand U7476 (N_7476,N_6512,N_6607);
or U7477 (N_7477,N_6596,N_6862);
nand U7478 (N_7478,N_6663,N_6887);
nand U7479 (N_7479,N_6704,N_6695);
xor U7480 (N_7480,N_6738,N_6862);
and U7481 (N_7481,N_6959,N_6622);
nor U7482 (N_7482,N_6519,N_6928);
nor U7483 (N_7483,N_6631,N_6843);
or U7484 (N_7484,N_6782,N_6524);
xor U7485 (N_7485,N_6707,N_6592);
and U7486 (N_7486,N_6927,N_6614);
or U7487 (N_7487,N_6740,N_6999);
or U7488 (N_7488,N_6894,N_6863);
or U7489 (N_7489,N_6561,N_6933);
or U7490 (N_7490,N_6746,N_6726);
nor U7491 (N_7491,N_6854,N_6523);
and U7492 (N_7492,N_6881,N_6653);
nor U7493 (N_7493,N_6506,N_6608);
nand U7494 (N_7494,N_6914,N_6876);
and U7495 (N_7495,N_6935,N_6563);
nor U7496 (N_7496,N_6752,N_6650);
nand U7497 (N_7497,N_6816,N_6780);
nand U7498 (N_7498,N_6884,N_6561);
and U7499 (N_7499,N_6876,N_6983);
or U7500 (N_7500,N_7226,N_7310);
xor U7501 (N_7501,N_7389,N_7448);
or U7502 (N_7502,N_7461,N_7081);
or U7503 (N_7503,N_7265,N_7267);
and U7504 (N_7504,N_7090,N_7318);
nand U7505 (N_7505,N_7385,N_7337);
nand U7506 (N_7506,N_7434,N_7296);
or U7507 (N_7507,N_7281,N_7011);
nand U7508 (N_7508,N_7051,N_7348);
nand U7509 (N_7509,N_7366,N_7167);
nand U7510 (N_7510,N_7333,N_7047);
or U7511 (N_7511,N_7153,N_7311);
nand U7512 (N_7512,N_7415,N_7041);
xnor U7513 (N_7513,N_7354,N_7302);
nor U7514 (N_7514,N_7493,N_7305);
xnor U7515 (N_7515,N_7183,N_7314);
or U7516 (N_7516,N_7382,N_7228);
nand U7517 (N_7517,N_7322,N_7138);
nor U7518 (N_7518,N_7271,N_7362);
nand U7519 (N_7519,N_7101,N_7156);
nand U7520 (N_7520,N_7331,N_7387);
and U7521 (N_7521,N_7490,N_7358);
nand U7522 (N_7522,N_7411,N_7221);
nor U7523 (N_7523,N_7406,N_7476);
nand U7524 (N_7524,N_7313,N_7251);
nor U7525 (N_7525,N_7238,N_7427);
and U7526 (N_7526,N_7008,N_7086);
xor U7527 (N_7527,N_7319,N_7034);
or U7528 (N_7528,N_7105,N_7112);
nand U7529 (N_7529,N_7222,N_7065);
or U7530 (N_7530,N_7037,N_7398);
xor U7531 (N_7531,N_7423,N_7060);
or U7532 (N_7532,N_7437,N_7270);
nor U7533 (N_7533,N_7405,N_7196);
nand U7534 (N_7534,N_7410,N_7005);
nand U7535 (N_7535,N_7071,N_7443);
nand U7536 (N_7536,N_7023,N_7345);
and U7537 (N_7537,N_7424,N_7367);
nand U7538 (N_7538,N_7031,N_7220);
nor U7539 (N_7539,N_7014,N_7022);
xnor U7540 (N_7540,N_7054,N_7492);
or U7541 (N_7541,N_7275,N_7092);
nand U7542 (N_7542,N_7069,N_7045);
or U7543 (N_7543,N_7338,N_7169);
nand U7544 (N_7544,N_7301,N_7203);
and U7545 (N_7545,N_7273,N_7095);
xnor U7546 (N_7546,N_7332,N_7481);
and U7547 (N_7547,N_7441,N_7306);
or U7548 (N_7548,N_7213,N_7312);
or U7549 (N_7549,N_7124,N_7059);
and U7550 (N_7550,N_7375,N_7370);
nor U7551 (N_7551,N_7479,N_7289);
nand U7552 (N_7552,N_7259,N_7297);
or U7553 (N_7553,N_7172,N_7159);
and U7554 (N_7554,N_7413,N_7335);
nand U7555 (N_7555,N_7098,N_7113);
xor U7556 (N_7556,N_7373,N_7082);
nand U7557 (N_7557,N_7119,N_7087);
nand U7558 (N_7558,N_7029,N_7056);
xor U7559 (N_7559,N_7452,N_7173);
nor U7560 (N_7560,N_7132,N_7482);
and U7561 (N_7561,N_7072,N_7147);
and U7562 (N_7562,N_7349,N_7395);
or U7563 (N_7563,N_7309,N_7459);
and U7564 (N_7564,N_7046,N_7036);
xnor U7565 (N_7565,N_7285,N_7280);
or U7566 (N_7566,N_7404,N_7039);
and U7567 (N_7567,N_7073,N_7379);
and U7568 (N_7568,N_7330,N_7080);
xor U7569 (N_7569,N_7152,N_7099);
xor U7570 (N_7570,N_7197,N_7118);
and U7571 (N_7571,N_7383,N_7300);
nor U7572 (N_7572,N_7384,N_7327);
or U7573 (N_7573,N_7177,N_7456);
or U7574 (N_7574,N_7211,N_7494);
and U7575 (N_7575,N_7170,N_7140);
nand U7576 (N_7576,N_7207,N_7006);
nand U7577 (N_7577,N_7368,N_7412);
and U7578 (N_7578,N_7209,N_7279);
nor U7579 (N_7579,N_7121,N_7328);
or U7580 (N_7580,N_7002,N_7290);
and U7581 (N_7581,N_7142,N_7103);
nand U7582 (N_7582,N_7055,N_7214);
and U7583 (N_7583,N_7117,N_7182);
and U7584 (N_7584,N_7438,N_7497);
nand U7585 (N_7585,N_7217,N_7148);
xnor U7586 (N_7586,N_7365,N_7272);
nand U7587 (N_7587,N_7288,N_7409);
nor U7588 (N_7588,N_7179,N_7061);
nor U7589 (N_7589,N_7143,N_7276);
nor U7590 (N_7590,N_7307,N_7012);
or U7591 (N_7591,N_7408,N_7477);
nor U7592 (N_7592,N_7193,N_7052);
or U7593 (N_7593,N_7397,N_7249);
nor U7594 (N_7594,N_7465,N_7115);
or U7595 (N_7595,N_7418,N_7131);
or U7596 (N_7596,N_7336,N_7450);
and U7597 (N_7597,N_7255,N_7346);
or U7598 (N_7598,N_7422,N_7356);
nor U7599 (N_7599,N_7262,N_7100);
nor U7600 (N_7600,N_7198,N_7467);
nand U7601 (N_7601,N_7096,N_7449);
xnor U7602 (N_7602,N_7471,N_7347);
nand U7603 (N_7603,N_7135,N_7453);
xor U7604 (N_7604,N_7257,N_7283);
nor U7605 (N_7605,N_7475,N_7208);
nand U7606 (N_7606,N_7161,N_7205);
xnor U7607 (N_7607,N_7341,N_7430);
xnor U7608 (N_7608,N_7454,N_7303);
nor U7609 (N_7609,N_7234,N_7166);
and U7610 (N_7610,N_7496,N_7458);
xnor U7611 (N_7611,N_7376,N_7308);
nand U7612 (N_7612,N_7067,N_7020);
or U7613 (N_7613,N_7266,N_7015);
or U7614 (N_7614,N_7189,N_7386);
or U7615 (N_7615,N_7457,N_7157);
and U7616 (N_7616,N_7190,N_7292);
and U7617 (N_7617,N_7250,N_7466);
nor U7618 (N_7618,N_7417,N_7446);
and U7619 (N_7619,N_7414,N_7224);
and U7620 (N_7620,N_7455,N_7294);
and U7621 (N_7621,N_7210,N_7261);
nand U7622 (N_7622,N_7218,N_7463);
xor U7623 (N_7623,N_7010,N_7164);
and U7624 (N_7624,N_7488,N_7237);
xnor U7625 (N_7625,N_7146,N_7195);
or U7626 (N_7626,N_7024,N_7174);
or U7627 (N_7627,N_7175,N_7363);
xnor U7628 (N_7628,N_7320,N_7044);
nand U7629 (N_7629,N_7339,N_7304);
or U7630 (N_7630,N_7009,N_7141);
or U7631 (N_7631,N_7013,N_7392);
nor U7632 (N_7632,N_7128,N_7248);
nor U7633 (N_7633,N_7378,N_7487);
or U7634 (N_7634,N_7125,N_7268);
or U7635 (N_7635,N_7160,N_7343);
xnor U7636 (N_7636,N_7106,N_7212);
or U7637 (N_7637,N_7050,N_7016);
xnor U7638 (N_7638,N_7491,N_7102);
nand U7639 (N_7639,N_7394,N_7342);
nand U7640 (N_7640,N_7278,N_7053);
and U7641 (N_7641,N_7233,N_7178);
or U7642 (N_7642,N_7478,N_7400);
nand U7643 (N_7643,N_7380,N_7393);
nor U7644 (N_7644,N_7133,N_7126);
and U7645 (N_7645,N_7240,N_7000);
nor U7646 (N_7646,N_7074,N_7287);
or U7647 (N_7647,N_7019,N_7245);
xnor U7648 (N_7648,N_7084,N_7359);
and U7649 (N_7649,N_7150,N_7277);
xnor U7650 (N_7650,N_7185,N_7246);
nand U7651 (N_7651,N_7078,N_7429);
or U7652 (N_7652,N_7460,N_7035);
nor U7653 (N_7653,N_7326,N_7155);
nor U7654 (N_7654,N_7269,N_7231);
or U7655 (N_7655,N_7192,N_7433);
and U7656 (N_7656,N_7130,N_7079);
or U7657 (N_7657,N_7144,N_7204);
and U7658 (N_7658,N_7134,N_7317);
and U7659 (N_7659,N_7033,N_7447);
nor U7660 (N_7660,N_7091,N_7388);
or U7661 (N_7661,N_7498,N_7236);
nand U7662 (N_7662,N_7371,N_7353);
xnor U7663 (N_7663,N_7361,N_7344);
nand U7664 (N_7664,N_7439,N_7426);
nand U7665 (N_7665,N_7032,N_7049);
xor U7666 (N_7666,N_7484,N_7485);
or U7667 (N_7667,N_7252,N_7176);
or U7668 (N_7668,N_7004,N_7377);
and U7669 (N_7669,N_7390,N_7444);
nor U7670 (N_7670,N_7110,N_7136);
or U7671 (N_7671,N_7070,N_7116);
or U7672 (N_7672,N_7064,N_7263);
xor U7673 (N_7673,N_7445,N_7235);
and U7674 (N_7674,N_7419,N_7191);
nor U7675 (N_7675,N_7139,N_7468);
xnor U7676 (N_7676,N_7089,N_7168);
and U7677 (N_7677,N_7165,N_7122);
xnor U7678 (N_7678,N_7293,N_7282);
nor U7679 (N_7679,N_7489,N_7470);
nor U7680 (N_7680,N_7062,N_7480);
nor U7681 (N_7681,N_7188,N_7027);
or U7682 (N_7682,N_7129,N_7316);
nand U7683 (N_7683,N_7432,N_7396);
nand U7684 (N_7684,N_7184,N_7186);
or U7685 (N_7685,N_7216,N_7352);
nand U7686 (N_7686,N_7180,N_7239);
nand U7687 (N_7687,N_7462,N_7431);
nand U7688 (N_7688,N_7154,N_7374);
nand U7689 (N_7689,N_7017,N_7063);
and U7690 (N_7690,N_7350,N_7127);
xor U7691 (N_7691,N_7123,N_7425);
or U7692 (N_7692,N_7030,N_7324);
or U7693 (N_7693,N_7325,N_7021);
and U7694 (N_7694,N_7025,N_7329);
nor U7695 (N_7695,N_7120,N_7472);
xor U7696 (N_7696,N_7007,N_7038);
nand U7697 (N_7697,N_7003,N_7299);
and U7698 (N_7698,N_7474,N_7321);
and U7699 (N_7699,N_7093,N_7094);
or U7700 (N_7700,N_7284,N_7372);
and U7701 (N_7701,N_7088,N_7163);
nand U7702 (N_7702,N_7215,N_7149);
xnor U7703 (N_7703,N_7158,N_7264);
and U7704 (N_7704,N_7421,N_7436);
and U7705 (N_7705,N_7440,N_7181);
and U7706 (N_7706,N_7058,N_7085);
nand U7707 (N_7707,N_7162,N_7243);
xor U7708 (N_7708,N_7247,N_7401);
nand U7709 (N_7709,N_7223,N_7355);
xor U7710 (N_7710,N_7076,N_7416);
nand U7711 (N_7711,N_7253,N_7286);
nor U7712 (N_7712,N_7403,N_7048);
and U7713 (N_7713,N_7254,N_7230);
nor U7714 (N_7714,N_7428,N_7258);
xnor U7715 (N_7715,N_7200,N_7360);
and U7716 (N_7716,N_7018,N_7227);
nor U7717 (N_7717,N_7114,N_7225);
or U7718 (N_7718,N_7402,N_7334);
and U7719 (N_7719,N_7351,N_7369);
or U7720 (N_7720,N_7256,N_7137);
nand U7721 (N_7721,N_7042,N_7083);
nor U7722 (N_7722,N_7242,N_7028);
or U7723 (N_7723,N_7219,N_7097);
or U7724 (N_7724,N_7001,N_7499);
or U7725 (N_7725,N_7464,N_7295);
nor U7726 (N_7726,N_7066,N_7068);
xnor U7727 (N_7727,N_7043,N_7111);
or U7728 (N_7728,N_7435,N_7202);
and U7729 (N_7729,N_7315,N_7206);
xor U7730 (N_7730,N_7407,N_7108);
or U7731 (N_7731,N_7145,N_7323);
or U7732 (N_7732,N_7229,N_7075);
nor U7733 (N_7733,N_7340,N_7495);
or U7734 (N_7734,N_7241,N_7260);
nand U7735 (N_7735,N_7077,N_7420);
and U7736 (N_7736,N_7469,N_7473);
xor U7737 (N_7737,N_7199,N_7357);
nand U7738 (N_7738,N_7298,N_7232);
nand U7739 (N_7739,N_7399,N_7171);
nor U7740 (N_7740,N_7381,N_7486);
nor U7741 (N_7741,N_7483,N_7187);
and U7742 (N_7742,N_7244,N_7291);
nor U7743 (N_7743,N_7107,N_7364);
nor U7744 (N_7744,N_7040,N_7194);
nand U7745 (N_7745,N_7026,N_7201);
nand U7746 (N_7746,N_7104,N_7109);
and U7747 (N_7747,N_7151,N_7274);
and U7748 (N_7748,N_7057,N_7391);
nor U7749 (N_7749,N_7451,N_7442);
nor U7750 (N_7750,N_7211,N_7149);
and U7751 (N_7751,N_7473,N_7124);
nand U7752 (N_7752,N_7035,N_7295);
xnor U7753 (N_7753,N_7466,N_7219);
or U7754 (N_7754,N_7067,N_7243);
and U7755 (N_7755,N_7126,N_7164);
nor U7756 (N_7756,N_7173,N_7240);
nand U7757 (N_7757,N_7478,N_7248);
and U7758 (N_7758,N_7287,N_7443);
nor U7759 (N_7759,N_7407,N_7128);
nand U7760 (N_7760,N_7301,N_7053);
and U7761 (N_7761,N_7110,N_7173);
or U7762 (N_7762,N_7311,N_7078);
nand U7763 (N_7763,N_7282,N_7426);
and U7764 (N_7764,N_7220,N_7290);
xnor U7765 (N_7765,N_7368,N_7180);
nand U7766 (N_7766,N_7325,N_7447);
xor U7767 (N_7767,N_7135,N_7031);
and U7768 (N_7768,N_7155,N_7301);
or U7769 (N_7769,N_7385,N_7406);
or U7770 (N_7770,N_7262,N_7227);
nand U7771 (N_7771,N_7209,N_7436);
or U7772 (N_7772,N_7284,N_7270);
xor U7773 (N_7773,N_7373,N_7068);
nand U7774 (N_7774,N_7471,N_7310);
nand U7775 (N_7775,N_7453,N_7029);
nor U7776 (N_7776,N_7354,N_7313);
and U7777 (N_7777,N_7077,N_7483);
and U7778 (N_7778,N_7265,N_7381);
xnor U7779 (N_7779,N_7089,N_7311);
nor U7780 (N_7780,N_7311,N_7334);
and U7781 (N_7781,N_7107,N_7137);
or U7782 (N_7782,N_7359,N_7312);
and U7783 (N_7783,N_7487,N_7407);
or U7784 (N_7784,N_7484,N_7340);
nor U7785 (N_7785,N_7464,N_7250);
nor U7786 (N_7786,N_7323,N_7464);
or U7787 (N_7787,N_7005,N_7379);
xor U7788 (N_7788,N_7203,N_7106);
and U7789 (N_7789,N_7285,N_7440);
or U7790 (N_7790,N_7161,N_7338);
nor U7791 (N_7791,N_7046,N_7347);
xor U7792 (N_7792,N_7250,N_7123);
and U7793 (N_7793,N_7145,N_7048);
nor U7794 (N_7794,N_7395,N_7323);
or U7795 (N_7795,N_7451,N_7385);
and U7796 (N_7796,N_7379,N_7306);
xnor U7797 (N_7797,N_7023,N_7452);
or U7798 (N_7798,N_7237,N_7145);
xor U7799 (N_7799,N_7276,N_7051);
xor U7800 (N_7800,N_7460,N_7041);
nor U7801 (N_7801,N_7322,N_7098);
nand U7802 (N_7802,N_7411,N_7266);
nand U7803 (N_7803,N_7006,N_7171);
and U7804 (N_7804,N_7209,N_7061);
and U7805 (N_7805,N_7467,N_7139);
or U7806 (N_7806,N_7244,N_7211);
xnor U7807 (N_7807,N_7417,N_7231);
nand U7808 (N_7808,N_7177,N_7024);
xor U7809 (N_7809,N_7354,N_7352);
and U7810 (N_7810,N_7023,N_7230);
xnor U7811 (N_7811,N_7076,N_7374);
or U7812 (N_7812,N_7352,N_7198);
nor U7813 (N_7813,N_7008,N_7404);
xnor U7814 (N_7814,N_7487,N_7071);
nor U7815 (N_7815,N_7097,N_7169);
nor U7816 (N_7816,N_7137,N_7241);
nor U7817 (N_7817,N_7405,N_7495);
xnor U7818 (N_7818,N_7391,N_7386);
nor U7819 (N_7819,N_7477,N_7172);
xor U7820 (N_7820,N_7317,N_7198);
nor U7821 (N_7821,N_7391,N_7354);
xor U7822 (N_7822,N_7477,N_7370);
or U7823 (N_7823,N_7154,N_7004);
and U7824 (N_7824,N_7374,N_7311);
and U7825 (N_7825,N_7302,N_7096);
or U7826 (N_7826,N_7040,N_7146);
or U7827 (N_7827,N_7280,N_7433);
xnor U7828 (N_7828,N_7433,N_7383);
nor U7829 (N_7829,N_7006,N_7038);
nand U7830 (N_7830,N_7261,N_7242);
nand U7831 (N_7831,N_7070,N_7325);
xnor U7832 (N_7832,N_7336,N_7249);
and U7833 (N_7833,N_7459,N_7212);
xor U7834 (N_7834,N_7085,N_7187);
or U7835 (N_7835,N_7052,N_7331);
or U7836 (N_7836,N_7127,N_7189);
nand U7837 (N_7837,N_7260,N_7495);
nor U7838 (N_7838,N_7372,N_7439);
and U7839 (N_7839,N_7134,N_7265);
xor U7840 (N_7840,N_7473,N_7149);
or U7841 (N_7841,N_7477,N_7126);
nand U7842 (N_7842,N_7278,N_7128);
nor U7843 (N_7843,N_7267,N_7461);
xor U7844 (N_7844,N_7275,N_7113);
nand U7845 (N_7845,N_7118,N_7296);
and U7846 (N_7846,N_7205,N_7361);
nand U7847 (N_7847,N_7120,N_7387);
and U7848 (N_7848,N_7344,N_7052);
nor U7849 (N_7849,N_7340,N_7164);
xnor U7850 (N_7850,N_7022,N_7000);
and U7851 (N_7851,N_7478,N_7323);
nand U7852 (N_7852,N_7436,N_7176);
and U7853 (N_7853,N_7184,N_7422);
nor U7854 (N_7854,N_7171,N_7374);
nor U7855 (N_7855,N_7093,N_7279);
or U7856 (N_7856,N_7132,N_7212);
nor U7857 (N_7857,N_7389,N_7496);
and U7858 (N_7858,N_7399,N_7013);
nand U7859 (N_7859,N_7171,N_7182);
xnor U7860 (N_7860,N_7171,N_7391);
xnor U7861 (N_7861,N_7381,N_7495);
xor U7862 (N_7862,N_7492,N_7279);
and U7863 (N_7863,N_7431,N_7195);
or U7864 (N_7864,N_7303,N_7100);
xor U7865 (N_7865,N_7313,N_7327);
and U7866 (N_7866,N_7464,N_7351);
xor U7867 (N_7867,N_7156,N_7206);
nor U7868 (N_7868,N_7219,N_7216);
and U7869 (N_7869,N_7160,N_7263);
or U7870 (N_7870,N_7013,N_7409);
and U7871 (N_7871,N_7323,N_7219);
xor U7872 (N_7872,N_7125,N_7447);
nand U7873 (N_7873,N_7064,N_7194);
nand U7874 (N_7874,N_7456,N_7095);
and U7875 (N_7875,N_7265,N_7427);
nor U7876 (N_7876,N_7393,N_7172);
or U7877 (N_7877,N_7205,N_7420);
or U7878 (N_7878,N_7486,N_7298);
nand U7879 (N_7879,N_7445,N_7416);
nand U7880 (N_7880,N_7317,N_7227);
or U7881 (N_7881,N_7083,N_7451);
or U7882 (N_7882,N_7216,N_7292);
nor U7883 (N_7883,N_7434,N_7117);
or U7884 (N_7884,N_7474,N_7486);
xnor U7885 (N_7885,N_7161,N_7474);
and U7886 (N_7886,N_7337,N_7291);
or U7887 (N_7887,N_7266,N_7187);
or U7888 (N_7888,N_7221,N_7407);
xor U7889 (N_7889,N_7274,N_7191);
nand U7890 (N_7890,N_7370,N_7083);
xor U7891 (N_7891,N_7335,N_7085);
and U7892 (N_7892,N_7356,N_7424);
xor U7893 (N_7893,N_7024,N_7003);
nand U7894 (N_7894,N_7216,N_7119);
nor U7895 (N_7895,N_7382,N_7362);
nor U7896 (N_7896,N_7403,N_7022);
or U7897 (N_7897,N_7310,N_7412);
nor U7898 (N_7898,N_7342,N_7100);
and U7899 (N_7899,N_7169,N_7118);
xnor U7900 (N_7900,N_7305,N_7455);
nor U7901 (N_7901,N_7045,N_7066);
and U7902 (N_7902,N_7405,N_7281);
nor U7903 (N_7903,N_7450,N_7211);
nor U7904 (N_7904,N_7439,N_7202);
and U7905 (N_7905,N_7189,N_7269);
and U7906 (N_7906,N_7116,N_7419);
and U7907 (N_7907,N_7327,N_7460);
nor U7908 (N_7908,N_7473,N_7150);
and U7909 (N_7909,N_7301,N_7224);
or U7910 (N_7910,N_7358,N_7198);
xnor U7911 (N_7911,N_7286,N_7265);
nor U7912 (N_7912,N_7184,N_7487);
or U7913 (N_7913,N_7499,N_7105);
or U7914 (N_7914,N_7437,N_7347);
xnor U7915 (N_7915,N_7359,N_7255);
nand U7916 (N_7916,N_7472,N_7038);
xor U7917 (N_7917,N_7062,N_7254);
and U7918 (N_7918,N_7246,N_7454);
xor U7919 (N_7919,N_7036,N_7137);
xor U7920 (N_7920,N_7042,N_7061);
nand U7921 (N_7921,N_7394,N_7371);
and U7922 (N_7922,N_7214,N_7205);
and U7923 (N_7923,N_7056,N_7024);
xor U7924 (N_7924,N_7148,N_7145);
nor U7925 (N_7925,N_7338,N_7157);
xnor U7926 (N_7926,N_7419,N_7082);
nor U7927 (N_7927,N_7144,N_7349);
xnor U7928 (N_7928,N_7171,N_7393);
xnor U7929 (N_7929,N_7312,N_7025);
nor U7930 (N_7930,N_7037,N_7429);
and U7931 (N_7931,N_7308,N_7080);
nand U7932 (N_7932,N_7185,N_7191);
and U7933 (N_7933,N_7479,N_7368);
and U7934 (N_7934,N_7058,N_7364);
xor U7935 (N_7935,N_7402,N_7157);
or U7936 (N_7936,N_7230,N_7458);
and U7937 (N_7937,N_7258,N_7138);
nor U7938 (N_7938,N_7311,N_7057);
or U7939 (N_7939,N_7458,N_7338);
or U7940 (N_7940,N_7278,N_7367);
nor U7941 (N_7941,N_7089,N_7109);
nor U7942 (N_7942,N_7229,N_7264);
and U7943 (N_7943,N_7210,N_7111);
or U7944 (N_7944,N_7232,N_7403);
nand U7945 (N_7945,N_7446,N_7378);
or U7946 (N_7946,N_7041,N_7470);
nor U7947 (N_7947,N_7111,N_7102);
xor U7948 (N_7948,N_7022,N_7209);
or U7949 (N_7949,N_7103,N_7489);
xor U7950 (N_7950,N_7320,N_7079);
xnor U7951 (N_7951,N_7414,N_7284);
xnor U7952 (N_7952,N_7126,N_7158);
xor U7953 (N_7953,N_7344,N_7472);
nor U7954 (N_7954,N_7346,N_7342);
nor U7955 (N_7955,N_7170,N_7111);
nand U7956 (N_7956,N_7317,N_7184);
xnor U7957 (N_7957,N_7438,N_7222);
or U7958 (N_7958,N_7099,N_7278);
and U7959 (N_7959,N_7308,N_7217);
or U7960 (N_7960,N_7474,N_7388);
nor U7961 (N_7961,N_7002,N_7198);
nor U7962 (N_7962,N_7162,N_7166);
nand U7963 (N_7963,N_7373,N_7181);
or U7964 (N_7964,N_7485,N_7009);
nor U7965 (N_7965,N_7300,N_7298);
and U7966 (N_7966,N_7164,N_7322);
nand U7967 (N_7967,N_7059,N_7241);
nand U7968 (N_7968,N_7491,N_7466);
nand U7969 (N_7969,N_7087,N_7160);
nor U7970 (N_7970,N_7054,N_7140);
nor U7971 (N_7971,N_7012,N_7332);
or U7972 (N_7972,N_7090,N_7371);
nor U7973 (N_7973,N_7372,N_7007);
and U7974 (N_7974,N_7302,N_7186);
nor U7975 (N_7975,N_7357,N_7370);
or U7976 (N_7976,N_7201,N_7448);
xnor U7977 (N_7977,N_7208,N_7450);
and U7978 (N_7978,N_7084,N_7013);
or U7979 (N_7979,N_7425,N_7302);
nor U7980 (N_7980,N_7376,N_7021);
and U7981 (N_7981,N_7130,N_7188);
xnor U7982 (N_7982,N_7063,N_7296);
xor U7983 (N_7983,N_7038,N_7235);
or U7984 (N_7984,N_7451,N_7234);
or U7985 (N_7985,N_7024,N_7147);
nand U7986 (N_7986,N_7388,N_7030);
nor U7987 (N_7987,N_7237,N_7317);
nand U7988 (N_7988,N_7099,N_7353);
or U7989 (N_7989,N_7100,N_7031);
xnor U7990 (N_7990,N_7307,N_7488);
nand U7991 (N_7991,N_7077,N_7084);
or U7992 (N_7992,N_7190,N_7003);
nor U7993 (N_7993,N_7340,N_7036);
nand U7994 (N_7994,N_7463,N_7346);
xnor U7995 (N_7995,N_7208,N_7077);
xnor U7996 (N_7996,N_7494,N_7326);
or U7997 (N_7997,N_7088,N_7184);
or U7998 (N_7998,N_7028,N_7371);
or U7999 (N_7999,N_7092,N_7311);
xor U8000 (N_8000,N_7834,N_7694);
or U8001 (N_8001,N_7727,N_7805);
nor U8002 (N_8002,N_7663,N_7649);
nand U8003 (N_8003,N_7511,N_7713);
nor U8004 (N_8004,N_7949,N_7558);
nor U8005 (N_8005,N_7809,N_7635);
or U8006 (N_8006,N_7785,N_7504);
nor U8007 (N_8007,N_7609,N_7795);
nor U8008 (N_8008,N_7913,N_7567);
nor U8009 (N_8009,N_7863,N_7573);
xor U8010 (N_8010,N_7963,N_7822);
and U8011 (N_8011,N_7682,N_7933);
xnor U8012 (N_8012,N_7641,N_7856);
or U8013 (N_8013,N_7736,N_7545);
and U8014 (N_8014,N_7651,N_7818);
and U8015 (N_8015,N_7642,N_7509);
nand U8016 (N_8016,N_7540,N_7537);
nand U8017 (N_8017,N_7574,N_7941);
xnor U8018 (N_8018,N_7895,N_7675);
and U8019 (N_8019,N_7897,N_7580);
and U8020 (N_8020,N_7684,N_7799);
and U8021 (N_8021,N_7846,N_7971);
and U8022 (N_8022,N_7615,N_7997);
xor U8023 (N_8023,N_7904,N_7938);
and U8024 (N_8024,N_7914,N_7668);
nor U8025 (N_8025,N_7690,N_7854);
nand U8026 (N_8026,N_7848,N_7508);
or U8027 (N_8027,N_7890,N_7951);
nand U8028 (N_8028,N_7581,N_7556);
nand U8029 (N_8029,N_7729,N_7894);
nor U8030 (N_8030,N_7717,N_7550);
xor U8031 (N_8031,N_7901,N_7975);
nand U8032 (N_8032,N_7525,N_7816);
xnor U8033 (N_8033,N_7853,N_7985);
xor U8034 (N_8034,N_7523,N_7746);
xor U8035 (N_8035,N_7942,N_7732);
nor U8036 (N_8036,N_7870,N_7921);
nor U8037 (N_8037,N_7990,N_7513);
and U8038 (N_8038,N_7843,N_7518);
and U8039 (N_8039,N_7903,N_7601);
nor U8040 (N_8040,N_7698,N_7801);
and U8041 (N_8041,N_7700,N_7959);
nor U8042 (N_8042,N_7950,N_7693);
or U8043 (N_8043,N_7503,N_7761);
xnor U8044 (N_8044,N_7733,N_7521);
or U8045 (N_8045,N_7589,N_7923);
or U8046 (N_8046,N_7578,N_7543);
xor U8047 (N_8047,N_7766,N_7747);
nor U8048 (N_8048,N_7630,N_7781);
nor U8049 (N_8049,N_7506,N_7881);
and U8050 (N_8050,N_7510,N_7815);
or U8051 (N_8051,N_7932,N_7899);
xor U8052 (N_8052,N_7887,N_7835);
xor U8053 (N_8053,N_7796,N_7632);
nand U8054 (N_8054,N_7687,N_7786);
and U8055 (N_8055,N_7628,N_7750);
nor U8056 (N_8056,N_7570,N_7878);
nor U8057 (N_8057,N_7844,N_7936);
or U8058 (N_8058,N_7531,N_7958);
or U8059 (N_8059,N_7869,N_7838);
nor U8060 (N_8060,N_7592,N_7871);
or U8061 (N_8061,N_7734,N_7626);
nor U8062 (N_8062,N_7885,N_7608);
or U8063 (N_8063,N_7538,N_7735);
and U8064 (N_8064,N_7535,N_7988);
and U8065 (N_8065,N_7876,N_7542);
nand U8066 (N_8066,N_7625,N_7820);
xor U8067 (N_8067,N_7745,N_7665);
or U8068 (N_8068,N_7962,N_7532);
nand U8069 (N_8069,N_7935,N_7814);
xor U8070 (N_8070,N_7644,N_7937);
xnor U8071 (N_8071,N_7502,N_7983);
or U8072 (N_8072,N_7945,N_7794);
and U8073 (N_8073,N_7652,N_7900);
and U8074 (N_8074,N_7517,N_7593);
and U8075 (N_8075,N_7884,N_7967);
nor U8076 (N_8076,N_7622,N_7998);
nor U8077 (N_8077,N_7519,N_7591);
or U8078 (N_8078,N_7619,N_7798);
xor U8079 (N_8079,N_7824,N_7823);
and U8080 (N_8080,N_7858,N_7765);
or U8081 (N_8081,N_7787,N_7563);
xnor U8082 (N_8082,N_7802,N_7947);
or U8083 (N_8083,N_7791,N_7516);
or U8084 (N_8084,N_7701,N_7992);
and U8085 (N_8085,N_7920,N_7548);
nor U8086 (N_8086,N_7623,N_7841);
nor U8087 (N_8087,N_7738,N_7520);
xnor U8088 (N_8088,N_7980,N_7554);
nor U8089 (N_8089,N_7678,N_7658);
nand U8090 (N_8090,N_7917,N_7655);
or U8091 (N_8091,N_7810,N_7769);
xnor U8092 (N_8092,N_7770,N_7891);
or U8093 (N_8093,N_7706,N_7879);
nor U8094 (N_8094,N_7851,N_7643);
xor U8095 (N_8095,N_7596,N_7926);
nor U8096 (N_8096,N_7565,N_7757);
xor U8097 (N_8097,N_7779,N_7832);
nor U8098 (N_8098,N_7780,N_7934);
and U8099 (N_8099,N_7603,N_7728);
xnor U8100 (N_8100,N_7893,N_7752);
nand U8101 (N_8101,N_7939,N_7915);
and U8102 (N_8102,N_7768,N_7753);
or U8103 (N_8103,N_7830,N_7528);
and U8104 (N_8104,N_7924,N_7569);
or U8105 (N_8105,N_7653,N_7677);
nor U8106 (N_8106,N_7696,N_7751);
or U8107 (N_8107,N_7555,N_7566);
and U8108 (N_8108,N_7892,N_7514);
and U8109 (N_8109,N_7600,N_7597);
and U8110 (N_8110,N_7737,N_7852);
xor U8111 (N_8111,N_7640,N_7562);
nand U8112 (N_8112,N_7703,N_7512);
nor U8113 (N_8113,N_7759,N_7704);
and U8114 (N_8114,N_7928,N_7999);
nand U8115 (N_8115,N_7866,N_7721);
nand U8116 (N_8116,N_7702,N_7788);
nand U8117 (N_8117,N_7515,N_7807);
xor U8118 (N_8118,N_7907,N_7961);
or U8119 (N_8119,N_7857,N_7719);
nand U8120 (N_8120,N_7862,N_7952);
nor U8121 (N_8121,N_7529,N_7575);
and U8122 (N_8122,N_7559,N_7875);
or U8123 (N_8123,N_7624,N_7716);
or U8124 (N_8124,N_7974,N_7964);
xor U8125 (N_8125,N_7782,N_7598);
and U8126 (N_8126,N_7731,N_7691);
xnor U8127 (N_8127,N_7507,N_7657);
nand U8128 (N_8128,N_7605,N_7916);
or U8129 (N_8129,N_7724,N_7647);
and U8130 (N_8130,N_7813,N_7965);
nor U8131 (N_8131,N_7636,N_7546);
xnor U8132 (N_8132,N_7621,N_7778);
or U8133 (N_8133,N_7760,N_7847);
or U8134 (N_8134,N_7861,N_7896);
or U8135 (N_8135,N_7995,N_7756);
or U8136 (N_8136,N_7976,N_7905);
xor U8137 (N_8137,N_7588,N_7888);
or U8138 (N_8138,N_7889,N_7973);
nor U8139 (N_8139,N_7966,N_7637);
nor U8140 (N_8140,N_7590,N_7908);
xor U8141 (N_8141,N_7882,N_7825);
or U8142 (N_8142,N_7708,N_7549);
nor U8143 (N_8143,N_7775,N_7730);
nand U8144 (N_8144,N_7577,N_7944);
or U8145 (N_8145,N_7720,N_7683);
nor U8146 (N_8146,N_7594,N_7648);
xnor U8147 (N_8147,N_7723,N_7929);
nand U8148 (N_8148,N_7533,N_7819);
xnor U8149 (N_8149,N_7855,N_7579);
nor U8150 (N_8150,N_7968,N_7777);
nand U8151 (N_8151,N_7912,N_7541);
or U8152 (N_8152,N_7804,N_7826);
xnor U8153 (N_8153,N_7501,N_7978);
nand U8154 (N_8154,N_7972,N_7634);
and U8155 (N_8155,N_7979,N_7910);
nand U8156 (N_8156,N_7865,N_7534);
xnor U8157 (N_8157,N_7638,N_7956);
nor U8158 (N_8158,N_7837,N_7650);
and U8159 (N_8159,N_7771,N_7874);
or U8160 (N_8160,N_7695,N_7705);
nand U8161 (N_8161,N_7919,N_7792);
nor U8162 (N_8162,N_7585,N_7612);
and U8163 (N_8163,N_7664,N_7987);
or U8164 (N_8164,N_7883,N_7880);
nand U8165 (N_8165,N_7860,N_7740);
or U8166 (N_8166,N_7551,N_7821);
nor U8167 (N_8167,N_7676,N_7829);
xor U8168 (N_8168,N_7714,N_7718);
nand U8169 (N_8169,N_7940,N_7654);
and U8170 (N_8170,N_7685,N_7722);
or U8171 (N_8171,N_7544,N_7697);
and U8172 (N_8172,N_7877,N_7681);
xor U8173 (N_8173,N_7726,N_7955);
xnor U8174 (N_8174,N_7828,N_7827);
nor U8175 (N_8175,N_7604,N_7868);
nor U8176 (N_8176,N_7500,N_7773);
nand U8177 (N_8177,N_7616,N_7833);
or U8178 (N_8178,N_7618,N_7557);
nor U8179 (N_8179,N_7789,N_7991);
and U8180 (N_8180,N_7595,N_7686);
nand U8181 (N_8181,N_7839,N_7748);
nand U8182 (N_8182,N_7560,N_7667);
xnor U8183 (N_8183,N_7661,N_7505);
or U8184 (N_8184,N_7969,N_7898);
xor U8185 (N_8185,N_7688,N_7536);
and U8186 (N_8186,N_7539,N_7553);
and U8187 (N_8187,N_7522,N_7859);
nor U8188 (N_8188,N_7599,N_7864);
nand U8189 (N_8189,N_7666,N_7960);
and U8190 (N_8190,N_7806,N_7755);
nand U8191 (N_8191,N_7849,N_7996);
xor U8192 (N_8192,N_7671,N_7783);
nand U8193 (N_8193,N_7572,N_7679);
and U8194 (N_8194,N_7840,N_7584);
nor U8195 (N_8195,N_7925,N_7922);
nand U8196 (N_8196,N_7711,N_7656);
xor U8197 (N_8197,N_7709,N_7743);
xnor U8198 (N_8198,N_7568,N_7571);
xnor U8199 (N_8199,N_7981,N_7930);
or U8200 (N_8200,N_7842,N_7631);
or U8201 (N_8201,N_7762,N_7524);
or U8202 (N_8202,N_7911,N_7530);
or U8203 (N_8203,N_7943,N_7547);
or U8204 (N_8204,N_7606,N_7772);
xnor U8205 (N_8205,N_7629,N_7872);
or U8206 (N_8206,N_7527,N_7715);
and U8207 (N_8207,N_7946,N_7583);
nor U8208 (N_8208,N_7909,N_7673);
nand U8209 (N_8209,N_7927,N_7957);
nand U8210 (N_8210,N_7776,N_7607);
and U8211 (N_8211,N_7582,N_7587);
or U8212 (N_8212,N_7873,N_7984);
or U8213 (N_8213,N_7639,N_7808);
or U8214 (N_8214,N_7948,N_7906);
and U8215 (N_8215,N_7749,N_7797);
xor U8216 (N_8216,N_7767,N_7672);
nor U8217 (N_8217,N_7977,N_7758);
or U8218 (N_8218,N_7602,N_7774);
nor U8219 (N_8219,N_7812,N_7803);
nor U8220 (N_8220,N_7744,N_7660);
nor U8221 (N_8221,N_7831,N_7561);
nand U8222 (N_8222,N_7611,N_7725);
nand U8223 (N_8223,N_7886,N_7627);
nor U8224 (N_8224,N_7564,N_7764);
nor U8225 (N_8225,N_7669,N_7982);
or U8226 (N_8226,N_7994,N_7953);
xnor U8227 (N_8227,N_7646,N_7845);
xor U8228 (N_8228,N_7680,N_7954);
or U8229 (N_8229,N_7692,N_7784);
nor U8230 (N_8230,N_7754,N_7902);
or U8231 (N_8231,N_7633,N_7970);
xor U8232 (N_8232,N_7850,N_7699);
and U8233 (N_8233,N_7836,N_7986);
and U8234 (N_8234,N_7526,N_7931);
xnor U8235 (N_8235,N_7793,N_7645);
and U8236 (N_8236,N_7993,N_7670);
and U8237 (N_8237,N_7739,N_7741);
or U8238 (N_8238,N_7614,N_7707);
nor U8239 (N_8239,N_7867,N_7817);
and U8240 (N_8240,N_7674,N_7576);
nand U8241 (N_8241,N_7763,N_7662);
or U8242 (N_8242,N_7613,N_7800);
nor U8243 (N_8243,N_7610,N_7617);
or U8244 (N_8244,N_7710,N_7989);
nor U8245 (N_8245,N_7689,N_7620);
or U8246 (N_8246,N_7659,N_7586);
nor U8247 (N_8247,N_7811,N_7712);
nor U8248 (N_8248,N_7790,N_7552);
or U8249 (N_8249,N_7742,N_7918);
nand U8250 (N_8250,N_7678,N_7686);
nor U8251 (N_8251,N_7881,N_7814);
xnor U8252 (N_8252,N_7724,N_7625);
nand U8253 (N_8253,N_7834,N_7505);
or U8254 (N_8254,N_7944,N_7593);
xor U8255 (N_8255,N_7735,N_7983);
xnor U8256 (N_8256,N_7507,N_7540);
and U8257 (N_8257,N_7969,N_7900);
xor U8258 (N_8258,N_7728,N_7752);
nand U8259 (N_8259,N_7564,N_7690);
or U8260 (N_8260,N_7761,N_7867);
nor U8261 (N_8261,N_7852,N_7670);
nor U8262 (N_8262,N_7996,N_7917);
xnor U8263 (N_8263,N_7623,N_7508);
or U8264 (N_8264,N_7623,N_7541);
nor U8265 (N_8265,N_7940,N_7934);
nand U8266 (N_8266,N_7631,N_7883);
xnor U8267 (N_8267,N_7555,N_7536);
or U8268 (N_8268,N_7924,N_7883);
nand U8269 (N_8269,N_7553,N_7547);
xor U8270 (N_8270,N_7632,N_7943);
and U8271 (N_8271,N_7503,N_7536);
xnor U8272 (N_8272,N_7998,N_7541);
and U8273 (N_8273,N_7954,N_7959);
or U8274 (N_8274,N_7679,N_7557);
nor U8275 (N_8275,N_7835,N_7779);
nand U8276 (N_8276,N_7534,N_7548);
nor U8277 (N_8277,N_7648,N_7723);
nor U8278 (N_8278,N_7643,N_7926);
and U8279 (N_8279,N_7856,N_7626);
nor U8280 (N_8280,N_7952,N_7797);
nor U8281 (N_8281,N_7614,N_7701);
or U8282 (N_8282,N_7636,N_7911);
nand U8283 (N_8283,N_7949,N_7528);
xnor U8284 (N_8284,N_7868,N_7690);
or U8285 (N_8285,N_7749,N_7983);
or U8286 (N_8286,N_7923,N_7831);
and U8287 (N_8287,N_7533,N_7692);
nor U8288 (N_8288,N_7825,N_7885);
nand U8289 (N_8289,N_7575,N_7739);
or U8290 (N_8290,N_7557,N_7563);
and U8291 (N_8291,N_7885,N_7679);
and U8292 (N_8292,N_7971,N_7570);
and U8293 (N_8293,N_7736,N_7768);
nand U8294 (N_8294,N_7664,N_7921);
and U8295 (N_8295,N_7607,N_7613);
or U8296 (N_8296,N_7555,N_7552);
nand U8297 (N_8297,N_7712,N_7841);
nand U8298 (N_8298,N_7951,N_7554);
nand U8299 (N_8299,N_7578,N_7557);
xnor U8300 (N_8300,N_7802,N_7890);
nand U8301 (N_8301,N_7847,N_7730);
xnor U8302 (N_8302,N_7689,N_7650);
xor U8303 (N_8303,N_7701,N_7656);
nand U8304 (N_8304,N_7645,N_7964);
xor U8305 (N_8305,N_7752,N_7855);
or U8306 (N_8306,N_7995,N_7968);
nor U8307 (N_8307,N_7585,N_7759);
nand U8308 (N_8308,N_7847,N_7861);
xor U8309 (N_8309,N_7904,N_7844);
and U8310 (N_8310,N_7983,N_7806);
nand U8311 (N_8311,N_7611,N_7855);
nand U8312 (N_8312,N_7732,N_7585);
nor U8313 (N_8313,N_7676,N_7762);
nor U8314 (N_8314,N_7784,N_7605);
xor U8315 (N_8315,N_7870,N_7695);
nor U8316 (N_8316,N_7551,N_7847);
xor U8317 (N_8317,N_7540,N_7744);
or U8318 (N_8318,N_7885,N_7769);
or U8319 (N_8319,N_7753,N_7795);
nand U8320 (N_8320,N_7737,N_7800);
nand U8321 (N_8321,N_7654,N_7556);
xor U8322 (N_8322,N_7679,N_7960);
and U8323 (N_8323,N_7650,N_7872);
nor U8324 (N_8324,N_7695,N_7630);
or U8325 (N_8325,N_7767,N_7884);
or U8326 (N_8326,N_7743,N_7796);
and U8327 (N_8327,N_7520,N_7787);
or U8328 (N_8328,N_7787,N_7544);
nor U8329 (N_8329,N_7741,N_7944);
xor U8330 (N_8330,N_7509,N_7501);
and U8331 (N_8331,N_7721,N_7737);
or U8332 (N_8332,N_7812,N_7763);
nor U8333 (N_8333,N_7542,N_7533);
nor U8334 (N_8334,N_7741,N_7710);
or U8335 (N_8335,N_7875,N_7753);
nor U8336 (N_8336,N_7599,N_7533);
nor U8337 (N_8337,N_7717,N_7618);
and U8338 (N_8338,N_7855,N_7517);
or U8339 (N_8339,N_7555,N_7514);
nand U8340 (N_8340,N_7924,N_7816);
nand U8341 (N_8341,N_7790,N_7721);
xor U8342 (N_8342,N_7581,N_7997);
nand U8343 (N_8343,N_7997,N_7870);
nand U8344 (N_8344,N_7780,N_7924);
nand U8345 (N_8345,N_7771,N_7595);
nand U8346 (N_8346,N_7628,N_7626);
nand U8347 (N_8347,N_7624,N_7776);
nor U8348 (N_8348,N_7700,N_7547);
nand U8349 (N_8349,N_7735,N_7819);
xnor U8350 (N_8350,N_7969,N_7858);
nor U8351 (N_8351,N_7671,N_7631);
and U8352 (N_8352,N_7807,N_7831);
nand U8353 (N_8353,N_7654,N_7984);
nor U8354 (N_8354,N_7926,N_7955);
and U8355 (N_8355,N_7745,N_7617);
xor U8356 (N_8356,N_7929,N_7830);
xor U8357 (N_8357,N_7703,N_7843);
and U8358 (N_8358,N_7713,N_7855);
nand U8359 (N_8359,N_7857,N_7508);
nand U8360 (N_8360,N_7976,N_7667);
xnor U8361 (N_8361,N_7593,N_7553);
and U8362 (N_8362,N_7894,N_7994);
or U8363 (N_8363,N_7993,N_7843);
nor U8364 (N_8364,N_7529,N_7666);
and U8365 (N_8365,N_7713,N_7643);
nand U8366 (N_8366,N_7721,N_7740);
xnor U8367 (N_8367,N_7882,N_7768);
and U8368 (N_8368,N_7674,N_7706);
nand U8369 (N_8369,N_7826,N_7776);
and U8370 (N_8370,N_7546,N_7569);
or U8371 (N_8371,N_7847,N_7965);
nand U8372 (N_8372,N_7757,N_7901);
xnor U8373 (N_8373,N_7762,N_7998);
xor U8374 (N_8374,N_7515,N_7732);
and U8375 (N_8375,N_7936,N_7619);
or U8376 (N_8376,N_7761,N_7562);
nand U8377 (N_8377,N_7761,N_7624);
nor U8378 (N_8378,N_7745,N_7720);
xor U8379 (N_8379,N_7632,N_7690);
or U8380 (N_8380,N_7938,N_7673);
or U8381 (N_8381,N_7948,N_7685);
and U8382 (N_8382,N_7823,N_7975);
or U8383 (N_8383,N_7717,N_7986);
or U8384 (N_8384,N_7849,N_7718);
nand U8385 (N_8385,N_7792,N_7749);
xnor U8386 (N_8386,N_7994,N_7905);
nor U8387 (N_8387,N_7863,N_7593);
nor U8388 (N_8388,N_7782,N_7587);
nand U8389 (N_8389,N_7509,N_7776);
and U8390 (N_8390,N_7875,N_7589);
or U8391 (N_8391,N_7629,N_7656);
xnor U8392 (N_8392,N_7702,N_7982);
and U8393 (N_8393,N_7542,N_7874);
xnor U8394 (N_8394,N_7743,N_7636);
nor U8395 (N_8395,N_7914,N_7853);
and U8396 (N_8396,N_7634,N_7655);
or U8397 (N_8397,N_7713,N_7895);
xnor U8398 (N_8398,N_7711,N_7789);
and U8399 (N_8399,N_7641,N_7886);
nor U8400 (N_8400,N_7970,N_7921);
and U8401 (N_8401,N_7684,N_7869);
nand U8402 (N_8402,N_7929,N_7961);
xnor U8403 (N_8403,N_7550,N_7729);
nor U8404 (N_8404,N_7583,N_7926);
or U8405 (N_8405,N_7996,N_7625);
nand U8406 (N_8406,N_7698,N_7791);
nor U8407 (N_8407,N_7573,N_7978);
and U8408 (N_8408,N_7602,N_7904);
nor U8409 (N_8409,N_7987,N_7611);
nand U8410 (N_8410,N_7801,N_7560);
nor U8411 (N_8411,N_7828,N_7873);
or U8412 (N_8412,N_7635,N_7798);
nand U8413 (N_8413,N_7876,N_7509);
xnor U8414 (N_8414,N_7778,N_7630);
nor U8415 (N_8415,N_7721,N_7524);
nand U8416 (N_8416,N_7868,N_7541);
and U8417 (N_8417,N_7567,N_7854);
xor U8418 (N_8418,N_7968,N_7563);
and U8419 (N_8419,N_7893,N_7787);
nor U8420 (N_8420,N_7866,N_7675);
nand U8421 (N_8421,N_7567,N_7595);
nor U8422 (N_8422,N_7516,N_7762);
xnor U8423 (N_8423,N_7700,N_7898);
nand U8424 (N_8424,N_7989,N_7871);
nand U8425 (N_8425,N_7951,N_7641);
nor U8426 (N_8426,N_7958,N_7761);
nor U8427 (N_8427,N_7673,N_7951);
xor U8428 (N_8428,N_7840,N_7796);
nor U8429 (N_8429,N_7579,N_7767);
nand U8430 (N_8430,N_7941,N_7640);
and U8431 (N_8431,N_7830,N_7527);
xor U8432 (N_8432,N_7782,N_7621);
or U8433 (N_8433,N_7722,N_7838);
xor U8434 (N_8434,N_7650,N_7767);
nand U8435 (N_8435,N_7911,N_7569);
nand U8436 (N_8436,N_7770,N_7791);
nor U8437 (N_8437,N_7759,N_7763);
and U8438 (N_8438,N_7899,N_7939);
or U8439 (N_8439,N_7912,N_7887);
or U8440 (N_8440,N_7884,N_7601);
xnor U8441 (N_8441,N_7860,N_7824);
xnor U8442 (N_8442,N_7668,N_7906);
nand U8443 (N_8443,N_7574,N_7673);
and U8444 (N_8444,N_7601,N_7667);
nor U8445 (N_8445,N_7769,N_7648);
nand U8446 (N_8446,N_7989,N_7720);
and U8447 (N_8447,N_7709,N_7990);
xor U8448 (N_8448,N_7569,N_7835);
and U8449 (N_8449,N_7543,N_7762);
or U8450 (N_8450,N_7993,N_7826);
xor U8451 (N_8451,N_7867,N_7509);
nand U8452 (N_8452,N_7794,N_7863);
xnor U8453 (N_8453,N_7648,N_7898);
xnor U8454 (N_8454,N_7575,N_7994);
and U8455 (N_8455,N_7908,N_7825);
nor U8456 (N_8456,N_7790,N_7837);
and U8457 (N_8457,N_7763,N_7786);
xor U8458 (N_8458,N_7550,N_7514);
nand U8459 (N_8459,N_7662,N_7605);
nand U8460 (N_8460,N_7781,N_7704);
and U8461 (N_8461,N_7781,N_7984);
nor U8462 (N_8462,N_7893,N_7958);
nand U8463 (N_8463,N_7657,N_7861);
nand U8464 (N_8464,N_7596,N_7632);
nand U8465 (N_8465,N_7749,N_7659);
or U8466 (N_8466,N_7848,N_7910);
or U8467 (N_8467,N_7774,N_7976);
nor U8468 (N_8468,N_7719,N_7978);
nor U8469 (N_8469,N_7642,N_7582);
or U8470 (N_8470,N_7795,N_7925);
xnor U8471 (N_8471,N_7796,N_7801);
xor U8472 (N_8472,N_7541,N_7567);
nor U8473 (N_8473,N_7706,N_7802);
and U8474 (N_8474,N_7819,N_7747);
xnor U8475 (N_8475,N_7510,N_7958);
or U8476 (N_8476,N_7548,N_7721);
xor U8477 (N_8477,N_7588,N_7610);
nand U8478 (N_8478,N_7791,N_7610);
and U8479 (N_8479,N_7825,N_7844);
nand U8480 (N_8480,N_7645,N_7557);
and U8481 (N_8481,N_7744,N_7560);
nand U8482 (N_8482,N_7527,N_7779);
or U8483 (N_8483,N_7778,N_7783);
or U8484 (N_8484,N_7613,N_7586);
or U8485 (N_8485,N_7601,N_7761);
nor U8486 (N_8486,N_7987,N_7706);
nor U8487 (N_8487,N_7757,N_7744);
xor U8488 (N_8488,N_7963,N_7570);
and U8489 (N_8489,N_7648,N_7764);
nor U8490 (N_8490,N_7833,N_7821);
nor U8491 (N_8491,N_7849,N_7514);
nor U8492 (N_8492,N_7509,N_7683);
nor U8493 (N_8493,N_7571,N_7911);
and U8494 (N_8494,N_7664,N_7949);
and U8495 (N_8495,N_7914,N_7595);
xnor U8496 (N_8496,N_7837,N_7900);
nand U8497 (N_8497,N_7850,N_7678);
or U8498 (N_8498,N_7551,N_7716);
nand U8499 (N_8499,N_7655,N_7961);
or U8500 (N_8500,N_8010,N_8441);
xor U8501 (N_8501,N_8257,N_8423);
nor U8502 (N_8502,N_8342,N_8496);
and U8503 (N_8503,N_8198,N_8160);
and U8504 (N_8504,N_8260,N_8458);
nand U8505 (N_8505,N_8226,N_8143);
xnor U8506 (N_8506,N_8339,N_8209);
or U8507 (N_8507,N_8492,N_8351);
nor U8508 (N_8508,N_8246,N_8466);
or U8509 (N_8509,N_8336,N_8296);
nor U8510 (N_8510,N_8448,N_8074);
nand U8511 (N_8511,N_8473,N_8359);
xnor U8512 (N_8512,N_8446,N_8028);
nor U8513 (N_8513,N_8371,N_8080);
or U8514 (N_8514,N_8460,N_8439);
nor U8515 (N_8515,N_8174,N_8271);
nor U8516 (N_8516,N_8258,N_8373);
nand U8517 (N_8517,N_8369,N_8155);
and U8518 (N_8518,N_8129,N_8150);
or U8519 (N_8519,N_8366,N_8071);
nor U8520 (N_8520,N_8130,N_8285);
or U8521 (N_8521,N_8135,N_8265);
or U8522 (N_8522,N_8292,N_8056);
nand U8523 (N_8523,N_8016,N_8240);
xor U8524 (N_8524,N_8133,N_8268);
and U8525 (N_8525,N_8344,N_8361);
xnor U8526 (N_8526,N_8352,N_8353);
and U8527 (N_8527,N_8485,N_8327);
and U8528 (N_8528,N_8462,N_8443);
nor U8529 (N_8529,N_8193,N_8430);
nand U8530 (N_8530,N_8020,N_8375);
nand U8531 (N_8531,N_8186,N_8166);
nand U8532 (N_8532,N_8293,N_8456);
xnor U8533 (N_8533,N_8329,N_8230);
and U8534 (N_8534,N_8228,N_8108);
nor U8535 (N_8535,N_8477,N_8343);
or U8536 (N_8536,N_8459,N_8383);
nor U8537 (N_8537,N_8414,N_8066);
xnor U8538 (N_8538,N_8461,N_8131);
and U8539 (N_8539,N_8086,N_8192);
and U8540 (N_8540,N_8031,N_8061);
nor U8541 (N_8541,N_8291,N_8057);
xnor U8542 (N_8542,N_8030,N_8280);
nand U8543 (N_8543,N_8404,N_8217);
nand U8544 (N_8544,N_8011,N_8349);
xnor U8545 (N_8545,N_8424,N_8249);
xor U8546 (N_8546,N_8043,N_8138);
or U8547 (N_8547,N_8019,N_8085);
and U8548 (N_8548,N_8163,N_8103);
or U8549 (N_8549,N_8137,N_8488);
nor U8550 (N_8550,N_8175,N_8451);
xnor U8551 (N_8551,N_8207,N_8070);
nor U8552 (N_8552,N_8204,N_8114);
nand U8553 (N_8553,N_8410,N_8440);
nand U8554 (N_8554,N_8241,N_8478);
nor U8555 (N_8555,N_8282,N_8310);
xor U8556 (N_8556,N_8153,N_8438);
xor U8557 (N_8557,N_8202,N_8255);
xor U8558 (N_8558,N_8127,N_8323);
xor U8559 (N_8559,N_8363,N_8376);
or U8560 (N_8560,N_8245,N_8356);
nor U8561 (N_8561,N_8382,N_8469);
nand U8562 (N_8562,N_8315,N_8001);
or U8563 (N_8563,N_8360,N_8279);
nand U8564 (N_8564,N_8232,N_8378);
xor U8565 (N_8565,N_8231,N_8038);
or U8566 (N_8566,N_8262,N_8183);
nand U8567 (N_8567,N_8158,N_8264);
xnor U8568 (N_8568,N_8152,N_8309);
xor U8569 (N_8569,N_8429,N_8453);
nor U8570 (N_8570,N_8128,N_8101);
or U8571 (N_8571,N_8076,N_8178);
and U8572 (N_8572,N_8023,N_8015);
or U8573 (N_8573,N_8092,N_8465);
nand U8574 (N_8574,N_8234,N_8391);
nand U8575 (N_8575,N_8390,N_8139);
nand U8576 (N_8576,N_8332,N_8165);
nor U8577 (N_8577,N_8215,N_8495);
nor U8578 (N_8578,N_8005,N_8433);
xnor U8579 (N_8579,N_8412,N_8384);
nand U8580 (N_8580,N_8381,N_8046);
and U8581 (N_8581,N_8110,N_8377);
and U8582 (N_8582,N_8340,N_8445);
nor U8583 (N_8583,N_8312,N_8027);
nand U8584 (N_8584,N_8077,N_8358);
and U8585 (N_8585,N_8078,N_8491);
nor U8586 (N_8586,N_8346,N_8029);
nor U8587 (N_8587,N_8051,N_8203);
nor U8588 (N_8588,N_8252,N_8059);
nor U8589 (N_8589,N_8302,N_8156);
xnor U8590 (N_8590,N_8251,N_8301);
or U8591 (N_8591,N_8179,N_8437);
nor U8592 (N_8592,N_8096,N_8483);
and U8593 (N_8593,N_8284,N_8069);
and U8594 (N_8594,N_8288,N_8393);
nor U8595 (N_8595,N_8317,N_8134);
nand U8596 (N_8596,N_8450,N_8106);
xor U8597 (N_8597,N_8300,N_8374);
or U8598 (N_8598,N_8159,N_8338);
or U8599 (N_8599,N_8233,N_8024);
nor U8600 (N_8600,N_8169,N_8331);
or U8601 (N_8601,N_8003,N_8012);
xnor U8602 (N_8602,N_8314,N_8164);
and U8603 (N_8603,N_8000,N_8102);
nand U8604 (N_8604,N_8125,N_8357);
nand U8605 (N_8605,N_8499,N_8425);
or U8606 (N_8606,N_8111,N_8455);
and U8607 (N_8607,N_8033,N_8224);
nand U8608 (N_8608,N_8487,N_8263);
nand U8609 (N_8609,N_8189,N_8321);
and U8610 (N_8610,N_8308,N_8354);
nand U8611 (N_8611,N_8136,N_8417);
or U8612 (N_8612,N_8259,N_8145);
nor U8613 (N_8613,N_8188,N_8047);
xnor U8614 (N_8614,N_8415,N_8093);
nand U8615 (N_8615,N_8398,N_8287);
and U8616 (N_8616,N_8432,N_8457);
and U8617 (N_8617,N_8431,N_8472);
nand U8618 (N_8618,N_8149,N_8079);
xnor U8619 (N_8619,N_8107,N_8118);
or U8620 (N_8620,N_8082,N_8148);
xor U8621 (N_8621,N_8008,N_8109);
nand U8622 (N_8622,N_8094,N_8442);
xor U8623 (N_8623,N_8223,N_8479);
nor U8624 (N_8624,N_8413,N_8176);
xnor U8625 (N_8625,N_8054,N_8277);
nor U8626 (N_8626,N_8269,N_8238);
and U8627 (N_8627,N_8042,N_8434);
or U8628 (N_8628,N_8062,N_8484);
and U8629 (N_8629,N_8403,N_8229);
xnor U8630 (N_8630,N_8050,N_8385);
xor U8631 (N_8631,N_8064,N_8147);
and U8632 (N_8632,N_8362,N_8196);
nor U8633 (N_8633,N_8368,N_8256);
nor U8634 (N_8634,N_8075,N_8225);
nand U8635 (N_8635,N_8348,N_8201);
or U8636 (N_8636,N_8489,N_8113);
xor U8637 (N_8637,N_8286,N_8290);
nand U8638 (N_8638,N_8182,N_8270);
nand U8639 (N_8639,N_8411,N_8266);
nand U8640 (N_8640,N_8401,N_8330);
nor U8641 (N_8641,N_8191,N_8272);
nand U8642 (N_8642,N_8387,N_8400);
xnor U8643 (N_8643,N_8180,N_8497);
nor U8644 (N_8644,N_8392,N_8243);
and U8645 (N_8645,N_8123,N_8091);
nor U8646 (N_8646,N_8289,N_8370);
or U8647 (N_8647,N_8476,N_8018);
or U8648 (N_8648,N_8017,N_8205);
or U8649 (N_8649,N_8173,N_8333);
and U8650 (N_8650,N_8426,N_8200);
or U8651 (N_8651,N_8090,N_8474);
and U8652 (N_8652,N_8299,N_8171);
xor U8653 (N_8653,N_8386,N_8151);
or U8654 (N_8654,N_8408,N_8002);
or U8655 (N_8655,N_8281,N_8420);
nor U8656 (N_8656,N_8195,N_8006);
and U8657 (N_8657,N_8480,N_8112);
and U8658 (N_8658,N_8117,N_8161);
xnor U8659 (N_8659,N_8427,N_8475);
and U8660 (N_8660,N_8222,N_8396);
xnor U8661 (N_8661,N_8388,N_8482);
and U8662 (N_8662,N_8493,N_8097);
and U8663 (N_8663,N_8212,N_8436);
or U8664 (N_8664,N_8468,N_8304);
and U8665 (N_8665,N_8157,N_8341);
xor U8666 (N_8666,N_8063,N_8334);
nand U8667 (N_8667,N_8444,N_8283);
and U8668 (N_8668,N_8126,N_8294);
nand U8669 (N_8669,N_8470,N_8072);
nand U8670 (N_8670,N_8058,N_8307);
xor U8671 (N_8671,N_8274,N_8303);
and U8672 (N_8672,N_8402,N_8247);
nor U8673 (N_8673,N_8372,N_8467);
nand U8674 (N_8674,N_8041,N_8248);
nand U8675 (N_8675,N_8380,N_8452);
and U8676 (N_8676,N_8276,N_8237);
xnor U8677 (N_8677,N_8124,N_8365);
and U8678 (N_8678,N_8236,N_8298);
nor U8679 (N_8679,N_8190,N_8405);
xnor U8680 (N_8680,N_8235,N_8407);
nand U8681 (N_8681,N_8490,N_8220);
or U8682 (N_8682,N_8034,N_8167);
and U8683 (N_8683,N_8239,N_8039);
nand U8684 (N_8684,N_8187,N_8142);
or U8685 (N_8685,N_8242,N_8214);
or U8686 (N_8686,N_8406,N_8140);
xor U8687 (N_8687,N_8267,N_8199);
xor U8688 (N_8688,N_8098,N_8449);
nand U8689 (N_8689,N_8170,N_8325);
xor U8690 (N_8690,N_8318,N_8185);
or U8691 (N_8691,N_8121,N_8087);
nor U8692 (N_8692,N_8115,N_8089);
xor U8693 (N_8693,N_8278,N_8014);
nor U8694 (N_8694,N_8211,N_8021);
nand U8695 (N_8695,N_8494,N_8146);
and U8696 (N_8696,N_8177,N_8026);
nand U8697 (N_8697,N_8421,N_8035);
nand U8698 (N_8698,N_8007,N_8168);
or U8699 (N_8699,N_8335,N_8454);
xor U8700 (N_8700,N_8037,N_8320);
and U8701 (N_8701,N_8295,N_8297);
nand U8702 (N_8702,N_8324,N_8206);
or U8703 (N_8703,N_8355,N_8254);
and U8704 (N_8704,N_8073,N_8316);
nor U8705 (N_8705,N_8227,N_8210);
and U8706 (N_8706,N_8218,N_8049);
or U8707 (N_8707,N_8221,N_8172);
or U8708 (N_8708,N_8498,N_8040);
or U8709 (N_8709,N_8162,N_8141);
nand U8710 (N_8710,N_8181,N_8144);
or U8711 (N_8711,N_8122,N_8194);
xnor U8712 (N_8712,N_8253,N_8464);
nor U8713 (N_8713,N_8032,N_8067);
nor U8714 (N_8714,N_8219,N_8463);
xor U8715 (N_8715,N_8347,N_8084);
and U8716 (N_8716,N_8306,N_8004);
nor U8717 (N_8717,N_8435,N_8013);
nand U8718 (N_8718,N_8104,N_8052);
xor U8719 (N_8719,N_8399,N_8081);
and U8720 (N_8720,N_8250,N_8313);
nor U8721 (N_8721,N_8060,N_8055);
nand U8722 (N_8722,N_8486,N_8244);
or U8723 (N_8723,N_8305,N_8044);
xnor U8724 (N_8724,N_8095,N_8120);
xnor U8725 (N_8725,N_8099,N_8481);
and U8726 (N_8726,N_8261,N_8065);
nand U8727 (N_8727,N_8022,N_8213);
or U8728 (N_8728,N_8328,N_8025);
nor U8729 (N_8729,N_8367,N_8119);
nor U8730 (N_8730,N_8273,N_8275);
and U8731 (N_8731,N_8326,N_8088);
nand U8732 (N_8732,N_8345,N_8428);
xnor U8733 (N_8733,N_8009,N_8053);
nor U8734 (N_8734,N_8395,N_8184);
xnor U8735 (N_8735,N_8389,N_8322);
xnor U8736 (N_8736,N_8036,N_8216);
nor U8737 (N_8737,N_8337,N_8154);
nand U8738 (N_8738,N_8422,N_8208);
or U8739 (N_8739,N_8364,N_8068);
nor U8740 (N_8740,N_8379,N_8100);
xor U8741 (N_8741,N_8045,N_8397);
nand U8742 (N_8742,N_8105,N_8350);
or U8743 (N_8743,N_8416,N_8197);
or U8744 (N_8744,N_8394,N_8418);
and U8745 (N_8745,N_8419,N_8319);
or U8746 (N_8746,N_8447,N_8409);
and U8747 (N_8747,N_8048,N_8132);
nor U8748 (N_8748,N_8311,N_8471);
nand U8749 (N_8749,N_8116,N_8083);
or U8750 (N_8750,N_8334,N_8335);
nand U8751 (N_8751,N_8455,N_8273);
nor U8752 (N_8752,N_8083,N_8428);
xnor U8753 (N_8753,N_8292,N_8451);
nand U8754 (N_8754,N_8134,N_8342);
or U8755 (N_8755,N_8331,N_8434);
nand U8756 (N_8756,N_8295,N_8144);
and U8757 (N_8757,N_8296,N_8395);
nand U8758 (N_8758,N_8146,N_8258);
nand U8759 (N_8759,N_8451,N_8101);
and U8760 (N_8760,N_8330,N_8296);
and U8761 (N_8761,N_8421,N_8389);
xor U8762 (N_8762,N_8236,N_8192);
xnor U8763 (N_8763,N_8197,N_8467);
and U8764 (N_8764,N_8296,N_8489);
nand U8765 (N_8765,N_8078,N_8195);
and U8766 (N_8766,N_8093,N_8382);
nand U8767 (N_8767,N_8302,N_8011);
xnor U8768 (N_8768,N_8386,N_8470);
and U8769 (N_8769,N_8462,N_8465);
xor U8770 (N_8770,N_8180,N_8231);
nor U8771 (N_8771,N_8394,N_8035);
nor U8772 (N_8772,N_8335,N_8251);
nor U8773 (N_8773,N_8495,N_8482);
or U8774 (N_8774,N_8457,N_8387);
xnor U8775 (N_8775,N_8282,N_8400);
nor U8776 (N_8776,N_8266,N_8126);
or U8777 (N_8777,N_8108,N_8457);
xnor U8778 (N_8778,N_8116,N_8260);
or U8779 (N_8779,N_8322,N_8220);
and U8780 (N_8780,N_8305,N_8473);
or U8781 (N_8781,N_8152,N_8086);
or U8782 (N_8782,N_8372,N_8336);
nand U8783 (N_8783,N_8140,N_8139);
and U8784 (N_8784,N_8150,N_8143);
xor U8785 (N_8785,N_8005,N_8103);
or U8786 (N_8786,N_8109,N_8221);
xnor U8787 (N_8787,N_8389,N_8328);
or U8788 (N_8788,N_8013,N_8231);
nand U8789 (N_8789,N_8144,N_8185);
xnor U8790 (N_8790,N_8120,N_8131);
or U8791 (N_8791,N_8488,N_8312);
nand U8792 (N_8792,N_8092,N_8143);
xor U8793 (N_8793,N_8100,N_8456);
or U8794 (N_8794,N_8415,N_8008);
or U8795 (N_8795,N_8489,N_8118);
nand U8796 (N_8796,N_8319,N_8367);
nor U8797 (N_8797,N_8162,N_8291);
nor U8798 (N_8798,N_8385,N_8012);
nor U8799 (N_8799,N_8309,N_8094);
and U8800 (N_8800,N_8486,N_8499);
xnor U8801 (N_8801,N_8409,N_8251);
or U8802 (N_8802,N_8236,N_8432);
xnor U8803 (N_8803,N_8493,N_8288);
nand U8804 (N_8804,N_8455,N_8317);
and U8805 (N_8805,N_8350,N_8496);
nor U8806 (N_8806,N_8453,N_8225);
and U8807 (N_8807,N_8188,N_8132);
and U8808 (N_8808,N_8425,N_8399);
xor U8809 (N_8809,N_8334,N_8262);
nor U8810 (N_8810,N_8224,N_8138);
xnor U8811 (N_8811,N_8210,N_8476);
or U8812 (N_8812,N_8045,N_8050);
nand U8813 (N_8813,N_8350,N_8036);
xor U8814 (N_8814,N_8433,N_8125);
or U8815 (N_8815,N_8030,N_8181);
nor U8816 (N_8816,N_8239,N_8456);
nor U8817 (N_8817,N_8425,N_8067);
nand U8818 (N_8818,N_8070,N_8375);
nand U8819 (N_8819,N_8282,N_8022);
and U8820 (N_8820,N_8225,N_8175);
nor U8821 (N_8821,N_8487,N_8309);
nand U8822 (N_8822,N_8196,N_8312);
xnor U8823 (N_8823,N_8117,N_8360);
and U8824 (N_8824,N_8179,N_8082);
and U8825 (N_8825,N_8377,N_8211);
xor U8826 (N_8826,N_8103,N_8165);
and U8827 (N_8827,N_8181,N_8241);
nand U8828 (N_8828,N_8320,N_8427);
or U8829 (N_8829,N_8400,N_8444);
nand U8830 (N_8830,N_8417,N_8076);
and U8831 (N_8831,N_8355,N_8147);
nor U8832 (N_8832,N_8165,N_8404);
or U8833 (N_8833,N_8032,N_8216);
or U8834 (N_8834,N_8061,N_8141);
xor U8835 (N_8835,N_8225,N_8150);
or U8836 (N_8836,N_8071,N_8394);
nor U8837 (N_8837,N_8321,N_8473);
or U8838 (N_8838,N_8348,N_8367);
nor U8839 (N_8839,N_8417,N_8234);
nand U8840 (N_8840,N_8269,N_8333);
and U8841 (N_8841,N_8461,N_8295);
or U8842 (N_8842,N_8341,N_8284);
xor U8843 (N_8843,N_8298,N_8353);
xnor U8844 (N_8844,N_8470,N_8466);
and U8845 (N_8845,N_8022,N_8246);
nor U8846 (N_8846,N_8289,N_8071);
or U8847 (N_8847,N_8263,N_8488);
or U8848 (N_8848,N_8106,N_8029);
nand U8849 (N_8849,N_8104,N_8352);
nor U8850 (N_8850,N_8151,N_8006);
nor U8851 (N_8851,N_8108,N_8432);
nand U8852 (N_8852,N_8190,N_8396);
or U8853 (N_8853,N_8002,N_8292);
nor U8854 (N_8854,N_8204,N_8333);
or U8855 (N_8855,N_8167,N_8124);
nand U8856 (N_8856,N_8128,N_8434);
or U8857 (N_8857,N_8243,N_8067);
nand U8858 (N_8858,N_8030,N_8229);
nor U8859 (N_8859,N_8405,N_8394);
or U8860 (N_8860,N_8224,N_8295);
nand U8861 (N_8861,N_8158,N_8276);
or U8862 (N_8862,N_8252,N_8130);
xor U8863 (N_8863,N_8396,N_8367);
or U8864 (N_8864,N_8328,N_8292);
and U8865 (N_8865,N_8052,N_8218);
or U8866 (N_8866,N_8400,N_8060);
xor U8867 (N_8867,N_8230,N_8156);
nor U8868 (N_8868,N_8195,N_8116);
and U8869 (N_8869,N_8051,N_8381);
or U8870 (N_8870,N_8106,N_8451);
xor U8871 (N_8871,N_8453,N_8043);
or U8872 (N_8872,N_8367,N_8082);
and U8873 (N_8873,N_8180,N_8388);
xor U8874 (N_8874,N_8274,N_8486);
and U8875 (N_8875,N_8353,N_8453);
xnor U8876 (N_8876,N_8235,N_8384);
xor U8877 (N_8877,N_8093,N_8322);
and U8878 (N_8878,N_8129,N_8278);
or U8879 (N_8879,N_8084,N_8213);
nand U8880 (N_8880,N_8323,N_8237);
nand U8881 (N_8881,N_8302,N_8052);
nand U8882 (N_8882,N_8229,N_8306);
nor U8883 (N_8883,N_8136,N_8039);
nand U8884 (N_8884,N_8010,N_8239);
nand U8885 (N_8885,N_8009,N_8016);
xor U8886 (N_8886,N_8255,N_8034);
or U8887 (N_8887,N_8330,N_8170);
nor U8888 (N_8888,N_8053,N_8375);
nor U8889 (N_8889,N_8175,N_8266);
nor U8890 (N_8890,N_8095,N_8068);
xnor U8891 (N_8891,N_8231,N_8448);
nor U8892 (N_8892,N_8173,N_8298);
or U8893 (N_8893,N_8462,N_8014);
nor U8894 (N_8894,N_8433,N_8070);
xnor U8895 (N_8895,N_8383,N_8472);
or U8896 (N_8896,N_8041,N_8028);
nor U8897 (N_8897,N_8139,N_8104);
xnor U8898 (N_8898,N_8404,N_8220);
nand U8899 (N_8899,N_8231,N_8238);
xnor U8900 (N_8900,N_8209,N_8206);
nor U8901 (N_8901,N_8083,N_8019);
xnor U8902 (N_8902,N_8000,N_8097);
or U8903 (N_8903,N_8388,N_8311);
xnor U8904 (N_8904,N_8174,N_8260);
or U8905 (N_8905,N_8091,N_8381);
and U8906 (N_8906,N_8031,N_8257);
xnor U8907 (N_8907,N_8059,N_8205);
and U8908 (N_8908,N_8165,N_8286);
and U8909 (N_8909,N_8300,N_8445);
xnor U8910 (N_8910,N_8454,N_8380);
xor U8911 (N_8911,N_8055,N_8313);
nor U8912 (N_8912,N_8411,N_8289);
nor U8913 (N_8913,N_8374,N_8079);
or U8914 (N_8914,N_8445,N_8106);
xnor U8915 (N_8915,N_8371,N_8168);
and U8916 (N_8916,N_8015,N_8364);
or U8917 (N_8917,N_8233,N_8022);
xnor U8918 (N_8918,N_8039,N_8186);
and U8919 (N_8919,N_8212,N_8119);
and U8920 (N_8920,N_8223,N_8036);
or U8921 (N_8921,N_8206,N_8391);
nand U8922 (N_8922,N_8414,N_8069);
or U8923 (N_8923,N_8202,N_8080);
nand U8924 (N_8924,N_8378,N_8035);
nor U8925 (N_8925,N_8301,N_8065);
and U8926 (N_8926,N_8182,N_8431);
or U8927 (N_8927,N_8160,N_8459);
nor U8928 (N_8928,N_8069,N_8115);
or U8929 (N_8929,N_8463,N_8242);
nor U8930 (N_8930,N_8131,N_8453);
and U8931 (N_8931,N_8154,N_8438);
nand U8932 (N_8932,N_8316,N_8157);
nor U8933 (N_8933,N_8279,N_8387);
xor U8934 (N_8934,N_8335,N_8039);
nor U8935 (N_8935,N_8083,N_8415);
xor U8936 (N_8936,N_8434,N_8288);
or U8937 (N_8937,N_8115,N_8132);
xor U8938 (N_8938,N_8398,N_8307);
or U8939 (N_8939,N_8255,N_8465);
or U8940 (N_8940,N_8346,N_8431);
nor U8941 (N_8941,N_8263,N_8290);
nor U8942 (N_8942,N_8298,N_8113);
nand U8943 (N_8943,N_8452,N_8123);
and U8944 (N_8944,N_8020,N_8235);
or U8945 (N_8945,N_8130,N_8434);
xnor U8946 (N_8946,N_8097,N_8024);
nor U8947 (N_8947,N_8463,N_8005);
or U8948 (N_8948,N_8141,N_8328);
nor U8949 (N_8949,N_8231,N_8210);
nand U8950 (N_8950,N_8315,N_8342);
nand U8951 (N_8951,N_8351,N_8458);
nand U8952 (N_8952,N_8111,N_8345);
and U8953 (N_8953,N_8318,N_8470);
and U8954 (N_8954,N_8126,N_8218);
nand U8955 (N_8955,N_8073,N_8002);
nor U8956 (N_8956,N_8219,N_8279);
and U8957 (N_8957,N_8245,N_8418);
and U8958 (N_8958,N_8318,N_8213);
and U8959 (N_8959,N_8043,N_8091);
nand U8960 (N_8960,N_8444,N_8314);
nand U8961 (N_8961,N_8182,N_8141);
nand U8962 (N_8962,N_8468,N_8097);
and U8963 (N_8963,N_8341,N_8224);
xnor U8964 (N_8964,N_8152,N_8321);
nor U8965 (N_8965,N_8458,N_8391);
xnor U8966 (N_8966,N_8418,N_8145);
and U8967 (N_8967,N_8113,N_8134);
nand U8968 (N_8968,N_8369,N_8012);
and U8969 (N_8969,N_8022,N_8320);
nor U8970 (N_8970,N_8166,N_8260);
and U8971 (N_8971,N_8245,N_8074);
nor U8972 (N_8972,N_8276,N_8242);
xor U8973 (N_8973,N_8005,N_8158);
xnor U8974 (N_8974,N_8346,N_8468);
or U8975 (N_8975,N_8113,N_8068);
and U8976 (N_8976,N_8170,N_8237);
or U8977 (N_8977,N_8002,N_8334);
nor U8978 (N_8978,N_8318,N_8079);
nor U8979 (N_8979,N_8026,N_8181);
and U8980 (N_8980,N_8241,N_8034);
nand U8981 (N_8981,N_8192,N_8442);
nand U8982 (N_8982,N_8261,N_8081);
or U8983 (N_8983,N_8485,N_8235);
nor U8984 (N_8984,N_8323,N_8147);
nor U8985 (N_8985,N_8012,N_8396);
and U8986 (N_8986,N_8496,N_8313);
or U8987 (N_8987,N_8480,N_8234);
xnor U8988 (N_8988,N_8070,N_8437);
or U8989 (N_8989,N_8285,N_8350);
xnor U8990 (N_8990,N_8122,N_8232);
xnor U8991 (N_8991,N_8123,N_8089);
nand U8992 (N_8992,N_8491,N_8124);
nor U8993 (N_8993,N_8077,N_8254);
or U8994 (N_8994,N_8295,N_8196);
xnor U8995 (N_8995,N_8386,N_8143);
nor U8996 (N_8996,N_8495,N_8321);
nor U8997 (N_8997,N_8368,N_8319);
xor U8998 (N_8998,N_8421,N_8493);
and U8999 (N_8999,N_8453,N_8263);
and U9000 (N_9000,N_8605,N_8828);
or U9001 (N_9001,N_8930,N_8973);
and U9002 (N_9002,N_8918,N_8618);
nor U9003 (N_9003,N_8691,N_8634);
or U9004 (N_9004,N_8633,N_8510);
nor U9005 (N_9005,N_8558,N_8699);
nor U9006 (N_9006,N_8928,N_8854);
nor U9007 (N_9007,N_8619,N_8886);
nor U9008 (N_9008,N_8945,N_8833);
nand U9009 (N_9009,N_8888,N_8884);
xnor U9010 (N_9010,N_8941,N_8529);
nor U9011 (N_9011,N_8920,N_8549);
and U9012 (N_9012,N_8859,N_8805);
or U9013 (N_9013,N_8848,N_8810);
nand U9014 (N_9014,N_8927,N_8915);
xor U9015 (N_9015,N_8522,N_8913);
or U9016 (N_9016,N_8844,N_8571);
xor U9017 (N_9017,N_8826,N_8507);
xnor U9018 (N_9018,N_8858,N_8591);
and U9019 (N_9019,N_8625,N_8840);
nor U9020 (N_9020,N_8789,N_8576);
nor U9021 (N_9021,N_8885,N_8792);
xnor U9022 (N_9022,N_8546,N_8984);
nor U9023 (N_9023,N_8539,N_8582);
nand U9024 (N_9024,N_8744,N_8501);
and U9025 (N_9025,N_8610,N_8845);
nor U9026 (N_9026,N_8550,N_8876);
and U9027 (N_9027,N_8819,N_8602);
xnor U9028 (N_9028,N_8584,N_8855);
xnor U9029 (N_9029,N_8748,N_8814);
xor U9030 (N_9030,N_8666,N_8512);
nor U9031 (N_9031,N_8574,N_8604);
nor U9032 (N_9032,N_8897,N_8993);
and U9033 (N_9033,N_8711,N_8516);
xor U9034 (N_9034,N_8745,N_8921);
and U9035 (N_9035,N_8873,N_8939);
nor U9036 (N_9036,N_8705,N_8503);
and U9037 (N_9037,N_8803,N_8670);
nor U9038 (N_9038,N_8590,N_8548);
nand U9039 (N_9039,N_8773,N_8615);
nor U9040 (N_9040,N_8698,N_8688);
and U9041 (N_9041,N_8685,N_8963);
xor U9042 (N_9042,N_8678,N_8836);
or U9043 (N_9043,N_8509,N_8635);
or U9044 (N_9044,N_8659,N_8924);
nand U9045 (N_9045,N_8946,N_8651);
nor U9046 (N_9046,N_8753,N_8552);
and U9047 (N_9047,N_8870,N_8820);
nor U9048 (N_9048,N_8646,N_8629);
or U9049 (N_9049,N_8746,N_8671);
and U9050 (N_9050,N_8543,N_8843);
or U9051 (N_9051,N_8975,N_8616);
and U9052 (N_9052,N_8764,N_8757);
and U9053 (N_9053,N_8761,N_8823);
nand U9054 (N_9054,N_8708,N_8637);
and U9055 (N_9055,N_8595,N_8813);
nor U9056 (N_9056,N_8923,N_8892);
nand U9057 (N_9057,N_8990,N_8573);
or U9058 (N_9058,N_8787,N_8658);
xor U9059 (N_9059,N_8955,N_8747);
nor U9060 (N_9060,N_8934,N_8555);
xnor U9061 (N_9061,N_8736,N_8500);
and U9062 (N_9062,N_8514,N_8566);
nor U9063 (N_9063,N_8725,N_8800);
or U9064 (N_9064,N_8891,N_8727);
or U9065 (N_9065,N_8648,N_8906);
nor U9066 (N_9066,N_8877,N_8758);
nand U9067 (N_9067,N_8653,N_8732);
nor U9068 (N_9068,N_8506,N_8889);
nand U9069 (N_9069,N_8812,N_8991);
or U9070 (N_9070,N_8718,N_8763);
or U9071 (N_9071,N_8997,N_8834);
xnor U9072 (N_9072,N_8720,N_8914);
nor U9073 (N_9073,N_8622,N_8562);
xnor U9074 (N_9074,N_8647,N_8739);
xor U9075 (N_9075,N_8904,N_8531);
and U9076 (N_9076,N_8545,N_8972);
nor U9077 (N_9077,N_8544,N_8690);
nor U9078 (N_9078,N_8650,N_8795);
and U9079 (N_9079,N_8687,N_8811);
or U9080 (N_9080,N_8774,N_8533);
xnor U9081 (N_9081,N_8655,N_8579);
nor U9082 (N_9082,N_8807,N_8933);
xor U9083 (N_9083,N_8673,N_8536);
xor U9084 (N_9084,N_8957,N_8560);
and U9085 (N_9085,N_8704,N_8983);
xnor U9086 (N_9086,N_8614,N_8722);
and U9087 (N_9087,N_8932,N_8701);
nor U9088 (N_9088,N_8970,N_8880);
nor U9089 (N_9089,N_8638,N_8808);
xor U9090 (N_9090,N_8917,N_8961);
nand U9091 (N_9091,N_8608,N_8559);
nor U9092 (N_9092,N_8598,N_8768);
xor U9093 (N_9093,N_8775,N_8741);
and U9094 (N_9094,N_8681,N_8759);
nand U9095 (N_9095,N_8527,N_8665);
nor U9096 (N_9096,N_8528,N_8692);
nand U9097 (N_9097,N_8717,N_8644);
xor U9098 (N_9098,N_8613,N_8967);
nor U9099 (N_9099,N_8860,N_8611);
and U9100 (N_9100,N_8627,N_8968);
nor U9101 (N_9101,N_8797,N_8903);
nand U9102 (N_9102,N_8733,N_8643);
and U9103 (N_9103,N_8847,N_8996);
nor U9104 (N_9104,N_8593,N_8657);
and U9105 (N_9105,N_8816,N_8824);
nor U9106 (N_9106,N_8632,N_8532);
nand U9107 (N_9107,N_8857,N_8989);
nand U9108 (N_9108,N_8964,N_8743);
nand U9109 (N_9109,N_8785,N_8935);
nor U9110 (N_9110,N_8538,N_8564);
or U9111 (N_9111,N_8907,N_8518);
or U9112 (N_9112,N_8667,N_8603);
nand U9113 (N_9113,N_8570,N_8977);
and U9114 (N_9114,N_8652,N_8976);
xor U9115 (N_9115,N_8992,N_8750);
nor U9116 (N_9116,N_8829,N_8583);
and U9117 (N_9117,N_8982,N_8675);
and U9118 (N_9118,N_8557,N_8664);
nor U9119 (N_9119,N_8922,N_8979);
xnor U9120 (N_9120,N_8954,N_8515);
nor U9121 (N_9121,N_8686,N_8542);
xor U9122 (N_9122,N_8995,N_8594);
nor U9123 (N_9123,N_8724,N_8909);
nand U9124 (N_9124,N_8796,N_8881);
xor U9125 (N_9125,N_8999,N_8709);
or U9126 (N_9126,N_8771,N_8521);
or U9127 (N_9127,N_8554,N_8537);
nand U9128 (N_9128,N_8953,N_8567);
xnor U9129 (N_9129,N_8798,N_8723);
nand U9130 (N_9130,N_8517,N_8872);
or U9131 (N_9131,N_8878,N_8809);
xor U9132 (N_9132,N_8730,N_8883);
and U9133 (N_9133,N_8871,N_8962);
or U9134 (N_9134,N_8700,N_8772);
and U9135 (N_9135,N_8609,N_8818);
or U9136 (N_9136,N_8817,N_8835);
xnor U9137 (N_9137,N_8988,N_8726);
nor U9138 (N_9138,N_8580,N_8766);
and U9139 (N_9139,N_8719,N_8682);
nor U9140 (N_9140,N_8985,N_8825);
xnor U9141 (N_9141,N_8656,N_8534);
or U9142 (N_9142,N_8965,N_8696);
and U9143 (N_9143,N_8765,N_8980);
xor U9144 (N_9144,N_8874,N_8944);
or U9145 (N_9145,N_8697,N_8721);
or U9146 (N_9146,N_8793,N_8535);
nor U9147 (N_9147,N_8754,N_8851);
nand U9148 (N_9148,N_8680,N_8940);
nor U9149 (N_9149,N_8863,N_8950);
nand U9150 (N_9150,N_8960,N_8879);
nand U9151 (N_9151,N_8601,N_8563);
nand U9152 (N_9152,N_8596,N_8641);
and U9153 (N_9153,N_8713,N_8861);
nand U9154 (N_9154,N_8827,N_8504);
nand U9155 (N_9155,N_8887,N_8790);
xnor U9156 (N_9156,N_8856,N_8791);
nor U9157 (N_9157,N_8842,N_8974);
and U9158 (N_9158,N_8752,N_8943);
and U9159 (N_9159,N_8735,N_8575);
and U9160 (N_9160,N_8662,N_8526);
or U9161 (N_9161,N_8606,N_8908);
nor U9162 (N_9162,N_8998,N_8931);
nor U9163 (N_9163,N_8617,N_8728);
nand U9164 (N_9164,N_8867,N_8645);
nand U9165 (N_9165,N_8868,N_8540);
nand U9166 (N_9166,N_8631,N_8952);
xor U9167 (N_9167,N_8640,N_8706);
or U9168 (N_9168,N_8951,N_8987);
xnor U9169 (N_9169,N_8734,N_8783);
and U9170 (N_9170,N_8737,N_8502);
nor U9171 (N_9171,N_8956,N_8949);
and U9172 (N_9172,N_8513,N_8551);
nor U9173 (N_9173,N_8929,N_8683);
and U9174 (N_9174,N_8942,N_8694);
or U9175 (N_9175,N_8779,N_8505);
and U9176 (N_9176,N_8839,N_8672);
or U9177 (N_9177,N_8519,N_8849);
nor U9178 (N_9178,N_8636,N_8893);
nor U9179 (N_9179,N_8882,N_8902);
xnor U9180 (N_9180,N_8780,N_8703);
nand U9181 (N_9181,N_8969,N_8898);
nor U9182 (N_9182,N_8801,N_8905);
and U9183 (N_9183,N_8896,N_8578);
or U9184 (N_9184,N_8778,N_8838);
and U9185 (N_9185,N_8702,N_8986);
or U9186 (N_9186,N_8804,N_8716);
nor U9187 (N_9187,N_8677,N_8523);
xnor U9188 (N_9188,N_8679,N_8668);
nor U9189 (N_9189,N_8815,N_8612);
and U9190 (N_9190,N_8948,N_8894);
or U9191 (N_9191,N_8715,N_8585);
or U9192 (N_9192,N_8832,N_8910);
or U9193 (N_9193,N_8926,N_8966);
or U9194 (N_9194,N_8577,N_8959);
and U9195 (N_9195,N_8553,N_8769);
nor U9196 (N_9196,N_8837,N_8831);
nand U9197 (N_9197,N_8654,N_8740);
nor U9198 (N_9198,N_8695,N_8572);
nand U9199 (N_9199,N_8588,N_8830);
and U9200 (N_9200,N_8742,N_8524);
or U9201 (N_9201,N_8788,N_8925);
xor U9202 (N_9202,N_8846,N_8581);
nand U9203 (N_9203,N_8630,N_8981);
nand U9204 (N_9204,N_8911,N_8895);
nand U9205 (N_9205,N_8869,N_8639);
or U9206 (N_9206,N_8731,N_8782);
nand U9207 (N_9207,N_8628,N_8541);
or U9208 (N_9208,N_8511,N_8669);
or U9209 (N_9209,N_8776,N_8770);
and U9210 (N_9210,N_8592,N_8806);
nor U9211 (N_9211,N_8508,N_8755);
and U9212 (N_9212,N_8802,N_8621);
or U9213 (N_9213,N_8589,N_8714);
or U9214 (N_9214,N_8561,N_8938);
xnor U9215 (N_9215,N_8597,N_8547);
nor U9216 (N_9216,N_8684,N_8799);
nand U9217 (N_9217,N_8749,N_8822);
or U9218 (N_9218,N_8899,N_8864);
or U9219 (N_9219,N_8676,N_8781);
xnor U9220 (N_9220,N_8568,N_8600);
or U9221 (N_9221,N_8994,N_8937);
nor U9222 (N_9222,N_8852,N_8663);
and U9223 (N_9223,N_8565,N_8794);
and U9224 (N_9224,N_8620,N_8916);
nand U9225 (N_9225,N_8569,N_8865);
and U9226 (N_9226,N_8919,N_8841);
and U9227 (N_9227,N_8623,N_8890);
and U9228 (N_9228,N_8912,N_8866);
nor U9229 (N_9229,N_8530,N_8821);
xor U9230 (N_9230,N_8756,N_8649);
xnor U9231 (N_9231,N_8710,N_8875);
and U9232 (N_9232,N_8520,N_8900);
and U9233 (N_9233,N_8738,N_8901);
nand U9234 (N_9234,N_8586,N_8971);
or U9235 (N_9235,N_8599,N_8587);
nand U9236 (N_9236,N_8674,N_8556);
or U9237 (N_9237,N_8958,N_8786);
and U9238 (N_9238,N_8693,N_8689);
xor U9239 (N_9239,N_8751,N_8712);
nand U9240 (N_9240,N_8642,N_8707);
and U9241 (N_9241,N_8525,N_8626);
and U9242 (N_9242,N_8767,N_8947);
or U9243 (N_9243,N_8862,N_8624);
xor U9244 (N_9244,N_8784,N_8978);
nor U9245 (N_9245,N_8853,N_8661);
nand U9246 (N_9246,N_8607,N_8777);
xor U9247 (N_9247,N_8660,N_8729);
nor U9248 (N_9248,N_8850,N_8760);
or U9249 (N_9249,N_8762,N_8936);
nand U9250 (N_9250,N_8723,N_8732);
or U9251 (N_9251,N_8921,N_8665);
xnor U9252 (N_9252,N_8562,N_8512);
or U9253 (N_9253,N_8797,N_8624);
nor U9254 (N_9254,N_8622,N_8767);
or U9255 (N_9255,N_8560,N_8894);
nor U9256 (N_9256,N_8999,N_8828);
xor U9257 (N_9257,N_8964,N_8665);
nor U9258 (N_9258,N_8662,N_8667);
or U9259 (N_9259,N_8614,N_8764);
and U9260 (N_9260,N_8793,N_8918);
and U9261 (N_9261,N_8782,N_8803);
nor U9262 (N_9262,N_8699,N_8963);
or U9263 (N_9263,N_8555,N_8827);
or U9264 (N_9264,N_8716,N_8926);
nand U9265 (N_9265,N_8940,N_8540);
nand U9266 (N_9266,N_8772,N_8535);
nor U9267 (N_9267,N_8627,N_8572);
and U9268 (N_9268,N_8967,N_8669);
and U9269 (N_9269,N_8873,N_8911);
xnor U9270 (N_9270,N_8639,N_8553);
and U9271 (N_9271,N_8587,N_8827);
or U9272 (N_9272,N_8733,N_8577);
nor U9273 (N_9273,N_8977,N_8719);
nor U9274 (N_9274,N_8717,N_8807);
and U9275 (N_9275,N_8953,N_8967);
and U9276 (N_9276,N_8675,N_8656);
and U9277 (N_9277,N_8737,N_8825);
nor U9278 (N_9278,N_8707,N_8660);
nand U9279 (N_9279,N_8945,N_8817);
nor U9280 (N_9280,N_8720,N_8594);
nor U9281 (N_9281,N_8502,N_8622);
nor U9282 (N_9282,N_8796,N_8992);
xor U9283 (N_9283,N_8613,N_8651);
nand U9284 (N_9284,N_8960,N_8606);
and U9285 (N_9285,N_8861,N_8732);
nor U9286 (N_9286,N_8966,N_8659);
xor U9287 (N_9287,N_8818,N_8837);
nor U9288 (N_9288,N_8976,N_8800);
xnor U9289 (N_9289,N_8901,N_8797);
nand U9290 (N_9290,N_8843,N_8504);
nand U9291 (N_9291,N_8766,N_8591);
or U9292 (N_9292,N_8817,N_8987);
and U9293 (N_9293,N_8890,N_8815);
nand U9294 (N_9294,N_8913,N_8586);
or U9295 (N_9295,N_8673,N_8794);
and U9296 (N_9296,N_8783,N_8511);
and U9297 (N_9297,N_8792,N_8949);
or U9298 (N_9298,N_8534,N_8719);
and U9299 (N_9299,N_8779,N_8960);
and U9300 (N_9300,N_8510,N_8690);
nor U9301 (N_9301,N_8947,N_8805);
and U9302 (N_9302,N_8590,N_8514);
and U9303 (N_9303,N_8941,N_8584);
nand U9304 (N_9304,N_8584,N_8506);
or U9305 (N_9305,N_8586,N_8530);
and U9306 (N_9306,N_8889,N_8887);
or U9307 (N_9307,N_8948,N_8876);
xor U9308 (N_9308,N_8620,N_8599);
and U9309 (N_9309,N_8605,N_8888);
and U9310 (N_9310,N_8767,N_8840);
xor U9311 (N_9311,N_8829,N_8644);
nor U9312 (N_9312,N_8582,N_8651);
nand U9313 (N_9313,N_8733,N_8535);
nand U9314 (N_9314,N_8773,N_8863);
xnor U9315 (N_9315,N_8866,N_8871);
xor U9316 (N_9316,N_8687,N_8798);
xor U9317 (N_9317,N_8619,N_8631);
and U9318 (N_9318,N_8947,N_8675);
xor U9319 (N_9319,N_8565,N_8879);
nor U9320 (N_9320,N_8948,N_8536);
and U9321 (N_9321,N_8959,N_8683);
xnor U9322 (N_9322,N_8689,N_8801);
nand U9323 (N_9323,N_8862,N_8836);
and U9324 (N_9324,N_8709,N_8640);
xor U9325 (N_9325,N_8501,N_8978);
nand U9326 (N_9326,N_8642,N_8882);
xor U9327 (N_9327,N_8635,N_8599);
and U9328 (N_9328,N_8643,N_8674);
nor U9329 (N_9329,N_8584,N_8968);
nor U9330 (N_9330,N_8865,N_8931);
xnor U9331 (N_9331,N_8726,N_8569);
nand U9332 (N_9332,N_8569,N_8987);
xnor U9333 (N_9333,N_8580,N_8724);
nand U9334 (N_9334,N_8912,N_8650);
nor U9335 (N_9335,N_8794,N_8505);
xnor U9336 (N_9336,N_8957,N_8879);
nand U9337 (N_9337,N_8873,N_8680);
and U9338 (N_9338,N_8935,N_8834);
and U9339 (N_9339,N_8914,N_8989);
nor U9340 (N_9340,N_8831,N_8783);
and U9341 (N_9341,N_8524,N_8849);
nor U9342 (N_9342,N_8980,N_8672);
nor U9343 (N_9343,N_8657,N_8975);
or U9344 (N_9344,N_8857,N_8710);
nand U9345 (N_9345,N_8954,N_8891);
nor U9346 (N_9346,N_8582,N_8994);
or U9347 (N_9347,N_8638,N_8876);
or U9348 (N_9348,N_8990,N_8861);
xor U9349 (N_9349,N_8845,N_8742);
and U9350 (N_9350,N_8816,N_8792);
nand U9351 (N_9351,N_8898,N_8805);
nand U9352 (N_9352,N_8766,N_8936);
nor U9353 (N_9353,N_8918,N_8983);
nand U9354 (N_9354,N_8991,N_8922);
and U9355 (N_9355,N_8959,N_8945);
or U9356 (N_9356,N_8627,N_8521);
nand U9357 (N_9357,N_8566,N_8976);
nand U9358 (N_9358,N_8538,N_8607);
xnor U9359 (N_9359,N_8953,N_8710);
nor U9360 (N_9360,N_8756,N_8949);
nor U9361 (N_9361,N_8549,N_8598);
or U9362 (N_9362,N_8784,N_8511);
xor U9363 (N_9363,N_8978,N_8890);
nor U9364 (N_9364,N_8708,N_8694);
nand U9365 (N_9365,N_8917,N_8597);
or U9366 (N_9366,N_8892,N_8613);
or U9367 (N_9367,N_8697,N_8666);
nand U9368 (N_9368,N_8508,N_8776);
xnor U9369 (N_9369,N_8700,N_8943);
and U9370 (N_9370,N_8987,N_8637);
and U9371 (N_9371,N_8829,N_8844);
xor U9372 (N_9372,N_8903,N_8693);
nor U9373 (N_9373,N_8645,N_8745);
nor U9374 (N_9374,N_8670,N_8931);
xor U9375 (N_9375,N_8814,N_8817);
or U9376 (N_9376,N_8505,N_8898);
and U9377 (N_9377,N_8612,N_8853);
xnor U9378 (N_9378,N_8713,N_8948);
nor U9379 (N_9379,N_8768,N_8664);
nor U9380 (N_9380,N_8868,N_8803);
nand U9381 (N_9381,N_8692,N_8803);
nor U9382 (N_9382,N_8792,N_8552);
nor U9383 (N_9383,N_8586,N_8599);
or U9384 (N_9384,N_8525,N_8628);
nor U9385 (N_9385,N_8569,N_8692);
nand U9386 (N_9386,N_8912,N_8522);
nand U9387 (N_9387,N_8641,N_8688);
and U9388 (N_9388,N_8986,N_8912);
nor U9389 (N_9389,N_8535,N_8611);
xnor U9390 (N_9390,N_8849,N_8730);
xor U9391 (N_9391,N_8985,N_8592);
nor U9392 (N_9392,N_8845,N_8884);
and U9393 (N_9393,N_8784,N_8530);
xor U9394 (N_9394,N_8547,N_8859);
nand U9395 (N_9395,N_8518,N_8589);
nor U9396 (N_9396,N_8756,N_8951);
nor U9397 (N_9397,N_8885,N_8799);
or U9398 (N_9398,N_8597,N_8700);
or U9399 (N_9399,N_8768,N_8783);
or U9400 (N_9400,N_8510,N_8620);
xnor U9401 (N_9401,N_8910,N_8523);
nand U9402 (N_9402,N_8807,N_8975);
and U9403 (N_9403,N_8998,N_8932);
and U9404 (N_9404,N_8534,N_8846);
and U9405 (N_9405,N_8970,N_8576);
nor U9406 (N_9406,N_8916,N_8538);
or U9407 (N_9407,N_8791,N_8858);
and U9408 (N_9408,N_8790,N_8548);
xnor U9409 (N_9409,N_8823,N_8877);
nand U9410 (N_9410,N_8903,N_8613);
nor U9411 (N_9411,N_8964,N_8812);
nor U9412 (N_9412,N_8865,N_8968);
or U9413 (N_9413,N_8767,N_8681);
nor U9414 (N_9414,N_8645,N_8876);
nand U9415 (N_9415,N_8812,N_8552);
nor U9416 (N_9416,N_8517,N_8692);
nor U9417 (N_9417,N_8620,N_8747);
nor U9418 (N_9418,N_8975,N_8932);
xnor U9419 (N_9419,N_8562,N_8711);
and U9420 (N_9420,N_8940,N_8810);
nor U9421 (N_9421,N_8968,N_8593);
nor U9422 (N_9422,N_8504,N_8838);
xor U9423 (N_9423,N_8686,N_8982);
or U9424 (N_9424,N_8958,N_8696);
xor U9425 (N_9425,N_8562,N_8933);
nand U9426 (N_9426,N_8794,N_8716);
and U9427 (N_9427,N_8645,N_8622);
nand U9428 (N_9428,N_8920,N_8961);
nand U9429 (N_9429,N_8843,N_8539);
or U9430 (N_9430,N_8640,N_8684);
nand U9431 (N_9431,N_8614,N_8954);
and U9432 (N_9432,N_8911,N_8751);
and U9433 (N_9433,N_8550,N_8572);
nor U9434 (N_9434,N_8902,N_8759);
nor U9435 (N_9435,N_8536,N_8628);
and U9436 (N_9436,N_8620,N_8567);
xnor U9437 (N_9437,N_8629,N_8753);
xnor U9438 (N_9438,N_8529,N_8531);
or U9439 (N_9439,N_8624,N_8589);
nand U9440 (N_9440,N_8734,N_8813);
nand U9441 (N_9441,N_8901,N_8713);
nor U9442 (N_9442,N_8931,N_8657);
or U9443 (N_9443,N_8885,N_8983);
or U9444 (N_9444,N_8677,N_8542);
and U9445 (N_9445,N_8644,N_8625);
xor U9446 (N_9446,N_8984,N_8882);
nor U9447 (N_9447,N_8699,N_8712);
or U9448 (N_9448,N_8949,N_8957);
nand U9449 (N_9449,N_8681,N_8995);
nand U9450 (N_9450,N_8848,N_8673);
and U9451 (N_9451,N_8603,N_8941);
or U9452 (N_9452,N_8834,N_8686);
nor U9453 (N_9453,N_8646,N_8616);
xor U9454 (N_9454,N_8693,N_8743);
xor U9455 (N_9455,N_8899,N_8703);
xnor U9456 (N_9456,N_8711,N_8789);
and U9457 (N_9457,N_8913,N_8618);
nor U9458 (N_9458,N_8524,N_8913);
nor U9459 (N_9459,N_8928,N_8612);
or U9460 (N_9460,N_8626,N_8919);
or U9461 (N_9461,N_8745,N_8802);
or U9462 (N_9462,N_8672,N_8669);
nor U9463 (N_9463,N_8741,N_8666);
nand U9464 (N_9464,N_8760,N_8896);
or U9465 (N_9465,N_8746,N_8546);
xor U9466 (N_9466,N_8900,N_8840);
xnor U9467 (N_9467,N_8919,N_8987);
nor U9468 (N_9468,N_8915,N_8510);
nor U9469 (N_9469,N_8542,N_8740);
or U9470 (N_9470,N_8852,N_8593);
or U9471 (N_9471,N_8669,N_8990);
nand U9472 (N_9472,N_8679,N_8818);
nor U9473 (N_9473,N_8612,N_8927);
xnor U9474 (N_9474,N_8928,N_8857);
nand U9475 (N_9475,N_8805,N_8506);
nand U9476 (N_9476,N_8690,N_8949);
and U9477 (N_9477,N_8764,N_8894);
xnor U9478 (N_9478,N_8835,N_8559);
nand U9479 (N_9479,N_8844,N_8501);
and U9480 (N_9480,N_8847,N_8658);
xor U9481 (N_9481,N_8641,N_8949);
or U9482 (N_9482,N_8865,N_8978);
and U9483 (N_9483,N_8882,N_8600);
and U9484 (N_9484,N_8501,N_8635);
xor U9485 (N_9485,N_8650,N_8596);
or U9486 (N_9486,N_8986,N_8661);
or U9487 (N_9487,N_8656,N_8876);
or U9488 (N_9488,N_8899,N_8911);
nand U9489 (N_9489,N_8716,N_8980);
and U9490 (N_9490,N_8529,N_8501);
nand U9491 (N_9491,N_8526,N_8835);
xor U9492 (N_9492,N_8886,N_8931);
nand U9493 (N_9493,N_8852,N_8529);
nand U9494 (N_9494,N_8896,N_8963);
nor U9495 (N_9495,N_8721,N_8640);
nand U9496 (N_9496,N_8762,N_8502);
and U9497 (N_9497,N_8624,N_8693);
or U9498 (N_9498,N_8656,N_8814);
nor U9499 (N_9499,N_8812,N_8997);
or U9500 (N_9500,N_9404,N_9004);
nor U9501 (N_9501,N_9419,N_9016);
nand U9502 (N_9502,N_9321,N_9093);
nand U9503 (N_9503,N_9086,N_9116);
and U9504 (N_9504,N_9352,N_9384);
xnor U9505 (N_9505,N_9395,N_9109);
and U9506 (N_9506,N_9166,N_9036);
nor U9507 (N_9507,N_9403,N_9486);
or U9508 (N_9508,N_9262,N_9148);
or U9509 (N_9509,N_9408,N_9247);
xor U9510 (N_9510,N_9153,N_9240);
nor U9511 (N_9511,N_9105,N_9013);
nor U9512 (N_9512,N_9470,N_9345);
xnor U9513 (N_9513,N_9229,N_9121);
nor U9514 (N_9514,N_9494,N_9103);
nor U9515 (N_9515,N_9149,N_9488);
nor U9516 (N_9516,N_9221,N_9396);
or U9517 (N_9517,N_9040,N_9054);
xor U9518 (N_9518,N_9442,N_9052);
and U9519 (N_9519,N_9219,N_9206);
nor U9520 (N_9520,N_9445,N_9382);
or U9521 (N_9521,N_9473,N_9430);
xor U9522 (N_9522,N_9208,N_9021);
nor U9523 (N_9523,N_9428,N_9122);
or U9524 (N_9524,N_9250,N_9427);
xnor U9525 (N_9525,N_9160,N_9475);
nor U9526 (N_9526,N_9235,N_9193);
xor U9527 (N_9527,N_9426,N_9058);
nor U9528 (N_9528,N_9253,N_9353);
or U9529 (N_9529,N_9409,N_9179);
and U9530 (N_9530,N_9306,N_9481);
nand U9531 (N_9531,N_9326,N_9406);
nor U9532 (N_9532,N_9386,N_9078);
or U9533 (N_9533,N_9362,N_9070);
and U9534 (N_9534,N_9331,N_9405);
nand U9535 (N_9535,N_9009,N_9150);
xnor U9536 (N_9536,N_9401,N_9059);
and U9537 (N_9537,N_9023,N_9022);
xnor U9538 (N_9538,N_9328,N_9100);
or U9539 (N_9539,N_9198,N_9459);
nand U9540 (N_9540,N_9271,N_9196);
or U9541 (N_9541,N_9480,N_9279);
xor U9542 (N_9542,N_9107,N_9090);
or U9543 (N_9543,N_9292,N_9431);
nor U9544 (N_9544,N_9187,N_9171);
and U9545 (N_9545,N_9195,N_9311);
nor U9546 (N_9546,N_9483,N_9260);
nor U9547 (N_9547,N_9172,N_9118);
nand U9548 (N_9548,N_9051,N_9334);
and U9549 (N_9549,N_9361,N_9478);
nor U9550 (N_9550,N_9266,N_9344);
and U9551 (N_9551,N_9393,N_9295);
and U9552 (N_9552,N_9019,N_9358);
or U9553 (N_9553,N_9413,N_9293);
or U9554 (N_9554,N_9484,N_9177);
and U9555 (N_9555,N_9389,N_9457);
nand U9556 (N_9556,N_9376,N_9068);
or U9557 (N_9557,N_9067,N_9239);
nand U9558 (N_9558,N_9324,N_9377);
and U9559 (N_9559,N_9290,N_9434);
xor U9560 (N_9560,N_9270,N_9178);
nor U9561 (N_9561,N_9071,N_9197);
xnor U9562 (N_9562,N_9460,N_9137);
nand U9563 (N_9563,N_9163,N_9463);
and U9564 (N_9564,N_9055,N_9447);
nand U9565 (N_9565,N_9073,N_9391);
nor U9566 (N_9566,N_9412,N_9299);
xnor U9567 (N_9567,N_9087,N_9053);
and U9568 (N_9568,N_9356,N_9210);
xnor U9569 (N_9569,N_9251,N_9001);
nand U9570 (N_9570,N_9330,N_9175);
and U9571 (N_9571,N_9225,N_9482);
nand U9572 (N_9572,N_9159,N_9114);
nor U9573 (N_9573,N_9038,N_9437);
and U9574 (N_9574,N_9283,N_9174);
xor U9575 (N_9575,N_9030,N_9056);
or U9576 (N_9576,N_9234,N_9307);
and U9577 (N_9577,N_9005,N_9258);
nand U9578 (N_9578,N_9048,N_9249);
nor U9579 (N_9579,N_9346,N_9259);
xor U9580 (N_9580,N_9216,N_9095);
nor U9581 (N_9581,N_9296,N_9144);
or U9582 (N_9582,N_9061,N_9242);
xnor U9583 (N_9583,N_9043,N_9433);
xor U9584 (N_9584,N_9367,N_9106);
nand U9585 (N_9585,N_9066,N_9398);
nand U9586 (N_9586,N_9257,N_9244);
nor U9587 (N_9587,N_9444,N_9273);
and U9588 (N_9588,N_9278,N_9026);
or U9589 (N_9589,N_9049,N_9161);
and U9590 (N_9590,N_9468,N_9372);
and U9591 (N_9591,N_9320,N_9065);
and U9592 (N_9592,N_9411,N_9044);
nor U9593 (N_9593,N_9131,N_9466);
nand U9594 (N_9594,N_9399,N_9017);
and U9595 (N_9595,N_9467,N_9498);
and U9596 (N_9596,N_9094,N_9471);
or U9597 (N_9597,N_9332,N_9135);
xnor U9598 (N_9598,N_9057,N_9209);
xnor U9599 (N_9599,N_9015,N_9223);
or U9600 (N_9600,N_9455,N_9339);
and U9601 (N_9601,N_9097,N_9085);
xor U9602 (N_9602,N_9380,N_9479);
nand U9603 (N_9603,N_9381,N_9316);
and U9604 (N_9604,N_9317,N_9034);
nor U9605 (N_9605,N_9343,N_9162);
or U9606 (N_9606,N_9452,N_9167);
xor U9607 (N_9607,N_9451,N_9485);
nand U9608 (N_9608,N_9421,N_9129);
nor U9609 (N_9609,N_9375,N_9072);
nand U9610 (N_9610,N_9336,N_9465);
nand U9611 (N_9611,N_9281,N_9374);
nor U9612 (N_9612,N_9417,N_9120);
xor U9613 (N_9613,N_9294,N_9300);
and U9614 (N_9614,N_9062,N_9327);
and U9615 (N_9615,N_9383,N_9370);
or U9616 (N_9616,N_9446,N_9314);
nand U9617 (N_9617,N_9269,N_9415);
xnor U9618 (N_9618,N_9154,N_9002);
xor U9619 (N_9619,N_9212,N_9474);
and U9620 (N_9620,N_9400,N_9138);
and U9621 (N_9621,N_9099,N_9369);
and U9622 (N_9622,N_9337,N_9201);
and U9623 (N_9623,N_9014,N_9477);
nand U9624 (N_9624,N_9499,N_9449);
and U9625 (N_9625,N_9082,N_9199);
nor U9626 (N_9626,N_9101,N_9289);
nor U9627 (N_9627,N_9441,N_9190);
nand U9628 (N_9628,N_9394,N_9132);
xnor U9629 (N_9629,N_9497,N_9489);
or U9630 (N_9630,N_9214,N_9211);
nand U9631 (N_9631,N_9156,N_9136);
nand U9632 (N_9632,N_9265,N_9063);
nor U9633 (N_9633,N_9047,N_9272);
nand U9634 (N_9634,N_9341,N_9487);
xor U9635 (N_9635,N_9350,N_9155);
and U9636 (N_9636,N_9464,N_9338);
nand U9637 (N_9637,N_9092,N_9333);
nor U9638 (N_9638,N_9123,N_9108);
xor U9639 (N_9639,N_9089,N_9165);
nor U9640 (N_9640,N_9207,N_9205);
and U9641 (N_9641,N_9491,N_9158);
xnor U9642 (N_9642,N_9139,N_9126);
and U9643 (N_9643,N_9079,N_9151);
or U9644 (N_9644,N_9102,N_9425);
and U9645 (N_9645,N_9416,N_9329);
and U9646 (N_9646,N_9371,N_9305);
xnor U9647 (N_9647,N_9228,N_9436);
nor U9648 (N_9648,N_9032,N_9186);
xnor U9649 (N_9649,N_9230,N_9322);
nor U9650 (N_9650,N_9182,N_9168);
nand U9651 (N_9651,N_9303,N_9077);
nand U9652 (N_9652,N_9111,N_9088);
xnor U9653 (N_9653,N_9390,N_9076);
nor U9654 (N_9654,N_9402,N_9349);
or U9655 (N_9655,N_9110,N_9096);
and U9656 (N_9656,N_9238,N_9011);
nor U9657 (N_9657,N_9181,N_9145);
xor U9658 (N_9658,N_9227,N_9191);
xor U9659 (N_9659,N_9288,N_9081);
xnor U9660 (N_9660,N_9276,N_9119);
nand U9661 (N_9661,N_9368,N_9098);
nor U9662 (N_9662,N_9218,N_9192);
xnor U9663 (N_9663,N_9232,N_9440);
or U9664 (N_9664,N_9313,N_9142);
and U9665 (N_9665,N_9462,N_9170);
nor U9666 (N_9666,N_9027,N_9157);
nand U9667 (N_9667,N_9046,N_9236);
and U9668 (N_9668,N_9008,N_9282);
nor U9669 (N_9669,N_9217,N_9037);
nor U9670 (N_9670,N_9185,N_9423);
nand U9671 (N_9671,N_9379,N_9202);
nand U9672 (N_9672,N_9133,N_9203);
nand U9673 (N_9673,N_9366,N_9490);
nor U9674 (N_9674,N_9256,N_9140);
xor U9675 (N_9675,N_9018,N_9176);
nand U9676 (N_9676,N_9439,N_9237);
and U9677 (N_9677,N_9435,N_9173);
or U9678 (N_9678,N_9115,N_9310);
or U9679 (N_9679,N_9143,N_9285);
nand U9680 (N_9680,N_9012,N_9064);
nand U9681 (N_9681,N_9496,N_9222);
nor U9682 (N_9682,N_9280,N_9297);
nor U9683 (N_9683,N_9277,N_9495);
and U9684 (N_9684,N_9388,N_9267);
and U9685 (N_9685,N_9308,N_9254);
nor U9686 (N_9686,N_9125,N_9233);
nand U9687 (N_9687,N_9113,N_9493);
nor U9688 (N_9688,N_9385,N_9104);
or U9689 (N_9689,N_9342,N_9152);
and U9690 (N_9690,N_9184,N_9028);
or U9691 (N_9691,N_9302,N_9450);
nor U9692 (N_9692,N_9365,N_9080);
or U9693 (N_9693,N_9291,N_9141);
or U9694 (N_9694,N_9252,N_9397);
nor U9695 (N_9695,N_9127,N_9422);
xnor U9696 (N_9696,N_9128,N_9215);
nor U9697 (N_9697,N_9351,N_9304);
and U9698 (N_9698,N_9245,N_9241);
and U9699 (N_9699,N_9169,N_9194);
nand U9700 (N_9700,N_9183,N_9274);
nand U9701 (N_9701,N_9204,N_9373);
xnor U9702 (N_9702,N_9407,N_9432);
nor U9703 (N_9703,N_9117,N_9246);
nor U9704 (N_9704,N_9354,N_9224);
nand U9705 (N_9705,N_9213,N_9042);
and U9706 (N_9706,N_9045,N_9325);
xor U9707 (N_9707,N_9024,N_9000);
or U9708 (N_9708,N_9006,N_9231);
and U9709 (N_9709,N_9033,N_9312);
and U9710 (N_9710,N_9248,N_9226);
or U9711 (N_9711,N_9472,N_9387);
nand U9712 (N_9712,N_9323,N_9130);
nand U9713 (N_9713,N_9284,N_9091);
nand U9714 (N_9714,N_9200,N_9360);
nand U9715 (N_9715,N_9335,N_9050);
and U9716 (N_9716,N_9264,N_9420);
and U9717 (N_9717,N_9364,N_9084);
or U9718 (N_9718,N_9458,N_9039);
xor U9719 (N_9719,N_9418,N_9456);
nand U9720 (N_9720,N_9355,N_9319);
or U9721 (N_9721,N_9020,N_9448);
nor U9722 (N_9722,N_9454,N_9029);
nor U9723 (N_9723,N_9189,N_9424);
nor U9724 (N_9724,N_9378,N_9083);
nand U9725 (N_9725,N_9359,N_9443);
and U9726 (N_9726,N_9069,N_9261);
or U9727 (N_9727,N_9429,N_9414);
or U9728 (N_9728,N_9003,N_9309);
nand U9729 (N_9729,N_9074,N_9124);
or U9730 (N_9730,N_9041,N_9243);
nand U9731 (N_9731,N_9492,N_9268);
xor U9732 (N_9732,N_9318,N_9340);
nand U9733 (N_9733,N_9031,N_9287);
or U9734 (N_9734,N_9220,N_9075);
or U9735 (N_9735,N_9188,N_9060);
nand U9736 (N_9736,N_9180,N_9146);
or U9737 (N_9737,N_9025,N_9315);
or U9738 (N_9738,N_9476,N_9286);
and U9739 (N_9739,N_9275,N_9461);
nor U9740 (N_9740,N_9255,N_9010);
or U9741 (N_9741,N_9410,N_9007);
nand U9742 (N_9742,N_9469,N_9392);
nand U9743 (N_9743,N_9147,N_9438);
and U9744 (N_9744,N_9363,N_9348);
and U9745 (N_9745,N_9298,N_9134);
and U9746 (N_9746,N_9347,N_9035);
nand U9747 (N_9747,N_9164,N_9453);
nor U9748 (N_9748,N_9112,N_9301);
nand U9749 (N_9749,N_9263,N_9357);
xnor U9750 (N_9750,N_9097,N_9326);
nor U9751 (N_9751,N_9001,N_9308);
or U9752 (N_9752,N_9418,N_9076);
and U9753 (N_9753,N_9399,N_9101);
and U9754 (N_9754,N_9174,N_9326);
nor U9755 (N_9755,N_9344,N_9179);
nor U9756 (N_9756,N_9133,N_9423);
and U9757 (N_9757,N_9370,N_9300);
xnor U9758 (N_9758,N_9410,N_9334);
or U9759 (N_9759,N_9031,N_9029);
or U9760 (N_9760,N_9385,N_9006);
nand U9761 (N_9761,N_9331,N_9309);
and U9762 (N_9762,N_9366,N_9111);
nand U9763 (N_9763,N_9018,N_9429);
nand U9764 (N_9764,N_9026,N_9224);
nor U9765 (N_9765,N_9203,N_9322);
nand U9766 (N_9766,N_9402,N_9343);
and U9767 (N_9767,N_9294,N_9137);
nand U9768 (N_9768,N_9054,N_9164);
or U9769 (N_9769,N_9376,N_9208);
nand U9770 (N_9770,N_9131,N_9199);
or U9771 (N_9771,N_9408,N_9153);
and U9772 (N_9772,N_9354,N_9068);
xor U9773 (N_9773,N_9281,N_9462);
xor U9774 (N_9774,N_9369,N_9490);
nand U9775 (N_9775,N_9169,N_9438);
and U9776 (N_9776,N_9475,N_9072);
nand U9777 (N_9777,N_9462,N_9227);
nand U9778 (N_9778,N_9327,N_9277);
nor U9779 (N_9779,N_9156,N_9073);
and U9780 (N_9780,N_9351,N_9407);
and U9781 (N_9781,N_9082,N_9383);
or U9782 (N_9782,N_9179,N_9011);
and U9783 (N_9783,N_9423,N_9479);
and U9784 (N_9784,N_9238,N_9054);
nand U9785 (N_9785,N_9344,N_9411);
or U9786 (N_9786,N_9263,N_9172);
and U9787 (N_9787,N_9113,N_9359);
nor U9788 (N_9788,N_9409,N_9462);
or U9789 (N_9789,N_9227,N_9331);
xor U9790 (N_9790,N_9434,N_9197);
xor U9791 (N_9791,N_9386,N_9481);
or U9792 (N_9792,N_9467,N_9302);
and U9793 (N_9793,N_9389,N_9383);
or U9794 (N_9794,N_9418,N_9289);
nor U9795 (N_9795,N_9168,N_9385);
nor U9796 (N_9796,N_9205,N_9139);
and U9797 (N_9797,N_9497,N_9251);
nor U9798 (N_9798,N_9127,N_9186);
nor U9799 (N_9799,N_9399,N_9178);
and U9800 (N_9800,N_9351,N_9472);
xor U9801 (N_9801,N_9357,N_9367);
or U9802 (N_9802,N_9489,N_9276);
or U9803 (N_9803,N_9408,N_9263);
or U9804 (N_9804,N_9166,N_9249);
and U9805 (N_9805,N_9401,N_9209);
nor U9806 (N_9806,N_9056,N_9147);
or U9807 (N_9807,N_9217,N_9448);
xnor U9808 (N_9808,N_9275,N_9278);
nand U9809 (N_9809,N_9074,N_9108);
and U9810 (N_9810,N_9340,N_9446);
nor U9811 (N_9811,N_9233,N_9370);
or U9812 (N_9812,N_9291,N_9452);
nor U9813 (N_9813,N_9253,N_9305);
nand U9814 (N_9814,N_9480,N_9306);
or U9815 (N_9815,N_9462,N_9456);
xor U9816 (N_9816,N_9400,N_9412);
nor U9817 (N_9817,N_9426,N_9371);
or U9818 (N_9818,N_9448,N_9093);
or U9819 (N_9819,N_9085,N_9445);
nand U9820 (N_9820,N_9059,N_9365);
or U9821 (N_9821,N_9496,N_9358);
nand U9822 (N_9822,N_9250,N_9479);
or U9823 (N_9823,N_9049,N_9436);
nand U9824 (N_9824,N_9494,N_9010);
nand U9825 (N_9825,N_9322,N_9052);
or U9826 (N_9826,N_9495,N_9087);
and U9827 (N_9827,N_9160,N_9408);
and U9828 (N_9828,N_9165,N_9069);
nor U9829 (N_9829,N_9391,N_9314);
and U9830 (N_9830,N_9329,N_9257);
nor U9831 (N_9831,N_9250,N_9365);
and U9832 (N_9832,N_9091,N_9383);
or U9833 (N_9833,N_9062,N_9442);
xor U9834 (N_9834,N_9346,N_9391);
nand U9835 (N_9835,N_9173,N_9002);
nand U9836 (N_9836,N_9173,N_9107);
or U9837 (N_9837,N_9490,N_9262);
or U9838 (N_9838,N_9030,N_9074);
nand U9839 (N_9839,N_9446,N_9488);
or U9840 (N_9840,N_9091,N_9070);
and U9841 (N_9841,N_9078,N_9315);
or U9842 (N_9842,N_9341,N_9035);
nand U9843 (N_9843,N_9006,N_9283);
xnor U9844 (N_9844,N_9478,N_9147);
nand U9845 (N_9845,N_9330,N_9229);
and U9846 (N_9846,N_9073,N_9284);
and U9847 (N_9847,N_9466,N_9325);
and U9848 (N_9848,N_9061,N_9469);
or U9849 (N_9849,N_9184,N_9461);
nand U9850 (N_9850,N_9492,N_9306);
and U9851 (N_9851,N_9042,N_9370);
xor U9852 (N_9852,N_9172,N_9154);
nand U9853 (N_9853,N_9315,N_9021);
xor U9854 (N_9854,N_9304,N_9014);
nor U9855 (N_9855,N_9066,N_9227);
nor U9856 (N_9856,N_9022,N_9018);
nand U9857 (N_9857,N_9297,N_9166);
nor U9858 (N_9858,N_9374,N_9268);
nand U9859 (N_9859,N_9208,N_9309);
nand U9860 (N_9860,N_9364,N_9147);
xnor U9861 (N_9861,N_9227,N_9341);
nand U9862 (N_9862,N_9097,N_9260);
xnor U9863 (N_9863,N_9277,N_9238);
and U9864 (N_9864,N_9078,N_9292);
and U9865 (N_9865,N_9250,N_9335);
nor U9866 (N_9866,N_9472,N_9405);
nand U9867 (N_9867,N_9192,N_9067);
or U9868 (N_9868,N_9139,N_9468);
xor U9869 (N_9869,N_9132,N_9049);
and U9870 (N_9870,N_9487,N_9294);
and U9871 (N_9871,N_9397,N_9171);
nor U9872 (N_9872,N_9471,N_9283);
and U9873 (N_9873,N_9219,N_9154);
nor U9874 (N_9874,N_9214,N_9473);
nor U9875 (N_9875,N_9194,N_9036);
nand U9876 (N_9876,N_9313,N_9022);
nor U9877 (N_9877,N_9476,N_9438);
nand U9878 (N_9878,N_9067,N_9415);
xor U9879 (N_9879,N_9149,N_9237);
nand U9880 (N_9880,N_9216,N_9041);
or U9881 (N_9881,N_9120,N_9078);
or U9882 (N_9882,N_9127,N_9421);
nand U9883 (N_9883,N_9341,N_9288);
and U9884 (N_9884,N_9106,N_9144);
xnor U9885 (N_9885,N_9398,N_9450);
nand U9886 (N_9886,N_9464,N_9075);
xor U9887 (N_9887,N_9033,N_9113);
nand U9888 (N_9888,N_9082,N_9009);
or U9889 (N_9889,N_9444,N_9498);
nand U9890 (N_9890,N_9073,N_9169);
nand U9891 (N_9891,N_9159,N_9241);
and U9892 (N_9892,N_9100,N_9317);
nand U9893 (N_9893,N_9472,N_9399);
and U9894 (N_9894,N_9244,N_9003);
nand U9895 (N_9895,N_9322,N_9295);
xor U9896 (N_9896,N_9061,N_9483);
and U9897 (N_9897,N_9259,N_9179);
nand U9898 (N_9898,N_9171,N_9466);
or U9899 (N_9899,N_9055,N_9083);
xnor U9900 (N_9900,N_9013,N_9451);
or U9901 (N_9901,N_9472,N_9161);
xnor U9902 (N_9902,N_9249,N_9009);
nor U9903 (N_9903,N_9241,N_9157);
and U9904 (N_9904,N_9272,N_9377);
nor U9905 (N_9905,N_9241,N_9347);
nand U9906 (N_9906,N_9110,N_9471);
xnor U9907 (N_9907,N_9230,N_9132);
nor U9908 (N_9908,N_9371,N_9255);
and U9909 (N_9909,N_9139,N_9247);
xnor U9910 (N_9910,N_9368,N_9047);
nor U9911 (N_9911,N_9246,N_9007);
nand U9912 (N_9912,N_9082,N_9038);
or U9913 (N_9913,N_9215,N_9078);
nor U9914 (N_9914,N_9428,N_9381);
nand U9915 (N_9915,N_9187,N_9455);
and U9916 (N_9916,N_9443,N_9331);
and U9917 (N_9917,N_9363,N_9226);
nand U9918 (N_9918,N_9333,N_9368);
xor U9919 (N_9919,N_9016,N_9161);
nand U9920 (N_9920,N_9472,N_9033);
xor U9921 (N_9921,N_9222,N_9172);
and U9922 (N_9922,N_9487,N_9424);
or U9923 (N_9923,N_9165,N_9258);
and U9924 (N_9924,N_9041,N_9265);
nor U9925 (N_9925,N_9165,N_9137);
xor U9926 (N_9926,N_9116,N_9069);
nand U9927 (N_9927,N_9026,N_9191);
nor U9928 (N_9928,N_9431,N_9412);
xor U9929 (N_9929,N_9223,N_9173);
and U9930 (N_9930,N_9197,N_9160);
nand U9931 (N_9931,N_9486,N_9317);
nor U9932 (N_9932,N_9050,N_9363);
xor U9933 (N_9933,N_9061,N_9487);
nand U9934 (N_9934,N_9044,N_9250);
xor U9935 (N_9935,N_9449,N_9285);
and U9936 (N_9936,N_9226,N_9076);
or U9937 (N_9937,N_9321,N_9069);
or U9938 (N_9938,N_9285,N_9305);
nor U9939 (N_9939,N_9183,N_9362);
or U9940 (N_9940,N_9130,N_9444);
nand U9941 (N_9941,N_9123,N_9322);
or U9942 (N_9942,N_9259,N_9204);
and U9943 (N_9943,N_9042,N_9019);
xor U9944 (N_9944,N_9087,N_9000);
nor U9945 (N_9945,N_9194,N_9423);
or U9946 (N_9946,N_9101,N_9320);
nand U9947 (N_9947,N_9296,N_9497);
xnor U9948 (N_9948,N_9470,N_9225);
nand U9949 (N_9949,N_9383,N_9217);
or U9950 (N_9950,N_9296,N_9091);
nand U9951 (N_9951,N_9468,N_9452);
nor U9952 (N_9952,N_9320,N_9204);
nand U9953 (N_9953,N_9484,N_9035);
nor U9954 (N_9954,N_9049,N_9317);
or U9955 (N_9955,N_9244,N_9036);
nor U9956 (N_9956,N_9230,N_9385);
nor U9957 (N_9957,N_9479,N_9145);
or U9958 (N_9958,N_9133,N_9086);
nor U9959 (N_9959,N_9354,N_9478);
xor U9960 (N_9960,N_9143,N_9306);
nor U9961 (N_9961,N_9488,N_9023);
nand U9962 (N_9962,N_9252,N_9439);
xor U9963 (N_9963,N_9438,N_9472);
xor U9964 (N_9964,N_9065,N_9176);
and U9965 (N_9965,N_9014,N_9005);
nand U9966 (N_9966,N_9297,N_9223);
nor U9967 (N_9967,N_9259,N_9114);
xor U9968 (N_9968,N_9353,N_9412);
and U9969 (N_9969,N_9308,N_9324);
xnor U9970 (N_9970,N_9305,N_9489);
and U9971 (N_9971,N_9408,N_9299);
or U9972 (N_9972,N_9435,N_9284);
and U9973 (N_9973,N_9261,N_9188);
nor U9974 (N_9974,N_9026,N_9120);
or U9975 (N_9975,N_9312,N_9230);
nand U9976 (N_9976,N_9413,N_9316);
nand U9977 (N_9977,N_9262,N_9185);
and U9978 (N_9978,N_9253,N_9487);
and U9979 (N_9979,N_9317,N_9219);
and U9980 (N_9980,N_9048,N_9297);
and U9981 (N_9981,N_9102,N_9393);
xor U9982 (N_9982,N_9159,N_9421);
nand U9983 (N_9983,N_9024,N_9435);
nand U9984 (N_9984,N_9440,N_9483);
xnor U9985 (N_9985,N_9309,N_9257);
nand U9986 (N_9986,N_9455,N_9274);
nor U9987 (N_9987,N_9207,N_9435);
or U9988 (N_9988,N_9478,N_9450);
xor U9989 (N_9989,N_9150,N_9472);
nand U9990 (N_9990,N_9147,N_9079);
xnor U9991 (N_9991,N_9130,N_9047);
or U9992 (N_9992,N_9443,N_9356);
xnor U9993 (N_9993,N_9161,N_9255);
nand U9994 (N_9994,N_9205,N_9237);
and U9995 (N_9995,N_9048,N_9128);
or U9996 (N_9996,N_9096,N_9145);
xnor U9997 (N_9997,N_9184,N_9335);
or U9998 (N_9998,N_9436,N_9269);
and U9999 (N_9999,N_9352,N_9188);
or U10000 (N_10000,N_9851,N_9754);
or U10001 (N_10001,N_9900,N_9890);
and U10002 (N_10002,N_9865,N_9596);
nor U10003 (N_10003,N_9970,N_9808);
or U10004 (N_10004,N_9902,N_9811);
xor U10005 (N_10005,N_9614,N_9783);
and U10006 (N_10006,N_9738,N_9776);
and U10007 (N_10007,N_9508,N_9501);
nor U10008 (N_10008,N_9521,N_9678);
xnor U10009 (N_10009,N_9536,N_9701);
nand U10010 (N_10010,N_9854,N_9682);
xnor U10011 (N_10011,N_9798,N_9564);
or U10012 (N_10012,N_9696,N_9601);
xnor U10013 (N_10013,N_9895,N_9660);
nor U10014 (N_10014,N_9936,N_9722);
nor U10015 (N_10015,N_9563,N_9575);
and U10016 (N_10016,N_9918,N_9937);
xor U10017 (N_10017,N_9848,N_9887);
or U10018 (N_10018,N_9824,N_9770);
xnor U10019 (N_10019,N_9619,N_9781);
and U10020 (N_10020,N_9989,N_9675);
nor U10021 (N_10021,N_9917,N_9637);
xnor U10022 (N_10022,N_9843,N_9567);
nand U10023 (N_10023,N_9646,N_9868);
nor U10024 (N_10024,N_9967,N_9551);
or U10025 (N_10025,N_9741,N_9993);
xnor U10026 (N_10026,N_9623,N_9642);
xnor U10027 (N_10027,N_9802,N_9991);
and U10028 (N_10028,N_9743,N_9663);
xnor U10029 (N_10029,N_9951,N_9830);
or U10030 (N_10030,N_9872,N_9800);
nand U10031 (N_10031,N_9946,N_9842);
xor U10032 (N_10032,N_9505,N_9524);
nand U10033 (N_10033,N_9537,N_9915);
nor U10034 (N_10034,N_9995,N_9554);
nor U10035 (N_10035,N_9700,N_9891);
nand U10036 (N_10036,N_9503,N_9958);
and U10037 (N_10037,N_9913,N_9736);
and U10038 (N_10038,N_9599,N_9870);
or U10039 (N_10039,N_9606,N_9806);
and U10040 (N_10040,N_9829,N_9681);
nand U10041 (N_10041,N_9799,N_9899);
xor U10042 (N_10042,N_9698,N_9661);
and U10043 (N_10043,N_9990,N_9558);
and U10044 (N_10044,N_9643,N_9685);
nand U10045 (N_10045,N_9767,N_9828);
and U10046 (N_10046,N_9620,N_9846);
xor U10047 (N_10047,N_9844,N_9534);
and U10048 (N_10048,N_9571,N_9655);
xnor U10049 (N_10049,N_9791,N_9539);
nor U10050 (N_10050,N_9657,N_9764);
nand U10051 (N_10051,N_9883,N_9768);
or U10052 (N_10052,N_9717,N_9595);
xnor U10053 (N_10053,N_9628,N_9971);
nor U10054 (N_10054,N_9742,N_9904);
and U10055 (N_10055,N_9629,N_9603);
or U10056 (N_10056,N_9912,N_9880);
or U10057 (N_10057,N_9672,N_9873);
xor U10058 (N_10058,N_9548,N_9938);
and U10059 (N_10059,N_9812,N_9697);
or U10060 (N_10060,N_9962,N_9907);
nand U10061 (N_10061,N_9562,N_9861);
xor U10062 (N_10062,N_9513,N_9901);
nor U10063 (N_10063,N_9641,N_9914);
xnor U10064 (N_10064,N_9592,N_9976);
and U10065 (N_10065,N_9598,N_9588);
nor U10066 (N_10066,N_9707,N_9602);
xor U10067 (N_10067,N_9691,N_9975);
or U10068 (N_10068,N_9862,N_9765);
nor U10069 (N_10069,N_9699,N_9780);
nand U10070 (N_10070,N_9705,N_9615);
and U10071 (N_10071,N_9528,N_9980);
xor U10072 (N_10072,N_9627,N_9788);
nor U10073 (N_10073,N_9787,N_9674);
or U10074 (N_10074,N_9866,N_9879);
nor U10075 (N_10075,N_9519,N_9624);
and U10076 (N_10076,N_9896,N_9504);
and U10077 (N_10077,N_9587,N_9546);
nor U10078 (N_10078,N_9834,N_9527);
xnor U10079 (N_10079,N_9723,N_9857);
and U10080 (N_10080,N_9929,N_9875);
and U10081 (N_10081,N_9827,N_9676);
nor U10082 (N_10082,N_9612,N_9784);
xnor U10083 (N_10083,N_9977,N_9838);
xnor U10084 (N_10084,N_9740,N_9797);
nor U10085 (N_10085,N_9773,N_9935);
nand U10086 (N_10086,N_9626,N_9925);
or U10087 (N_10087,N_9998,N_9909);
or U10088 (N_10088,N_9777,N_9545);
nor U10089 (N_10089,N_9718,N_9953);
xor U10090 (N_10090,N_9745,N_9502);
or U10091 (N_10091,N_9910,N_9968);
nor U10092 (N_10092,N_9613,N_9943);
or U10093 (N_10093,N_9583,N_9923);
or U10094 (N_10094,N_9758,N_9724);
and U10095 (N_10095,N_9955,N_9852);
xor U10096 (N_10096,N_9749,N_9530);
nor U10097 (N_10097,N_9826,N_9529);
xnor U10098 (N_10098,N_9730,N_9704);
and U10099 (N_10099,N_9631,N_9541);
nor U10100 (N_10100,N_9618,N_9919);
and U10101 (N_10101,N_9856,N_9982);
and U10102 (N_10102,N_9898,N_9974);
nand U10103 (N_10103,N_9589,N_9559);
and U10104 (N_10104,N_9570,N_9978);
and U10105 (N_10105,N_9930,N_9855);
nor U10106 (N_10106,N_9669,N_9825);
nand U10107 (N_10107,N_9579,N_9638);
nand U10108 (N_10108,N_9771,N_9600);
xor U10109 (N_10109,N_9966,N_9533);
nor U10110 (N_10110,N_9805,N_9684);
xor U10111 (N_10111,N_9874,N_9858);
nand U10112 (N_10112,N_9963,N_9869);
xor U10113 (N_10113,N_9511,N_9610);
nand U10114 (N_10114,N_9934,N_9702);
nand U10115 (N_10115,N_9514,N_9756);
xnor U10116 (N_10116,N_9926,N_9867);
and U10117 (N_10117,N_9817,N_9737);
and U10118 (N_10118,N_9731,N_9590);
and U10119 (N_10119,N_9645,N_9574);
nand U10120 (N_10120,N_9594,N_9709);
xnor U10121 (N_10121,N_9630,N_9656);
or U10122 (N_10122,N_9959,N_9840);
nand U10123 (N_10123,N_9782,N_9597);
nor U10124 (N_10124,N_9755,N_9762);
and U10125 (N_10125,N_9747,N_9665);
nand U10126 (N_10126,N_9894,N_9803);
and U10127 (N_10127,N_9761,N_9994);
xnor U10128 (N_10128,N_9997,N_9651);
nor U10129 (N_10129,N_9703,N_9807);
xnor U10130 (N_10130,N_9653,N_9833);
nand U10131 (N_10131,N_9985,N_9821);
nor U10132 (N_10132,N_9734,N_9969);
or U10133 (N_10133,N_9549,N_9778);
and U10134 (N_10134,N_9832,N_9987);
nor U10135 (N_10135,N_9779,N_9635);
nor U10136 (N_10136,N_9711,N_9555);
xor U10137 (N_10137,N_9720,N_9786);
and U10138 (N_10138,N_9956,N_9560);
xor U10139 (N_10139,N_9582,N_9877);
and U10140 (N_10140,N_9690,N_9526);
nor U10141 (N_10141,N_9772,N_9584);
nor U10142 (N_10142,N_9729,N_9726);
and U10143 (N_10143,N_9948,N_9591);
nor U10144 (N_10144,N_9577,N_9608);
and U10145 (N_10145,N_9813,N_9816);
and U10146 (N_10146,N_9659,N_9552);
xor U10147 (N_10147,N_9622,N_9979);
xnor U10148 (N_10148,N_9728,N_9666);
nor U10149 (N_10149,N_9725,N_9905);
and U10150 (N_10150,N_9658,N_9760);
xor U10151 (N_10151,N_9878,N_9580);
or U10152 (N_10152,N_9820,N_9632);
xnor U10153 (N_10153,N_9836,N_9538);
nand U10154 (N_10154,N_9794,N_9540);
and U10155 (N_10155,N_9522,N_9517);
nor U10156 (N_10156,N_9815,N_9680);
or U10157 (N_10157,N_9954,N_9999);
nand U10158 (N_10158,N_9604,N_9565);
nand U10159 (N_10159,N_9947,N_9992);
nand U10160 (N_10160,N_9897,N_9739);
or U10161 (N_10161,N_9908,N_9735);
nor U10162 (N_10162,N_9692,N_9727);
or U10163 (N_10163,N_9689,N_9984);
xor U10164 (N_10164,N_9532,N_9906);
nor U10165 (N_10165,N_9759,N_9810);
and U10166 (N_10166,N_9550,N_9662);
nand U10167 (N_10167,N_9924,N_9860);
nor U10168 (N_10168,N_9616,N_9694);
and U10169 (N_10169,N_9965,N_9876);
and U10170 (N_10170,N_9667,N_9647);
or U10171 (N_10171,N_9634,N_9586);
or U10172 (N_10172,N_9751,N_9795);
or U10173 (N_10173,N_9774,N_9520);
and U10174 (N_10174,N_9839,N_9719);
nor U10175 (N_10175,N_9940,N_9687);
and U10176 (N_10176,N_9957,N_9686);
xnor U10177 (N_10177,N_9920,N_9819);
and U10178 (N_10178,N_9964,N_9516);
and U10179 (N_10179,N_9581,N_9983);
xnor U10180 (N_10180,N_9605,N_9973);
nor U10181 (N_10181,N_9790,N_9853);
or U10182 (N_10182,N_9556,N_9886);
nand U10183 (N_10183,N_9921,N_9708);
and U10184 (N_10184,N_9892,N_9847);
and U10185 (N_10185,N_9649,N_9945);
and U10186 (N_10186,N_9793,N_9688);
xor U10187 (N_10187,N_9933,N_9944);
nand U10188 (N_10188,N_9916,N_9668);
xor U10189 (N_10189,N_9617,N_9673);
nor U10190 (N_10190,N_9535,N_9510);
nor U10191 (N_10191,N_9952,N_9542);
nor U10192 (N_10192,N_9523,N_9850);
or U10193 (N_10193,N_9931,N_9713);
and U10194 (N_10194,N_9515,N_9512);
nor U10195 (N_10195,N_9573,N_9835);
and U10196 (N_10196,N_9644,N_9561);
or U10197 (N_10197,N_9972,N_9531);
nor U10198 (N_10198,N_9706,N_9721);
or U10199 (N_10199,N_9746,N_9569);
nor U10200 (N_10200,N_9670,N_9607);
and U10201 (N_10201,N_9789,N_9942);
xor U10202 (N_10202,N_9809,N_9593);
xor U10203 (N_10203,N_9544,N_9949);
xnor U10204 (N_10204,N_9748,N_9712);
nor U10205 (N_10205,N_9792,N_9625);
nand U10206 (N_10206,N_9814,N_9566);
nand U10207 (N_10207,N_9652,N_9859);
nand U10208 (N_10208,N_9543,N_9671);
and U10209 (N_10209,N_9547,N_9888);
or U10210 (N_10210,N_9884,N_9961);
xnor U10211 (N_10211,N_9796,N_9903);
or U10212 (N_10212,N_9716,N_9831);
and U10213 (N_10213,N_9664,N_9753);
or U10214 (N_10214,N_9823,N_9766);
xnor U10215 (N_10215,N_9763,N_9525);
or U10216 (N_10216,N_9845,N_9801);
xor U10217 (N_10217,N_9732,N_9769);
nand U10218 (N_10218,N_9871,N_9863);
and U10219 (N_10219,N_9633,N_9988);
xnor U10220 (N_10220,N_9960,N_9733);
xnor U10221 (N_10221,N_9928,N_9553);
nor U10222 (N_10222,N_9500,N_9981);
xor U10223 (N_10223,N_9609,N_9578);
and U10224 (N_10224,N_9677,N_9996);
nand U10225 (N_10225,N_9911,N_9585);
or U10226 (N_10226,N_9557,N_9882);
and U10227 (N_10227,N_9893,N_9648);
nor U10228 (N_10228,N_9695,N_9693);
and U10229 (N_10229,N_9679,N_9804);
or U10230 (N_10230,N_9654,N_9785);
nor U10231 (N_10231,N_9941,N_9822);
and U10232 (N_10232,N_9752,N_9714);
or U10233 (N_10233,N_9986,N_9841);
and U10234 (N_10234,N_9927,N_9775);
and U10235 (N_10235,N_9922,N_9506);
nor U10236 (N_10236,N_9837,N_9576);
xnor U10237 (N_10237,N_9849,N_9710);
and U10238 (N_10238,N_9939,N_9611);
xor U10239 (N_10239,N_9572,N_9881);
and U10240 (N_10240,N_9744,N_9621);
or U10241 (N_10241,N_9650,N_9568);
and U10242 (N_10242,N_9885,N_9889);
and U10243 (N_10243,N_9640,N_9683);
nand U10244 (N_10244,N_9864,N_9950);
and U10245 (N_10245,N_9507,N_9932);
and U10246 (N_10246,N_9509,N_9757);
or U10247 (N_10247,N_9715,N_9639);
and U10248 (N_10248,N_9750,N_9518);
or U10249 (N_10249,N_9636,N_9818);
nand U10250 (N_10250,N_9768,N_9669);
nor U10251 (N_10251,N_9587,N_9588);
or U10252 (N_10252,N_9561,N_9558);
nand U10253 (N_10253,N_9983,N_9562);
nand U10254 (N_10254,N_9971,N_9725);
and U10255 (N_10255,N_9981,N_9573);
nand U10256 (N_10256,N_9757,N_9700);
or U10257 (N_10257,N_9810,N_9788);
nand U10258 (N_10258,N_9671,N_9988);
nand U10259 (N_10259,N_9850,N_9973);
or U10260 (N_10260,N_9641,N_9863);
or U10261 (N_10261,N_9852,N_9926);
nor U10262 (N_10262,N_9834,N_9724);
and U10263 (N_10263,N_9784,N_9789);
xnor U10264 (N_10264,N_9963,N_9605);
xor U10265 (N_10265,N_9736,N_9506);
xor U10266 (N_10266,N_9667,N_9824);
xor U10267 (N_10267,N_9798,N_9932);
xor U10268 (N_10268,N_9820,N_9633);
nand U10269 (N_10269,N_9734,N_9708);
xor U10270 (N_10270,N_9784,N_9874);
xnor U10271 (N_10271,N_9547,N_9568);
xor U10272 (N_10272,N_9875,N_9980);
and U10273 (N_10273,N_9680,N_9806);
and U10274 (N_10274,N_9781,N_9758);
nand U10275 (N_10275,N_9516,N_9904);
xor U10276 (N_10276,N_9574,N_9812);
xor U10277 (N_10277,N_9587,N_9686);
nand U10278 (N_10278,N_9907,N_9707);
nand U10279 (N_10279,N_9663,N_9856);
xor U10280 (N_10280,N_9534,N_9767);
nand U10281 (N_10281,N_9882,N_9784);
nand U10282 (N_10282,N_9875,N_9740);
xnor U10283 (N_10283,N_9542,N_9662);
xnor U10284 (N_10284,N_9810,N_9990);
or U10285 (N_10285,N_9794,N_9586);
or U10286 (N_10286,N_9987,N_9877);
or U10287 (N_10287,N_9957,N_9743);
nand U10288 (N_10288,N_9749,N_9692);
nor U10289 (N_10289,N_9863,N_9570);
or U10290 (N_10290,N_9659,N_9501);
nand U10291 (N_10291,N_9563,N_9691);
nand U10292 (N_10292,N_9679,N_9891);
nand U10293 (N_10293,N_9893,N_9754);
nand U10294 (N_10294,N_9542,N_9533);
and U10295 (N_10295,N_9583,N_9777);
nor U10296 (N_10296,N_9656,N_9944);
nor U10297 (N_10297,N_9841,N_9546);
nor U10298 (N_10298,N_9961,N_9720);
nand U10299 (N_10299,N_9572,N_9836);
or U10300 (N_10300,N_9524,N_9725);
and U10301 (N_10301,N_9982,N_9924);
xor U10302 (N_10302,N_9673,N_9871);
and U10303 (N_10303,N_9682,N_9811);
nor U10304 (N_10304,N_9613,N_9823);
and U10305 (N_10305,N_9779,N_9552);
and U10306 (N_10306,N_9824,N_9814);
nor U10307 (N_10307,N_9532,N_9637);
and U10308 (N_10308,N_9594,N_9615);
or U10309 (N_10309,N_9982,N_9998);
nand U10310 (N_10310,N_9752,N_9732);
nand U10311 (N_10311,N_9626,N_9901);
xnor U10312 (N_10312,N_9862,N_9507);
and U10313 (N_10313,N_9828,N_9953);
nor U10314 (N_10314,N_9681,N_9617);
nand U10315 (N_10315,N_9695,N_9883);
and U10316 (N_10316,N_9807,N_9687);
or U10317 (N_10317,N_9523,N_9859);
xnor U10318 (N_10318,N_9635,N_9758);
nor U10319 (N_10319,N_9525,N_9577);
nand U10320 (N_10320,N_9899,N_9517);
nand U10321 (N_10321,N_9709,N_9970);
xnor U10322 (N_10322,N_9516,N_9707);
nand U10323 (N_10323,N_9840,N_9654);
nor U10324 (N_10324,N_9932,N_9578);
or U10325 (N_10325,N_9575,N_9656);
xnor U10326 (N_10326,N_9551,N_9973);
nand U10327 (N_10327,N_9758,N_9707);
nor U10328 (N_10328,N_9585,N_9678);
or U10329 (N_10329,N_9870,N_9937);
nand U10330 (N_10330,N_9996,N_9779);
xnor U10331 (N_10331,N_9980,N_9970);
or U10332 (N_10332,N_9891,N_9641);
nand U10333 (N_10333,N_9759,N_9899);
xnor U10334 (N_10334,N_9978,N_9758);
xnor U10335 (N_10335,N_9744,N_9916);
and U10336 (N_10336,N_9957,N_9824);
or U10337 (N_10337,N_9865,N_9703);
nor U10338 (N_10338,N_9956,N_9965);
or U10339 (N_10339,N_9931,N_9880);
or U10340 (N_10340,N_9855,N_9958);
xor U10341 (N_10341,N_9897,N_9798);
nor U10342 (N_10342,N_9705,N_9675);
nor U10343 (N_10343,N_9723,N_9876);
nor U10344 (N_10344,N_9924,N_9629);
xor U10345 (N_10345,N_9799,N_9824);
xor U10346 (N_10346,N_9910,N_9926);
and U10347 (N_10347,N_9755,N_9545);
nor U10348 (N_10348,N_9915,N_9745);
xnor U10349 (N_10349,N_9620,N_9859);
xnor U10350 (N_10350,N_9848,N_9817);
or U10351 (N_10351,N_9539,N_9832);
nor U10352 (N_10352,N_9567,N_9629);
or U10353 (N_10353,N_9707,N_9971);
or U10354 (N_10354,N_9665,N_9943);
and U10355 (N_10355,N_9530,N_9995);
nor U10356 (N_10356,N_9646,N_9677);
or U10357 (N_10357,N_9862,N_9506);
and U10358 (N_10358,N_9783,N_9760);
nor U10359 (N_10359,N_9838,N_9687);
xnor U10360 (N_10360,N_9900,N_9979);
xor U10361 (N_10361,N_9644,N_9759);
nor U10362 (N_10362,N_9763,N_9658);
and U10363 (N_10363,N_9845,N_9627);
nand U10364 (N_10364,N_9779,N_9521);
and U10365 (N_10365,N_9683,N_9704);
and U10366 (N_10366,N_9958,N_9649);
xor U10367 (N_10367,N_9541,N_9872);
xnor U10368 (N_10368,N_9613,N_9798);
nand U10369 (N_10369,N_9661,N_9824);
nor U10370 (N_10370,N_9684,N_9607);
xnor U10371 (N_10371,N_9866,N_9820);
nor U10372 (N_10372,N_9795,N_9765);
nand U10373 (N_10373,N_9948,N_9934);
or U10374 (N_10374,N_9634,N_9809);
nand U10375 (N_10375,N_9950,N_9936);
and U10376 (N_10376,N_9824,N_9716);
or U10377 (N_10377,N_9631,N_9969);
xor U10378 (N_10378,N_9620,N_9614);
xnor U10379 (N_10379,N_9953,N_9997);
nor U10380 (N_10380,N_9526,N_9873);
xnor U10381 (N_10381,N_9689,N_9740);
xor U10382 (N_10382,N_9945,N_9814);
and U10383 (N_10383,N_9596,N_9752);
xnor U10384 (N_10384,N_9604,N_9929);
and U10385 (N_10385,N_9638,N_9507);
nand U10386 (N_10386,N_9904,N_9721);
nand U10387 (N_10387,N_9533,N_9617);
nand U10388 (N_10388,N_9776,N_9700);
xor U10389 (N_10389,N_9783,N_9841);
nand U10390 (N_10390,N_9826,N_9733);
nand U10391 (N_10391,N_9966,N_9702);
or U10392 (N_10392,N_9740,N_9910);
nand U10393 (N_10393,N_9979,N_9827);
nand U10394 (N_10394,N_9752,N_9906);
xor U10395 (N_10395,N_9831,N_9907);
nor U10396 (N_10396,N_9711,N_9659);
or U10397 (N_10397,N_9624,N_9856);
or U10398 (N_10398,N_9707,N_9691);
or U10399 (N_10399,N_9578,N_9846);
and U10400 (N_10400,N_9594,N_9720);
or U10401 (N_10401,N_9953,N_9689);
nand U10402 (N_10402,N_9533,N_9877);
or U10403 (N_10403,N_9652,N_9606);
and U10404 (N_10404,N_9960,N_9976);
nor U10405 (N_10405,N_9670,N_9698);
nor U10406 (N_10406,N_9860,N_9748);
xor U10407 (N_10407,N_9697,N_9827);
xnor U10408 (N_10408,N_9596,N_9595);
nand U10409 (N_10409,N_9932,N_9664);
xnor U10410 (N_10410,N_9938,N_9997);
xnor U10411 (N_10411,N_9572,N_9636);
nand U10412 (N_10412,N_9678,N_9786);
and U10413 (N_10413,N_9666,N_9882);
nand U10414 (N_10414,N_9878,N_9882);
xor U10415 (N_10415,N_9659,N_9647);
nor U10416 (N_10416,N_9520,N_9530);
xnor U10417 (N_10417,N_9991,N_9625);
xor U10418 (N_10418,N_9598,N_9825);
xnor U10419 (N_10419,N_9633,N_9830);
nand U10420 (N_10420,N_9859,N_9894);
nor U10421 (N_10421,N_9504,N_9529);
and U10422 (N_10422,N_9883,N_9978);
xor U10423 (N_10423,N_9736,N_9842);
and U10424 (N_10424,N_9530,N_9973);
nor U10425 (N_10425,N_9667,N_9658);
and U10426 (N_10426,N_9860,N_9704);
nand U10427 (N_10427,N_9948,N_9518);
xor U10428 (N_10428,N_9846,N_9684);
nor U10429 (N_10429,N_9565,N_9533);
nor U10430 (N_10430,N_9867,N_9762);
xor U10431 (N_10431,N_9812,N_9997);
nand U10432 (N_10432,N_9545,N_9848);
or U10433 (N_10433,N_9625,N_9872);
or U10434 (N_10434,N_9823,N_9535);
nand U10435 (N_10435,N_9552,N_9928);
nand U10436 (N_10436,N_9947,N_9554);
nand U10437 (N_10437,N_9606,N_9706);
xnor U10438 (N_10438,N_9837,N_9764);
xnor U10439 (N_10439,N_9743,N_9846);
and U10440 (N_10440,N_9665,N_9772);
nor U10441 (N_10441,N_9983,N_9596);
xnor U10442 (N_10442,N_9610,N_9935);
xor U10443 (N_10443,N_9525,N_9519);
nor U10444 (N_10444,N_9883,N_9832);
or U10445 (N_10445,N_9645,N_9736);
and U10446 (N_10446,N_9991,N_9586);
xor U10447 (N_10447,N_9840,N_9507);
and U10448 (N_10448,N_9609,N_9611);
nand U10449 (N_10449,N_9660,N_9970);
nand U10450 (N_10450,N_9614,N_9885);
or U10451 (N_10451,N_9871,N_9502);
and U10452 (N_10452,N_9656,N_9728);
or U10453 (N_10453,N_9573,N_9779);
xnor U10454 (N_10454,N_9617,N_9530);
or U10455 (N_10455,N_9911,N_9929);
nand U10456 (N_10456,N_9982,N_9532);
nand U10457 (N_10457,N_9541,N_9875);
or U10458 (N_10458,N_9749,N_9562);
and U10459 (N_10459,N_9733,N_9749);
or U10460 (N_10460,N_9715,N_9904);
nor U10461 (N_10461,N_9682,N_9657);
nor U10462 (N_10462,N_9516,N_9543);
nand U10463 (N_10463,N_9840,N_9752);
or U10464 (N_10464,N_9995,N_9536);
nor U10465 (N_10465,N_9946,N_9980);
and U10466 (N_10466,N_9704,N_9824);
or U10467 (N_10467,N_9917,N_9923);
or U10468 (N_10468,N_9940,N_9997);
and U10469 (N_10469,N_9877,N_9775);
nand U10470 (N_10470,N_9767,N_9991);
and U10471 (N_10471,N_9713,N_9710);
and U10472 (N_10472,N_9844,N_9695);
nand U10473 (N_10473,N_9561,N_9833);
nor U10474 (N_10474,N_9637,N_9640);
or U10475 (N_10475,N_9545,N_9634);
and U10476 (N_10476,N_9511,N_9661);
xor U10477 (N_10477,N_9806,N_9964);
or U10478 (N_10478,N_9600,N_9548);
and U10479 (N_10479,N_9849,N_9940);
nand U10480 (N_10480,N_9544,N_9616);
and U10481 (N_10481,N_9759,N_9675);
nor U10482 (N_10482,N_9805,N_9519);
or U10483 (N_10483,N_9854,N_9793);
nor U10484 (N_10484,N_9751,N_9949);
or U10485 (N_10485,N_9996,N_9801);
xor U10486 (N_10486,N_9822,N_9532);
xor U10487 (N_10487,N_9743,N_9540);
and U10488 (N_10488,N_9601,N_9670);
nand U10489 (N_10489,N_9753,N_9957);
or U10490 (N_10490,N_9548,N_9603);
xor U10491 (N_10491,N_9802,N_9703);
xor U10492 (N_10492,N_9936,N_9528);
and U10493 (N_10493,N_9748,N_9793);
nand U10494 (N_10494,N_9977,N_9704);
nand U10495 (N_10495,N_9740,N_9820);
or U10496 (N_10496,N_9847,N_9551);
and U10497 (N_10497,N_9913,N_9800);
or U10498 (N_10498,N_9792,N_9789);
and U10499 (N_10499,N_9794,N_9869);
nor U10500 (N_10500,N_10310,N_10302);
nand U10501 (N_10501,N_10049,N_10379);
and U10502 (N_10502,N_10220,N_10184);
nand U10503 (N_10503,N_10145,N_10135);
xor U10504 (N_10504,N_10185,N_10139);
and U10505 (N_10505,N_10419,N_10098);
xor U10506 (N_10506,N_10240,N_10385);
xnor U10507 (N_10507,N_10369,N_10437);
or U10508 (N_10508,N_10000,N_10335);
xnor U10509 (N_10509,N_10111,N_10477);
xor U10510 (N_10510,N_10440,N_10328);
nand U10511 (N_10511,N_10412,N_10390);
or U10512 (N_10512,N_10435,N_10360);
and U10513 (N_10513,N_10093,N_10094);
nand U10514 (N_10514,N_10048,N_10023);
and U10515 (N_10515,N_10449,N_10339);
or U10516 (N_10516,N_10167,N_10337);
or U10517 (N_10517,N_10485,N_10469);
or U10518 (N_10518,N_10002,N_10027);
or U10519 (N_10519,N_10192,N_10365);
nor U10520 (N_10520,N_10248,N_10333);
and U10521 (N_10521,N_10095,N_10007);
xor U10522 (N_10522,N_10151,N_10253);
xnor U10523 (N_10523,N_10482,N_10439);
nand U10524 (N_10524,N_10186,N_10112);
nand U10525 (N_10525,N_10164,N_10232);
nor U10526 (N_10526,N_10236,N_10173);
nand U10527 (N_10527,N_10085,N_10043);
nand U10528 (N_10528,N_10036,N_10193);
nand U10529 (N_10529,N_10046,N_10309);
nand U10530 (N_10530,N_10357,N_10096);
and U10531 (N_10531,N_10190,N_10075);
nor U10532 (N_10532,N_10138,N_10426);
and U10533 (N_10533,N_10380,N_10057);
or U10534 (N_10534,N_10037,N_10320);
and U10535 (N_10535,N_10129,N_10176);
or U10536 (N_10536,N_10022,N_10345);
and U10537 (N_10537,N_10104,N_10494);
or U10538 (N_10538,N_10457,N_10197);
nand U10539 (N_10539,N_10080,N_10131);
or U10540 (N_10540,N_10355,N_10463);
nand U10541 (N_10541,N_10406,N_10019);
nand U10542 (N_10542,N_10327,N_10281);
nand U10543 (N_10543,N_10126,N_10142);
or U10544 (N_10544,N_10246,N_10227);
and U10545 (N_10545,N_10404,N_10398);
or U10546 (N_10546,N_10191,N_10231);
or U10547 (N_10547,N_10493,N_10341);
and U10548 (N_10548,N_10330,N_10351);
and U10549 (N_10549,N_10265,N_10148);
xor U10550 (N_10550,N_10307,N_10225);
and U10551 (N_10551,N_10376,N_10051);
and U10552 (N_10552,N_10206,N_10137);
nor U10553 (N_10553,N_10492,N_10081);
nand U10554 (N_10554,N_10389,N_10498);
or U10555 (N_10555,N_10155,N_10268);
and U10556 (N_10556,N_10004,N_10461);
nor U10557 (N_10557,N_10045,N_10450);
xnor U10558 (N_10558,N_10067,N_10063);
and U10559 (N_10559,N_10420,N_10241);
nor U10560 (N_10560,N_10103,N_10047);
and U10561 (N_10561,N_10034,N_10024);
or U10562 (N_10562,N_10316,N_10226);
nand U10563 (N_10563,N_10203,N_10286);
or U10564 (N_10564,N_10405,N_10251);
nand U10565 (N_10565,N_10417,N_10099);
xor U10566 (N_10566,N_10234,N_10446);
and U10567 (N_10567,N_10260,N_10179);
and U10568 (N_10568,N_10041,N_10213);
and U10569 (N_10569,N_10064,N_10323);
nor U10570 (N_10570,N_10490,N_10211);
xnor U10571 (N_10571,N_10212,N_10074);
nor U10572 (N_10572,N_10101,N_10486);
nor U10573 (N_10573,N_10267,N_10395);
and U10574 (N_10574,N_10278,N_10006);
nor U10575 (N_10575,N_10361,N_10218);
xnor U10576 (N_10576,N_10242,N_10352);
xnor U10577 (N_10577,N_10090,N_10257);
nor U10578 (N_10578,N_10154,N_10035);
nor U10579 (N_10579,N_10358,N_10243);
nand U10580 (N_10580,N_10445,N_10172);
and U10581 (N_10581,N_10038,N_10296);
nand U10582 (N_10582,N_10366,N_10367);
nor U10583 (N_10583,N_10165,N_10315);
and U10584 (N_10584,N_10195,N_10336);
and U10585 (N_10585,N_10318,N_10247);
and U10586 (N_10586,N_10429,N_10387);
or U10587 (N_10587,N_10427,N_10059);
or U10588 (N_10588,N_10263,N_10269);
nor U10589 (N_10589,N_10329,N_10201);
xnor U10590 (N_10590,N_10487,N_10144);
nand U10591 (N_10591,N_10146,N_10354);
nand U10592 (N_10592,N_10187,N_10065);
and U10593 (N_10593,N_10421,N_10411);
and U10594 (N_10594,N_10194,N_10216);
and U10595 (N_10595,N_10181,N_10244);
and U10596 (N_10596,N_10384,N_10326);
nor U10597 (N_10597,N_10344,N_10386);
nand U10598 (N_10598,N_10465,N_10061);
nand U10599 (N_10599,N_10013,N_10130);
and U10600 (N_10600,N_10219,N_10478);
and U10601 (N_10601,N_10128,N_10350);
and U10602 (N_10602,N_10393,N_10270);
nor U10603 (N_10603,N_10343,N_10015);
and U10604 (N_10604,N_10282,N_10430);
xnor U10605 (N_10605,N_10056,N_10223);
xnor U10606 (N_10606,N_10118,N_10293);
nor U10607 (N_10607,N_10418,N_10136);
and U10608 (N_10608,N_10356,N_10169);
xor U10609 (N_10609,N_10324,N_10495);
nor U10610 (N_10610,N_10455,N_10143);
and U10611 (N_10611,N_10070,N_10434);
and U10612 (N_10612,N_10189,N_10346);
nand U10613 (N_10613,N_10025,N_10105);
or U10614 (N_10614,N_10082,N_10140);
or U10615 (N_10615,N_10483,N_10353);
xnor U10616 (N_10616,N_10292,N_10416);
nand U10617 (N_10617,N_10259,N_10030);
xnor U10618 (N_10618,N_10071,N_10397);
xnor U10619 (N_10619,N_10062,N_10170);
nand U10620 (N_10620,N_10338,N_10459);
and U10621 (N_10621,N_10392,N_10238);
or U10622 (N_10622,N_10077,N_10290);
and U10623 (N_10623,N_10467,N_10011);
or U10624 (N_10624,N_10252,N_10003);
nand U10625 (N_10625,N_10381,N_10403);
xor U10626 (N_10626,N_10488,N_10442);
nand U10627 (N_10627,N_10413,N_10147);
and U10628 (N_10628,N_10141,N_10497);
nor U10629 (N_10629,N_10311,N_10221);
or U10630 (N_10630,N_10300,N_10150);
nor U10631 (N_10631,N_10363,N_10414);
or U10632 (N_10632,N_10444,N_10266);
or U10633 (N_10633,N_10297,N_10097);
or U10634 (N_10634,N_10438,N_10382);
nor U10635 (N_10635,N_10110,N_10399);
xor U10636 (N_10636,N_10271,N_10291);
or U10637 (N_10637,N_10092,N_10298);
nor U10638 (N_10638,N_10076,N_10375);
and U10639 (N_10639,N_10275,N_10202);
and U10640 (N_10640,N_10084,N_10204);
and U10641 (N_10641,N_10016,N_10012);
xnor U10642 (N_10642,N_10134,N_10331);
nand U10643 (N_10643,N_10072,N_10162);
xor U10644 (N_10644,N_10371,N_10304);
or U10645 (N_10645,N_10156,N_10254);
xnor U10646 (N_10646,N_10055,N_10370);
xnor U10647 (N_10647,N_10250,N_10317);
or U10648 (N_10648,N_10456,N_10471);
xnor U10649 (N_10649,N_10157,N_10009);
nand U10650 (N_10650,N_10332,N_10088);
or U10651 (N_10651,N_10039,N_10479);
and U10652 (N_10652,N_10453,N_10233);
or U10653 (N_10653,N_10454,N_10228);
xnor U10654 (N_10654,N_10272,N_10410);
or U10655 (N_10655,N_10264,N_10305);
or U10656 (N_10656,N_10078,N_10441);
xnor U10657 (N_10657,N_10239,N_10102);
or U10658 (N_10658,N_10209,N_10308);
or U10659 (N_10659,N_10159,N_10001);
and U10660 (N_10660,N_10447,N_10086);
xnor U10661 (N_10661,N_10347,N_10010);
nand U10662 (N_10662,N_10113,N_10031);
nor U10663 (N_10663,N_10364,N_10277);
nand U10664 (N_10664,N_10106,N_10091);
nor U10665 (N_10665,N_10208,N_10119);
or U10666 (N_10666,N_10472,N_10499);
nor U10667 (N_10667,N_10443,N_10287);
nor U10668 (N_10668,N_10100,N_10127);
nand U10669 (N_10669,N_10188,N_10132);
nor U10670 (N_10670,N_10174,N_10273);
nor U10671 (N_10671,N_10029,N_10042);
nor U10672 (N_10672,N_10462,N_10026);
xnor U10673 (N_10673,N_10117,N_10033);
or U10674 (N_10674,N_10237,N_10249);
nor U10675 (N_10675,N_10149,N_10284);
or U10676 (N_10676,N_10295,N_10050);
or U10677 (N_10677,N_10448,N_10205);
and U10678 (N_10678,N_10044,N_10217);
xor U10679 (N_10679,N_10152,N_10391);
nand U10680 (N_10680,N_10073,N_10303);
xnor U10681 (N_10681,N_10359,N_10422);
nor U10682 (N_10682,N_10415,N_10222);
xnor U10683 (N_10683,N_10121,N_10198);
nor U10684 (N_10684,N_10400,N_10423);
nor U10685 (N_10685,N_10255,N_10052);
nand U10686 (N_10686,N_10163,N_10294);
and U10687 (N_10687,N_10373,N_10068);
xor U10688 (N_10688,N_10464,N_10374);
or U10689 (N_10689,N_10409,N_10183);
xnor U10690 (N_10690,N_10109,N_10325);
and U10691 (N_10691,N_10388,N_10340);
xor U10692 (N_10692,N_10377,N_10285);
nand U10693 (N_10693,N_10476,N_10491);
nor U10694 (N_10694,N_10408,N_10362);
or U10695 (N_10695,N_10180,N_10177);
xor U10696 (N_10696,N_10394,N_10460);
and U10697 (N_10697,N_10224,N_10288);
and U10698 (N_10698,N_10262,N_10060);
or U10699 (N_10699,N_10175,N_10171);
xor U10700 (N_10700,N_10452,N_10474);
xor U10701 (N_10701,N_10207,N_10306);
nand U10702 (N_10702,N_10158,N_10018);
or U10703 (N_10703,N_10032,N_10160);
nand U10704 (N_10704,N_10276,N_10066);
nor U10705 (N_10705,N_10424,N_10199);
nor U10706 (N_10706,N_10168,N_10178);
or U10707 (N_10707,N_10040,N_10312);
and U10708 (N_10708,N_10182,N_10484);
xor U10709 (N_10709,N_10480,N_10079);
or U10710 (N_10710,N_10210,N_10431);
nor U10711 (N_10711,N_10299,N_10349);
and U10712 (N_10712,N_10342,N_10314);
nand U10713 (N_10713,N_10017,N_10235);
nor U10714 (N_10714,N_10468,N_10083);
and U10715 (N_10715,N_10115,N_10058);
or U10716 (N_10716,N_10114,N_10458);
nand U10717 (N_10717,N_10425,N_10005);
and U10718 (N_10718,N_10215,N_10166);
and U10719 (N_10719,N_10321,N_10283);
nand U10720 (N_10720,N_10028,N_10496);
nor U10721 (N_10721,N_10125,N_10289);
nor U10722 (N_10722,N_10214,N_10279);
nor U10723 (N_10723,N_10313,N_10451);
xor U10724 (N_10724,N_10473,N_10108);
nor U10725 (N_10725,N_10402,N_10466);
and U10726 (N_10726,N_10122,N_10020);
and U10727 (N_10727,N_10319,N_10200);
nand U10728 (N_10728,N_10433,N_10383);
or U10729 (N_10729,N_10008,N_10123);
xnor U10730 (N_10730,N_10322,N_10069);
or U10731 (N_10731,N_10280,N_10470);
and U10732 (N_10732,N_10116,N_10107);
xnor U10733 (N_10733,N_10014,N_10396);
xor U10734 (N_10734,N_10230,N_10021);
or U10735 (N_10735,N_10229,N_10245);
xor U10736 (N_10736,N_10258,N_10120);
or U10737 (N_10737,N_10261,N_10196);
nor U10738 (N_10738,N_10378,N_10475);
xnor U10739 (N_10739,N_10124,N_10161);
or U10740 (N_10740,N_10348,N_10432);
and U10741 (N_10741,N_10436,N_10401);
xnor U10742 (N_10742,N_10274,N_10053);
or U10743 (N_10743,N_10368,N_10089);
nand U10744 (N_10744,N_10301,N_10054);
nand U10745 (N_10745,N_10489,N_10256);
nand U10746 (N_10746,N_10481,N_10087);
nor U10747 (N_10747,N_10153,N_10133);
xnor U10748 (N_10748,N_10372,N_10407);
and U10749 (N_10749,N_10428,N_10334);
or U10750 (N_10750,N_10358,N_10176);
or U10751 (N_10751,N_10210,N_10496);
nand U10752 (N_10752,N_10013,N_10218);
and U10753 (N_10753,N_10484,N_10075);
xnor U10754 (N_10754,N_10431,N_10327);
and U10755 (N_10755,N_10097,N_10399);
and U10756 (N_10756,N_10277,N_10436);
nor U10757 (N_10757,N_10364,N_10467);
and U10758 (N_10758,N_10441,N_10265);
and U10759 (N_10759,N_10176,N_10172);
xor U10760 (N_10760,N_10350,N_10322);
nand U10761 (N_10761,N_10198,N_10042);
xor U10762 (N_10762,N_10183,N_10019);
nor U10763 (N_10763,N_10013,N_10167);
or U10764 (N_10764,N_10177,N_10458);
or U10765 (N_10765,N_10145,N_10244);
xnor U10766 (N_10766,N_10261,N_10027);
nor U10767 (N_10767,N_10315,N_10239);
nor U10768 (N_10768,N_10409,N_10481);
xor U10769 (N_10769,N_10483,N_10204);
xor U10770 (N_10770,N_10355,N_10430);
nand U10771 (N_10771,N_10108,N_10317);
xor U10772 (N_10772,N_10349,N_10317);
or U10773 (N_10773,N_10362,N_10168);
nand U10774 (N_10774,N_10405,N_10332);
or U10775 (N_10775,N_10050,N_10328);
or U10776 (N_10776,N_10458,N_10312);
nand U10777 (N_10777,N_10442,N_10374);
nand U10778 (N_10778,N_10406,N_10035);
nor U10779 (N_10779,N_10031,N_10391);
and U10780 (N_10780,N_10250,N_10092);
nand U10781 (N_10781,N_10363,N_10057);
and U10782 (N_10782,N_10344,N_10039);
nor U10783 (N_10783,N_10316,N_10208);
xnor U10784 (N_10784,N_10472,N_10289);
nand U10785 (N_10785,N_10070,N_10029);
nor U10786 (N_10786,N_10337,N_10194);
xnor U10787 (N_10787,N_10011,N_10122);
or U10788 (N_10788,N_10379,N_10298);
nand U10789 (N_10789,N_10130,N_10489);
nor U10790 (N_10790,N_10227,N_10036);
xnor U10791 (N_10791,N_10012,N_10175);
xor U10792 (N_10792,N_10429,N_10224);
or U10793 (N_10793,N_10203,N_10363);
and U10794 (N_10794,N_10122,N_10260);
xor U10795 (N_10795,N_10456,N_10103);
or U10796 (N_10796,N_10183,N_10493);
and U10797 (N_10797,N_10069,N_10152);
or U10798 (N_10798,N_10287,N_10022);
xor U10799 (N_10799,N_10188,N_10002);
nor U10800 (N_10800,N_10421,N_10094);
xnor U10801 (N_10801,N_10173,N_10057);
nand U10802 (N_10802,N_10103,N_10024);
nand U10803 (N_10803,N_10023,N_10077);
nor U10804 (N_10804,N_10392,N_10050);
and U10805 (N_10805,N_10350,N_10059);
nor U10806 (N_10806,N_10302,N_10473);
and U10807 (N_10807,N_10200,N_10339);
or U10808 (N_10808,N_10326,N_10202);
and U10809 (N_10809,N_10275,N_10419);
nor U10810 (N_10810,N_10384,N_10128);
and U10811 (N_10811,N_10091,N_10170);
or U10812 (N_10812,N_10137,N_10264);
nor U10813 (N_10813,N_10176,N_10065);
and U10814 (N_10814,N_10008,N_10028);
or U10815 (N_10815,N_10104,N_10041);
nor U10816 (N_10816,N_10162,N_10484);
and U10817 (N_10817,N_10149,N_10434);
nand U10818 (N_10818,N_10463,N_10190);
xnor U10819 (N_10819,N_10173,N_10479);
nor U10820 (N_10820,N_10057,N_10495);
nand U10821 (N_10821,N_10101,N_10477);
nand U10822 (N_10822,N_10321,N_10165);
and U10823 (N_10823,N_10401,N_10047);
or U10824 (N_10824,N_10292,N_10193);
xor U10825 (N_10825,N_10259,N_10093);
xor U10826 (N_10826,N_10301,N_10112);
or U10827 (N_10827,N_10497,N_10338);
nand U10828 (N_10828,N_10497,N_10224);
xnor U10829 (N_10829,N_10294,N_10080);
nor U10830 (N_10830,N_10426,N_10051);
nor U10831 (N_10831,N_10262,N_10202);
nand U10832 (N_10832,N_10242,N_10421);
or U10833 (N_10833,N_10454,N_10170);
nor U10834 (N_10834,N_10283,N_10187);
nand U10835 (N_10835,N_10244,N_10123);
xnor U10836 (N_10836,N_10440,N_10140);
xnor U10837 (N_10837,N_10302,N_10314);
nor U10838 (N_10838,N_10295,N_10142);
nand U10839 (N_10839,N_10238,N_10034);
xnor U10840 (N_10840,N_10376,N_10152);
nor U10841 (N_10841,N_10189,N_10012);
nand U10842 (N_10842,N_10486,N_10018);
and U10843 (N_10843,N_10132,N_10295);
or U10844 (N_10844,N_10053,N_10426);
nand U10845 (N_10845,N_10123,N_10273);
or U10846 (N_10846,N_10112,N_10270);
or U10847 (N_10847,N_10231,N_10113);
and U10848 (N_10848,N_10422,N_10115);
nor U10849 (N_10849,N_10392,N_10260);
or U10850 (N_10850,N_10386,N_10417);
xor U10851 (N_10851,N_10408,N_10296);
xnor U10852 (N_10852,N_10020,N_10282);
and U10853 (N_10853,N_10396,N_10422);
xor U10854 (N_10854,N_10479,N_10006);
xnor U10855 (N_10855,N_10064,N_10137);
and U10856 (N_10856,N_10431,N_10074);
nor U10857 (N_10857,N_10379,N_10254);
and U10858 (N_10858,N_10085,N_10002);
nand U10859 (N_10859,N_10431,N_10241);
and U10860 (N_10860,N_10360,N_10232);
xor U10861 (N_10861,N_10163,N_10201);
xnor U10862 (N_10862,N_10290,N_10102);
nor U10863 (N_10863,N_10346,N_10411);
and U10864 (N_10864,N_10158,N_10457);
nand U10865 (N_10865,N_10313,N_10302);
and U10866 (N_10866,N_10346,N_10017);
nor U10867 (N_10867,N_10070,N_10192);
nand U10868 (N_10868,N_10325,N_10195);
or U10869 (N_10869,N_10301,N_10011);
nand U10870 (N_10870,N_10129,N_10290);
and U10871 (N_10871,N_10431,N_10276);
nand U10872 (N_10872,N_10271,N_10393);
or U10873 (N_10873,N_10129,N_10473);
and U10874 (N_10874,N_10392,N_10234);
or U10875 (N_10875,N_10443,N_10239);
nor U10876 (N_10876,N_10455,N_10012);
nor U10877 (N_10877,N_10271,N_10354);
nand U10878 (N_10878,N_10168,N_10020);
nand U10879 (N_10879,N_10140,N_10021);
nand U10880 (N_10880,N_10352,N_10189);
and U10881 (N_10881,N_10262,N_10133);
nor U10882 (N_10882,N_10410,N_10115);
and U10883 (N_10883,N_10381,N_10266);
or U10884 (N_10884,N_10218,N_10190);
nand U10885 (N_10885,N_10381,N_10149);
and U10886 (N_10886,N_10255,N_10337);
nand U10887 (N_10887,N_10178,N_10032);
and U10888 (N_10888,N_10265,N_10254);
xnor U10889 (N_10889,N_10341,N_10398);
or U10890 (N_10890,N_10376,N_10125);
nand U10891 (N_10891,N_10095,N_10417);
nand U10892 (N_10892,N_10171,N_10081);
nand U10893 (N_10893,N_10072,N_10319);
nand U10894 (N_10894,N_10377,N_10043);
or U10895 (N_10895,N_10252,N_10083);
or U10896 (N_10896,N_10434,N_10425);
xor U10897 (N_10897,N_10024,N_10015);
or U10898 (N_10898,N_10309,N_10086);
and U10899 (N_10899,N_10420,N_10170);
nand U10900 (N_10900,N_10362,N_10178);
or U10901 (N_10901,N_10329,N_10021);
or U10902 (N_10902,N_10484,N_10431);
xnor U10903 (N_10903,N_10459,N_10375);
nand U10904 (N_10904,N_10327,N_10033);
nor U10905 (N_10905,N_10298,N_10093);
and U10906 (N_10906,N_10220,N_10241);
xnor U10907 (N_10907,N_10117,N_10228);
and U10908 (N_10908,N_10417,N_10182);
nor U10909 (N_10909,N_10191,N_10133);
or U10910 (N_10910,N_10111,N_10432);
nor U10911 (N_10911,N_10138,N_10472);
xor U10912 (N_10912,N_10035,N_10448);
nand U10913 (N_10913,N_10245,N_10006);
nand U10914 (N_10914,N_10234,N_10225);
and U10915 (N_10915,N_10422,N_10055);
xnor U10916 (N_10916,N_10232,N_10004);
and U10917 (N_10917,N_10014,N_10313);
nand U10918 (N_10918,N_10288,N_10233);
xor U10919 (N_10919,N_10340,N_10115);
nor U10920 (N_10920,N_10199,N_10376);
xnor U10921 (N_10921,N_10223,N_10007);
xnor U10922 (N_10922,N_10463,N_10496);
xor U10923 (N_10923,N_10236,N_10432);
nand U10924 (N_10924,N_10120,N_10306);
nand U10925 (N_10925,N_10377,N_10401);
nor U10926 (N_10926,N_10174,N_10038);
nand U10927 (N_10927,N_10261,N_10331);
or U10928 (N_10928,N_10213,N_10090);
nand U10929 (N_10929,N_10439,N_10056);
nor U10930 (N_10930,N_10392,N_10215);
or U10931 (N_10931,N_10378,N_10496);
xor U10932 (N_10932,N_10403,N_10092);
xnor U10933 (N_10933,N_10415,N_10452);
and U10934 (N_10934,N_10496,N_10058);
nand U10935 (N_10935,N_10496,N_10114);
nor U10936 (N_10936,N_10261,N_10404);
xor U10937 (N_10937,N_10441,N_10341);
or U10938 (N_10938,N_10376,N_10334);
nor U10939 (N_10939,N_10284,N_10492);
nand U10940 (N_10940,N_10419,N_10042);
and U10941 (N_10941,N_10162,N_10314);
and U10942 (N_10942,N_10468,N_10073);
nor U10943 (N_10943,N_10232,N_10023);
and U10944 (N_10944,N_10444,N_10147);
xor U10945 (N_10945,N_10336,N_10057);
nor U10946 (N_10946,N_10230,N_10198);
nand U10947 (N_10947,N_10035,N_10265);
or U10948 (N_10948,N_10184,N_10042);
nor U10949 (N_10949,N_10214,N_10466);
xnor U10950 (N_10950,N_10225,N_10494);
and U10951 (N_10951,N_10359,N_10001);
xor U10952 (N_10952,N_10209,N_10386);
or U10953 (N_10953,N_10003,N_10340);
nor U10954 (N_10954,N_10149,N_10008);
nand U10955 (N_10955,N_10205,N_10249);
xor U10956 (N_10956,N_10124,N_10242);
nand U10957 (N_10957,N_10025,N_10123);
nand U10958 (N_10958,N_10226,N_10148);
xnor U10959 (N_10959,N_10369,N_10420);
nor U10960 (N_10960,N_10308,N_10023);
nor U10961 (N_10961,N_10115,N_10124);
and U10962 (N_10962,N_10286,N_10108);
nand U10963 (N_10963,N_10410,N_10427);
or U10964 (N_10964,N_10045,N_10365);
or U10965 (N_10965,N_10373,N_10247);
nand U10966 (N_10966,N_10358,N_10094);
and U10967 (N_10967,N_10150,N_10010);
nand U10968 (N_10968,N_10110,N_10404);
nor U10969 (N_10969,N_10004,N_10175);
nand U10970 (N_10970,N_10423,N_10254);
xor U10971 (N_10971,N_10157,N_10113);
or U10972 (N_10972,N_10339,N_10082);
and U10973 (N_10973,N_10130,N_10179);
and U10974 (N_10974,N_10078,N_10253);
nor U10975 (N_10975,N_10441,N_10003);
nor U10976 (N_10976,N_10117,N_10398);
and U10977 (N_10977,N_10432,N_10134);
xnor U10978 (N_10978,N_10308,N_10309);
nand U10979 (N_10979,N_10191,N_10224);
nor U10980 (N_10980,N_10473,N_10446);
nand U10981 (N_10981,N_10495,N_10388);
and U10982 (N_10982,N_10418,N_10262);
nor U10983 (N_10983,N_10011,N_10062);
nand U10984 (N_10984,N_10194,N_10050);
nor U10985 (N_10985,N_10002,N_10400);
nor U10986 (N_10986,N_10338,N_10360);
nand U10987 (N_10987,N_10160,N_10485);
xnor U10988 (N_10988,N_10196,N_10343);
or U10989 (N_10989,N_10214,N_10304);
nor U10990 (N_10990,N_10348,N_10483);
nand U10991 (N_10991,N_10027,N_10250);
xnor U10992 (N_10992,N_10393,N_10465);
nand U10993 (N_10993,N_10336,N_10271);
xnor U10994 (N_10994,N_10257,N_10017);
nand U10995 (N_10995,N_10481,N_10318);
or U10996 (N_10996,N_10363,N_10304);
nor U10997 (N_10997,N_10469,N_10259);
and U10998 (N_10998,N_10267,N_10217);
or U10999 (N_10999,N_10177,N_10361);
and U11000 (N_11000,N_10523,N_10573);
nor U11001 (N_11001,N_10647,N_10673);
or U11002 (N_11002,N_10782,N_10519);
nor U11003 (N_11003,N_10643,N_10876);
or U11004 (N_11004,N_10735,N_10669);
and U11005 (N_11005,N_10741,N_10863);
nand U11006 (N_11006,N_10727,N_10815);
nand U11007 (N_11007,N_10611,N_10682);
xor U11008 (N_11008,N_10506,N_10587);
and U11009 (N_11009,N_10999,N_10685);
xnor U11010 (N_11010,N_10770,N_10839);
nand U11011 (N_11011,N_10914,N_10942);
nand U11012 (N_11012,N_10624,N_10882);
xor U11013 (N_11013,N_10631,N_10531);
nor U11014 (N_11014,N_10500,N_10540);
xnor U11015 (N_11015,N_10802,N_10684);
or U11016 (N_11016,N_10671,N_10964);
nor U11017 (N_11017,N_10695,N_10891);
xor U11018 (N_11018,N_10849,N_10790);
xnor U11019 (N_11019,N_10653,N_10869);
nand U11020 (N_11020,N_10772,N_10524);
xnor U11021 (N_11021,N_10608,N_10638);
nor U11022 (N_11022,N_10726,N_10640);
nand U11023 (N_11023,N_10875,N_10689);
xor U11024 (N_11024,N_10541,N_10976);
xor U11025 (N_11025,N_10562,N_10621);
nor U11026 (N_11026,N_10829,N_10992);
and U11027 (N_11027,N_10796,N_10950);
nand U11028 (N_11028,N_10502,N_10730);
nor U11029 (N_11029,N_10605,N_10873);
xor U11030 (N_11030,N_10901,N_10517);
nor U11031 (N_11031,N_10812,N_10819);
and U11032 (N_11032,N_10826,N_10632);
or U11033 (N_11033,N_10574,N_10538);
or U11034 (N_11034,N_10745,N_10867);
nor U11035 (N_11035,N_10855,N_10748);
xnor U11036 (N_11036,N_10586,N_10791);
nor U11037 (N_11037,N_10533,N_10995);
nor U11038 (N_11038,N_10902,N_10807);
nor U11039 (N_11039,N_10732,N_10967);
and U11040 (N_11040,N_10532,N_10527);
and U11041 (N_11041,N_10809,N_10751);
or U11042 (N_11042,N_10639,N_10700);
nand U11043 (N_11043,N_10825,N_10589);
nor U11044 (N_11044,N_10559,N_10549);
and U11045 (N_11045,N_10868,N_10686);
nor U11046 (N_11046,N_10958,N_10646);
and U11047 (N_11047,N_10762,N_10957);
xor U11048 (N_11048,N_10593,N_10924);
and U11049 (N_11049,N_10652,N_10966);
and U11050 (N_11050,N_10920,N_10766);
or U11051 (N_11051,N_10814,N_10936);
and U11052 (N_11052,N_10596,N_10721);
or U11053 (N_11053,N_10838,N_10597);
and U11054 (N_11054,N_10656,N_10630);
nand U11055 (N_11055,N_10680,N_10548);
or U11056 (N_11056,N_10827,N_10921);
nand U11057 (N_11057,N_10832,N_10581);
nor U11058 (N_11058,N_10828,N_10811);
and U11059 (N_11059,N_10717,N_10505);
nor U11060 (N_11060,N_10607,N_10723);
nand U11061 (N_11061,N_10842,N_10883);
nand U11062 (N_11062,N_10692,N_10663);
nor U11063 (N_11063,N_10767,N_10906);
and U11064 (N_11064,N_10918,N_10810);
and U11065 (N_11065,N_10895,N_10637);
and U11066 (N_11066,N_10856,N_10709);
and U11067 (N_11067,N_10785,N_10951);
nand U11068 (N_11068,N_10623,N_10563);
nand U11069 (N_11069,N_10705,N_10558);
nor U11070 (N_11070,N_10986,N_10853);
nor U11071 (N_11071,N_10620,N_10716);
nor U11072 (N_11072,N_10679,N_10687);
nand U11073 (N_11073,N_10744,N_10820);
nor U11074 (N_11074,N_10696,N_10897);
nor U11075 (N_11075,N_10534,N_10583);
nor U11076 (N_11076,N_10889,N_10569);
nor U11077 (N_11077,N_10953,N_10850);
nand U11078 (N_11078,N_10552,N_10779);
and U11079 (N_11079,N_10893,N_10601);
nor U11080 (N_11080,N_10852,N_10940);
or U11081 (N_11081,N_10930,N_10715);
nand U11082 (N_11082,N_10834,N_10746);
and U11083 (N_11083,N_10645,N_10778);
or U11084 (N_11084,N_10719,N_10606);
or U11085 (N_11085,N_10994,N_10675);
xor U11086 (N_11086,N_10773,N_10835);
nand U11087 (N_11087,N_10823,N_10511);
nand U11088 (N_11088,N_10763,N_10555);
or U11089 (N_11089,N_10960,N_10602);
nand U11090 (N_11090,N_10818,N_10697);
and U11091 (N_11091,N_10981,N_10968);
nor U11092 (N_11092,N_10514,N_10703);
or U11093 (N_11093,N_10961,N_10526);
nor U11094 (N_11094,N_10765,N_10948);
or U11095 (N_11095,N_10604,N_10707);
or U11096 (N_11096,N_10939,N_10972);
and U11097 (N_11097,N_10592,N_10668);
and U11098 (N_11098,N_10963,N_10641);
nor U11099 (N_11099,N_10793,N_10676);
and U11100 (N_11100,N_10616,N_10561);
nor U11101 (N_11101,N_10844,N_10898);
nand U11102 (N_11102,N_10980,N_10702);
xnor U11103 (N_11103,N_10714,N_10996);
and U11104 (N_11104,N_10613,N_10911);
and U11105 (N_11105,N_10938,N_10629);
xnor U11106 (N_11106,N_10781,N_10739);
nor U11107 (N_11107,N_10708,N_10733);
or U11108 (N_11108,N_10545,N_10642);
nand U11109 (N_11109,N_10947,N_10881);
xor U11110 (N_11110,N_10657,N_10627);
nand U11111 (N_11111,N_10982,N_10988);
and U11112 (N_11112,N_10927,N_10965);
or U11113 (N_11113,N_10774,N_10915);
or U11114 (N_11114,N_10580,N_10858);
and U11115 (N_11115,N_10599,N_10833);
xnor U11116 (N_11116,N_10694,N_10879);
nand U11117 (N_11117,N_10722,N_10542);
xor U11118 (N_11118,N_10576,N_10822);
nor U11119 (N_11119,N_10567,N_10738);
nand U11120 (N_11120,N_10990,N_10507);
and U11121 (N_11121,N_10768,N_10720);
or U11122 (N_11122,N_10670,N_10614);
nor U11123 (N_11123,N_10677,N_10813);
and U11124 (N_11124,N_10859,N_10848);
nand U11125 (N_11125,N_10530,N_10655);
nor U11126 (N_11126,N_10619,N_10794);
or U11127 (N_11127,N_10931,N_10634);
or U11128 (N_11128,N_10956,N_10536);
and U11129 (N_11129,N_10887,N_10740);
and U11130 (N_11130,N_10821,N_10591);
xor U11131 (N_11131,N_10520,N_10556);
or U11132 (N_11132,N_10909,N_10760);
nand U11133 (N_11133,N_10649,N_10575);
xor U11134 (N_11134,N_10713,N_10905);
nand U11135 (N_11135,N_10952,N_10513);
xor U11136 (N_11136,N_10518,N_10870);
or U11137 (N_11137,N_10725,N_10789);
or U11138 (N_11138,N_10554,N_10550);
and U11139 (N_11139,N_10626,N_10742);
and U11140 (N_11140,N_10805,N_10525);
and U11141 (N_11141,N_10515,N_10547);
nand U11142 (N_11142,N_10622,N_10764);
nor U11143 (N_11143,N_10658,N_10831);
xor U11144 (N_11144,N_10864,N_10955);
nand U11145 (N_11145,N_10934,N_10737);
nor U11146 (N_11146,N_10880,N_10866);
xnor U11147 (N_11147,N_10944,N_10937);
xnor U11148 (N_11148,N_10628,N_10512);
and U11149 (N_11149,N_10516,N_10693);
xor U11150 (N_11150,N_10816,N_10617);
or U11151 (N_11151,N_10691,N_10557);
xor U11152 (N_11152,N_10800,N_10706);
and U11153 (N_11153,N_10836,N_10878);
and U11154 (N_11154,N_10754,N_10598);
xnor U11155 (N_11155,N_10749,N_10798);
xor U11156 (N_11156,N_10943,N_10734);
nand U11157 (N_11157,N_10929,N_10681);
xnor U11158 (N_11158,N_10997,N_10989);
or U11159 (N_11159,N_10962,N_10568);
and U11160 (N_11160,N_10872,N_10894);
and U11161 (N_11161,N_10886,N_10933);
xnor U11162 (N_11162,N_10651,N_10660);
xnor U11163 (N_11163,N_10570,N_10854);
or U11164 (N_11164,N_10945,N_10664);
or U11165 (N_11165,N_10701,N_10539);
nor U11166 (N_11166,N_10600,N_10806);
or U11167 (N_11167,N_10690,N_10529);
nand U11168 (N_11168,N_10970,N_10871);
or U11169 (N_11169,N_10577,N_10729);
nand U11170 (N_11170,N_10851,N_10743);
nor U11171 (N_11171,N_10799,N_10916);
or U11172 (N_11172,N_10588,N_10801);
nand U11173 (N_11173,N_10769,N_10877);
nand U11174 (N_11174,N_10578,N_10824);
or U11175 (N_11175,N_10925,N_10503);
nand U11176 (N_11176,N_10508,N_10932);
and U11177 (N_11177,N_10712,N_10792);
nor U11178 (N_11178,N_10625,N_10987);
or U11179 (N_11179,N_10797,N_10564);
or U11180 (N_11180,N_10991,N_10609);
xor U11181 (N_11181,N_10718,N_10688);
xor U11182 (N_11182,N_10803,N_10843);
and U11183 (N_11183,N_10666,N_10857);
xnor U11184 (N_11184,N_10846,N_10662);
nand U11185 (N_11185,N_10946,N_10636);
or U11186 (N_11186,N_10674,N_10923);
nand U11187 (N_11187,N_10584,N_10845);
nand U11188 (N_11188,N_10777,N_10750);
and U11189 (N_11189,N_10775,N_10973);
nor U11190 (N_11190,N_10941,N_10566);
or U11191 (N_11191,N_10665,N_10635);
nand U11192 (N_11192,N_10678,N_10710);
and U11193 (N_11193,N_10585,N_10683);
nor U11194 (N_11194,N_10998,N_10753);
xor U11195 (N_11195,N_10786,N_10919);
or U11196 (N_11196,N_10904,N_10757);
or U11197 (N_11197,N_10565,N_10771);
xnor U11198 (N_11198,N_10892,N_10975);
and U11199 (N_11199,N_10747,N_10603);
nand U11200 (N_11200,N_10926,N_10908);
nand U11201 (N_11201,N_10704,N_10837);
nand U11202 (N_11202,N_10928,N_10874);
nor U11203 (N_11203,N_10935,N_10731);
and U11204 (N_11204,N_10978,N_10659);
nand U11205 (N_11205,N_10537,N_10644);
or U11206 (N_11206,N_10612,N_10535);
nor U11207 (N_11207,N_10654,N_10787);
nor U11208 (N_11208,N_10900,N_10724);
xor U11209 (N_11209,N_10840,N_10817);
or U11210 (N_11210,N_10756,N_10594);
nor U11211 (N_11211,N_10865,N_10788);
nand U11212 (N_11212,N_10841,N_10830);
xnor U11213 (N_11213,N_10755,N_10985);
and U11214 (N_11214,N_10862,N_10521);
and U11215 (N_11215,N_10504,N_10903);
nand U11216 (N_11216,N_10860,N_10590);
xor U11217 (N_11217,N_10912,N_10913);
and U11218 (N_11218,N_10808,N_10780);
nor U11219 (N_11219,N_10667,N_10672);
and U11220 (N_11220,N_10759,N_10633);
and U11221 (N_11221,N_10661,N_10551);
nor U11222 (N_11222,N_10917,N_10553);
or U11223 (N_11223,N_10579,N_10969);
nor U11224 (N_11224,N_10784,N_10544);
and U11225 (N_11225,N_10907,N_10650);
xnor U11226 (N_11226,N_10910,N_10528);
and U11227 (N_11227,N_10698,N_10776);
nand U11228 (N_11228,N_10648,N_10595);
nand U11229 (N_11229,N_10509,N_10959);
or U11230 (N_11230,N_10501,N_10977);
and U11231 (N_11231,N_10522,N_10752);
and U11232 (N_11232,N_10783,N_10949);
or U11233 (N_11233,N_10560,N_10899);
nand U11234 (N_11234,N_10983,N_10699);
or U11235 (N_11235,N_10971,N_10979);
and U11236 (N_11236,N_10572,N_10543);
xor U11237 (N_11237,N_10615,N_10546);
and U11238 (N_11238,N_10888,N_10711);
and U11239 (N_11239,N_10610,N_10954);
xor U11240 (N_11240,N_10571,N_10885);
nor U11241 (N_11241,N_10804,N_10896);
or U11242 (N_11242,N_10993,N_10984);
nand U11243 (N_11243,N_10884,N_10618);
xor U11244 (N_11244,N_10582,N_10728);
xor U11245 (N_11245,N_10974,N_10758);
xnor U11246 (N_11246,N_10795,N_10736);
xnor U11247 (N_11247,N_10761,N_10890);
nand U11248 (N_11248,N_10861,N_10922);
xnor U11249 (N_11249,N_10847,N_10510);
xnor U11250 (N_11250,N_10503,N_10987);
or U11251 (N_11251,N_10584,N_10548);
and U11252 (N_11252,N_10960,N_10646);
and U11253 (N_11253,N_10599,N_10588);
nor U11254 (N_11254,N_10939,N_10510);
nand U11255 (N_11255,N_10609,N_10900);
and U11256 (N_11256,N_10560,N_10866);
or U11257 (N_11257,N_10766,N_10662);
and U11258 (N_11258,N_10811,N_10997);
or U11259 (N_11259,N_10663,N_10968);
nand U11260 (N_11260,N_10854,N_10806);
nand U11261 (N_11261,N_10675,N_10865);
nand U11262 (N_11262,N_10566,N_10538);
and U11263 (N_11263,N_10987,N_10917);
and U11264 (N_11264,N_10859,N_10627);
or U11265 (N_11265,N_10552,N_10857);
xor U11266 (N_11266,N_10847,N_10972);
nor U11267 (N_11267,N_10781,N_10600);
nor U11268 (N_11268,N_10682,N_10866);
nand U11269 (N_11269,N_10905,N_10850);
nand U11270 (N_11270,N_10609,N_10675);
or U11271 (N_11271,N_10633,N_10864);
nand U11272 (N_11272,N_10593,N_10928);
and U11273 (N_11273,N_10838,N_10888);
and U11274 (N_11274,N_10642,N_10952);
nor U11275 (N_11275,N_10699,N_10730);
or U11276 (N_11276,N_10721,N_10578);
xor U11277 (N_11277,N_10665,N_10720);
xnor U11278 (N_11278,N_10751,N_10957);
or U11279 (N_11279,N_10710,N_10546);
nand U11280 (N_11280,N_10679,N_10964);
xnor U11281 (N_11281,N_10752,N_10538);
or U11282 (N_11282,N_10677,N_10734);
and U11283 (N_11283,N_10812,N_10766);
xor U11284 (N_11284,N_10720,N_10731);
xor U11285 (N_11285,N_10563,N_10769);
or U11286 (N_11286,N_10507,N_10789);
xnor U11287 (N_11287,N_10947,N_10853);
nand U11288 (N_11288,N_10729,N_10827);
and U11289 (N_11289,N_10769,N_10793);
or U11290 (N_11290,N_10977,N_10885);
and U11291 (N_11291,N_10584,N_10928);
xnor U11292 (N_11292,N_10950,N_10655);
or U11293 (N_11293,N_10717,N_10808);
nand U11294 (N_11294,N_10553,N_10576);
and U11295 (N_11295,N_10955,N_10671);
nand U11296 (N_11296,N_10956,N_10620);
nor U11297 (N_11297,N_10598,N_10911);
and U11298 (N_11298,N_10899,N_10580);
or U11299 (N_11299,N_10580,N_10509);
xor U11300 (N_11300,N_10689,N_10527);
or U11301 (N_11301,N_10516,N_10514);
nand U11302 (N_11302,N_10613,N_10869);
or U11303 (N_11303,N_10875,N_10655);
xnor U11304 (N_11304,N_10679,N_10937);
nor U11305 (N_11305,N_10830,N_10708);
nor U11306 (N_11306,N_10664,N_10930);
nand U11307 (N_11307,N_10753,N_10978);
xor U11308 (N_11308,N_10692,N_10852);
nor U11309 (N_11309,N_10680,N_10759);
or U11310 (N_11310,N_10989,N_10893);
and U11311 (N_11311,N_10804,N_10531);
nor U11312 (N_11312,N_10609,N_10969);
nor U11313 (N_11313,N_10827,N_10710);
or U11314 (N_11314,N_10954,N_10850);
nand U11315 (N_11315,N_10952,N_10538);
or U11316 (N_11316,N_10703,N_10518);
or U11317 (N_11317,N_10975,N_10645);
and U11318 (N_11318,N_10501,N_10578);
xor U11319 (N_11319,N_10992,N_10918);
and U11320 (N_11320,N_10843,N_10567);
and U11321 (N_11321,N_10685,N_10908);
nand U11322 (N_11322,N_10821,N_10808);
and U11323 (N_11323,N_10828,N_10672);
or U11324 (N_11324,N_10864,N_10629);
and U11325 (N_11325,N_10622,N_10709);
and U11326 (N_11326,N_10549,N_10741);
xnor U11327 (N_11327,N_10671,N_10855);
or U11328 (N_11328,N_10515,N_10789);
xor U11329 (N_11329,N_10984,N_10950);
nand U11330 (N_11330,N_10861,N_10816);
nand U11331 (N_11331,N_10763,N_10853);
or U11332 (N_11332,N_10512,N_10726);
xnor U11333 (N_11333,N_10861,N_10813);
or U11334 (N_11334,N_10737,N_10887);
xnor U11335 (N_11335,N_10540,N_10933);
nor U11336 (N_11336,N_10926,N_10875);
and U11337 (N_11337,N_10665,N_10845);
nor U11338 (N_11338,N_10807,N_10965);
nand U11339 (N_11339,N_10619,N_10910);
and U11340 (N_11340,N_10830,N_10729);
and U11341 (N_11341,N_10609,N_10589);
and U11342 (N_11342,N_10677,N_10575);
xnor U11343 (N_11343,N_10906,N_10796);
nand U11344 (N_11344,N_10983,N_10533);
and U11345 (N_11345,N_10825,N_10862);
and U11346 (N_11346,N_10882,N_10811);
or U11347 (N_11347,N_10624,N_10978);
nand U11348 (N_11348,N_10616,N_10859);
and U11349 (N_11349,N_10799,N_10687);
and U11350 (N_11350,N_10853,N_10945);
nor U11351 (N_11351,N_10874,N_10810);
xnor U11352 (N_11352,N_10766,N_10955);
xor U11353 (N_11353,N_10933,N_10928);
or U11354 (N_11354,N_10735,N_10967);
and U11355 (N_11355,N_10879,N_10731);
and U11356 (N_11356,N_10566,N_10578);
xnor U11357 (N_11357,N_10627,N_10507);
and U11358 (N_11358,N_10539,N_10506);
nand U11359 (N_11359,N_10900,N_10541);
xor U11360 (N_11360,N_10965,N_10530);
and U11361 (N_11361,N_10826,N_10668);
xnor U11362 (N_11362,N_10835,N_10880);
nor U11363 (N_11363,N_10746,N_10566);
and U11364 (N_11364,N_10621,N_10792);
and U11365 (N_11365,N_10986,N_10955);
nand U11366 (N_11366,N_10655,N_10967);
or U11367 (N_11367,N_10903,N_10968);
or U11368 (N_11368,N_10833,N_10561);
xor U11369 (N_11369,N_10588,N_10997);
nor U11370 (N_11370,N_10978,N_10976);
xor U11371 (N_11371,N_10654,N_10891);
nor U11372 (N_11372,N_10809,N_10683);
nand U11373 (N_11373,N_10673,N_10668);
nor U11374 (N_11374,N_10808,N_10750);
or U11375 (N_11375,N_10799,N_10525);
xnor U11376 (N_11376,N_10870,N_10580);
xor U11377 (N_11377,N_10502,N_10622);
or U11378 (N_11378,N_10550,N_10507);
nor U11379 (N_11379,N_10990,N_10522);
nand U11380 (N_11380,N_10937,N_10622);
nor U11381 (N_11381,N_10503,N_10790);
xnor U11382 (N_11382,N_10932,N_10887);
xor U11383 (N_11383,N_10611,N_10932);
nor U11384 (N_11384,N_10879,N_10661);
nor U11385 (N_11385,N_10855,N_10951);
nand U11386 (N_11386,N_10670,N_10773);
and U11387 (N_11387,N_10870,N_10591);
nand U11388 (N_11388,N_10989,N_10980);
xor U11389 (N_11389,N_10604,N_10718);
nand U11390 (N_11390,N_10683,N_10510);
nor U11391 (N_11391,N_10622,N_10584);
or U11392 (N_11392,N_10597,N_10903);
nor U11393 (N_11393,N_10504,N_10723);
xnor U11394 (N_11394,N_10590,N_10551);
or U11395 (N_11395,N_10506,N_10781);
and U11396 (N_11396,N_10939,N_10611);
or U11397 (N_11397,N_10817,N_10700);
and U11398 (N_11398,N_10802,N_10623);
or U11399 (N_11399,N_10762,N_10999);
nor U11400 (N_11400,N_10589,N_10809);
nand U11401 (N_11401,N_10686,N_10505);
or U11402 (N_11402,N_10786,N_10931);
nor U11403 (N_11403,N_10651,N_10588);
and U11404 (N_11404,N_10667,N_10954);
and U11405 (N_11405,N_10798,N_10815);
xor U11406 (N_11406,N_10514,N_10607);
and U11407 (N_11407,N_10986,N_10782);
and U11408 (N_11408,N_10845,N_10675);
and U11409 (N_11409,N_10639,N_10797);
xnor U11410 (N_11410,N_10748,N_10765);
xnor U11411 (N_11411,N_10571,N_10575);
nand U11412 (N_11412,N_10815,N_10998);
nor U11413 (N_11413,N_10828,N_10666);
or U11414 (N_11414,N_10538,N_10596);
nand U11415 (N_11415,N_10861,N_10530);
nand U11416 (N_11416,N_10608,N_10933);
and U11417 (N_11417,N_10965,N_10629);
xor U11418 (N_11418,N_10521,N_10956);
xnor U11419 (N_11419,N_10739,N_10799);
nand U11420 (N_11420,N_10993,N_10754);
nor U11421 (N_11421,N_10828,N_10860);
xor U11422 (N_11422,N_10640,N_10549);
xnor U11423 (N_11423,N_10875,N_10864);
or U11424 (N_11424,N_10881,N_10798);
xor U11425 (N_11425,N_10941,N_10756);
or U11426 (N_11426,N_10943,N_10976);
xor U11427 (N_11427,N_10591,N_10859);
nor U11428 (N_11428,N_10871,N_10931);
nor U11429 (N_11429,N_10929,N_10562);
nand U11430 (N_11430,N_10628,N_10983);
nor U11431 (N_11431,N_10966,N_10511);
xor U11432 (N_11432,N_10871,N_10581);
nor U11433 (N_11433,N_10933,N_10918);
nand U11434 (N_11434,N_10630,N_10680);
or U11435 (N_11435,N_10966,N_10623);
or U11436 (N_11436,N_10539,N_10740);
nand U11437 (N_11437,N_10503,N_10538);
nor U11438 (N_11438,N_10962,N_10912);
nor U11439 (N_11439,N_10952,N_10955);
or U11440 (N_11440,N_10848,N_10943);
or U11441 (N_11441,N_10809,N_10578);
and U11442 (N_11442,N_10747,N_10568);
and U11443 (N_11443,N_10903,N_10527);
nand U11444 (N_11444,N_10810,N_10805);
xor U11445 (N_11445,N_10989,N_10917);
nand U11446 (N_11446,N_10721,N_10828);
nor U11447 (N_11447,N_10720,N_10761);
or U11448 (N_11448,N_10784,N_10622);
nor U11449 (N_11449,N_10976,N_10794);
xor U11450 (N_11450,N_10904,N_10659);
and U11451 (N_11451,N_10692,N_10735);
nand U11452 (N_11452,N_10945,N_10569);
nand U11453 (N_11453,N_10765,N_10662);
or U11454 (N_11454,N_10874,N_10582);
xor U11455 (N_11455,N_10809,N_10973);
xnor U11456 (N_11456,N_10545,N_10979);
xnor U11457 (N_11457,N_10579,N_10782);
nand U11458 (N_11458,N_10940,N_10559);
or U11459 (N_11459,N_10727,N_10867);
nor U11460 (N_11460,N_10833,N_10971);
nand U11461 (N_11461,N_10946,N_10877);
and U11462 (N_11462,N_10620,N_10651);
nand U11463 (N_11463,N_10676,N_10524);
nor U11464 (N_11464,N_10695,N_10571);
nor U11465 (N_11465,N_10634,N_10646);
or U11466 (N_11466,N_10592,N_10672);
and U11467 (N_11467,N_10913,N_10506);
and U11468 (N_11468,N_10805,N_10655);
and U11469 (N_11469,N_10827,N_10949);
nand U11470 (N_11470,N_10655,N_10873);
nor U11471 (N_11471,N_10694,N_10572);
and U11472 (N_11472,N_10660,N_10981);
or U11473 (N_11473,N_10555,N_10560);
or U11474 (N_11474,N_10965,N_10887);
and U11475 (N_11475,N_10864,N_10905);
xor U11476 (N_11476,N_10614,N_10778);
xor U11477 (N_11477,N_10992,N_10501);
nand U11478 (N_11478,N_10803,N_10813);
nor U11479 (N_11479,N_10787,N_10975);
and U11480 (N_11480,N_10801,N_10782);
nand U11481 (N_11481,N_10970,N_10853);
xor U11482 (N_11482,N_10838,N_10602);
xor U11483 (N_11483,N_10736,N_10836);
nand U11484 (N_11484,N_10578,N_10645);
nand U11485 (N_11485,N_10803,N_10611);
or U11486 (N_11486,N_10928,N_10961);
or U11487 (N_11487,N_10712,N_10747);
nand U11488 (N_11488,N_10929,N_10871);
nor U11489 (N_11489,N_10921,N_10524);
nand U11490 (N_11490,N_10746,N_10559);
nand U11491 (N_11491,N_10983,N_10991);
nor U11492 (N_11492,N_10946,N_10954);
xor U11493 (N_11493,N_10859,N_10617);
nor U11494 (N_11494,N_10633,N_10601);
or U11495 (N_11495,N_10701,N_10865);
nor U11496 (N_11496,N_10978,N_10931);
xor U11497 (N_11497,N_10931,N_10712);
or U11498 (N_11498,N_10675,N_10530);
nand U11499 (N_11499,N_10558,N_10507);
nor U11500 (N_11500,N_11157,N_11047);
nand U11501 (N_11501,N_11362,N_11076);
or U11502 (N_11502,N_11200,N_11368);
nand U11503 (N_11503,N_11271,N_11168);
xor U11504 (N_11504,N_11459,N_11172);
or U11505 (N_11505,N_11310,N_11451);
or U11506 (N_11506,N_11306,N_11301);
or U11507 (N_11507,N_11446,N_11018);
or U11508 (N_11508,N_11461,N_11097);
or U11509 (N_11509,N_11242,N_11291);
nor U11510 (N_11510,N_11014,N_11186);
nor U11511 (N_11511,N_11262,N_11385);
and U11512 (N_11512,N_11475,N_11119);
xnor U11513 (N_11513,N_11479,N_11332);
and U11514 (N_11514,N_11474,N_11419);
nor U11515 (N_11515,N_11095,N_11135);
and U11516 (N_11516,N_11358,N_11082);
xor U11517 (N_11517,N_11438,N_11366);
nor U11518 (N_11518,N_11276,N_11452);
xnor U11519 (N_11519,N_11233,N_11110);
nor U11520 (N_11520,N_11062,N_11315);
or U11521 (N_11521,N_11013,N_11052);
and U11522 (N_11522,N_11465,N_11123);
or U11523 (N_11523,N_11122,N_11004);
and U11524 (N_11524,N_11435,N_11484);
and U11525 (N_11525,N_11216,N_11169);
xor U11526 (N_11526,N_11182,N_11287);
or U11527 (N_11527,N_11305,N_11090);
or U11528 (N_11528,N_11179,N_11031);
nor U11529 (N_11529,N_11083,N_11250);
nor U11530 (N_11530,N_11388,N_11241);
and U11531 (N_11531,N_11458,N_11313);
or U11532 (N_11532,N_11338,N_11214);
nand U11533 (N_11533,N_11491,N_11273);
or U11534 (N_11534,N_11382,N_11220);
or U11535 (N_11535,N_11371,N_11333);
and U11536 (N_11536,N_11345,N_11208);
or U11537 (N_11537,N_11483,N_11405);
xor U11538 (N_11538,N_11225,N_11360);
xnor U11539 (N_11539,N_11425,N_11493);
xnor U11540 (N_11540,N_11196,N_11104);
or U11541 (N_11541,N_11245,N_11312);
xor U11542 (N_11542,N_11354,N_11327);
and U11543 (N_11543,N_11159,N_11392);
and U11544 (N_11544,N_11422,N_11290);
and U11545 (N_11545,N_11207,N_11117);
and U11546 (N_11546,N_11285,N_11228);
and U11547 (N_11547,N_11275,N_11028);
nor U11548 (N_11548,N_11416,N_11361);
and U11549 (N_11549,N_11486,N_11340);
nor U11550 (N_11550,N_11295,N_11341);
nand U11551 (N_11551,N_11077,N_11440);
or U11552 (N_11552,N_11330,N_11384);
or U11553 (N_11553,N_11442,N_11467);
or U11554 (N_11554,N_11150,N_11115);
nor U11555 (N_11555,N_11078,N_11443);
and U11556 (N_11556,N_11215,N_11421);
or U11557 (N_11557,N_11490,N_11365);
or U11558 (N_11558,N_11266,N_11041);
nor U11559 (N_11559,N_11171,N_11155);
nand U11560 (N_11560,N_11068,N_11012);
or U11561 (N_11561,N_11380,N_11434);
or U11562 (N_11562,N_11217,N_11057);
and U11563 (N_11563,N_11205,N_11302);
nand U11564 (N_11564,N_11218,N_11387);
nand U11565 (N_11565,N_11254,N_11370);
nor U11566 (N_11566,N_11274,N_11349);
nor U11567 (N_11567,N_11134,N_11386);
nor U11568 (N_11568,N_11269,N_11036);
nand U11569 (N_11569,N_11194,N_11282);
xnor U11570 (N_11570,N_11105,N_11042);
nand U11571 (N_11571,N_11178,N_11283);
or U11572 (N_11572,N_11255,N_11089);
nand U11573 (N_11573,N_11470,N_11058);
nand U11574 (N_11574,N_11297,N_11065);
and U11575 (N_11575,N_11079,N_11433);
nand U11576 (N_11576,N_11293,N_11067);
or U11577 (N_11577,N_11137,N_11001);
or U11578 (N_11578,N_11230,N_11267);
xnor U11579 (N_11579,N_11026,N_11175);
and U11580 (N_11580,N_11107,N_11351);
xor U11581 (N_11581,N_11292,N_11131);
nand U11582 (N_11582,N_11010,N_11053);
or U11583 (N_11583,N_11289,N_11002);
and U11584 (N_11584,N_11399,N_11303);
xnor U11585 (N_11585,N_11347,N_11198);
nand U11586 (N_11586,N_11396,N_11096);
nor U11587 (N_11587,N_11112,N_11211);
and U11588 (N_11588,N_11298,N_11085);
nor U11589 (N_11589,N_11258,N_11143);
or U11590 (N_11590,N_11174,N_11418);
or U11591 (N_11591,N_11180,N_11165);
or U11592 (N_11592,N_11232,N_11492);
xor U11593 (N_11593,N_11160,N_11444);
and U11594 (N_11594,N_11304,N_11049);
or U11595 (N_11595,N_11436,N_11356);
nor U11596 (N_11596,N_11447,N_11163);
or U11597 (N_11597,N_11206,N_11323);
xor U11598 (N_11598,N_11482,N_11229);
xor U11599 (N_11599,N_11209,N_11379);
nor U11600 (N_11600,N_11034,N_11322);
and U11601 (N_11601,N_11397,N_11035);
xor U11602 (N_11602,N_11264,N_11429);
xor U11603 (N_11603,N_11240,N_11226);
xnor U11604 (N_11604,N_11466,N_11191);
and U11605 (N_11605,N_11145,N_11251);
nor U11606 (N_11606,N_11268,N_11391);
nor U11607 (N_11607,N_11201,N_11390);
nor U11608 (N_11608,N_11183,N_11263);
nand U11609 (N_11609,N_11025,N_11389);
or U11610 (N_11610,N_11431,N_11044);
and U11611 (N_11611,N_11103,N_11128);
and U11612 (N_11612,N_11037,N_11480);
or U11613 (N_11613,N_11441,N_11113);
nand U11614 (N_11614,N_11412,N_11363);
nand U11615 (N_11615,N_11448,N_11496);
nand U11616 (N_11616,N_11093,N_11234);
and U11617 (N_11617,N_11005,N_11468);
nand U11618 (N_11618,N_11326,N_11141);
nor U11619 (N_11619,N_11087,N_11343);
xor U11620 (N_11620,N_11106,N_11202);
nor U11621 (N_11621,N_11478,N_11073);
nor U11622 (N_11622,N_11488,N_11350);
nand U11623 (N_11623,N_11147,N_11348);
nand U11624 (N_11624,N_11210,N_11063);
and U11625 (N_11625,N_11108,N_11040);
nor U11626 (N_11626,N_11219,N_11193);
and U11627 (N_11627,N_11265,N_11432);
xor U11628 (N_11628,N_11296,N_11092);
nor U11629 (N_11629,N_11158,N_11499);
and U11630 (N_11630,N_11357,N_11060);
xor U11631 (N_11631,N_11455,N_11235);
nor U11632 (N_11632,N_11056,N_11376);
xnor U11633 (N_11633,N_11006,N_11378);
nor U11634 (N_11634,N_11334,N_11227);
or U11635 (N_11635,N_11415,N_11142);
nand U11636 (N_11636,N_11102,N_11473);
nand U11637 (N_11637,N_11420,N_11030);
or U11638 (N_11638,N_11139,N_11055);
xor U11639 (N_11639,N_11253,N_11342);
and U11640 (N_11640,N_11329,N_11148);
nor U11641 (N_11641,N_11243,N_11111);
or U11642 (N_11642,N_11054,N_11279);
nand U11643 (N_11643,N_11048,N_11127);
nor U11644 (N_11644,N_11064,N_11314);
nor U11645 (N_11645,N_11395,N_11288);
or U11646 (N_11646,N_11213,N_11476);
nand U11647 (N_11647,N_11043,N_11080);
nor U11648 (N_11648,N_11430,N_11437);
xnor U11649 (N_11649,N_11132,N_11066);
and U11650 (N_11650,N_11318,N_11231);
and U11651 (N_11651,N_11339,N_11244);
nor U11652 (N_11652,N_11109,N_11469);
nand U11653 (N_11653,N_11317,N_11099);
xnor U11654 (N_11654,N_11003,N_11187);
nand U11655 (N_11655,N_11406,N_11411);
nor U11656 (N_11656,N_11221,N_11101);
or U11657 (N_11657,N_11404,N_11407);
or U11658 (N_11658,N_11118,N_11197);
nor U11659 (N_11659,N_11125,N_11324);
nor U11660 (N_11660,N_11427,N_11007);
nor U11661 (N_11661,N_11185,N_11033);
nor U11662 (N_11662,N_11015,N_11477);
nand U11663 (N_11663,N_11328,N_11204);
nand U11664 (N_11664,N_11029,N_11454);
nand U11665 (N_11665,N_11199,N_11166);
and U11666 (N_11666,N_11114,N_11249);
or U11667 (N_11667,N_11402,N_11272);
and U11668 (N_11668,N_11337,N_11375);
xor U11669 (N_11669,N_11364,N_11176);
or U11670 (N_11670,N_11321,N_11428);
nor U11671 (N_11671,N_11286,N_11481);
and U11672 (N_11672,N_11124,N_11236);
nand U11673 (N_11673,N_11355,N_11181);
nor U11674 (N_11674,N_11011,N_11140);
or U11675 (N_11675,N_11410,N_11032);
and U11676 (N_11676,N_11498,N_11038);
xor U11677 (N_11677,N_11335,N_11126);
and U11678 (N_11678,N_11472,N_11247);
xor U11679 (N_11679,N_11022,N_11116);
nor U11680 (N_11680,N_11308,N_11450);
xor U11681 (N_11681,N_11456,N_11462);
xor U11682 (N_11682,N_11426,N_11151);
xor U11683 (N_11683,N_11192,N_11280);
xor U11684 (N_11684,N_11203,N_11120);
or U11685 (N_11685,N_11189,N_11346);
and U11686 (N_11686,N_11069,N_11460);
nand U11687 (N_11687,N_11084,N_11146);
nor U11688 (N_11688,N_11374,N_11223);
or U11689 (N_11689,N_11161,N_11094);
and U11690 (N_11690,N_11091,N_11173);
xor U11691 (N_11691,N_11401,N_11445);
or U11692 (N_11692,N_11294,N_11130);
nor U11693 (N_11693,N_11284,N_11224);
nand U11694 (N_11694,N_11152,N_11495);
xnor U11695 (N_11695,N_11331,N_11400);
xnor U11696 (N_11696,N_11072,N_11403);
nor U11697 (N_11697,N_11256,N_11162);
or U11698 (N_11698,N_11381,N_11372);
nand U11699 (N_11699,N_11471,N_11023);
xnor U11700 (N_11700,N_11320,N_11020);
nand U11701 (N_11701,N_11136,N_11039);
nand U11702 (N_11702,N_11489,N_11121);
or U11703 (N_11703,N_11367,N_11252);
nand U11704 (N_11704,N_11177,N_11248);
nand U11705 (N_11705,N_11417,N_11463);
nand U11706 (N_11706,N_11156,N_11046);
or U11707 (N_11707,N_11222,N_11494);
and U11708 (N_11708,N_11074,N_11008);
or U11709 (N_11709,N_11019,N_11021);
or U11710 (N_11710,N_11423,N_11149);
and U11711 (N_11711,N_11016,N_11188);
nor U11712 (N_11712,N_11449,N_11414);
nor U11713 (N_11713,N_11259,N_11394);
nand U11714 (N_11714,N_11051,N_11133);
xor U11715 (N_11715,N_11373,N_11281);
nand U11716 (N_11716,N_11138,N_11344);
or U11717 (N_11717,N_11316,N_11352);
nand U11718 (N_11718,N_11000,N_11027);
and U11719 (N_11719,N_11024,N_11086);
or U11720 (N_11720,N_11195,N_11325);
nand U11721 (N_11721,N_11424,N_11319);
or U11722 (N_11722,N_11071,N_11359);
or U11723 (N_11723,N_11246,N_11045);
nor U11724 (N_11724,N_11353,N_11369);
and U11725 (N_11725,N_11278,N_11307);
or U11726 (N_11726,N_11184,N_11144);
nand U11727 (N_11727,N_11261,N_11167);
or U11728 (N_11728,N_11277,N_11088);
xnor U11729 (N_11729,N_11260,N_11300);
nand U11730 (N_11730,N_11164,N_11413);
or U11731 (N_11731,N_11070,N_11270);
nor U11732 (N_11732,N_11017,N_11098);
nor U11733 (N_11733,N_11439,N_11383);
nor U11734 (N_11734,N_11393,N_11311);
nor U11735 (N_11735,N_11239,N_11100);
and U11736 (N_11736,N_11408,N_11190);
or U11737 (N_11737,N_11009,N_11497);
xnor U11738 (N_11738,N_11075,N_11336);
nand U11739 (N_11739,N_11061,N_11170);
and U11740 (N_11740,N_11238,N_11237);
xor U11741 (N_11741,N_11377,N_11457);
nor U11742 (N_11742,N_11257,N_11309);
nand U11743 (N_11743,N_11464,N_11409);
and U11744 (N_11744,N_11299,N_11059);
nor U11745 (N_11745,N_11453,N_11485);
nand U11746 (N_11746,N_11154,N_11129);
nand U11747 (N_11747,N_11487,N_11081);
nor U11748 (N_11748,N_11050,N_11153);
nand U11749 (N_11749,N_11398,N_11212);
or U11750 (N_11750,N_11267,N_11313);
or U11751 (N_11751,N_11062,N_11099);
and U11752 (N_11752,N_11120,N_11017);
nor U11753 (N_11753,N_11085,N_11354);
nand U11754 (N_11754,N_11201,N_11316);
xor U11755 (N_11755,N_11001,N_11161);
xnor U11756 (N_11756,N_11437,N_11078);
nor U11757 (N_11757,N_11258,N_11033);
nand U11758 (N_11758,N_11447,N_11394);
xnor U11759 (N_11759,N_11004,N_11447);
xor U11760 (N_11760,N_11171,N_11126);
nor U11761 (N_11761,N_11443,N_11192);
nor U11762 (N_11762,N_11209,N_11048);
nor U11763 (N_11763,N_11246,N_11184);
and U11764 (N_11764,N_11366,N_11222);
nor U11765 (N_11765,N_11156,N_11101);
nand U11766 (N_11766,N_11045,N_11360);
or U11767 (N_11767,N_11039,N_11249);
nor U11768 (N_11768,N_11051,N_11238);
nor U11769 (N_11769,N_11064,N_11350);
nor U11770 (N_11770,N_11279,N_11028);
or U11771 (N_11771,N_11062,N_11452);
or U11772 (N_11772,N_11099,N_11435);
nand U11773 (N_11773,N_11022,N_11185);
and U11774 (N_11774,N_11392,N_11002);
nand U11775 (N_11775,N_11131,N_11411);
nand U11776 (N_11776,N_11262,N_11107);
nand U11777 (N_11777,N_11234,N_11214);
nor U11778 (N_11778,N_11202,N_11412);
xnor U11779 (N_11779,N_11442,N_11184);
nand U11780 (N_11780,N_11100,N_11041);
or U11781 (N_11781,N_11190,N_11029);
or U11782 (N_11782,N_11117,N_11001);
and U11783 (N_11783,N_11036,N_11275);
xor U11784 (N_11784,N_11476,N_11017);
nor U11785 (N_11785,N_11390,N_11413);
and U11786 (N_11786,N_11483,N_11017);
or U11787 (N_11787,N_11165,N_11448);
xor U11788 (N_11788,N_11202,N_11081);
or U11789 (N_11789,N_11423,N_11133);
or U11790 (N_11790,N_11357,N_11038);
nor U11791 (N_11791,N_11094,N_11423);
nand U11792 (N_11792,N_11169,N_11392);
or U11793 (N_11793,N_11269,N_11183);
and U11794 (N_11794,N_11285,N_11325);
nor U11795 (N_11795,N_11281,N_11279);
nand U11796 (N_11796,N_11201,N_11109);
or U11797 (N_11797,N_11107,N_11066);
nand U11798 (N_11798,N_11086,N_11409);
or U11799 (N_11799,N_11303,N_11104);
nor U11800 (N_11800,N_11132,N_11093);
nand U11801 (N_11801,N_11455,N_11448);
or U11802 (N_11802,N_11372,N_11044);
nor U11803 (N_11803,N_11069,N_11409);
and U11804 (N_11804,N_11204,N_11062);
nor U11805 (N_11805,N_11406,N_11175);
nand U11806 (N_11806,N_11111,N_11322);
xnor U11807 (N_11807,N_11423,N_11405);
nand U11808 (N_11808,N_11028,N_11040);
xor U11809 (N_11809,N_11002,N_11109);
and U11810 (N_11810,N_11221,N_11447);
nand U11811 (N_11811,N_11063,N_11196);
nor U11812 (N_11812,N_11289,N_11285);
or U11813 (N_11813,N_11396,N_11005);
nor U11814 (N_11814,N_11139,N_11021);
and U11815 (N_11815,N_11107,N_11208);
xnor U11816 (N_11816,N_11352,N_11484);
xor U11817 (N_11817,N_11488,N_11459);
xor U11818 (N_11818,N_11095,N_11157);
nand U11819 (N_11819,N_11286,N_11358);
and U11820 (N_11820,N_11099,N_11121);
or U11821 (N_11821,N_11143,N_11149);
and U11822 (N_11822,N_11406,N_11333);
or U11823 (N_11823,N_11087,N_11045);
and U11824 (N_11824,N_11301,N_11106);
nor U11825 (N_11825,N_11141,N_11305);
nand U11826 (N_11826,N_11130,N_11110);
nor U11827 (N_11827,N_11034,N_11318);
nand U11828 (N_11828,N_11451,N_11196);
xnor U11829 (N_11829,N_11236,N_11313);
and U11830 (N_11830,N_11234,N_11490);
nand U11831 (N_11831,N_11234,N_11126);
xor U11832 (N_11832,N_11340,N_11259);
xor U11833 (N_11833,N_11487,N_11004);
nand U11834 (N_11834,N_11105,N_11375);
nand U11835 (N_11835,N_11355,N_11477);
or U11836 (N_11836,N_11013,N_11261);
nand U11837 (N_11837,N_11188,N_11449);
nand U11838 (N_11838,N_11260,N_11325);
xnor U11839 (N_11839,N_11334,N_11265);
or U11840 (N_11840,N_11385,N_11074);
xor U11841 (N_11841,N_11313,N_11478);
xor U11842 (N_11842,N_11132,N_11462);
nand U11843 (N_11843,N_11317,N_11101);
nor U11844 (N_11844,N_11283,N_11236);
nand U11845 (N_11845,N_11262,N_11295);
nor U11846 (N_11846,N_11365,N_11228);
xnor U11847 (N_11847,N_11109,N_11304);
or U11848 (N_11848,N_11043,N_11166);
and U11849 (N_11849,N_11499,N_11239);
xor U11850 (N_11850,N_11277,N_11454);
and U11851 (N_11851,N_11352,N_11046);
or U11852 (N_11852,N_11331,N_11384);
nand U11853 (N_11853,N_11166,N_11061);
and U11854 (N_11854,N_11178,N_11241);
xor U11855 (N_11855,N_11465,N_11278);
xor U11856 (N_11856,N_11456,N_11415);
or U11857 (N_11857,N_11034,N_11012);
and U11858 (N_11858,N_11291,N_11239);
xor U11859 (N_11859,N_11142,N_11273);
xor U11860 (N_11860,N_11319,N_11450);
or U11861 (N_11861,N_11115,N_11331);
nor U11862 (N_11862,N_11006,N_11026);
or U11863 (N_11863,N_11119,N_11233);
xor U11864 (N_11864,N_11200,N_11256);
and U11865 (N_11865,N_11096,N_11330);
and U11866 (N_11866,N_11176,N_11012);
xnor U11867 (N_11867,N_11256,N_11059);
nor U11868 (N_11868,N_11234,N_11034);
nand U11869 (N_11869,N_11483,N_11274);
nor U11870 (N_11870,N_11082,N_11173);
and U11871 (N_11871,N_11190,N_11205);
or U11872 (N_11872,N_11469,N_11140);
nand U11873 (N_11873,N_11341,N_11078);
nor U11874 (N_11874,N_11287,N_11175);
xnor U11875 (N_11875,N_11071,N_11395);
nor U11876 (N_11876,N_11128,N_11172);
nand U11877 (N_11877,N_11384,N_11455);
nand U11878 (N_11878,N_11068,N_11438);
or U11879 (N_11879,N_11439,N_11238);
or U11880 (N_11880,N_11250,N_11415);
nand U11881 (N_11881,N_11344,N_11028);
or U11882 (N_11882,N_11204,N_11271);
xor U11883 (N_11883,N_11419,N_11195);
and U11884 (N_11884,N_11230,N_11310);
and U11885 (N_11885,N_11174,N_11486);
nand U11886 (N_11886,N_11141,N_11334);
and U11887 (N_11887,N_11128,N_11197);
xor U11888 (N_11888,N_11274,N_11219);
and U11889 (N_11889,N_11209,N_11413);
and U11890 (N_11890,N_11115,N_11434);
nand U11891 (N_11891,N_11471,N_11088);
nor U11892 (N_11892,N_11242,N_11088);
nand U11893 (N_11893,N_11417,N_11015);
or U11894 (N_11894,N_11053,N_11060);
nor U11895 (N_11895,N_11298,N_11433);
and U11896 (N_11896,N_11156,N_11307);
xor U11897 (N_11897,N_11195,N_11249);
or U11898 (N_11898,N_11050,N_11182);
or U11899 (N_11899,N_11232,N_11330);
nand U11900 (N_11900,N_11226,N_11080);
nand U11901 (N_11901,N_11444,N_11007);
and U11902 (N_11902,N_11188,N_11048);
nor U11903 (N_11903,N_11066,N_11001);
or U11904 (N_11904,N_11172,N_11111);
and U11905 (N_11905,N_11381,N_11309);
and U11906 (N_11906,N_11300,N_11038);
xor U11907 (N_11907,N_11321,N_11457);
xnor U11908 (N_11908,N_11449,N_11485);
nor U11909 (N_11909,N_11096,N_11317);
nor U11910 (N_11910,N_11071,N_11090);
and U11911 (N_11911,N_11360,N_11095);
nor U11912 (N_11912,N_11088,N_11014);
or U11913 (N_11913,N_11407,N_11084);
nor U11914 (N_11914,N_11202,N_11280);
and U11915 (N_11915,N_11103,N_11248);
nand U11916 (N_11916,N_11354,N_11180);
or U11917 (N_11917,N_11072,N_11165);
xor U11918 (N_11918,N_11441,N_11085);
xnor U11919 (N_11919,N_11200,N_11325);
xor U11920 (N_11920,N_11247,N_11105);
xor U11921 (N_11921,N_11475,N_11122);
and U11922 (N_11922,N_11453,N_11415);
and U11923 (N_11923,N_11244,N_11050);
and U11924 (N_11924,N_11295,N_11467);
xor U11925 (N_11925,N_11317,N_11400);
xor U11926 (N_11926,N_11166,N_11102);
or U11927 (N_11927,N_11315,N_11187);
nand U11928 (N_11928,N_11387,N_11477);
xnor U11929 (N_11929,N_11468,N_11484);
and U11930 (N_11930,N_11218,N_11359);
xor U11931 (N_11931,N_11149,N_11014);
nor U11932 (N_11932,N_11256,N_11051);
or U11933 (N_11933,N_11081,N_11481);
nand U11934 (N_11934,N_11089,N_11013);
and U11935 (N_11935,N_11372,N_11377);
xnor U11936 (N_11936,N_11098,N_11316);
xnor U11937 (N_11937,N_11051,N_11307);
xor U11938 (N_11938,N_11192,N_11370);
xor U11939 (N_11939,N_11333,N_11124);
nor U11940 (N_11940,N_11458,N_11409);
or U11941 (N_11941,N_11075,N_11376);
nor U11942 (N_11942,N_11414,N_11462);
and U11943 (N_11943,N_11367,N_11184);
nand U11944 (N_11944,N_11464,N_11037);
nor U11945 (N_11945,N_11381,N_11399);
nor U11946 (N_11946,N_11404,N_11402);
or U11947 (N_11947,N_11140,N_11123);
xor U11948 (N_11948,N_11494,N_11389);
nor U11949 (N_11949,N_11254,N_11202);
nor U11950 (N_11950,N_11202,N_11120);
nor U11951 (N_11951,N_11356,N_11357);
or U11952 (N_11952,N_11169,N_11076);
or U11953 (N_11953,N_11171,N_11389);
or U11954 (N_11954,N_11337,N_11204);
and U11955 (N_11955,N_11449,N_11381);
xnor U11956 (N_11956,N_11458,N_11333);
xnor U11957 (N_11957,N_11023,N_11357);
or U11958 (N_11958,N_11499,N_11218);
nand U11959 (N_11959,N_11221,N_11496);
xor U11960 (N_11960,N_11438,N_11003);
nand U11961 (N_11961,N_11258,N_11473);
or U11962 (N_11962,N_11371,N_11112);
nand U11963 (N_11963,N_11080,N_11359);
xor U11964 (N_11964,N_11449,N_11104);
nor U11965 (N_11965,N_11145,N_11318);
nor U11966 (N_11966,N_11278,N_11071);
xor U11967 (N_11967,N_11277,N_11094);
and U11968 (N_11968,N_11015,N_11458);
and U11969 (N_11969,N_11433,N_11475);
xnor U11970 (N_11970,N_11397,N_11041);
and U11971 (N_11971,N_11324,N_11284);
xor U11972 (N_11972,N_11486,N_11044);
or U11973 (N_11973,N_11258,N_11177);
nand U11974 (N_11974,N_11376,N_11348);
and U11975 (N_11975,N_11123,N_11483);
xor U11976 (N_11976,N_11203,N_11326);
and U11977 (N_11977,N_11236,N_11480);
or U11978 (N_11978,N_11484,N_11333);
nor U11979 (N_11979,N_11259,N_11226);
or U11980 (N_11980,N_11282,N_11251);
or U11981 (N_11981,N_11492,N_11225);
and U11982 (N_11982,N_11372,N_11272);
nand U11983 (N_11983,N_11135,N_11252);
nand U11984 (N_11984,N_11106,N_11188);
or U11985 (N_11985,N_11004,N_11251);
xnor U11986 (N_11986,N_11292,N_11262);
nand U11987 (N_11987,N_11474,N_11398);
xor U11988 (N_11988,N_11186,N_11484);
nand U11989 (N_11989,N_11327,N_11468);
nor U11990 (N_11990,N_11231,N_11369);
nand U11991 (N_11991,N_11210,N_11235);
or U11992 (N_11992,N_11221,N_11172);
xnor U11993 (N_11993,N_11104,N_11099);
nor U11994 (N_11994,N_11163,N_11475);
nor U11995 (N_11995,N_11226,N_11144);
and U11996 (N_11996,N_11011,N_11040);
and U11997 (N_11997,N_11470,N_11412);
and U11998 (N_11998,N_11311,N_11142);
and U11999 (N_11999,N_11034,N_11100);
nor U12000 (N_12000,N_11514,N_11830);
nand U12001 (N_12001,N_11528,N_11766);
and U12002 (N_12002,N_11535,N_11936);
nor U12003 (N_12003,N_11629,N_11961);
and U12004 (N_12004,N_11713,N_11626);
or U12005 (N_12005,N_11693,N_11703);
or U12006 (N_12006,N_11988,N_11680);
xor U12007 (N_12007,N_11771,N_11633);
xor U12008 (N_12008,N_11933,N_11710);
xor U12009 (N_12009,N_11920,N_11530);
or U12010 (N_12010,N_11863,N_11947);
nand U12011 (N_12011,N_11910,N_11704);
nor U12012 (N_12012,N_11675,N_11513);
and U12013 (N_12013,N_11751,N_11511);
xor U12014 (N_12014,N_11662,N_11873);
nand U12015 (N_12015,N_11911,N_11974);
or U12016 (N_12016,N_11568,N_11864);
nand U12017 (N_12017,N_11869,N_11534);
xor U12018 (N_12018,N_11912,N_11652);
or U12019 (N_12019,N_11828,N_11654);
nor U12020 (N_12020,N_11667,N_11931);
and U12021 (N_12021,N_11708,N_11905);
xor U12022 (N_12022,N_11990,N_11915);
nand U12023 (N_12023,N_11749,N_11850);
nor U12024 (N_12024,N_11757,N_11849);
and U12025 (N_12025,N_11590,N_11997);
and U12026 (N_12026,N_11764,N_11950);
nor U12027 (N_12027,N_11999,N_11502);
nand U12028 (N_12028,N_11759,N_11963);
nor U12029 (N_12029,N_11921,N_11670);
or U12030 (N_12030,N_11983,N_11519);
nor U12031 (N_12031,N_11781,N_11734);
nor U12032 (N_12032,N_11518,N_11929);
xor U12033 (N_12033,N_11743,N_11982);
nor U12034 (N_12034,N_11733,N_11688);
nand U12035 (N_12035,N_11878,N_11524);
or U12036 (N_12036,N_11602,N_11934);
or U12037 (N_12037,N_11575,N_11976);
xnor U12038 (N_12038,N_11701,N_11539);
and U12039 (N_12039,N_11711,N_11672);
or U12040 (N_12040,N_11817,N_11532);
nor U12041 (N_12041,N_11541,N_11943);
xor U12042 (N_12042,N_11612,N_11619);
nand U12043 (N_12043,N_11698,N_11940);
nand U12044 (N_12044,N_11526,N_11861);
xnor U12045 (N_12045,N_11832,N_11696);
xnor U12046 (N_12046,N_11617,N_11560);
and U12047 (N_12047,N_11607,N_11674);
nor U12048 (N_12048,N_11635,N_11648);
nor U12049 (N_12049,N_11977,N_11777);
nand U12050 (N_12050,N_11702,N_11706);
and U12051 (N_12051,N_11538,N_11883);
xor U12052 (N_12052,N_11681,N_11577);
nor U12053 (N_12053,N_11664,N_11862);
nand U12054 (N_12054,N_11797,N_11896);
and U12055 (N_12055,N_11956,N_11650);
xor U12056 (N_12056,N_11782,N_11826);
xnor U12057 (N_12057,N_11601,N_11754);
nand U12058 (N_12058,N_11952,N_11813);
nor U12059 (N_12059,N_11755,N_11770);
nand U12060 (N_12060,N_11835,N_11890);
xnor U12061 (N_12061,N_11622,N_11747);
or U12062 (N_12062,N_11882,N_11647);
nor U12063 (N_12063,N_11914,N_11948);
nand U12064 (N_12064,N_11840,N_11899);
xnor U12065 (N_12065,N_11721,N_11561);
xor U12066 (N_12066,N_11957,N_11837);
or U12067 (N_12067,N_11859,N_11520);
xor U12068 (N_12068,N_11968,N_11897);
or U12069 (N_12069,N_11555,N_11892);
nor U12070 (N_12070,N_11844,N_11776);
and U12071 (N_12071,N_11671,N_11705);
nand U12072 (N_12072,N_11803,N_11768);
or U12073 (N_12073,N_11825,N_11984);
nor U12074 (N_12074,N_11854,N_11877);
xnor U12075 (N_12075,N_11725,N_11669);
nor U12076 (N_12076,N_11769,N_11506);
nand U12077 (N_12077,N_11636,N_11603);
xnor U12078 (N_12078,N_11531,N_11529);
and U12079 (N_12079,N_11658,N_11549);
nor U12080 (N_12080,N_11596,N_11762);
or U12081 (N_12081,N_11512,N_11536);
xnor U12082 (N_12082,N_11924,N_11595);
and U12083 (N_12083,N_11913,N_11690);
nor U12084 (N_12084,N_11614,N_11919);
nor U12085 (N_12085,N_11966,N_11935);
nor U12086 (N_12086,N_11951,N_11611);
xnor U12087 (N_12087,N_11904,N_11683);
or U12088 (N_12088,N_11620,N_11716);
xnor U12089 (N_12089,N_11673,N_11839);
nor U12090 (N_12090,N_11730,N_11889);
and U12091 (N_12091,N_11756,N_11739);
and U12092 (N_12092,N_11738,N_11876);
nand U12093 (N_12093,N_11820,N_11867);
nand U12094 (N_12094,N_11745,N_11744);
xor U12095 (N_12095,N_11939,N_11763);
and U12096 (N_12096,N_11548,N_11623);
nand U12097 (N_12097,N_11656,N_11558);
or U12098 (N_12098,N_11898,N_11509);
xnor U12099 (N_12099,N_11804,N_11679);
xor U12100 (N_12100,N_11556,N_11836);
or U12101 (N_12101,N_11578,N_11818);
xnor U12102 (N_12102,N_11563,N_11846);
or U12103 (N_12103,N_11774,N_11576);
nand U12104 (N_12104,N_11608,N_11564);
nand U12105 (N_12105,N_11712,N_11908);
and U12106 (N_12106,N_11980,N_11923);
nand U12107 (N_12107,N_11857,N_11613);
nand U12108 (N_12108,N_11579,N_11917);
xnor U12109 (N_12109,N_11599,N_11634);
or U12110 (N_12110,N_11586,N_11895);
nand U12111 (N_12111,N_11510,N_11565);
nand U12112 (N_12112,N_11885,N_11969);
nand U12113 (N_12113,N_11942,N_11790);
or U12114 (N_12114,N_11870,N_11842);
xnor U12115 (N_12115,N_11545,N_11573);
or U12116 (N_12116,N_11838,N_11814);
nor U12117 (N_12117,N_11587,N_11525);
xor U12118 (N_12118,N_11752,N_11845);
nor U12119 (N_12119,N_11993,N_11802);
xnor U12120 (N_12120,N_11597,N_11979);
and U12121 (N_12121,N_11808,N_11925);
or U12122 (N_12122,N_11559,N_11659);
nor U12123 (N_12123,N_11843,N_11954);
or U12124 (N_12124,N_11801,N_11799);
nand U12125 (N_12125,N_11784,N_11624);
nand U12126 (N_12126,N_11741,N_11780);
nand U12127 (N_12127,N_11959,N_11930);
nand U12128 (N_12128,N_11909,N_11775);
nor U12129 (N_12129,N_11550,N_11894);
and U12130 (N_12130,N_11717,N_11593);
or U12131 (N_12131,N_11588,N_11697);
xor U12132 (N_12132,N_11687,N_11724);
nor U12133 (N_12133,N_11748,N_11865);
xnor U12134 (N_12134,N_11750,N_11886);
and U12135 (N_12135,N_11821,N_11589);
nand U12136 (N_12136,N_11727,N_11643);
and U12137 (N_12137,N_11855,N_11900);
nand U12138 (N_12138,N_11812,N_11958);
or U12139 (N_12139,N_11848,N_11884);
nor U12140 (N_12140,N_11965,N_11584);
and U12141 (N_12141,N_11552,N_11960);
nand U12142 (N_12142,N_11605,N_11783);
xnor U12143 (N_12143,N_11786,N_11973);
nand U12144 (N_12144,N_11872,N_11606);
xnor U12145 (N_12145,N_11718,N_11938);
and U12146 (N_12146,N_11628,N_11932);
or U12147 (N_12147,N_11574,N_11926);
or U12148 (N_12148,N_11753,N_11946);
and U12149 (N_12149,N_11789,N_11823);
and U12150 (N_12150,N_11767,N_11728);
nand U12151 (N_12151,N_11798,N_11971);
xnor U12152 (N_12152,N_11665,N_11742);
nor U12153 (N_12153,N_11554,N_11795);
nand U12154 (N_12154,N_11815,N_11682);
xor U12155 (N_12155,N_11995,N_11949);
xor U12156 (N_12156,N_11507,N_11642);
xnor U12157 (N_12157,N_11737,N_11686);
or U12158 (N_12158,N_11962,N_11685);
or U12159 (N_12159,N_11772,N_11691);
and U12160 (N_12160,N_11726,N_11785);
nand U12161 (N_12161,N_11707,N_11794);
and U12162 (N_12162,N_11805,N_11879);
xor U12163 (N_12163,N_11720,N_11736);
nor U12164 (N_12164,N_11562,N_11591);
xnor U12165 (N_12165,N_11874,N_11981);
nor U12166 (N_12166,N_11632,N_11907);
nor U12167 (N_12167,N_11505,N_11918);
or U12168 (N_12168,N_11553,N_11880);
nor U12169 (N_12169,N_11645,N_11996);
xnor U12170 (N_12170,N_11504,N_11592);
nand U12171 (N_12171,N_11501,N_11941);
nor U12172 (N_12172,N_11903,N_11699);
nand U12173 (N_12173,N_11523,N_11991);
nor U12174 (N_12174,N_11955,N_11819);
nand U12175 (N_12175,N_11594,N_11809);
or U12176 (N_12176,N_11779,N_11975);
nor U12177 (N_12177,N_11668,N_11807);
or U12178 (N_12178,N_11871,N_11722);
and U12179 (N_12179,N_11902,N_11834);
or U12180 (N_12180,N_11901,N_11922);
nand U12181 (N_12181,N_11989,N_11700);
nand U12182 (N_12182,N_11663,N_11551);
xor U12183 (N_12183,N_11853,N_11831);
xnor U12184 (N_12184,N_11661,N_11928);
and U12185 (N_12185,N_11994,N_11967);
and U12186 (N_12186,N_11972,N_11657);
or U12187 (N_12187,N_11638,N_11944);
xor U12188 (N_12188,N_11824,N_11816);
nand U12189 (N_12189,N_11793,N_11806);
or U12190 (N_12190,N_11740,N_11945);
nand U12191 (N_12191,N_11694,N_11598);
and U12192 (N_12192,N_11765,N_11860);
xor U12193 (N_12193,N_11609,N_11571);
and U12194 (N_12194,N_11787,N_11858);
nor U12195 (N_12195,N_11600,N_11585);
xor U12196 (N_12196,N_11649,N_11500);
and U12197 (N_12197,N_11646,N_11856);
xor U12198 (N_12198,N_11875,N_11758);
and U12199 (N_12199,N_11630,N_11676);
nor U12200 (N_12200,N_11540,N_11572);
and U12201 (N_12201,N_11678,N_11732);
and U12202 (N_12202,N_11615,N_11543);
nor U12203 (N_12203,N_11618,N_11508);
and U12204 (N_12204,N_11810,N_11731);
and U12205 (N_12205,N_11714,N_11978);
or U12206 (N_12206,N_11841,N_11517);
and U12207 (N_12207,N_11621,N_11527);
and U12208 (N_12208,N_11964,N_11723);
or U12209 (N_12209,N_11887,N_11761);
or U12210 (N_12210,N_11522,N_11610);
xnor U12211 (N_12211,N_11569,N_11891);
nor U12212 (N_12212,N_11760,N_11537);
or U12213 (N_12213,N_11637,N_11677);
nand U12214 (N_12214,N_11625,N_11970);
xor U12215 (N_12215,N_11616,N_11986);
nor U12216 (N_12216,N_11644,N_11515);
nand U12217 (N_12217,N_11833,N_11692);
or U12218 (N_12218,N_11778,N_11811);
nand U12219 (N_12219,N_11533,N_11655);
and U12220 (N_12220,N_11746,N_11985);
or U12221 (N_12221,N_11916,N_11544);
and U12222 (N_12222,N_11829,N_11992);
and U12223 (N_12223,N_11640,N_11666);
xor U12224 (N_12224,N_11639,N_11791);
nor U12225 (N_12225,N_11684,N_11888);
nand U12226 (N_12226,N_11581,N_11660);
and U12227 (N_12227,N_11566,N_11719);
nor U12228 (N_12228,N_11580,N_11852);
nor U12229 (N_12229,N_11827,N_11631);
xnor U12230 (N_12230,N_11792,N_11735);
xnor U12231 (N_12231,N_11953,N_11557);
xor U12232 (N_12232,N_11773,N_11604);
xnor U12233 (N_12233,N_11570,N_11800);
xor U12234 (N_12234,N_11868,N_11516);
and U12235 (N_12235,N_11546,N_11822);
xnor U12236 (N_12236,N_11542,N_11893);
nor U12237 (N_12237,N_11851,N_11641);
nor U12238 (N_12238,N_11583,N_11847);
nor U12239 (N_12239,N_11503,N_11906);
and U12240 (N_12240,N_11715,N_11987);
xor U12241 (N_12241,N_11881,N_11689);
and U12242 (N_12242,N_11521,N_11651);
nand U12243 (N_12243,N_11866,N_11937);
nor U12244 (N_12244,N_11653,N_11547);
or U12245 (N_12245,N_11695,N_11788);
nand U12246 (N_12246,N_11709,N_11998);
xnor U12247 (N_12247,N_11567,N_11796);
or U12248 (N_12248,N_11927,N_11582);
xor U12249 (N_12249,N_11729,N_11627);
or U12250 (N_12250,N_11985,N_11966);
xnor U12251 (N_12251,N_11836,N_11536);
and U12252 (N_12252,N_11586,N_11814);
or U12253 (N_12253,N_11801,N_11713);
and U12254 (N_12254,N_11575,N_11665);
or U12255 (N_12255,N_11753,N_11720);
xnor U12256 (N_12256,N_11640,N_11628);
and U12257 (N_12257,N_11836,N_11811);
nand U12258 (N_12258,N_11516,N_11562);
xor U12259 (N_12259,N_11903,N_11559);
nor U12260 (N_12260,N_11523,N_11829);
nand U12261 (N_12261,N_11564,N_11937);
xnor U12262 (N_12262,N_11833,N_11874);
xor U12263 (N_12263,N_11592,N_11880);
and U12264 (N_12264,N_11830,N_11524);
or U12265 (N_12265,N_11636,N_11645);
xor U12266 (N_12266,N_11772,N_11670);
nor U12267 (N_12267,N_11592,N_11633);
nor U12268 (N_12268,N_11642,N_11898);
nor U12269 (N_12269,N_11962,N_11828);
and U12270 (N_12270,N_11741,N_11622);
nand U12271 (N_12271,N_11910,N_11756);
xnor U12272 (N_12272,N_11900,N_11752);
or U12273 (N_12273,N_11930,N_11908);
and U12274 (N_12274,N_11739,N_11557);
nand U12275 (N_12275,N_11739,N_11707);
xnor U12276 (N_12276,N_11975,N_11696);
or U12277 (N_12277,N_11774,N_11819);
xnor U12278 (N_12278,N_11982,N_11749);
xnor U12279 (N_12279,N_11772,N_11537);
and U12280 (N_12280,N_11886,N_11837);
or U12281 (N_12281,N_11847,N_11759);
or U12282 (N_12282,N_11908,N_11831);
nand U12283 (N_12283,N_11952,N_11520);
nand U12284 (N_12284,N_11955,N_11587);
or U12285 (N_12285,N_11774,N_11740);
xnor U12286 (N_12286,N_11772,N_11880);
and U12287 (N_12287,N_11939,N_11648);
nand U12288 (N_12288,N_11824,N_11897);
nand U12289 (N_12289,N_11675,N_11707);
nand U12290 (N_12290,N_11824,N_11711);
nor U12291 (N_12291,N_11964,N_11642);
nand U12292 (N_12292,N_11783,N_11520);
and U12293 (N_12293,N_11558,N_11799);
nand U12294 (N_12294,N_11842,N_11633);
nor U12295 (N_12295,N_11536,N_11743);
xor U12296 (N_12296,N_11769,N_11562);
nor U12297 (N_12297,N_11547,N_11941);
or U12298 (N_12298,N_11734,N_11733);
nor U12299 (N_12299,N_11956,N_11680);
nand U12300 (N_12300,N_11669,N_11537);
and U12301 (N_12301,N_11665,N_11529);
xor U12302 (N_12302,N_11934,N_11788);
and U12303 (N_12303,N_11971,N_11786);
xnor U12304 (N_12304,N_11573,N_11527);
xor U12305 (N_12305,N_11683,N_11942);
xor U12306 (N_12306,N_11856,N_11879);
xor U12307 (N_12307,N_11983,N_11798);
nand U12308 (N_12308,N_11931,N_11549);
or U12309 (N_12309,N_11578,N_11934);
and U12310 (N_12310,N_11518,N_11509);
xnor U12311 (N_12311,N_11762,N_11648);
nor U12312 (N_12312,N_11593,N_11791);
nor U12313 (N_12313,N_11940,N_11980);
xnor U12314 (N_12314,N_11573,N_11630);
nor U12315 (N_12315,N_11851,N_11776);
nand U12316 (N_12316,N_11929,N_11571);
xnor U12317 (N_12317,N_11697,N_11894);
xor U12318 (N_12318,N_11758,N_11940);
or U12319 (N_12319,N_11692,N_11936);
nor U12320 (N_12320,N_11775,N_11656);
nor U12321 (N_12321,N_11809,N_11651);
xor U12322 (N_12322,N_11567,N_11600);
and U12323 (N_12323,N_11710,N_11749);
or U12324 (N_12324,N_11980,N_11583);
or U12325 (N_12325,N_11666,N_11900);
xnor U12326 (N_12326,N_11690,N_11570);
nand U12327 (N_12327,N_11969,N_11740);
and U12328 (N_12328,N_11681,N_11904);
xor U12329 (N_12329,N_11657,N_11599);
nand U12330 (N_12330,N_11836,N_11614);
or U12331 (N_12331,N_11970,N_11504);
xnor U12332 (N_12332,N_11570,N_11803);
and U12333 (N_12333,N_11850,N_11644);
or U12334 (N_12334,N_11522,N_11573);
nand U12335 (N_12335,N_11509,N_11511);
or U12336 (N_12336,N_11876,N_11533);
and U12337 (N_12337,N_11549,N_11935);
nand U12338 (N_12338,N_11567,N_11642);
or U12339 (N_12339,N_11958,N_11762);
or U12340 (N_12340,N_11720,N_11890);
xor U12341 (N_12341,N_11667,N_11900);
nor U12342 (N_12342,N_11505,N_11936);
or U12343 (N_12343,N_11740,N_11791);
nor U12344 (N_12344,N_11832,N_11685);
or U12345 (N_12345,N_11553,N_11971);
xor U12346 (N_12346,N_11840,N_11748);
and U12347 (N_12347,N_11891,N_11733);
or U12348 (N_12348,N_11573,N_11640);
nor U12349 (N_12349,N_11750,N_11829);
nand U12350 (N_12350,N_11561,N_11749);
nor U12351 (N_12351,N_11886,N_11859);
or U12352 (N_12352,N_11994,N_11691);
nand U12353 (N_12353,N_11583,N_11567);
nand U12354 (N_12354,N_11839,N_11593);
xnor U12355 (N_12355,N_11980,N_11774);
nor U12356 (N_12356,N_11749,N_11879);
and U12357 (N_12357,N_11537,N_11514);
nor U12358 (N_12358,N_11621,N_11927);
and U12359 (N_12359,N_11745,N_11962);
nor U12360 (N_12360,N_11506,N_11528);
nand U12361 (N_12361,N_11846,N_11930);
or U12362 (N_12362,N_11692,N_11818);
nor U12363 (N_12363,N_11917,N_11954);
nand U12364 (N_12364,N_11695,N_11588);
nor U12365 (N_12365,N_11576,N_11843);
or U12366 (N_12366,N_11572,N_11993);
or U12367 (N_12367,N_11870,N_11882);
xor U12368 (N_12368,N_11584,N_11862);
and U12369 (N_12369,N_11973,N_11675);
and U12370 (N_12370,N_11514,N_11515);
nor U12371 (N_12371,N_11535,N_11765);
or U12372 (N_12372,N_11644,N_11953);
and U12373 (N_12373,N_11819,N_11803);
or U12374 (N_12374,N_11918,N_11876);
or U12375 (N_12375,N_11756,N_11992);
or U12376 (N_12376,N_11958,N_11830);
nor U12377 (N_12377,N_11668,N_11835);
nand U12378 (N_12378,N_11887,N_11603);
nand U12379 (N_12379,N_11770,N_11815);
and U12380 (N_12380,N_11682,N_11645);
xnor U12381 (N_12381,N_11900,N_11698);
nand U12382 (N_12382,N_11921,N_11566);
and U12383 (N_12383,N_11505,N_11828);
or U12384 (N_12384,N_11936,N_11639);
and U12385 (N_12385,N_11961,N_11934);
and U12386 (N_12386,N_11974,N_11918);
nor U12387 (N_12387,N_11655,N_11885);
nand U12388 (N_12388,N_11938,N_11725);
or U12389 (N_12389,N_11966,N_11934);
nor U12390 (N_12390,N_11823,N_11676);
nor U12391 (N_12391,N_11896,N_11730);
nand U12392 (N_12392,N_11643,N_11736);
xnor U12393 (N_12393,N_11858,N_11553);
and U12394 (N_12394,N_11580,N_11988);
or U12395 (N_12395,N_11747,N_11609);
or U12396 (N_12396,N_11614,N_11832);
nand U12397 (N_12397,N_11541,N_11950);
nor U12398 (N_12398,N_11658,N_11613);
or U12399 (N_12399,N_11587,N_11514);
xor U12400 (N_12400,N_11902,N_11964);
nor U12401 (N_12401,N_11620,N_11606);
nor U12402 (N_12402,N_11751,N_11608);
nand U12403 (N_12403,N_11865,N_11555);
nor U12404 (N_12404,N_11967,N_11972);
and U12405 (N_12405,N_11982,N_11606);
nor U12406 (N_12406,N_11672,N_11980);
nor U12407 (N_12407,N_11635,N_11661);
or U12408 (N_12408,N_11823,N_11785);
nand U12409 (N_12409,N_11604,N_11862);
or U12410 (N_12410,N_11804,N_11503);
nand U12411 (N_12411,N_11774,N_11699);
nor U12412 (N_12412,N_11648,N_11510);
or U12413 (N_12413,N_11898,N_11779);
xnor U12414 (N_12414,N_11534,N_11966);
nand U12415 (N_12415,N_11604,N_11810);
nand U12416 (N_12416,N_11621,N_11799);
and U12417 (N_12417,N_11825,N_11510);
and U12418 (N_12418,N_11872,N_11732);
and U12419 (N_12419,N_11797,N_11926);
nor U12420 (N_12420,N_11822,N_11508);
xnor U12421 (N_12421,N_11962,N_11865);
nor U12422 (N_12422,N_11781,N_11974);
nor U12423 (N_12423,N_11538,N_11791);
and U12424 (N_12424,N_11890,N_11921);
xnor U12425 (N_12425,N_11893,N_11825);
nor U12426 (N_12426,N_11619,N_11526);
nor U12427 (N_12427,N_11902,N_11753);
xnor U12428 (N_12428,N_11880,N_11652);
and U12429 (N_12429,N_11758,N_11613);
xor U12430 (N_12430,N_11737,N_11675);
nor U12431 (N_12431,N_11710,N_11551);
xnor U12432 (N_12432,N_11716,N_11547);
xor U12433 (N_12433,N_11646,N_11785);
xnor U12434 (N_12434,N_11870,N_11928);
and U12435 (N_12435,N_11798,N_11911);
xnor U12436 (N_12436,N_11556,N_11613);
and U12437 (N_12437,N_11920,N_11521);
nand U12438 (N_12438,N_11550,N_11614);
or U12439 (N_12439,N_11730,N_11553);
and U12440 (N_12440,N_11810,N_11631);
nand U12441 (N_12441,N_11734,N_11732);
xnor U12442 (N_12442,N_11602,N_11790);
nor U12443 (N_12443,N_11783,N_11905);
or U12444 (N_12444,N_11932,N_11945);
xor U12445 (N_12445,N_11884,N_11604);
nand U12446 (N_12446,N_11972,N_11715);
nand U12447 (N_12447,N_11805,N_11803);
nor U12448 (N_12448,N_11937,N_11568);
nor U12449 (N_12449,N_11611,N_11832);
and U12450 (N_12450,N_11655,N_11870);
or U12451 (N_12451,N_11897,N_11637);
or U12452 (N_12452,N_11706,N_11619);
nor U12453 (N_12453,N_11782,N_11849);
nor U12454 (N_12454,N_11909,N_11780);
nand U12455 (N_12455,N_11552,N_11711);
nor U12456 (N_12456,N_11871,N_11665);
and U12457 (N_12457,N_11545,N_11751);
xnor U12458 (N_12458,N_11542,N_11732);
or U12459 (N_12459,N_11947,N_11995);
nor U12460 (N_12460,N_11914,N_11611);
and U12461 (N_12461,N_11872,N_11838);
and U12462 (N_12462,N_11949,N_11826);
nand U12463 (N_12463,N_11546,N_11541);
nand U12464 (N_12464,N_11685,N_11913);
or U12465 (N_12465,N_11648,N_11846);
and U12466 (N_12466,N_11506,N_11982);
xor U12467 (N_12467,N_11557,N_11938);
nand U12468 (N_12468,N_11597,N_11908);
nor U12469 (N_12469,N_11619,N_11871);
nor U12470 (N_12470,N_11828,N_11615);
xnor U12471 (N_12471,N_11869,N_11934);
and U12472 (N_12472,N_11544,N_11996);
and U12473 (N_12473,N_11616,N_11620);
nand U12474 (N_12474,N_11745,N_11736);
nor U12475 (N_12475,N_11515,N_11592);
nor U12476 (N_12476,N_11989,N_11795);
xor U12477 (N_12477,N_11783,N_11925);
nand U12478 (N_12478,N_11608,N_11923);
nor U12479 (N_12479,N_11724,N_11942);
and U12480 (N_12480,N_11903,N_11782);
nor U12481 (N_12481,N_11722,N_11674);
and U12482 (N_12482,N_11588,N_11971);
nor U12483 (N_12483,N_11836,N_11537);
nor U12484 (N_12484,N_11985,N_11789);
xor U12485 (N_12485,N_11742,N_11932);
xnor U12486 (N_12486,N_11974,N_11695);
or U12487 (N_12487,N_11688,N_11560);
nand U12488 (N_12488,N_11823,N_11623);
or U12489 (N_12489,N_11554,N_11659);
nand U12490 (N_12490,N_11725,N_11862);
nor U12491 (N_12491,N_11801,N_11997);
nor U12492 (N_12492,N_11984,N_11781);
nand U12493 (N_12493,N_11894,N_11932);
or U12494 (N_12494,N_11990,N_11505);
nor U12495 (N_12495,N_11793,N_11612);
xnor U12496 (N_12496,N_11876,N_11689);
nor U12497 (N_12497,N_11866,N_11608);
xnor U12498 (N_12498,N_11590,N_11895);
nand U12499 (N_12499,N_11886,N_11935);
or U12500 (N_12500,N_12459,N_12281);
xnor U12501 (N_12501,N_12127,N_12255);
or U12502 (N_12502,N_12138,N_12365);
or U12503 (N_12503,N_12376,N_12322);
nand U12504 (N_12504,N_12337,N_12286);
xnor U12505 (N_12505,N_12397,N_12387);
or U12506 (N_12506,N_12406,N_12317);
nor U12507 (N_12507,N_12001,N_12458);
and U12508 (N_12508,N_12282,N_12124);
and U12509 (N_12509,N_12071,N_12269);
nand U12510 (N_12510,N_12099,N_12457);
and U12511 (N_12511,N_12130,N_12328);
nor U12512 (N_12512,N_12123,N_12232);
nand U12513 (N_12513,N_12155,N_12113);
xnor U12514 (N_12514,N_12145,N_12329);
nor U12515 (N_12515,N_12167,N_12366);
xnor U12516 (N_12516,N_12093,N_12343);
or U12517 (N_12517,N_12469,N_12222);
nand U12518 (N_12518,N_12190,N_12098);
or U12519 (N_12519,N_12035,N_12235);
nand U12520 (N_12520,N_12416,N_12236);
or U12521 (N_12521,N_12291,N_12132);
xnor U12522 (N_12522,N_12298,N_12120);
and U12523 (N_12523,N_12193,N_12492);
xnor U12524 (N_12524,N_12196,N_12181);
nand U12525 (N_12525,N_12010,N_12108);
or U12526 (N_12526,N_12392,N_12074);
xor U12527 (N_12527,N_12359,N_12103);
or U12528 (N_12528,N_12191,N_12162);
nand U12529 (N_12529,N_12425,N_12465);
nand U12530 (N_12530,N_12381,N_12379);
or U12531 (N_12531,N_12067,N_12385);
or U12532 (N_12532,N_12079,N_12351);
and U12533 (N_12533,N_12426,N_12302);
nor U12534 (N_12534,N_12441,N_12306);
and U12535 (N_12535,N_12195,N_12354);
or U12536 (N_12536,N_12046,N_12148);
and U12537 (N_12537,N_12154,N_12070);
nand U12538 (N_12538,N_12021,N_12263);
nor U12539 (N_12539,N_12331,N_12065);
xor U12540 (N_12540,N_12445,N_12198);
nor U12541 (N_12541,N_12422,N_12128);
nand U12542 (N_12542,N_12361,N_12234);
or U12543 (N_12543,N_12399,N_12184);
nand U12544 (N_12544,N_12327,N_12086);
and U12545 (N_12545,N_12452,N_12491);
or U12546 (N_12546,N_12000,N_12407);
nor U12547 (N_12547,N_12477,N_12319);
nor U12548 (N_12548,N_12131,N_12034);
nor U12549 (N_12549,N_12398,N_12052);
xor U12550 (N_12550,N_12402,N_12220);
nand U12551 (N_12551,N_12212,N_12495);
nor U12552 (N_12552,N_12428,N_12077);
nor U12553 (N_12553,N_12178,N_12369);
nand U12554 (N_12554,N_12166,N_12434);
xnor U12555 (N_12555,N_12456,N_12216);
xnor U12556 (N_12556,N_12016,N_12436);
xnor U12557 (N_12557,N_12481,N_12227);
and U12558 (N_12558,N_12279,N_12403);
nor U12559 (N_12559,N_12210,N_12423);
xor U12560 (N_12560,N_12174,N_12028);
xnor U12561 (N_12561,N_12064,N_12454);
and U12562 (N_12562,N_12400,N_12483);
or U12563 (N_12563,N_12047,N_12151);
and U12564 (N_12564,N_12371,N_12228);
xor U12565 (N_12565,N_12041,N_12304);
and U12566 (N_12566,N_12325,N_12499);
or U12567 (N_12567,N_12299,N_12150);
and U12568 (N_12568,N_12200,N_12078);
nor U12569 (N_12569,N_12036,N_12039);
nand U12570 (N_12570,N_12069,N_12002);
nor U12571 (N_12571,N_12223,N_12006);
nand U12572 (N_12572,N_12187,N_12336);
or U12573 (N_12573,N_12380,N_12312);
and U12574 (N_12574,N_12126,N_12346);
or U12575 (N_12575,N_12262,N_12109);
or U12576 (N_12576,N_12122,N_12453);
xnor U12577 (N_12577,N_12350,N_12107);
nand U12578 (N_12578,N_12294,N_12023);
nor U12579 (N_12579,N_12231,N_12146);
nand U12580 (N_12580,N_12247,N_12498);
nor U12581 (N_12581,N_12244,N_12118);
xor U12582 (N_12582,N_12180,N_12242);
or U12583 (N_12583,N_12240,N_12153);
and U12584 (N_12584,N_12476,N_12435);
nand U12585 (N_12585,N_12163,N_12374);
or U12586 (N_12586,N_12060,N_12049);
nor U12587 (N_12587,N_12179,N_12221);
nor U12588 (N_12588,N_12037,N_12288);
and U12589 (N_12589,N_12159,N_12011);
xor U12590 (N_12590,N_12097,N_12012);
and U12591 (N_12591,N_12349,N_12061);
nand U12592 (N_12592,N_12233,N_12280);
nor U12593 (N_12593,N_12117,N_12348);
and U12594 (N_12594,N_12413,N_12264);
xor U12595 (N_12595,N_12488,N_12363);
nand U12596 (N_12596,N_12217,N_12250);
xnor U12597 (N_12597,N_12185,N_12278);
and U12598 (N_12598,N_12014,N_12192);
and U12599 (N_12599,N_12142,N_12352);
xnor U12600 (N_12600,N_12063,N_12489);
and U12601 (N_12601,N_12214,N_12496);
nand U12602 (N_12602,N_12472,N_12115);
or U12603 (N_12603,N_12493,N_12292);
nor U12604 (N_12604,N_12438,N_12333);
or U12605 (N_12605,N_12075,N_12475);
and U12606 (N_12606,N_12055,N_12275);
and U12607 (N_12607,N_12451,N_12135);
xor U12608 (N_12608,N_12090,N_12321);
nor U12609 (N_12609,N_12168,N_12199);
nor U12610 (N_12610,N_12054,N_12252);
and U12611 (N_12611,N_12478,N_12018);
or U12612 (N_12612,N_12463,N_12025);
or U12613 (N_12613,N_12088,N_12040);
and U12614 (N_12614,N_12165,N_12089);
or U12615 (N_12615,N_12433,N_12033);
xor U12616 (N_12616,N_12101,N_12203);
or U12617 (N_12617,N_12309,N_12443);
xnor U12618 (N_12618,N_12301,N_12170);
or U12619 (N_12619,N_12189,N_12225);
nand U12620 (N_12620,N_12091,N_12266);
xor U12621 (N_12621,N_12332,N_12133);
or U12622 (N_12622,N_12019,N_12156);
or U12623 (N_12623,N_12338,N_12470);
or U12624 (N_12624,N_12270,N_12417);
nor U12625 (N_12625,N_12026,N_12125);
nand U12626 (N_12626,N_12431,N_12076);
xor U12627 (N_12627,N_12169,N_12256);
nand U12628 (N_12628,N_12013,N_12355);
and U12629 (N_12629,N_12056,N_12134);
or U12630 (N_12630,N_12172,N_12081);
or U12631 (N_12631,N_12296,N_12137);
nand U12632 (N_12632,N_12057,N_12290);
xor U12633 (N_12633,N_12257,N_12258);
nor U12634 (N_12634,N_12437,N_12267);
nor U12635 (N_12635,N_12050,N_12393);
nand U12636 (N_12636,N_12186,N_12015);
xor U12637 (N_12637,N_12485,N_12377);
or U12638 (N_12638,N_12430,N_12418);
nand U12639 (N_12639,N_12318,N_12215);
nand U12640 (N_12640,N_12136,N_12284);
and U12641 (N_12641,N_12066,N_12206);
xnor U12642 (N_12642,N_12188,N_12211);
and U12643 (N_12643,N_12271,N_12415);
or U12644 (N_12644,N_12110,N_12114);
nor U12645 (N_12645,N_12253,N_12412);
xnor U12646 (N_12646,N_12388,N_12408);
xnor U12647 (N_12647,N_12238,N_12390);
and U12648 (N_12648,N_12080,N_12100);
or U12649 (N_12649,N_12283,N_12224);
xor U12650 (N_12650,N_12357,N_12273);
or U12651 (N_12651,N_12020,N_12031);
nand U12652 (N_12652,N_12111,N_12072);
xor U12653 (N_12653,N_12062,N_12313);
and U12654 (N_12654,N_12486,N_12446);
and U12655 (N_12655,N_12395,N_12116);
xnor U12656 (N_12656,N_12411,N_12339);
xor U12657 (N_12657,N_12043,N_12048);
nand U12658 (N_12658,N_12440,N_12102);
nor U12659 (N_12659,N_12276,N_12375);
xnor U12660 (N_12660,N_12378,N_12143);
and U12661 (N_12661,N_12414,N_12295);
nor U12662 (N_12662,N_12194,N_12461);
nor U12663 (N_12663,N_12209,N_12095);
nor U12664 (N_12664,N_12173,N_12042);
nor U12665 (N_12665,N_12314,N_12429);
xnor U12666 (N_12666,N_12382,N_12082);
xor U12667 (N_12667,N_12310,N_12007);
xor U12668 (N_12668,N_12201,N_12335);
xor U12669 (N_12669,N_12183,N_12347);
xor U12670 (N_12670,N_12094,N_12106);
xnor U12671 (N_12671,N_12368,N_12372);
nand U12672 (N_12672,N_12432,N_12259);
and U12673 (N_12673,N_12289,N_12241);
or U12674 (N_12674,N_12229,N_12038);
or U12675 (N_12675,N_12112,N_12141);
and U12676 (N_12676,N_12249,N_12389);
nand U12677 (N_12677,N_12176,N_12129);
nor U12678 (N_12678,N_12449,N_12139);
and U12679 (N_12679,N_12386,N_12497);
and U12680 (N_12680,N_12004,N_12083);
and U12681 (N_12681,N_12480,N_12009);
nand U12682 (N_12682,N_12030,N_12474);
nor U12683 (N_12683,N_12410,N_12032);
or U12684 (N_12684,N_12391,N_12239);
nor U12685 (N_12685,N_12344,N_12326);
nand U12686 (N_12686,N_12300,N_12274);
and U12687 (N_12687,N_12421,N_12008);
or U12688 (N_12688,N_12261,N_12045);
or U12689 (N_12689,N_12308,N_12265);
or U12690 (N_12690,N_12424,N_12029);
or U12691 (N_12691,N_12405,N_12362);
xnor U12692 (N_12692,N_12085,N_12364);
and U12693 (N_12693,N_12466,N_12208);
nand U12694 (N_12694,N_12268,N_12315);
xor U12695 (N_12695,N_12447,N_12053);
and U12696 (N_12696,N_12468,N_12420);
or U12697 (N_12697,N_12394,N_12419);
xnor U12698 (N_12698,N_12360,N_12059);
nor U12699 (N_12699,N_12442,N_12104);
or U12700 (N_12700,N_12367,N_12490);
and U12701 (N_12701,N_12149,N_12197);
nand U12702 (N_12702,N_12330,N_12334);
nand U12703 (N_12703,N_12311,N_12345);
and U12704 (N_12704,N_12439,N_12207);
or U12705 (N_12705,N_12277,N_12058);
nor U12706 (N_12706,N_12084,N_12464);
nand U12707 (N_12707,N_12254,N_12341);
or U12708 (N_12708,N_12462,N_12237);
or U12709 (N_12709,N_12320,N_12353);
nor U12710 (N_12710,N_12383,N_12324);
and U12711 (N_12711,N_12024,N_12342);
xnor U12712 (N_12712,N_12005,N_12204);
or U12713 (N_12713,N_12450,N_12087);
nand U12714 (N_12714,N_12409,N_12448);
nand U12715 (N_12715,N_12119,N_12404);
nor U12716 (N_12716,N_12487,N_12305);
nand U12717 (N_12717,N_12297,N_12484);
xnor U12718 (N_12718,N_12356,N_12160);
nand U12719 (N_12719,N_12401,N_12230);
nand U12720 (N_12720,N_12285,N_12370);
nand U12721 (N_12721,N_12396,N_12158);
and U12722 (N_12722,N_12051,N_12044);
nand U12723 (N_12723,N_12251,N_12171);
nor U12724 (N_12724,N_12455,N_12460);
and U12725 (N_12725,N_12140,N_12157);
nor U12726 (N_12726,N_12003,N_12482);
and U12727 (N_12727,N_12022,N_12293);
and U12728 (N_12728,N_12205,N_12384);
and U12729 (N_12729,N_12444,N_12177);
and U12730 (N_12730,N_12218,N_12358);
and U12731 (N_12731,N_12373,N_12017);
nor U12732 (N_12732,N_12340,N_12272);
and U12733 (N_12733,N_12105,N_12248);
and U12734 (N_12734,N_12471,N_12316);
nor U12735 (N_12735,N_12152,N_12175);
or U12736 (N_12736,N_12323,N_12479);
nor U12737 (N_12737,N_12219,N_12202);
nand U12738 (N_12738,N_12307,N_12245);
or U12739 (N_12739,N_12164,N_12121);
and U12740 (N_12740,N_12161,N_12473);
and U12741 (N_12741,N_12246,N_12144);
nor U12742 (N_12742,N_12287,N_12182);
and U12743 (N_12743,N_12092,N_12494);
nor U12744 (N_12744,N_12467,N_12226);
or U12745 (N_12745,N_12027,N_12068);
nor U12746 (N_12746,N_12096,N_12073);
or U12747 (N_12747,N_12303,N_12213);
or U12748 (N_12748,N_12243,N_12427);
or U12749 (N_12749,N_12260,N_12147);
nand U12750 (N_12750,N_12490,N_12150);
or U12751 (N_12751,N_12217,N_12351);
and U12752 (N_12752,N_12392,N_12110);
nor U12753 (N_12753,N_12295,N_12127);
xor U12754 (N_12754,N_12269,N_12367);
and U12755 (N_12755,N_12272,N_12455);
nor U12756 (N_12756,N_12252,N_12049);
and U12757 (N_12757,N_12269,N_12297);
or U12758 (N_12758,N_12343,N_12391);
nand U12759 (N_12759,N_12450,N_12318);
nand U12760 (N_12760,N_12465,N_12123);
xnor U12761 (N_12761,N_12145,N_12283);
or U12762 (N_12762,N_12378,N_12040);
nor U12763 (N_12763,N_12492,N_12371);
or U12764 (N_12764,N_12366,N_12084);
xnor U12765 (N_12765,N_12007,N_12422);
nor U12766 (N_12766,N_12012,N_12489);
nand U12767 (N_12767,N_12184,N_12101);
nand U12768 (N_12768,N_12137,N_12204);
nand U12769 (N_12769,N_12275,N_12276);
nand U12770 (N_12770,N_12274,N_12298);
and U12771 (N_12771,N_12346,N_12328);
or U12772 (N_12772,N_12286,N_12078);
and U12773 (N_12773,N_12073,N_12211);
nor U12774 (N_12774,N_12142,N_12452);
nor U12775 (N_12775,N_12322,N_12433);
xnor U12776 (N_12776,N_12495,N_12291);
nand U12777 (N_12777,N_12191,N_12471);
nor U12778 (N_12778,N_12019,N_12086);
and U12779 (N_12779,N_12360,N_12067);
or U12780 (N_12780,N_12308,N_12480);
or U12781 (N_12781,N_12229,N_12056);
nand U12782 (N_12782,N_12392,N_12129);
and U12783 (N_12783,N_12413,N_12383);
nand U12784 (N_12784,N_12205,N_12440);
xor U12785 (N_12785,N_12010,N_12486);
nand U12786 (N_12786,N_12338,N_12381);
nor U12787 (N_12787,N_12023,N_12412);
xnor U12788 (N_12788,N_12141,N_12185);
xnor U12789 (N_12789,N_12453,N_12259);
xor U12790 (N_12790,N_12085,N_12345);
xor U12791 (N_12791,N_12297,N_12279);
nor U12792 (N_12792,N_12151,N_12053);
nor U12793 (N_12793,N_12331,N_12418);
xor U12794 (N_12794,N_12011,N_12330);
xnor U12795 (N_12795,N_12313,N_12476);
xnor U12796 (N_12796,N_12376,N_12081);
xnor U12797 (N_12797,N_12468,N_12213);
nor U12798 (N_12798,N_12229,N_12352);
nand U12799 (N_12799,N_12044,N_12200);
or U12800 (N_12800,N_12345,N_12323);
nor U12801 (N_12801,N_12449,N_12365);
or U12802 (N_12802,N_12054,N_12333);
nand U12803 (N_12803,N_12497,N_12459);
xnor U12804 (N_12804,N_12196,N_12446);
or U12805 (N_12805,N_12255,N_12452);
nand U12806 (N_12806,N_12144,N_12117);
or U12807 (N_12807,N_12150,N_12331);
and U12808 (N_12808,N_12333,N_12128);
nand U12809 (N_12809,N_12466,N_12282);
xor U12810 (N_12810,N_12465,N_12442);
and U12811 (N_12811,N_12493,N_12247);
or U12812 (N_12812,N_12286,N_12121);
nand U12813 (N_12813,N_12356,N_12451);
nand U12814 (N_12814,N_12118,N_12328);
and U12815 (N_12815,N_12305,N_12062);
xnor U12816 (N_12816,N_12244,N_12437);
xor U12817 (N_12817,N_12086,N_12076);
and U12818 (N_12818,N_12333,N_12430);
xnor U12819 (N_12819,N_12277,N_12291);
or U12820 (N_12820,N_12256,N_12281);
nor U12821 (N_12821,N_12155,N_12335);
or U12822 (N_12822,N_12225,N_12043);
nor U12823 (N_12823,N_12183,N_12393);
nand U12824 (N_12824,N_12073,N_12402);
or U12825 (N_12825,N_12499,N_12230);
nor U12826 (N_12826,N_12154,N_12120);
nand U12827 (N_12827,N_12338,N_12244);
nor U12828 (N_12828,N_12432,N_12288);
nand U12829 (N_12829,N_12235,N_12003);
nand U12830 (N_12830,N_12047,N_12002);
and U12831 (N_12831,N_12356,N_12108);
nor U12832 (N_12832,N_12126,N_12132);
or U12833 (N_12833,N_12074,N_12444);
or U12834 (N_12834,N_12294,N_12005);
and U12835 (N_12835,N_12074,N_12399);
xor U12836 (N_12836,N_12140,N_12039);
xor U12837 (N_12837,N_12306,N_12311);
nand U12838 (N_12838,N_12448,N_12218);
nor U12839 (N_12839,N_12465,N_12446);
xnor U12840 (N_12840,N_12454,N_12246);
and U12841 (N_12841,N_12374,N_12148);
xor U12842 (N_12842,N_12394,N_12014);
nand U12843 (N_12843,N_12332,N_12384);
or U12844 (N_12844,N_12199,N_12435);
nand U12845 (N_12845,N_12075,N_12021);
or U12846 (N_12846,N_12412,N_12076);
or U12847 (N_12847,N_12412,N_12001);
nand U12848 (N_12848,N_12463,N_12020);
or U12849 (N_12849,N_12158,N_12163);
and U12850 (N_12850,N_12046,N_12341);
nand U12851 (N_12851,N_12270,N_12234);
xor U12852 (N_12852,N_12151,N_12374);
nand U12853 (N_12853,N_12250,N_12138);
or U12854 (N_12854,N_12203,N_12447);
and U12855 (N_12855,N_12279,N_12001);
nand U12856 (N_12856,N_12098,N_12354);
nor U12857 (N_12857,N_12402,N_12110);
or U12858 (N_12858,N_12152,N_12027);
or U12859 (N_12859,N_12328,N_12046);
nand U12860 (N_12860,N_12165,N_12244);
nor U12861 (N_12861,N_12022,N_12378);
nand U12862 (N_12862,N_12039,N_12309);
and U12863 (N_12863,N_12186,N_12353);
xnor U12864 (N_12864,N_12141,N_12202);
or U12865 (N_12865,N_12113,N_12078);
nand U12866 (N_12866,N_12187,N_12081);
nand U12867 (N_12867,N_12157,N_12070);
nor U12868 (N_12868,N_12020,N_12021);
nor U12869 (N_12869,N_12373,N_12108);
nor U12870 (N_12870,N_12296,N_12259);
xor U12871 (N_12871,N_12290,N_12470);
and U12872 (N_12872,N_12369,N_12280);
and U12873 (N_12873,N_12319,N_12202);
xor U12874 (N_12874,N_12163,N_12494);
and U12875 (N_12875,N_12294,N_12437);
xnor U12876 (N_12876,N_12178,N_12181);
xor U12877 (N_12877,N_12355,N_12143);
nand U12878 (N_12878,N_12017,N_12335);
nor U12879 (N_12879,N_12154,N_12098);
nor U12880 (N_12880,N_12380,N_12004);
and U12881 (N_12881,N_12293,N_12229);
nor U12882 (N_12882,N_12118,N_12253);
or U12883 (N_12883,N_12044,N_12466);
nand U12884 (N_12884,N_12413,N_12483);
nor U12885 (N_12885,N_12002,N_12386);
nor U12886 (N_12886,N_12477,N_12016);
nor U12887 (N_12887,N_12338,N_12358);
xnor U12888 (N_12888,N_12058,N_12358);
and U12889 (N_12889,N_12025,N_12340);
nand U12890 (N_12890,N_12412,N_12462);
nor U12891 (N_12891,N_12452,N_12160);
or U12892 (N_12892,N_12465,N_12016);
xnor U12893 (N_12893,N_12460,N_12199);
and U12894 (N_12894,N_12112,N_12162);
nand U12895 (N_12895,N_12365,N_12047);
nor U12896 (N_12896,N_12117,N_12400);
xnor U12897 (N_12897,N_12083,N_12150);
nand U12898 (N_12898,N_12225,N_12246);
and U12899 (N_12899,N_12046,N_12235);
and U12900 (N_12900,N_12388,N_12458);
nand U12901 (N_12901,N_12262,N_12056);
nor U12902 (N_12902,N_12202,N_12387);
or U12903 (N_12903,N_12140,N_12231);
and U12904 (N_12904,N_12337,N_12018);
xnor U12905 (N_12905,N_12097,N_12235);
xor U12906 (N_12906,N_12102,N_12094);
nor U12907 (N_12907,N_12088,N_12082);
nand U12908 (N_12908,N_12085,N_12432);
nand U12909 (N_12909,N_12169,N_12441);
nor U12910 (N_12910,N_12215,N_12311);
xor U12911 (N_12911,N_12133,N_12037);
nand U12912 (N_12912,N_12290,N_12398);
or U12913 (N_12913,N_12243,N_12051);
xnor U12914 (N_12914,N_12236,N_12005);
nand U12915 (N_12915,N_12390,N_12365);
xnor U12916 (N_12916,N_12081,N_12173);
nand U12917 (N_12917,N_12065,N_12053);
and U12918 (N_12918,N_12441,N_12474);
nor U12919 (N_12919,N_12027,N_12137);
or U12920 (N_12920,N_12038,N_12094);
and U12921 (N_12921,N_12236,N_12463);
nor U12922 (N_12922,N_12254,N_12405);
nand U12923 (N_12923,N_12042,N_12287);
nand U12924 (N_12924,N_12417,N_12183);
or U12925 (N_12925,N_12463,N_12395);
xor U12926 (N_12926,N_12036,N_12174);
nor U12927 (N_12927,N_12169,N_12383);
xor U12928 (N_12928,N_12377,N_12101);
nand U12929 (N_12929,N_12412,N_12263);
nand U12930 (N_12930,N_12162,N_12462);
nand U12931 (N_12931,N_12106,N_12362);
nor U12932 (N_12932,N_12279,N_12376);
nand U12933 (N_12933,N_12094,N_12300);
nor U12934 (N_12934,N_12498,N_12307);
xnor U12935 (N_12935,N_12197,N_12012);
or U12936 (N_12936,N_12002,N_12221);
nand U12937 (N_12937,N_12375,N_12116);
or U12938 (N_12938,N_12191,N_12318);
and U12939 (N_12939,N_12435,N_12245);
and U12940 (N_12940,N_12291,N_12061);
nand U12941 (N_12941,N_12460,N_12255);
or U12942 (N_12942,N_12181,N_12352);
nor U12943 (N_12943,N_12059,N_12294);
nor U12944 (N_12944,N_12063,N_12289);
and U12945 (N_12945,N_12208,N_12021);
and U12946 (N_12946,N_12095,N_12267);
nor U12947 (N_12947,N_12016,N_12172);
and U12948 (N_12948,N_12343,N_12493);
or U12949 (N_12949,N_12064,N_12089);
or U12950 (N_12950,N_12158,N_12272);
xnor U12951 (N_12951,N_12384,N_12128);
or U12952 (N_12952,N_12153,N_12338);
and U12953 (N_12953,N_12363,N_12022);
nand U12954 (N_12954,N_12379,N_12257);
xor U12955 (N_12955,N_12135,N_12071);
nand U12956 (N_12956,N_12336,N_12390);
nand U12957 (N_12957,N_12245,N_12152);
xor U12958 (N_12958,N_12388,N_12230);
nor U12959 (N_12959,N_12266,N_12232);
nand U12960 (N_12960,N_12289,N_12208);
xnor U12961 (N_12961,N_12356,N_12389);
nand U12962 (N_12962,N_12328,N_12065);
or U12963 (N_12963,N_12353,N_12310);
or U12964 (N_12964,N_12225,N_12291);
or U12965 (N_12965,N_12194,N_12085);
nor U12966 (N_12966,N_12006,N_12342);
nand U12967 (N_12967,N_12279,N_12253);
nand U12968 (N_12968,N_12253,N_12174);
or U12969 (N_12969,N_12384,N_12072);
nor U12970 (N_12970,N_12009,N_12349);
or U12971 (N_12971,N_12258,N_12376);
nand U12972 (N_12972,N_12126,N_12227);
or U12973 (N_12973,N_12269,N_12227);
nand U12974 (N_12974,N_12132,N_12094);
and U12975 (N_12975,N_12010,N_12228);
or U12976 (N_12976,N_12227,N_12465);
or U12977 (N_12977,N_12386,N_12092);
nor U12978 (N_12978,N_12023,N_12436);
nand U12979 (N_12979,N_12123,N_12040);
xnor U12980 (N_12980,N_12431,N_12205);
nand U12981 (N_12981,N_12226,N_12233);
and U12982 (N_12982,N_12067,N_12045);
and U12983 (N_12983,N_12460,N_12216);
xor U12984 (N_12984,N_12336,N_12397);
xnor U12985 (N_12985,N_12443,N_12015);
nor U12986 (N_12986,N_12495,N_12122);
or U12987 (N_12987,N_12392,N_12318);
nor U12988 (N_12988,N_12378,N_12412);
nand U12989 (N_12989,N_12460,N_12104);
xor U12990 (N_12990,N_12245,N_12491);
nor U12991 (N_12991,N_12461,N_12243);
nor U12992 (N_12992,N_12344,N_12411);
nor U12993 (N_12993,N_12120,N_12468);
nand U12994 (N_12994,N_12244,N_12413);
nand U12995 (N_12995,N_12244,N_12134);
xnor U12996 (N_12996,N_12071,N_12420);
nand U12997 (N_12997,N_12424,N_12050);
nand U12998 (N_12998,N_12079,N_12494);
nor U12999 (N_12999,N_12105,N_12419);
or U13000 (N_13000,N_12904,N_12716);
and U13001 (N_13001,N_12771,N_12621);
or U13002 (N_13002,N_12786,N_12737);
xnor U13003 (N_13003,N_12501,N_12962);
nor U13004 (N_13004,N_12964,N_12511);
and U13005 (N_13005,N_12997,N_12687);
nand U13006 (N_13006,N_12577,N_12730);
nand U13007 (N_13007,N_12895,N_12767);
or U13008 (N_13008,N_12925,N_12533);
or U13009 (N_13009,N_12700,N_12884);
or U13010 (N_13010,N_12978,N_12571);
and U13011 (N_13011,N_12833,N_12512);
and U13012 (N_13012,N_12957,N_12672);
and U13013 (N_13013,N_12627,N_12788);
or U13014 (N_13014,N_12747,N_12597);
xnor U13015 (N_13015,N_12675,N_12686);
nor U13016 (N_13016,N_12709,N_12924);
nand U13017 (N_13017,N_12845,N_12612);
nand U13018 (N_13018,N_12732,N_12685);
nand U13019 (N_13019,N_12509,N_12541);
xor U13020 (N_13020,N_12914,N_12699);
and U13021 (N_13021,N_12857,N_12664);
nor U13022 (N_13022,N_12630,N_12937);
or U13023 (N_13023,N_12979,N_12929);
and U13024 (N_13024,N_12795,N_12837);
and U13025 (N_13025,N_12559,N_12696);
nor U13026 (N_13026,N_12887,N_12564);
xnor U13027 (N_13027,N_12897,N_12774);
xnor U13028 (N_13028,N_12622,N_12866);
xor U13029 (N_13029,N_12817,N_12872);
and U13030 (N_13030,N_12603,N_12618);
nor U13031 (N_13031,N_12635,N_12575);
xor U13032 (N_13032,N_12799,N_12764);
and U13033 (N_13033,N_12827,N_12809);
nand U13034 (N_13034,N_12915,N_12530);
and U13035 (N_13035,N_12835,N_12873);
nor U13036 (N_13036,N_12824,N_12531);
xor U13037 (N_13037,N_12840,N_12593);
nand U13038 (N_13038,N_12901,N_12846);
xor U13039 (N_13039,N_12549,N_12877);
or U13040 (N_13040,N_12665,N_12981);
nand U13041 (N_13041,N_12663,N_12992);
nor U13042 (N_13042,N_12503,N_12582);
nor U13043 (N_13043,N_12898,N_12996);
nor U13044 (N_13044,N_12982,N_12602);
or U13045 (N_13045,N_12615,N_12763);
or U13046 (N_13046,N_12619,N_12752);
and U13047 (N_13047,N_12868,N_12975);
nor U13048 (N_13048,N_12820,N_12894);
nand U13049 (N_13049,N_12911,N_12762);
xnor U13050 (N_13050,N_12540,N_12959);
nand U13051 (N_13051,N_12811,N_12655);
and U13052 (N_13052,N_12885,N_12576);
or U13053 (N_13053,N_12573,N_12639);
nor U13054 (N_13054,N_12591,N_12669);
or U13055 (N_13055,N_12798,N_12725);
xnor U13056 (N_13056,N_12688,N_12754);
nand U13057 (N_13057,N_12768,N_12727);
or U13058 (N_13058,N_12753,N_12584);
and U13059 (N_13059,N_12706,N_12526);
or U13060 (N_13060,N_12759,N_12710);
and U13061 (N_13061,N_12968,N_12967);
nand U13062 (N_13062,N_12773,N_12938);
and U13063 (N_13063,N_12613,N_12947);
nor U13064 (N_13064,N_12524,N_12604);
nor U13065 (N_13065,N_12547,N_12505);
or U13066 (N_13066,N_12864,N_12538);
xor U13067 (N_13067,N_12607,N_12670);
nor U13068 (N_13068,N_12698,N_12916);
and U13069 (N_13069,N_12965,N_12870);
xnor U13070 (N_13070,N_12985,N_12579);
xnor U13071 (N_13071,N_12632,N_12739);
and U13072 (N_13072,N_12896,N_12831);
nand U13073 (N_13073,N_12535,N_12515);
or U13074 (N_13074,N_12590,N_12761);
xor U13075 (N_13075,N_12802,N_12674);
or U13076 (N_13076,N_12955,N_12879);
xor U13077 (N_13077,N_12713,N_12646);
xnor U13078 (N_13078,N_12797,N_12942);
or U13079 (N_13079,N_12594,N_12726);
or U13080 (N_13080,N_12500,N_12731);
or U13081 (N_13081,N_12527,N_12690);
or U13082 (N_13082,N_12828,N_12645);
nand U13083 (N_13083,N_12766,N_12949);
nor U13084 (N_13084,N_12550,N_12912);
and U13085 (N_13085,N_12769,N_12510);
and U13086 (N_13086,N_12728,N_12789);
and U13087 (N_13087,N_12717,N_12810);
nand U13088 (N_13088,N_12702,N_12814);
nor U13089 (N_13089,N_12909,N_12544);
nand U13090 (N_13090,N_12936,N_12553);
xor U13091 (N_13091,N_12601,N_12654);
nand U13092 (N_13092,N_12636,N_12583);
or U13093 (N_13093,N_12660,N_12623);
nor U13094 (N_13094,N_12973,N_12958);
xor U13095 (N_13095,N_12528,N_12647);
and U13096 (N_13096,N_12869,N_12792);
or U13097 (N_13097,N_12841,N_12933);
xor U13098 (N_13098,N_12542,N_12922);
or U13099 (N_13099,N_12668,N_12609);
nand U13100 (N_13100,N_12520,N_12961);
or U13101 (N_13101,N_12880,N_12863);
or U13102 (N_13102,N_12539,N_12614);
nand U13103 (N_13103,N_12755,N_12948);
and U13104 (N_13104,N_12923,N_12977);
nand U13105 (N_13105,N_12850,N_12781);
nor U13106 (N_13106,N_12677,N_12648);
nor U13107 (N_13107,N_12637,N_12718);
or U13108 (N_13108,N_12858,N_12723);
nor U13109 (N_13109,N_12756,N_12859);
xnor U13110 (N_13110,N_12998,N_12839);
nand U13111 (N_13111,N_12946,N_12643);
and U13112 (N_13112,N_12765,N_12680);
nand U13113 (N_13113,N_12989,N_12740);
xor U13114 (N_13114,N_12954,N_12504);
and U13115 (N_13115,N_12729,N_12681);
xor U13116 (N_13116,N_12860,N_12852);
or U13117 (N_13117,N_12715,N_12694);
nand U13118 (N_13118,N_12558,N_12746);
nor U13119 (N_13119,N_12777,N_12722);
or U13120 (N_13120,N_12628,N_12776);
or U13121 (N_13121,N_12823,N_12930);
and U13122 (N_13122,N_12679,N_12598);
xnor U13123 (N_13123,N_12745,N_12805);
or U13124 (N_13124,N_12804,N_12758);
nor U13125 (N_13125,N_12812,N_12704);
or U13126 (N_13126,N_12658,N_12775);
xnor U13127 (N_13127,N_12748,N_12890);
nor U13128 (N_13128,N_12760,N_12794);
and U13129 (N_13129,N_12691,N_12529);
and U13130 (N_13130,N_12659,N_12662);
xor U13131 (N_13131,N_12641,N_12712);
and U13132 (N_13132,N_12651,N_12711);
nor U13133 (N_13133,N_12692,N_12834);
nor U13134 (N_13134,N_12772,N_12803);
xnor U13135 (N_13135,N_12703,N_12871);
xor U13136 (N_13136,N_12854,N_12517);
and U13137 (N_13137,N_12851,N_12617);
nand U13138 (N_13138,N_12552,N_12525);
and U13139 (N_13139,N_12782,N_12506);
nor U13140 (N_13140,N_12983,N_12631);
or U13141 (N_13141,N_12900,N_12984);
and U13142 (N_13142,N_12838,N_12578);
nand U13143 (N_13143,N_12932,N_12832);
nor U13144 (N_13144,N_12910,N_12689);
and U13145 (N_13145,N_12861,N_12656);
and U13146 (N_13146,N_12653,N_12652);
xnor U13147 (N_13147,N_12951,N_12707);
xor U13148 (N_13148,N_12620,N_12970);
and U13149 (N_13149,N_12642,N_12701);
nand U13150 (N_13150,N_12638,N_12826);
and U13151 (N_13151,N_12574,N_12518);
xor U13152 (N_13152,N_12836,N_12939);
nor U13153 (N_13153,N_12567,N_12757);
and U13154 (N_13154,N_12588,N_12822);
and U13155 (N_13155,N_12565,N_12551);
xnor U13156 (N_13156,N_12561,N_12848);
xnor U13157 (N_13157,N_12796,N_12994);
and U13158 (N_13158,N_12546,N_12523);
nand U13159 (N_13159,N_12891,N_12741);
xor U13160 (N_13160,N_12956,N_12719);
nor U13161 (N_13161,N_12563,N_12963);
xor U13162 (N_13162,N_12750,N_12980);
xnor U13163 (N_13163,N_12855,N_12650);
or U13164 (N_13164,N_12592,N_12875);
nand U13165 (N_13165,N_12986,N_12534);
nor U13166 (N_13166,N_12724,N_12581);
xnor U13167 (N_13167,N_12883,N_12847);
nand U13168 (N_13168,N_12749,N_12736);
and U13169 (N_13169,N_12993,N_12783);
or U13170 (N_13170,N_12508,N_12566);
or U13171 (N_13171,N_12522,N_12626);
xnor U13172 (N_13172,N_12844,N_12537);
nor U13173 (N_13173,N_12589,N_12743);
xor U13174 (N_13174,N_12676,N_12905);
nand U13175 (N_13175,N_12972,N_12807);
nor U13176 (N_13176,N_12634,N_12562);
or U13177 (N_13177,N_12849,N_12610);
or U13178 (N_13178,N_12580,N_12999);
or U13179 (N_13179,N_12640,N_12734);
nand U13180 (N_13180,N_12543,N_12507);
xor U13181 (N_13181,N_12666,N_12587);
and U13182 (N_13182,N_12976,N_12842);
nand U13183 (N_13183,N_12806,N_12867);
and U13184 (N_13184,N_12596,N_12953);
and U13185 (N_13185,N_12819,N_12926);
nor U13186 (N_13186,N_12952,N_12818);
or U13187 (N_13187,N_12536,N_12555);
nand U13188 (N_13188,N_12892,N_12899);
nor U13189 (N_13189,N_12931,N_12673);
xor U13190 (N_13190,N_12876,N_12742);
or U13191 (N_13191,N_12790,N_12893);
xnor U13192 (N_13192,N_12945,N_12557);
nor U13193 (N_13193,N_12682,N_12878);
nor U13194 (N_13194,N_12940,N_12586);
or U13195 (N_13195,N_12865,N_12720);
nor U13196 (N_13196,N_12950,N_12902);
nand U13197 (N_13197,N_12667,N_12695);
nor U13198 (N_13198,N_12570,N_12644);
nand U13199 (N_13199,N_12751,N_12793);
and U13200 (N_13200,N_12502,N_12625);
nand U13201 (N_13201,N_12800,N_12988);
xnor U13202 (N_13202,N_12516,N_12572);
or U13203 (N_13203,N_12974,N_12960);
nand U13204 (N_13204,N_12569,N_12843);
xor U13205 (N_13205,N_12600,N_12991);
xor U13206 (N_13206,N_12825,N_12684);
nor U13207 (N_13207,N_12554,N_12966);
nor U13208 (N_13208,N_12918,N_12599);
and U13209 (N_13209,N_12683,N_12556);
and U13210 (N_13210,N_12605,N_12714);
or U13211 (N_13211,N_12738,N_12791);
xor U13212 (N_13212,N_12521,N_12513);
nand U13213 (N_13213,N_12920,N_12862);
and U13214 (N_13214,N_12815,N_12816);
xnor U13215 (N_13215,N_12770,N_12697);
or U13216 (N_13216,N_12785,N_12995);
and U13217 (N_13217,N_12830,N_12611);
or U13218 (N_13218,N_12990,N_12629);
or U13219 (N_13219,N_12969,N_12548);
or U13220 (N_13220,N_12808,N_12921);
or U13221 (N_13221,N_12928,N_12568);
nand U13222 (N_13222,N_12560,N_12721);
and U13223 (N_13223,N_12943,N_12616);
and U13224 (N_13224,N_12917,N_12661);
xnor U13225 (N_13225,N_12944,N_12608);
nand U13226 (N_13226,N_12801,N_12906);
or U13227 (N_13227,N_12874,N_12780);
or U13228 (N_13228,N_12829,N_12705);
and U13229 (N_13229,N_12735,N_12934);
nor U13230 (N_13230,N_12693,N_12856);
nor U13231 (N_13231,N_12935,N_12881);
or U13232 (N_13232,N_12813,N_12733);
nor U13233 (N_13233,N_12708,N_12821);
nand U13234 (N_13234,N_12882,N_12907);
xnor U13235 (N_13235,N_12657,N_12927);
nand U13236 (N_13236,N_12678,N_12649);
nand U13237 (N_13237,N_12888,N_12941);
or U13238 (N_13238,N_12595,N_12778);
nor U13239 (N_13239,N_12919,N_12784);
nand U13240 (N_13240,N_12532,N_12908);
and U13241 (N_13241,N_12971,N_12545);
or U13242 (N_13242,N_12633,N_12519);
and U13243 (N_13243,N_12987,N_12606);
nand U13244 (N_13244,N_12779,N_12744);
xnor U13245 (N_13245,N_12903,N_12886);
and U13246 (N_13246,N_12787,N_12514);
and U13247 (N_13247,N_12585,N_12853);
or U13248 (N_13248,N_12624,N_12889);
or U13249 (N_13249,N_12913,N_12671);
and U13250 (N_13250,N_12954,N_12579);
nor U13251 (N_13251,N_12619,N_12606);
nand U13252 (N_13252,N_12601,N_12784);
and U13253 (N_13253,N_12958,N_12733);
or U13254 (N_13254,N_12731,N_12557);
or U13255 (N_13255,N_12560,N_12689);
nand U13256 (N_13256,N_12808,N_12766);
or U13257 (N_13257,N_12721,N_12750);
xnor U13258 (N_13258,N_12581,N_12788);
xor U13259 (N_13259,N_12568,N_12827);
or U13260 (N_13260,N_12659,N_12706);
xnor U13261 (N_13261,N_12565,N_12847);
and U13262 (N_13262,N_12516,N_12951);
and U13263 (N_13263,N_12636,N_12658);
or U13264 (N_13264,N_12666,N_12973);
or U13265 (N_13265,N_12922,N_12755);
or U13266 (N_13266,N_12725,N_12566);
nor U13267 (N_13267,N_12626,N_12758);
nand U13268 (N_13268,N_12962,N_12880);
and U13269 (N_13269,N_12810,N_12968);
nand U13270 (N_13270,N_12646,N_12507);
nor U13271 (N_13271,N_12999,N_12653);
nand U13272 (N_13272,N_12906,N_12721);
or U13273 (N_13273,N_12641,N_12753);
or U13274 (N_13274,N_12626,N_12900);
or U13275 (N_13275,N_12790,N_12705);
and U13276 (N_13276,N_12622,N_12756);
nand U13277 (N_13277,N_12776,N_12793);
or U13278 (N_13278,N_12656,N_12866);
xor U13279 (N_13279,N_12511,N_12578);
nand U13280 (N_13280,N_12551,N_12571);
and U13281 (N_13281,N_12631,N_12947);
xor U13282 (N_13282,N_12582,N_12674);
xor U13283 (N_13283,N_12682,N_12954);
nand U13284 (N_13284,N_12806,N_12972);
or U13285 (N_13285,N_12821,N_12677);
xor U13286 (N_13286,N_12631,N_12813);
and U13287 (N_13287,N_12647,N_12724);
and U13288 (N_13288,N_12823,N_12928);
nand U13289 (N_13289,N_12616,N_12792);
nor U13290 (N_13290,N_12526,N_12681);
or U13291 (N_13291,N_12563,N_12862);
nand U13292 (N_13292,N_12611,N_12509);
nand U13293 (N_13293,N_12568,N_12854);
nand U13294 (N_13294,N_12969,N_12785);
xor U13295 (N_13295,N_12956,N_12774);
and U13296 (N_13296,N_12773,N_12777);
or U13297 (N_13297,N_12651,N_12547);
or U13298 (N_13298,N_12740,N_12671);
and U13299 (N_13299,N_12804,N_12556);
nand U13300 (N_13300,N_12712,N_12925);
and U13301 (N_13301,N_12534,N_12788);
nand U13302 (N_13302,N_12899,N_12603);
xor U13303 (N_13303,N_12863,N_12736);
xor U13304 (N_13304,N_12892,N_12727);
nand U13305 (N_13305,N_12555,N_12986);
or U13306 (N_13306,N_12891,N_12972);
nand U13307 (N_13307,N_12667,N_12687);
or U13308 (N_13308,N_12910,N_12645);
nor U13309 (N_13309,N_12610,N_12820);
xnor U13310 (N_13310,N_12905,N_12882);
and U13311 (N_13311,N_12820,N_12825);
xor U13312 (N_13312,N_12531,N_12990);
or U13313 (N_13313,N_12930,N_12985);
nand U13314 (N_13314,N_12814,N_12691);
nand U13315 (N_13315,N_12880,N_12862);
nand U13316 (N_13316,N_12535,N_12582);
nor U13317 (N_13317,N_12517,N_12571);
or U13318 (N_13318,N_12536,N_12651);
nand U13319 (N_13319,N_12831,N_12623);
nand U13320 (N_13320,N_12946,N_12695);
xor U13321 (N_13321,N_12988,N_12614);
or U13322 (N_13322,N_12646,N_12775);
nor U13323 (N_13323,N_12938,N_12631);
or U13324 (N_13324,N_12698,N_12884);
xnor U13325 (N_13325,N_12797,N_12643);
xnor U13326 (N_13326,N_12537,N_12593);
xor U13327 (N_13327,N_12733,N_12707);
xor U13328 (N_13328,N_12520,N_12601);
nor U13329 (N_13329,N_12874,N_12623);
and U13330 (N_13330,N_12503,N_12548);
or U13331 (N_13331,N_12938,N_12903);
xor U13332 (N_13332,N_12584,N_12687);
or U13333 (N_13333,N_12745,N_12986);
or U13334 (N_13334,N_12670,N_12806);
and U13335 (N_13335,N_12741,N_12500);
nor U13336 (N_13336,N_12972,N_12589);
nand U13337 (N_13337,N_12724,N_12874);
nand U13338 (N_13338,N_12623,N_12724);
xor U13339 (N_13339,N_12774,N_12923);
or U13340 (N_13340,N_12673,N_12827);
or U13341 (N_13341,N_12522,N_12873);
nor U13342 (N_13342,N_12619,N_12660);
and U13343 (N_13343,N_12561,N_12633);
nor U13344 (N_13344,N_12717,N_12505);
and U13345 (N_13345,N_12710,N_12532);
xor U13346 (N_13346,N_12962,N_12749);
nor U13347 (N_13347,N_12542,N_12630);
nand U13348 (N_13348,N_12826,N_12543);
nand U13349 (N_13349,N_12849,N_12735);
and U13350 (N_13350,N_12510,N_12910);
and U13351 (N_13351,N_12771,N_12899);
xor U13352 (N_13352,N_12714,N_12607);
xnor U13353 (N_13353,N_12709,N_12912);
xnor U13354 (N_13354,N_12656,N_12933);
and U13355 (N_13355,N_12583,N_12506);
and U13356 (N_13356,N_12599,N_12675);
and U13357 (N_13357,N_12872,N_12689);
or U13358 (N_13358,N_12933,N_12517);
xnor U13359 (N_13359,N_12875,N_12695);
nor U13360 (N_13360,N_12841,N_12770);
xor U13361 (N_13361,N_12605,N_12856);
xor U13362 (N_13362,N_12954,N_12692);
nand U13363 (N_13363,N_12509,N_12711);
nand U13364 (N_13364,N_12561,N_12810);
or U13365 (N_13365,N_12645,N_12737);
nand U13366 (N_13366,N_12760,N_12543);
xnor U13367 (N_13367,N_12838,N_12664);
and U13368 (N_13368,N_12908,N_12615);
xor U13369 (N_13369,N_12631,N_12740);
or U13370 (N_13370,N_12666,N_12724);
nand U13371 (N_13371,N_12796,N_12631);
xnor U13372 (N_13372,N_12816,N_12758);
and U13373 (N_13373,N_12836,N_12822);
xor U13374 (N_13374,N_12950,N_12563);
xor U13375 (N_13375,N_12921,N_12939);
and U13376 (N_13376,N_12622,N_12669);
and U13377 (N_13377,N_12510,N_12558);
nor U13378 (N_13378,N_12717,N_12796);
nor U13379 (N_13379,N_12501,N_12937);
xor U13380 (N_13380,N_12659,N_12912);
nor U13381 (N_13381,N_12667,N_12656);
or U13382 (N_13382,N_12910,N_12868);
or U13383 (N_13383,N_12845,N_12543);
or U13384 (N_13384,N_12856,N_12947);
and U13385 (N_13385,N_12548,N_12978);
xnor U13386 (N_13386,N_12901,N_12570);
or U13387 (N_13387,N_12994,N_12630);
xnor U13388 (N_13388,N_12604,N_12964);
nand U13389 (N_13389,N_12832,N_12870);
and U13390 (N_13390,N_12827,N_12943);
nor U13391 (N_13391,N_12790,N_12797);
xnor U13392 (N_13392,N_12854,N_12792);
nand U13393 (N_13393,N_12929,N_12915);
and U13394 (N_13394,N_12541,N_12800);
xnor U13395 (N_13395,N_12695,N_12981);
nor U13396 (N_13396,N_12804,N_12578);
and U13397 (N_13397,N_12691,N_12786);
nor U13398 (N_13398,N_12553,N_12544);
nand U13399 (N_13399,N_12907,N_12710);
and U13400 (N_13400,N_12544,N_12743);
or U13401 (N_13401,N_12593,N_12993);
xor U13402 (N_13402,N_12908,N_12903);
nor U13403 (N_13403,N_12503,N_12956);
nand U13404 (N_13404,N_12951,N_12688);
and U13405 (N_13405,N_12864,N_12632);
or U13406 (N_13406,N_12972,N_12510);
or U13407 (N_13407,N_12604,N_12516);
nand U13408 (N_13408,N_12652,N_12548);
nand U13409 (N_13409,N_12848,N_12940);
and U13410 (N_13410,N_12947,N_12687);
or U13411 (N_13411,N_12656,N_12869);
xor U13412 (N_13412,N_12598,N_12906);
xor U13413 (N_13413,N_12803,N_12620);
nor U13414 (N_13414,N_12799,N_12970);
nor U13415 (N_13415,N_12651,N_12662);
or U13416 (N_13416,N_12564,N_12552);
nand U13417 (N_13417,N_12773,N_12533);
nand U13418 (N_13418,N_12763,N_12956);
and U13419 (N_13419,N_12790,N_12603);
nor U13420 (N_13420,N_12819,N_12659);
xor U13421 (N_13421,N_12695,N_12927);
nand U13422 (N_13422,N_12624,N_12540);
or U13423 (N_13423,N_12708,N_12834);
nor U13424 (N_13424,N_12570,N_12799);
xnor U13425 (N_13425,N_12558,N_12596);
nor U13426 (N_13426,N_12913,N_12935);
nor U13427 (N_13427,N_12766,N_12740);
nand U13428 (N_13428,N_12545,N_12563);
and U13429 (N_13429,N_12585,N_12836);
or U13430 (N_13430,N_12724,N_12700);
nand U13431 (N_13431,N_12771,N_12876);
xnor U13432 (N_13432,N_12640,N_12785);
or U13433 (N_13433,N_12662,N_12918);
nor U13434 (N_13434,N_12556,N_12931);
xnor U13435 (N_13435,N_12787,N_12897);
nor U13436 (N_13436,N_12868,N_12692);
nand U13437 (N_13437,N_12576,N_12803);
xnor U13438 (N_13438,N_12814,N_12795);
nor U13439 (N_13439,N_12713,N_12843);
nand U13440 (N_13440,N_12865,N_12626);
or U13441 (N_13441,N_12753,N_12629);
and U13442 (N_13442,N_12839,N_12566);
nand U13443 (N_13443,N_12902,N_12911);
or U13444 (N_13444,N_12769,N_12847);
xor U13445 (N_13445,N_12773,N_12842);
xnor U13446 (N_13446,N_12890,N_12711);
nand U13447 (N_13447,N_12653,N_12852);
xnor U13448 (N_13448,N_12817,N_12691);
nor U13449 (N_13449,N_12661,N_12719);
xor U13450 (N_13450,N_12678,N_12858);
nor U13451 (N_13451,N_12959,N_12532);
nand U13452 (N_13452,N_12960,N_12667);
or U13453 (N_13453,N_12643,N_12873);
or U13454 (N_13454,N_12823,N_12970);
or U13455 (N_13455,N_12871,N_12823);
nand U13456 (N_13456,N_12691,N_12794);
xor U13457 (N_13457,N_12731,N_12946);
and U13458 (N_13458,N_12909,N_12555);
xnor U13459 (N_13459,N_12688,N_12971);
xnor U13460 (N_13460,N_12979,N_12692);
or U13461 (N_13461,N_12707,N_12594);
nor U13462 (N_13462,N_12575,N_12922);
nor U13463 (N_13463,N_12866,N_12786);
and U13464 (N_13464,N_12923,N_12826);
nand U13465 (N_13465,N_12928,N_12818);
xor U13466 (N_13466,N_12877,N_12906);
nand U13467 (N_13467,N_12996,N_12986);
nand U13468 (N_13468,N_12792,N_12631);
nor U13469 (N_13469,N_12554,N_12744);
or U13470 (N_13470,N_12797,N_12640);
nor U13471 (N_13471,N_12781,N_12765);
nor U13472 (N_13472,N_12752,N_12668);
or U13473 (N_13473,N_12822,N_12941);
and U13474 (N_13474,N_12624,N_12592);
or U13475 (N_13475,N_12716,N_12728);
xor U13476 (N_13476,N_12834,N_12563);
xnor U13477 (N_13477,N_12718,N_12765);
nor U13478 (N_13478,N_12504,N_12888);
xor U13479 (N_13479,N_12661,N_12869);
xnor U13480 (N_13480,N_12783,N_12532);
or U13481 (N_13481,N_12793,N_12500);
and U13482 (N_13482,N_12859,N_12991);
and U13483 (N_13483,N_12976,N_12998);
and U13484 (N_13484,N_12817,N_12744);
xnor U13485 (N_13485,N_12752,N_12962);
xnor U13486 (N_13486,N_12983,N_12823);
and U13487 (N_13487,N_12926,N_12586);
nor U13488 (N_13488,N_12534,N_12590);
nand U13489 (N_13489,N_12660,N_12540);
xor U13490 (N_13490,N_12884,N_12563);
nor U13491 (N_13491,N_12535,N_12887);
and U13492 (N_13492,N_12566,N_12754);
and U13493 (N_13493,N_12899,N_12588);
or U13494 (N_13494,N_12945,N_12787);
nor U13495 (N_13495,N_12562,N_12608);
or U13496 (N_13496,N_12988,N_12556);
nand U13497 (N_13497,N_12846,N_12948);
or U13498 (N_13498,N_12848,N_12892);
xnor U13499 (N_13499,N_12764,N_12989);
nor U13500 (N_13500,N_13399,N_13341);
and U13501 (N_13501,N_13490,N_13374);
xor U13502 (N_13502,N_13079,N_13058);
or U13503 (N_13503,N_13092,N_13190);
nor U13504 (N_13504,N_13276,N_13155);
nand U13505 (N_13505,N_13274,N_13157);
nand U13506 (N_13506,N_13458,N_13060);
nand U13507 (N_13507,N_13169,N_13351);
xor U13508 (N_13508,N_13259,N_13459);
xor U13509 (N_13509,N_13313,N_13487);
nand U13510 (N_13510,N_13446,N_13448);
or U13511 (N_13511,N_13204,N_13476);
and U13512 (N_13512,N_13095,N_13427);
nor U13513 (N_13513,N_13415,N_13452);
xor U13514 (N_13514,N_13425,N_13054);
nor U13515 (N_13515,N_13408,N_13188);
and U13516 (N_13516,N_13260,N_13349);
nor U13517 (N_13517,N_13442,N_13432);
and U13518 (N_13518,N_13353,N_13307);
or U13519 (N_13519,N_13499,N_13175);
or U13520 (N_13520,N_13347,N_13239);
nand U13521 (N_13521,N_13395,N_13311);
or U13522 (N_13522,N_13163,N_13382);
and U13523 (N_13523,N_13479,N_13215);
xor U13524 (N_13524,N_13370,N_13118);
or U13525 (N_13525,N_13271,N_13394);
and U13526 (N_13526,N_13363,N_13390);
or U13527 (N_13527,N_13352,N_13191);
or U13528 (N_13528,N_13158,N_13318);
xor U13529 (N_13529,N_13142,N_13401);
or U13530 (N_13530,N_13127,N_13102);
nor U13531 (N_13531,N_13094,N_13321);
nor U13532 (N_13532,N_13410,N_13391);
nor U13533 (N_13533,N_13430,N_13482);
and U13534 (N_13534,N_13231,N_13081);
or U13535 (N_13535,N_13251,N_13019);
xnor U13536 (N_13536,N_13316,N_13460);
xnor U13537 (N_13537,N_13290,N_13134);
or U13538 (N_13538,N_13380,N_13372);
nor U13539 (N_13539,N_13420,N_13084);
and U13540 (N_13540,N_13138,N_13133);
or U13541 (N_13541,N_13017,N_13419);
xnor U13542 (N_13542,N_13197,N_13464);
and U13543 (N_13543,N_13379,N_13113);
nand U13544 (N_13544,N_13069,N_13146);
nor U13545 (N_13545,N_13404,N_13129);
nand U13546 (N_13546,N_13020,N_13108);
xor U13547 (N_13547,N_13164,N_13210);
nor U13548 (N_13548,N_13320,N_13039);
nor U13549 (N_13549,N_13350,N_13240);
xor U13550 (N_13550,N_13193,N_13185);
or U13551 (N_13551,N_13326,N_13368);
or U13552 (N_13552,N_13270,N_13196);
nor U13553 (N_13553,N_13236,N_13145);
and U13554 (N_13554,N_13284,N_13120);
and U13555 (N_13555,N_13337,N_13428);
nand U13556 (N_13556,N_13227,N_13214);
nand U13557 (N_13557,N_13021,N_13469);
nor U13558 (N_13558,N_13243,N_13346);
or U13559 (N_13559,N_13160,N_13254);
nand U13560 (N_13560,N_13421,N_13480);
and U13561 (N_13561,N_13258,N_13264);
nand U13562 (N_13562,N_13206,N_13180);
xnor U13563 (N_13563,N_13063,N_13319);
and U13564 (N_13564,N_13070,N_13198);
xor U13565 (N_13565,N_13362,N_13001);
nand U13566 (N_13566,N_13250,N_13280);
and U13567 (N_13567,N_13167,N_13181);
or U13568 (N_13568,N_13219,N_13008);
and U13569 (N_13569,N_13493,N_13298);
and U13570 (N_13570,N_13287,N_13241);
and U13571 (N_13571,N_13025,N_13444);
and U13572 (N_13572,N_13300,N_13463);
or U13573 (N_13573,N_13100,N_13011);
or U13574 (N_13574,N_13327,N_13360);
nand U13575 (N_13575,N_13348,N_13494);
and U13576 (N_13576,N_13221,N_13333);
xnor U13577 (N_13577,N_13447,N_13294);
or U13578 (N_13578,N_13149,N_13230);
and U13579 (N_13579,N_13050,N_13246);
xnor U13580 (N_13580,N_13159,N_13179);
nor U13581 (N_13581,N_13114,N_13166);
xor U13582 (N_13582,N_13301,N_13140);
and U13583 (N_13583,N_13006,N_13066);
nor U13584 (N_13584,N_13378,N_13106);
xnor U13585 (N_13585,N_13109,N_13441);
and U13586 (N_13586,N_13199,N_13402);
and U13587 (N_13587,N_13031,N_13309);
nor U13588 (N_13588,N_13339,N_13137);
and U13589 (N_13589,N_13211,N_13338);
xor U13590 (N_13590,N_13073,N_13484);
and U13591 (N_13591,N_13183,N_13291);
nand U13592 (N_13592,N_13176,N_13229);
or U13593 (N_13593,N_13397,N_13304);
and U13594 (N_13594,N_13310,N_13451);
nand U13595 (N_13595,N_13289,N_13373);
and U13596 (N_13596,N_13010,N_13409);
nor U13597 (N_13597,N_13356,N_13007);
xor U13598 (N_13598,N_13178,N_13147);
nand U13599 (N_13599,N_13002,N_13381);
nor U13600 (N_13600,N_13096,N_13068);
and U13601 (N_13601,N_13201,N_13288);
xnor U13602 (N_13602,N_13152,N_13266);
and U13603 (N_13603,N_13483,N_13467);
and U13604 (N_13604,N_13189,N_13150);
nand U13605 (N_13605,N_13209,N_13237);
or U13606 (N_13606,N_13044,N_13004);
xnor U13607 (N_13607,N_13042,N_13295);
xnor U13608 (N_13608,N_13141,N_13099);
and U13609 (N_13609,N_13216,N_13473);
xnor U13610 (N_13610,N_13470,N_13117);
nand U13611 (N_13611,N_13226,N_13389);
nand U13612 (N_13612,N_13000,N_13220);
xnor U13613 (N_13613,N_13282,N_13302);
nand U13614 (N_13614,N_13426,N_13027);
or U13615 (N_13615,N_13022,N_13485);
nand U13616 (N_13616,N_13116,N_13080);
or U13617 (N_13617,N_13342,N_13332);
xnor U13618 (N_13618,N_13435,N_13387);
nor U13619 (N_13619,N_13093,N_13385);
nand U13620 (N_13620,N_13105,N_13376);
or U13621 (N_13621,N_13103,N_13277);
and U13622 (N_13622,N_13354,N_13110);
or U13623 (N_13623,N_13411,N_13043);
nor U13624 (N_13624,N_13305,N_13052);
nor U13625 (N_13625,N_13045,N_13440);
nand U13626 (N_13626,N_13121,N_13015);
nand U13627 (N_13627,N_13064,N_13281);
xnor U13628 (N_13628,N_13489,N_13014);
and U13629 (N_13629,N_13224,N_13055);
nor U13630 (N_13630,N_13085,N_13322);
xnor U13631 (N_13631,N_13268,N_13187);
nor U13632 (N_13632,N_13016,N_13456);
xor U13633 (N_13633,N_13242,N_13125);
xor U13634 (N_13634,N_13488,N_13192);
or U13635 (N_13635,N_13172,N_13371);
nand U13636 (N_13636,N_13091,N_13393);
and U13637 (N_13637,N_13213,N_13495);
and U13638 (N_13638,N_13296,N_13122);
or U13639 (N_13639,N_13194,N_13028);
or U13640 (N_13640,N_13072,N_13478);
and U13641 (N_13641,N_13088,N_13367);
nor U13642 (N_13642,N_13471,N_13171);
and U13643 (N_13643,N_13323,N_13089);
nand U13644 (N_13644,N_13388,N_13184);
xor U13645 (N_13645,N_13344,N_13267);
nor U13646 (N_13646,N_13156,N_13355);
or U13647 (N_13647,N_13462,N_13437);
nor U13648 (N_13648,N_13104,N_13217);
or U13649 (N_13649,N_13369,N_13030);
and U13650 (N_13650,N_13059,N_13203);
and U13651 (N_13651,N_13256,N_13076);
or U13652 (N_13652,N_13297,N_13174);
or U13653 (N_13653,N_13018,N_13465);
nand U13654 (N_13654,N_13496,N_13112);
nor U13655 (N_13655,N_13238,N_13357);
or U13656 (N_13656,N_13083,N_13005);
nor U13657 (N_13657,N_13033,N_13173);
or U13658 (N_13658,N_13299,N_13486);
and U13659 (N_13659,N_13461,N_13082);
or U13660 (N_13660,N_13269,N_13262);
nand U13661 (N_13661,N_13498,N_13400);
nand U13662 (N_13662,N_13392,N_13433);
and U13663 (N_13663,N_13038,N_13205);
or U13664 (N_13664,N_13115,N_13265);
nor U13665 (N_13665,N_13416,N_13041);
nor U13666 (N_13666,N_13200,N_13165);
or U13667 (N_13667,N_13407,N_13023);
xor U13668 (N_13668,N_13074,N_13170);
nand U13669 (N_13669,N_13275,N_13003);
nor U13670 (N_13670,N_13132,N_13423);
nand U13671 (N_13671,N_13126,N_13417);
nand U13672 (N_13672,N_13324,N_13477);
or U13673 (N_13673,N_13406,N_13049);
nor U13674 (N_13674,N_13143,N_13481);
nand U13675 (N_13675,N_13013,N_13336);
and U13676 (N_13676,N_13466,N_13012);
or U13677 (N_13677,N_13361,N_13233);
and U13678 (N_13678,N_13414,N_13398);
nor U13679 (N_13679,N_13090,N_13453);
and U13680 (N_13680,N_13283,N_13450);
xor U13681 (N_13681,N_13228,N_13443);
or U13682 (N_13682,N_13024,N_13148);
nand U13683 (N_13683,N_13384,N_13056);
nor U13684 (N_13684,N_13405,N_13439);
nor U13685 (N_13685,N_13154,N_13272);
xnor U13686 (N_13686,N_13247,N_13474);
nand U13687 (N_13687,N_13062,N_13308);
nand U13688 (N_13688,N_13051,N_13047);
nand U13689 (N_13689,N_13386,N_13075);
or U13690 (N_13690,N_13273,N_13087);
nand U13691 (N_13691,N_13424,N_13334);
nand U13692 (N_13692,N_13314,N_13312);
nor U13693 (N_13693,N_13067,N_13071);
and U13694 (N_13694,N_13135,N_13162);
nand U13695 (N_13695,N_13131,N_13218);
nor U13696 (N_13696,N_13413,N_13449);
or U13697 (N_13697,N_13383,N_13119);
xor U13698 (N_13698,N_13124,N_13078);
and U13699 (N_13699,N_13345,N_13136);
nand U13700 (N_13700,N_13182,N_13037);
nand U13701 (N_13701,N_13365,N_13292);
xnor U13702 (N_13702,N_13429,N_13123);
xor U13703 (N_13703,N_13098,N_13285);
nor U13704 (N_13704,N_13223,N_13331);
xor U13705 (N_13705,N_13235,N_13497);
nor U13706 (N_13706,N_13358,N_13329);
nor U13707 (N_13707,N_13151,N_13340);
nor U13708 (N_13708,N_13186,N_13202);
and U13709 (N_13709,N_13232,N_13222);
and U13710 (N_13710,N_13086,N_13279);
nor U13711 (N_13711,N_13107,N_13455);
nand U13712 (N_13712,N_13111,N_13252);
or U13713 (N_13713,N_13177,N_13364);
nor U13714 (N_13714,N_13472,N_13491);
nor U13715 (N_13715,N_13245,N_13097);
or U13716 (N_13716,N_13445,N_13139);
nand U13717 (N_13717,N_13035,N_13168);
and U13718 (N_13718,N_13438,N_13195);
nand U13719 (N_13719,N_13418,N_13328);
or U13720 (N_13720,N_13212,N_13026);
xnor U13721 (N_13721,N_13325,N_13454);
nand U13722 (N_13722,N_13330,N_13034);
nor U13723 (N_13723,N_13036,N_13101);
nor U13724 (N_13724,N_13396,N_13130);
or U13725 (N_13725,N_13366,N_13434);
nor U13726 (N_13726,N_13208,N_13248);
xnor U13727 (N_13727,N_13359,N_13293);
xnor U13728 (N_13728,N_13377,N_13128);
nor U13729 (N_13729,N_13457,N_13412);
and U13730 (N_13730,N_13244,N_13343);
or U13731 (N_13731,N_13032,N_13009);
xor U13732 (N_13732,N_13234,N_13249);
or U13733 (N_13733,N_13422,N_13257);
nor U13734 (N_13734,N_13431,N_13077);
nand U13735 (N_13735,N_13492,N_13375);
nand U13736 (N_13736,N_13335,N_13475);
xnor U13737 (N_13737,N_13403,N_13153);
xnor U13738 (N_13738,N_13278,N_13057);
nand U13739 (N_13739,N_13255,N_13161);
xor U13740 (N_13740,N_13061,N_13306);
or U13741 (N_13741,N_13144,N_13286);
nor U13742 (N_13742,N_13436,N_13053);
nand U13743 (N_13743,N_13048,N_13040);
and U13744 (N_13744,N_13315,N_13046);
xnor U13745 (N_13745,N_13317,N_13261);
nor U13746 (N_13746,N_13263,N_13303);
xnor U13747 (N_13747,N_13065,N_13225);
nor U13748 (N_13748,N_13029,N_13468);
xnor U13749 (N_13749,N_13253,N_13207);
nand U13750 (N_13750,N_13384,N_13223);
nand U13751 (N_13751,N_13227,N_13159);
and U13752 (N_13752,N_13204,N_13354);
or U13753 (N_13753,N_13056,N_13104);
or U13754 (N_13754,N_13409,N_13097);
and U13755 (N_13755,N_13156,N_13323);
nor U13756 (N_13756,N_13368,N_13239);
nor U13757 (N_13757,N_13253,N_13415);
and U13758 (N_13758,N_13246,N_13294);
or U13759 (N_13759,N_13001,N_13287);
and U13760 (N_13760,N_13130,N_13462);
or U13761 (N_13761,N_13026,N_13014);
nand U13762 (N_13762,N_13340,N_13444);
xnor U13763 (N_13763,N_13274,N_13053);
nor U13764 (N_13764,N_13325,N_13347);
and U13765 (N_13765,N_13493,N_13382);
or U13766 (N_13766,N_13279,N_13346);
nand U13767 (N_13767,N_13123,N_13048);
or U13768 (N_13768,N_13231,N_13173);
nand U13769 (N_13769,N_13070,N_13192);
xnor U13770 (N_13770,N_13148,N_13017);
xnor U13771 (N_13771,N_13037,N_13160);
nand U13772 (N_13772,N_13194,N_13376);
xnor U13773 (N_13773,N_13464,N_13195);
or U13774 (N_13774,N_13191,N_13238);
and U13775 (N_13775,N_13087,N_13260);
nand U13776 (N_13776,N_13073,N_13408);
and U13777 (N_13777,N_13247,N_13010);
nand U13778 (N_13778,N_13292,N_13353);
or U13779 (N_13779,N_13140,N_13110);
nand U13780 (N_13780,N_13232,N_13098);
nor U13781 (N_13781,N_13220,N_13016);
nor U13782 (N_13782,N_13008,N_13473);
nand U13783 (N_13783,N_13210,N_13078);
nor U13784 (N_13784,N_13009,N_13241);
nor U13785 (N_13785,N_13448,N_13246);
nand U13786 (N_13786,N_13252,N_13173);
nand U13787 (N_13787,N_13457,N_13024);
or U13788 (N_13788,N_13497,N_13384);
nor U13789 (N_13789,N_13154,N_13249);
nand U13790 (N_13790,N_13177,N_13266);
nor U13791 (N_13791,N_13452,N_13326);
or U13792 (N_13792,N_13302,N_13474);
nand U13793 (N_13793,N_13399,N_13294);
and U13794 (N_13794,N_13442,N_13176);
xor U13795 (N_13795,N_13391,N_13134);
and U13796 (N_13796,N_13047,N_13098);
nor U13797 (N_13797,N_13497,N_13029);
nor U13798 (N_13798,N_13039,N_13034);
nand U13799 (N_13799,N_13414,N_13202);
nand U13800 (N_13800,N_13011,N_13086);
or U13801 (N_13801,N_13081,N_13164);
nand U13802 (N_13802,N_13121,N_13098);
or U13803 (N_13803,N_13436,N_13276);
and U13804 (N_13804,N_13093,N_13432);
nand U13805 (N_13805,N_13191,N_13468);
xor U13806 (N_13806,N_13311,N_13175);
or U13807 (N_13807,N_13264,N_13139);
and U13808 (N_13808,N_13348,N_13132);
or U13809 (N_13809,N_13368,N_13480);
nand U13810 (N_13810,N_13162,N_13244);
nor U13811 (N_13811,N_13225,N_13381);
nand U13812 (N_13812,N_13083,N_13454);
or U13813 (N_13813,N_13369,N_13439);
nand U13814 (N_13814,N_13058,N_13155);
xor U13815 (N_13815,N_13175,N_13202);
and U13816 (N_13816,N_13439,N_13356);
and U13817 (N_13817,N_13010,N_13123);
or U13818 (N_13818,N_13485,N_13030);
nand U13819 (N_13819,N_13419,N_13253);
and U13820 (N_13820,N_13070,N_13015);
nor U13821 (N_13821,N_13336,N_13335);
or U13822 (N_13822,N_13476,N_13133);
or U13823 (N_13823,N_13272,N_13051);
and U13824 (N_13824,N_13139,N_13183);
xnor U13825 (N_13825,N_13050,N_13351);
xnor U13826 (N_13826,N_13344,N_13085);
nor U13827 (N_13827,N_13442,N_13317);
or U13828 (N_13828,N_13066,N_13447);
xnor U13829 (N_13829,N_13150,N_13233);
or U13830 (N_13830,N_13039,N_13158);
xor U13831 (N_13831,N_13129,N_13461);
or U13832 (N_13832,N_13017,N_13400);
xnor U13833 (N_13833,N_13078,N_13214);
or U13834 (N_13834,N_13110,N_13050);
xnor U13835 (N_13835,N_13216,N_13435);
nand U13836 (N_13836,N_13163,N_13045);
xnor U13837 (N_13837,N_13052,N_13340);
and U13838 (N_13838,N_13141,N_13040);
nor U13839 (N_13839,N_13035,N_13466);
xor U13840 (N_13840,N_13450,N_13135);
or U13841 (N_13841,N_13152,N_13260);
xnor U13842 (N_13842,N_13052,N_13369);
nor U13843 (N_13843,N_13260,N_13231);
nand U13844 (N_13844,N_13333,N_13415);
nand U13845 (N_13845,N_13051,N_13425);
nor U13846 (N_13846,N_13482,N_13172);
nand U13847 (N_13847,N_13138,N_13493);
xor U13848 (N_13848,N_13362,N_13162);
or U13849 (N_13849,N_13315,N_13099);
nor U13850 (N_13850,N_13385,N_13425);
xor U13851 (N_13851,N_13064,N_13383);
and U13852 (N_13852,N_13394,N_13035);
nor U13853 (N_13853,N_13218,N_13165);
and U13854 (N_13854,N_13430,N_13259);
nor U13855 (N_13855,N_13157,N_13113);
xor U13856 (N_13856,N_13021,N_13352);
nor U13857 (N_13857,N_13218,N_13446);
nor U13858 (N_13858,N_13183,N_13361);
xnor U13859 (N_13859,N_13472,N_13270);
nand U13860 (N_13860,N_13263,N_13248);
nor U13861 (N_13861,N_13233,N_13251);
or U13862 (N_13862,N_13277,N_13424);
nor U13863 (N_13863,N_13104,N_13482);
or U13864 (N_13864,N_13037,N_13354);
nand U13865 (N_13865,N_13217,N_13144);
nor U13866 (N_13866,N_13004,N_13395);
nand U13867 (N_13867,N_13422,N_13326);
nor U13868 (N_13868,N_13399,N_13453);
xor U13869 (N_13869,N_13149,N_13414);
nor U13870 (N_13870,N_13430,N_13350);
xor U13871 (N_13871,N_13468,N_13158);
nor U13872 (N_13872,N_13087,N_13182);
xor U13873 (N_13873,N_13429,N_13085);
nor U13874 (N_13874,N_13473,N_13242);
xor U13875 (N_13875,N_13438,N_13149);
xor U13876 (N_13876,N_13439,N_13220);
nor U13877 (N_13877,N_13285,N_13448);
nor U13878 (N_13878,N_13429,N_13118);
nor U13879 (N_13879,N_13202,N_13481);
or U13880 (N_13880,N_13165,N_13095);
and U13881 (N_13881,N_13265,N_13229);
nor U13882 (N_13882,N_13426,N_13407);
and U13883 (N_13883,N_13123,N_13155);
nand U13884 (N_13884,N_13282,N_13470);
xor U13885 (N_13885,N_13272,N_13171);
nor U13886 (N_13886,N_13161,N_13000);
or U13887 (N_13887,N_13156,N_13295);
nand U13888 (N_13888,N_13147,N_13357);
and U13889 (N_13889,N_13322,N_13301);
nand U13890 (N_13890,N_13413,N_13291);
xor U13891 (N_13891,N_13414,N_13477);
xnor U13892 (N_13892,N_13289,N_13135);
and U13893 (N_13893,N_13490,N_13435);
nand U13894 (N_13894,N_13261,N_13466);
or U13895 (N_13895,N_13279,N_13330);
nand U13896 (N_13896,N_13270,N_13217);
xnor U13897 (N_13897,N_13381,N_13401);
xnor U13898 (N_13898,N_13082,N_13356);
and U13899 (N_13899,N_13219,N_13003);
xnor U13900 (N_13900,N_13472,N_13136);
nor U13901 (N_13901,N_13259,N_13209);
nor U13902 (N_13902,N_13248,N_13002);
nor U13903 (N_13903,N_13400,N_13068);
nand U13904 (N_13904,N_13449,N_13069);
and U13905 (N_13905,N_13095,N_13034);
xor U13906 (N_13906,N_13263,N_13417);
or U13907 (N_13907,N_13282,N_13477);
and U13908 (N_13908,N_13162,N_13229);
or U13909 (N_13909,N_13292,N_13012);
or U13910 (N_13910,N_13151,N_13458);
nand U13911 (N_13911,N_13348,N_13166);
nor U13912 (N_13912,N_13008,N_13451);
or U13913 (N_13913,N_13411,N_13277);
xor U13914 (N_13914,N_13357,N_13483);
nor U13915 (N_13915,N_13458,N_13197);
nor U13916 (N_13916,N_13088,N_13174);
and U13917 (N_13917,N_13203,N_13497);
and U13918 (N_13918,N_13145,N_13389);
nand U13919 (N_13919,N_13224,N_13260);
nand U13920 (N_13920,N_13307,N_13404);
nor U13921 (N_13921,N_13096,N_13484);
xor U13922 (N_13922,N_13217,N_13319);
or U13923 (N_13923,N_13022,N_13010);
or U13924 (N_13924,N_13120,N_13378);
or U13925 (N_13925,N_13478,N_13468);
or U13926 (N_13926,N_13467,N_13381);
or U13927 (N_13927,N_13155,N_13219);
nor U13928 (N_13928,N_13483,N_13243);
or U13929 (N_13929,N_13336,N_13302);
nand U13930 (N_13930,N_13104,N_13013);
nor U13931 (N_13931,N_13010,N_13490);
nand U13932 (N_13932,N_13417,N_13284);
nor U13933 (N_13933,N_13320,N_13248);
or U13934 (N_13934,N_13471,N_13214);
nor U13935 (N_13935,N_13310,N_13102);
and U13936 (N_13936,N_13275,N_13188);
nand U13937 (N_13937,N_13109,N_13280);
nor U13938 (N_13938,N_13399,N_13301);
or U13939 (N_13939,N_13419,N_13272);
xnor U13940 (N_13940,N_13463,N_13108);
nand U13941 (N_13941,N_13191,N_13362);
or U13942 (N_13942,N_13208,N_13032);
or U13943 (N_13943,N_13366,N_13111);
or U13944 (N_13944,N_13097,N_13372);
and U13945 (N_13945,N_13360,N_13446);
nand U13946 (N_13946,N_13048,N_13386);
and U13947 (N_13947,N_13464,N_13441);
or U13948 (N_13948,N_13356,N_13408);
or U13949 (N_13949,N_13050,N_13209);
nand U13950 (N_13950,N_13155,N_13117);
nand U13951 (N_13951,N_13243,N_13314);
xnor U13952 (N_13952,N_13499,N_13416);
nor U13953 (N_13953,N_13375,N_13070);
or U13954 (N_13954,N_13404,N_13064);
xor U13955 (N_13955,N_13338,N_13161);
and U13956 (N_13956,N_13246,N_13442);
xor U13957 (N_13957,N_13095,N_13090);
nor U13958 (N_13958,N_13180,N_13269);
nor U13959 (N_13959,N_13280,N_13032);
and U13960 (N_13960,N_13050,N_13135);
xnor U13961 (N_13961,N_13053,N_13109);
xnor U13962 (N_13962,N_13422,N_13256);
nand U13963 (N_13963,N_13320,N_13014);
nand U13964 (N_13964,N_13258,N_13083);
or U13965 (N_13965,N_13444,N_13029);
nor U13966 (N_13966,N_13273,N_13079);
or U13967 (N_13967,N_13236,N_13217);
nand U13968 (N_13968,N_13469,N_13296);
nor U13969 (N_13969,N_13266,N_13433);
nand U13970 (N_13970,N_13091,N_13074);
nor U13971 (N_13971,N_13020,N_13193);
xnor U13972 (N_13972,N_13007,N_13027);
nand U13973 (N_13973,N_13430,N_13485);
and U13974 (N_13974,N_13179,N_13055);
or U13975 (N_13975,N_13344,N_13465);
or U13976 (N_13976,N_13204,N_13232);
or U13977 (N_13977,N_13404,N_13168);
nor U13978 (N_13978,N_13435,N_13334);
nand U13979 (N_13979,N_13072,N_13053);
and U13980 (N_13980,N_13434,N_13025);
nand U13981 (N_13981,N_13168,N_13233);
xnor U13982 (N_13982,N_13292,N_13396);
and U13983 (N_13983,N_13024,N_13497);
xor U13984 (N_13984,N_13381,N_13349);
or U13985 (N_13985,N_13403,N_13110);
xnor U13986 (N_13986,N_13049,N_13414);
xnor U13987 (N_13987,N_13028,N_13100);
nand U13988 (N_13988,N_13377,N_13354);
xnor U13989 (N_13989,N_13430,N_13314);
nor U13990 (N_13990,N_13127,N_13190);
and U13991 (N_13991,N_13474,N_13401);
nand U13992 (N_13992,N_13136,N_13271);
nor U13993 (N_13993,N_13206,N_13447);
xnor U13994 (N_13994,N_13213,N_13255);
xnor U13995 (N_13995,N_13467,N_13002);
nor U13996 (N_13996,N_13003,N_13205);
or U13997 (N_13997,N_13454,N_13082);
and U13998 (N_13998,N_13433,N_13127);
nor U13999 (N_13999,N_13216,N_13332);
nand U14000 (N_14000,N_13641,N_13690);
or U14001 (N_14001,N_13979,N_13817);
or U14002 (N_14002,N_13624,N_13598);
and U14003 (N_14003,N_13737,N_13844);
nor U14004 (N_14004,N_13961,N_13813);
and U14005 (N_14005,N_13509,N_13670);
xor U14006 (N_14006,N_13889,N_13604);
nand U14007 (N_14007,N_13526,N_13619);
nand U14008 (N_14008,N_13674,N_13689);
nor U14009 (N_14009,N_13822,N_13995);
or U14010 (N_14010,N_13515,N_13934);
nand U14011 (N_14011,N_13643,N_13572);
nor U14012 (N_14012,N_13603,N_13880);
nand U14013 (N_14013,N_13917,N_13649);
nor U14014 (N_14014,N_13591,N_13857);
or U14015 (N_14015,N_13521,N_13790);
xor U14016 (N_14016,N_13673,N_13658);
nor U14017 (N_14017,N_13664,N_13660);
or U14018 (N_14018,N_13721,N_13996);
or U14019 (N_14019,N_13640,N_13621);
and U14020 (N_14020,N_13590,N_13759);
xor U14021 (N_14021,N_13628,N_13545);
xnor U14022 (N_14022,N_13778,N_13744);
xor U14023 (N_14023,N_13748,N_13648);
nand U14024 (N_14024,N_13559,N_13907);
nand U14025 (N_14025,N_13529,N_13717);
and U14026 (N_14026,N_13718,N_13579);
nor U14027 (N_14027,N_13825,N_13903);
nor U14028 (N_14028,N_13663,N_13882);
or U14029 (N_14029,N_13945,N_13588);
and U14030 (N_14030,N_13821,N_13766);
nand U14031 (N_14031,N_13676,N_13706);
nor U14032 (N_14032,N_13781,N_13806);
nor U14033 (N_14033,N_13680,N_13966);
nor U14034 (N_14034,N_13523,N_13539);
or U14035 (N_14035,N_13682,N_13876);
and U14036 (N_14036,N_13738,N_13926);
nor U14037 (N_14037,N_13727,N_13542);
xnor U14038 (N_14038,N_13988,N_13511);
xor U14039 (N_14039,N_13911,N_13575);
nor U14040 (N_14040,N_13853,N_13839);
nand U14041 (N_14041,N_13623,N_13816);
and U14042 (N_14042,N_13700,N_13894);
and U14043 (N_14043,N_13524,N_13634);
or U14044 (N_14044,N_13855,N_13602);
nand U14045 (N_14045,N_13600,N_13993);
nand U14046 (N_14046,N_13667,N_13863);
and U14047 (N_14047,N_13779,N_13789);
or U14048 (N_14048,N_13609,N_13708);
and U14049 (N_14049,N_13973,N_13848);
nor U14050 (N_14050,N_13638,N_13944);
and U14051 (N_14051,N_13586,N_13841);
nand U14052 (N_14052,N_13583,N_13653);
and U14053 (N_14053,N_13796,N_13842);
xor U14054 (N_14054,N_13878,N_13845);
xnor U14055 (N_14055,N_13512,N_13750);
nor U14056 (N_14056,N_13998,N_13981);
nor U14057 (N_14057,N_13893,N_13686);
or U14058 (N_14058,N_13854,N_13608);
xor U14059 (N_14059,N_13895,N_13508);
xnor U14060 (N_14060,N_13942,N_13935);
or U14061 (N_14061,N_13525,N_13518);
nand U14062 (N_14062,N_13601,N_13709);
nor U14063 (N_14063,N_13930,N_13976);
or U14064 (N_14064,N_13777,N_13818);
or U14065 (N_14065,N_13954,N_13832);
nor U14066 (N_14066,N_13991,N_13540);
xnor U14067 (N_14067,N_13587,N_13885);
and U14068 (N_14068,N_13571,N_13868);
or U14069 (N_14069,N_13925,N_13932);
or U14070 (N_14070,N_13666,N_13705);
nor U14071 (N_14071,N_13910,N_13929);
xnor U14072 (N_14072,N_13951,N_13560);
or U14073 (N_14073,N_13754,N_13888);
nand U14074 (N_14074,N_13793,N_13782);
or U14075 (N_14075,N_13537,N_13724);
xnor U14076 (N_14076,N_13612,N_13859);
nor U14077 (N_14077,N_13568,N_13768);
and U14078 (N_14078,N_13558,N_13714);
nor U14079 (N_14079,N_13772,N_13740);
nand U14080 (N_14080,N_13651,N_13865);
or U14081 (N_14081,N_13804,N_13760);
and U14082 (N_14082,N_13985,N_13574);
or U14083 (N_14083,N_13616,N_13656);
or U14084 (N_14084,N_13513,N_13968);
xnor U14085 (N_14085,N_13502,N_13928);
or U14086 (N_14086,N_13869,N_13629);
nand U14087 (N_14087,N_13742,N_13639);
or U14088 (N_14088,N_13946,N_13803);
nor U14089 (N_14089,N_13688,N_13982);
nand U14090 (N_14090,N_13522,N_13884);
nor U14091 (N_14091,N_13916,N_13657);
xor U14092 (N_14092,N_13546,N_13983);
nor U14093 (N_14093,N_13831,N_13729);
nand U14094 (N_14094,N_13684,N_13655);
xor U14095 (N_14095,N_13899,N_13947);
nand U14096 (N_14096,N_13883,N_13549);
nor U14097 (N_14097,N_13570,N_13711);
or U14098 (N_14098,N_13798,N_13728);
xnor U14099 (N_14099,N_13987,N_13920);
or U14100 (N_14100,N_13720,N_13683);
xnor U14101 (N_14101,N_13918,N_13891);
nand U14102 (N_14102,N_13584,N_13722);
nor U14103 (N_14103,N_13758,N_13791);
xor U14104 (N_14104,N_13696,N_13541);
nand U14105 (N_14105,N_13678,N_13715);
nand U14106 (N_14106,N_13902,N_13900);
xor U14107 (N_14107,N_13703,N_13784);
and U14108 (N_14108,N_13610,N_13811);
and U14109 (N_14109,N_13501,N_13555);
and U14110 (N_14110,N_13593,N_13685);
nor U14111 (N_14111,N_13662,N_13625);
or U14112 (N_14112,N_13636,N_13956);
nand U14113 (N_14113,N_13828,N_13719);
xor U14114 (N_14114,N_13736,N_13805);
nor U14115 (N_14115,N_13861,N_13978);
nor U14116 (N_14116,N_13800,N_13971);
and U14117 (N_14117,N_13815,N_13614);
nand U14118 (N_14118,N_13516,N_13536);
nor U14119 (N_14119,N_13553,N_13573);
or U14120 (N_14120,N_13972,N_13810);
or U14121 (N_14121,N_13989,N_13617);
and U14122 (N_14122,N_13637,N_13746);
nand U14123 (N_14123,N_13723,N_13699);
or U14124 (N_14124,N_13654,N_13826);
nand U14125 (N_14125,N_13792,N_13783);
xnor U14126 (N_14126,N_13950,N_13892);
xnor U14127 (N_14127,N_13531,N_13802);
nor U14128 (N_14128,N_13952,N_13829);
or U14129 (N_14129,N_13730,N_13770);
nor U14130 (N_14130,N_13974,N_13589);
nor U14131 (N_14131,N_13836,N_13970);
xnor U14132 (N_14132,N_13901,N_13812);
and U14133 (N_14133,N_13922,N_13999);
nor U14134 (N_14134,N_13733,N_13938);
xor U14135 (N_14135,N_13533,N_13615);
and U14136 (N_14136,N_13780,N_13906);
xor U14137 (N_14137,N_13503,N_13940);
nand U14138 (N_14138,N_13606,N_13618);
xor U14139 (N_14139,N_13691,N_13967);
xor U14140 (N_14140,N_13843,N_13599);
nor U14141 (N_14141,N_13924,N_13771);
nand U14142 (N_14142,N_13908,N_13626);
nor U14143 (N_14143,N_13692,N_13607);
nor U14144 (N_14144,N_13550,N_13679);
and U14145 (N_14145,N_13795,N_13646);
xnor U14146 (N_14146,N_13786,N_13990);
and U14147 (N_14147,N_13927,N_13847);
nand U14148 (N_14148,N_13915,N_13919);
nand U14149 (N_14149,N_13797,N_13630);
nor U14150 (N_14150,N_13677,N_13694);
and U14151 (N_14151,N_13527,N_13544);
or U14152 (N_14152,N_13814,N_13704);
nor U14153 (N_14153,N_13563,N_13548);
nand U14154 (N_14154,N_13994,N_13962);
xor U14155 (N_14155,N_13931,N_13505);
nand U14156 (N_14156,N_13933,N_13941);
or U14157 (N_14157,N_13774,N_13776);
and U14158 (N_14158,N_13734,N_13867);
and U14159 (N_14159,N_13631,N_13862);
or U14160 (N_14160,N_13870,N_13898);
and U14161 (N_14161,N_13528,N_13939);
nor U14162 (N_14162,N_13581,N_13948);
or U14163 (N_14163,N_13785,N_13534);
xnor U14164 (N_14164,N_13960,N_13578);
and U14165 (N_14165,N_13823,N_13735);
or U14166 (N_14166,N_13596,N_13824);
xnor U14167 (N_14167,N_13788,N_13852);
xnor U14168 (N_14168,N_13984,N_13794);
and U14169 (N_14169,N_13672,N_13535);
xnor U14170 (N_14170,N_13840,N_13731);
xnor U14171 (N_14171,N_13500,N_13712);
nor U14172 (N_14172,N_13890,N_13661);
nand U14173 (N_14173,N_13977,N_13873);
nor U14174 (N_14174,N_13665,N_13532);
or U14175 (N_14175,N_13507,N_13547);
nor U14176 (N_14176,N_13773,N_13846);
and U14177 (N_14177,N_13580,N_13702);
or U14178 (N_14178,N_13992,N_13921);
or U14179 (N_14179,N_13605,N_13755);
or U14180 (N_14180,N_13556,N_13576);
or U14181 (N_14181,N_13504,N_13752);
nand U14182 (N_14182,N_13567,N_13959);
and U14183 (N_14183,N_13799,N_13613);
nor U14184 (N_14184,N_13896,N_13582);
nor U14185 (N_14185,N_13749,N_13936);
nand U14186 (N_14186,N_13937,N_13675);
and U14187 (N_14187,N_13732,N_13904);
and U14188 (N_14188,N_13695,N_13986);
nor U14189 (N_14189,N_13969,N_13762);
and U14190 (N_14190,N_13949,N_13808);
and U14191 (N_14191,N_13963,N_13850);
or U14192 (N_14192,N_13765,N_13764);
and U14193 (N_14193,N_13726,N_13801);
and U14194 (N_14194,N_13860,N_13851);
nor U14195 (N_14195,N_13632,N_13520);
nand U14196 (N_14196,N_13997,N_13964);
nand U14197 (N_14197,N_13566,N_13569);
and U14198 (N_14198,N_13538,N_13652);
nor U14199 (N_14199,N_13807,N_13953);
nor U14200 (N_14200,N_13592,N_13597);
nor U14201 (N_14201,N_13725,N_13943);
xor U14202 (N_14202,N_13769,N_13757);
nand U14203 (N_14203,N_13905,N_13879);
nand U14204 (N_14204,N_13872,N_13669);
xor U14205 (N_14205,N_13698,N_13835);
or U14206 (N_14206,N_13681,N_13633);
or U14207 (N_14207,N_13787,N_13647);
xnor U14208 (N_14208,N_13693,N_13761);
nor U14209 (N_14209,N_13595,N_13965);
nand U14210 (N_14210,N_13517,N_13849);
nand U14211 (N_14211,N_13611,N_13552);
or U14212 (N_14212,N_13886,N_13697);
nor U14213 (N_14213,N_13775,N_13627);
or U14214 (N_14214,N_13912,N_13833);
and U14215 (N_14215,N_13875,N_13510);
xor U14216 (N_14216,N_13741,N_13756);
or U14217 (N_14217,N_13557,N_13881);
or U14218 (N_14218,N_13622,N_13659);
nand U14219 (N_14219,N_13747,N_13864);
and U14220 (N_14220,N_13763,N_13564);
xor U14221 (N_14221,N_13519,N_13650);
nor U14222 (N_14222,N_13620,N_13980);
xnor U14223 (N_14223,N_13745,N_13909);
or U14224 (N_14224,N_13585,N_13838);
xnor U14225 (N_14225,N_13957,N_13561);
nor U14226 (N_14226,N_13887,N_13858);
nand U14227 (N_14227,N_13837,N_13753);
and U14228 (N_14228,N_13687,N_13897);
nand U14229 (N_14229,N_13743,N_13819);
nor U14230 (N_14230,N_13767,N_13739);
xor U14231 (N_14231,N_13874,N_13577);
nand U14232 (N_14232,N_13671,N_13551);
xnor U14233 (N_14233,N_13856,N_13644);
or U14234 (N_14234,N_13975,N_13594);
and U14235 (N_14235,N_13830,N_13820);
and U14236 (N_14236,N_13827,N_13834);
and U14237 (N_14237,N_13543,N_13707);
or U14238 (N_14238,N_13562,N_13871);
xor U14239 (N_14239,N_13877,N_13506);
xnor U14240 (N_14240,N_13716,N_13668);
or U14241 (N_14241,N_13635,N_13955);
and U14242 (N_14242,N_13958,N_13642);
or U14243 (N_14243,N_13751,N_13913);
or U14244 (N_14244,N_13914,N_13701);
and U14245 (N_14245,N_13710,N_13514);
nor U14246 (N_14246,N_13866,N_13923);
or U14247 (N_14247,N_13530,N_13554);
or U14248 (N_14248,N_13565,N_13809);
xnor U14249 (N_14249,N_13645,N_13713);
and U14250 (N_14250,N_13615,N_13648);
or U14251 (N_14251,N_13682,N_13595);
nor U14252 (N_14252,N_13930,N_13767);
nor U14253 (N_14253,N_13549,N_13662);
nand U14254 (N_14254,N_13802,N_13575);
and U14255 (N_14255,N_13967,N_13785);
xnor U14256 (N_14256,N_13586,N_13531);
nand U14257 (N_14257,N_13526,N_13611);
nor U14258 (N_14258,N_13832,N_13726);
xor U14259 (N_14259,N_13904,N_13940);
or U14260 (N_14260,N_13617,N_13697);
or U14261 (N_14261,N_13852,N_13967);
and U14262 (N_14262,N_13799,N_13617);
xnor U14263 (N_14263,N_13979,N_13553);
xor U14264 (N_14264,N_13959,N_13698);
nor U14265 (N_14265,N_13958,N_13937);
and U14266 (N_14266,N_13904,N_13512);
nand U14267 (N_14267,N_13730,N_13831);
xnor U14268 (N_14268,N_13896,N_13731);
xnor U14269 (N_14269,N_13607,N_13536);
or U14270 (N_14270,N_13934,N_13513);
nor U14271 (N_14271,N_13990,N_13731);
nor U14272 (N_14272,N_13688,N_13713);
and U14273 (N_14273,N_13852,N_13616);
or U14274 (N_14274,N_13566,N_13848);
xor U14275 (N_14275,N_13798,N_13974);
nor U14276 (N_14276,N_13924,N_13633);
nor U14277 (N_14277,N_13548,N_13818);
and U14278 (N_14278,N_13976,N_13856);
or U14279 (N_14279,N_13543,N_13768);
or U14280 (N_14280,N_13775,N_13997);
or U14281 (N_14281,N_13813,N_13911);
or U14282 (N_14282,N_13504,N_13892);
and U14283 (N_14283,N_13817,N_13583);
or U14284 (N_14284,N_13577,N_13960);
and U14285 (N_14285,N_13957,N_13923);
nor U14286 (N_14286,N_13551,N_13731);
and U14287 (N_14287,N_13981,N_13983);
and U14288 (N_14288,N_13729,N_13965);
or U14289 (N_14289,N_13827,N_13566);
or U14290 (N_14290,N_13568,N_13573);
and U14291 (N_14291,N_13981,N_13554);
nand U14292 (N_14292,N_13855,N_13930);
or U14293 (N_14293,N_13724,N_13656);
and U14294 (N_14294,N_13708,N_13635);
nor U14295 (N_14295,N_13562,N_13624);
nor U14296 (N_14296,N_13734,N_13686);
xor U14297 (N_14297,N_13994,N_13886);
nor U14298 (N_14298,N_13964,N_13691);
nand U14299 (N_14299,N_13654,N_13940);
nand U14300 (N_14300,N_13794,N_13538);
nor U14301 (N_14301,N_13798,N_13895);
xor U14302 (N_14302,N_13781,N_13699);
and U14303 (N_14303,N_13733,N_13744);
and U14304 (N_14304,N_13997,N_13988);
or U14305 (N_14305,N_13656,N_13756);
xnor U14306 (N_14306,N_13885,N_13828);
nand U14307 (N_14307,N_13824,N_13506);
xor U14308 (N_14308,N_13528,N_13601);
nand U14309 (N_14309,N_13764,N_13921);
and U14310 (N_14310,N_13861,N_13954);
nor U14311 (N_14311,N_13697,N_13694);
xnor U14312 (N_14312,N_13865,N_13563);
or U14313 (N_14313,N_13904,N_13803);
nand U14314 (N_14314,N_13973,N_13643);
and U14315 (N_14315,N_13909,N_13807);
or U14316 (N_14316,N_13957,N_13662);
nor U14317 (N_14317,N_13842,N_13739);
nor U14318 (N_14318,N_13908,N_13516);
xor U14319 (N_14319,N_13981,N_13967);
and U14320 (N_14320,N_13710,N_13757);
nand U14321 (N_14321,N_13557,N_13697);
nor U14322 (N_14322,N_13600,N_13778);
and U14323 (N_14323,N_13736,N_13532);
and U14324 (N_14324,N_13867,N_13588);
nor U14325 (N_14325,N_13541,N_13767);
xor U14326 (N_14326,N_13727,N_13636);
and U14327 (N_14327,N_13749,N_13748);
nor U14328 (N_14328,N_13759,N_13935);
or U14329 (N_14329,N_13943,N_13917);
nand U14330 (N_14330,N_13660,N_13662);
xor U14331 (N_14331,N_13835,N_13514);
xnor U14332 (N_14332,N_13579,N_13917);
xnor U14333 (N_14333,N_13792,N_13734);
or U14334 (N_14334,N_13841,N_13703);
nor U14335 (N_14335,N_13719,N_13851);
nand U14336 (N_14336,N_13736,N_13759);
or U14337 (N_14337,N_13640,N_13986);
nor U14338 (N_14338,N_13557,N_13977);
xor U14339 (N_14339,N_13753,N_13925);
and U14340 (N_14340,N_13955,N_13611);
or U14341 (N_14341,N_13739,N_13768);
nand U14342 (N_14342,N_13693,N_13930);
and U14343 (N_14343,N_13504,N_13578);
xnor U14344 (N_14344,N_13532,N_13776);
nand U14345 (N_14345,N_13954,N_13982);
xor U14346 (N_14346,N_13617,N_13841);
nand U14347 (N_14347,N_13677,N_13549);
nor U14348 (N_14348,N_13959,N_13911);
and U14349 (N_14349,N_13561,N_13916);
and U14350 (N_14350,N_13707,N_13961);
nand U14351 (N_14351,N_13807,N_13887);
nand U14352 (N_14352,N_13924,N_13500);
nor U14353 (N_14353,N_13746,N_13980);
nor U14354 (N_14354,N_13697,N_13676);
nor U14355 (N_14355,N_13770,N_13925);
xor U14356 (N_14356,N_13586,N_13877);
or U14357 (N_14357,N_13672,N_13865);
and U14358 (N_14358,N_13785,N_13806);
nor U14359 (N_14359,N_13544,N_13505);
or U14360 (N_14360,N_13680,N_13587);
or U14361 (N_14361,N_13581,N_13556);
or U14362 (N_14362,N_13831,N_13904);
nor U14363 (N_14363,N_13675,N_13736);
xor U14364 (N_14364,N_13659,N_13575);
nand U14365 (N_14365,N_13697,N_13562);
nor U14366 (N_14366,N_13514,N_13945);
xnor U14367 (N_14367,N_13604,N_13735);
nand U14368 (N_14368,N_13520,N_13691);
nand U14369 (N_14369,N_13510,N_13857);
nand U14370 (N_14370,N_13661,N_13600);
or U14371 (N_14371,N_13818,N_13866);
or U14372 (N_14372,N_13933,N_13563);
nand U14373 (N_14373,N_13871,N_13727);
xnor U14374 (N_14374,N_13868,N_13662);
nand U14375 (N_14375,N_13779,N_13709);
or U14376 (N_14376,N_13505,N_13890);
and U14377 (N_14377,N_13749,N_13590);
nor U14378 (N_14378,N_13661,N_13873);
or U14379 (N_14379,N_13869,N_13849);
xor U14380 (N_14380,N_13654,N_13555);
nor U14381 (N_14381,N_13927,N_13909);
or U14382 (N_14382,N_13959,N_13785);
and U14383 (N_14383,N_13738,N_13973);
and U14384 (N_14384,N_13773,N_13888);
xor U14385 (N_14385,N_13572,N_13548);
or U14386 (N_14386,N_13987,N_13918);
xnor U14387 (N_14387,N_13817,N_13667);
xnor U14388 (N_14388,N_13926,N_13649);
nor U14389 (N_14389,N_13538,N_13895);
xnor U14390 (N_14390,N_13936,N_13698);
nor U14391 (N_14391,N_13916,N_13726);
or U14392 (N_14392,N_13769,N_13594);
nor U14393 (N_14393,N_13782,N_13678);
xor U14394 (N_14394,N_13847,N_13979);
nand U14395 (N_14395,N_13961,N_13692);
nor U14396 (N_14396,N_13610,N_13960);
xnor U14397 (N_14397,N_13982,N_13578);
and U14398 (N_14398,N_13666,N_13956);
nor U14399 (N_14399,N_13669,N_13705);
xnor U14400 (N_14400,N_13974,N_13562);
or U14401 (N_14401,N_13817,N_13932);
and U14402 (N_14402,N_13507,N_13694);
nor U14403 (N_14403,N_13935,N_13993);
and U14404 (N_14404,N_13665,N_13909);
nand U14405 (N_14405,N_13886,N_13653);
nor U14406 (N_14406,N_13811,N_13612);
and U14407 (N_14407,N_13595,N_13772);
and U14408 (N_14408,N_13818,N_13981);
and U14409 (N_14409,N_13844,N_13559);
nand U14410 (N_14410,N_13770,N_13958);
and U14411 (N_14411,N_13892,N_13833);
and U14412 (N_14412,N_13533,N_13535);
nor U14413 (N_14413,N_13935,N_13906);
and U14414 (N_14414,N_13891,N_13763);
nand U14415 (N_14415,N_13641,N_13640);
xnor U14416 (N_14416,N_13721,N_13738);
and U14417 (N_14417,N_13621,N_13822);
nand U14418 (N_14418,N_13529,N_13715);
and U14419 (N_14419,N_13770,N_13525);
nand U14420 (N_14420,N_13631,N_13558);
nand U14421 (N_14421,N_13951,N_13866);
or U14422 (N_14422,N_13839,N_13948);
nor U14423 (N_14423,N_13828,N_13820);
or U14424 (N_14424,N_13651,N_13646);
or U14425 (N_14425,N_13785,N_13866);
nor U14426 (N_14426,N_13599,N_13888);
nor U14427 (N_14427,N_13560,N_13814);
xnor U14428 (N_14428,N_13977,N_13771);
and U14429 (N_14429,N_13978,N_13638);
nor U14430 (N_14430,N_13659,N_13516);
nand U14431 (N_14431,N_13980,N_13538);
or U14432 (N_14432,N_13869,N_13766);
nand U14433 (N_14433,N_13944,N_13505);
nand U14434 (N_14434,N_13887,N_13688);
and U14435 (N_14435,N_13610,N_13608);
and U14436 (N_14436,N_13881,N_13713);
or U14437 (N_14437,N_13987,N_13813);
nor U14438 (N_14438,N_13554,N_13609);
and U14439 (N_14439,N_13624,N_13828);
nor U14440 (N_14440,N_13692,N_13506);
and U14441 (N_14441,N_13639,N_13703);
xor U14442 (N_14442,N_13588,N_13652);
or U14443 (N_14443,N_13984,N_13942);
nand U14444 (N_14444,N_13925,N_13569);
nor U14445 (N_14445,N_13777,N_13909);
or U14446 (N_14446,N_13853,N_13772);
nor U14447 (N_14447,N_13501,N_13637);
or U14448 (N_14448,N_13746,N_13711);
xnor U14449 (N_14449,N_13769,N_13776);
nand U14450 (N_14450,N_13981,N_13533);
nor U14451 (N_14451,N_13932,N_13709);
nand U14452 (N_14452,N_13870,N_13588);
nand U14453 (N_14453,N_13884,N_13611);
nor U14454 (N_14454,N_13581,N_13923);
nor U14455 (N_14455,N_13917,N_13916);
nor U14456 (N_14456,N_13896,N_13753);
or U14457 (N_14457,N_13984,N_13922);
xnor U14458 (N_14458,N_13885,N_13913);
nand U14459 (N_14459,N_13743,N_13515);
nand U14460 (N_14460,N_13578,N_13587);
nand U14461 (N_14461,N_13811,N_13734);
xor U14462 (N_14462,N_13801,N_13566);
and U14463 (N_14463,N_13508,N_13946);
xor U14464 (N_14464,N_13840,N_13711);
and U14465 (N_14465,N_13931,N_13854);
and U14466 (N_14466,N_13752,N_13695);
and U14467 (N_14467,N_13638,N_13883);
and U14468 (N_14468,N_13733,N_13550);
or U14469 (N_14469,N_13818,N_13625);
and U14470 (N_14470,N_13708,N_13522);
nor U14471 (N_14471,N_13919,N_13957);
xnor U14472 (N_14472,N_13667,N_13947);
nor U14473 (N_14473,N_13760,N_13960);
or U14474 (N_14474,N_13976,N_13725);
or U14475 (N_14475,N_13855,N_13551);
or U14476 (N_14476,N_13855,N_13728);
nand U14477 (N_14477,N_13857,N_13994);
nor U14478 (N_14478,N_13556,N_13615);
xnor U14479 (N_14479,N_13921,N_13990);
nor U14480 (N_14480,N_13648,N_13684);
and U14481 (N_14481,N_13579,N_13852);
nand U14482 (N_14482,N_13629,N_13783);
xnor U14483 (N_14483,N_13812,N_13735);
nand U14484 (N_14484,N_13507,N_13599);
xnor U14485 (N_14485,N_13652,N_13610);
or U14486 (N_14486,N_13984,N_13925);
nand U14487 (N_14487,N_13550,N_13753);
xnor U14488 (N_14488,N_13716,N_13705);
or U14489 (N_14489,N_13716,N_13902);
xnor U14490 (N_14490,N_13838,N_13653);
nor U14491 (N_14491,N_13700,N_13842);
nand U14492 (N_14492,N_13738,N_13658);
nand U14493 (N_14493,N_13826,N_13995);
and U14494 (N_14494,N_13822,N_13954);
xor U14495 (N_14495,N_13818,N_13572);
or U14496 (N_14496,N_13883,N_13932);
nand U14497 (N_14497,N_13741,N_13641);
nand U14498 (N_14498,N_13858,N_13717);
or U14499 (N_14499,N_13964,N_13665);
nor U14500 (N_14500,N_14102,N_14314);
xnor U14501 (N_14501,N_14275,N_14341);
or U14502 (N_14502,N_14016,N_14020);
nor U14503 (N_14503,N_14088,N_14045);
xor U14504 (N_14504,N_14445,N_14465);
and U14505 (N_14505,N_14343,N_14018);
and U14506 (N_14506,N_14210,N_14139);
xnor U14507 (N_14507,N_14048,N_14281);
or U14508 (N_14508,N_14359,N_14134);
nor U14509 (N_14509,N_14356,N_14234);
nand U14510 (N_14510,N_14253,N_14093);
and U14511 (N_14511,N_14410,N_14217);
and U14512 (N_14512,N_14489,N_14418);
xor U14513 (N_14513,N_14366,N_14317);
or U14514 (N_14514,N_14362,N_14334);
and U14515 (N_14515,N_14125,N_14376);
nand U14516 (N_14516,N_14447,N_14474);
or U14517 (N_14517,N_14196,N_14370);
or U14518 (N_14518,N_14326,N_14029);
nand U14519 (N_14519,N_14254,N_14215);
nand U14520 (N_14520,N_14096,N_14014);
or U14521 (N_14521,N_14371,N_14060);
xor U14522 (N_14522,N_14319,N_14122);
and U14523 (N_14523,N_14218,N_14170);
nand U14524 (N_14524,N_14069,N_14034);
or U14525 (N_14525,N_14167,N_14270);
or U14526 (N_14526,N_14479,N_14041);
or U14527 (N_14527,N_14394,N_14100);
nor U14528 (N_14528,N_14459,N_14178);
and U14529 (N_14529,N_14432,N_14222);
or U14530 (N_14530,N_14420,N_14345);
xor U14531 (N_14531,N_14415,N_14441);
and U14532 (N_14532,N_14409,N_14193);
nand U14533 (N_14533,N_14309,N_14203);
xnor U14534 (N_14534,N_14119,N_14239);
nor U14535 (N_14535,N_14230,N_14017);
nor U14536 (N_14536,N_14220,N_14351);
nand U14537 (N_14537,N_14276,N_14400);
xor U14538 (N_14538,N_14397,N_14083);
or U14539 (N_14539,N_14169,N_14171);
or U14540 (N_14540,N_14392,N_14427);
and U14541 (N_14541,N_14201,N_14130);
or U14542 (N_14542,N_14472,N_14111);
or U14543 (N_14543,N_14377,N_14492);
nor U14544 (N_14544,N_14338,N_14259);
and U14545 (N_14545,N_14464,N_14227);
or U14546 (N_14546,N_14375,N_14223);
and U14547 (N_14547,N_14293,N_14488);
or U14548 (N_14548,N_14142,N_14145);
and U14549 (N_14549,N_14063,N_14274);
or U14550 (N_14550,N_14398,N_14114);
nand U14551 (N_14551,N_14391,N_14112);
nor U14552 (N_14552,N_14312,N_14085);
and U14553 (N_14553,N_14135,N_14342);
or U14554 (N_14554,N_14458,N_14174);
xor U14555 (N_14555,N_14204,N_14187);
nand U14556 (N_14556,N_14363,N_14473);
nand U14557 (N_14557,N_14067,N_14129);
nor U14558 (N_14558,N_14156,N_14221);
xnor U14559 (N_14559,N_14148,N_14089);
nand U14560 (N_14560,N_14225,N_14015);
and U14561 (N_14561,N_14138,N_14168);
or U14562 (N_14562,N_14298,N_14010);
or U14563 (N_14563,N_14353,N_14261);
nor U14564 (N_14564,N_14143,N_14283);
and U14565 (N_14565,N_14315,N_14277);
nand U14566 (N_14566,N_14379,N_14497);
nand U14567 (N_14567,N_14411,N_14477);
nor U14568 (N_14568,N_14146,N_14381);
nand U14569 (N_14569,N_14327,N_14491);
xnor U14570 (N_14570,N_14357,N_14296);
and U14571 (N_14571,N_14158,N_14213);
or U14572 (N_14572,N_14393,N_14438);
and U14573 (N_14573,N_14316,N_14249);
and U14574 (N_14574,N_14443,N_14303);
nor U14575 (N_14575,N_14452,N_14003);
or U14576 (N_14576,N_14074,N_14332);
or U14577 (N_14577,N_14499,N_14435);
or U14578 (N_14578,N_14344,N_14109);
or U14579 (N_14579,N_14416,N_14264);
or U14580 (N_14580,N_14121,N_14434);
xor U14581 (N_14581,N_14133,N_14080);
and U14582 (N_14582,N_14105,N_14198);
nor U14583 (N_14583,N_14448,N_14077);
or U14584 (N_14584,N_14176,N_14446);
or U14585 (N_14585,N_14440,N_14248);
or U14586 (N_14586,N_14384,N_14395);
xnor U14587 (N_14587,N_14128,N_14373);
xnor U14588 (N_14588,N_14461,N_14190);
nand U14589 (N_14589,N_14047,N_14322);
nor U14590 (N_14590,N_14487,N_14090);
or U14591 (N_14591,N_14262,N_14182);
nand U14592 (N_14592,N_14437,N_14406);
nand U14593 (N_14593,N_14401,N_14044);
and U14594 (N_14594,N_14228,N_14049);
nor U14595 (N_14595,N_14470,N_14131);
xnor U14596 (N_14596,N_14216,N_14032);
and U14597 (N_14597,N_14429,N_14475);
nor U14598 (N_14598,N_14388,N_14329);
nor U14599 (N_14599,N_14449,N_14118);
or U14600 (N_14600,N_14076,N_14064);
or U14601 (N_14601,N_14059,N_14426);
nor U14602 (N_14602,N_14483,N_14000);
and U14603 (N_14603,N_14185,N_14242);
and U14604 (N_14604,N_14233,N_14246);
or U14605 (N_14605,N_14269,N_14022);
or U14606 (N_14606,N_14005,N_14478);
and U14607 (N_14607,N_14365,N_14278);
xor U14608 (N_14608,N_14117,N_14493);
or U14609 (N_14609,N_14403,N_14368);
and U14610 (N_14610,N_14383,N_14037);
or U14611 (N_14611,N_14051,N_14350);
or U14612 (N_14612,N_14374,N_14271);
nand U14613 (N_14613,N_14232,N_14323);
nand U14614 (N_14614,N_14157,N_14414);
nand U14615 (N_14615,N_14197,N_14144);
nor U14616 (N_14616,N_14476,N_14295);
xnor U14617 (N_14617,N_14006,N_14250);
or U14618 (N_14618,N_14071,N_14101);
or U14619 (N_14619,N_14177,N_14207);
nand U14620 (N_14620,N_14290,N_14120);
xor U14621 (N_14621,N_14147,N_14288);
and U14622 (N_14622,N_14455,N_14495);
or U14623 (N_14623,N_14137,N_14252);
xnor U14624 (N_14624,N_14444,N_14436);
or U14625 (N_14625,N_14282,N_14162);
xor U14626 (N_14626,N_14094,N_14107);
nor U14627 (N_14627,N_14172,N_14200);
or U14628 (N_14628,N_14042,N_14304);
nand U14629 (N_14629,N_14033,N_14301);
and U14630 (N_14630,N_14219,N_14013);
nand U14631 (N_14631,N_14354,N_14325);
xnor U14632 (N_14632,N_14019,N_14468);
xnor U14633 (N_14633,N_14021,N_14424);
or U14634 (N_14634,N_14419,N_14245);
and U14635 (N_14635,N_14481,N_14463);
nor U14636 (N_14636,N_14369,N_14040);
and U14637 (N_14637,N_14428,N_14199);
nor U14638 (N_14638,N_14348,N_14358);
nor U14639 (N_14639,N_14484,N_14123);
nand U14640 (N_14640,N_14072,N_14031);
nand U14641 (N_14641,N_14136,N_14066);
nor U14642 (N_14642,N_14056,N_14266);
and U14643 (N_14643,N_14442,N_14036);
or U14644 (N_14644,N_14462,N_14372);
or U14645 (N_14645,N_14194,N_14291);
nor U14646 (N_14646,N_14405,N_14106);
xnor U14647 (N_14647,N_14412,N_14108);
nand U14648 (N_14648,N_14333,N_14231);
and U14649 (N_14649,N_14404,N_14320);
xnor U14650 (N_14650,N_14104,N_14211);
nand U14651 (N_14651,N_14055,N_14163);
and U14652 (N_14652,N_14183,N_14399);
or U14653 (N_14653,N_14098,N_14453);
nand U14654 (N_14654,N_14302,N_14058);
nand U14655 (N_14655,N_14155,N_14127);
nor U14656 (N_14656,N_14299,N_14425);
xnor U14657 (N_14657,N_14087,N_14046);
and U14658 (N_14658,N_14268,N_14001);
and U14659 (N_14659,N_14456,N_14439);
or U14660 (N_14660,N_14161,N_14116);
nand U14661 (N_14661,N_14244,N_14318);
nor U14662 (N_14662,N_14361,N_14339);
or U14663 (N_14663,N_14280,N_14141);
and U14664 (N_14664,N_14160,N_14279);
nor U14665 (N_14665,N_14265,N_14494);
nor U14666 (N_14666,N_14097,N_14212);
xor U14667 (N_14667,N_14173,N_14454);
and U14668 (N_14668,N_14229,N_14335);
and U14669 (N_14669,N_14113,N_14039);
or U14670 (N_14670,N_14214,N_14025);
nor U14671 (N_14671,N_14011,N_14390);
or U14672 (N_14672,N_14272,N_14030);
nor U14673 (N_14673,N_14466,N_14402);
nor U14674 (N_14674,N_14306,N_14347);
nand U14675 (N_14675,N_14349,N_14256);
or U14676 (N_14676,N_14038,N_14054);
xor U14677 (N_14677,N_14257,N_14243);
nand U14678 (N_14678,N_14386,N_14260);
nand U14679 (N_14679,N_14297,N_14068);
or U14680 (N_14680,N_14337,N_14287);
and U14681 (N_14681,N_14159,N_14367);
nand U14682 (N_14682,N_14175,N_14189);
xnor U14683 (N_14683,N_14417,N_14050);
or U14684 (N_14684,N_14009,N_14235);
xnor U14685 (N_14685,N_14286,N_14328);
nand U14686 (N_14686,N_14292,N_14086);
xnor U14687 (N_14687,N_14153,N_14004);
nand U14688 (N_14688,N_14313,N_14099);
nor U14689 (N_14689,N_14450,N_14413);
nand U14690 (N_14690,N_14273,N_14092);
nand U14691 (N_14691,N_14289,N_14007);
nand U14692 (N_14692,N_14070,N_14103);
nand U14693 (N_14693,N_14188,N_14065);
xnor U14694 (N_14694,N_14340,N_14352);
and U14695 (N_14695,N_14294,N_14430);
and U14696 (N_14696,N_14181,N_14095);
or U14697 (N_14697,N_14081,N_14061);
or U14698 (N_14698,N_14467,N_14457);
nor U14699 (N_14699,N_14091,N_14382);
nand U14700 (N_14700,N_14150,N_14084);
nand U14701 (N_14701,N_14237,N_14180);
xnor U14702 (N_14702,N_14026,N_14205);
nand U14703 (N_14703,N_14310,N_14431);
xnor U14704 (N_14704,N_14132,N_14285);
nor U14705 (N_14705,N_14284,N_14179);
nor U14706 (N_14706,N_14154,N_14151);
or U14707 (N_14707,N_14241,N_14396);
and U14708 (N_14708,N_14421,N_14469);
or U14709 (N_14709,N_14023,N_14002);
and U14710 (N_14710,N_14126,N_14209);
nor U14711 (N_14711,N_14008,N_14027);
nand U14712 (N_14712,N_14308,N_14378);
nand U14713 (N_14713,N_14195,N_14191);
or U14714 (N_14714,N_14075,N_14300);
xor U14715 (N_14715,N_14433,N_14408);
nor U14716 (N_14716,N_14311,N_14166);
nand U14717 (N_14717,N_14078,N_14258);
nor U14718 (N_14718,N_14226,N_14236);
nand U14719 (N_14719,N_14385,N_14028);
and U14720 (N_14720,N_14496,N_14389);
nor U14721 (N_14721,N_14422,N_14486);
and U14722 (N_14722,N_14110,N_14192);
nor U14723 (N_14723,N_14202,N_14330);
nand U14724 (N_14724,N_14263,N_14380);
xor U14725 (N_14725,N_14082,N_14485);
or U14726 (N_14726,N_14124,N_14208);
nand U14727 (N_14727,N_14307,N_14115);
nor U14728 (N_14728,N_14043,N_14255);
or U14729 (N_14729,N_14186,N_14331);
xnor U14730 (N_14730,N_14480,N_14053);
xnor U14731 (N_14731,N_14206,N_14240);
or U14732 (N_14732,N_14324,N_14062);
or U14733 (N_14733,N_14387,N_14149);
or U14734 (N_14734,N_14360,N_14267);
xor U14735 (N_14735,N_14451,N_14305);
xor U14736 (N_14736,N_14224,N_14407);
nor U14737 (N_14737,N_14057,N_14423);
and U14738 (N_14738,N_14073,N_14052);
nand U14739 (N_14739,N_14364,N_14346);
or U14740 (N_14740,N_14336,N_14079);
nand U14741 (N_14741,N_14035,N_14184);
nor U14742 (N_14742,N_14251,N_14140);
xnor U14743 (N_14743,N_14471,N_14012);
or U14744 (N_14744,N_14165,N_14482);
or U14745 (N_14745,N_14024,N_14247);
nor U14746 (N_14746,N_14355,N_14238);
nor U14747 (N_14747,N_14498,N_14321);
and U14748 (N_14748,N_14152,N_14490);
nand U14749 (N_14749,N_14164,N_14460);
xor U14750 (N_14750,N_14277,N_14138);
xor U14751 (N_14751,N_14087,N_14442);
nor U14752 (N_14752,N_14416,N_14497);
or U14753 (N_14753,N_14051,N_14055);
or U14754 (N_14754,N_14477,N_14075);
nand U14755 (N_14755,N_14385,N_14414);
nor U14756 (N_14756,N_14043,N_14019);
xnor U14757 (N_14757,N_14255,N_14346);
nor U14758 (N_14758,N_14066,N_14043);
or U14759 (N_14759,N_14373,N_14484);
and U14760 (N_14760,N_14071,N_14051);
xnor U14761 (N_14761,N_14178,N_14495);
nor U14762 (N_14762,N_14226,N_14204);
nand U14763 (N_14763,N_14071,N_14383);
and U14764 (N_14764,N_14205,N_14100);
or U14765 (N_14765,N_14093,N_14035);
nor U14766 (N_14766,N_14094,N_14401);
nand U14767 (N_14767,N_14437,N_14313);
nor U14768 (N_14768,N_14184,N_14199);
xor U14769 (N_14769,N_14475,N_14196);
xnor U14770 (N_14770,N_14172,N_14001);
or U14771 (N_14771,N_14097,N_14373);
nand U14772 (N_14772,N_14269,N_14029);
xnor U14773 (N_14773,N_14170,N_14270);
nand U14774 (N_14774,N_14057,N_14283);
nand U14775 (N_14775,N_14097,N_14491);
nor U14776 (N_14776,N_14150,N_14438);
xnor U14777 (N_14777,N_14239,N_14165);
nand U14778 (N_14778,N_14457,N_14292);
or U14779 (N_14779,N_14107,N_14423);
nor U14780 (N_14780,N_14475,N_14293);
nand U14781 (N_14781,N_14184,N_14168);
nor U14782 (N_14782,N_14056,N_14379);
or U14783 (N_14783,N_14152,N_14050);
xnor U14784 (N_14784,N_14162,N_14472);
or U14785 (N_14785,N_14346,N_14206);
or U14786 (N_14786,N_14305,N_14362);
nor U14787 (N_14787,N_14482,N_14048);
and U14788 (N_14788,N_14491,N_14079);
xnor U14789 (N_14789,N_14460,N_14044);
or U14790 (N_14790,N_14328,N_14154);
nand U14791 (N_14791,N_14455,N_14072);
and U14792 (N_14792,N_14240,N_14480);
xnor U14793 (N_14793,N_14076,N_14444);
nor U14794 (N_14794,N_14413,N_14182);
nor U14795 (N_14795,N_14054,N_14032);
nand U14796 (N_14796,N_14431,N_14102);
or U14797 (N_14797,N_14484,N_14375);
or U14798 (N_14798,N_14269,N_14162);
nand U14799 (N_14799,N_14047,N_14117);
nor U14800 (N_14800,N_14148,N_14158);
and U14801 (N_14801,N_14145,N_14469);
or U14802 (N_14802,N_14205,N_14101);
or U14803 (N_14803,N_14094,N_14351);
and U14804 (N_14804,N_14252,N_14209);
nor U14805 (N_14805,N_14445,N_14286);
xor U14806 (N_14806,N_14391,N_14285);
nand U14807 (N_14807,N_14354,N_14038);
or U14808 (N_14808,N_14287,N_14435);
xor U14809 (N_14809,N_14083,N_14247);
xor U14810 (N_14810,N_14485,N_14270);
or U14811 (N_14811,N_14487,N_14484);
nor U14812 (N_14812,N_14107,N_14170);
and U14813 (N_14813,N_14256,N_14039);
and U14814 (N_14814,N_14463,N_14008);
and U14815 (N_14815,N_14187,N_14340);
nor U14816 (N_14816,N_14373,N_14461);
nor U14817 (N_14817,N_14393,N_14379);
nand U14818 (N_14818,N_14176,N_14217);
nand U14819 (N_14819,N_14393,N_14459);
nand U14820 (N_14820,N_14471,N_14050);
nand U14821 (N_14821,N_14075,N_14116);
or U14822 (N_14822,N_14377,N_14345);
nand U14823 (N_14823,N_14209,N_14384);
nor U14824 (N_14824,N_14473,N_14231);
or U14825 (N_14825,N_14066,N_14378);
xor U14826 (N_14826,N_14456,N_14336);
or U14827 (N_14827,N_14465,N_14472);
or U14828 (N_14828,N_14240,N_14211);
nor U14829 (N_14829,N_14029,N_14263);
and U14830 (N_14830,N_14394,N_14485);
or U14831 (N_14831,N_14029,N_14461);
and U14832 (N_14832,N_14115,N_14499);
xnor U14833 (N_14833,N_14408,N_14338);
and U14834 (N_14834,N_14122,N_14497);
and U14835 (N_14835,N_14407,N_14246);
xor U14836 (N_14836,N_14220,N_14055);
nand U14837 (N_14837,N_14420,N_14434);
and U14838 (N_14838,N_14197,N_14055);
nor U14839 (N_14839,N_14445,N_14335);
xnor U14840 (N_14840,N_14153,N_14281);
nor U14841 (N_14841,N_14300,N_14474);
xnor U14842 (N_14842,N_14482,N_14064);
and U14843 (N_14843,N_14384,N_14170);
or U14844 (N_14844,N_14486,N_14445);
nor U14845 (N_14845,N_14498,N_14105);
or U14846 (N_14846,N_14430,N_14104);
xor U14847 (N_14847,N_14450,N_14354);
or U14848 (N_14848,N_14060,N_14237);
or U14849 (N_14849,N_14175,N_14156);
xor U14850 (N_14850,N_14301,N_14339);
xnor U14851 (N_14851,N_14062,N_14305);
and U14852 (N_14852,N_14440,N_14339);
and U14853 (N_14853,N_14145,N_14085);
xnor U14854 (N_14854,N_14071,N_14343);
nand U14855 (N_14855,N_14160,N_14267);
nand U14856 (N_14856,N_14107,N_14012);
nand U14857 (N_14857,N_14132,N_14326);
and U14858 (N_14858,N_14410,N_14151);
nand U14859 (N_14859,N_14283,N_14444);
and U14860 (N_14860,N_14185,N_14223);
or U14861 (N_14861,N_14252,N_14315);
xnor U14862 (N_14862,N_14278,N_14109);
nand U14863 (N_14863,N_14048,N_14403);
nand U14864 (N_14864,N_14081,N_14220);
xnor U14865 (N_14865,N_14161,N_14108);
nor U14866 (N_14866,N_14224,N_14400);
xnor U14867 (N_14867,N_14214,N_14322);
and U14868 (N_14868,N_14126,N_14022);
nor U14869 (N_14869,N_14002,N_14057);
and U14870 (N_14870,N_14201,N_14017);
nand U14871 (N_14871,N_14232,N_14415);
and U14872 (N_14872,N_14215,N_14165);
nand U14873 (N_14873,N_14239,N_14244);
nor U14874 (N_14874,N_14464,N_14440);
or U14875 (N_14875,N_14445,N_14127);
and U14876 (N_14876,N_14264,N_14484);
xor U14877 (N_14877,N_14305,N_14225);
or U14878 (N_14878,N_14221,N_14072);
nand U14879 (N_14879,N_14397,N_14089);
and U14880 (N_14880,N_14468,N_14460);
xor U14881 (N_14881,N_14384,N_14084);
nand U14882 (N_14882,N_14008,N_14195);
and U14883 (N_14883,N_14379,N_14358);
and U14884 (N_14884,N_14427,N_14034);
xnor U14885 (N_14885,N_14241,N_14110);
nand U14886 (N_14886,N_14291,N_14238);
nor U14887 (N_14887,N_14005,N_14443);
and U14888 (N_14888,N_14409,N_14492);
or U14889 (N_14889,N_14124,N_14082);
xor U14890 (N_14890,N_14310,N_14197);
xor U14891 (N_14891,N_14298,N_14177);
or U14892 (N_14892,N_14066,N_14141);
and U14893 (N_14893,N_14324,N_14455);
xnor U14894 (N_14894,N_14408,N_14222);
nand U14895 (N_14895,N_14220,N_14322);
xor U14896 (N_14896,N_14454,N_14377);
xnor U14897 (N_14897,N_14413,N_14277);
xnor U14898 (N_14898,N_14097,N_14485);
xnor U14899 (N_14899,N_14154,N_14211);
xor U14900 (N_14900,N_14463,N_14070);
nor U14901 (N_14901,N_14268,N_14423);
nor U14902 (N_14902,N_14160,N_14312);
nand U14903 (N_14903,N_14469,N_14407);
nor U14904 (N_14904,N_14138,N_14226);
nor U14905 (N_14905,N_14306,N_14152);
xor U14906 (N_14906,N_14407,N_14133);
nand U14907 (N_14907,N_14229,N_14057);
or U14908 (N_14908,N_14068,N_14138);
and U14909 (N_14909,N_14435,N_14152);
xor U14910 (N_14910,N_14266,N_14310);
or U14911 (N_14911,N_14399,N_14490);
and U14912 (N_14912,N_14304,N_14439);
or U14913 (N_14913,N_14389,N_14163);
xnor U14914 (N_14914,N_14359,N_14313);
nor U14915 (N_14915,N_14289,N_14108);
xnor U14916 (N_14916,N_14311,N_14221);
xnor U14917 (N_14917,N_14378,N_14032);
and U14918 (N_14918,N_14300,N_14141);
xor U14919 (N_14919,N_14443,N_14111);
xnor U14920 (N_14920,N_14350,N_14354);
and U14921 (N_14921,N_14010,N_14475);
nor U14922 (N_14922,N_14350,N_14061);
or U14923 (N_14923,N_14268,N_14313);
xor U14924 (N_14924,N_14375,N_14176);
and U14925 (N_14925,N_14496,N_14275);
or U14926 (N_14926,N_14000,N_14468);
or U14927 (N_14927,N_14112,N_14189);
and U14928 (N_14928,N_14093,N_14398);
xnor U14929 (N_14929,N_14151,N_14156);
nor U14930 (N_14930,N_14375,N_14161);
nand U14931 (N_14931,N_14372,N_14188);
xnor U14932 (N_14932,N_14250,N_14370);
xor U14933 (N_14933,N_14413,N_14228);
xor U14934 (N_14934,N_14302,N_14405);
xor U14935 (N_14935,N_14452,N_14048);
nand U14936 (N_14936,N_14220,N_14194);
or U14937 (N_14937,N_14345,N_14340);
and U14938 (N_14938,N_14421,N_14007);
and U14939 (N_14939,N_14177,N_14335);
nor U14940 (N_14940,N_14107,N_14124);
nand U14941 (N_14941,N_14095,N_14069);
nand U14942 (N_14942,N_14459,N_14065);
or U14943 (N_14943,N_14113,N_14104);
nor U14944 (N_14944,N_14341,N_14293);
xnor U14945 (N_14945,N_14448,N_14177);
nand U14946 (N_14946,N_14344,N_14420);
nor U14947 (N_14947,N_14175,N_14262);
xnor U14948 (N_14948,N_14297,N_14304);
and U14949 (N_14949,N_14220,N_14047);
and U14950 (N_14950,N_14417,N_14084);
xor U14951 (N_14951,N_14268,N_14372);
nor U14952 (N_14952,N_14156,N_14399);
nor U14953 (N_14953,N_14355,N_14391);
and U14954 (N_14954,N_14387,N_14050);
xor U14955 (N_14955,N_14316,N_14119);
or U14956 (N_14956,N_14466,N_14418);
xnor U14957 (N_14957,N_14026,N_14214);
and U14958 (N_14958,N_14429,N_14493);
xnor U14959 (N_14959,N_14358,N_14461);
and U14960 (N_14960,N_14221,N_14434);
nor U14961 (N_14961,N_14326,N_14379);
or U14962 (N_14962,N_14388,N_14484);
nor U14963 (N_14963,N_14099,N_14154);
xnor U14964 (N_14964,N_14439,N_14360);
and U14965 (N_14965,N_14453,N_14251);
xnor U14966 (N_14966,N_14134,N_14426);
nand U14967 (N_14967,N_14447,N_14274);
xor U14968 (N_14968,N_14101,N_14146);
nor U14969 (N_14969,N_14233,N_14188);
nand U14970 (N_14970,N_14112,N_14471);
and U14971 (N_14971,N_14303,N_14055);
nand U14972 (N_14972,N_14311,N_14051);
or U14973 (N_14973,N_14220,N_14392);
or U14974 (N_14974,N_14033,N_14223);
and U14975 (N_14975,N_14476,N_14084);
nand U14976 (N_14976,N_14278,N_14057);
or U14977 (N_14977,N_14126,N_14441);
nand U14978 (N_14978,N_14472,N_14445);
nor U14979 (N_14979,N_14005,N_14102);
and U14980 (N_14980,N_14269,N_14274);
nor U14981 (N_14981,N_14297,N_14110);
or U14982 (N_14982,N_14396,N_14065);
xnor U14983 (N_14983,N_14336,N_14407);
or U14984 (N_14984,N_14464,N_14406);
and U14985 (N_14985,N_14038,N_14059);
xnor U14986 (N_14986,N_14277,N_14318);
and U14987 (N_14987,N_14027,N_14044);
xor U14988 (N_14988,N_14323,N_14337);
nand U14989 (N_14989,N_14186,N_14442);
nor U14990 (N_14990,N_14063,N_14086);
xnor U14991 (N_14991,N_14374,N_14130);
or U14992 (N_14992,N_14427,N_14059);
or U14993 (N_14993,N_14432,N_14144);
xnor U14994 (N_14994,N_14186,N_14360);
nor U14995 (N_14995,N_14417,N_14433);
and U14996 (N_14996,N_14231,N_14424);
xnor U14997 (N_14997,N_14187,N_14175);
xor U14998 (N_14998,N_14375,N_14081);
and U14999 (N_14999,N_14038,N_14499);
or U15000 (N_15000,N_14613,N_14650);
nand U15001 (N_15001,N_14892,N_14719);
nor U15002 (N_15002,N_14758,N_14837);
or U15003 (N_15003,N_14874,N_14673);
nor U15004 (N_15004,N_14510,N_14718);
and U15005 (N_15005,N_14964,N_14503);
and U15006 (N_15006,N_14654,N_14971);
and U15007 (N_15007,N_14596,N_14771);
nor U15008 (N_15008,N_14560,N_14949);
nor U15009 (N_15009,N_14842,N_14559);
nand U15010 (N_15010,N_14626,N_14521);
and U15011 (N_15011,N_14506,N_14936);
or U15012 (N_15012,N_14751,N_14672);
nor U15013 (N_15013,N_14772,N_14921);
and U15014 (N_15014,N_14708,N_14863);
or U15015 (N_15015,N_14856,N_14818);
or U15016 (N_15016,N_14900,N_14760);
xor U15017 (N_15017,N_14757,N_14594);
xor U15018 (N_15018,N_14514,N_14529);
or U15019 (N_15019,N_14530,N_14883);
or U15020 (N_15020,N_14759,N_14545);
xnor U15021 (N_15021,N_14828,N_14937);
and U15022 (N_15022,N_14962,N_14695);
and U15023 (N_15023,N_14819,N_14601);
and U15024 (N_15024,N_14666,N_14821);
or U15025 (N_15025,N_14925,N_14676);
xor U15026 (N_15026,N_14661,N_14720);
xor U15027 (N_15027,N_14912,N_14508);
or U15028 (N_15028,N_14558,N_14552);
or U15029 (N_15029,N_14574,N_14788);
xnor U15030 (N_15030,N_14903,N_14645);
nand U15031 (N_15031,N_14777,N_14569);
nand U15032 (N_15032,N_14512,N_14527);
nor U15033 (N_15033,N_14966,N_14638);
xnor U15034 (N_15034,N_14605,N_14977);
xor U15035 (N_15035,N_14968,N_14565);
nor U15036 (N_15036,N_14524,N_14523);
xor U15037 (N_15037,N_14905,N_14740);
xnor U15038 (N_15038,N_14860,N_14704);
nand U15039 (N_15039,N_14745,N_14683);
nand U15040 (N_15040,N_14911,N_14698);
and U15041 (N_15041,N_14792,N_14754);
xnor U15042 (N_15042,N_14826,N_14781);
or U15043 (N_15043,N_14778,N_14848);
nor U15044 (N_15044,N_14855,N_14554);
and U15045 (N_15045,N_14710,N_14840);
and U15046 (N_15046,N_14736,N_14542);
xor U15047 (N_15047,N_14696,N_14768);
nor U15048 (N_15048,N_14501,N_14763);
xnor U15049 (N_15049,N_14904,N_14595);
nand U15050 (N_15050,N_14733,N_14582);
or U15051 (N_15051,N_14711,N_14959);
and U15052 (N_15052,N_14616,N_14847);
or U15053 (N_15053,N_14592,N_14767);
or U15054 (N_15054,N_14651,N_14539);
and U15055 (N_15055,N_14697,N_14952);
and U15056 (N_15056,N_14998,N_14954);
or U15057 (N_15057,N_14603,N_14598);
or U15058 (N_15058,N_14774,N_14556);
and U15059 (N_15059,N_14928,N_14924);
nor U15060 (N_15060,N_14681,N_14532);
nand U15061 (N_15061,N_14862,N_14817);
nand U15062 (N_15062,N_14707,N_14914);
and U15063 (N_15063,N_14541,N_14806);
or U15064 (N_15064,N_14983,N_14907);
and U15065 (N_15065,N_14607,N_14726);
xnor U15066 (N_15066,N_14667,N_14656);
xor U15067 (N_15067,N_14816,N_14713);
nand U15068 (N_15068,N_14967,N_14563);
nand U15069 (N_15069,N_14742,N_14618);
nand U15070 (N_15070,N_14665,N_14899);
xnor U15071 (N_15071,N_14987,N_14868);
or U15072 (N_15072,N_14734,N_14980);
and U15073 (N_15073,N_14858,N_14991);
and U15074 (N_15074,N_14876,N_14864);
xor U15075 (N_15075,N_14787,N_14910);
nor U15076 (N_15076,N_14625,N_14573);
xnor U15077 (N_15077,N_14641,N_14835);
nand U15078 (N_15078,N_14504,N_14852);
or U15079 (N_15079,N_14802,N_14875);
nand U15080 (N_15080,N_14690,N_14873);
and U15081 (N_15081,N_14931,N_14688);
nor U15082 (N_15082,N_14827,N_14941);
nor U15083 (N_15083,N_14775,N_14623);
nor U15084 (N_15084,N_14606,N_14640);
or U15085 (N_15085,N_14632,N_14615);
or U15086 (N_15086,N_14660,N_14857);
and U15087 (N_15087,N_14536,N_14674);
and U15088 (N_15088,N_14744,N_14790);
xnor U15089 (N_15089,N_14584,N_14943);
and U15090 (N_15090,N_14890,N_14786);
nor U15091 (N_15091,N_14551,N_14649);
and U15092 (N_15092,N_14628,N_14516);
and U15093 (N_15093,N_14624,N_14915);
or U15094 (N_15094,N_14940,N_14561);
xor U15095 (N_15095,N_14534,N_14990);
nor U15096 (N_15096,N_14716,N_14981);
or U15097 (N_15097,N_14648,N_14526);
xnor U15098 (N_15098,N_14955,N_14549);
or U15099 (N_15099,N_14870,N_14557);
and U15100 (N_15100,N_14811,N_14965);
and U15101 (N_15101,N_14597,N_14702);
nor U15102 (N_15102,N_14942,N_14723);
nor U15103 (N_15103,N_14764,N_14583);
xor U15104 (N_15104,N_14762,N_14995);
nand U15105 (N_15105,N_14933,N_14620);
nand U15106 (N_15106,N_14974,N_14520);
and U15107 (N_15107,N_14916,N_14579);
nand U15108 (N_15108,N_14999,N_14570);
xnor U15109 (N_15109,N_14838,N_14895);
xnor U15110 (N_15110,N_14783,N_14963);
nand U15111 (N_15111,N_14580,N_14988);
xnor U15112 (N_15112,N_14658,N_14957);
or U15113 (N_15113,N_14951,N_14646);
or U15114 (N_15114,N_14973,N_14538);
or U15115 (N_15115,N_14678,N_14630);
nand U15116 (N_15116,N_14642,N_14861);
nor U15117 (N_15117,N_14752,N_14970);
nand U15118 (N_15118,N_14800,N_14635);
or U15119 (N_15119,N_14587,N_14629);
nor U15120 (N_15120,N_14555,N_14839);
nor U15121 (N_15121,N_14923,N_14715);
nor U15122 (N_15122,N_14636,N_14770);
or U15123 (N_15123,N_14691,N_14714);
nand U15124 (N_15124,N_14884,N_14647);
nor U15125 (N_15125,N_14608,N_14515);
and U15126 (N_15126,N_14902,N_14637);
nor U15127 (N_15127,N_14631,N_14577);
nor U15128 (N_15128,N_14797,N_14805);
nor U15129 (N_15129,N_14982,N_14908);
nor U15130 (N_15130,N_14897,N_14865);
xor U15131 (N_15131,N_14706,N_14578);
and U15132 (N_15132,N_14680,N_14547);
or U15133 (N_15133,N_14929,N_14617);
nor U15134 (N_15134,N_14668,N_14544);
nor U15135 (N_15135,N_14765,N_14675);
or U15136 (N_15136,N_14815,N_14502);
nor U15137 (N_15137,N_14913,N_14602);
nand U15138 (N_15138,N_14693,N_14992);
nor U15139 (N_15139,N_14894,N_14830);
nor U15140 (N_15140,N_14801,N_14945);
nand U15141 (N_15141,N_14849,N_14750);
and U15142 (N_15142,N_14985,N_14591);
and U15143 (N_15143,N_14731,N_14960);
nor U15144 (N_15144,N_14956,N_14834);
nor U15145 (N_15145,N_14938,N_14677);
or U15146 (N_15146,N_14585,N_14548);
xnor U15147 (N_15147,N_14671,N_14776);
xnor U15148 (N_15148,N_14589,N_14738);
and U15149 (N_15149,N_14853,N_14896);
and U15150 (N_15150,N_14824,N_14746);
nand U15151 (N_15151,N_14798,N_14562);
and U15152 (N_15152,N_14619,N_14872);
nand U15153 (N_15153,N_14918,N_14748);
and U15154 (N_15154,N_14947,N_14909);
nor U15155 (N_15155,N_14513,N_14946);
xnor U15156 (N_15156,N_14851,N_14845);
nand U15157 (N_15157,N_14784,N_14749);
nor U15158 (N_15158,N_14934,N_14730);
nand U15159 (N_15159,N_14511,N_14922);
or U15160 (N_15160,N_14993,N_14887);
xor U15161 (N_15161,N_14808,N_14567);
xor U15162 (N_15162,N_14935,N_14659);
nor U15163 (N_15163,N_14846,N_14901);
nor U15164 (N_15164,N_14878,N_14886);
nor U15165 (N_15165,N_14810,N_14881);
xor U15166 (N_15166,N_14871,N_14709);
and U15167 (N_15167,N_14793,N_14885);
nor U15168 (N_15168,N_14682,N_14739);
or U15169 (N_15169,N_14888,N_14796);
xnor U15170 (N_15170,N_14729,N_14590);
nand U15171 (N_15171,N_14564,N_14753);
nand U15172 (N_15172,N_14893,N_14535);
and U15173 (N_15173,N_14930,N_14932);
nor U15174 (N_15174,N_14586,N_14572);
nor U15175 (N_15175,N_14531,N_14571);
or U15176 (N_15176,N_14721,N_14780);
nor U15177 (N_15177,N_14722,N_14737);
nor U15178 (N_15178,N_14814,N_14822);
nand U15179 (N_15179,N_14939,N_14841);
or U15180 (N_15180,N_14779,N_14703);
nor U15181 (N_15181,N_14794,N_14755);
xnor U15182 (N_15182,N_14517,N_14553);
xnor U15183 (N_15183,N_14525,N_14880);
xor U15184 (N_15184,N_14699,N_14537);
xnor U15185 (N_15185,N_14773,N_14568);
xnor U15186 (N_15186,N_14576,N_14741);
and U15187 (N_15187,N_14543,N_14614);
and U15188 (N_15188,N_14882,N_14877);
or U15189 (N_15189,N_14728,N_14789);
xnor U15190 (N_15190,N_14593,N_14621);
and U15191 (N_15191,N_14969,N_14989);
xnor U15192 (N_15192,N_14700,N_14509);
and U15193 (N_15193,N_14727,N_14664);
xnor U15194 (N_15194,N_14831,N_14743);
and U15195 (N_15195,N_14994,N_14604);
xor U15196 (N_15196,N_14979,N_14581);
nor U15197 (N_15197,N_14953,N_14799);
nor U15198 (N_15198,N_14919,N_14528);
nand U15199 (N_15199,N_14725,N_14735);
nor U15200 (N_15200,N_14825,N_14519);
xnor U15201 (N_15201,N_14747,N_14609);
and U15202 (N_15202,N_14782,N_14701);
or U15203 (N_15203,N_14518,N_14652);
nor U15204 (N_15204,N_14976,N_14687);
or U15205 (N_15205,N_14889,N_14972);
xor U15206 (N_15206,N_14948,N_14705);
nor U15207 (N_15207,N_14823,N_14653);
or U15208 (N_15208,N_14769,N_14975);
and U15209 (N_15209,N_14766,N_14958);
xnor U15210 (N_15210,N_14599,N_14869);
and U15211 (N_15211,N_14575,N_14996);
and U15212 (N_15212,N_14732,N_14906);
and U15213 (N_15213,N_14984,N_14655);
nor U15214 (N_15214,N_14926,N_14540);
or U15215 (N_15215,N_14550,N_14920);
nor U15216 (N_15216,N_14669,N_14644);
or U15217 (N_15217,N_14761,N_14600);
and U15218 (N_15218,N_14807,N_14566);
xnor U15219 (N_15219,N_14867,N_14997);
and U15220 (N_15220,N_14866,N_14643);
or U15221 (N_15221,N_14812,N_14679);
or U15222 (N_15222,N_14986,N_14507);
nor U15223 (N_15223,N_14756,N_14634);
xnor U15224 (N_15224,N_14836,N_14879);
xnor U15225 (N_15225,N_14610,N_14917);
nor U15226 (N_15226,N_14717,N_14791);
nand U15227 (N_15227,N_14692,N_14859);
or U15228 (N_15228,N_14712,N_14612);
or U15229 (N_15229,N_14533,N_14670);
nand U15230 (N_15230,N_14854,N_14663);
nor U15231 (N_15231,N_14961,N_14844);
nor U15232 (N_15232,N_14891,N_14500);
and U15233 (N_15233,N_14820,N_14622);
nand U15234 (N_15234,N_14522,N_14611);
xnor U15235 (N_15235,N_14809,N_14804);
and U15236 (N_15236,N_14694,N_14662);
nand U15237 (N_15237,N_14785,N_14944);
and U15238 (N_15238,N_14833,N_14832);
nor U15239 (N_15239,N_14689,N_14546);
and U15240 (N_15240,N_14657,N_14813);
and U15241 (N_15241,N_14803,N_14627);
or U15242 (N_15242,N_14850,N_14505);
nor U15243 (N_15243,N_14843,N_14795);
and U15244 (N_15244,N_14950,N_14978);
nor U15245 (N_15245,N_14927,N_14686);
and U15246 (N_15246,N_14639,N_14685);
xor U15247 (N_15247,N_14633,N_14684);
xnor U15248 (N_15248,N_14724,N_14898);
or U15249 (N_15249,N_14829,N_14588);
nor U15250 (N_15250,N_14638,N_14574);
or U15251 (N_15251,N_14614,N_14584);
nand U15252 (N_15252,N_14928,N_14817);
nor U15253 (N_15253,N_14687,N_14832);
and U15254 (N_15254,N_14830,N_14720);
nand U15255 (N_15255,N_14978,N_14636);
nor U15256 (N_15256,N_14908,N_14886);
nand U15257 (N_15257,N_14533,N_14858);
nand U15258 (N_15258,N_14706,N_14549);
nand U15259 (N_15259,N_14895,N_14606);
nor U15260 (N_15260,N_14674,N_14621);
nor U15261 (N_15261,N_14939,N_14829);
xnor U15262 (N_15262,N_14908,N_14545);
xor U15263 (N_15263,N_14619,N_14625);
nor U15264 (N_15264,N_14556,N_14997);
xor U15265 (N_15265,N_14852,N_14830);
xor U15266 (N_15266,N_14815,N_14957);
and U15267 (N_15267,N_14724,N_14587);
or U15268 (N_15268,N_14547,N_14770);
nand U15269 (N_15269,N_14587,N_14881);
xor U15270 (N_15270,N_14761,N_14655);
nor U15271 (N_15271,N_14772,N_14848);
xnor U15272 (N_15272,N_14757,N_14667);
xnor U15273 (N_15273,N_14805,N_14729);
or U15274 (N_15274,N_14999,N_14871);
nor U15275 (N_15275,N_14548,N_14671);
and U15276 (N_15276,N_14874,N_14902);
or U15277 (N_15277,N_14910,N_14686);
or U15278 (N_15278,N_14587,N_14607);
nand U15279 (N_15279,N_14917,N_14861);
and U15280 (N_15280,N_14815,N_14735);
or U15281 (N_15281,N_14750,N_14810);
xnor U15282 (N_15282,N_14865,N_14804);
nand U15283 (N_15283,N_14633,N_14950);
xor U15284 (N_15284,N_14865,N_14666);
or U15285 (N_15285,N_14749,N_14585);
nand U15286 (N_15286,N_14656,N_14594);
nor U15287 (N_15287,N_14848,N_14931);
and U15288 (N_15288,N_14638,N_14668);
and U15289 (N_15289,N_14659,N_14761);
xor U15290 (N_15290,N_14749,N_14702);
nand U15291 (N_15291,N_14783,N_14980);
nor U15292 (N_15292,N_14869,N_14950);
or U15293 (N_15293,N_14806,N_14610);
and U15294 (N_15294,N_14910,N_14656);
and U15295 (N_15295,N_14653,N_14538);
nand U15296 (N_15296,N_14730,N_14541);
and U15297 (N_15297,N_14744,N_14522);
xnor U15298 (N_15298,N_14638,N_14940);
nand U15299 (N_15299,N_14948,N_14505);
or U15300 (N_15300,N_14735,N_14945);
nand U15301 (N_15301,N_14657,N_14903);
and U15302 (N_15302,N_14802,N_14955);
nor U15303 (N_15303,N_14883,N_14999);
or U15304 (N_15304,N_14545,N_14838);
xor U15305 (N_15305,N_14987,N_14846);
nand U15306 (N_15306,N_14674,N_14743);
xor U15307 (N_15307,N_14556,N_14715);
xnor U15308 (N_15308,N_14636,N_14621);
nand U15309 (N_15309,N_14789,N_14602);
nor U15310 (N_15310,N_14704,N_14564);
xor U15311 (N_15311,N_14702,N_14846);
nand U15312 (N_15312,N_14824,N_14626);
nand U15313 (N_15313,N_14664,N_14740);
and U15314 (N_15314,N_14972,N_14755);
xor U15315 (N_15315,N_14889,N_14586);
nand U15316 (N_15316,N_14660,N_14978);
nor U15317 (N_15317,N_14957,N_14530);
xor U15318 (N_15318,N_14900,N_14810);
nor U15319 (N_15319,N_14522,N_14577);
nor U15320 (N_15320,N_14871,N_14879);
and U15321 (N_15321,N_14880,N_14867);
nand U15322 (N_15322,N_14528,N_14987);
xor U15323 (N_15323,N_14790,N_14520);
and U15324 (N_15324,N_14933,N_14926);
or U15325 (N_15325,N_14735,N_14642);
nand U15326 (N_15326,N_14742,N_14654);
nand U15327 (N_15327,N_14566,N_14652);
and U15328 (N_15328,N_14875,N_14877);
nand U15329 (N_15329,N_14833,N_14743);
nor U15330 (N_15330,N_14746,N_14993);
nor U15331 (N_15331,N_14892,N_14740);
xor U15332 (N_15332,N_14649,N_14865);
nand U15333 (N_15333,N_14813,N_14951);
or U15334 (N_15334,N_14891,N_14588);
xnor U15335 (N_15335,N_14854,N_14665);
nand U15336 (N_15336,N_14854,N_14548);
nand U15337 (N_15337,N_14692,N_14966);
or U15338 (N_15338,N_14855,N_14887);
nand U15339 (N_15339,N_14834,N_14844);
xor U15340 (N_15340,N_14660,N_14900);
xnor U15341 (N_15341,N_14532,N_14791);
nor U15342 (N_15342,N_14553,N_14877);
and U15343 (N_15343,N_14624,N_14747);
nand U15344 (N_15344,N_14744,N_14800);
nor U15345 (N_15345,N_14882,N_14615);
and U15346 (N_15346,N_14732,N_14887);
or U15347 (N_15347,N_14916,N_14927);
nand U15348 (N_15348,N_14542,N_14742);
and U15349 (N_15349,N_14824,N_14879);
or U15350 (N_15350,N_14818,N_14787);
or U15351 (N_15351,N_14629,N_14532);
xor U15352 (N_15352,N_14647,N_14772);
or U15353 (N_15353,N_14612,N_14633);
or U15354 (N_15354,N_14923,N_14725);
and U15355 (N_15355,N_14938,N_14547);
nand U15356 (N_15356,N_14512,N_14785);
nor U15357 (N_15357,N_14923,N_14781);
and U15358 (N_15358,N_14685,N_14801);
and U15359 (N_15359,N_14648,N_14540);
xnor U15360 (N_15360,N_14745,N_14542);
nor U15361 (N_15361,N_14898,N_14742);
nand U15362 (N_15362,N_14954,N_14597);
or U15363 (N_15363,N_14961,N_14779);
nand U15364 (N_15364,N_14768,N_14618);
or U15365 (N_15365,N_14819,N_14816);
xnor U15366 (N_15366,N_14619,N_14760);
or U15367 (N_15367,N_14726,N_14679);
nand U15368 (N_15368,N_14897,N_14601);
nor U15369 (N_15369,N_14569,N_14507);
nand U15370 (N_15370,N_14618,N_14898);
xor U15371 (N_15371,N_14706,N_14762);
nor U15372 (N_15372,N_14883,N_14507);
nor U15373 (N_15373,N_14728,N_14605);
xor U15374 (N_15374,N_14640,N_14864);
or U15375 (N_15375,N_14549,N_14598);
or U15376 (N_15376,N_14785,N_14877);
xor U15377 (N_15377,N_14949,N_14730);
xnor U15378 (N_15378,N_14921,N_14938);
or U15379 (N_15379,N_14883,N_14633);
nor U15380 (N_15380,N_14666,N_14585);
or U15381 (N_15381,N_14971,N_14669);
xor U15382 (N_15382,N_14863,N_14755);
and U15383 (N_15383,N_14644,N_14700);
nor U15384 (N_15384,N_14695,N_14762);
nand U15385 (N_15385,N_14981,N_14938);
xor U15386 (N_15386,N_14807,N_14989);
xor U15387 (N_15387,N_14596,N_14997);
and U15388 (N_15388,N_14755,N_14884);
xnor U15389 (N_15389,N_14503,N_14581);
or U15390 (N_15390,N_14581,N_14786);
nand U15391 (N_15391,N_14891,N_14585);
nand U15392 (N_15392,N_14507,N_14845);
xnor U15393 (N_15393,N_14659,N_14720);
or U15394 (N_15394,N_14949,N_14661);
xnor U15395 (N_15395,N_14675,N_14845);
xor U15396 (N_15396,N_14865,N_14584);
xnor U15397 (N_15397,N_14594,N_14695);
nand U15398 (N_15398,N_14604,N_14530);
or U15399 (N_15399,N_14596,N_14793);
and U15400 (N_15400,N_14983,N_14531);
xor U15401 (N_15401,N_14722,N_14983);
nand U15402 (N_15402,N_14802,N_14998);
and U15403 (N_15403,N_14785,N_14515);
or U15404 (N_15404,N_14782,N_14834);
xor U15405 (N_15405,N_14828,N_14503);
and U15406 (N_15406,N_14566,N_14654);
or U15407 (N_15407,N_14631,N_14907);
nor U15408 (N_15408,N_14631,N_14534);
nand U15409 (N_15409,N_14932,N_14830);
nor U15410 (N_15410,N_14962,N_14539);
and U15411 (N_15411,N_14921,N_14869);
xnor U15412 (N_15412,N_14627,N_14886);
xnor U15413 (N_15413,N_14853,N_14568);
or U15414 (N_15414,N_14650,N_14705);
xor U15415 (N_15415,N_14669,N_14972);
nor U15416 (N_15416,N_14776,N_14697);
nand U15417 (N_15417,N_14907,N_14704);
and U15418 (N_15418,N_14876,N_14742);
or U15419 (N_15419,N_14538,N_14748);
nor U15420 (N_15420,N_14785,N_14814);
nand U15421 (N_15421,N_14713,N_14533);
nand U15422 (N_15422,N_14893,N_14792);
nand U15423 (N_15423,N_14844,N_14995);
xnor U15424 (N_15424,N_14939,N_14893);
nand U15425 (N_15425,N_14501,N_14837);
or U15426 (N_15426,N_14970,N_14961);
xor U15427 (N_15427,N_14988,N_14953);
and U15428 (N_15428,N_14701,N_14654);
nor U15429 (N_15429,N_14941,N_14636);
xor U15430 (N_15430,N_14945,N_14950);
or U15431 (N_15431,N_14879,N_14688);
nand U15432 (N_15432,N_14601,N_14675);
nand U15433 (N_15433,N_14562,N_14821);
or U15434 (N_15434,N_14937,N_14740);
and U15435 (N_15435,N_14678,N_14736);
and U15436 (N_15436,N_14886,N_14951);
nor U15437 (N_15437,N_14797,N_14648);
nand U15438 (N_15438,N_14704,N_14571);
or U15439 (N_15439,N_14606,N_14805);
and U15440 (N_15440,N_14585,N_14524);
or U15441 (N_15441,N_14740,N_14731);
or U15442 (N_15442,N_14562,N_14847);
nor U15443 (N_15443,N_14910,N_14781);
and U15444 (N_15444,N_14546,N_14657);
xor U15445 (N_15445,N_14779,N_14878);
and U15446 (N_15446,N_14830,N_14861);
and U15447 (N_15447,N_14575,N_14932);
or U15448 (N_15448,N_14634,N_14834);
nor U15449 (N_15449,N_14981,N_14564);
nor U15450 (N_15450,N_14528,N_14890);
or U15451 (N_15451,N_14697,N_14636);
nor U15452 (N_15452,N_14752,N_14544);
xnor U15453 (N_15453,N_14675,N_14534);
and U15454 (N_15454,N_14593,N_14694);
and U15455 (N_15455,N_14673,N_14781);
and U15456 (N_15456,N_14614,N_14770);
nand U15457 (N_15457,N_14637,N_14956);
xnor U15458 (N_15458,N_14533,N_14884);
nor U15459 (N_15459,N_14744,N_14922);
nor U15460 (N_15460,N_14944,N_14842);
or U15461 (N_15461,N_14572,N_14766);
nor U15462 (N_15462,N_14728,N_14633);
nor U15463 (N_15463,N_14848,N_14784);
nor U15464 (N_15464,N_14693,N_14849);
and U15465 (N_15465,N_14769,N_14945);
xnor U15466 (N_15466,N_14510,N_14869);
and U15467 (N_15467,N_14749,N_14632);
and U15468 (N_15468,N_14844,N_14781);
nand U15469 (N_15469,N_14730,N_14713);
nand U15470 (N_15470,N_14864,N_14613);
nand U15471 (N_15471,N_14651,N_14999);
or U15472 (N_15472,N_14854,N_14999);
nand U15473 (N_15473,N_14853,N_14610);
nand U15474 (N_15474,N_14604,N_14539);
and U15475 (N_15475,N_14816,N_14909);
nor U15476 (N_15476,N_14536,N_14525);
nor U15477 (N_15477,N_14751,N_14512);
xnor U15478 (N_15478,N_14969,N_14515);
nor U15479 (N_15479,N_14846,N_14924);
nand U15480 (N_15480,N_14941,N_14573);
xor U15481 (N_15481,N_14738,N_14530);
and U15482 (N_15482,N_14972,N_14931);
or U15483 (N_15483,N_14804,N_14660);
nor U15484 (N_15484,N_14647,N_14746);
or U15485 (N_15485,N_14746,N_14745);
xnor U15486 (N_15486,N_14955,N_14874);
or U15487 (N_15487,N_14559,N_14515);
xnor U15488 (N_15488,N_14576,N_14587);
nor U15489 (N_15489,N_14773,N_14882);
nand U15490 (N_15490,N_14905,N_14595);
nand U15491 (N_15491,N_14948,N_14756);
nor U15492 (N_15492,N_14850,N_14935);
nand U15493 (N_15493,N_14921,N_14870);
nand U15494 (N_15494,N_14760,N_14757);
and U15495 (N_15495,N_14763,N_14975);
and U15496 (N_15496,N_14629,N_14632);
nand U15497 (N_15497,N_14614,N_14858);
nor U15498 (N_15498,N_14834,N_14507);
nand U15499 (N_15499,N_14767,N_14797);
or U15500 (N_15500,N_15324,N_15471);
nor U15501 (N_15501,N_15013,N_15047);
xor U15502 (N_15502,N_15095,N_15210);
and U15503 (N_15503,N_15259,N_15096);
or U15504 (N_15504,N_15314,N_15078);
and U15505 (N_15505,N_15483,N_15338);
xnor U15506 (N_15506,N_15045,N_15212);
xor U15507 (N_15507,N_15003,N_15348);
nor U15508 (N_15508,N_15129,N_15151);
nand U15509 (N_15509,N_15159,N_15235);
xnor U15510 (N_15510,N_15111,N_15406);
xnor U15511 (N_15511,N_15457,N_15164);
nor U15512 (N_15512,N_15354,N_15146);
nor U15513 (N_15513,N_15200,N_15100);
nor U15514 (N_15514,N_15413,N_15296);
xor U15515 (N_15515,N_15463,N_15228);
or U15516 (N_15516,N_15071,N_15394);
or U15517 (N_15517,N_15479,N_15224);
xor U15518 (N_15518,N_15052,N_15222);
and U15519 (N_15519,N_15020,N_15009);
and U15520 (N_15520,N_15171,N_15079);
or U15521 (N_15521,N_15350,N_15410);
nor U15522 (N_15522,N_15482,N_15018);
nor U15523 (N_15523,N_15173,N_15082);
nand U15524 (N_15524,N_15172,N_15105);
or U15525 (N_15525,N_15325,N_15230);
nor U15526 (N_15526,N_15431,N_15110);
and U15527 (N_15527,N_15498,N_15250);
and U15528 (N_15528,N_15415,N_15213);
and U15529 (N_15529,N_15084,N_15391);
xor U15530 (N_15530,N_15035,N_15373);
nand U15531 (N_15531,N_15279,N_15055);
or U15532 (N_15532,N_15321,N_15201);
or U15533 (N_15533,N_15420,N_15025);
nor U15534 (N_15534,N_15118,N_15365);
nor U15535 (N_15535,N_15179,N_15496);
xor U15536 (N_15536,N_15480,N_15134);
or U15537 (N_15537,N_15476,N_15438);
nand U15538 (N_15538,N_15466,N_15097);
or U15539 (N_15539,N_15252,N_15458);
nor U15540 (N_15540,N_15298,N_15019);
nand U15541 (N_15541,N_15390,N_15232);
nor U15542 (N_15542,N_15441,N_15166);
xnor U15543 (N_15543,N_15322,N_15051);
or U15544 (N_15544,N_15137,N_15323);
nor U15545 (N_15545,N_15284,N_15157);
or U15546 (N_15546,N_15209,N_15405);
nand U15547 (N_15547,N_15380,N_15238);
xor U15548 (N_15548,N_15447,N_15233);
and U15549 (N_15549,N_15178,N_15089);
xor U15550 (N_15550,N_15419,N_15026);
or U15551 (N_15551,N_15087,N_15266);
xor U15552 (N_15552,N_15142,N_15468);
nand U15553 (N_15553,N_15368,N_15067);
xor U15554 (N_15554,N_15149,N_15421);
and U15555 (N_15555,N_15192,N_15214);
nor U15556 (N_15556,N_15370,N_15006);
nor U15557 (N_15557,N_15063,N_15371);
nand U15558 (N_15558,N_15372,N_15357);
nor U15559 (N_15559,N_15318,N_15221);
and U15560 (N_15560,N_15248,N_15046);
nand U15561 (N_15561,N_15456,N_15080);
and U15562 (N_15562,N_15285,N_15276);
or U15563 (N_15563,N_15043,N_15465);
nor U15564 (N_15564,N_15287,N_15231);
nand U15565 (N_15565,N_15351,N_15469);
nand U15566 (N_15566,N_15181,N_15029);
nor U15567 (N_15567,N_15448,N_15091);
nand U15568 (N_15568,N_15382,N_15244);
nand U15569 (N_15569,N_15211,N_15075);
xnor U15570 (N_15570,N_15311,N_15358);
nor U15571 (N_15571,N_15104,N_15384);
nand U15572 (N_15572,N_15281,N_15132);
nand U15573 (N_15573,N_15396,N_15360);
xnor U15574 (N_15574,N_15054,N_15195);
and U15575 (N_15575,N_15345,N_15467);
nand U15576 (N_15576,N_15455,N_15131);
or U15577 (N_15577,N_15460,N_15107);
xnor U15578 (N_15578,N_15305,N_15056);
nor U15579 (N_15579,N_15304,N_15088);
or U15580 (N_15580,N_15258,N_15387);
xor U15581 (N_15581,N_15416,N_15176);
nand U15582 (N_15582,N_15032,N_15265);
nor U15583 (N_15583,N_15359,N_15170);
or U15584 (N_15584,N_15484,N_15334);
or U15585 (N_15585,N_15106,N_15263);
and U15586 (N_15586,N_15388,N_15123);
or U15587 (N_15587,N_15090,N_15393);
and U15588 (N_15588,N_15422,N_15464);
or U15589 (N_15589,N_15016,N_15128);
xnor U15590 (N_15590,N_15340,N_15494);
and U15591 (N_15591,N_15307,N_15041);
or U15592 (N_15592,N_15008,N_15040);
nor U15593 (N_15593,N_15150,N_15445);
or U15594 (N_15594,N_15256,N_15499);
nand U15595 (N_15595,N_15439,N_15050);
xnor U15596 (N_15596,N_15001,N_15058);
xor U15597 (N_15597,N_15411,N_15335);
xor U15598 (N_15598,N_15000,N_15218);
nand U15599 (N_15599,N_15076,N_15452);
and U15600 (N_15600,N_15486,N_15169);
nor U15601 (N_15601,N_15034,N_15103);
nand U15602 (N_15602,N_15364,N_15376);
nor U15603 (N_15603,N_15207,N_15154);
and U15604 (N_15604,N_15074,N_15036);
or U15605 (N_15605,N_15136,N_15140);
nand U15606 (N_15606,N_15234,N_15434);
nand U15607 (N_15607,N_15361,N_15124);
nor U15608 (N_15608,N_15004,N_15148);
and U15609 (N_15609,N_15062,N_15301);
xnor U15610 (N_15610,N_15282,N_15108);
nor U15611 (N_15611,N_15342,N_15186);
nor U15612 (N_15612,N_15353,N_15240);
nand U15613 (N_15613,N_15064,N_15261);
xor U15614 (N_15614,N_15440,N_15061);
nand U15615 (N_15615,N_15239,N_15474);
nor U15616 (N_15616,N_15490,N_15116);
nand U15617 (N_15617,N_15428,N_15152);
xor U15618 (N_15618,N_15433,N_15291);
or U15619 (N_15619,N_15241,N_15488);
or U15620 (N_15620,N_15070,N_15189);
nor U15621 (N_15621,N_15475,N_15492);
or U15622 (N_15622,N_15030,N_15255);
and U15623 (N_15623,N_15269,N_15031);
and U15624 (N_15624,N_15010,N_15251);
nand U15625 (N_15625,N_15369,N_15168);
xor U15626 (N_15626,N_15022,N_15328);
nor U15627 (N_15627,N_15024,N_15306);
nand U15628 (N_15628,N_15115,N_15346);
or U15629 (N_15629,N_15081,N_15401);
and U15630 (N_15630,N_15144,N_15120);
nand U15631 (N_15631,N_15461,N_15094);
or U15632 (N_15632,N_15011,N_15145);
nor U15633 (N_15633,N_15264,N_15086);
and U15634 (N_15634,N_15014,N_15085);
or U15635 (N_15635,N_15229,N_15194);
nand U15636 (N_15636,N_15288,N_15427);
or U15637 (N_15637,N_15048,N_15092);
xor U15638 (N_15638,N_15319,N_15253);
nand U15639 (N_15639,N_15473,N_15190);
nand U15640 (N_15640,N_15143,N_15226);
nor U15641 (N_15641,N_15156,N_15133);
nand U15642 (N_15642,N_15112,N_15363);
nand U15643 (N_15643,N_15180,N_15320);
or U15644 (N_15644,N_15450,N_15139);
or U15645 (N_15645,N_15444,N_15037);
and U15646 (N_15646,N_15442,N_15158);
nand U15647 (N_15647,N_15313,N_15012);
nor U15648 (N_15648,N_15122,N_15098);
xnor U15649 (N_15649,N_15188,N_15023);
and U15650 (N_15650,N_15449,N_15163);
or U15651 (N_15651,N_15242,N_15332);
xnor U15652 (N_15652,N_15275,N_15027);
or U15653 (N_15653,N_15042,N_15293);
nor U15654 (N_15654,N_15446,N_15408);
or U15655 (N_15655,N_15039,N_15336);
or U15656 (N_15656,N_15491,N_15299);
nor U15657 (N_15657,N_15102,N_15472);
xnor U15658 (N_15658,N_15196,N_15290);
and U15659 (N_15659,N_15247,N_15206);
xor U15660 (N_15660,N_15217,N_15451);
nor U15661 (N_15661,N_15385,N_15177);
nand U15662 (N_15662,N_15292,N_15199);
nor U15663 (N_15663,N_15470,N_15099);
and U15664 (N_15664,N_15005,N_15268);
nand U15665 (N_15665,N_15147,N_15356);
nor U15666 (N_15666,N_15068,N_15021);
xor U15667 (N_15667,N_15141,N_15073);
nand U15668 (N_15668,N_15057,N_15495);
and U15669 (N_15669,N_15493,N_15202);
xor U15670 (N_15670,N_15381,N_15267);
and U15671 (N_15671,N_15038,N_15278);
xnor U15672 (N_15672,N_15402,N_15349);
and U15673 (N_15673,N_15205,N_15254);
xnor U15674 (N_15674,N_15412,N_15453);
or U15675 (N_15675,N_15236,N_15262);
and U15676 (N_15676,N_15383,N_15283);
and U15677 (N_15677,N_15400,N_15302);
and U15678 (N_15678,N_15017,N_15286);
nand U15679 (N_15679,N_15294,N_15223);
and U15680 (N_15680,N_15007,N_15191);
or U15681 (N_15681,N_15225,N_15430);
or U15682 (N_15682,N_15330,N_15109);
or U15683 (N_15683,N_15127,N_15274);
xnor U15684 (N_15684,N_15386,N_15125);
or U15685 (N_15685,N_15077,N_15060);
or U15686 (N_15686,N_15341,N_15423);
xnor U15687 (N_15687,N_15160,N_15246);
and U15688 (N_15688,N_15398,N_15183);
or U15689 (N_15689,N_15015,N_15317);
and U15690 (N_15690,N_15316,N_15489);
and U15691 (N_15691,N_15331,N_15426);
and U15692 (N_15692,N_15404,N_15271);
nor U15693 (N_15693,N_15033,N_15187);
nand U15694 (N_15694,N_15002,N_15315);
or U15695 (N_15695,N_15409,N_15049);
xor U15696 (N_15696,N_15310,N_15289);
nor U15697 (N_15697,N_15425,N_15114);
and U15698 (N_15698,N_15367,N_15337);
and U15699 (N_15699,N_15072,N_15297);
and U15700 (N_15700,N_15478,N_15477);
xnor U15701 (N_15701,N_15497,N_15215);
and U15702 (N_15702,N_15208,N_15155);
or U15703 (N_15703,N_15414,N_15203);
xnor U15704 (N_15704,N_15135,N_15272);
nand U15705 (N_15705,N_15227,N_15204);
nand U15706 (N_15706,N_15355,N_15407);
nand U15707 (N_15707,N_15344,N_15362);
nand U15708 (N_15708,N_15113,N_15101);
or U15709 (N_15709,N_15198,N_15403);
and U15710 (N_15710,N_15378,N_15277);
xor U15711 (N_15711,N_15459,N_15308);
xnor U15712 (N_15712,N_15069,N_15161);
and U15713 (N_15713,N_15333,N_15126);
nand U15714 (N_15714,N_15165,N_15300);
nand U15715 (N_15715,N_15053,N_15329);
or U15716 (N_15716,N_15193,N_15309);
nor U15717 (N_15717,N_15339,N_15280);
xnor U15718 (N_15718,N_15395,N_15216);
nand U15719 (N_15719,N_15028,N_15220);
and U15720 (N_15720,N_15245,N_15379);
xnor U15721 (N_15721,N_15429,N_15424);
or U15722 (N_15722,N_15182,N_15377);
xor U15723 (N_15723,N_15417,N_15312);
and U15724 (N_15724,N_15352,N_15249);
or U15725 (N_15725,N_15397,N_15117);
and U15726 (N_15726,N_15454,N_15065);
nand U15727 (N_15727,N_15260,N_15437);
nand U15728 (N_15728,N_15295,N_15343);
or U15729 (N_15729,N_15044,N_15167);
nand U15730 (N_15730,N_15418,N_15389);
nand U15731 (N_15731,N_15443,N_15162);
nand U15732 (N_15732,N_15130,N_15197);
nand U15733 (N_15733,N_15392,N_15174);
nand U15734 (N_15734,N_15435,N_15237);
and U15735 (N_15735,N_15374,N_15485);
nand U15736 (N_15736,N_15119,N_15219);
or U15737 (N_15737,N_15326,N_15366);
nand U15738 (N_15738,N_15303,N_15399);
xor U15739 (N_15739,N_15347,N_15243);
nor U15740 (N_15740,N_15436,N_15066);
and U15741 (N_15741,N_15138,N_15257);
xnor U15742 (N_15742,N_15083,N_15432);
xnor U15743 (N_15743,N_15487,N_15481);
and U15744 (N_15744,N_15327,N_15059);
xnor U15745 (N_15745,N_15121,N_15462);
nand U15746 (N_15746,N_15185,N_15273);
or U15747 (N_15747,N_15184,N_15175);
nor U15748 (N_15748,N_15153,N_15270);
nor U15749 (N_15749,N_15093,N_15375);
xor U15750 (N_15750,N_15278,N_15230);
nor U15751 (N_15751,N_15448,N_15457);
or U15752 (N_15752,N_15146,N_15317);
and U15753 (N_15753,N_15062,N_15337);
and U15754 (N_15754,N_15235,N_15228);
or U15755 (N_15755,N_15271,N_15460);
and U15756 (N_15756,N_15486,N_15043);
or U15757 (N_15757,N_15188,N_15273);
nor U15758 (N_15758,N_15333,N_15141);
xor U15759 (N_15759,N_15152,N_15457);
and U15760 (N_15760,N_15360,N_15462);
and U15761 (N_15761,N_15102,N_15049);
xnor U15762 (N_15762,N_15488,N_15326);
and U15763 (N_15763,N_15317,N_15114);
and U15764 (N_15764,N_15296,N_15018);
xor U15765 (N_15765,N_15498,N_15437);
or U15766 (N_15766,N_15410,N_15097);
nor U15767 (N_15767,N_15355,N_15309);
xor U15768 (N_15768,N_15149,N_15391);
nand U15769 (N_15769,N_15319,N_15402);
nor U15770 (N_15770,N_15027,N_15159);
nor U15771 (N_15771,N_15000,N_15009);
and U15772 (N_15772,N_15136,N_15119);
nor U15773 (N_15773,N_15365,N_15285);
nand U15774 (N_15774,N_15144,N_15023);
nand U15775 (N_15775,N_15388,N_15421);
xnor U15776 (N_15776,N_15444,N_15380);
xor U15777 (N_15777,N_15423,N_15286);
nor U15778 (N_15778,N_15398,N_15203);
nor U15779 (N_15779,N_15187,N_15209);
nor U15780 (N_15780,N_15301,N_15035);
nand U15781 (N_15781,N_15395,N_15347);
xnor U15782 (N_15782,N_15050,N_15019);
xnor U15783 (N_15783,N_15266,N_15284);
nor U15784 (N_15784,N_15253,N_15361);
and U15785 (N_15785,N_15462,N_15168);
and U15786 (N_15786,N_15212,N_15247);
and U15787 (N_15787,N_15451,N_15336);
nor U15788 (N_15788,N_15020,N_15066);
nor U15789 (N_15789,N_15492,N_15176);
and U15790 (N_15790,N_15115,N_15458);
or U15791 (N_15791,N_15413,N_15285);
and U15792 (N_15792,N_15100,N_15450);
and U15793 (N_15793,N_15147,N_15149);
and U15794 (N_15794,N_15201,N_15441);
xnor U15795 (N_15795,N_15477,N_15432);
nor U15796 (N_15796,N_15036,N_15052);
or U15797 (N_15797,N_15299,N_15497);
or U15798 (N_15798,N_15369,N_15003);
or U15799 (N_15799,N_15419,N_15050);
nor U15800 (N_15800,N_15166,N_15480);
xor U15801 (N_15801,N_15256,N_15176);
nand U15802 (N_15802,N_15226,N_15239);
nand U15803 (N_15803,N_15240,N_15059);
nand U15804 (N_15804,N_15377,N_15381);
and U15805 (N_15805,N_15376,N_15262);
nor U15806 (N_15806,N_15338,N_15101);
nand U15807 (N_15807,N_15340,N_15420);
and U15808 (N_15808,N_15019,N_15186);
or U15809 (N_15809,N_15396,N_15497);
and U15810 (N_15810,N_15429,N_15077);
or U15811 (N_15811,N_15038,N_15270);
nand U15812 (N_15812,N_15185,N_15097);
xor U15813 (N_15813,N_15382,N_15449);
and U15814 (N_15814,N_15162,N_15078);
or U15815 (N_15815,N_15161,N_15118);
and U15816 (N_15816,N_15286,N_15392);
and U15817 (N_15817,N_15460,N_15207);
or U15818 (N_15818,N_15493,N_15461);
or U15819 (N_15819,N_15089,N_15480);
and U15820 (N_15820,N_15362,N_15275);
and U15821 (N_15821,N_15033,N_15403);
nor U15822 (N_15822,N_15272,N_15389);
or U15823 (N_15823,N_15480,N_15390);
xor U15824 (N_15824,N_15334,N_15093);
xnor U15825 (N_15825,N_15007,N_15430);
nor U15826 (N_15826,N_15456,N_15295);
xor U15827 (N_15827,N_15263,N_15012);
xor U15828 (N_15828,N_15065,N_15466);
nor U15829 (N_15829,N_15169,N_15204);
nor U15830 (N_15830,N_15083,N_15039);
and U15831 (N_15831,N_15370,N_15105);
xnor U15832 (N_15832,N_15273,N_15110);
or U15833 (N_15833,N_15082,N_15194);
nor U15834 (N_15834,N_15436,N_15242);
xnor U15835 (N_15835,N_15365,N_15357);
xnor U15836 (N_15836,N_15023,N_15481);
or U15837 (N_15837,N_15219,N_15006);
xor U15838 (N_15838,N_15204,N_15124);
nor U15839 (N_15839,N_15188,N_15097);
and U15840 (N_15840,N_15254,N_15409);
and U15841 (N_15841,N_15217,N_15388);
nor U15842 (N_15842,N_15226,N_15227);
nor U15843 (N_15843,N_15032,N_15287);
nand U15844 (N_15844,N_15385,N_15218);
and U15845 (N_15845,N_15373,N_15239);
xnor U15846 (N_15846,N_15331,N_15230);
and U15847 (N_15847,N_15091,N_15133);
xor U15848 (N_15848,N_15349,N_15353);
or U15849 (N_15849,N_15460,N_15278);
nor U15850 (N_15850,N_15438,N_15131);
and U15851 (N_15851,N_15490,N_15421);
xnor U15852 (N_15852,N_15005,N_15065);
nor U15853 (N_15853,N_15246,N_15356);
or U15854 (N_15854,N_15080,N_15362);
xnor U15855 (N_15855,N_15490,N_15070);
or U15856 (N_15856,N_15241,N_15489);
xnor U15857 (N_15857,N_15166,N_15428);
and U15858 (N_15858,N_15244,N_15059);
or U15859 (N_15859,N_15391,N_15485);
and U15860 (N_15860,N_15121,N_15207);
nand U15861 (N_15861,N_15401,N_15099);
nand U15862 (N_15862,N_15272,N_15308);
xor U15863 (N_15863,N_15149,N_15256);
xor U15864 (N_15864,N_15082,N_15362);
nand U15865 (N_15865,N_15356,N_15079);
nor U15866 (N_15866,N_15025,N_15371);
xnor U15867 (N_15867,N_15492,N_15340);
or U15868 (N_15868,N_15177,N_15411);
nor U15869 (N_15869,N_15417,N_15236);
nor U15870 (N_15870,N_15423,N_15050);
or U15871 (N_15871,N_15301,N_15226);
or U15872 (N_15872,N_15351,N_15188);
nand U15873 (N_15873,N_15188,N_15446);
and U15874 (N_15874,N_15330,N_15113);
and U15875 (N_15875,N_15259,N_15366);
and U15876 (N_15876,N_15247,N_15449);
xnor U15877 (N_15877,N_15229,N_15395);
or U15878 (N_15878,N_15311,N_15215);
or U15879 (N_15879,N_15242,N_15071);
nand U15880 (N_15880,N_15109,N_15232);
nand U15881 (N_15881,N_15346,N_15495);
nand U15882 (N_15882,N_15396,N_15405);
nor U15883 (N_15883,N_15471,N_15333);
nand U15884 (N_15884,N_15196,N_15232);
or U15885 (N_15885,N_15034,N_15039);
and U15886 (N_15886,N_15365,N_15297);
xor U15887 (N_15887,N_15450,N_15182);
or U15888 (N_15888,N_15229,N_15316);
and U15889 (N_15889,N_15068,N_15408);
and U15890 (N_15890,N_15154,N_15377);
nor U15891 (N_15891,N_15344,N_15172);
nor U15892 (N_15892,N_15016,N_15399);
nor U15893 (N_15893,N_15385,N_15060);
or U15894 (N_15894,N_15447,N_15451);
nor U15895 (N_15895,N_15201,N_15357);
xor U15896 (N_15896,N_15425,N_15388);
and U15897 (N_15897,N_15139,N_15074);
or U15898 (N_15898,N_15348,N_15222);
xnor U15899 (N_15899,N_15150,N_15417);
or U15900 (N_15900,N_15223,N_15468);
xnor U15901 (N_15901,N_15426,N_15277);
nor U15902 (N_15902,N_15277,N_15328);
nand U15903 (N_15903,N_15261,N_15385);
xor U15904 (N_15904,N_15078,N_15073);
nor U15905 (N_15905,N_15145,N_15009);
nor U15906 (N_15906,N_15011,N_15370);
nand U15907 (N_15907,N_15180,N_15085);
nand U15908 (N_15908,N_15040,N_15070);
and U15909 (N_15909,N_15379,N_15197);
nor U15910 (N_15910,N_15001,N_15385);
or U15911 (N_15911,N_15080,N_15246);
and U15912 (N_15912,N_15099,N_15365);
xor U15913 (N_15913,N_15337,N_15034);
or U15914 (N_15914,N_15324,N_15305);
nor U15915 (N_15915,N_15467,N_15121);
xnor U15916 (N_15916,N_15067,N_15310);
xnor U15917 (N_15917,N_15210,N_15014);
nor U15918 (N_15918,N_15354,N_15062);
nor U15919 (N_15919,N_15085,N_15335);
and U15920 (N_15920,N_15150,N_15183);
nor U15921 (N_15921,N_15169,N_15083);
nor U15922 (N_15922,N_15180,N_15413);
nand U15923 (N_15923,N_15480,N_15129);
xnor U15924 (N_15924,N_15073,N_15202);
xor U15925 (N_15925,N_15359,N_15466);
and U15926 (N_15926,N_15372,N_15491);
or U15927 (N_15927,N_15099,N_15072);
nand U15928 (N_15928,N_15162,N_15089);
xor U15929 (N_15929,N_15024,N_15016);
xor U15930 (N_15930,N_15077,N_15017);
xnor U15931 (N_15931,N_15129,N_15360);
nor U15932 (N_15932,N_15053,N_15253);
and U15933 (N_15933,N_15297,N_15384);
nand U15934 (N_15934,N_15136,N_15322);
or U15935 (N_15935,N_15065,N_15189);
nand U15936 (N_15936,N_15153,N_15339);
xnor U15937 (N_15937,N_15201,N_15104);
and U15938 (N_15938,N_15403,N_15292);
nor U15939 (N_15939,N_15132,N_15156);
and U15940 (N_15940,N_15419,N_15049);
nand U15941 (N_15941,N_15194,N_15425);
and U15942 (N_15942,N_15041,N_15315);
or U15943 (N_15943,N_15371,N_15202);
nor U15944 (N_15944,N_15000,N_15423);
or U15945 (N_15945,N_15307,N_15257);
or U15946 (N_15946,N_15452,N_15093);
nor U15947 (N_15947,N_15123,N_15209);
and U15948 (N_15948,N_15444,N_15410);
nand U15949 (N_15949,N_15340,N_15189);
and U15950 (N_15950,N_15041,N_15158);
xor U15951 (N_15951,N_15276,N_15310);
nor U15952 (N_15952,N_15135,N_15139);
nor U15953 (N_15953,N_15231,N_15338);
or U15954 (N_15954,N_15413,N_15406);
or U15955 (N_15955,N_15199,N_15215);
xnor U15956 (N_15956,N_15004,N_15328);
nor U15957 (N_15957,N_15125,N_15289);
nor U15958 (N_15958,N_15352,N_15487);
nand U15959 (N_15959,N_15367,N_15228);
or U15960 (N_15960,N_15253,N_15164);
nor U15961 (N_15961,N_15356,N_15131);
nand U15962 (N_15962,N_15396,N_15018);
nor U15963 (N_15963,N_15319,N_15471);
xor U15964 (N_15964,N_15378,N_15473);
nand U15965 (N_15965,N_15407,N_15132);
nand U15966 (N_15966,N_15161,N_15245);
or U15967 (N_15967,N_15187,N_15458);
xnor U15968 (N_15968,N_15171,N_15179);
nor U15969 (N_15969,N_15261,N_15102);
and U15970 (N_15970,N_15336,N_15196);
nand U15971 (N_15971,N_15108,N_15486);
or U15972 (N_15972,N_15162,N_15015);
xor U15973 (N_15973,N_15216,N_15059);
or U15974 (N_15974,N_15105,N_15201);
and U15975 (N_15975,N_15420,N_15228);
xor U15976 (N_15976,N_15465,N_15394);
xor U15977 (N_15977,N_15116,N_15294);
nand U15978 (N_15978,N_15365,N_15069);
nand U15979 (N_15979,N_15233,N_15442);
nand U15980 (N_15980,N_15493,N_15463);
or U15981 (N_15981,N_15187,N_15164);
nor U15982 (N_15982,N_15090,N_15209);
nand U15983 (N_15983,N_15479,N_15448);
xor U15984 (N_15984,N_15123,N_15028);
or U15985 (N_15985,N_15232,N_15471);
nor U15986 (N_15986,N_15327,N_15068);
xor U15987 (N_15987,N_15267,N_15441);
nor U15988 (N_15988,N_15407,N_15024);
and U15989 (N_15989,N_15005,N_15399);
xnor U15990 (N_15990,N_15351,N_15185);
or U15991 (N_15991,N_15441,N_15004);
xor U15992 (N_15992,N_15113,N_15143);
or U15993 (N_15993,N_15198,N_15279);
xnor U15994 (N_15994,N_15401,N_15360);
or U15995 (N_15995,N_15085,N_15141);
and U15996 (N_15996,N_15148,N_15388);
or U15997 (N_15997,N_15168,N_15025);
nand U15998 (N_15998,N_15359,N_15353);
and U15999 (N_15999,N_15116,N_15434);
or U16000 (N_16000,N_15711,N_15809);
and U16001 (N_16001,N_15559,N_15771);
and U16002 (N_16002,N_15694,N_15787);
xor U16003 (N_16003,N_15586,N_15639);
xnor U16004 (N_16004,N_15732,N_15858);
or U16005 (N_16005,N_15981,N_15561);
nor U16006 (N_16006,N_15661,N_15897);
nor U16007 (N_16007,N_15828,N_15812);
nor U16008 (N_16008,N_15999,N_15529);
nor U16009 (N_16009,N_15862,N_15595);
and U16010 (N_16010,N_15650,N_15912);
nor U16011 (N_16011,N_15686,N_15930);
and U16012 (N_16012,N_15986,N_15863);
nor U16013 (N_16013,N_15870,N_15721);
xnor U16014 (N_16014,N_15868,N_15923);
xnor U16015 (N_16015,N_15502,N_15903);
nor U16016 (N_16016,N_15937,N_15767);
xnor U16017 (N_16017,N_15844,N_15867);
xor U16018 (N_16018,N_15548,N_15904);
or U16019 (N_16019,N_15552,N_15616);
xnor U16020 (N_16020,N_15683,N_15663);
nand U16021 (N_16021,N_15672,N_15971);
nand U16022 (N_16022,N_15608,N_15703);
and U16023 (N_16023,N_15582,N_15806);
nand U16024 (N_16024,N_15519,N_15525);
and U16025 (N_16025,N_15564,N_15871);
nor U16026 (N_16026,N_15766,N_15651);
nand U16027 (N_16027,N_15562,N_15827);
or U16028 (N_16028,N_15964,N_15638);
or U16029 (N_16029,N_15501,N_15509);
or U16030 (N_16030,N_15810,N_15983);
or U16031 (N_16031,N_15852,N_15697);
and U16032 (N_16032,N_15829,N_15953);
nand U16033 (N_16033,N_15647,N_15584);
xnor U16034 (N_16034,N_15790,N_15688);
or U16035 (N_16035,N_15706,N_15585);
and U16036 (N_16036,N_15955,N_15624);
nor U16037 (N_16037,N_15774,N_15982);
or U16038 (N_16038,N_15795,N_15611);
xnor U16039 (N_16039,N_15883,N_15918);
nand U16040 (N_16040,N_15554,N_15682);
and U16041 (N_16041,N_15752,N_15521);
nand U16042 (N_16042,N_15635,N_15792);
or U16043 (N_16043,N_15640,N_15784);
nor U16044 (N_16044,N_15832,N_15908);
or U16045 (N_16045,N_15876,N_15615);
or U16046 (N_16046,N_15880,N_15737);
xnor U16047 (N_16047,N_15833,N_15655);
nor U16048 (N_16048,N_15807,N_15726);
and U16049 (N_16049,N_15882,N_15736);
xnor U16050 (N_16050,N_15541,N_15928);
and U16051 (N_16051,N_15596,N_15756);
nand U16052 (N_16052,N_15765,N_15836);
xnor U16053 (N_16053,N_15580,N_15602);
xnor U16054 (N_16054,N_15619,N_15546);
nand U16055 (N_16055,N_15738,N_15961);
nor U16056 (N_16056,N_15909,N_15759);
xnor U16057 (N_16057,N_15991,N_15948);
or U16058 (N_16058,N_15947,N_15779);
nand U16059 (N_16059,N_15671,N_15536);
or U16060 (N_16060,N_15796,N_15594);
nor U16061 (N_16061,N_15527,N_15845);
nand U16062 (N_16062,N_15704,N_15893);
xor U16063 (N_16063,N_15593,N_15646);
nand U16064 (N_16064,N_15813,N_15530);
nor U16065 (N_16065,N_15659,N_15621);
or U16066 (N_16066,N_15718,N_15926);
xnor U16067 (N_16067,N_15811,N_15526);
nor U16068 (N_16068,N_15735,N_15895);
and U16069 (N_16069,N_15588,N_15547);
nand U16070 (N_16070,N_15850,N_15700);
and U16071 (N_16071,N_15653,N_15920);
nor U16072 (N_16072,N_15570,N_15549);
nand U16073 (N_16073,N_15855,N_15587);
nor U16074 (N_16074,N_15965,N_15834);
xnor U16075 (N_16075,N_15943,N_15872);
nor U16076 (N_16076,N_15719,N_15709);
xnor U16077 (N_16077,N_15517,N_15627);
nand U16078 (N_16078,N_15927,N_15949);
nor U16079 (N_16079,N_15980,N_15932);
nand U16080 (N_16080,N_15710,N_15819);
nor U16081 (N_16081,N_15538,N_15601);
xor U16082 (N_16082,N_15695,N_15881);
or U16083 (N_16083,N_15551,N_15696);
nand U16084 (N_16084,N_15540,N_15757);
and U16085 (N_16085,N_15625,N_15618);
nor U16086 (N_16086,N_15569,N_15575);
or U16087 (N_16087,N_15960,N_15783);
nor U16088 (N_16088,N_15905,N_15693);
nor U16089 (N_16089,N_15523,N_15793);
and U16090 (N_16090,N_15591,N_15839);
xnor U16091 (N_16091,N_15684,N_15959);
nand U16092 (N_16092,N_15919,N_15861);
and U16093 (N_16093,N_15555,N_15531);
xor U16094 (N_16094,N_15702,N_15885);
nor U16095 (N_16095,N_15835,N_15542);
nor U16096 (N_16096,N_15707,N_15817);
or U16097 (N_16097,N_15823,N_15579);
nor U16098 (N_16098,N_15724,N_15689);
nor U16099 (N_16099,N_15984,N_15634);
nand U16100 (N_16100,N_15990,N_15853);
nand U16101 (N_16101,N_15749,N_15713);
or U16102 (N_16102,N_15950,N_15856);
or U16103 (N_16103,N_15753,N_15632);
nand U16104 (N_16104,N_15763,N_15637);
nor U16105 (N_16105,N_15565,N_15864);
nand U16106 (N_16106,N_15667,N_15566);
nand U16107 (N_16107,N_15642,N_15681);
nand U16108 (N_16108,N_15644,N_15906);
or U16109 (N_16109,N_15989,N_15875);
and U16110 (N_16110,N_15788,N_15645);
or U16111 (N_16111,N_15613,N_15831);
xnor U16112 (N_16112,N_15929,N_15623);
nor U16113 (N_16113,N_15946,N_15820);
nor U16114 (N_16114,N_15939,N_15915);
nor U16115 (N_16115,N_15717,N_15781);
or U16116 (N_16116,N_15972,N_15922);
nor U16117 (N_16117,N_15898,N_15544);
nor U16118 (N_16118,N_15612,N_15680);
xor U16119 (N_16119,N_15901,N_15600);
xor U16120 (N_16120,N_15968,N_15698);
and U16121 (N_16121,N_15957,N_15954);
nor U16122 (N_16122,N_15803,N_15974);
or U16123 (N_16123,N_15840,N_15510);
or U16124 (N_16124,N_15670,N_15533);
and U16125 (N_16125,N_15979,N_15687);
nand U16126 (N_16126,N_15516,N_15677);
nand U16127 (N_16127,N_15617,N_15630);
and U16128 (N_16128,N_15535,N_15992);
or U16129 (N_16129,N_15818,N_15805);
and U16130 (N_16130,N_15631,N_15679);
or U16131 (N_16131,N_15673,N_15592);
and U16132 (N_16132,N_15537,N_15761);
or U16133 (N_16133,N_15748,N_15925);
or U16134 (N_16134,N_15857,N_15899);
nor U16135 (N_16135,N_15648,N_15916);
and U16136 (N_16136,N_15628,N_15520);
or U16137 (N_16137,N_15951,N_15636);
and U16138 (N_16138,N_15866,N_15692);
or U16139 (N_16139,N_15626,N_15825);
nand U16140 (N_16140,N_15914,N_15824);
nand U16141 (N_16141,N_15902,N_15567);
nand U16142 (N_16142,N_15607,N_15800);
xor U16143 (N_16143,N_15599,N_15690);
or U16144 (N_16144,N_15515,N_15563);
nand U16145 (N_16145,N_15892,N_15878);
xor U16146 (N_16146,N_15782,N_15814);
nor U16147 (N_16147,N_15775,N_15723);
xnor U16148 (N_16148,N_15963,N_15791);
nand U16149 (N_16149,N_15604,N_15851);
xor U16150 (N_16150,N_15772,N_15854);
and U16151 (N_16151,N_15750,N_15553);
nand U16152 (N_16152,N_15797,N_15712);
xnor U16153 (N_16153,N_15799,N_15708);
and U16154 (N_16154,N_15973,N_15747);
xnor U16155 (N_16155,N_15879,N_15933);
xor U16156 (N_16156,N_15610,N_15508);
xnor U16157 (N_16157,N_15940,N_15729);
nor U16158 (N_16158,N_15865,N_15576);
and U16159 (N_16159,N_15841,N_15597);
and U16160 (N_16160,N_15622,N_15745);
or U16161 (N_16161,N_15847,N_15921);
nor U16162 (N_16162,N_15573,N_15913);
xnor U16163 (N_16163,N_15746,N_15987);
nand U16164 (N_16164,N_15997,N_15741);
nand U16165 (N_16165,N_15666,N_15568);
xnor U16166 (N_16166,N_15603,N_15975);
nor U16167 (N_16167,N_15822,N_15837);
and U16168 (N_16168,N_15518,N_15821);
and U16169 (N_16169,N_15994,N_15534);
and U16170 (N_16170,N_15924,N_15804);
and U16171 (N_16171,N_15641,N_15764);
xnor U16172 (N_16172,N_15649,N_15891);
xor U16173 (N_16173,N_15993,N_15941);
and U16174 (N_16174,N_15558,N_15578);
nor U16175 (N_16175,N_15557,N_15846);
and U16176 (N_16176,N_15614,N_15751);
or U16177 (N_16177,N_15877,N_15572);
nand U16178 (N_16178,N_15522,N_15869);
nand U16179 (N_16179,N_15755,N_15900);
or U16180 (N_16180,N_15896,N_15571);
or U16181 (N_16181,N_15577,N_15581);
xnor U16182 (N_16182,N_15754,N_15938);
and U16183 (N_16183,N_15590,N_15785);
xnor U16184 (N_16184,N_15705,N_15716);
nor U16185 (N_16185,N_15652,N_15816);
nor U16186 (N_16186,N_15894,N_15727);
nand U16187 (N_16187,N_15715,N_15760);
xor U16188 (N_16188,N_15956,N_15773);
and U16189 (N_16189,N_15633,N_15660);
and U16190 (N_16190,N_15911,N_15794);
nor U16191 (N_16191,N_15998,N_15675);
nand U16192 (N_16192,N_15665,N_15886);
xnor U16193 (N_16193,N_15976,N_15743);
or U16194 (N_16194,N_15731,N_15643);
and U16195 (N_16195,N_15656,N_15815);
or U16196 (N_16196,N_15884,N_15550);
nand U16197 (N_16197,N_15931,N_15777);
nand U16198 (N_16198,N_15744,N_15657);
or U16199 (N_16199,N_15668,N_15511);
nor U16200 (N_16200,N_15978,N_15967);
and U16201 (N_16201,N_15539,N_15532);
nor U16202 (N_16202,N_15917,N_15504);
nand U16203 (N_16203,N_15560,N_15942);
xor U16204 (N_16204,N_15730,N_15770);
or U16205 (N_16205,N_15583,N_15514);
and U16206 (N_16206,N_15739,N_15740);
nor U16207 (N_16207,N_15524,N_15944);
or U16208 (N_16208,N_15969,N_15988);
xnor U16209 (N_16209,N_15620,N_15658);
xor U16210 (N_16210,N_15888,N_15685);
or U16211 (N_16211,N_15733,N_15699);
and U16212 (N_16212,N_15606,N_15889);
xnor U16213 (N_16213,N_15500,N_15503);
nand U16214 (N_16214,N_15936,N_15589);
and U16215 (N_16215,N_15506,N_15662);
nor U16216 (N_16216,N_15890,N_15776);
nor U16217 (N_16217,N_15762,N_15664);
nand U16218 (N_16218,N_15691,N_15808);
nor U16219 (N_16219,N_15966,N_15722);
and U16220 (N_16220,N_15801,N_15874);
and U16221 (N_16221,N_15678,N_15742);
nor U16222 (N_16222,N_15545,N_15676);
xor U16223 (N_16223,N_15907,N_15887);
or U16224 (N_16224,N_15843,N_15505);
xor U16225 (N_16225,N_15977,N_15654);
xor U16226 (N_16226,N_15728,N_15945);
and U16227 (N_16227,N_15669,N_15720);
or U16228 (N_16228,N_15802,N_15838);
nor U16229 (N_16229,N_15725,N_15789);
or U16230 (N_16230,N_15512,N_15935);
and U16231 (N_16231,N_15556,N_15786);
or U16232 (N_16232,N_15970,N_15701);
or U16233 (N_16233,N_15958,N_15985);
xnor U16234 (N_16234,N_15848,N_15768);
and U16235 (N_16235,N_15996,N_15910);
nor U16236 (N_16236,N_15605,N_15528);
nor U16237 (N_16237,N_15873,N_15629);
nand U16238 (N_16238,N_15609,N_15962);
or U16239 (N_16239,N_15598,N_15842);
and U16240 (N_16240,N_15758,N_15859);
and U16241 (N_16241,N_15798,N_15826);
nand U16242 (N_16242,N_15769,N_15860);
nor U16243 (N_16243,N_15734,N_15674);
nand U16244 (N_16244,N_15714,N_15513);
xnor U16245 (N_16245,N_15507,N_15934);
and U16246 (N_16246,N_15849,N_15780);
or U16247 (N_16247,N_15778,N_15830);
nand U16248 (N_16248,N_15995,N_15574);
or U16249 (N_16249,N_15543,N_15952);
and U16250 (N_16250,N_15884,N_15558);
nor U16251 (N_16251,N_15573,N_15622);
or U16252 (N_16252,N_15519,N_15621);
or U16253 (N_16253,N_15913,N_15681);
xor U16254 (N_16254,N_15823,N_15959);
nor U16255 (N_16255,N_15709,N_15850);
nor U16256 (N_16256,N_15685,N_15629);
xor U16257 (N_16257,N_15623,N_15632);
and U16258 (N_16258,N_15998,N_15514);
xnor U16259 (N_16259,N_15735,N_15809);
or U16260 (N_16260,N_15560,N_15500);
nand U16261 (N_16261,N_15680,N_15884);
and U16262 (N_16262,N_15889,N_15551);
or U16263 (N_16263,N_15773,N_15731);
xor U16264 (N_16264,N_15701,N_15536);
xor U16265 (N_16265,N_15911,N_15960);
and U16266 (N_16266,N_15883,N_15851);
xnor U16267 (N_16267,N_15889,N_15883);
nand U16268 (N_16268,N_15686,N_15611);
xnor U16269 (N_16269,N_15793,N_15783);
nor U16270 (N_16270,N_15847,N_15533);
nor U16271 (N_16271,N_15554,N_15690);
xor U16272 (N_16272,N_15634,N_15518);
xor U16273 (N_16273,N_15728,N_15869);
nand U16274 (N_16274,N_15843,N_15894);
and U16275 (N_16275,N_15836,N_15594);
nor U16276 (N_16276,N_15828,N_15945);
or U16277 (N_16277,N_15808,N_15835);
xor U16278 (N_16278,N_15524,N_15766);
nor U16279 (N_16279,N_15706,N_15934);
xnor U16280 (N_16280,N_15648,N_15626);
xnor U16281 (N_16281,N_15553,N_15867);
nor U16282 (N_16282,N_15912,N_15713);
or U16283 (N_16283,N_15502,N_15760);
nor U16284 (N_16284,N_15892,N_15662);
xor U16285 (N_16285,N_15932,N_15548);
xnor U16286 (N_16286,N_15948,N_15732);
xor U16287 (N_16287,N_15991,N_15573);
xnor U16288 (N_16288,N_15591,N_15532);
and U16289 (N_16289,N_15941,N_15667);
xor U16290 (N_16290,N_15664,N_15612);
nand U16291 (N_16291,N_15797,N_15745);
nand U16292 (N_16292,N_15709,N_15570);
and U16293 (N_16293,N_15646,N_15633);
xnor U16294 (N_16294,N_15513,N_15734);
xor U16295 (N_16295,N_15777,N_15853);
nand U16296 (N_16296,N_15598,N_15622);
xor U16297 (N_16297,N_15761,N_15828);
nor U16298 (N_16298,N_15834,N_15652);
nand U16299 (N_16299,N_15690,N_15729);
and U16300 (N_16300,N_15529,N_15670);
xor U16301 (N_16301,N_15685,N_15543);
or U16302 (N_16302,N_15653,N_15716);
xnor U16303 (N_16303,N_15841,N_15742);
nor U16304 (N_16304,N_15872,N_15618);
and U16305 (N_16305,N_15550,N_15624);
and U16306 (N_16306,N_15646,N_15658);
nor U16307 (N_16307,N_15864,N_15702);
nor U16308 (N_16308,N_15970,N_15816);
xor U16309 (N_16309,N_15641,N_15961);
nand U16310 (N_16310,N_15601,N_15508);
or U16311 (N_16311,N_15976,N_15608);
nand U16312 (N_16312,N_15574,N_15958);
and U16313 (N_16313,N_15893,N_15781);
xor U16314 (N_16314,N_15876,N_15767);
xnor U16315 (N_16315,N_15969,N_15992);
nand U16316 (N_16316,N_15973,N_15716);
nor U16317 (N_16317,N_15584,N_15874);
xnor U16318 (N_16318,N_15781,N_15549);
nor U16319 (N_16319,N_15671,N_15990);
nor U16320 (N_16320,N_15813,N_15843);
nand U16321 (N_16321,N_15926,N_15976);
xor U16322 (N_16322,N_15586,N_15799);
xnor U16323 (N_16323,N_15542,N_15696);
or U16324 (N_16324,N_15509,N_15879);
nand U16325 (N_16325,N_15615,N_15669);
xor U16326 (N_16326,N_15516,N_15851);
nand U16327 (N_16327,N_15769,N_15993);
xnor U16328 (N_16328,N_15808,N_15667);
nand U16329 (N_16329,N_15703,N_15508);
nor U16330 (N_16330,N_15952,N_15659);
and U16331 (N_16331,N_15881,N_15620);
or U16332 (N_16332,N_15683,N_15636);
or U16333 (N_16333,N_15797,N_15943);
nand U16334 (N_16334,N_15519,N_15666);
or U16335 (N_16335,N_15967,N_15837);
or U16336 (N_16336,N_15549,N_15801);
and U16337 (N_16337,N_15661,N_15781);
or U16338 (N_16338,N_15727,N_15556);
or U16339 (N_16339,N_15997,N_15515);
and U16340 (N_16340,N_15790,N_15751);
xor U16341 (N_16341,N_15972,N_15599);
nor U16342 (N_16342,N_15642,N_15721);
and U16343 (N_16343,N_15521,N_15568);
xor U16344 (N_16344,N_15815,N_15757);
and U16345 (N_16345,N_15726,N_15541);
nand U16346 (N_16346,N_15841,N_15944);
nand U16347 (N_16347,N_15938,N_15714);
xor U16348 (N_16348,N_15925,N_15766);
nand U16349 (N_16349,N_15692,N_15519);
nor U16350 (N_16350,N_15574,N_15867);
and U16351 (N_16351,N_15801,N_15512);
nand U16352 (N_16352,N_15938,N_15748);
xnor U16353 (N_16353,N_15634,N_15654);
and U16354 (N_16354,N_15560,N_15979);
xnor U16355 (N_16355,N_15699,N_15937);
nand U16356 (N_16356,N_15566,N_15786);
and U16357 (N_16357,N_15921,N_15844);
xor U16358 (N_16358,N_15729,N_15784);
and U16359 (N_16359,N_15834,N_15536);
nor U16360 (N_16360,N_15869,N_15576);
and U16361 (N_16361,N_15842,N_15571);
and U16362 (N_16362,N_15522,N_15801);
and U16363 (N_16363,N_15818,N_15769);
or U16364 (N_16364,N_15808,N_15544);
nand U16365 (N_16365,N_15516,N_15779);
and U16366 (N_16366,N_15796,N_15821);
or U16367 (N_16367,N_15968,N_15947);
and U16368 (N_16368,N_15921,N_15894);
xor U16369 (N_16369,N_15831,N_15646);
and U16370 (N_16370,N_15841,N_15521);
nand U16371 (N_16371,N_15603,N_15565);
and U16372 (N_16372,N_15890,N_15962);
nor U16373 (N_16373,N_15725,N_15648);
xor U16374 (N_16374,N_15913,N_15861);
nor U16375 (N_16375,N_15921,N_15660);
or U16376 (N_16376,N_15562,N_15925);
and U16377 (N_16377,N_15683,N_15773);
nand U16378 (N_16378,N_15821,N_15736);
xor U16379 (N_16379,N_15978,N_15540);
xor U16380 (N_16380,N_15926,N_15605);
nand U16381 (N_16381,N_15655,N_15550);
or U16382 (N_16382,N_15894,N_15866);
xor U16383 (N_16383,N_15576,N_15647);
xnor U16384 (N_16384,N_15507,N_15804);
nand U16385 (N_16385,N_15970,N_15629);
nand U16386 (N_16386,N_15701,N_15835);
or U16387 (N_16387,N_15803,N_15548);
or U16388 (N_16388,N_15607,N_15627);
or U16389 (N_16389,N_15636,N_15518);
nor U16390 (N_16390,N_15706,N_15889);
xnor U16391 (N_16391,N_15866,N_15671);
nor U16392 (N_16392,N_15500,N_15811);
nand U16393 (N_16393,N_15635,N_15706);
nor U16394 (N_16394,N_15649,N_15752);
nand U16395 (N_16395,N_15593,N_15938);
or U16396 (N_16396,N_15888,N_15905);
nand U16397 (N_16397,N_15765,N_15698);
nor U16398 (N_16398,N_15915,N_15944);
nand U16399 (N_16399,N_15717,N_15563);
or U16400 (N_16400,N_15899,N_15708);
nand U16401 (N_16401,N_15826,N_15809);
nand U16402 (N_16402,N_15894,N_15979);
and U16403 (N_16403,N_15877,N_15953);
xnor U16404 (N_16404,N_15665,N_15509);
and U16405 (N_16405,N_15626,N_15628);
nand U16406 (N_16406,N_15829,N_15606);
nor U16407 (N_16407,N_15661,N_15806);
nand U16408 (N_16408,N_15873,N_15661);
or U16409 (N_16409,N_15705,N_15540);
and U16410 (N_16410,N_15573,N_15786);
xnor U16411 (N_16411,N_15642,N_15816);
xor U16412 (N_16412,N_15756,N_15508);
nor U16413 (N_16413,N_15793,N_15626);
or U16414 (N_16414,N_15682,N_15511);
nor U16415 (N_16415,N_15704,N_15599);
xnor U16416 (N_16416,N_15525,N_15672);
nand U16417 (N_16417,N_15720,N_15709);
xnor U16418 (N_16418,N_15532,N_15503);
and U16419 (N_16419,N_15520,N_15908);
and U16420 (N_16420,N_15534,N_15825);
nor U16421 (N_16421,N_15760,N_15518);
xnor U16422 (N_16422,N_15567,N_15501);
or U16423 (N_16423,N_15566,N_15515);
xor U16424 (N_16424,N_15847,N_15934);
xnor U16425 (N_16425,N_15954,N_15535);
nor U16426 (N_16426,N_15938,N_15540);
xor U16427 (N_16427,N_15850,N_15785);
nor U16428 (N_16428,N_15980,N_15930);
xnor U16429 (N_16429,N_15675,N_15864);
or U16430 (N_16430,N_15600,N_15618);
xnor U16431 (N_16431,N_15793,N_15680);
nor U16432 (N_16432,N_15795,N_15538);
nand U16433 (N_16433,N_15770,N_15872);
xnor U16434 (N_16434,N_15941,N_15699);
xnor U16435 (N_16435,N_15900,N_15881);
nand U16436 (N_16436,N_15922,N_15648);
nand U16437 (N_16437,N_15743,N_15996);
and U16438 (N_16438,N_15657,N_15738);
nand U16439 (N_16439,N_15778,N_15982);
nor U16440 (N_16440,N_15752,N_15749);
nor U16441 (N_16441,N_15545,N_15916);
and U16442 (N_16442,N_15895,N_15807);
and U16443 (N_16443,N_15923,N_15792);
nand U16444 (N_16444,N_15878,N_15766);
nand U16445 (N_16445,N_15903,N_15546);
xor U16446 (N_16446,N_15694,N_15730);
nand U16447 (N_16447,N_15777,N_15996);
or U16448 (N_16448,N_15914,N_15809);
or U16449 (N_16449,N_15668,N_15808);
nor U16450 (N_16450,N_15685,N_15660);
nor U16451 (N_16451,N_15782,N_15502);
and U16452 (N_16452,N_15654,N_15528);
xnor U16453 (N_16453,N_15916,N_15882);
and U16454 (N_16454,N_15723,N_15690);
xnor U16455 (N_16455,N_15590,N_15711);
and U16456 (N_16456,N_15908,N_15531);
nand U16457 (N_16457,N_15698,N_15586);
xnor U16458 (N_16458,N_15881,N_15877);
and U16459 (N_16459,N_15583,N_15746);
xor U16460 (N_16460,N_15969,N_15983);
nand U16461 (N_16461,N_15714,N_15987);
xor U16462 (N_16462,N_15534,N_15852);
nor U16463 (N_16463,N_15728,N_15861);
or U16464 (N_16464,N_15847,N_15739);
or U16465 (N_16465,N_15764,N_15505);
xor U16466 (N_16466,N_15543,N_15740);
and U16467 (N_16467,N_15887,N_15894);
nand U16468 (N_16468,N_15636,N_15801);
nor U16469 (N_16469,N_15884,N_15693);
xor U16470 (N_16470,N_15961,N_15542);
nor U16471 (N_16471,N_15557,N_15760);
nor U16472 (N_16472,N_15668,N_15924);
xnor U16473 (N_16473,N_15871,N_15695);
nor U16474 (N_16474,N_15721,N_15727);
xor U16475 (N_16475,N_15548,N_15955);
xor U16476 (N_16476,N_15978,N_15656);
nand U16477 (N_16477,N_15579,N_15782);
xor U16478 (N_16478,N_15516,N_15774);
and U16479 (N_16479,N_15941,N_15773);
xnor U16480 (N_16480,N_15729,N_15934);
nand U16481 (N_16481,N_15698,N_15869);
xor U16482 (N_16482,N_15746,N_15761);
nand U16483 (N_16483,N_15650,N_15829);
and U16484 (N_16484,N_15714,N_15876);
nor U16485 (N_16485,N_15522,N_15999);
nand U16486 (N_16486,N_15779,N_15988);
and U16487 (N_16487,N_15824,N_15801);
xnor U16488 (N_16488,N_15837,N_15667);
xor U16489 (N_16489,N_15808,N_15678);
nor U16490 (N_16490,N_15723,N_15569);
xor U16491 (N_16491,N_15806,N_15748);
or U16492 (N_16492,N_15993,N_15551);
or U16493 (N_16493,N_15801,N_15711);
nand U16494 (N_16494,N_15770,N_15930);
and U16495 (N_16495,N_15533,N_15942);
nor U16496 (N_16496,N_15539,N_15725);
nand U16497 (N_16497,N_15531,N_15850);
or U16498 (N_16498,N_15941,N_15760);
nand U16499 (N_16499,N_15768,N_15807);
nand U16500 (N_16500,N_16140,N_16282);
nor U16501 (N_16501,N_16236,N_16286);
and U16502 (N_16502,N_16135,N_16494);
xor U16503 (N_16503,N_16249,N_16237);
nor U16504 (N_16504,N_16288,N_16052);
nand U16505 (N_16505,N_16074,N_16318);
xor U16506 (N_16506,N_16424,N_16376);
or U16507 (N_16507,N_16014,N_16253);
xor U16508 (N_16508,N_16324,N_16361);
nand U16509 (N_16509,N_16468,N_16363);
or U16510 (N_16510,N_16228,N_16146);
and U16511 (N_16511,N_16188,N_16438);
and U16512 (N_16512,N_16484,N_16496);
nand U16513 (N_16513,N_16099,N_16442);
or U16514 (N_16514,N_16157,N_16113);
or U16515 (N_16515,N_16230,N_16061);
xor U16516 (N_16516,N_16184,N_16243);
or U16517 (N_16517,N_16434,N_16202);
nand U16518 (N_16518,N_16083,N_16490);
nor U16519 (N_16519,N_16463,N_16458);
or U16520 (N_16520,N_16109,N_16275);
nor U16521 (N_16521,N_16255,N_16080);
and U16522 (N_16522,N_16136,N_16160);
nor U16523 (N_16523,N_16030,N_16142);
and U16524 (N_16524,N_16345,N_16467);
and U16525 (N_16525,N_16077,N_16343);
and U16526 (N_16526,N_16280,N_16180);
xor U16527 (N_16527,N_16312,N_16357);
xor U16528 (N_16528,N_16290,N_16491);
or U16529 (N_16529,N_16398,N_16394);
nor U16530 (N_16530,N_16093,N_16384);
nand U16531 (N_16531,N_16443,N_16487);
xnor U16532 (N_16532,N_16067,N_16094);
and U16533 (N_16533,N_16486,N_16265);
and U16534 (N_16534,N_16181,N_16322);
or U16535 (N_16535,N_16276,N_16219);
nor U16536 (N_16536,N_16015,N_16214);
xor U16537 (N_16537,N_16153,N_16409);
or U16538 (N_16538,N_16155,N_16303);
and U16539 (N_16539,N_16241,N_16270);
and U16540 (N_16540,N_16017,N_16063);
nand U16541 (N_16541,N_16207,N_16375);
xnor U16542 (N_16542,N_16182,N_16003);
xnor U16543 (N_16543,N_16302,N_16267);
xnor U16544 (N_16544,N_16386,N_16464);
xor U16545 (N_16545,N_16366,N_16441);
or U16546 (N_16546,N_16308,N_16450);
or U16547 (N_16547,N_16435,N_16341);
and U16548 (N_16548,N_16478,N_16189);
nor U16549 (N_16549,N_16006,N_16119);
or U16550 (N_16550,N_16277,N_16232);
nor U16551 (N_16551,N_16351,N_16473);
and U16552 (N_16552,N_16414,N_16362);
and U16553 (N_16553,N_16165,N_16066);
xor U16554 (N_16554,N_16416,N_16148);
nor U16555 (N_16555,N_16060,N_16129);
nor U16556 (N_16556,N_16258,N_16498);
nor U16557 (N_16557,N_16321,N_16381);
xnor U16558 (N_16558,N_16462,N_16400);
nor U16559 (N_16559,N_16021,N_16311);
or U16560 (N_16560,N_16242,N_16370);
nor U16561 (N_16561,N_16102,N_16421);
xor U16562 (N_16562,N_16070,N_16103);
nor U16563 (N_16563,N_16296,N_16143);
or U16564 (N_16564,N_16340,N_16183);
xnor U16565 (N_16565,N_16372,N_16257);
nor U16566 (N_16566,N_16331,N_16396);
nor U16567 (N_16567,N_16088,N_16195);
xnor U16568 (N_16568,N_16037,N_16062);
or U16569 (N_16569,N_16256,N_16047);
xnor U16570 (N_16570,N_16447,N_16069);
and U16571 (N_16571,N_16422,N_16344);
nand U16572 (N_16572,N_16432,N_16065);
xor U16573 (N_16573,N_16029,N_16134);
nand U16574 (N_16574,N_16440,N_16389);
and U16575 (N_16575,N_16115,N_16141);
and U16576 (N_16576,N_16173,N_16378);
xor U16577 (N_16577,N_16128,N_16336);
xor U16578 (N_16578,N_16012,N_16335);
nand U16579 (N_16579,N_16114,N_16079);
xnor U16580 (N_16580,N_16299,N_16263);
nor U16581 (N_16581,N_16055,N_16091);
nand U16582 (N_16582,N_16377,N_16216);
nand U16583 (N_16583,N_16224,N_16225);
xnor U16584 (N_16584,N_16198,N_16399);
and U16585 (N_16585,N_16315,N_16050);
nand U16586 (N_16586,N_16108,N_16352);
nor U16587 (N_16587,N_16279,N_16385);
or U16588 (N_16588,N_16368,N_16301);
nand U16589 (N_16589,N_16338,N_16185);
nor U16590 (N_16590,N_16412,N_16053);
or U16591 (N_16591,N_16456,N_16110);
nand U16592 (N_16592,N_16425,N_16085);
xnor U16593 (N_16593,N_16056,N_16204);
nand U16594 (N_16594,N_16127,N_16126);
nor U16595 (N_16595,N_16426,N_16310);
or U16596 (N_16596,N_16297,N_16035);
nand U16597 (N_16597,N_16223,N_16164);
xnor U16598 (N_16598,N_16227,N_16167);
or U16599 (N_16599,N_16367,N_16355);
or U16600 (N_16600,N_16213,N_16316);
or U16601 (N_16601,N_16120,N_16009);
xnor U16602 (N_16602,N_16457,N_16293);
and U16603 (N_16603,N_16098,N_16347);
or U16604 (N_16604,N_16323,N_16350);
xnor U16605 (N_16605,N_16139,N_16395);
xnor U16606 (N_16606,N_16268,N_16187);
or U16607 (N_16607,N_16097,N_16123);
and U16608 (N_16608,N_16031,N_16452);
or U16609 (N_16609,N_16483,N_16479);
and U16610 (N_16610,N_16049,N_16383);
nand U16611 (N_16611,N_16033,N_16392);
or U16612 (N_16612,N_16419,N_16229);
and U16613 (N_16613,N_16481,N_16446);
nand U16614 (N_16614,N_16169,N_16266);
and U16615 (N_16615,N_16238,N_16106);
or U16616 (N_16616,N_16292,N_16489);
and U16617 (N_16617,N_16272,N_16420);
nor U16618 (N_16618,N_16281,N_16240);
nor U16619 (N_16619,N_16057,N_16154);
and U16620 (N_16620,N_16246,N_16245);
nand U16621 (N_16621,N_16171,N_16313);
and U16622 (N_16622,N_16453,N_16048);
xnor U16623 (N_16623,N_16449,N_16125);
and U16624 (N_16624,N_16177,N_16284);
xnor U16625 (N_16625,N_16193,N_16418);
xor U16626 (N_16626,N_16178,N_16101);
or U16627 (N_16627,N_16248,N_16360);
nand U16628 (N_16628,N_16333,N_16273);
or U16629 (N_16629,N_16170,N_16118);
xnor U16630 (N_16630,N_16051,N_16064);
xnor U16631 (N_16631,N_16317,N_16078);
nor U16632 (N_16632,N_16095,N_16206);
or U16633 (N_16633,N_16320,N_16104);
nor U16634 (N_16634,N_16482,N_16469);
xnor U16635 (N_16635,N_16024,N_16010);
and U16636 (N_16636,N_16151,N_16111);
and U16637 (N_16637,N_16190,N_16495);
and U16638 (N_16638,N_16081,N_16158);
nor U16639 (N_16639,N_16349,N_16013);
nand U16640 (N_16640,N_16005,N_16445);
nand U16641 (N_16641,N_16027,N_16201);
nand U16642 (N_16642,N_16427,N_16209);
nand U16643 (N_16643,N_16304,N_16326);
and U16644 (N_16644,N_16235,N_16300);
or U16645 (N_16645,N_16234,N_16466);
or U16646 (N_16646,N_16451,N_16019);
nor U16647 (N_16647,N_16461,N_16174);
nor U16648 (N_16648,N_16168,N_16166);
nand U16649 (N_16649,N_16105,N_16334);
and U16650 (N_16650,N_16208,N_16149);
nor U16651 (N_16651,N_16261,N_16000);
nor U16652 (N_16652,N_16329,N_16084);
nor U16653 (N_16653,N_16004,N_16194);
xnor U16654 (N_16654,N_16150,N_16072);
xnor U16655 (N_16655,N_16455,N_16410);
and U16656 (N_16656,N_16474,N_16161);
or U16657 (N_16657,N_16390,N_16122);
nor U16658 (N_16658,N_16133,N_16045);
xnor U16659 (N_16659,N_16071,N_16274);
or U16660 (N_16660,N_16089,N_16262);
nand U16661 (N_16661,N_16096,N_16138);
nand U16662 (N_16662,N_16411,N_16374);
and U16663 (N_16663,N_16359,N_16159);
nand U16664 (N_16664,N_16497,N_16233);
or U16665 (N_16665,N_16036,N_16417);
or U16666 (N_16666,N_16295,N_16391);
nand U16667 (N_16667,N_16200,N_16382);
nor U16668 (N_16668,N_16252,N_16309);
or U16669 (N_16669,N_16470,N_16287);
nor U16670 (N_16670,N_16402,N_16254);
xnor U16671 (N_16671,N_16429,N_16239);
nand U16672 (N_16672,N_16332,N_16371);
nor U16673 (N_16673,N_16059,N_16145);
and U16674 (N_16674,N_16147,N_16217);
nor U16675 (N_16675,N_16131,N_16020);
nand U16676 (N_16676,N_16028,N_16026);
nor U16677 (N_16677,N_16407,N_16087);
xnor U16678 (N_16678,N_16132,N_16250);
or U16679 (N_16679,N_16197,N_16488);
and U16680 (N_16680,N_16058,N_16205);
nor U16681 (N_16681,N_16471,N_16075);
or U16682 (N_16682,N_16325,N_16401);
or U16683 (N_16683,N_16365,N_16346);
xnor U16684 (N_16684,N_16144,N_16413);
nor U16685 (N_16685,N_16007,N_16068);
nand U16686 (N_16686,N_16305,N_16393);
nand U16687 (N_16687,N_16259,N_16480);
or U16688 (N_16688,N_16043,N_16244);
nor U16689 (N_16689,N_16212,N_16405);
xnor U16690 (N_16690,N_16218,N_16289);
nor U16691 (N_16691,N_16403,N_16086);
nand U16692 (N_16692,N_16199,N_16387);
or U16693 (N_16693,N_16222,N_16226);
and U16694 (N_16694,N_16196,N_16016);
or U16695 (N_16695,N_16465,N_16082);
nor U16696 (N_16696,N_16454,N_16162);
nand U16697 (N_16697,N_16191,N_16269);
or U16698 (N_16698,N_16448,N_16054);
and U16699 (N_16699,N_16439,N_16092);
or U16700 (N_16700,N_16404,N_16018);
xor U16701 (N_16701,N_16220,N_16328);
and U16702 (N_16702,N_16011,N_16476);
and U16703 (N_16703,N_16117,N_16152);
nor U16704 (N_16704,N_16264,N_16319);
nand U16705 (N_16705,N_16492,N_16428);
or U16706 (N_16706,N_16042,N_16388);
or U16707 (N_16707,N_16116,N_16348);
and U16708 (N_16708,N_16415,N_16001);
nor U16709 (N_16709,N_16431,N_16038);
and U16710 (N_16710,N_16008,N_16475);
xor U16711 (N_16711,N_16291,N_16231);
nor U16712 (N_16712,N_16285,N_16459);
and U16713 (N_16713,N_16025,N_16221);
nand U16714 (N_16714,N_16186,N_16436);
xor U16715 (N_16715,N_16460,N_16437);
xor U16716 (N_16716,N_16121,N_16369);
nor U16717 (N_16717,N_16339,N_16342);
nand U16718 (N_16718,N_16039,N_16397);
nor U16719 (N_16719,N_16179,N_16477);
xnor U16720 (N_16720,N_16124,N_16423);
or U16721 (N_16721,N_16251,N_16327);
nand U16722 (N_16722,N_16364,N_16176);
nand U16723 (N_16723,N_16032,N_16373);
nor U16724 (N_16724,N_16472,N_16211);
nor U16725 (N_16725,N_16408,N_16100);
or U16726 (N_16726,N_16210,N_16175);
or U16727 (N_16727,N_16041,N_16112);
and U16728 (N_16728,N_16046,N_16203);
nor U16729 (N_16729,N_16260,N_16002);
nand U16730 (N_16730,N_16278,N_16379);
or U16731 (N_16731,N_16192,N_16294);
or U16732 (N_16732,N_16380,N_16406);
nand U16733 (N_16733,N_16306,N_16215);
nor U16734 (N_16734,N_16073,N_16247);
nor U16735 (N_16735,N_16356,N_16444);
and U16736 (N_16736,N_16271,N_16107);
nand U16737 (N_16737,N_16156,N_16034);
nand U16738 (N_16738,N_16337,N_16090);
nand U16739 (N_16739,N_16137,N_16130);
nand U16740 (N_16740,N_16298,N_16493);
nor U16741 (N_16741,N_16044,N_16430);
or U16742 (N_16742,N_16023,N_16307);
or U16743 (N_16743,N_16330,N_16076);
xor U16744 (N_16744,N_16499,N_16353);
or U16745 (N_16745,N_16485,N_16358);
or U16746 (N_16746,N_16433,N_16354);
xor U16747 (N_16747,N_16040,N_16172);
xor U16748 (N_16748,N_16314,N_16283);
nand U16749 (N_16749,N_16163,N_16022);
xor U16750 (N_16750,N_16396,N_16318);
nor U16751 (N_16751,N_16286,N_16400);
xor U16752 (N_16752,N_16259,N_16303);
or U16753 (N_16753,N_16091,N_16078);
and U16754 (N_16754,N_16192,N_16149);
or U16755 (N_16755,N_16111,N_16021);
nor U16756 (N_16756,N_16215,N_16268);
and U16757 (N_16757,N_16342,N_16149);
or U16758 (N_16758,N_16216,N_16354);
and U16759 (N_16759,N_16066,N_16048);
or U16760 (N_16760,N_16061,N_16290);
xnor U16761 (N_16761,N_16447,N_16115);
and U16762 (N_16762,N_16438,N_16097);
nand U16763 (N_16763,N_16412,N_16469);
nand U16764 (N_16764,N_16442,N_16024);
nand U16765 (N_16765,N_16312,N_16071);
or U16766 (N_16766,N_16228,N_16429);
xor U16767 (N_16767,N_16276,N_16496);
nand U16768 (N_16768,N_16366,N_16212);
nand U16769 (N_16769,N_16259,N_16324);
and U16770 (N_16770,N_16323,N_16186);
nor U16771 (N_16771,N_16373,N_16124);
nand U16772 (N_16772,N_16057,N_16238);
xor U16773 (N_16773,N_16480,N_16267);
xor U16774 (N_16774,N_16458,N_16453);
and U16775 (N_16775,N_16095,N_16019);
xor U16776 (N_16776,N_16470,N_16241);
xnor U16777 (N_16777,N_16446,N_16034);
nand U16778 (N_16778,N_16380,N_16256);
nor U16779 (N_16779,N_16125,N_16062);
nor U16780 (N_16780,N_16075,N_16110);
xnor U16781 (N_16781,N_16107,N_16496);
or U16782 (N_16782,N_16040,N_16086);
nor U16783 (N_16783,N_16248,N_16458);
xnor U16784 (N_16784,N_16178,N_16406);
nor U16785 (N_16785,N_16027,N_16078);
and U16786 (N_16786,N_16224,N_16121);
nor U16787 (N_16787,N_16424,N_16395);
and U16788 (N_16788,N_16404,N_16314);
or U16789 (N_16789,N_16351,N_16150);
nor U16790 (N_16790,N_16127,N_16179);
nor U16791 (N_16791,N_16372,N_16112);
or U16792 (N_16792,N_16396,N_16249);
xor U16793 (N_16793,N_16343,N_16458);
xnor U16794 (N_16794,N_16463,N_16441);
and U16795 (N_16795,N_16482,N_16304);
or U16796 (N_16796,N_16057,N_16162);
or U16797 (N_16797,N_16004,N_16463);
xnor U16798 (N_16798,N_16303,N_16091);
nor U16799 (N_16799,N_16210,N_16486);
xor U16800 (N_16800,N_16268,N_16192);
nor U16801 (N_16801,N_16416,N_16087);
xnor U16802 (N_16802,N_16013,N_16179);
nor U16803 (N_16803,N_16398,N_16255);
nor U16804 (N_16804,N_16114,N_16083);
and U16805 (N_16805,N_16248,N_16480);
or U16806 (N_16806,N_16031,N_16432);
nand U16807 (N_16807,N_16121,N_16356);
nor U16808 (N_16808,N_16148,N_16378);
or U16809 (N_16809,N_16030,N_16439);
and U16810 (N_16810,N_16123,N_16171);
nand U16811 (N_16811,N_16485,N_16284);
xor U16812 (N_16812,N_16151,N_16431);
nand U16813 (N_16813,N_16167,N_16110);
nor U16814 (N_16814,N_16429,N_16329);
nand U16815 (N_16815,N_16275,N_16395);
nand U16816 (N_16816,N_16423,N_16171);
xor U16817 (N_16817,N_16276,N_16084);
xor U16818 (N_16818,N_16055,N_16006);
or U16819 (N_16819,N_16427,N_16099);
and U16820 (N_16820,N_16414,N_16432);
nor U16821 (N_16821,N_16429,N_16224);
and U16822 (N_16822,N_16158,N_16465);
and U16823 (N_16823,N_16247,N_16259);
nand U16824 (N_16824,N_16399,N_16253);
xor U16825 (N_16825,N_16496,N_16089);
and U16826 (N_16826,N_16128,N_16358);
nand U16827 (N_16827,N_16041,N_16096);
nand U16828 (N_16828,N_16353,N_16308);
or U16829 (N_16829,N_16066,N_16130);
nor U16830 (N_16830,N_16238,N_16229);
or U16831 (N_16831,N_16385,N_16222);
nor U16832 (N_16832,N_16342,N_16233);
nand U16833 (N_16833,N_16388,N_16010);
nand U16834 (N_16834,N_16176,N_16450);
nand U16835 (N_16835,N_16014,N_16038);
or U16836 (N_16836,N_16291,N_16205);
nor U16837 (N_16837,N_16373,N_16036);
or U16838 (N_16838,N_16405,N_16443);
nor U16839 (N_16839,N_16085,N_16201);
and U16840 (N_16840,N_16382,N_16466);
and U16841 (N_16841,N_16042,N_16264);
nand U16842 (N_16842,N_16201,N_16291);
xor U16843 (N_16843,N_16131,N_16492);
nand U16844 (N_16844,N_16229,N_16236);
nor U16845 (N_16845,N_16179,N_16049);
nor U16846 (N_16846,N_16152,N_16362);
and U16847 (N_16847,N_16426,N_16383);
or U16848 (N_16848,N_16169,N_16315);
xor U16849 (N_16849,N_16474,N_16465);
xor U16850 (N_16850,N_16444,N_16068);
nand U16851 (N_16851,N_16372,N_16338);
or U16852 (N_16852,N_16058,N_16171);
and U16853 (N_16853,N_16076,N_16071);
nand U16854 (N_16854,N_16420,N_16217);
xor U16855 (N_16855,N_16190,N_16414);
nand U16856 (N_16856,N_16373,N_16268);
xor U16857 (N_16857,N_16325,N_16299);
or U16858 (N_16858,N_16429,N_16116);
and U16859 (N_16859,N_16110,N_16354);
nor U16860 (N_16860,N_16078,N_16311);
xnor U16861 (N_16861,N_16213,N_16402);
nand U16862 (N_16862,N_16056,N_16416);
nand U16863 (N_16863,N_16381,N_16092);
and U16864 (N_16864,N_16472,N_16203);
and U16865 (N_16865,N_16319,N_16402);
and U16866 (N_16866,N_16453,N_16030);
nor U16867 (N_16867,N_16228,N_16409);
xor U16868 (N_16868,N_16109,N_16182);
and U16869 (N_16869,N_16437,N_16200);
or U16870 (N_16870,N_16214,N_16191);
xor U16871 (N_16871,N_16210,N_16459);
or U16872 (N_16872,N_16264,N_16041);
and U16873 (N_16873,N_16412,N_16159);
nand U16874 (N_16874,N_16219,N_16393);
nor U16875 (N_16875,N_16112,N_16222);
nor U16876 (N_16876,N_16037,N_16393);
and U16877 (N_16877,N_16169,N_16360);
xnor U16878 (N_16878,N_16356,N_16200);
and U16879 (N_16879,N_16109,N_16491);
and U16880 (N_16880,N_16307,N_16177);
nor U16881 (N_16881,N_16476,N_16430);
and U16882 (N_16882,N_16452,N_16441);
xnor U16883 (N_16883,N_16206,N_16404);
nand U16884 (N_16884,N_16053,N_16059);
nor U16885 (N_16885,N_16447,N_16079);
nor U16886 (N_16886,N_16097,N_16154);
and U16887 (N_16887,N_16251,N_16352);
nand U16888 (N_16888,N_16318,N_16300);
nand U16889 (N_16889,N_16013,N_16404);
nor U16890 (N_16890,N_16475,N_16007);
nand U16891 (N_16891,N_16389,N_16005);
and U16892 (N_16892,N_16207,N_16058);
xor U16893 (N_16893,N_16485,N_16259);
nand U16894 (N_16894,N_16257,N_16107);
nor U16895 (N_16895,N_16146,N_16128);
or U16896 (N_16896,N_16020,N_16167);
xnor U16897 (N_16897,N_16488,N_16034);
xnor U16898 (N_16898,N_16015,N_16291);
nor U16899 (N_16899,N_16452,N_16330);
nand U16900 (N_16900,N_16354,N_16183);
nand U16901 (N_16901,N_16190,N_16469);
or U16902 (N_16902,N_16210,N_16296);
or U16903 (N_16903,N_16495,N_16173);
or U16904 (N_16904,N_16250,N_16016);
or U16905 (N_16905,N_16472,N_16206);
or U16906 (N_16906,N_16139,N_16337);
nor U16907 (N_16907,N_16499,N_16129);
and U16908 (N_16908,N_16305,N_16094);
nand U16909 (N_16909,N_16230,N_16235);
nor U16910 (N_16910,N_16360,N_16349);
nor U16911 (N_16911,N_16445,N_16407);
nor U16912 (N_16912,N_16464,N_16270);
or U16913 (N_16913,N_16401,N_16457);
nand U16914 (N_16914,N_16070,N_16156);
and U16915 (N_16915,N_16100,N_16119);
xnor U16916 (N_16916,N_16458,N_16238);
nor U16917 (N_16917,N_16247,N_16455);
and U16918 (N_16918,N_16084,N_16497);
nor U16919 (N_16919,N_16371,N_16080);
and U16920 (N_16920,N_16473,N_16482);
xor U16921 (N_16921,N_16142,N_16106);
xnor U16922 (N_16922,N_16334,N_16252);
nor U16923 (N_16923,N_16044,N_16366);
or U16924 (N_16924,N_16171,N_16151);
nand U16925 (N_16925,N_16100,N_16351);
or U16926 (N_16926,N_16293,N_16446);
nand U16927 (N_16927,N_16458,N_16317);
or U16928 (N_16928,N_16405,N_16229);
and U16929 (N_16929,N_16122,N_16437);
nand U16930 (N_16930,N_16061,N_16082);
nand U16931 (N_16931,N_16334,N_16047);
or U16932 (N_16932,N_16320,N_16135);
xnor U16933 (N_16933,N_16205,N_16351);
xnor U16934 (N_16934,N_16168,N_16283);
xor U16935 (N_16935,N_16196,N_16235);
nor U16936 (N_16936,N_16071,N_16353);
and U16937 (N_16937,N_16209,N_16101);
nor U16938 (N_16938,N_16064,N_16104);
and U16939 (N_16939,N_16406,N_16404);
xnor U16940 (N_16940,N_16302,N_16088);
nand U16941 (N_16941,N_16268,N_16309);
nor U16942 (N_16942,N_16262,N_16415);
xor U16943 (N_16943,N_16301,N_16202);
nand U16944 (N_16944,N_16188,N_16256);
xnor U16945 (N_16945,N_16059,N_16311);
or U16946 (N_16946,N_16150,N_16091);
xor U16947 (N_16947,N_16386,N_16444);
and U16948 (N_16948,N_16395,N_16322);
or U16949 (N_16949,N_16386,N_16484);
nor U16950 (N_16950,N_16059,N_16491);
nor U16951 (N_16951,N_16348,N_16424);
nor U16952 (N_16952,N_16307,N_16497);
and U16953 (N_16953,N_16453,N_16064);
nand U16954 (N_16954,N_16280,N_16209);
nand U16955 (N_16955,N_16063,N_16036);
nor U16956 (N_16956,N_16151,N_16443);
xnor U16957 (N_16957,N_16275,N_16342);
nand U16958 (N_16958,N_16285,N_16289);
or U16959 (N_16959,N_16377,N_16047);
xor U16960 (N_16960,N_16468,N_16280);
nor U16961 (N_16961,N_16494,N_16445);
nor U16962 (N_16962,N_16283,N_16297);
nor U16963 (N_16963,N_16214,N_16144);
xor U16964 (N_16964,N_16467,N_16060);
and U16965 (N_16965,N_16220,N_16293);
xor U16966 (N_16966,N_16286,N_16361);
xnor U16967 (N_16967,N_16271,N_16288);
nor U16968 (N_16968,N_16062,N_16399);
and U16969 (N_16969,N_16212,N_16470);
and U16970 (N_16970,N_16169,N_16207);
xor U16971 (N_16971,N_16220,N_16298);
xnor U16972 (N_16972,N_16229,N_16437);
nor U16973 (N_16973,N_16082,N_16388);
nor U16974 (N_16974,N_16214,N_16138);
or U16975 (N_16975,N_16202,N_16412);
or U16976 (N_16976,N_16047,N_16027);
xnor U16977 (N_16977,N_16036,N_16401);
nand U16978 (N_16978,N_16003,N_16300);
nand U16979 (N_16979,N_16403,N_16483);
nor U16980 (N_16980,N_16491,N_16395);
or U16981 (N_16981,N_16314,N_16458);
nor U16982 (N_16982,N_16291,N_16079);
and U16983 (N_16983,N_16199,N_16347);
or U16984 (N_16984,N_16115,N_16225);
or U16985 (N_16985,N_16492,N_16027);
xor U16986 (N_16986,N_16047,N_16447);
nor U16987 (N_16987,N_16189,N_16022);
nand U16988 (N_16988,N_16130,N_16222);
nand U16989 (N_16989,N_16216,N_16394);
nor U16990 (N_16990,N_16248,N_16003);
xnor U16991 (N_16991,N_16146,N_16293);
or U16992 (N_16992,N_16044,N_16133);
nor U16993 (N_16993,N_16313,N_16462);
and U16994 (N_16994,N_16362,N_16012);
xor U16995 (N_16995,N_16305,N_16411);
nand U16996 (N_16996,N_16007,N_16140);
nor U16997 (N_16997,N_16292,N_16006);
xor U16998 (N_16998,N_16062,N_16396);
nor U16999 (N_16999,N_16258,N_16425);
nor U17000 (N_17000,N_16581,N_16503);
xnor U17001 (N_17001,N_16754,N_16557);
xnor U17002 (N_17002,N_16975,N_16751);
nand U17003 (N_17003,N_16521,N_16767);
nand U17004 (N_17004,N_16505,N_16747);
nand U17005 (N_17005,N_16864,N_16980);
nor U17006 (N_17006,N_16946,N_16591);
or U17007 (N_17007,N_16504,N_16652);
nor U17008 (N_17008,N_16892,N_16685);
nand U17009 (N_17009,N_16550,N_16909);
or U17010 (N_17010,N_16809,N_16618);
nand U17011 (N_17011,N_16533,N_16737);
xor U17012 (N_17012,N_16871,N_16776);
xnor U17013 (N_17013,N_16831,N_16880);
or U17014 (N_17014,N_16819,N_16610);
and U17015 (N_17015,N_16915,N_16796);
or U17016 (N_17016,N_16606,N_16905);
nor U17017 (N_17017,N_16537,N_16609);
nor U17018 (N_17018,N_16710,N_16781);
and U17019 (N_17019,N_16692,N_16735);
and U17020 (N_17020,N_16518,N_16567);
nand U17021 (N_17021,N_16563,N_16999);
nand U17022 (N_17022,N_16811,N_16956);
and U17023 (N_17023,N_16532,N_16862);
nand U17024 (N_17024,N_16935,N_16608);
and U17025 (N_17025,N_16649,N_16719);
nor U17026 (N_17026,N_16939,N_16502);
nand U17027 (N_17027,N_16839,N_16788);
nand U17028 (N_17028,N_16854,N_16808);
and U17029 (N_17029,N_16714,N_16799);
nand U17030 (N_17030,N_16955,N_16711);
and U17031 (N_17031,N_16965,N_16583);
xor U17032 (N_17032,N_16589,N_16912);
nor U17033 (N_17033,N_16893,N_16682);
xor U17034 (N_17034,N_16662,N_16549);
and U17035 (N_17035,N_16742,N_16868);
nor U17036 (N_17036,N_16522,N_16593);
and U17037 (N_17037,N_16827,N_16923);
xnor U17038 (N_17038,N_16793,N_16655);
nor U17039 (N_17039,N_16640,N_16953);
nand U17040 (N_17040,N_16829,N_16744);
nand U17041 (N_17041,N_16680,N_16562);
nand U17042 (N_17042,N_16646,N_16607);
nor U17043 (N_17043,N_16543,N_16579);
nand U17044 (N_17044,N_16968,N_16990);
nand U17045 (N_17045,N_16508,N_16906);
and U17046 (N_17046,N_16875,N_16643);
nor U17047 (N_17047,N_16706,N_16555);
and U17048 (N_17048,N_16930,N_16852);
nor U17049 (N_17049,N_16560,N_16654);
or U17050 (N_17050,N_16826,N_16604);
nand U17051 (N_17051,N_16559,N_16985);
nand U17052 (N_17052,N_16869,N_16536);
nor U17053 (N_17053,N_16668,N_16840);
nor U17054 (N_17054,N_16770,N_16592);
or U17055 (N_17055,N_16671,N_16667);
nor U17056 (N_17056,N_16895,N_16613);
or U17057 (N_17057,N_16628,N_16763);
xor U17058 (N_17058,N_16701,N_16988);
or U17059 (N_17059,N_16899,N_16860);
and U17060 (N_17060,N_16683,N_16526);
nor U17061 (N_17061,N_16994,N_16630);
nor U17062 (N_17062,N_16568,N_16524);
xor U17063 (N_17063,N_16542,N_16716);
or U17064 (N_17064,N_16547,N_16556);
nor U17065 (N_17065,N_16972,N_16723);
xnor U17066 (N_17066,N_16700,N_16582);
and U17067 (N_17067,N_16566,N_16684);
or U17068 (N_17068,N_16870,N_16539);
nor U17069 (N_17069,N_16952,N_16725);
and U17070 (N_17070,N_16883,N_16746);
and U17071 (N_17071,N_16535,N_16509);
xor U17072 (N_17072,N_16861,N_16850);
or U17073 (N_17073,N_16983,N_16689);
nand U17074 (N_17074,N_16670,N_16941);
nand U17075 (N_17075,N_16734,N_16901);
nand U17076 (N_17076,N_16832,N_16573);
xnor U17077 (N_17077,N_16847,N_16812);
and U17078 (N_17078,N_16639,N_16707);
xnor U17079 (N_17079,N_16715,N_16515);
nand U17080 (N_17080,N_16674,N_16998);
xor U17081 (N_17081,N_16529,N_16511);
and U17082 (N_17082,N_16506,N_16704);
or U17083 (N_17083,N_16718,N_16645);
xnor U17084 (N_17084,N_16791,N_16756);
or U17085 (N_17085,N_16678,N_16825);
xor U17086 (N_17086,N_16748,N_16631);
xnor U17087 (N_17087,N_16545,N_16903);
and U17088 (N_17088,N_16884,N_16777);
nand U17089 (N_17089,N_16815,N_16814);
and U17090 (N_17090,N_16614,N_16943);
xor U17091 (N_17091,N_16789,N_16888);
and U17092 (N_17092,N_16865,N_16836);
nor U17093 (N_17093,N_16922,N_16576);
nor U17094 (N_17094,N_16838,N_16779);
and U17095 (N_17095,N_16920,N_16585);
nor U17096 (N_17096,N_16695,N_16616);
and U17097 (N_17097,N_16802,N_16992);
xor U17098 (N_17098,N_16797,N_16774);
xnor U17099 (N_17099,N_16690,N_16786);
nor U17100 (N_17100,N_16970,N_16558);
or U17101 (N_17101,N_16936,N_16771);
or U17102 (N_17102,N_16958,N_16790);
nor U17103 (N_17103,N_16580,N_16876);
xor U17104 (N_17104,N_16782,N_16553);
xnor U17105 (N_17105,N_16733,N_16743);
and U17106 (N_17106,N_16961,N_16863);
and U17107 (N_17107,N_16507,N_16708);
xor U17108 (N_17108,N_16621,N_16816);
nand U17109 (N_17109,N_16996,N_16633);
nand U17110 (N_17110,N_16561,N_16926);
nand U17111 (N_17111,N_16612,N_16800);
nand U17112 (N_17112,N_16709,N_16913);
xor U17113 (N_17113,N_16638,N_16969);
or U17114 (N_17114,N_16773,N_16931);
and U17115 (N_17115,N_16750,N_16534);
nand U17116 (N_17116,N_16967,N_16887);
xor U17117 (N_17117,N_16531,N_16702);
nor U17118 (N_17118,N_16823,N_16552);
and U17119 (N_17119,N_16745,N_16927);
nand U17120 (N_17120,N_16530,N_16554);
nand U17121 (N_17121,N_16886,N_16605);
or U17122 (N_17122,N_16548,N_16921);
and U17123 (N_17123,N_16760,N_16803);
nand U17124 (N_17124,N_16962,N_16993);
and U17125 (N_17125,N_16938,N_16986);
xnor U17126 (N_17126,N_16694,N_16792);
xnor U17127 (N_17127,N_16660,N_16721);
nor U17128 (N_17128,N_16785,N_16635);
nand U17129 (N_17129,N_16977,N_16590);
or U17130 (N_17130,N_16642,N_16873);
and U17131 (N_17131,N_16594,N_16724);
nand U17132 (N_17132,N_16712,N_16765);
and U17133 (N_17133,N_16769,N_16757);
xor U17134 (N_17134,N_16699,N_16948);
nand U17135 (N_17135,N_16540,N_16749);
nand U17136 (N_17136,N_16720,N_16705);
or U17137 (N_17137,N_16966,N_16738);
or U17138 (N_17138,N_16947,N_16626);
xor U17139 (N_17139,N_16902,N_16984);
xnor U17140 (N_17140,N_16571,N_16885);
nor U17141 (N_17141,N_16805,N_16665);
nor U17142 (N_17142,N_16625,N_16527);
nand U17143 (N_17143,N_16960,N_16634);
nand U17144 (N_17144,N_16577,N_16783);
nand U17145 (N_17145,N_16991,N_16917);
or U17146 (N_17146,N_16647,N_16525);
or U17147 (N_17147,N_16663,N_16950);
nor U17148 (N_17148,N_16882,N_16795);
or U17149 (N_17149,N_16780,N_16603);
or U17150 (N_17150,N_16857,N_16835);
or U17151 (N_17151,N_16807,N_16601);
and U17152 (N_17152,N_16517,N_16928);
nand U17153 (N_17153,N_16866,N_16964);
nand U17154 (N_17154,N_16820,N_16904);
and U17155 (N_17155,N_16676,N_16973);
and U17156 (N_17156,N_16672,N_16907);
and U17157 (N_17157,N_16673,N_16954);
and U17158 (N_17158,N_16622,N_16794);
and U17159 (N_17159,N_16801,N_16908);
and U17160 (N_17160,N_16806,N_16600);
xor U17161 (N_17161,N_16989,N_16787);
and U17162 (N_17162,N_16810,N_16910);
and U17163 (N_17163,N_16637,N_16636);
nor U17164 (N_17164,N_16874,N_16500);
xnor U17165 (N_17165,N_16698,N_16858);
or U17166 (N_17166,N_16848,N_16981);
nand U17167 (N_17167,N_16932,N_16942);
and U17168 (N_17168,N_16741,N_16804);
or U17169 (N_17169,N_16584,N_16818);
or U17170 (N_17170,N_16987,N_16872);
and U17171 (N_17171,N_16546,N_16541);
xor U17172 (N_17172,N_16653,N_16828);
nor U17173 (N_17173,N_16681,N_16978);
xor U17174 (N_17174,N_16564,N_16528);
and U17175 (N_17175,N_16813,N_16615);
nand U17176 (N_17176,N_16619,N_16891);
nand U17177 (N_17177,N_16916,N_16971);
or U17178 (N_17178,N_16824,N_16523);
nand U17179 (N_17179,N_16696,N_16659);
and U17180 (N_17180,N_16516,N_16859);
xnor U17181 (N_17181,N_16597,N_16775);
and U17182 (N_17182,N_16669,N_16798);
xor U17183 (N_17183,N_16664,N_16768);
and U17184 (N_17184,N_16879,N_16934);
nand U17185 (N_17185,N_16572,N_16599);
or U17186 (N_17186,N_16817,N_16570);
or U17187 (N_17187,N_16675,N_16940);
nand U17188 (N_17188,N_16551,N_16846);
nand U17189 (N_17189,N_16717,N_16762);
xnor U17190 (N_17190,N_16679,N_16588);
nor U17191 (N_17191,N_16849,N_16951);
xor U17192 (N_17192,N_16666,N_16844);
or U17193 (N_17193,N_16519,N_16687);
and U17194 (N_17194,N_16924,N_16833);
nor U17195 (N_17195,N_16501,N_16620);
xnor U17196 (N_17196,N_16753,N_16761);
and U17197 (N_17197,N_16764,N_16656);
or U17198 (N_17198,N_16834,N_16778);
xor U17199 (N_17199,N_16569,N_16595);
or U17200 (N_17200,N_16851,N_16586);
xor U17201 (N_17201,N_16755,N_16730);
or U17202 (N_17202,N_16611,N_16841);
nand U17203 (N_17203,N_16945,N_16898);
and U17204 (N_17204,N_16784,N_16726);
nor U17205 (N_17205,N_16867,N_16658);
nand U17206 (N_17206,N_16878,N_16837);
xor U17207 (N_17207,N_16772,N_16575);
xor U17208 (N_17208,N_16544,N_16644);
or U17209 (N_17209,N_16732,N_16739);
or U17210 (N_17210,N_16914,N_16979);
xnor U17211 (N_17211,N_16661,N_16513);
nand U17212 (N_17212,N_16623,N_16959);
and U17213 (N_17213,N_16758,N_16703);
and U17214 (N_17214,N_16937,N_16565);
xor U17215 (N_17215,N_16911,N_16520);
xor U17216 (N_17216,N_16731,N_16890);
nand U17217 (N_17217,N_16729,N_16881);
xor U17218 (N_17218,N_16512,N_16693);
nor U17219 (N_17219,N_16997,N_16995);
nand U17220 (N_17220,N_16657,N_16752);
xnor U17221 (N_17221,N_16845,N_16957);
or U17222 (N_17222,N_16822,N_16821);
and U17223 (N_17223,N_16722,N_16736);
nand U17224 (N_17224,N_16624,N_16919);
or U17225 (N_17225,N_16918,N_16842);
and U17226 (N_17226,N_16587,N_16598);
xnor U17227 (N_17227,N_16686,N_16974);
nand U17228 (N_17228,N_16728,N_16830);
or U17229 (N_17229,N_16538,N_16944);
nand U17230 (N_17230,N_16677,N_16650);
and U17231 (N_17231,N_16713,N_16697);
nor U17232 (N_17232,N_16976,N_16925);
xnor U17233 (N_17233,N_16632,N_16510);
or U17234 (N_17234,N_16629,N_16617);
nor U17235 (N_17235,N_16949,N_16963);
and U17236 (N_17236,N_16897,N_16933);
nor U17237 (N_17237,N_16877,N_16574);
xnor U17238 (N_17238,N_16843,N_16740);
nor U17239 (N_17239,N_16514,N_16894);
or U17240 (N_17240,N_16759,N_16727);
and U17241 (N_17241,N_16766,N_16627);
nand U17242 (N_17242,N_16651,N_16889);
xnor U17243 (N_17243,N_16982,N_16648);
or U17244 (N_17244,N_16578,N_16691);
or U17245 (N_17245,N_16900,N_16641);
nor U17246 (N_17246,N_16929,N_16596);
nor U17247 (N_17247,N_16853,N_16688);
xor U17248 (N_17248,N_16855,N_16856);
xor U17249 (N_17249,N_16602,N_16896);
nor U17250 (N_17250,N_16841,N_16827);
xor U17251 (N_17251,N_16583,N_16719);
and U17252 (N_17252,N_16744,N_16541);
xnor U17253 (N_17253,N_16649,N_16680);
xnor U17254 (N_17254,N_16999,N_16936);
nor U17255 (N_17255,N_16766,N_16909);
or U17256 (N_17256,N_16995,N_16641);
nor U17257 (N_17257,N_16519,N_16596);
and U17258 (N_17258,N_16830,N_16754);
or U17259 (N_17259,N_16798,N_16688);
nand U17260 (N_17260,N_16728,N_16640);
xor U17261 (N_17261,N_16526,N_16594);
nand U17262 (N_17262,N_16979,N_16849);
or U17263 (N_17263,N_16757,N_16610);
xnor U17264 (N_17264,N_16697,N_16591);
xnor U17265 (N_17265,N_16971,N_16871);
or U17266 (N_17266,N_16585,N_16721);
nor U17267 (N_17267,N_16723,N_16963);
nand U17268 (N_17268,N_16842,N_16833);
xnor U17269 (N_17269,N_16966,N_16856);
or U17270 (N_17270,N_16504,N_16900);
nor U17271 (N_17271,N_16906,N_16888);
and U17272 (N_17272,N_16672,N_16505);
nor U17273 (N_17273,N_16512,N_16672);
xnor U17274 (N_17274,N_16749,N_16719);
nor U17275 (N_17275,N_16967,N_16818);
or U17276 (N_17276,N_16879,N_16831);
or U17277 (N_17277,N_16667,N_16568);
nand U17278 (N_17278,N_16564,N_16764);
nor U17279 (N_17279,N_16658,N_16936);
nand U17280 (N_17280,N_16920,N_16998);
or U17281 (N_17281,N_16902,N_16512);
nand U17282 (N_17282,N_16913,N_16926);
nor U17283 (N_17283,N_16928,N_16726);
nand U17284 (N_17284,N_16918,N_16539);
and U17285 (N_17285,N_16625,N_16537);
xnor U17286 (N_17286,N_16690,N_16953);
or U17287 (N_17287,N_16673,N_16992);
and U17288 (N_17288,N_16503,N_16688);
xnor U17289 (N_17289,N_16827,N_16901);
nand U17290 (N_17290,N_16847,N_16500);
or U17291 (N_17291,N_16662,N_16737);
nor U17292 (N_17292,N_16910,N_16921);
nand U17293 (N_17293,N_16730,N_16656);
xor U17294 (N_17294,N_16787,N_16944);
nor U17295 (N_17295,N_16751,N_16573);
nand U17296 (N_17296,N_16981,N_16763);
xnor U17297 (N_17297,N_16721,N_16703);
xnor U17298 (N_17298,N_16973,N_16540);
nor U17299 (N_17299,N_16509,N_16614);
or U17300 (N_17300,N_16836,N_16551);
nand U17301 (N_17301,N_16537,N_16614);
or U17302 (N_17302,N_16568,N_16936);
or U17303 (N_17303,N_16577,N_16823);
xor U17304 (N_17304,N_16828,N_16623);
xor U17305 (N_17305,N_16556,N_16704);
nor U17306 (N_17306,N_16967,N_16820);
nand U17307 (N_17307,N_16978,N_16875);
and U17308 (N_17308,N_16614,N_16998);
or U17309 (N_17309,N_16724,N_16849);
and U17310 (N_17310,N_16510,N_16974);
nor U17311 (N_17311,N_16740,N_16958);
and U17312 (N_17312,N_16671,N_16799);
nand U17313 (N_17313,N_16688,N_16818);
or U17314 (N_17314,N_16981,N_16682);
and U17315 (N_17315,N_16555,N_16737);
xor U17316 (N_17316,N_16559,N_16910);
nand U17317 (N_17317,N_16764,N_16953);
and U17318 (N_17318,N_16814,N_16950);
xnor U17319 (N_17319,N_16902,N_16788);
nor U17320 (N_17320,N_16695,N_16987);
nand U17321 (N_17321,N_16834,N_16975);
and U17322 (N_17322,N_16640,N_16539);
nor U17323 (N_17323,N_16841,N_16967);
nand U17324 (N_17324,N_16637,N_16803);
nor U17325 (N_17325,N_16814,N_16683);
nand U17326 (N_17326,N_16656,N_16755);
nor U17327 (N_17327,N_16712,N_16866);
xnor U17328 (N_17328,N_16508,N_16595);
nand U17329 (N_17329,N_16767,N_16968);
and U17330 (N_17330,N_16599,N_16855);
nand U17331 (N_17331,N_16638,N_16985);
nand U17332 (N_17332,N_16722,N_16513);
nor U17333 (N_17333,N_16984,N_16627);
xnor U17334 (N_17334,N_16608,N_16827);
and U17335 (N_17335,N_16567,N_16790);
xnor U17336 (N_17336,N_16716,N_16549);
or U17337 (N_17337,N_16622,N_16699);
xor U17338 (N_17338,N_16610,N_16865);
xor U17339 (N_17339,N_16829,N_16701);
and U17340 (N_17340,N_16979,N_16981);
nor U17341 (N_17341,N_16795,N_16927);
or U17342 (N_17342,N_16857,N_16986);
nor U17343 (N_17343,N_16797,N_16585);
nor U17344 (N_17344,N_16814,N_16824);
nand U17345 (N_17345,N_16888,N_16647);
xor U17346 (N_17346,N_16512,N_16664);
xnor U17347 (N_17347,N_16788,N_16773);
nor U17348 (N_17348,N_16902,N_16802);
xnor U17349 (N_17349,N_16590,N_16814);
and U17350 (N_17350,N_16544,N_16719);
nand U17351 (N_17351,N_16546,N_16563);
xor U17352 (N_17352,N_16834,N_16888);
nand U17353 (N_17353,N_16930,N_16742);
nor U17354 (N_17354,N_16873,N_16815);
and U17355 (N_17355,N_16820,N_16564);
xor U17356 (N_17356,N_16761,N_16631);
nand U17357 (N_17357,N_16853,N_16517);
and U17358 (N_17358,N_16506,N_16773);
nand U17359 (N_17359,N_16543,N_16980);
and U17360 (N_17360,N_16639,N_16696);
nor U17361 (N_17361,N_16659,N_16753);
or U17362 (N_17362,N_16664,N_16913);
or U17363 (N_17363,N_16542,N_16603);
or U17364 (N_17364,N_16951,N_16946);
xnor U17365 (N_17365,N_16868,N_16605);
nor U17366 (N_17366,N_16669,N_16828);
nand U17367 (N_17367,N_16617,N_16599);
nand U17368 (N_17368,N_16732,N_16798);
nand U17369 (N_17369,N_16775,N_16570);
and U17370 (N_17370,N_16978,N_16884);
or U17371 (N_17371,N_16674,N_16744);
nor U17372 (N_17372,N_16658,N_16868);
nor U17373 (N_17373,N_16990,N_16907);
xnor U17374 (N_17374,N_16858,N_16752);
xor U17375 (N_17375,N_16839,N_16924);
xnor U17376 (N_17376,N_16635,N_16885);
and U17377 (N_17377,N_16885,N_16702);
and U17378 (N_17378,N_16836,N_16882);
nor U17379 (N_17379,N_16833,N_16912);
nand U17380 (N_17380,N_16676,N_16882);
nor U17381 (N_17381,N_16803,N_16991);
or U17382 (N_17382,N_16945,N_16786);
or U17383 (N_17383,N_16824,N_16599);
nand U17384 (N_17384,N_16641,N_16529);
xor U17385 (N_17385,N_16856,N_16892);
xor U17386 (N_17386,N_16709,N_16893);
and U17387 (N_17387,N_16712,N_16733);
nor U17388 (N_17388,N_16793,N_16769);
or U17389 (N_17389,N_16892,N_16995);
xor U17390 (N_17390,N_16550,N_16645);
and U17391 (N_17391,N_16635,N_16719);
xnor U17392 (N_17392,N_16598,N_16806);
xor U17393 (N_17393,N_16708,N_16802);
nand U17394 (N_17394,N_16913,N_16943);
nor U17395 (N_17395,N_16632,N_16514);
xor U17396 (N_17396,N_16712,N_16936);
and U17397 (N_17397,N_16779,N_16649);
or U17398 (N_17398,N_16731,N_16559);
xnor U17399 (N_17399,N_16772,N_16905);
xor U17400 (N_17400,N_16860,N_16777);
or U17401 (N_17401,N_16604,N_16846);
nand U17402 (N_17402,N_16897,N_16873);
nand U17403 (N_17403,N_16919,N_16851);
or U17404 (N_17404,N_16898,N_16993);
and U17405 (N_17405,N_16673,N_16996);
and U17406 (N_17406,N_16699,N_16849);
nor U17407 (N_17407,N_16763,N_16607);
xnor U17408 (N_17408,N_16548,N_16500);
and U17409 (N_17409,N_16575,N_16694);
nor U17410 (N_17410,N_16661,N_16917);
or U17411 (N_17411,N_16706,N_16592);
and U17412 (N_17412,N_16545,N_16678);
xor U17413 (N_17413,N_16736,N_16655);
or U17414 (N_17414,N_16590,N_16827);
nor U17415 (N_17415,N_16705,N_16556);
xor U17416 (N_17416,N_16893,N_16613);
and U17417 (N_17417,N_16823,N_16938);
or U17418 (N_17418,N_16716,N_16702);
or U17419 (N_17419,N_16613,N_16962);
or U17420 (N_17420,N_16587,N_16676);
or U17421 (N_17421,N_16500,N_16666);
nand U17422 (N_17422,N_16671,N_16976);
xnor U17423 (N_17423,N_16553,N_16941);
or U17424 (N_17424,N_16944,N_16814);
and U17425 (N_17425,N_16702,N_16654);
xor U17426 (N_17426,N_16731,N_16693);
or U17427 (N_17427,N_16849,N_16962);
xnor U17428 (N_17428,N_16951,N_16916);
nand U17429 (N_17429,N_16679,N_16716);
and U17430 (N_17430,N_16944,N_16522);
and U17431 (N_17431,N_16691,N_16753);
xor U17432 (N_17432,N_16882,N_16883);
or U17433 (N_17433,N_16866,N_16583);
nor U17434 (N_17434,N_16967,N_16570);
and U17435 (N_17435,N_16838,N_16568);
and U17436 (N_17436,N_16813,N_16948);
nor U17437 (N_17437,N_16820,N_16531);
nand U17438 (N_17438,N_16696,N_16760);
nor U17439 (N_17439,N_16772,N_16824);
nand U17440 (N_17440,N_16849,N_16516);
nand U17441 (N_17441,N_16684,N_16851);
nor U17442 (N_17442,N_16614,N_16939);
xor U17443 (N_17443,N_16677,N_16980);
nand U17444 (N_17444,N_16960,N_16753);
and U17445 (N_17445,N_16801,N_16720);
or U17446 (N_17446,N_16784,N_16791);
nor U17447 (N_17447,N_16968,N_16701);
or U17448 (N_17448,N_16573,N_16814);
nor U17449 (N_17449,N_16777,N_16539);
nor U17450 (N_17450,N_16511,N_16919);
nand U17451 (N_17451,N_16619,N_16883);
nand U17452 (N_17452,N_16819,N_16614);
xnor U17453 (N_17453,N_16856,N_16726);
nor U17454 (N_17454,N_16604,N_16676);
nor U17455 (N_17455,N_16783,N_16806);
nor U17456 (N_17456,N_16507,N_16689);
nor U17457 (N_17457,N_16832,N_16772);
nor U17458 (N_17458,N_16594,N_16711);
nand U17459 (N_17459,N_16551,N_16852);
nor U17460 (N_17460,N_16809,N_16578);
xor U17461 (N_17461,N_16798,N_16921);
nand U17462 (N_17462,N_16973,N_16733);
or U17463 (N_17463,N_16949,N_16522);
nor U17464 (N_17464,N_16732,N_16560);
xor U17465 (N_17465,N_16691,N_16582);
nand U17466 (N_17466,N_16598,N_16654);
nand U17467 (N_17467,N_16638,N_16971);
nand U17468 (N_17468,N_16712,N_16518);
nor U17469 (N_17469,N_16930,N_16758);
nand U17470 (N_17470,N_16707,N_16718);
xnor U17471 (N_17471,N_16956,N_16641);
nand U17472 (N_17472,N_16805,N_16704);
nand U17473 (N_17473,N_16834,N_16881);
or U17474 (N_17474,N_16667,N_16526);
or U17475 (N_17475,N_16763,N_16814);
nor U17476 (N_17476,N_16625,N_16991);
or U17477 (N_17477,N_16869,N_16708);
and U17478 (N_17478,N_16766,N_16739);
or U17479 (N_17479,N_16500,N_16530);
and U17480 (N_17480,N_16998,N_16636);
xnor U17481 (N_17481,N_16963,N_16836);
nor U17482 (N_17482,N_16628,N_16856);
xnor U17483 (N_17483,N_16957,N_16798);
or U17484 (N_17484,N_16890,N_16633);
nor U17485 (N_17485,N_16642,N_16813);
and U17486 (N_17486,N_16896,N_16626);
xnor U17487 (N_17487,N_16993,N_16754);
and U17488 (N_17488,N_16669,N_16676);
nor U17489 (N_17489,N_16632,N_16735);
nand U17490 (N_17490,N_16830,N_16709);
nand U17491 (N_17491,N_16742,N_16990);
nor U17492 (N_17492,N_16547,N_16951);
nor U17493 (N_17493,N_16934,N_16800);
nand U17494 (N_17494,N_16623,N_16803);
nor U17495 (N_17495,N_16961,N_16870);
or U17496 (N_17496,N_16787,N_16535);
or U17497 (N_17497,N_16988,N_16758);
nor U17498 (N_17498,N_16987,N_16990);
nand U17499 (N_17499,N_16980,N_16670);
xor U17500 (N_17500,N_17381,N_17388);
xnor U17501 (N_17501,N_17297,N_17422);
xor U17502 (N_17502,N_17368,N_17064);
and U17503 (N_17503,N_17233,N_17162);
xor U17504 (N_17504,N_17014,N_17081);
or U17505 (N_17505,N_17439,N_17328);
and U17506 (N_17506,N_17481,N_17232);
nor U17507 (N_17507,N_17462,N_17456);
or U17508 (N_17508,N_17478,N_17370);
and U17509 (N_17509,N_17337,N_17257);
nand U17510 (N_17510,N_17311,N_17461);
and U17511 (N_17511,N_17256,N_17354);
or U17512 (N_17512,N_17334,N_17121);
or U17513 (N_17513,N_17196,N_17054);
or U17514 (N_17514,N_17405,N_17383);
or U17515 (N_17515,N_17124,N_17067);
nor U17516 (N_17516,N_17276,N_17105);
xnor U17517 (N_17517,N_17473,N_17321);
xor U17518 (N_17518,N_17069,N_17062);
or U17519 (N_17519,N_17187,N_17415);
or U17520 (N_17520,N_17469,N_17406);
nor U17521 (N_17521,N_17397,N_17443);
nor U17522 (N_17522,N_17491,N_17013);
nor U17523 (N_17523,N_17213,N_17129);
and U17524 (N_17524,N_17326,N_17211);
or U17525 (N_17525,N_17202,N_17155);
or U17526 (N_17526,N_17270,N_17079);
xor U17527 (N_17527,N_17269,N_17194);
nand U17528 (N_17528,N_17059,N_17109);
and U17529 (N_17529,N_17010,N_17208);
nand U17530 (N_17530,N_17045,N_17240);
or U17531 (N_17531,N_17253,N_17179);
nand U17532 (N_17532,N_17477,N_17131);
nand U17533 (N_17533,N_17167,N_17459);
and U17534 (N_17534,N_17214,N_17363);
nand U17535 (N_17535,N_17025,N_17031);
nand U17536 (N_17536,N_17409,N_17258);
and U17537 (N_17537,N_17386,N_17078);
and U17538 (N_17538,N_17329,N_17317);
and U17539 (N_17539,N_17086,N_17437);
or U17540 (N_17540,N_17490,N_17482);
or U17541 (N_17541,N_17138,N_17222);
xnor U17542 (N_17542,N_17177,N_17040);
or U17543 (N_17543,N_17352,N_17003);
nor U17544 (N_17544,N_17396,N_17418);
and U17545 (N_17545,N_17082,N_17038);
and U17546 (N_17546,N_17362,N_17034);
nor U17547 (N_17547,N_17466,N_17331);
xnor U17548 (N_17548,N_17008,N_17313);
and U17549 (N_17549,N_17055,N_17113);
and U17550 (N_17550,N_17351,N_17309);
nand U17551 (N_17551,N_17002,N_17450);
or U17552 (N_17552,N_17367,N_17268);
xnor U17553 (N_17553,N_17250,N_17189);
nand U17554 (N_17554,N_17181,N_17301);
or U17555 (N_17555,N_17403,N_17102);
nor U17556 (N_17556,N_17001,N_17154);
or U17557 (N_17557,N_17420,N_17020);
xnor U17558 (N_17558,N_17350,N_17076);
and U17559 (N_17559,N_17310,N_17114);
nand U17560 (N_17560,N_17330,N_17149);
xnor U17561 (N_17561,N_17251,N_17077);
and U17562 (N_17562,N_17359,N_17335);
xor U17563 (N_17563,N_17434,N_17246);
nand U17564 (N_17564,N_17380,N_17412);
xor U17565 (N_17565,N_17265,N_17223);
xnor U17566 (N_17566,N_17424,N_17042);
and U17567 (N_17567,N_17293,N_17135);
or U17568 (N_17568,N_17188,N_17063);
and U17569 (N_17569,N_17080,N_17186);
and U17570 (N_17570,N_17339,N_17230);
xor U17571 (N_17571,N_17428,N_17170);
and U17572 (N_17572,N_17304,N_17302);
and U17573 (N_17573,N_17197,N_17207);
and U17574 (N_17574,N_17185,N_17349);
xor U17575 (N_17575,N_17387,N_17404);
or U17576 (N_17576,N_17163,N_17123);
and U17577 (N_17577,N_17474,N_17345);
nand U17578 (N_17578,N_17382,N_17125);
nand U17579 (N_17579,N_17238,N_17432);
nand U17580 (N_17580,N_17091,N_17264);
and U17581 (N_17581,N_17066,N_17441);
nand U17582 (N_17582,N_17291,N_17361);
or U17583 (N_17583,N_17216,N_17005);
xor U17584 (N_17584,N_17004,N_17389);
and U17585 (N_17585,N_17324,N_17183);
or U17586 (N_17586,N_17485,N_17308);
xor U17587 (N_17587,N_17200,N_17252);
or U17588 (N_17588,N_17495,N_17262);
and U17589 (N_17589,N_17116,N_17006);
xnor U17590 (N_17590,N_17390,N_17152);
or U17591 (N_17591,N_17377,N_17488);
or U17592 (N_17592,N_17140,N_17413);
nand U17593 (N_17593,N_17333,N_17053);
and U17594 (N_17594,N_17212,N_17206);
xnor U17595 (N_17595,N_17033,N_17322);
or U17596 (N_17596,N_17289,N_17058);
nor U17597 (N_17597,N_17391,N_17127);
nor U17598 (N_17598,N_17104,N_17433);
nor U17599 (N_17599,N_17134,N_17278);
and U17600 (N_17600,N_17411,N_17373);
nand U17601 (N_17601,N_17316,N_17201);
xnor U17602 (N_17602,N_17087,N_17344);
xor U17603 (N_17603,N_17126,N_17342);
nor U17604 (N_17604,N_17294,N_17153);
nand U17605 (N_17605,N_17193,N_17015);
nor U17606 (N_17606,N_17052,N_17487);
and U17607 (N_17607,N_17041,N_17011);
and U17608 (N_17608,N_17271,N_17384);
xnor U17609 (N_17609,N_17047,N_17340);
or U17610 (N_17610,N_17470,N_17347);
nand U17611 (N_17611,N_17247,N_17022);
and U17612 (N_17612,N_17272,N_17353);
nor U17613 (N_17613,N_17472,N_17072);
nor U17614 (N_17614,N_17307,N_17281);
or U17615 (N_17615,N_17327,N_17492);
xnor U17616 (N_17616,N_17493,N_17184);
nand U17617 (N_17617,N_17379,N_17220);
and U17618 (N_17618,N_17036,N_17239);
xor U17619 (N_17619,N_17044,N_17249);
and U17620 (N_17620,N_17132,N_17463);
or U17621 (N_17621,N_17032,N_17090);
nand U17622 (N_17622,N_17095,N_17267);
xnor U17623 (N_17623,N_17017,N_17400);
and U17624 (N_17624,N_17235,N_17115);
nand U17625 (N_17625,N_17137,N_17205);
nand U17626 (N_17626,N_17435,N_17332);
nand U17627 (N_17627,N_17288,N_17071);
xnor U17628 (N_17628,N_17260,N_17180);
nand U17629 (N_17629,N_17101,N_17451);
nand U17630 (N_17630,N_17401,N_17275);
or U17631 (N_17631,N_17242,N_17173);
or U17632 (N_17632,N_17467,N_17171);
nand U17633 (N_17633,N_17225,N_17369);
nor U17634 (N_17634,N_17489,N_17343);
xnor U17635 (N_17635,N_17292,N_17145);
nor U17636 (N_17636,N_17431,N_17007);
and U17637 (N_17637,N_17446,N_17112);
nor U17638 (N_17638,N_17374,N_17217);
nor U17639 (N_17639,N_17073,N_17417);
xnor U17640 (N_17640,N_17442,N_17164);
xnor U17641 (N_17641,N_17144,N_17098);
and U17642 (N_17642,N_17346,N_17049);
xnor U17643 (N_17643,N_17438,N_17111);
or U17644 (N_17644,N_17471,N_17141);
and U17645 (N_17645,N_17426,N_17423);
and U17646 (N_17646,N_17449,N_17050);
xor U17647 (N_17647,N_17110,N_17224);
nand U17648 (N_17648,N_17160,N_17133);
nand U17649 (N_17649,N_17355,N_17051);
and U17650 (N_17650,N_17299,N_17290);
nor U17651 (N_17651,N_17084,N_17429);
or U17652 (N_17652,N_17348,N_17283);
nand U17653 (N_17653,N_17023,N_17277);
xnor U17654 (N_17654,N_17475,N_17108);
xor U17655 (N_17655,N_17097,N_17046);
and U17656 (N_17656,N_17009,N_17158);
or U17657 (N_17657,N_17458,N_17476);
nor U17658 (N_17658,N_17016,N_17416);
and U17659 (N_17659,N_17394,N_17018);
nand U17660 (N_17660,N_17026,N_17306);
xor U17661 (N_17661,N_17336,N_17305);
and U17662 (N_17662,N_17312,N_17139);
nand U17663 (N_17663,N_17393,N_17496);
nor U17664 (N_17664,N_17146,N_17150);
nor U17665 (N_17665,N_17447,N_17303);
nor U17666 (N_17666,N_17430,N_17147);
xnor U17667 (N_17667,N_17378,N_17148);
and U17668 (N_17668,N_17479,N_17280);
or U17669 (N_17669,N_17364,N_17103);
nor U17670 (N_17670,N_17284,N_17012);
nand U17671 (N_17671,N_17143,N_17088);
xnor U17672 (N_17672,N_17096,N_17122);
xnor U17673 (N_17673,N_17445,N_17024);
or U17674 (N_17674,N_17168,N_17427);
or U17675 (N_17675,N_17100,N_17402);
nor U17676 (N_17676,N_17236,N_17157);
nand U17677 (N_17677,N_17234,N_17392);
nand U17678 (N_17678,N_17440,N_17237);
nor U17679 (N_17679,N_17410,N_17372);
nand U17680 (N_17680,N_17419,N_17480);
nand U17681 (N_17681,N_17019,N_17421);
nor U17682 (N_17682,N_17065,N_17274);
nor U17683 (N_17683,N_17497,N_17151);
or U17684 (N_17684,N_17178,N_17255);
nand U17685 (N_17685,N_17159,N_17092);
and U17686 (N_17686,N_17182,N_17169);
nand U17687 (N_17687,N_17323,N_17120);
nor U17688 (N_17688,N_17128,N_17228);
xnor U17689 (N_17689,N_17254,N_17375);
or U17690 (N_17690,N_17494,N_17425);
xnor U17691 (N_17691,N_17166,N_17360);
and U17692 (N_17692,N_17085,N_17021);
nand U17693 (N_17693,N_17460,N_17407);
or U17694 (N_17694,N_17030,N_17320);
and U17695 (N_17695,N_17093,N_17338);
and U17696 (N_17696,N_17498,N_17273);
and U17697 (N_17697,N_17165,N_17191);
or U17698 (N_17698,N_17074,N_17341);
xor U17699 (N_17699,N_17043,N_17465);
or U17700 (N_17700,N_17035,N_17039);
xor U17701 (N_17701,N_17203,N_17027);
or U17702 (N_17702,N_17298,N_17204);
nor U17703 (N_17703,N_17259,N_17070);
nand U17704 (N_17704,N_17028,N_17356);
nand U17705 (N_17705,N_17192,N_17315);
nor U17706 (N_17706,N_17385,N_17231);
nor U17707 (N_17707,N_17117,N_17499);
or U17708 (N_17708,N_17226,N_17089);
nand U17709 (N_17709,N_17452,N_17454);
nand U17710 (N_17710,N_17279,N_17414);
xor U17711 (N_17711,N_17219,N_17398);
xor U17712 (N_17712,N_17029,N_17000);
xor U17713 (N_17713,N_17172,N_17325);
and U17714 (N_17714,N_17295,N_17483);
and U17715 (N_17715,N_17061,N_17266);
and U17716 (N_17716,N_17068,N_17486);
and U17717 (N_17717,N_17057,N_17318);
and U17718 (N_17718,N_17198,N_17209);
nor U17719 (N_17719,N_17119,N_17408);
xor U17720 (N_17720,N_17118,N_17083);
or U17721 (N_17721,N_17319,N_17484);
nor U17722 (N_17722,N_17376,N_17176);
nand U17723 (N_17723,N_17244,N_17136);
nor U17724 (N_17724,N_17453,N_17468);
nand U17725 (N_17725,N_17161,N_17357);
nand U17726 (N_17726,N_17199,N_17056);
xor U17727 (N_17727,N_17060,N_17210);
and U17728 (N_17728,N_17142,N_17156);
nand U17729 (N_17729,N_17037,N_17261);
nand U17730 (N_17730,N_17190,N_17444);
nor U17731 (N_17731,N_17366,N_17358);
nor U17732 (N_17732,N_17174,N_17248);
nand U17733 (N_17733,N_17287,N_17227);
and U17734 (N_17734,N_17221,N_17245);
or U17735 (N_17735,N_17106,N_17107);
xor U17736 (N_17736,N_17243,N_17094);
xnor U17737 (N_17737,N_17296,N_17314);
xnor U17738 (N_17738,N_17365,N_17286);
xnor U17739 (N_17739,N_17048,N_17241);
and U17740 (N_17740,N_17285,N_17195);
xnor U17741 (N_17741,N_17282,N_17436);
or U17742 (N_17742,N_17263,N_17448);
or U17743 (N_17743,N_17229,N_17464);
nor U17744 (N_17744,N_17399,N_17300);
xor U17745 (N_17745,N_17215,N_17175);
xor U17746 (N_17746,N_17099,N_17075);
xnor U17747 (N_17747,N_17395,N_17218);
nor U17748 (N_17748,N_17457,N_17130);
nor U17749 (N_17749,N_17371,N_17455);
and U17750 (N_17750,N_17235,N_17011);
or U17751 (N_17751,N_17266,N_17442);
or U17752 (N_17752,N_17250,N_17021);
nand U17753 (N_17753,N_17333,N_17151);
and U17754 (N_17754,N_17348,N_17146);
nand U17755 (N_17755,N_17323,N_17200);
nor U17756 (N_17756,N_17447,N_17182);
nand U17757 (N_17757,N_17440,N_17051);
nor U17758 (N_17758,N_17355,N_17450);
nor U17759 (N_17759,N_17385,N_17192);
nor U17760 (N_17760,N_17041,N_17478);
xnor U17761 (N_17761,N_17279,N_17172);
and U17762 (N_17762,N_17181,N_17051);
nor U17763 (N_17763,N_17153,N_17323);
nor U17764 (N_17764,N_17091,N_17305);
xnor U17765 (N_17765,N_17031,N_17361);
nor U17766 (N_17766,N_17045,N_17075);
xnor U17767 (N_17767,N_17228,N_17446);
nor U17768 (N_17768,N_17293,N_17144);
nand U17769 (N_17769,N_17339,N_17063);
xnor U17770 (N_17770,N_17480,N_17350);
and U17771 (N_17771,N_17361,N_17001);
xor U17772 (N_17772,N_17278,N_17246);
nand U17773 (N_17773,N_17364,N_17380);
xor U17774 (N_17774,N_17282,N_17315);
or U17775 (N_17775,N_17330,N_17138);
or U17776 (N_17776,N_17009,N_17208);
xor U17777 (N_17777,N_17118,N_17300);
xor U17778 (N_17778,N_17412,N_17487);
and U17779 (N_17779,N_17378,N_17097);
and U17780 (N_17780,N_17305,N_17129);
or U17781 (N_17781,N_17257,N_17250);
or U17782 (N_17782,N_17030,N_17369);
nor U17783 (N_17783,N_17258,N_17229);
or U17784 (N_17784,N_17311,N_17431);
nor U17785 (N_17785,N_17297,N_17410);
and U17786 (N_17786,N_17267,N_17311);
or U17787 (N_17787,N_17305,N_17286);
nor U17788 (N_17788,N_17171,N_17378);
or U17789 (N_17789,N_17314,N_17427);
nor U17790 (N_17790,N_17329,N_17036);
nor U17791 (N_17791,N_17235,N_17295);
nand U17792 (N_17792,N_17089,N_17229);
and U17793 (N_17793,N_17448,N_17245);
nand U17794 (N_17794,N_17170,N_17185);
and U17795 (N_17795,N_17238,N_17252);
nor U17796 (N_17796,N_17046,N_17498);
nor U17797 (N_17797,N_17015,N_17494);
and U17798 (N_17798,N_17004,N_17370);
or U17799 (N_17799,N_17374,N_17236);
or U17800 (N_17800,N_17158,N_17005);
nand U17801 (N_17801,N_17488,N_17359);
or U17802 (N_17802,N_17061,N_17337);
and U17803 (N_17803,N_17124,N_17424);
and U17804 (N_17804,N_17312,N_17343);
nand U17805 (N_17805,N_17470,N_17398);
nand U17806 (N_17806,N_17165,N_17294);
xor U17807 (N_17807,N_17049,N_17202);
nor U17808 (N_17808,N_17203,N_17428);
or U17809 (N_17809,N_17192,N_17040);
nor U17810 (N_17810,N_17005,N_17254);
xor U17811 (N_17811,N_17399,N_17194);
nand U17812 (N_17812,N_17104,N_17368);
nor U17813 (N_17813,N_17255,N_17080);
nor U17814 (N_17814,N_17321,N_17162);
nor U17815 (N_17815,N_17356,N_17388);
xor U17816 (N_17816,N_17031,N_17327);
and U17817 (N_17817,N_17384,N_17449);
and U17818 (N_17818,N_17366,N_17203);
and U17819 (N_17819,N_17211,N_17196);
xor U17820 (N_17820,N_17336,N_17187);
and U17821 (N_17821,N_17110,N_17176);
xnor U17822 (N_17822,N_17348,N_17097);
or U17823 (N_17823,N_17329,N_17469);
or U17824 (N_17824,N_17159,N_17317);
or U17825 (N_17825,N_17490,N_17180);
nand U17826 (N_17826,N_17194,N_17056);
xnor U17827 (N_17827,N_17306,N_17222);
and U17828 (N_17828,N_17070,N_17322);
or U17829 (N_17829,N_17020,N_17068);
and U17830 (N_17830,N_17093,N_17387);
nor U17831 (N_17831,N_17095,N_17496);
nor U17832 (N_17832,N_17128,N_17375);
and U17833 (N_17833,N_17033,N_17499);
nor U17834 (N_17834,N_17115,N_17474);
xor U17835 (N_17835,N_17234,N_17129);
nor U17836 (N_17836,N_17247,N_17082);
nor U17837 (N_17837,N_17143,N_17475);
and U17838 (N_17838,N_17471,N_17336);
and U17839 (N_17839,N_17433,N_17393);
and U17840 (N_17840,N_17181,N_17326);
nand U17841 (N_17841,N_17480,N_17460);
nand U17842 (N_17842,N_17039,N_17231);
nand U17843 (N_17843,N_17407,N_17223);
xor U17844 (N_17844,N_17072,N_17450);
and U17845 (N_17845,N_17281,N_17381);
or U17846 (N_17846,N_17449,N_17274);
xnor U17847 (N_17847,N_17398,N_17165);
and U17848 (N_17848,N_17081,N_17382);
nand U17849 (N_17849,N_17382,N_17466);
nor U17850 (N_17850,N_17127,N_17227);
xor U17851 (N_17851,N_17068,N_17199);
nor U17852 (N_17852,N_17238,N_17353);
or U17853 (N_17853,N_17393,N_17382);
xnor U17854 (N_17854,N_17378,N_17435);
xor U17855 (N_17855,N_17160,N_17159);
nand U17856 (N_17856,N_17460,N_17418);
or U17857 (N_17857,N_17218,N_17159);
xor U17858 (N_17858,N_17067,N_17402);
nand U17859 (N_17859,N_17340,N_17184);
or U17860 (N_17860,N_17045,N_17194);
and U17861 (N_17861,N_17215,N_17133);
or U17862 (N_17862,N_17441,N_17311);
xor U17863 (N_17863,N_17053,N_17349);
nand U17864 (N_17864,N_17157,N_17365);
nand U17865 (N_17865,N_17482,N_17492);
xor U17866 (N_17866,N_17456,N_17287);
and U17867 (N_17867,N_17170,N_17429);
and U17868 (N_17868,N_17351,N_17348);
xor U17869 (N_17869,N_17150,N_17305);
nand U17870 (N_17870,N_17241,N_17092);
nand U17871 (N_17871,N_17331,N_17436);
and U17872 (N_17872,N_17422,N_17051);
nor U17873 (N_17873,N_17358,N_17363);
nor U17874 (N_17874,N_17425,N_17364);
nand U17875 (N_17875,N_17253,N_17157);
xor U17876 (N_17876,N_17288,N_17122);
nand U17877 (N_17877,N_17186,N_17002);
or U17878 (N_17878,N_17026,N_17124);
and U17879 (N_17879,N_17279,N_17053);
nor U17880 (N_17880,N_17093,N_17070);
nor U17881 (N_17881,N_17196,N_17345);
nor U17882 (N_17882,N_17320,N_17054);
or U17883 (N_17883,N_17442,N_17012);
nor U17884 (N_17884,N_17141,N_17053);
or U17885 (N_17885,N_17194,N_17143);
nor U17886 (N_17886,N_17237,N_17432);
or U17887 (N_17887,N_17311,N_17065);
and U17888 (N_17888,N_17059,N_17197);
nor U17889 (N_17889,N_17447,N_17322);
xor U17890 (N_17890,N_17449,N_17393);
nand U17891 (N_17891,N_17228,N_17301);
or U17892 (N_17892,N_17036,N_17392);
and U17893 (N_17893,N_17202,N_17278);
and U17894 (N_17894,N_17480,N_17389);
or U17895 (N_17895,N_17084,N_17037);
nand U17896 (N_17896,N_17281,N_17249);
nor U17897 (N_17897,N_17426,N_17416);
nor U17898 (N_17898,N_17146,N_17455);
nand U17899 (N_17899,N_17151,N_17005);
or U17900 (N_17900,N_17436,N_17151);
nand U17901 (N_17901,N_17130,N_17369);
nand U17902 (N_17902,N_17176,N_17324);
xnor U17903 (N_17903,N_17302,N_17403);
nand U17904 (N_17904,N_17410,N_17302);
and U17905 (N_17905,N_17064,N_17092);
xor U17906 (N_17906,N_17208,N_17317);
or U17907 (N_17907,N_17105,N_17040);
and U17908 (N_17908,N_17136,N_17316);
xor U17909 (N_17909,N_17164,N_17398);
nand U17910 (N_17910,N_17358,N_17454);
xnor U17911 (N_17911,N_17435,N_17329);
xnor U17912 (N_17912,N_17156,N_17417);
nand U17913 (N_17913,N_17388,N_17209);
and U17914 (N_17914,N_17413,N_17261);
nor U17915 (N_17915,N_17278,N_17044);
nand U17916 (N_17916,N_17290,N_17175);
nand U17917 (N_17917,N_17073,N_17330);
or U17918 (N_17918,N_17216,N_17411);
xor U17919 (N_17919,N_17181,N_17307);
or U17920 (N_17920,N_17475,N_17139);
nand U17921 (N_17921,N_17115,N_17250);
or U17922 (N_17922,N_17085,N_17382);
and U17923 (N_17923,N_17146,N_17181);
nand U17924 (N_17924,N_17126,N_17495);
xnor U17925 (N_17925,N_17476,N_17039);
xnor U17926 (N_17926,N_17153,N_17337);
and U17927 (N_17927,N_17113,N_17354);
nor U17928 (N_17928,N_17233,N_17189);
nand U17929 (N_17929,N_17124,N_17050);
nand U17930 (N_17930,N_17213,N_17194);
or U17931 (N_17931,N_17210,N_17404);
xor U17932 (N_17932,N_17266,N_17315);
and U17933 (N_17933,N_17342,N_17414);
nand U17934 (N_17934,N_17287,N_17171);
nand U17935 (N_17935,N_17118,N_17123);
or U17936 (N_17936,N_17224,N_17122);
nor U17937 (N_17937,N_17234,N_17199);
nand U17938 (N_17938,N_17000,N_17087);
xnor U17939 (N_17939,N_17035,N_17406);
nor U17940 (N_17940,N_17323,N_17365);
nor U17941 (N_17941,N_17283,N_17158);
nor U17942 (N_17942,N_17398,N_17159);
or U17943 (N_17943,N_17281,N_17274);
nor U17944 (N_17944,N_17052,N_17033);
and U17945 (N_17945,N_17229,N_17411);
xor U17946 (N_17946,N_17405,N_17310);
nand U17947 (N_17947,N_17180,N_17431);
xnor U17948 (N_17948,N_17155,N_17120);
nor U17949 (N_17949,N_17103,N_17462);
nand U17950 (N_17950,N_17256,N_17177);
nor U17951 (N_17951,N_17353,N_17412);
xor U17952 (N_17952,N_17110,N_17248);
xnor U17953 (N_17953,N_17285,N_17376);
or U17954 (N_17954,N_17434,N_17142);
nand U17955 (N_17955,N_17495,N_17354);
or U17956 (N_17956,N_17077,N_17194);
and U17957 (N_17957,N_17112,N_17462);
and U17958 (N_17958,N_17105,N_17336);
and U17959 (N_17959,N_17288,N_17037);
nor U17960 (N_17960,N_17191,N_17337);
nand U17961 (N_17961,N_17293,N_17467);
and U17962 (N_17962,N_17063,N_17167);
or U17963 (N_17963,N_17201,N_17205);
xor U17964 (N_17964,N_17264,N_17028);
nor U17965 (N_17965,N_17402,N_17128);
nand U17966 (N_17966,N_17272,N_17133);
or U17967 (N_17967,N_17107,N_17318);
and U17968 (N_17968,N_17044,N_17257);
nand U17969 (N_17969,N_17251,N_17148);
or U17970 (N_17970,N_17323,N_17367);
or U17971 (N_17971,N_17496,N_17355);
and U17972 (N_17972,N_17254,N_17048);
nand U17973 (N_17973,N_17157,N_17295);
or U17974 (N_17974,N_17305,N_17192);
xnor U17975 (N_17975,N_17004,N_17219);
nand U17976 (N_17976,N_17404,N_17151);
or U17977 (N_17977,N_17229,N_17005);
nand U17978 (N_17978,N_17050,N_17152);
nand U17979 (N_17979,N_17400,N_17060);
nor U17980 (N_17980,N_17432,N_17164);
or U17981 (N_17981,N_17444,N_17305);
or U17982 (N_17982,N_17406,N_17012);
or U17983 (N_17983,N_17000,N_17242);
and U17984 (N_17984,N_17354,N_17216);
nand U17985 (N_17985,N_17055,N_17050);
nand U17986 (N_17986,N_17293,N_17081);
xnor U17987 (N_17987,N_17103,N_17162);
or U17988 (N_17988,N_17353,N_17361);
nor U17989 (N_17989,N_17421,N_17388);
xor U17990 (N_17990,N_17113,N_17375);
and U17991 (N_17991,N_17201,N_17387);
nand U17992 (N_17992,N_17117,N_17481);
or U17993 (N_17993,N_17301,N_17293);
nand U17994 (N_17994,N_17086,N_17224);
and U17995 (N_17995,N_17481,N_17061);
or U17996 (N_17996,N_17105,N_17056);
xor U17997 (N_17997,N_17369,N_17079);
and U17998 (N_17998,N_17056,N_17355);
xnor U17999 (N_17999,N_17060,N_17198);
and U18000 (N_18000,N_17511,N_17869);
xnor U18001 (N_18001,N_17853,N_17964);
and U18002 (N_18002,N_17927,N_17648);
and U18003 (N_18003,N_17737,N_17647);
or U18004 (N_18004,N_17980,N_17658);
xnor U18005 (N_18005,N_17947,N_17973);
nand U18006 (N_18006,N_17761,N_17575);
nor U18007 (N_18007,N_17940,N_17549);
and U18008 (N_18008,N_17969,N_17729);
and U18009 (N_18009,N_17736,N_17856);
nand U18010 (N_18010,N_17509,N_17991);
nand U18011 (N_18011,N_17829,N_17556);
or U18012 (N_18012,N_17816,N_17982);
nor U18013 (N_18013,N_17653,N_17772);
or U18014 (N_18014,N_17855,N_17941);
or U18015 (N_18015,N_17907,N_17974);
xnor U18016 (N_18016,N_17608,N_17680);
nor U18017 (N_18017,N_17847,N_17850);
or U18018 (N_18018,N_17779,N_17603);
xnor U18019 (N_18019,N_17713,N_17780);
nand U18020 (N_18020,N_17600,N_17985);
nor U18021 (N_18021,N_17815,N_17615);
or U18022 (N_18022,N_17983,N_17895);
and U18023 (N_18023,N_17684,N_17687);
and U18024 (N_18024,N_17611,N_17538);
or U18025 (N_18025,N_17748,N_17958);
nand U18026 (N_18026,N_17832,N_17609);
and U18027 (N_18027,N_17759,N_17524);
xnor U18028 (N_18028,N_17763,N_17764);
and U18029 (N_18029,N_17630,N_17614);
nor U18030 (N_18030,N_17904,N_17861);
or U18031 (N_18031,N_17786,N_17837);
nor U18032 (N_18032,N_17826,N_17714);
and U18033 (N_18033,N_17698,N_17688);
and U18034 (N_18034,N_17507,N_17744);
or U18035 (N_18035,N_17915,N_17866);
nand U18036 (N_18036,N_17734,N_17751);
xor U18037 (N_18037,N_17757,N_17876);
or U18038 (N_18038,N_17552,N_17694);
xor U18039 (N_18039,N_17703,N_17732);
and U18040 (N_18040,N_17650,N_17702);
xnor U18041 (N_18041,N_17811,N_17889);
nor U18042 (N_18042,N_17669,N_17957);
and U18043 (N_18043,N_17929,N_17508);
or U18044 (N_18044,N_17785,N_17537);
nand U18045 (N_18045,N_17840,N_17818);
xnor U18046 (N_18046,N_17994,N_17890);
and U18047 (N_18047,N_17674,N_17776);
xor U18048 (N_18048,N_17920,N_17789);
nand U18049 (N_18049,N_17717,N_17733);
xnor U18050 (N_18050,N_17823,N_17749);
nor U18051 (N_18051,N_17635,N_17543);
and U18052 (N_18052,N_17835,N_17949);
nand U18053 (N_18053,N_17705,N_17926);
and U18054 (N_18054,N_17622,N_17555);
xor U18055 (N_18055,N_17760,N_17607);
and U18056 (N_18056,N_17930,N_17762);
nor U18057 (N_18057,N_17577,N_17953);
xnor U18058 (N_18058,N_17978,N_17629);
and U18059 (N_18059,N_17682,N_17659);
nand U18060 (N_18060,N_17743,N_17568);
nor U18061 (N_18061,N_17945,N_17546);
and U18062 (N_18062,N_17649,N_17988);
nor U18063 (N_18063,N_17894,N_17578);
and U18064 (N_18064,N_17886,N_17725);
or U18065 (N_18065,N_17710,N_17916);
nand U18066 (N_18066,N_17867,N_17989);
and U18067 (N_18067,N_17673,N_17632);
and U18068 (N_18068,N_17986,N_17881);
xor U18069 (N_18069,N_17672,N_17571);
xnor U18070 (N_18070,N_17750,N_17505);
or U18071 (N_18071,N_17686,N_17944);
nor U18072 (N_18072,N_17821,N_17896);
and U18073 (N_18073,N_17868,N_17726);
nor U18074 (N_18074,N_17767,N_17828);
nor U18075 (N_18075,N_17951,N_17965);
and U18076 (N_18076,N_17846,N_17962);
nand U18077 (N_18077,N_17919,N_17665);
nor U18078 (N_18078,N_17553,N_17690);
nor U18079 (N_18079,N_17917,N_17834);
or U18080 (N_18080,N_17641,N_17996);
nor U18081 (N_18081,N_17654,N_17778);
nor U18082 (N_18082,N_17851,N_17643);
xor U18083 (N_18083,N_17583,N_17668);
and U18084 (N_18084,N_17848,N_17874);
nand U18085 (N_18085,N_17987,N_17602);
nor U18086 (N_18086,N_17955,N_17598);
nand U18087 (N_18087,N_17731,N_17975);
nor U18088 (N_18088,N_17746,N_17597);
or U18089 (N_18089,N_17822,N_17783);
xor U18090 (N_18090,N_17715,N_17679);
xor U18091 (N_18091,N_17681,N_17753);
xnor U18092 (N_18092,N_17937,N_17970);
xnor U18093 (N_18093,N_17616,N_17662);
and U18094 (N_18094,N_17666,N_17843);
and U18095 (N_18095,N_17845,N_17661);
nor U18096 (N_18096,N_17706,N_17569);
xor U18097 (N_18097,N_17923,N_17745);
and U18098 (N_18098,N_17638,N_17685);
or U18099 (N_18099,N_17993,N_17925);
or U18100 (N_18100,N_17592,N_17799);
and U18101 (N_18101,N_17901,N_17908);
or U18102 (N_18102,N_17839,N_17523);
nand U18103 (N_18103,N_17747,N_17884);
xnor U18104 (N_18104,N_17900,N_17514);
nor U18105 (N_18105,N_17977,N_17961);
nor U18106 (N_18106,N_17708,N_17527);
nor U18107 (N_18107,N_17709,N_17660);
and U18108 (N_18108,N_17513,N_17581);
xor U18109 (N_18109,N_17879,N_17652);
and U18110 (N_18110,N_17812,N_17551);
nand U18111 (N_18111,N_17590,N_17824);
or U18112 (N_18112,N_17701,N_17781);
xnor U18113 (N_18113,N_17677,N_17536);
nand U18114 (N_18114,N_17863,N_17515);
or U18115 (N_18115,N_17601,N_17981);
and U18116 (N_18116,N_17535,N_17898);
nor U18117 (N_18117,N_17612,N_17695);
or U18118 (N_18118,N_17588,N_17586);
nand U18119 (N_18119,N_17642,N_17932);
xor U18120 (N_18120,N_17563,N_17992);
nor U18121 (N_18121,N_17872,N_17939);
and U18122 (N_18122,N_17921,N_17624);
and U18123 (N_18123,N_17959,N_17864);
xnor U18124 (N_18124,N_17842,N_17885);
nor U18125 (N_18125,N_17873,N_17663);
nand U18126 (N_18126,N_17558,N_17765);
xnor U18127 (N_18127,N_17548,N_17880);
nor U18128 (N_18128,N_17903,N_17712);
and U18129 (N_18129,N_17999,N_17802);
or U18130 (N_18130,N_17860,N_17503);
or U18131 (N_18131,N_17865,N_17678);
or U18132 (N_18132,N_17591,N_17722);
or U18133 (N_18133,N_17562,N_17573);
nor U18134 (N_18134,N_17526,N_17979);
or U18135 (N_18135,N_17596,N_17814);
nand U18136 (N_18136,N_17567,N_17516);
nand U18137 (N_18137,N_17631,N_17777);
xor U18138 (N_18138,N_17956,N_17875);
xor U18139 (N_18139,N_17950,N_17912);
nor U18140 (N_18140,N_17773,N_17887);
nand U18141 (N_18141,N_17792,N_17948);
nor U18142 (N_18142,N_17617,N_17878);
nand U18143 (N_18143,N_17531,N_17984);
and U18144 (N_18144,N_17740,N_17905);
nor U18145 (N_18145,N_17530,N_17730);
nand U18146 (N_18146,N_17707,N_17911);
nand U18147 (N_18147,N_17877,N_17582);
or U18148 (N_18148,N_17522,N_17804);
or U18149 (N_18149,N_17532,N_17599);
and U18150 (N_18150,N_17791,N_17692);
nor U18151 (N_18151,N_17790,N_17796);
nor U18152 (N_18152,N_17933,N_17914);
xor U18153 (N_18153,N_17998,N_17613);
or U18154 (N_18154,N_17623,N_17805);
and U18155 (N_18155,N_17644,N_17836);
xor U18156 (N_18156,N_17554,N_17724);
nand U18157 (N_18157,N_17892,N_17794);
xnor U18158 (N_18158,N_17542,N_17931);
and U18159 (N_18159,N_17807,N_17620);
or U18160 (N_18160,N_17651,N_17852);
nor U18161 (N_18161,N_17938,N_17766);
nor U18162 (N_18162,N_17533,N_17954);
nand U18163 (N_18163,N_17589,N_17817);
or U18164 (N_18164,N_17723,N_17990);
or U18165 (N_18165,N_17606,N_17858);
nand U18166 (N_18166,N_17557,N_17906);
nor U18167 (N_18167,N_17946,N_17528);
xor U18168 (N_18168,N_17995,N_17691);
xor U18169 (N_18169,N_17518,N_17891);
nor U18170 (N_18170,N_17899,N_17711);
nor U18171 (N_18171,N_17547,N_17771);
and U18172 (N_18172,N_17689,N_17803);
nand U18173 (N_18173,N_17539,N_17862);
nor U18174 (N_18174,N_17909,N_17593);
nor U18175 (N_18175,N_17883,N_17605);
or U18176 (N_18176,N_17810,N_17844);
xnor U18177 (N_18177,N_17699,N_17645);
and U18178 (N_18178,N_17768,N_17667);
nor U18179 (N_18179,N_17519,N_17693);
xor U18180 (N_18180,N_17512,N_17676);
nand U18181 (N_18181,N_17838,N_17727);
nor U18182 (N_18182,N_17656,N_17797);
and U18183 (N_18183,N_17870,N_17640);
nor U18184 (N_18184,N_17774,N_17570);
or U18185 (N_18185,N_17627,N_17968);
nand U18186 (N_18186,N_17700,N_17566);
and U18187 (N_18187,N_17902,N_17756);
nand U18188 (N_18188,N_17752,N_17997);
xor U18189 (N_18189,N_17971,N_17500);
nor U18190 (N_18190,N_17718,N_17888);
or U18191 (N_18191,N_17739,N_17960);
or U18192 (N_18192,N_17859,N_17897);
xnor U18193 (N_18193,N_17913,N_17720);
and U18194 (N_18194,N_17545,N_17671);
xnor U18195 (N_18195,N_17541,N_17857);
or U18196 (N_18196,N_17936,N_17664);
and U18197 (N_18197,N_17626,N_17741);
nand U18198 (N_18198,N_17621,N_17830);
nand U18199 (N_18199,N_17935,N_17738);
nand U18200 (N_18200,N_17910,N_17587);
nor U18201 (N_18201,N_17560,N_17628);
and U18202 (N_18202,N_17625,N_17572);
nand U18203 (N_18203,N_17634,N_17809);
xor U18204 (N_18204,N_17517,N_17934);
xnor U18205 (N_18205,N_17924,N_17800);
nand U18206 (N_18206,N_17893,N_17520);
nand U18207 (N_18207,N_17976,N_17928);
or U18208 (N_18208,N_17882,N_17683);
or U18209 (N_18209,N_17559,N_17637);
and U18210 (N_18210,N_17827,N_17579);
xnor U18211 (N_18211,N_17550,N_17521);
xnor U18212 (N_18212,N_17604,N_17501);
xnor U18213 (N_18213,N_17833,N_17655);
or U18214 (N_18214,N_17716,N_17967);
nor U18215 (N_18215,N_17854,N_17825);
xor U18216 (N_18216,N_17952,N_17942);
nor U18217 (N_18217,N_17584,N_17704);
nor U18218 (N_18218,N_17849,N_17831);
nand U18219 (N_18219,N_17788,N_17742);
nor U18220 (N_18220,N_17534,N_17639);
xnor U18221 (N_18221,N_17594,N_17721);
and U18222 (N_18222,N_17793,N_17574);
and U18223 (N_18223,N_17782,N_17755);
and U18224 (N_18224,N_17697,N_17610);
or U18225 (N_18225,N_17719,N_17544);
nand U18226 (N_18226,N_17580,N_17696);
nor U18227 (N_18227,N_17670,N_17775);
nor U18228 (N_18228,N_17922,N_17595);
nor U18229 (N_18229,N_17529,N_17758);
or U18230 (N_18230,N_17564,N_17841);
nor U18231 (N_18231,N_17798,N_17795);
xnor U18232 (N_18232,N_17769,N_17728);
and U18233 (N_18233,N_17806,N_17506);
and U18234 (N_18234,N_17871,N_17675);
and U18235 (N_18235,N_17633,N_17813);
nand U18236 (N_18236,N_17754,N_17618);
nor U18237 (N_18237,N_17801,N_17502);
nor U18238 (N_18238,N_17504,N_17808);
nor U18239 (N_18239,N_17585,N_17943);
and U18240 (N_18240,N_17619,N_17565);
and U18241 (N_18241,N_17784,N_17525);
nand U18242 (N_18242,N_17770,N_17787);
nor U18243 (N_18243,N_17576,N_17820);
nor U18244 (N_18244,N_17657,N_17918);
xnor U18245 (N_18245,N_17561,N_17972);
nand U18246 (N_18246,N_17735,N_17646);
nand U18247 (N_18247,N_17819,N_17636);
and U18248 (N_18248,N_17966,N_17540);
nand U18249 (N_18249,N_17510,N_17963);
nand U18250 (N_18250,N_17991,N_17874);
and U18251 (N_18251,N_17962,N_17604);
xor U18252 (N_18252,N_17951,N_17789);
xnor U18253 (N_18253,N_17676,N_17627);
nand U18254 (N_18254,N_17996,N_17743);
nor U18255 (N_18255,N_17653,N_17604);
nand U18256 (N_18256,N_17955,N_17762);
nand U18257 (N_18257,N_17945,N_17750);
and U18258 (N_18258,N_17567,N_17853);
nand U18259 (N_18259,N_17773,N_17552);
nor U18260 (N_18260,N_17501,N_17695);
and U18261 (N_18261,N_17686,N_17649);
nand U18262 (N_18262,N_17797,N_17775);
and U18263 (N_18263,N_17999,N_17526);
nand U18264 (N_18264,N_17947,N_17912);
nor U18265 (N_18265,N_17518,N_17924);
xnor U18266 (N_18266,N_17624,N_17928);
nor U18267 (N_18267,N_17703,N_17576);
nor U18268 (N_18268,N_17616,N_17736);
or U18269 (N_18269,N_17795,N_17609);
nor U18270 (N_18270,N_17550,N_17912);
and U18271 (N_18271,N_17619,N_17516);
and U18272 (N_18272,N_17843,N_17955);
nor U18273 (N_18273,N_17573,N_17717);
nor U18274 (N_18274,N_17929,N_17706);
and U18275 (N_18275,N_17519,N_17902);
nand U18276 (N_18276,N_17572,N_17604);
nor U18277 (N_18277,N_17761,N_17794);
or U18278 (N_18278,N_17587,N_17893);
nand U18279 (N_18279,N_17910,N_17755);
nor U18280 (N_18280,N_17653,N_17640);
nor U18281 (N_18281,N_17773,N_17781);
xor U18282 (N_18282,N_17572,N_17833);
nor U18283 (N_18283,N_17776,N_17954);
nor U18284 (N_18284,N_17735,N_17849);
nor U18285 (N_18285,N_17658,N_17817);
nand U18286 (N_18286,N_17600,N_17579);
nor U18287 (N_18287,N_17702,N_17891);
and U18288 (N_18288,N_17803,N_17545);
and U18289 (N_18289,N_17947,N_17893);
nor U18290 (N_18290,N_17572,N_17658);
xnor U18291 (N_18291,N_17501,N_17738);
or U18292 (N_18292,N_17515,N_17585);
nand U18293 (N_18293,N_17681,N_17876);
and U18294 (N_18294,N_17747,N_17656);
nor U18295 (N_18295,N_17825,N_17999);
or U18296 (N_18296,N_17684,N_17805);
or U18297 (N_18297,N_17650,N_17786);
and U18298 (N_18298,N_17828,N_17715);
nor U18299 (N_18299,N_17666,N_17625);
nand U18300 (N_18300,N_17880,N_17993);
nand U18301 (N_18301,N_17927,N_17617);
nand U18302 (N_18302,N_17884,N_17603);
nor U18303 (N_18303,N_17675,N_17980);
nand U18304 (N_18304,N_17937,N_17580);
and U18305 (N_18305,N_17608,N_17765);
xor U18306 (N_18306,N_17934,N_17859);
and U18307 (N_18307,N_17569,N_17774);
nand U18308 (N_18308,N_17804,N_17686);
and U18309 (N_18309,N_17797,N_17846);
and U18310 (N_18310,N_17784,N_17816);
nand U18311 (N_18311,N_17861,N_17731);
nor U18312 (N_18312,N_17667,N_17731);
and U18313 (N_18313,N_17995,N_17746);
or U18314 (N_18314,N_17721,N_17933);
or U18315 (N_18315,N_17997,N_17949);
xnor U18316 (N_18316,N_17756,N_17989);
nor U18317 (N_18317,N_17874,N_17841);
nor U18318 (N_18318,N_17611,N_17698);
or U18319 (N_18319,N_17958,N_17728);
and U18320 (N_18320,N_17758,N_17514);
and U18321 (N_18321,N_17762,N_17995);
and U18322 (N_18322,N_17523,N_17518);
nand U18323 (N_18323,N_17627,N_17639);
nor U18324 (N_18324,N_17849,N_17975);
and U18325 (N_18325,N_17557,N_17699);
or U18326 (N_18326,N_17930,N_17810);
and U18327 (N_18327,N_17950,N_17581);
xnor U18328 (N_18328,N_17717,N_17581);
nor U18329 (N_18329,N_17506,N_17655);
xnor U18330 (N_18330,N_17757,N_17893);
and U18331 (N_18331,N_17934,N_17804);
or U18332 (N_18332,N_17783,N_17877);
nand U18333 (N_18333,N_17815,N_17967);
nor U18334 (N_18334,N_17887,N_17714);
and U18335 (N_18335,N_17807,N_17693);
and U18336 (N_18336,N_17547,N_17663);
or U18337 (N_18337,N_17852,N_17888);
or U18338 (N_18338,N_17899,N_17753);
and U18339 (N_18339,N_17861,N_17863);
nor U18340 (N_18340,N_17961,N_17844);
or U18341 (N_18341,N_17760,N_17828);
xnor U18342 (N_18342,N_17651,N_17923);
xnor U18343 (N_18343,N_17796,N_17972);
or U18344 (N_18344,N_17853,N_17903);
nor U18345 (N_18345,N_17871,N_17757);
or U18346 (N_18346,N_17790,N_17552);
and U18347 (N_18347,N_17897,N_17656);
and U18348 (N_18348,N_17786,N_17651);
or U18349 (N_18349,N_17888,N_17561);
or U18350 (N_18350,N_17502,N_17828);
nand U18351 (N_18351,N_17603,N_17502);
nand U18352 (N_18352,N_17581,N_17561);
xor U18353 (N_18353,N_17538,N_17573);
nand U18354 (N_18354,N_17572,N_17518);
or U18355 (N_18355,N_17914,N_17937);
or U18356 (N_18356,N_17862,N_17637);
or U18357 (N_18357,N_17882,N_17607);
nand U18358 (N_18358,N_17615,N_17589);
nand U18359 (N_18359,N_17982,N_17963);
xnor U18360 (N_18360,N_17825,N_17626);
and U18361 (N_18361,N_17639,N_17817);
or U18362 (N_18362,N_17542,N_17539);
nor U18363 (N_18363,N_17689,N_17970);
and U18364 (N_18364,N_17945,N_17899);
xnor U18365 (N_18365,N_17979,N_17764);
nand U18366 (N_18366,N_17892,N_17987);
xor U18367 (N_18367,N_17840,N_17585);
xnor U18368 (N_18368,N_17909,N_17730);
or U18369 (N_18369,N_17575,N_17915);
or U18370 (N_18370,N_17630,N_17652);
nor U18371 (N_18371,N_17765,N_17824);
or U18372 (N_18372,N_17969,N_17662);
nor U18373 (N_18373,N_17612,N_17571);
xnor U18374 (N_18374,N_17833,N_17807);
xnor U18375 (N_18375,N_17668,N_17660);
nor U18376 (N_18376,N_17832,N_17999);
nor U18377 (N_18377,N_17771,N_17503);
and U18378 (N_18378,N_17988,N_17578);
nor U18379 (N_18379,N_17567,N_17575);
and U18380 (N_18380,N_17904,N_17926);
nor U18381 (N_18381,N_17672,N_17938);
nand U18382 (N_18382,N_17633,N_17759);
xor U18383 (N_18383,N_17550,N_17730);
xnor U18384 (N_18384,N_17626,N_17952);
xor U18385 (N_18385,N_17631,N_17913);
xor U18386 (N_18386,N_17952,N_17871);
and U18387 (N_18387,N_17981,N_17534);
nand U18388 (N_18388,N_17647,N_17868);
nor U18389 (N_18389,N_17799,N_17895);
nor U18390 (N_18390,N_17986,N_17717);
nand U18391 (N_18391,N_17858,N_17847);
or U18392 (N_18392,N_17902,N_17811);
and U18393 (N_18393,N_17708,N_17659);
nand U18394 (N_18394,N_17576,N_17885);
nand U18395 (N_18395,N_17718,N_17855);
and U18396 (N_18396,N_17885,N_17913);
nor U18397 (N_18397,N_17536,N_17604);
nor U18398 (N_18398,N_17501,N_17674);
or U18399 (N_18399,N_17969,N_17839);
nor U18400 (N_18400,N_17920,N_17626);
or U18401 (N_18401,N_17689,N_17702);
nor U18402 (N_18402,N_17665,N_17570);
xnor U18403 (N_18403,N_17930,N_17669);
or U18404 (N_18404,N_17966,N_17775);
and U18405 (N_18405,N_17894,N_17807);
xor U18406 (N_18406,N_17588,N_17851);
xnor U18407 (N_18407,N_17685,N_17641);
or U18408 (N_18408,N_17550,N_17902);
xnor U18409 (N_18409,N_17976,N_17753);
nand U18410 (N_18410,N_17548,N_17749);
xor U18411 (N_18411,N_17785,N_17761);
or U18412 (N_18412,N_17806,N_17893);
nand U18413 (N_18413,N_17502,N_17706);
and U18414 (N_18414,N_17743,N_17727);
xnor U18415 (N_18415,N_17703,N_17730);
or U18416 (N_18416,N_17914,N_17765);
nand U18417 (N_18417,N_17676,N_17574);
xnor U18418 (N_18418,N_17749,N_17995);
or U18419 (N_18419,N_17764,N_17749);
xor U18420 (N_18420,N_17591,N_17766);
and U18421 (N_18421,N_17727,N_17661);
nor U18422 (N_18422,N_17783,N_17608);
and U18423 (N_18423,N_17504,N_17519);
or U18424 (N_18424,N_17929,N_17703);
xor U18425 (N_18425,N_17892,N_17809);
and U18426 (N_18426,N_17543,N_17958);
nor U18427 (N_18427,N_17926,N_17776);
nand U18428 (N_18428,N_17841,N_17916);
and U18429 (N_18429,N_17958,N_17707);
or U18430 (N_18430,N_17824,N_17763);
and U18431 (N_18431,N_17801,N_17712);
nand U18432 (N_18432,N_17559,N_17877);
and U18433 (N_18433,N_17739,N_17677);
and U18434 (N_18434,N_17931,N_17582);
xnor U18435 (N_18435,N_17681,N_17881);
nor U18436 (N_18436,N_17793,N_17588);
xnor U18437 (N_18437,N_17800,N_17860);
nand U18438 (N_18438,N_17611,N_17861);
nor U18439 (N_18439,N_17715,N_17856);
and U18440 (N_18440,N_17987,N_17718);
nor U18441 (N_18441,N_17783,N_17687);
xor U18442 (N_18442,N_17870,N_17522);
nor U18443 (N_18443,N_17659,N_17770);
nor U18444 (N_18444,N_17968,N_17911);
and U18445 (N_18445,N_17946,N_17989);
or U18446 (N_18446,N_17538,N_17586);
and U18447 (N_18447,N_17616,N_17948);
nor U18448 (N_18448,N_17646,N_17854);
and U18449 (N_18449,N_17868,N_17834);
xnor U18450 (N_18450,N_17858,N_17546);
or U18451 (N_18451,N_17726,N_17906);
or U18452 (N_18452,N_17856,N_17843);
nor U18453 (N_18453,N_17658,N_17637);
and U18454 (N_18454,N_17596,N_17750);
nand U18455 (N_18455,N_17734,N_17828);
or U18456 (N_18456,N_17681,N_17603);
nand U18457 (N_18457,N_17791,N_17515);
nor U18458 (N_18458,N_17987,N_17656);
nor U18459 (N_18459,N_17632,N_17799);
xor U18460 (N_18460,N_17678,N_17636);
nor U18461 (N_18461,N_17592,N_17996);
nor U18462 (N_18462,N_17508,N_17819);
nor U18463 (N_18463,N_17861,N_17640);
xor U18464 (N_18464,N_17766,N_17709);
xor U18465 (N_18465,N_17981,N_17795);
and U18466 (N_18466,N_17815,N_17766);
and U18467 (N_18467,N_17884,N_17546);
nor U18468 (N_18468,N_17525,N_17616);
or U18469 (N_18469,N_17746,N_17885);
nand U18470 (N_18470,N_17911,N_17712);
nor U18471 (N_18471,N_17659,N_17623);
and U18472 (N_18472,N_17519,N_17927);
xnor U18473 (N_18473,N_17937,N_17659);
and U18474 (N_18474,N_17873,N_17960);
nand U18475 (N_18475,N_17560,N_17906);
or U18476 (N_18476,N_17770,N_17548);
xnor U18477 (N_18477,N_17934,N_17978);
and U18478 (N_18478,N_17836,N_17843);
nor U18479 (N_18479,N_17989,N_17795);
and U18480 (N_18480,N_17826,N_17588);
nor U18481 (N_18481,N_17871,N_17710);
xnor U18482 (N_18482,N_17823,N_17954);
nand U18483 (N_18483,N_17701,N_17688);
and U18484 (N_18484,N_17585,N_17615);
or U18485 (N_18485,N_17852,N_17596);
nand U18486 (N_18486,N_17982,N_17967);
nand U18487 (N_18487,N_17613,N_17843);
and U18488 (N_18488,N_17747,N_17897);
xor U18489 (N_18489,N_17847,N_17862);
and U18490 (N_18490,N_17520,N_17697);
and U18491 (N_18491,N_17634,N_17733);
and U18492 (N_18492,N_17757,N_17937);
xnor U18493 (N_18493,N_17735,N_17957);
and U18494 (N_18494,N_17835,N_17776);
nor U18495 (N_18495,N_17893,N_17656);
xor U18496 (N_18496,N_17724,N_17927);
or U18497 (N_18497,N_17562,N_17770);
or U18498 (N_18498,N_17604,N_17999);
or U18499 (N_18499,N_17963,N_17700);
or U18500 (N_18500,N_18368,N_18202);
or U18501 (N_18501,N_18379,N_18410);
or U18502 (N_18502,N_18355,N_18424);
nor U18503 (N_18503,N_18108,N_18405);
nor U18504 (N_18504,N_18026,N_18011);
nand U18505 (N_18505,N_18012,N_18003);
or U18506 (N_18506,N_18371,N_18065);
xnor U18507 (N_18507,N_18138,N_18354);
and U18508 (N_18508,N_18177,N_18269);
xnor U18509 (N_18509,N_18334,N_18459);
nand U18510 (N_18510,N_18057,N_18312);
and U18511 (N_18511,N_18275,N_18062);
nand U18512 (N_18512,N_18159,N_18282);
or U18513 (N_18513,N_18315,N_18021);
nor U18514 (N_18514,N_18325,N_18238);
or U18515 (N_18515,N_18236,N_18245);
nor U18516 (N_18516,N_18305,N_18316);
and U18517 (N_18517,N_18147,N_18456);
and U18518 (N_18518,N_18426,N_18001);
and U18519 (N_18519,N_18425,N_18149);
xnor U18520 (N_18520,N_18078,N_18358);
and U18521 (N_18521,N_18215,N_18232);
and U18522 (N_18522,N_18383,N_18076);
xor U18523 (N_18523,N_18034,N_18234);
or U18524 (N_18524,N_18349,N_18223);
xor U18525 (N_18525,N_18242,N_18435);
nand U18526 (N_18526,N_18491,N_18303);
or U18527 (N_18527,N_18109,N_18407);
nand U18528 (N_18528,N_18276,N_18472);
or U18529 (N_18529,N_18098,N_18219);
nand U18530 (N_18530,N_18196,N_18350);
and U18531 (N_18531,N_18007,N_18366);
or U18532 (N_18532,N_18018,N_18211);
xnor U18533 (N_18533,N_18281,N_18356);
xor U18534 (N_18534,N_18233,N_18489);
or U18535 (N_18535,N_18307,N_18048);
and U18536 (N_18536,N_18169,N_18106);
nand U18537 (N_18537,N_18037,N_18227);
xor U18538 (N_18538,N_18360,N_18450);
nor U18539 (N_18539,N_18440,N_18474);
xnor U18540 (N_18540,N_18056,N_18042);
and U18541 (N_18541,N_18168,N_18362);
or U18542 (N_18542,N_18051,N_18403);
nand U18543 (N_18543,N_18071,N_18104);
nand U18544 (N_18544,N_18398,N_18086);
nand U18545 (N_18545,N_18128,N_18191);
nand U18546 (N_18546,N_18326,N_18493);
nand U18547 (N_18547,N_18045,N_18420);
nand U18548 (N_18548,N_18402,N_18218);
or U18549 (N_18549,N_18213,N_18016);
nor U18550 (N_18550,N_18170,N_18421);
or U18551 (N_18551,N_18391,N_18005);
or U18552 (N_18552,N_18330,N_18301);
or U18553 (N_18553,N_18067,N_18473);
xnor U18554 (N_18554,N_18388,N_18295);
xor U18555 (N_18555,N_18417,N_18247);
nand U18556 (N_18556,N_18033,N_18460);
or U18557 (N_18557,N_18436,N_18404);
or U18558 (N_18558,N_18284,N_18271);
or U18559 (N_18559,N_18338,N_18201);
or U18560 (N_18560,N_18431,N_18449);
or U18561 (N_18561,N_18451,N_18343);
xor U18562 (N_18562,N_18100,N_18323);
and U18563 (N_18563,N_18013,N_18454);
nand U18564 (N_18564,N_18142,N_18453);
and U18565 (N_18565,N_18126,N_18118);
xor U18566 (N_18566,N_18277,N_18495);
and U18567 (N_18567,N_18455,N_18114);
nor U18568 (N_18568,N_18162,N_18110);
nor U18569 (N_18569,N_18442,N_18397);
nor U18570 (N_18570,N_18441,N_18035);
xor U18571 (N_18571,N_18310,N_18029);
and U18572 (N_18572,N_18023,N_18116);
nand U18573 (N_18573,N_18380,N_18304);
or U18574 (N_18574,N_18199,N_18422);
nor U18575 (N_18575,N_18193,N_18494);
or U18576 (N_18576,N_18146,N_18187);
nand U18577 (N_18577,N_18317,N_18097);
nand U18578 (N_18578,N_18123,N_18387);
nor U18579 (N_18579,N_18476,N_18393);
nor U18580 (N_18580,N_18471,N_18153);
nand U18581 (N_18581,N_18363,N_18220);
nor U18582 (N_18582,N_18480,N_18073);
nor U18583 (N_18583,N_18179,N_18024);
nand U18584 (N_18584,N_18143,N_18302);
and U18585 (N_18585,N_18216,N_18306);
or U18586 (N_18586,N_18423,N_18337);
xor U18587 (N_18587,N_18102,N_18158);
nand U18588 (N_18588,N_18228,N_18198);
and U18589 (N_18589,N_18414,N_18053);
nand U18590 (N_18590,N_18250,N_18127);
nand U18591 (N_18591,N_18009,N_18478);
nand U18592 (N_18592,N_18214,N_18135);
nand U18593 (N_18593,N_18463,N_18099);
nor U18594 (N_18594,N_18115,N_18186);
and U18595 (N_18595,N_18049,N_18208);
and U18596 (N_18596,N_18176,N_18438);
or U18597 (N_18597,N_18195,N_18265);
or U18598 (N_18598,N_18167,N_18210);
or U18599 (N_18599,N_18339,N_18020);
nor U18600 (N_18600,N_18376,N_18047);
nor U18601 (N_18601,N_18130,N_18486);
nand U18602 (N_18602,N_18446,N_18212);
and U18603 (N_18603,N_18032,N_18031);
xnor U18604 (N_18604,N_18027,N_18178);
or U18605 (N_18605,N_18419,N_18381);
nand U18606 (N_18606,N_18103,N_18010);
nand U18607 (N_18607,N_18248,N_18386);
nand U18608 (N_18608,N_18239,N_18164);
xor U18609 (N_18609,N_18481,N_18006);
nor U18610 (N_18610,N_18240,N_18293);
or U18611 (N_18611,N_18299,N_18092);
xnor U18612 (N_18612,N_18160,N_18144);
or U18613 (N_18613,N_18230,N_18095);
nor U18614 (N_18614,N_18319,N_18372);
nand U18615 (N_18615,N_18496,N_18352);
nand U18616 (N_18616,N_18415,N_18241);
xnor U18617 (N_18617,N_18036,N_18263);
xnor U18618 (N_18618,N_18445,N_18184);
or U18619 (N_18619,N_18452,N_18467);
nand U18620 (N_18620,N_18043,N_18175);
nand U18621 (N_18621,N_18336,N_18185);
xor U18622 (N_18622,N_18261,N_18040);
xnor U18623 (N_18623,N_18427,N_18041);
xnor U18624 (N_18624,N_18353,N_18133);
or U18625 (N_18625,N_18030,N_18163);
or U18626 (N_18626,N_18072,N_18087);
or U18627 (N_18627,N_18059,N_18348);
xnor U18628 (N_18628,N_18485,N_18140);
nand U18629 (N_18629,N_18151,N_18061);
and U18630 (N_18630,N_18361,N_18054);
and U18631 (N_18631,N_18457,N_18229);
nand U18632 (N_18632,N_18434,N_18409);
nand U18633 (N_18633,N_18161,N_18283);
nand U18634 (N_18634,N_18082,N_18292);
nor U18635 (N_18635,N_18131,N_18318);
nand U18636 (N_18636,N_18401,N_18329);
xnor U18637 (N_18637,N_18406,N_18145);
nor U18638 (N_18638,N_18433,N_18468);
or U18639 (N_18639,N_18039,N_18134);
nand U18640 (N_18640,N_18136,N_18389);
nor U18641 (N_18641,N_18447,N_18462);
or U18642 (N_18642,N_18272,N_18038);
nor U18643 (N_18643,N_18477,N_18412);
or U18644 (N_18644,N_18080,N_18017);
xnor U18645 (N_18645,N_18152,N_18296);
nand U18646 (N_18646,N_18313,N_18287);
xnor U18647 (N_18647,N_18254,N_18458);
or U18648 (N_18648,N_18188,N_18429);
xnor U18649 (N_18649,N_18111,N_18112);
nor U18650 (N_18650,N_18249,N_18081);
or U18651 (N_18651,N_18000,N_18091);
nor U18652 (N_18652,N_18200,N_18331);
and U18653 (N_18653,N_18079,N_18224);
nor U18654 (N_18654,N_18088,N_18235);
xor U18655 (N_18655,N_18492,N_18324);
or U18656 (N_18656,N_18157,N_18014);
xor U18657 (N_18657,N_18390,N_18257);
and U18658 (N_18658,N_18139,N_18259);
xor U18659 (N_18659,N_18221,N_18411);
and U18660 (N_18660,N_18165,N_18244);
nor U18661 (N_18661,N_18192,N_18385);
xor U18662 (N_18662,N_18278,N_18066);
and U18663 (N_18663,N_18328,N_18205);
xor U18664 (N_18664,N_18430,N_18279);
nor U18665 (N_18665,N_18084,N_18222);
and U18666 (N_18666,N_18268,N_18085);
and U18667 (N_18667,N_18096,N_18231);
and U18668 (N_18668,N_18365,N_18068);
nor U18669 (N_18669,N_18137,N_18264);
nor U18670 (N_18670,N_18347,N_18487);
nand U18671 (N_18671,N_18197,N_18322);
or U18672 (N_18672,N_18369,N_18344);
or U18673 (N_18673,N_18443,N_18416);
nor U18674 (N_18674,N_18439,N_18378);
xnor U18675 (N_18675,N_18357,N_18174);
or U18676 (N_18676,N_18470,N_18173);
nand U18677 (N_18677,N_18243,N_18124);
nand U18678 (N_18678,N_18129,N_18117);
or U18679 (N_18679,N_18267,N_18364);
nand U18680 (N_18680,N_18141,N_18015);
and U18681 (N_18681,N_18055,N_18274);
and U18682 (N_18682,N_18022,N_18497);
nand U18683 (N_18683,N_18204,N_18070);
and U18684 (N_18684,N_18050,N_18107);
xor U18685 (N_18685,N_18448,N_18340);
and U18686 (N_18686,N_18294,N_18028);
or U18687 (N_18687,N_18237,N_18252);
or U18688 (N_18688,N_18428,N_18101);
nor U18689 (N_18689,N_18413,N_18209);
or U18690 (N_18690,N_18119,N_18342);
xnor U18691 (N_18691,N_18154,N_18260);
nor U18692 (N_18692,N_18311,N_18399);
nand U18693 (N_18693,N_18125,N_18408);
xnor U18694 (N_18694,N_18190,N_18090);
or U18695 (N_18695,N_18002,N_18172);
xor U18696 (N_18696,N_18359,N_18004);
nand U18697 (N_18697,N_18203,N_18488);
nand U18698 (N_18698,N_18113,N_18255);
nand U18699 (N_18699,N_18308,N_18121);
nor U18700 (N_18700,N_18156,N_18370);
nor U18701 (N_18701,N_18466,N_18309);
xnor U18702 (N_18702,N_18171,N_18289);
nand U18703 (N_18703,N_18183,N_18418);
nand U18704 (N_18704,N_18335,N_18075);
nand U18705 (N_18705,N_18064,N_18266);
or U18706 (N_18706,N_18194,N_18345);
nand U18707 (N_18707,N_18189,N_18483);
xor U18708 (N_18708,N_18074,N_18333);
xor U18709 (N_18709,N_18063,N_18246);
or U18710 (N_18710,N_18346,N_18132);
nor U18711 (N_18711,N_18206,N_18226);
xnor U18712 (N_18712,N_18332,N_18498);
xnor U18713 (N_18713,N_18225,N_18251);
nor U18714 (N_18714,N_18093,N_18046);
nand U18715 (N_18715,N_18298,N_18150);
nand U18716 (N_18716,N_18475,N_18288);
or U18717 (N_18717,N_18437,N_18382);
or U18718 (N_18718,N_18320,N_18469);
xor U18719 (N_18719,N_18285,N_18351);
xnor U18720 (N_18720,N_18482,N_18148);
xnor U18721 (N_18721,N_18069,N_18182);
nor U18722 (N_18722,N_18166,N_18394);
and U18723 (N_18723,N_18180,N_18155);
and U18724 (N_18724,N_18367,N_18060);
xor U18725 (N_18725,N_18253,N_18262);
or U18726 (N_18726,N_18019,N_18058);
nand U18727 (N_18727,N_18384,N_18044);
nand U18728 (N_18728,N_18392,N_18052);
nor U18729 (N_18729,N_18484,N_18432);
or U18730 (N_18730,N_18089,N_18461);
nor U18731 (N_18731,N_18105,N_18490);
nand U18732 (N_18732,N_18290,N_18400);
nor U18733 (N_18733,N_18273,N_18300);
and U18734 (N_18734,N_18120,N_18181);
or U18735 (N_18735,N_18286,N_18327);
or U18736 (N_18736,N_18025,N_18077);
and U18737 (N_18737,N_18297,N_18321);
and U18738 (N_18738,N_18280,N_18373);
nand U18739 (N_18739,N_18314,N_18396);
xnor U18740 (N_18740,N_18444,N_18499);
xnor U18741 (N_18741,N_18374,N_18395);
xor U18742 (N_18742,N_18464,N_18377);
nor U18743 (N_18743,N_18291,N_18094);
nor U18744 (N_18744,N_18479,N_18465);
xor U18745 (N_18745,N_18375,N_18207);
or U18746 (N_18746,N_18217,N_18122);
nand U18747 (N_18747,N_18083,N_18256);
nand U18748 (N_18748,N_18008,N_18341);
and U18749 (N_18749,N_18270,N_18258);
nand U18750 (N_18750,N_18244,N_18297);
xnor U18751 (N_18751,N_18344,N_18096);
nor U18752 (N_18752,N_18282,N_18328);
nor U18753 (N_18753,N_18397,N_18287);
nor U18754 (N_18754,N_18163,N_18476);
and U18755 (N_18755,N_18048,N_18273);
nor U18756 (N_18756,N_18339,N_18363);
and U18757 (N_18757,N_18114,N_18269);
xor U18758 (N_18758,N_18177,N_18329);
or U18759 (N_18759,N_18369,N_18443);
and U18760 (N_18760,N_18443,N_18144);
xor U18761 (N_18761,N_18168,N_18101);
nor U18762 (N_18762,N_18101,N_18376);
nand U18763 (N_18763,N_18213,N_18397);
nand U18764 (N_18764,N_18329,N_18496);
xor U18765 (N_18765,N_18452,N_18304);
nand U18766 (N_18766,N_18115,N_18024);
and U18767 (N_18767,N_18062,N_18258);
xor U18768 (N_18768,N_18496,N_18361);
and U18769 (N_18769,N_18378,N_18239);
and U18770 (N_18770,N_18420,N_18098);
and U18771 (N_18771,N_18496,N_18055);
nor U18772 (N_18772,N_18123,N_18396);
nor U18773 (N_18773,N_18060,N_18191);
nor U18774 (N_18774,N_18380,N_18475);
and U18775 (N_18775,N_18248,N_18327);
nand U18776 (N_18776,N_18060,N_18265);
nand U18777 (N_18777,N_18233,N_18134);
or U18778 (N_18778,N_18358,N_18222);
xor U18779 (N_18779,N_18027,N_18244);
nand U18780 (N_18780,N_18034,N_18216);
or U18781 (N_18781,N_18177,N_18233);
xnor U18782 (N_18782,N_18098,N_18036);
nor U18783 (N_18783,N_18186,N_18100);
xnor U18784 (N_18784,N_18142,N_18465);
xnor U18785 (N_18785,N_18444,N_18072);
and U18786 (N_18786,N_18014,N_18123);
or U18787 (N_18787,N_18202,N_18408);
and U18788 (N_18788,N_18167,N_18292);
and U18789 (N_18789,N_18253,N_18081);
nor U18790 (N_18790,N_18365,N_18131);
and U18791 (N_18791,N_18454,N_18241);
and U18792 (N_18792,N_18261,N_18140);
or U18793 (N_18793,N_18000,N_18186);
nor U18794 (N_18794,N_18324,N_18441);
or U18795 (N_18795,N_18163,N_18058);
xnor U18796 (N_18796,N_18418,N_18200);
or U18797 (N_18797,N_18099,N_18092);
xor U18798 (N_18798,N_18481,N_18139);
nor U18799 (N_18799,N_18287,N_18189);
xor U18800 (N_18800,N_18080,N_18092);
or U18801 (N_18801,N_18108,N_18173);
nor U18802 (N_18802,N_18450,N_18106);
nand U18803 (N_18803,N_18378,N_18312);
nand U18804 (N_18804,N_18031,N_18244);
xor U18805 (N_18805,N_18130,N_18355);
xnor U18806 (N_18806,N_18058,N_18251);
nor U18807 (N_18807,N_18378,N_18277);
and U18808 (N_18808,N_18064,N_18159);
xnor U18809 (N_18809,N_18066,N_18217);
nor U18810 (N_18810,N_18317,N_18189);
nand U18811 (N_18811,N_18439,N_18426);
nor U18812 (N_18812,N_18185,N_18127);
or U18813 (N_18813,N_18182,N_18400);
xor U18814 (N_18814,N_18017,N_18024);
xnor U18815 (N_18815,N_18119,N_18472);
nand U18816 (N_18816,N_18096,N_18131);
nor U18817 (N_18817,N_18199,N_18184);
nand U18818 (N_18818,N_18108,N_18211);
nor U18819 (N_18819,N_18128,N_18475);
nand U18820 (N_18820,N_18236,N_18027);
nor U18821 (N_18821,N_18088,N_18257);
nor U18822 (N_18822,N_18288,N_18067);
nand U18823 (N_18823,N_18138,N_18302);
nor U18824 (N_18824,N_18487,N_18084);
xnor U18825 (N_18825,N_18082,N_18153);
xor U18826 (N_18826,N_18228,N_18231);
and U18827 (N_18827,N_18462,N_18263);
xnor U18828 (N_18828,N_18416,N_18159);
and U18829 (N_18829,N_18490,N_18018);
nor U18830 (N_18830,N_18093,N_18261);
or U18831 (N_18831,N_18055,N_18227);
or U18832 (N_18832,N_18186,N_18472);
or U18833 (N_18833,N_18446,N_18296);
or U18834 (N_18834,N_18374,N_18323);
xnor U18835 (N_18835,N_18191,N_18228);
nand U18836 (N_18836,N_18326,N_18172);
nand U18837 (N_18837,N_18410,N_18039);
xor U18838 (N_18838,N_18088,N_18037);
or U18839 (N_18839,N_18281,N_18344);
and U18840 (N_18840,N_18249,N_18063);
or U18841 (N_18841,N_18019,N_18487);
or U18842 (N_18842,N_18337,N_18201);
nand U18843 (N_18843,N_18280,N_18152);
nor U18844 (N_18844,N_18420,N_18397);
nor U18845 (N_18845,N_18464,N_18091);
nor U18846 (N_18846,N_18359,N_18284);
nor U18847 (N_18847,N_18193,N_18177);
or U18848 (N_18848,N_18291,N_18120);
nor U18849 (N_18849,N_18158,N_18060);
nand U18850 (N_18850,N_18055,N_18359);
nand U18851 (N_18851,N_18349,N_18177);
nor U18852 (N_18852,N_18186,N_18232);
nand U18853 (N_18853,N_18240,N_18472);
and U18854 (N_18854,N_18481,N_18364);
nand U18855 (N_18855,N_18182,N_18283);
xor U18856 (N_18856,N_18118,N_18197);
xor U18857 (N_18857,N_18378,N_18127);
nor U18858 (N_18858,N_18280,N_18270);
and U18859 (N_18859,N_18383,N_18121);
nor U18860 (N_18860,N_18113,N_18171);
nor U18861 (N_18861,N_18343,N_18071);
or U18862 (N_18862,N_18278,N_18275);
nor U18863 (N_18863,N_18129,N_18280);
or U18864 (N_18864,N_18059,N_18172);
xor U18865 (N_18865,N_18245,N_18206);
xor U18866 (N_18866,N_18375,N_18116);
or U18867 (N_18867,N_18144,N_18363);
or U18868 (N_18868,N_18255,N_18164);
and U18869 (N_18869,N_18012,N_18115);
nor U18870 (N_18870,N_18240,N_18411);
and U18871 (N_18871,N_18461,N_18098);
and U18872 (N_18872,N_18320,N_18353);
xnor U18873 (N_18873,N_18448,N_18337);
nor U18874 (N_18874,N_18106,N_18372);
and U18875 (N_18875,N_18345,N_18105);
or U18876 (N_18876,N_18052,N_18061);
and U18877 (N_18877,N_18379,N_18176);
or U18878 (N_18878,N_18319,N_18153);
nand U18879 (N_18879,N_18116,N_18340);
nand U18880 (N_18880,N_18398,N_18221);
nor U18881 (N_18881,N_18121,N_18355);
nand U18882 (N_18882,N_18444,N_18378);
or U18883 (N_18883,N_18223,N_18286);
or U18884 (N_18884,N_18149,N_18110);
xnor U18885 (N_18885,N_18210,N_18244);
and U18886 (N_18886,N_18319,N_18488);
nand U18887 (N_18887,N_18423,N_18468);
or U18888 (N_18888,N_18247,N_18285);
or U18889 (N_18889,N_18350,N_18081);
nor U18890 (N_18890,N_18201,N_18085);
nand U18891 (N_18891,N_18093,N_18058);
nor U18892 (N_18892,N_18312,N_18283);
or U18893 (N_18893,N_18019,N_18497);
nor U18894 (N_18894,N_18224,N_18390);
or U18895 (N_18895,N_18380,N_18057);
or U18896 (N_18896,N_18098,N_18033);
nand U18897 (N_18897,N_18199,N_18064);
nor U18898 (N_18898,N_18219,N_18484);
xor U18899 (N_18899,N_18245,N_18317);
or U18900 (N_18900,N_18138,N_18464);
xnor U18901 (N_18901,N_18454,N_18239);
nor U18902 (N_18902,N_18365,N_18105);
and U18903 (N_18903,N_18326,N_18485);
and U18904 (N_18904,N_18362,N_18364);
xor U18905 (N_18905,N_18042,N_18114);
xnor U18906 (N_18906,N_18094,N_18319);
nand U18907 (N_18907,N_18239,N_18273);
nor U18908 (N_18908,N_18485,N_18099);
xnor U18909 (N_18909,N_18473,N_18289);
xor U18910 (N_18910,N_18191,N_18382);
nand U18911 (N_18911,N_18394,N_18430);
or U18912 (N_18912,N_18326,N_18475);
xor U18913 (N_18913,N_18258,N_18321);
and U18914 (N_18914,N_18251,N_18437);
xor U18915 (N_18915,N_18062,N_18450);
or U18916 (N_18916,N_18051,N_18217);
and U18917 (N_18917,N_18427,N_18377);
nor U18918 (N_18918,N_18173,N_18352);
nand U18919 (N_18919,N_18049,N_18465);
nor U18920 (N_18920,N_18143,N_18482);
nor U18921 (N_18921,N_18182,N_18001);
and U18922 (N_18922,N_18444,N_18256);
or U18923 (N_18923,N_18447,N_18494);
nand U18924 (N_18924,N_18007,N_18209);
nand U18925 (N_18925,N_18339,N_18414);
nand U18926 (N_18926,N_18477,N_18168);
xnor U18927 (N_18927,N_18473,N_18171);
xnor U18928 (N_18928,N_18455,N_18089);
nor U18929 (N_18929,N_18130,N_18187);
nand U18930 (N_18930,N_18280,N_18475);
xor U18931 (N_18931,N_18205,N_18303);
nor U18932 (N_18932,N_18207,N_18211);
xnor U18933 (N_18933,N_18119,N_18393);
and U18934 (N_18934,N_18097,N_18022);
nand U18935 (N_18935,N_18074,N_18095);
nand U18936 (N_18936,N_18143,N_18343);
nor U18937 (N_18937,N_18014,N_18344);
and U18938 (N_18938,N_18181,N_18294);
xnor U18939 (N_18939,N_18115,N_18215);
and U18940 (N_18940,N_18248,N_18291);
xor U18941 (N_18941,N_18468,N_18255);
nand U18942 (N_18942,N_18398,N_18460);
and U18943 (N_18943,N_18022,N_18194);
nand U18944 (N_18944,N_18347,N_18209);
and U18945 (N_18945,N_18075,N_18236);
or U18946 (N_18946,N_18070,N_18071);
xnor U18947 (N_18947,N_18210,N_18259);
nand U18948 (N_18948,N_18037,N_18166);
nand U18949 (N_18949,N_18181,N_18076);
nand U18950 (N_18950,N_18024,N_18355);
and U18951 (N_18951,N_18376,N_18442);
nand U18952 (N_18952,N_18482,N_18209);
nand U18953 (N_18953,N_18245,N_18011);
or U18954 (N_18954,N_18018,N_18338);
nand U18955 (N_18955,N_18214,N_18454);
nor U18956 (N_18956,N_18398,N_18294);
and U18957 (N_18957,N_18028,N_18431);
xor U18958 (N_18958,N_18494,N_18468);
and U18959 (N_18959,N_18172,N_18067);
nor U18960 (N_18960,N_18039,N_18278);
xnor U18961 (N_18961,N_18144,N_18439);
and U18962 (N_18962,N_18453,N_18410);
or U18963 (N_18963,N_18311,N_18178);
nor U18964 (N_18964,N_18064,N_18020);
nand U18965 (N_18965,N_18019,N_18185);
xor U18966 (N_18966,N_18083,N_18299);
or U18967 (N_18967,N_18167,N_18301);
or U18968 (N_18968,N_18161,N_18369);
nor U18969 (N_18969,N_18107,N_18041);
or U18970 (N_18970,N_18417,N_18482);
nand U18971 (N_18971,N_18308,N_18362);
nand U18972 (N_18972,N_18331,N_18393);
nor U18973 (N_18973,N_18259,N_18408);
and U18974 (N_18974,N_18265,N_18128);
and U18975 (N_18975,N_18286,N_18494);
and U18976 (N_18976,N_18199,N_18168);
xnor U18977 (N_18977,N_18174,N_18390);
nor U18978 (N_18978,N_18365,N_18315);
and U18979 (N_18979,N_18116,N_18096);
and U18980 (N_18980,N_18142,N_18225);
nor U18981 (N_18981,N_18008,N_18058);
xor U18982 (N_18982,N_18237,N_18256);
nor U18983 (N_18983,N_18230,N_18152);
xnor U18984 (N_18984,N_18305,N_18231);
nor U18985 (N_18985,N_18371,N_18079);
nor U18986 (N_18986,N_18066,N_18024);
nor U18987 (N_18987,N_18242,N_18018);
and U18988 (N_18988,N_18346,N_18476);
xor U18989 (N_18989,N_18345,N_18443);
xor U18990 (N_18990,N_18237,N_18049);
nor U18991 (N_18991,N_18037,N_18473);
or U18992 (N_18992,N_18159,N_18218);
and U18993 (N_18993,N_18452,N_18329);
nand U18994 (N_18994,N_18118,N_18009);
nor U18995 (N_18995,N_18477,N_18182);
nor U18996 (N_18996,N_18398,N_18428);
or U18997 (N_18997,N_18454,N_18251);
nand U18998 (N_18998,N_18056,N_18200);
and U18999 (N_18999,N_18071,N_18206);
xnor U19000 (N_19000,N_18662,N_18528);
and U19001 (N_19001,N_18983,N_18881);
and U19002 (N_19002,N_18601,N_18993);
or U19003 (N_19003,N_18802,N_18959);
nor U19004 (N_19004,N_18512,N_18578);
xor U19005 (N_19005,N_18902,N_18692);
nand U19006 (N_19006,N_18500,N_18771);
xnor U19007 (N_19007,N_18774,N_18855);
or U19008 (N_19008,N_18981,N_18527);
xor U19009 (N_19009,N_18600,N_18519);
nor U19010 (N_19010,N_18569,N_18714);
xnor U19011 (N_19011,N_18803,N_18645);
or U19012 (N_19012,N_18675,N_18523);
and U19013 (N_19013,N_18904,N_18951);
nand U19014 (N_19014,N_18935,N_18599);
nand U19015 (N_19015,N_18788,N_18579);
and U19016 (N_19016,N_18734,N_18844);
nand U19017 (N_19017,N_18572,N_18558);
and U19018 (N_19018,N_18938,N_18680);
and U19019 (N_19019,N_18622,N_18857);
nor U19020 (N_19020,N_18638,N_18652);
nor U19021 (N_19021,N_18838,N_18962);
xor U19022 (N_19022,N_18866,N_18754);
nor U19023 (N_19023,N_18748,N_18811);
nand U19024 (N_19024,N_18603,N_18884);
xor U19025 (N_19025,N_18980,N_18909);
and U19026 (N_19026,N_18618,N_18710);
xor U19027 (N_19027,N_18963,N_18661);
and U19028 (N_19028,N_18597,N_18913);
xnor U19029 (N_19029,N_18725,N_18997);
or U19030 (N_19030,N_18534,N_18691);
nand U19031 (N_19031,N_18780,N_18713);
nand U19032 (N_19032,N_18787,N_18712);
nor U19033 (N_19033,N_18945,N_18669);
nand U19034 (N_19034,N_18860,N_18849);
xnor U19035 (N_19035,N_18593,N_18605);
nand U19036 (N_19036,N_18635,N_18695);
or U19037 (N_19037,N_18567,N_18944);
xor U19038 (N_19038,N_18954,N_18539);
and U19039 (N_19039,N_18629,N_18984);
and U19040 (N_19040,N_18611,N_18503);
nor U19041 (N_19041,N_18765,N_18960);
or U19042 (N_19042,N_18955,N_18637);
nor U19043 (N_19043,N_18843,N_18687);
nand U19044 (N_19044,N_18737,N_18782);
or U19045 (N_19045,N_18893,N_18950);
nand U19046 (N_19046,N_18856,N_18819);
or U19047 (N_19047,N_18685,N_18776);
nand U19048 (N_19048,N_18628,N_18910);
nand U19049 (N_19049,N_18553,N_18510);
nand U19050 (N_19050,N_18670,N_18831);
and U19051 (N_19051,N_18508,N_18973);
or U19052 (N_19052,N_18943,N_18870);
xnor U19053 (N_19053,N_18898,N_18990);
nand U19054 (N_19054,N_18756,N_18625);
nand U19055 (N_19055,N_18681,N_18892);
nor U19056 (N_19056,N_18786,N_18835);
xor U19057 (N_19057,N_18609,N_18650);
nand U19058 (N_19058,N_18524,N_18889);
nand U19059 (N_19059,N_18651,N_18663);
and U19060 (N_19060,N_18877,N_18975);
xnor U19061 (N_19061,N_18833,N_18672);
and U19062 (N_19062,N_18919,N_18864);
xor U19063 (N_19063,N_18850,N_18509);
and U19064 (N_19064,N_18632,N_18683);
nor U19065 (N_19065,N_18530,N_18789);
xor U19066 (N_19066,N_18667,N_18773);
and U19067 (N_19067,N_18542,N_18688);
nand U19068 (N_19068,N_18595,N_18658);
and U19069 (N_19069,N_18738,N_18747);
nor U19070 (N_19070,N_18920,N_18521);
nand U19071 (N_19071,N_18607,N_18654);
and U19072 (N_19072,N_18940,N_18809);
xor U19073 (N_19073,N_18548,N_18694);
nand U19074 (N_19074,N_18656,N_18813);
or U19075 (N_19075,N_18999,N_18582);
and U19076 (N_19076,N_18676,N_18770);
or U19077 (N_19077,N_18964,N_18757);
or U19078 (N_19078,N_18633,N_18987);
xnor U19079 (N_19079,N_18924,N_18852);
xor U19080 (N_19080,N_18794,N_18772);
nand U19081 (N_19081,N_18804,N_18549);
nand U19082 (N_19082,N_18736,N_18532);
nor U19083 (N_19083,N_18862,N_18921);
and U19084 (N_19084,N_18859,N_18846);
or U19085 (N_19085,N_18965,N_18653);
or U19086 (N_19086,N_18867,N_18798);
nor U19087 (N_19087,N_18896,N_18942);
and U19088 (N_19088,N_18674,N_18907);
or U19089 (N_19089,N_18887,N_18808);
nand U19090 (N_19090,N_18777,N_18931);
nor U19091 (N_19091,N_18761,N_18568);
and U19092 (N_19092,N_18668,N_18948);
and U19093 (N_19093,N_18636,N_18589);
xnor U19094 (N_19094,N_18778,N_18576);
xnor U19095 (N_19095,N_18923,N_18711);
nand U19096 (N_19096,N_18995,N_18801);
nand U19097 (N_19097,N_18810,N_18785);
or U19098 (N_19098,N_18513,N_18586);
or U19099 (N_19099,N_18511,N_18957);
and U19100 (N_19100,N_18630,N_18643);
nand U19101 (N_19101,N_18851,N_18516);
nand U19102 (N_19102,N_18739,N_18895);
xor U19103 (N_19103,N_18974,N_18565);
and U19104 (N_19104,N_18551,N_18735);
or U19105 (N_19105,N_18580,N_18925);
and U19106 (N_19106,N_18918,N_18886);
nand U19107 (N_19107,N_18613,N_18868);
nor U19108 (N_19108,N_18875,N_18564);
and U19109 (N_19109,N_18936,N_18905);
xor U19110 (N_19110,N_18665,N_18836);
xor U19111 (N_19111,N_18543,N_18614);
and U19112 (N_19112,N_18552,N_18561);
or U19113 (N_19113,N_18894,N_18827);
and U19114 (N_19114,N_18679,N_18820);
or U19115 (N_19115,N_18563,N_18514);
nor U19116 (N_19116,N_18590,N_18571);
xor U19117 (N_19117,N_18506,N_18546);
nand U19118 (N_19118,N_18750,N_18556);
or U19119 (N_19119,N_18817,N_18649);
nand U19120 (N_19120,N_18847,N_18930);
nor U19121 (N_19121,N_18715,N_18766);
nor U19122 (N_19122,N_18823,N_18644);
or U19123 (N_19123,N_18807,N_18744);
or U19124 (N_19124,N_18915,N_18879);
nand U19125 (N_19125,N_18555,N_18709);
and U19126 (N_19126,N_18826,N_18861);
or U19127 (N_19127,N_18928,N_18912);
xor U19128 (N_19128,N_18966,N_18818);
and U19129 (N_19129,N_18719,N_18805);
xor U19130 (N_19130,N_18626,N_18627);
nor U19131 (N_19131,N_18976,N_18538);
or U19132 (N_19132,N_18704,N_18972);
nand U19133 (N_19133,N_18793,N_18620);
or U19134 (N_19134,N_18869,N_18806);
and U19135 (N_19135,N_18906,N_18970);
xnor U19136 (N_19136,N_18927,N_18608);
xor U19137 (N_19137,N_18730,N_18594);
nor U19138 (N_19138,N_18746,N_18723);
xnor U19139 (N_19139,N_18876,N_18791);
and U19140 (N_19140,N_18502,N_18520);
nor U19141 (N_19141,N_18588,N_18979);
nand U19142 (N_19142,N_18677,N_18795);
xor U19143 (N_19143,N_18751,N_18941);
nor U19144 (N_19144,N_18504,N_18678);
xnor U19145 (N_19145,N_18557,N_18853);
or U19146 (N_19146,N_18947,N_18891);
xnor U19147 (N_19147,N_18996,N_18764);
and U19148 (N_19148,N_18880,N_18647);
and U19149 (N_19149,N_18562,N_18937);
nand U19150 (N_19150,N_18900,N_18529);
xor U19151 (N_19151,N_18830,N_18958);
or U19152 (N_19152,N_18897,N_18854);
nor U19153 (N_19153,N_18540,N_18671);
or U19154 (N_19154,N_18624,N_18535);
and U19155 (N_19155,N_18575,N_18716);
xor U19156 (N_19156,N_18584,N_18901);
or U19157 (N_19157,N_18544,N_18812);
xor U19158 (N_19158,N_18890,N_18655);
nand U19159 (N_19159,N_18641,N_18648);
nor U19160 (N_19160,N_18956,N_18606);
nand U19161 (N_19161,N_18952,N_18926);
xor U19162 (N_19162,N_18961,N_18690);
and U19163 (N_19163,N_18517,N_18783);
or U19164 (N_19164,N_18696,N_18932);
nand U19165 (N_19165,N_18845,N_18899);
or U19166 (N_19166,N_18825,N_18969);
and U19167 (N_19167,N_18610,N_18616);
and U19168 (N_19168,N_18721,N_18664);
or U19169 (N_19169,N_18612,N_18934);
or U19170 (N_19170,N_18699,N_18989);
xor U19171 (N_19171,N_18848,N_18740);
xor U19172 (N_19172,N_18752,N_18684);
or U19173 (N_19173,N_18686,N_18749);
xnor U19174 (N_19174,N_18768,N_18968);
and U19175 (N_19175,N_18871,N_18917);
and U19176 (N_19176,N_18505,N_18596);
or U19177 (N_19177,N_18903,N_18779);
xnor U19178 (N_19178,N_18767,N_18797);
nand U19179 (N_19179,N_18731,N_18729);
and U19180 (N_19180,N_18554,N_18988);
or U19181 (N_19181,N_18873,N_18537);
or U19182 (N_19182,N_18982,N_18971);
nor U19183 (N_19183,N_18559,N_18623);
xor U19184 (N_19184,N_18939,N_18728);
nor U19185 (N_19185,N_18732,N_18911);
nand U19186 (N_19186,N_18619,N_18781);
nand U19187 (N_19187,N_18742,N_18800);
xor U19188 (N_19188,N_18745,N_18703);
xnor U19189 (N_19189,N_18587,N_18615);
nor U19190 (N_19190,N_18883,N_18790);
nand U19191 (N_19191,N_18642,N_18837);
and U19192 (N_19192,N_18560,N_18824);
nor U19193 (N_19193,N_18829,N_18840);
or U19194 (N_19194,N_18998,N_18828);
nor U19195 (N_19195,N_18698,N_18531);
and U19196 (N_19196,N_18885,N_18585);
or U19197 (N_19197,N_18657,N_18753);
or U19198 (N_19198,N_18922,N_18727);
nand U19199 (N_19199,N_18763,N_18758);
and U19200 (N_19200,N_18700,N_18659);
xnor U19201 (N_19201,N_18536,N_18547);
nor U19202 (N_19202,N_18566,N_18697);
nor U19203 (N_19203,N_18796,N_18929);
nor U19204 (N_19204,N_18977,N_18741);
xnor U19205 (N_19205,N_18762,N_18839);
xor U19206 (N_19206,N_18515,N_18946);
or U19207 (N_19207,N_18631,N_18722);
and U19208 (N_19208,N_18573,N_18522);
nand U19209 (N_19209,N_18832,N_18707);
and U19210 (N_19210,N_18646,N_18816);
xnor U19211 (N_19211,N_18878,N_18933);
nor U19212 (N_19212,N_18822,N_18545);
or U19213 (N_19213,N_18660,N_18874);
and U19214 (N_19214,N_18792,N_18991);
nor U19215 (N_19215,N_18705,N_18949);
nor U19216 (N_19216,N_18759,N_18604);
and U19217 (N_19217,N_18914,N_18865);
nor U19218 (N_19218,N_18863,N_18550);
nand U19219 (N_19219,N_18621,N_18743);
nand U19220 (N_19220,N_18821,N_18994);
nand U19221 (N_19221,N_18592,N_18639);
xnor U19222 (N_19222,N_18888,N_18717);
nand U19223 (N_19223,N_18755,N_18689);
nand U19224 (N_19224,N_18872,N_18581);
nor U19225 (N_19225,N_18673,N_18916);
nor U19226 (N_19226,N_18583,N_18602);
nand U19227 (N_19227,N_18775,N_18682);
nand U19228 (N_19228,N_18726,N_18702);
or U19229 (N_19229,N_18708,N_18953);
or U19230 (N_19230,N_18598,N_18858);
or U19231 (N_19231,N_18978,N_18501);
or U19232 (N_19232,N_18799,N_18986);
or U19233 (N_19233,N_18815,N_18507);
and U19234 (N_19234,N_18574,N_18541);
nand U19235 (N_19235,N_18617,N_18814);
nand U19236 (N_19236,N_18733,N_18701);
or U19237 (N_19237,N_18992,N_18518);
nor U19238 (N_19238,N_18842,N_18718);
or U19239 (N_19239,N_18640,N_18570);
and U19240 (N_19240,N_18985,N_18526);
or U19241 (N_19241,N_18882,N_18533);
nor U19242 (N_19242,N_18769,N_18784);
nor U19243 (N_19243,N_18908,N_18666);
nand U19244 (N_19244,N_18841,N_18834);
nand U19245 (N_19245,N_18591,N_18760);
and U19246 (N_19246,N_18634,N_18693);
and U19247 (N_19247,N_18577,N_18706);
and U19248 (N_19248,N_18724,N_18720);
nand U19249 (N_19249,N_18967,N_18525);
nor U19250 (N_19250,N_18830,N_18747);
nor U19251 (N_19251,N_18921,N_18619);
nor U19252 (N_19252,N_18809,N_18622);
xor U19253 (N_19253,N_18843,N_18972);
or U19254 (N_19254,N_18786,N_18940);
nand U19255 (N_19255,N_18703,N_18641);
xor U19256 (N_19256,N_18876,N_18964);
xnor U19257 (N_19257,N_18629,N_18639);
nand U19258 (N_19258,N_18688,N_18928);
and U19259 (N_19259,N_18700,N_18972);
nand U19260 (N_19260,N_18807,N_18974);
nor U19261 (N_19261,N_18976,N_18586);
or U19262 (N_19262,N_18688,N_18908);
and U19263 (N_19263,N_18994,N_18555);
nand U19264 (N_19264,N_18797,N_18701);
xor U19265 (N_19265,N_18612,N_18517);
nand U19266 (N_19266,N_18686,N_18890);
nand U19267 (N_19267,N_18626,N_18860);
xor U19268 (N_19268,N_18697,N_18968);
nand U19269 (N_19269,N_18806,N_18996);
xor U19270 (N_19270,N_18822,N_18860);
xnor U19271 (N_19271,N_18756,N_18673);
and U19272 (N_19272,N_18962,N_18812);
nand U19273 (N_19273,N_18982,N_18666);
or U19274 (N_19274,N_18602,N_18563);
and U19275 (N_19275,N_18598,N_18760);
nand U19276 (N_19276,N_18900,N_18754);
and U19277 (N_19277,N_18736,N_18661);
nand U19278 (N_19278,N_18835,N_18850);
nor U19279 (N_19279,N_18692,N_18612);
xnor U19280 (N_19280,N_18541,N_18898);
nor U19281 (N_19281,N_18820,N_18600);
or U19282 (N_19282,N_18901,N_18551);
and U19283 (N_19283,N_18635,N_18609);
and U19284 (N_19284,N_18716,N_18888);
or U19285 (N_19285,N_18989,N_18626);
and U19286 (N_19286,N_18910,N_18720);
nand U19287 (N_19287,N_18731,N_18984);
nand U19288 (N_19288,N_18549,N_18730);
xor U19289 (N_19289,N_18920,N_18782);
xor U19290 (N_19290,N_18654,N_18813);
xnor U19291 (N_19291,N_18999,N_18912);
nor U19292 (N_19292,N_18824,N_18553);
nor U19293 (N_19293,N_18527,N_18984);
nand U19294 (N_19294,N_18799,N_18937);
xnor U19295 (N_19295,N_18649,N_18975);
nor U19296 (N_19296,N_18822,N_18511);
and U19297 (N_19297,N_18876,N_18883);
and U19298 (N_19298,N_18698,N_18992);
nor U19299 (N_19299,N_18518,N_18933);
xnor U19300 (N_19300,N_18802,N_18929);
nor U19301 (N_19301,N_18784,N_18966);
nor U19302 (N_19302,N_18542,N_18839);
xor U19303 (N_19303,N_18987,N_18760);
nor U19304 (N_19304,N_18988,N_18934);
xnor U19305 (N_19305,N_18694,N_18904);
and U19306 (N_19306,N_18986,N_18873);
nor U19307 (N_19307,N_18681,N_18571);
or U19308 (N_19308,N_18911,N_18812);
nor U19309 (N_19309,N_18673,N_18978);
or U19310 (N_19310,N_18996,N_18847);
or U19311 (N_19311,N_18870,N_18816);
xnor U19312 (N_19312,N_18736,N_18867);
xor U19313 (N_19313,N_18511,N_18885);
or U19314 (N_19314,N_18732,N_18596);
xor U19315 (N_19315,N_18977,N_18929);
xnor U19316 (N_19316,N_18957,N_18994);
nor U19317 (N_19317,N_18647,N_18843);
nor U19318 (N_19318,N_18920,N_18783);
xor U19319 (N_19319,N_18760,N_18988);
nor U19320 (N_19320,N_18876,N_18974);
nand U19321 (N_19321,N_18637,N_18954);
or U19322 (N_19322,N_18701,N_18644);
nor U19323 (N_19323,N_18950,N_18803);
or U19324 (N_19324,N_18691,N_18759);
nor U19325 (N_19325,N_18994,N_18786);
nand U19326 (N_19326,N_18984,N_18908);
or U19327 (N_19327,N_18968,N_18522);
nor U19328 (N_19328,N_18683,N_18913);
nor U19329 (N_19329,N_18514,N_18865);
nand U19330 (N_19330,N_18904,N_18581);
nand U19331 (N_19331,N_18927,N_18762);
nand U19332 (N_19332,N_18864,N_18719);
or U19333 (N_19333,N_18589,N_18559);
or U19334 (N_19334,N_18591,N_18892);
nor U19335 (N_19335,N_18544,N_18540);
and U19336 (N_19336,N_18794,N_18899);
xor U19337 (N_19337,N_18779,N_18535);
nand U19338 (N_19338,N_18906,N_18759);
nand U19339 (N_19339,N_18837,N_18721);
and U19340 (N_19340,N_18989,N_18972);
nor U19341 (N_19341,N_18938,N_18878);
nor U19342 (N_19342,N_18664,N_18777);
nor U19343 (N_19343,N_18761,N_18930);
or U19344 (N_19344,N_18806,N_18801);
xor U19345 (N_19345,N_18836,N_18529);
xnor U19346 (N_19346,N_18755,N_18870);
and U19347 (N_19347,N_18822,N_18864);
nand U19348 (N_19348,N_18548,N_18544);
nand U19349 (N_19349,N_18978,N_18963);
or U19350 (N_19350,N_18859,N_18970);
xnor U19351 (N_19351,N_18887,N_18758);
or U19352 (N_19352,N_18849,N_18628);
xnor U19353 (N_19353,N_18527,N_18614);
nand U19354 (N_19354,N_18807,N_18854);
xnor U19355 (N_19355,N_18634,N_18526);
or U19356 (N_19356,N_18549,N_18555);
xor U19357 (N_19357,N_18609,N_18877);
nor U19358 (N_19358,N_18802,N_18584);
nor U19359 (N_19359,N_18559,N_18859);
nand U19360 (N_19360,N_18610,N_18889);
xnor U19361 (N_19361,N_18573,N_18561);
xnor U19362 (N_19362,N_18874,N_18572);
or U19363 (N_19363,N_18524,N_18940);
nor U19364 (N_19364,N_18540,N_18733);
xor U19365 (N_19365,N_18688,N_18987);
or U19366 (N_19366,N_18929,N_18506);
or U19367 (N_19367,N_18880,N_18812);
nor U19368 (N_19368,N_18749,N_18965);
and U19369 (N_19369,N_18628,N_18957);
nor U19370 (N_19370,N_18868,N_18939);
nor U19371 (N_19371,N_18537,N_18502);
and U19372 (N_19372,N_18651,N_18763);
or U19373 (N_19373,N_18665,N_18586);
nand U19374 (N_19374,N_18922,N_18576);
xor U19375 (N_19375,N_18986,N_18975);
xor U19376 (N_19376,N_18838,N_18903);
and U19377 (N_19377,N_18948,N_18876);
nor U19378 (N_19378,N_18520,N_18825);
xnor U19379 (N_19379,N_18964,N_18910);
nor U19380 (N_19380,N_18750,N_18999);
nor U19381 (N_19381,N_18600,N_18811);
nor U19382 (N_19382,N_18753,N_18526);
xnor U19383 (N_19383,N_18649,N_18929);
or U19384 (N_19384,N_18686,N_18560);
xor U19385 (N_19385,N_18979,N_18925);
and U19386 (N_19386,N_18765,N_18512);
or U19387 (N_19387,N_18749,N_18750);
xor U19388 (N_19388,N_18769,N_18645);
and U19389 (N_19389,N_18839,N_18554);
nor U19390 (N_19390,N_18961,N_18721);
and U19391 (N_19391,N_18623,N_18640);
xnor U19392 (N_19392,N_18925,N_18830);
xor U19393 (N_19393,N_18870,N_18916);
or U19394 (N_19394,N_18884,N_18563);
nor U19395 (N_19395,N_18515,N_18797);
nand U19396 (N_19396,N_18809,N_18842);
and U19397 (N_19397,N_18855,N_18635);
nor U19398 (N_19398,N_18788,N_18653);
or U19399 (N_19399,N_18633,N_18823);
or U19400 (N_19400,N_18627,N_18937);
nand U19401 (N_19401,N_18556,N_18738);
or U19402 (N_19402,N_18815,N_18719);
xnor U19403 (N_19403,N_18832,N_18611);
or U19404 (N_19404,N_18834,N_18664);
or U19405 (N_19405,N_18620,N_18839);
nand U19406 (N_19406,N_18910,N_18584);
and U19407 (N_19407,N_18875,N_18680);
or U19408 (N_19408,N_18602,N_18936);
or U19409 (N_19409,N_18578,N_18956);
xor U19410 (N_19410,N_18707,N_18866);
and U19411 (N_19411,N_18736,N_18749);
and U19412 (N_19412,N_18605,N_18866);
nand U19413 (N_19413,N_18658,N_18932);
xnor U19414 (N_19414,N_18998,N_18708);
xnor U19415 (N_19415,N_18870,N_18812);
nor U19416 (N_19416,N_18830,N_18739);
or U19417 (N_19417,N_18801,N_18818);
xnor U19418 (N_19418,N_18927,N_18516);
and U19419 (N_19419,N_18778,N_18962);
and U19420 (N_19420,N_18824,N_18712);
or U19421 (N_19421,N_18620,N_18608);
nor U19422 (N_19422,N_18643,N_18615);
or U19423 (N_19423,N_18800,N_18754);
and U19424 (N_19424,N_18784,N_18582);
and U19425 (N_19425,N_18687,N_18637);
nor U19426 (N_19426,N_18958,N_18930);
nor U19427 (N_19427,N_18703,N_18552);
nand U19428 (N_19428,N_18714,N_18633);
xor U19429 (N_19429,N_18578,N_18545);
nand U19430 (N_19430,N_18708,N_18741);
and U19431 (N_19431,N_18696,N_18655);
and U19432 (N_19432,N_18960,N_18809);
nand U19433 (N_19433,N_18882,N_18548);
nor U19434 (N_19434,N_18685,N_18725);
and U19435 (N_19435,N_18831,N_18991);
xnor U19436 (N_19436,N_18518,N_18623);
nor U19437 (N_19437,N_18959,N_18594);
and U19438 (N_19438,N_18833,N_18574);
nand U19439 (N_19439,N_18698,N_18931);
and U19440 (N_19440,N_18761,N_18744);
or U19441 (N_19441,N_18827,N_18760);
and U19442 (N_19442,N_18797,N_18832);
or U19443 (N_19443,N_18729,N_18550);
or U19444 (N_19444,N_18798,N_18610);
xor U19445 (N_19445,N_18681,N_18931);
nand U19446 (N_19446,N_18851,N_18661);
nor U19447 (N_19447,N_18861,N_18750);
and U19448 (N_19448,N_18859,N_18508);
nor U19449 (N_19449,N_18628,N_18538);
and U19450 (N_19450,N_18996,N_18563);
xnor U19451 (N_19451,N_18748,N_18756);
and U19452 (N_19452,N_18935,N_18819);
nor U19453 (N_19453,N_18617,N_18979);
and U19454 (N_19454,N_18762,N_18964);
or U19455 (N_19455,N_18707,N_18858);
nor U19456 (N_19456,N_18864,N_18821);
xnor U19457 (N_19457,N_18908,N_18999);
nand U19458 (N_19458,N_18580,N_18559);
nor U19459 (N_19459,N_18648,N_18931);
nand U19460 (N_19460,N_18532,N_18686);
or U19461 (N_19461,N_18854,N_18534);
nand U19462 (N_19462,N_18997,N_18993);
nand U19463 (N_19463,N_18671,N_18811);
or U19464 (N_19464,N_18852,N_18936);
or U19465 (N_19465,N_18577,N_18954);
and U19466 (N_19466,N_18910,N_18875);
and U19467 (N_19467,N_18690,N_18940);
or U19468 (N_19468,N_18549,N_18573);
nor U19469 (N_19469,N_18882,N_18708);
or U19470 (N_19470,N_18516,N_18777);
xor U19471 (N_19471,N_18999,N_18886);
nor U19472 (N_19472,N_18948,N_18975);
xor U19473 (N_19473,N_18679,N_18852);
or U19474 (N_19474,N_18948,N_18657);
xnor U19475 (N_19475,N_18590,N_18814);
and U19476 (N_19476,N_18785,N_18965);
or U19477 (N_19477,N_18883,N_18540);
nor U19478 (N_19478,N_18668,N_18776);
xnor U19479 (N_19479,N_18979,N_18852);
nand U19480 (N_19480,N_18516,N_18723);
and U19481 (N_19481,N_18929,N_18502);
xnor U19482 (N_19482,N_18827,N_18634);
and U19483 (N_19483,N_18925,N_18656);
or U19484 (N_19484,N_18615,N_18732);
nand U19485 (N_19485,N_18917,N_18802);
nand U19486 (N_19486,N_18618,N_18839);
xor U19487 (N_19487,N_18631,N_18595);
nor U19488 (N_19488,N_18541,N_18974);
nor U19489 (N_19489,N_18781,N_18955);
nand U19490 (N_19490,N_18721,N_18677);
xnor U19491 (N_19491,N_18616,N_18905);
or U19492 (N_19492,N_18711,N_18807);
and U19493 (N_19493,N_18914,N_18532);
or U19494 (N_19494,N_18869,N_18584);
xnor U19495 (N_19495,N_18953,N_18516);
or U19496 (N_19496,N_18617,N_18892);
nand U19497 (N_19497,N_18695,N_18686);
nand U19498 (N_19498,N_18593,N_18718);
nor U19499 (N_19499,N_18726,N_18960);
and U19500 (N_19500,N_19337,N_19237);
nor U19501 (N_19501,N_19271,N_19484);
or U19502 (N_19502,N_19178,N_19233);
or U19503 (N_19503,N_19136,N_19048);
nor U19504 (N_19504,N_19309,N_19464);
and U19505 (N_19505,N_19344,N_19357);
or U19506 (N_19506,N_19373,N_19084);
nor U19507 (N_19507,N_19481,N_19314);
nand U19508 (N_19508,N_19386,N_19370);
or U19509 (N_19509,N_19135,N_19066);
nor U19510 (N_19510,N_19226,N_19022);
or U19511 (N_19511,N_19418,N_19041);
nand U19512 (N_19512,N_19438,N_19243);
xnor U19513 (N_19513,N_19017,N_19258);
or U19514 (N_19514,N_19212,N_19432);
or U19515 (N_19515,N_19261,N_19087);
and U19516 (N_19516,N_19256,N_19191);
nand U19517 (N_19517,N_19369,N_19074);
or U19518 (N_19518,N_19211,N_19238);
nand U19519 (N_19519,N_19359,N_19329);
xnor U19520 (N_19520,N_19296,N_19094);
nand U19521 (N_19521,N_19001,N_19196);
nor U19522 (N_19522,N_19322,N_19448);
and U19523 (N_19523,N_19060,N_19098);
or U19524 (N_19524,N_19132,N_19478);
nor U19525 (N_19525,N_19206,N_19489);
or U19526 (N_19526,N_19303,N_19086);
nand U19527 (N_19527,N_19100,N_19073);
nor U19528 (N_19528,N_19002,N_19106);
or U19529 (N_19529,N_19378,N_19148);
or U19530 (N_19530,N_19065,N_19328);
nor U19531 (N_19531,N_19468,N_19323);
xor U19532 (N_19532,N_19056,N_19031);
nor U19533 (N_19533,N_19277,N_19442);
or U19534 (N_19534,N_19294,N_19003);
nand U19535 (N_19535,N_19187,N_19299);
xor U19536 (N_19536,N_19388,N_19078);
nand U19537 (N_19537,N_19466,N_19321);
xor U19538 (N_19538,N_19488,N_19429);
or U19539 (N_19539,N_19397,N_19366);
nand U19540 (N_19540,N_19179,N_19394);
or U19541 (N_19541,N_19381,N_19401);
nor U19542 (N_19542,N_19362,N_19014);
and U19543 (N_19543,N_19114,N_19459);
nand U19544 (N_19544,N_19019,N_19199);
nor U19545 (N_19545,N_19312,N_19472);
and U19546 (N_19546,N_19159,N_19333);
xor U19547 (N_19547,N_19389,N_19101);
nor U19548 (N_19548,N_19130,N_19404);
nand U19549 (N_19549,N_19380,N_19324);
nor U19550 (N_19550,N_19213,N_19278);
or U19551 (N_19551,N_19456,N_19012);
or U19552 (N_19552,N_19234,N_19411);
xnor U19553 (N_19553,N_19257,N_19005);
and U19554 (N_19554,N_19255,N_19387);
nand U19555 (N_19555,N_19252,N_19058);
and U19556 (N_19556,N_19254,N_19368);
nor U19557 (N_19557,N_19482,N_19050);
nand U19558 (N_19558,N_19088,N_19280);
xnor U19559 (N_19559,N_19289,N_19297);
or U19560 (N_19560,N_19232,N_19108);
xor U19561 (N_19561,N_19247,N_19218);
and U19562 (N_19562,N_19485,N_19200);
and U19563 (N_19563,N_19365,N_19497);
and U19564 (N_19564,N_19245,N_19047);
nor U19565 (N_19565,N_19051,N_19240);
nor U19566 (N_19566,N_19209,N_19061);
and U19567 (N_19567,N_19391,N_19334);
xor U19568 (N_19568,N_19339,N_19253);
xor U19569 (N_19569,N_19099,N_19295);
nor U19570 (N_19570,N_19142,N_19119);
and U19571 (N_19571,N_19204,N_19096);
nor U19572 (N_19572,N_19110,N_19330);
xnor U19573 (N_19573,N_19076,N_19029);
xnor U19574 (N_19574,N_19157,N_19189);
xor U19575 (N_19575,N_19044,N_19140);
nor U19576 (N_19576,N_19180,N_19230);
or U19577 (N_19577,N_19393,N_19379);
nand U19578 (N_19578,N_19037,N_19340);
xor U19579 (N_19579,N_19267,N_19409);
and U19580 (N_19580,N_19195,N_19287);
and U19581 (N_19581,N_19040,N_19053);
and U19582 (N_19582,N_19461,N_19275);
xor U19583 (N_19583,N_19281,N_19118);
nand U19584 (N_19584,N_19355,N_19408);
nor U19585 (N_19585,N_19122,N_19049);
and U19586 (N_19586,N_19239,N_19385);
or U19587 (N_19587,N_19131,N_19090);
and U19588 (N_19588,N_19374,N_19483);
nor U19589 (N_19589,N_19134,N_19172);
nor U19590 (N_19590,N_19062,N_19499);
nor U19591 (N_19591,N_19462,N_19176);
and U19592 (N_19592,N_19476,N_19460);
and U19593 (N_19593,N_19085,N_19165);
nor U19594 (N_19594,N_19444,N_19128);
and U19595 (N_19595,N_19479,N_19197);
xnor U19596 (N_19596,N_19000,N_19454);
xor U19597 (N_19597,N_19080,N_19198);
or U19598 (N_19598,N_19354,N_19072);
nor U19599 (N_19599,N_19112,N_19302);
nor U19600 (N_19600,N_19286,N_19124);
xor U19601 (N_19601,N_19470,N_19015);
and U19602 (N_19602,N_19054,N_19282);
and U19603 (N_19603,N_19417,N_19202);
and U19604 (N_19604,N_19452,N_19268);
and U19605 (N_19605,N_19270,N_19467);
nand U19606 (N_19606,N_19445,N_19376);
nand U19607 (N_19607,N_19225,N_19463);
nand U19608 (N_19608,N_19071,N_19350);
or U19609 (N_19609,N_19410,N_19293);
nand U19610 (N_19610,N_19447,N_19127);
and U19611 (N_19611,N_19011,N_19347);
and U19612 (N_19612,N_19116,N_19325);
xnor U19613 (N_19613,N_19009,N_19228);
nand U19614 (N_19614,N_19210,N_19190);
and U19615 (N_19615,N_19120,N_19193);
nor U19616 (N_19616,N_19244,N_19251);
or U19617 (N_19617,N_19338,N_19398);
and U19618 (N_19618,N_19371,N_19335);
and U19619 (N_19619,N_19317,N_19490);
xor U19620 (N_19620,N_19104,N_19351);
nand U19621 (N_19621,N_19182,N_19349);
or U19622 (N_19622,N_19064,N_19138);
nand U19623 (N_19623,N_19471,N_19346);
and U19624 (N_19624,N_19079,N_19208);
nand U19625 (N_19625,N_19423,N_19006);
and U19626 (N_19626,N_19276,N_19183);
xnor U19627 (N_19627,N_19420,N_19095);
nor U19628 (N_19628,N_19327,N_19181);
nand U19629 (N_19629,N_19262,N_19169);
or U19630 (N_19630,N_19400,N_19161);
xor U19631 (N_19631,N_19004,N_19020);
xnor U19632 (N_19632,N_19170,N_19434);
or U19633 (N_19633,N_19168,N_19216);
or U19634 (N_19634,N_19077,N_19046);
or U19635 (N_19635,N_19144,N_19083);
xnor U19636 (N_19636,N_19129,N_19111);
nand U19637 (N_19637,N_19487,N_19052);
or U19638 (N_19638,N_19057,N_19318);
or U19639 (N_19639,N_19115,N_19407);
nor U19640 (N_19640,N_19364,N_19455);
nand U19641 (N_19641,N_19160,N_19308);
nand U19642 (N_19642,N_19320,N_19474);
nor U19643 (N_19643,N_19345,N_19413);
nor U19644 (N_19644,N_19185,N_19173);
and U19645 (N_19645,N_19439,N_19477);
xor U19646 (N_19646,N_19032,N_19224);
nor U19647 (N_19647,N_19028,N_19375);
or U19648 (N_19648,N_19141,N_19306);
xor U19649 (N_19649,N_19227,N_19026);
nand U19650 (N_19650,N_19266,N_19203);
xor U19651 (N_19651,N_19008,N_19291);
nor U19652 (N_19652,N_19465,N_19236);
nand U19653 (N_19653,N_19486,N_19310);
nor U19654 (N_19654,N_19133,N_19450);
nor U19655 (N_19655,N_19194,N_19038);
or U19656 (N_19656,N_19153,N_19360);
and U19657 (N_19657,N_19403,N_19356);
or U19658 (N_19658,N_19363,N_19152);
nor U19659 (N_19659,N_19125,N_19395);
and U19660 (N_19660,N_19042,N_19214);
nor U19661 (N_19661,N_19425,N_19146);
and U19662 (N_19662,N_19348,N_19428);
nor U19663 (N_19663,N_19025,N_19343);
xor U19664 (N_19664,N_19081,N_19402);
nand U19665 (N_19665,N_19443,N_19021);
xnor U19666 (N_19666,N_19219,N_19436);
nor U19667 (N_19667,N_19033,N_19092);
xnor U19668 (N_19668,N_19188,N_19039);
xnor U19669 (N_19669,N_19121,N_19301);
nand U19670 (N_19670,N_19155,N_19451);
nor U19671 (N_19671,N_19435,N_19298);
nand U19672 (N_19672,N_19458,N_19264);
nand U19673 (N_19673,N_19184,N_19024);
nor U19674 (N_19674,N_19269,N_19035);
nand U19675 (N_19675,N_19067,N_19272);
nand U19676 (N_19676,N_19105,N_19384);
and U19677 (N_19677,N_19171,N_19126);
or U19678 (N_19678,N_19068,N_19300);
and U19679 (N_19679,N_19036,N_19186);
xor U19680 (N_19680,N_19361,N_19235);
nand U19681 (N_19681,N_19358,N_19290);
and U19682 (N_19682,N_19283,N_19336);
xor U19683 (N_19683,N_19010,N_19332);
or U19684 (N_19684,N_19241,N_19396);
nor U19685 (N_19685,N_19475,N_19150);
xnor U19686 (N_19686,N_19063,N_19457);
or U19687 (N_19687,N_19311,N_19034);
nand U19688 (N_19688,N_19422,N_19201);
xor U19689 (N_19689,N_19163,N_19285);
xor U19690 (N_19690,N_19491,N_19453);
nor U19691 (N_19691,N_19151,N_19431);
nand U19692 (N_19692,N_19223,N_19433);
or U19693 (N_19693,N_19059,N_19082);
nor U19694 (N_19694,N_19414,N_19249);
xor U19695 (N_19695,N_19158,N_19440);
nor U19696 (N_19696,N_19390,N_19473);
and U19697 (N_19697,N_19229,N_19259);
or U19698 (N_19698,N_19217,N_19016);
or U19699 (N_19699,N_19156,N_19342);
xnor U19700 (N_19700,N_19273,N_19449);
or U19701 (N_19701,N_19246,N_19313);
nand U19702 (N_19702,N_19341,N_19372);
and U19703 (N_19703,N_19089,N_19167);
xor U19704 (N_19704,N_19419,N_19288);
xnor U19705 (N_19705,N_19207,N_19353);
or U19706 (N_19706,N_19107,N_19027);
xnor U19707 (N_19707,N_19139,N_19304);
and U19708 (N_19708,N_19215,N_19030);
and U19709 (N_19709,N_19284,N_19043);
xor U19710 (N_19710,N_19307,N_19424);
xor U19711 (N_19711,N_19430,N_19143);
xor U19712 (N_19712,N_19437,N_19222);
nand U19713 (N_19713,N_19495,N_19469);
and U19714 (N_19714,N_19292,N_19205);
nor U19715 (N_19715,N_19279,N_19498);
nor U19716 (N_19716,N_19315,N_19441);
nor U19717 (N_19717,N_19421,N_19352);
or U19718 (N_19718,N_19109,N_19177);
nand U19719 (N_19719,N_19263,N_19416);
nor U19720 (N_19720,N_19007,N_19174);
and U19721 (N_19721,N_19166,N_19274);
nand U19722 (N_19722,N_19162,N_19221);
and U19723 (N_19723,N_19117,N_19392);
or U19724 (N_19724,N_19316,N_19137);
nand U19725 (N_19725,N_19220,N_19097);
xnor U19726 (N_19726,N_19480,N_19415);
nor U19727 (N_19727,N_19147,N_19248);
nand U19728 (N_19728,N_19427,N_19493);
nand U19729 (N_19729,N_19494,N_19164);
and U19730 (N_19730,N_19069,N_19382);
and U19731 (N_19731,N_19013,N_19145);
nor U19732 (N_19732,N_19250,N_19102);
and U19733 (N_19733,N_19070,N_19260);
nor U19734 (N_19734,N_19075,N_19383);
nor U19735 (N_19735,N_19192,N_19496);
nand U19736 (N_19736,N_19319,N_19149);
nand U19737 (N_19737,N_19055,N_19093);
xnor U19738 (N_19738,N_19399,N_19175);
or U19739 (N_19739,N_19406,N_19123);
nor U19740 (N_19740,N_19446,N_19377);
nor U19741 (N_19741,N_19412,N_19113);
or U19742 (N_19742,N_19091,N_19331);
and U19743 (N_19743,N_19231,N_19426);
nand U19744 (N_19744,N_19326,N_19154);
nor U19745 (N_19745,N_19018,N_19405);
or U19746 (N_19746,N_19103,N_19367);
and U19747 (N_19747,N_19242,N_19305);
nor U19748 (N_19748,N_19045,N_19023);
or U19749 (N_19749,N_19492,N_19265);
nor U19750 (N_19750,N_19449,N_19387);
nand U19751 (N_19751,N_19375,N_19291);
nor U19752 (N_19752,N_19221,N_19000);
xor U19753 (N_19753,N_19481,N_19020);
or U19754 (N_19754,N_19333,N_19312);
or U19755 (N_19755,N_19073,N_19078);
and U19756 (N_19756,N_19295,N_19133);
and U19757 (N_19757,N_19158,N_19339);
nand U19758 (N_19758,N_19154,N_19240);
or U19759 (N_19759,N_19173,N_19456);
nor U19760 (N_19760,N_19124,N_19448);
nor U19761 (N_19761,N_19036,N_19297);
nand U19762 (N_19762,N_19137,N_19059);
or U19763 (N_19763,N_19319,N_19092);
and U19764 (N_19764,N_19409,N_19013);
nand U19765 (N_19765,N_19068,N_19235);
and U19766 (N_19766,N_19177,N_19252);
xor U19767 (N_19767,N_19465,N_19135);
nor U19768 (N_19768,N_19096,N_19169);
nor U19769 (N_19769,N_19255,N_19332);
and U19770 (N_19770,N_19178,N_19311);
xor U19771 (N_19771,N_19262,N_19301);
or U19772 (N_19772,N_19411,N_19041);
or U19773 (N_19773,N_19289,N_19202);
or U19774 (N_19774,N_19276,N_19176);
xnor U19775 (N_19775,N_19481,N_19258);
and U19776 (N_19776,N_19170,N_19258);
xor U19777 (N_19777,N_19456,N_19313);
xnor U19778 (N_19778,N_19094,N_19279);
nand U19779 (N_19779,N_19458,N_19457);
nor U19780 (N_19780,N_19161,N_19490);
nand U19781 (N_19781,N_19431,N_19209);
nand U19782 (N_19782,N_19000,N_19141);
xor U19783 (N_19783,N_19117,N_19406);
nand U19784 (N_19784,N_19155,N_19447);
xor U19785 (N_19785,N_19004,N_19016);
xnor U19786 (N_19786,N_19145,N_19404);
and U19787 (N_19787,N_19459,N_19334);
xnor U19788 (N_19788,N_19478,N_19048);
nor U19789 (N_19789,N_19068,N_19213);
or U19790 (N_19790,N_19365,N_19064);
nand U19791 (N_19791,N_19317,N_19083);
nor U19792 (N_19792,N_19343,N_19349);
and U19793 (N_19793,N_19110,N_19208);
and U19794 (N_19794,N_19389,N_19017);
or U19795 (N_19795,N_19387,N_19213);
nand U19796 (N_19796,N_19452,N_19005);
or U19797 (N_19797,N_19211,N_19439);
and U19798 (N_19798,N_19115,N_19435);
or U19799 (N_19799,N_19129,N_19127);
or U19800 (N_19800,N_19284,N_19031);
nor U19801 (N_19801,N_19276,N_19150);
nand U19802 (N_19802,N_19360,N_19252);
xor U19803 (N_19803,N_19029,N_19261);
and U19804 (N_19804,N_19130,N_19235);
nor U19805 (N_19805,N_19078,N_19235);
and U19806 (N_19806,N_19491,N_19331);
nand U19807 (N_19807,N_19154,N_19440);
nor U19808 (N_19808,N_19190,N_19371);
xor U19809 (N_19809,N_19193,N_19103);
nor U19810 (N_19810,N_19088,N_19409);
nand U19811 (N_19811,N_19168,N_19369);
nor U19812 (N_19812,N_19012,N_19000);
nand U19813 (N_19813,N_19028,N_19452);
nor U19814 (N_19814,N_19257,N_19171);
and U19815 (N_19815,N_19203,N_19179);
and U19816 (N_19816,N_19362,N_19403);
nor U19817 (N_19817,N_19181,N_19434);
nor U19818 (N_19818,N_19147,N_19412);
xnor U19819 (N_19819,N_19219,N_19399);
and U19820 (N_19820,N_19157,N_19004);
nor U19821 (N_19821,N_19221,N_19475);
and U19822 (N_19822,N_19022,N_19471);
nand U19823 (N_19823,N_19125,N_19423);
and U19824 (N_19824,N_19430,N_19421);
and U19825 (N_19825,N_19460,N_19025);
nor U19826 (N_19826,N_19319,N_19296);
xor U19827 (N_19827,N_19333,N_19120);
nor U19828 (N_19828,N_19471,N_19099);
nand U19829 (N_19829,N_19371,N_19318);
xor U19830 (N_19830,N_19472,N_19146);
xor U19831 (N_19831,N_19466,N_19085);
nor U19832 (N_19832,N_19442,N_19070);
xnor U19833 (N_19833,N_19416,N_19015);
xor U19834 (N_19834,N_19215,N_19489);
xnor U19835 (N_19835,N_19371,N_19450);
nand U19836 (N_19836,N_19132,N_19092);
nor U19837 (N_19837,N_19136,N_19200);
and U19838 (N_19838,N_19090,N_19378);
xor U19839 (N_19839,N_19225,N_19178);
xor U19840 (N_19840,N_19290,N_19269);
or U19841 (N_19841,N_19059,N_19488);
or U19842 (N_19842,N_19143,N_19013);
nand U19843 (N_19843,N_19328,N_19235);
nand U19844 (N_19844,N_19217,N_19238);
xnor U19845 (N_19845,N_19192,N_19265);
and U19846 (N_19846,N_19223,N_19312);
or U19847 (N_19847,N_19348,N_19281);
or U19848 (N_19848,N_19046,N_19326);
nand U19849 (N_19849,N_19017,N_19454);
xor U19850 (N_19850,N_19220,N_19319);
or U19851 (N_19851,N_19019,N_19214);
nand U19852 (N_19852,N_19297,N_19157);
and U19853 (N_19853,N_19146,N_19109);
or U19854 (N_19854,N_19416,N_19482);
and U19855 (N_19855,N_19464,N_19075);
or U19856 (N_19856,N_19142,N_19096);
and U19857 (N_19857,N_19070,N_19160);
and U19858 (N_19858,N_19425,N_19270);
nor U19859 (N_19859,N_19108,N_19438);
xor U19860 (N_19860,N_19280,N_19467);
or U19861 (N_19861,N_19233,N_19172);
and U19862 (N_19862,N_19314,N_19174);
or U19863 (N_19863,N_19088,N_19243);
or U19864 (N_19864,N_19319,N_19013);
nand U19865 (N_19865,N_19337,N_19399);
nand U19866 (N_19866,N_19475,N_19152);
and U19867 (N_19867,N_19229,N_19267);
xnor U19868 (N_19868,N_19123,N_19255);
or U19869 (N_19869,N_19437,N_19372);
xor U19870 (N_19870,N_19349,N_19172);
nor U19871 (N_19871,N_19055,N_19164);
xor U19872 (N_19872,N_19265,N_19109);
nand U19873 (N_19873,N_19433,N_19361);
or U19874 (N_19874,N_19031,N_19047);
nor U19875 (N_19875,N_19053,N_19266);
and U19876 (N_19876,N_19209,N_19223);
nor U19877 (N_19877,N_19267,N_19319);
or U19878 (N_19878,N_19068,N_19190);
nand U19879 (N_19879,N_19045,N_19220);
nand U19880 (N_19880,N_19274,N_19361);
nor U19881 (N_19881,N_19107,N_19323);
and U19882 (N_19882,N_19484,N_19032);
xor U19883 (N_19883,N_19232,N_19497);
or U19884 (N_19884,N_19034,N_19255);
xnor U19885 (N_19885,N_19097,N_19207);
and U19886 (N_19886,N_19082,N_19157);
xor U19887 (N_19887,N_19244,N_19365);
nand U19888 (N_19888,N_19219,N_19083);
xor U19889 (N_19889,N_19210,N_19213);
xnor U19890 (N_19890,N_19123,N_19407);
xnor U19891 (N_19891,N_19215,N_19243);
and U19892 (N_19892,N_19001,N_19088);
xor U19893 (N_19893,N_19161,N_19358);
or U19894 (N_19894,N_19130,N_19115);
nand U19895 (N_19895,N_19413,N_19034);
nand U19896 (N_19896,N_19292,N_19222);
nand U19897 (N_19897,N_19181,N_19118);
or U19898 (N_19898,N_19494,N_19014);
or U19899 (N_19899,N_19279,N_19384);
nand U19900 (N_19900,N_19009,N_19208);
nor U19901 (N_19901,N_19013,N_19140);
nand U19902 (N_19902,N_19295,N_19288);
and U19903 (N_19903,N_19486,N_19460);
xnor U19904 (N_19904,N_19492,N_19328);
nor U19905 (N_19905,N_19154,N_19401);
xnor U19906 (N_19906,N_19413,N_19454);
nand U19907 (N_19907,N_19009,N_19268);
nand U19908 (N_19908,N_19306,N_19491);
nor U19909 (N_19909,N_19424,N_19402);
and U19910 (N_19910,N_19266,N_19127);
and U19911 (N_19911,N_19383,N_19406);
or U19912 (N_19912,N_19101,N_19158);
nor U19913 (N_19913,N_19134,N_19225);
and U19914 (N_19914,N_19182,N_19488);
xnor U19915 (N_19915,N_19037,N_19278);
xnor U19916 (N_19916,N_19006,N_19067);
nand U19917 (N_19917,N_19291,N_19128);
or U19918 (N_19918,N_19204,N_19114);
or U19919 (N_19919,N_19251,N_19315);
xor U19920 (N_19920,N_19416,N_19101);
or U19921 (N_19921,N_19365,N_19124);
nand U19922 (N_19922,N_19426,N_19161);
and U19923 (N_19923,N_19015,N_19050);
nand U19924 (N_19924,N_19487,N_19076);
or U19925 (N_19925,N_19123,N_19475);
xnor U19926 (N_19926,N_19290,N_19096);
nor U19927 (N_19927,N_19339,N_19233);
xor U19928 (N_19928,N_19377,N_19056);
nand U19929 (N_19929,N_19382,N_19288);
nand U19930 (N_19930,N_19466,N_19110);
nor U19931 (N_19931,N_19054,N_19255);
and U19932 (N_19932,N_19297,N_19029);
and U19933 (N_19933,N_19271,N_19066);
nand U19934 (N_19934,N_19467,N_19404);
nor U19935 (N_19935,N_19267,N_19153);
and U19936 (N_19936,N_19292,N_19437);
or U19937 (N_19937,N_19025,N_19483);
or U19938 (N_19938,N_19350,N_19407);
xor U19939 (N_19939,N_19092,N_19017);
xor U19940 (N_19940,N_19198,N_19095);
and U19941 (N_19941,N_19096,N_19114);
nor U19942 (N_19942,N_19295,N_19430);
nor U19943 (N_19943,N_19082,N_19056);
nor U19944 (N_19944,N_19023,N_19189);
nand U19945 (N_19945,N_19124,N_19195);
nor U19946 (N_19946,N_19120,N_19115);
nand U19947 (N_19947,N_19256,N_19008);
nand U19948 (N_19948,N_19193,N_19100);
nor U19949 (N_19949,N_19432,N_19232);
or U19950 (N_19950,N_19030,N_19177);
xor U19951 (N_19951,N_19243,N_19496);
and U19952 (N_19952,N_19175,N_19216);
or U19953 (N_19953,N_19316,N_19177);
or U19954 (N_19954,N_19073,N_19010);
nor U19955 (N_19955,N_19196,N_19063);
nand U19956 (N_19956,N_19021,N_19166);
or U19957 (N_19957,N_19096,N_19199);
nor U19958 (N_19958,N_19279,N_19454);
and U19959 (N_19959,N_19153,N_19323);
nor U19960 (N_19960,N_19118,N_19267);
nand U19961 (N_19961,N_19303,N_19177);
or U19962 (N_19962,N_19260,N_19313);
and U19963 (N_19963,N_19096,N_19094);
xnor U19964 (N_19964,N_19031,N_19113);
nor U19965 (N_19965,N_19291,N_19313);
and U19966 (N_19966,N_19243,N_19285);
and U19967 (N_19967,N_19292,N_19127);
xnor U19968 (N_19968,N_19122,N_19482);
xor U19969 (N_19969,N_19397,N_19052);
and U19970 (N_19970,N_19356,N_19380);
or U19971 (N_19971,N_19147,N_19230);
xor U19972 (N_19972,N_19365,N_19166);
nand U19973 (N_19973,N_19002,N_19353);
xnor U19974 (N_19974,N_19292,N_19125);
nand U19975 (N_19975,N_19147,N_19117);
nand U19976 (N_19976,N_19027,N_19466);
and U19977 (N_19977,N_19168,N_19062);
xor U19978 (N_19978,N_19312,N_19259);
or U19979 (N_19979,N_19216,N_19239);
and U19980 (N_19980,N_19486,N_19125);
xor U19981 (N_19981,N_19019,N_19446);
nor U19982 (N_19982,N_19118,N_19184);
nor U19983 (N_19983,N_19032,N_19293);
nor U19984 (N_19984,N_19085,N_19408);
xnor U19985 (N_19985,N_19474,N_19447);
and U19986 (N_19986,N_19426,N_19247);
xnor U19987 (N_19987,N_19015,N_19199);
nand U19988 (N_19988,N_19420,N_19401);
or U19989 (N_19989,N_19033,N_19155);
nor U19990 (N_19990,N_19344,N_19216);
or U19991 (N_19991,N_19068,N_19168);
nor U19992 (N_19992,N_19258,N_19437);
or U19993 (N_19993,N_19471,N_19053);
and U19994 (N_19994,N_19169,N_19198);
nand U19995 (N_19995,N_19243,N_19130);
and U19996 (N_19996,N_19088,N_19470);
or U19997 (N_19997,N_19370,N_19237);
xor U19998 (N_19998,N_19275,N_19167);
or U19999 (N_19999,N_19456,N_19164);
nor U20000 (N_20000,N_19692,N_19869);
xnor U20001 (N_20001,N_19826,N_19661);
and U20002 (N_20002,N_19996,N_19884);
or U20003 (N_20003,N_19964,N_19715);
xor U20004 (N_20004,N_19740,N_19594);
nand U20005 (N_20005,N_19879,N_19545);
nor U20006 (N_20006,N_19628,N_19749);
nand U20007 (N_20007,N_19702,N_19755);
or U20008 (N_20008,N_19639,N_19575);
or U20009 (N_20009,N_19974,N_19941);
xnor U20010 (N_20010,N_19846,N_19560);
xor U20011 (N_20011,N_19588,N_19958);
nor U20012 (N_20012,N_19712,N_19893);
nand U20013 (N_20013,N_19946,N_19921);
or U20014 (N_20014,N_19744,N_19577);
xor U20015 (N_20015,N_19798,N_19728);
and U20016 (N_20016,N_19844,N_19993);
nand U20017 (N_20017,N_19595,N_19885);
nor U20018 (N_20018,N_19512,N_19932);
xor U20019 (N_20019,N_19853,N_19883);
nand U20020 (N_20020,N_19587,N_19697);
and U20021 (N_20021,N_19904,N_19979);
nor U20022 (N_20022,N_19854,N_19604);
or U20023 (N_20023,N_19813,N_19818);
nor U20024 (N_20024,N_19583,N_19747);
or U20025 (N_20025,N_19616,N_19934);
nand U20026 (N_20026,N_19589,N_19930);
nor U20027 (N_20027,N_19637,N_19889);
nand U20028 (N_20028,N_19732,N_19614);
or U20029 (N_20029,N_19647,N_19871);
nor U20030 (N_20030,N_19986,N_19901);
nand U20031 (N_20031,N_19551,N_19806);
and U20032 (N_20032,N_19668,N_19786);
nand U20033 (N_20033,N_19693,N_19772);
nand U20034 (N_20034,N_19805,N_19836);
and U20035 (N_20035,N_19540,N_19924);
or U20036 (N_20036,N_19507,N_19689);
nor U20037 (N_20037,N_19601,N_19652);
or U20038 (N_20038,N_19635,N_19925);
nand U20039 (N_20039,N_19777,N_19988);
nor U20040 (N_20040,N_19723,N_19566);
and U20041 (N_20041,N_19721,N_19593);
and U20042 (N_20042,N_19963,N_19664);
and U20043 (N_20043,N_19649,N_19838);
xor U20044 (N_20044,N_19841,N_19731);
nor U20045 (N_20045,N_19817,N_19768);
xnor U20046 (N_20046,N_19994,N_19918);
nor U20047 (N_20047,N_19691,N_19896);
nor U20048 (N_20048,N_19665,N_19726);
nor U20049 (N_20049,N_19790,N_19951);
xnor U20050 (N_20050,N_19567,N_19686);
nor U20051 (N_20051,N_19807,N_19950);
and U20052 (N_20052,N_19849,N_19799);
or U20053 (N_20053,N_19761,N_19876);
xor U20054 (N_20054,N_19770,N_19877);
xor U20055 (N_20055,N_19984,N_19911);
xnor U20056 (N_20056,N_19511,N_19792);
nor U20057 (N_20057,N_19831,N_19961);
or U20058 (N_20058,N_19613,N_19793);
nor U20059 (N_20059,N_19645,N_19662);
nand U20060 (N_20060,N_19959,N_19558);
nand U20061 (N_20061,N_19833,N_19561);
xor U20062 (N_20062,N_19821,N_19825);
or U20063 (N_20063,N_19698,N_19823);
or U20064 (N_20064,N_19590,N_19940);
nand U20065 (N_20065,N_19573,N_19928);
xnor U20066 (N_20066,N_19773,N_19520);
xor U20067 (N_20067,N_19724,N_19529);
nor U20068 (N_20068,N_19743,N_19803);
nor U20069 (N_20069,N_19975,N_19978);
and U20070 (N_20070,N_19982,N_19801);
nand U20071 (N_20071,N_19788,N_19919);
or U20072 (N_20072,N_19555,N_19537);
xnor U20073 (N_20073,N_19960,N_19699);
and U20074 (N_20074,N_19685,N_19987);
xor U20075 (N_20075,N_19864,N_19599);
and U20076 (N_20076,N_19542,N_19630);
and U20077 (N_20077,N_19525,N_19952);
nand U20078 (N_20078,N_19648,N_19582);
nand U20079 (N_20079,N_19868,N_19912);
nor U20080 (N_20080,N_19535,N_19569);
or U20081 (N_20081,N_19713,N_19842);
and U20082 (N_20082,N_19553,N_19625);
xnor U20083 (N_20083,N_19830,N_19631);
and U20084 (N_20084,N_19920,N_19766);
nor U20085 (N_20085,N_19977,N_19654);
xor U20086 (N_20086,N_19727,N_19804);
xnor U20087 (N_20087,N_19722,N_19969);
nand U20088 (N_20088,N_19967,N_19612);
nand U20089 (N_20089,N_19579,N_19906);
xnor U20090 (N_20090,N_19784,N_19863);
or U20091 (N_20091,N_19767,N_19633);
and U20092 (N_20092,N_19684,N_19933);
nand U20093 (N_20093,N_19531,N_19550);
nor U20094 (N_20094,N_19745,N_19910);
xor U20095 (N_20095,N_19903,N_19942);
and U20096 (N_20096,N_19992,N_19694);
and U20097 (N_20097,N_19900,N_19897);
nand U20098 (N_20098,N_19541,N_19629);
nand U20099 (N_20099,N_19638,N_19819);
and U20100 (N_20100,N_19677,N_19608);
nor U20101 (N_20101,N_19509,N_19563);
xor U20102 (N_20102,N_19929,N_19999);
xor U20103 (N_20103,N_19789,N_19576);
and U20104 (N_20104,N_19760,N_19927);
nor U20105 (N_20105,N_19701,N_19711);
nand U20106 (N_20106,N_19667,N_19671);
nor U20107 (N_20107,N_19778,N_19559);
xnor U20108 (N_20108,N_19687,N_19754);
or U20109 (N_20109,N_19843,N_19568);
nor U20110 (N_20110,N_19953,N_19794);
xnor U20111 (N_20111,N_19973,N_19503);
and U20112 (N_20112,N_19516,N_19617);
or U20113 (N_20113,N_19748,N_19666);
and U20114 (N_20114,N_19522,N_19533);
xor U20115 (N_20115,N_19966,N_19624);
and U20116 (N_20116,N_19815,N_19640);
nand U20117 (N_20117,N_19539,N_19812);
xor U20118 (N_20118,N_19546,N_19899);
nand U20119 (N_20119,N_19873,N_19673);
nor U20120 (N_20120,N_19787,N_19584);
or U20121 (N_20121,N_19502,N_19945);
and U20122 (N_20122,N_19622,N_19554);
or U20123 (N_20123,N_19870,N_19898);
nand U20124 (N_20124,N_19644,N_19949);
or U20125 (N_20125,N_19508,N_19556);
xnor U20126 (N_20126,N_19970,N_19890);
nor U20127 (N_20127,N_19954,N_19695);
nand U20128 (N_20128,N_19971,N_19678);
xnor U20129 (N_20129,N_19562,N_19708);
nor U20130 (N_20130,N_19549,N_19866);
and U20131 (N_20131,N_19659,N_19922);
or U20132 (N_20132,N_19943,N_19565);
and U20133 (N_20133,N_19600,N_19504);
or U20134 (N_20134,N_19814,N_19956);
or U20135 (N_20135,N_19995,N_19874);
or U20136 (N_20136,N_19705,N_19968);
nor U20137 (N_20137,N_19962,N_19634);
and U20138 (N_20138,N_19626,N_19811);
xnor U20139 (N_20139,N_19653,N_19780);
nand U20140 (N_20140,N_19886,N_19643);
nor U20141 (N_20141,N_19672,N_19730);
and U20142 (N_20142,N_19517,N_19704);
or U20143 (N_20143,N_19955,N_19658);
or U20144 (N_20144,N_19936,N_19717);
nand U20145 (N_20145,N_19750,N_19719);
nor U20146 (N_20146,N_19742,N_19603);
xor U20147 (N_20147,N_19720,N_19738);
or U20148 (N_20148,N_19769,N_19515);
or U20149 (N_20149,N_19574,N_19675);
and U20150 (N_20150,N_19669,N_19880);
xor U20151 (N_20151,N_19636,N_19981);
nand U20152 (N_20152,N_19564,N_19845);
or U20153 (N_20153,N_19592,N_19707);
and U20154 (N_20154,N_19598,N_19827);
nand U20155 (N_20155,N_19894,N_19581);
or U20156 (N_20156,N_19983,N_19552);
and U20157 (N_20157,N_19544,N_19532);
xnor U20158 (N_20158,N_19802,N_19834);
and U20159 (N_20159,N_19783,N_19623);
xor U20160 (N_20160,N_19824,N_19641);
nor U20161 (N_20161,N_19736,N_19944);
nand U20162 (N_20162,N_19580,N_19865);
and U20163 (N_20163,N_19935,N_19781);
or U20164 (N_20164,N_19500,N_19729);
and U20165 (N_20165,N_19670,N_19602);
or U20166 (N_20166,N_19538,N_19828);
xor U20167 (N_20167,N_19615,N_19548);
and U20168 (N_20168,N_19985,N_19850);
nand U20169 (N_20169,N_19820,N_19907);
or U20170 (N_20170,N_19696,N_19609);
nor U20171 (N_20171,N_19976,N_19752);
nand U20172 (N_20172,N_19832,N_19937);
nand U20173 (N_20173,N_19610,N_19611);
nor U20174 (N_20174,N_19570,N_19980);
nor U20175 (N_20175,N_19585,N_19757);
and U20176 (N_20176,N_19764,N_19632);
nor U20177 (N_20177,N_19578,N_19855);
nor U20178 (N_20178,N_19858,N_19605);
nand U20179 (N_20179,N_19680,N_19725);
or U20180 (N_20180,N_19856,N_19571);
nand U20181 (N_20181,N_19646,N_19829);
xnor U20182 (N_20182,N_19859,N_19779);
nor U20183 (N_20183,N_19867,N_19735);
xor U20184 (N_20184,N_19716,N_19771);
and U20185 (N_20185,N_19957,N_19683);
xor U20186 (N_20186,N_19872,N_19536);
nor U20187 (N_20187,N_19923,N_19796);
xor U20188 (N_20188,N_19762,N_19948);
nor U20189 (N_20189,N_19709,N_19892);
xnor U20190 (N_20190,N_19989,N_19753);
nor U20191 (N_20191,N_19875,N_19700);
nand U20192 (N_20192,N_19851,N_19913);
or U20193 (N_20193,N_19763,N_19857);
nor U20194 (N_20194,N_19656,N_19882);
nor U20195 (N_20195,N_19676,N_19916);
and U20196 (N_20196,N_19606,N_19690);
or U20197 (N_20197,N_19682,N_19914);
and U20198 (N_20198,N_19619,N_19751);
xor U20199 (N_20199,N_19908,N_19627);
nand U20200 (N_20200,N_19765,N_19607);
nor U20201 (N_20201,N_19674,N_19510);
and U20202 (N_20202,N_19852,N_19543);
or U20203 (N_20203,N_19746,N_19972);
xnor U20204 (N_20204,N_19990,N_19905);
and U20205 (N_20205,N_19513,N_19775);
xor U20206 (N_20206,N_19547,N_19997);
nand U20207 (N_20207,N_19862,N_19718);
nand U20208 (N_20208,N_19785,N_19518);
nor U20209 (N_20209,N_19759,N_19521);
and U20210 (N_20210,N_19909,N_19847);
nand U20211 (N_20211,N_19706,N_19642);
nor U20212 (N_20212,N_19505,N_19939);
xnor U20213 (N_20213,N_19557,N_19650);
nor U20214 (N_20214,N_19991,N_19837);
and U20215 (N_20215,N_19917,N_19931);
nor U20216 (N_20216,N_19938,N_19506);
and U20217 (N_20217,N_19572,N_19663);
nor U20218 (N_20218,N_19808,N_19688);
or U20219 (N_20219,N_19891,N_19527);
nand U20220 (N_20220,N_19887,N_19782);
or U20221 (N_20221,N_19530,N_19965);
nand U20222 (N_20222,N_19655,N_19878);
xnor U20223 (N_20223,N_19651,N_19620);
or U20224 (N_20224,N_19816,N_19947);
nand U20225 (N_20225,N_19758,N_19998);
and U20226 (N_20226,N_19881,N_19774);
xor U20227 (N_20227,N_19586,N_19519);
xnor U20228 (N_20228,N_19791,N_19657);
or U20229 (N_20229,N_19809,N_19741);
or U20230 (N_20230,N_19618,N_19756);
nand U20231 (N_20231,N_19848,N_19861);
xor U20232 (N_20232,N_19795,N_19733);
nor U20233 (N_20233,N_19902,N_19797);
nor U20234 (N_20234,N_19810,N_19926);
and U20235 (N_20235,N_19895,N_19523);
nand U20236 (N_20236,N_19915,N_19528);
xnor U20237 (N_20237,N_19714,N_19739);
and U20238 (N_20238,N_19591,N_19734);
nor U20239 (N_20239,N_19860,N_19597);
and U20240 (N_20240,N_19660,N_19835);
or U20241 (N_20241,N_19737,N_19524);
nand U20242 (N_20242,N_19776,N_19840);
and U20243 (N_20243,N_19526,N_19501);
or U20244 (N_20244,N_19888,N_19621);
nor U20245 (N_20245,N_19839,N_19534);
nand U20246 (N_20246,N_19514,N_19822);
and U20247 (N_20247,N_19800,N_19710);
and U20248 (N_20248,N_19703,N_19679);
or U20249 (N_20249,N_19681,N_19596);
nand U20250 (N_20250,N_19713,N_19962);
xor U20251 (N_20251,N_19603,N_19612);
nand U20252 (N_20252,N_19937,N_19882);
and U20253 (N_20253,N_19647,N_19737);
and U20254 (N_20254,N_19581,N_19862);
xor U20255 (N_20255,N_19552,N_19571);
or U20256 (N_20256,N_19731,N_19802);
nor U20257 (N_20257,N_19554,N_19899);
nand U20258 (N_20258,N_19762,N_19521);
or U20259 (N_20259,N_19940,N_19541);
nand U20260 (N_20260,N_19585,N_19912);
and U20261 (N_20261,N_19978,N_19904);
or U20262 (N_20262,N_19680,N_19988);
or U20263 (N_20263,N_19952,N_19824);
xnor U20264 (N_20264,N_19648,N_19669);
nor U20265 (N_20265,N_19785,N_19525);
xor U20266 (N_20266,N_19642,N_19875);
xnor U20267 (N_20267,N_19688,N_19638);
xnor U20268 (N_20268,N_19582,N_19690);
nor U20269 (N_20269,N_19627,N_19962);
and U20270 (N_20270,N_19576,N_19530);
nand U20271 (N_20271,N_19944,N_19793);
and U20272 (N_20272,N_19720,N_19867);
nand U20273 (N_20273,N_19793,N_19639);
nand U20274 (N_20274,N_19507,N_19979);
nor U20275 (N_20275,N_19722,N_19768);
xor U20276 (N_20276,N_19703,N_19814);
and U20277 (N_20277,N_19643,N_19992);
nor U20278 (N_20278,N_19550,N_19868);
xnor U20279 (N_20279,N_19836,N_19574);
nor U20280 (N_20280,N_19930,N_19840);
and U20281 (N_20281,N_19717,N_19590);
nor U20282 (N_20282,N_19590,N_19753);
nor U20283 (N_20283,N_19763,N_19526);
and U20284 (N_20284,N_19996,N_19991);
or U20285 (N_20285,N_19583,N_19993);
and U20286 (N_20286,N_19949,N_19724);
and U20287 (N_20287,N_19631,N_19780);
and U20288 (N_20288,N_19690,N_19781);
and U20289 (N_20289,N_19958,N_19653);
nor U20290 (N_20290,N_19608,N_19669);
nand U20291 (N_20291,N_19663,N_19600);
xnor U20292 (N_20292,N_19759,N_19671);
and U20293 (N_20293,N_19652,N_19537);
or U20294 (N_20294,N_19673,N_19847);
and U20295 (N_20295,N_19770,N_19842);
and U20296 (N_20296,N_19813,N_19765);
nand U20297 (N_20297,N_19502,N_19834);
and U20298 (N_20298,N_19996,N_19662);
xor U20299 (N_20299,N_19849,N_19670);
or U20300 (N_20300,N_19722,N_19555);
xor U20301 (N_20301,N_19525,N_19837);
or U20302 (N_20302,N_19950,N_19913);
or U20303 (N_20303,N_19966,N_19539);
nand U20304 (N_20304,N_19591,N_19722);
xnor U20305 (N_20305,N_19708,N_19938);
xor U20306 (N_20306,N_19945,N_19855);
or U20307 (N_20307,N_19556,N_19574);
or U20308 (N_20308,N_19517,N_19762);
or U20309 (N_20309,N_19778,N_19770);
nand U20310 (N_20310,N_19790,N_19747);
nand U20311 (N_20311,N_19675,N_19767);
or U20312 (N_20312,N_19838,N_19926);
nor U20313 (N_20313,N_19702,N_19918);
xnor U20314 (N_20314,N_19548,N_19893);
nor U20315 (N_20315,N_19731,N_19661);
nor U20316 (N_20316,N_19977,N_19910);
xnor U20317 (N_20317,N_19971,N_19961);
and U20318 (N_20318,N_19897,N_19759);
or U20319 (N_20319,N_19990,N_19985);
xnor U20320 (N_20320,N_19894,N_19748);
nand U20321 (N_20321,N_19936,N_19550);
nor U20322 (N_20322,N_19769,N_19968);
and U20323 (N_20323,N_19948,N_19994);
and U20324 (N_20324,N_19752,N_19944);
xor U20325 (N_20325,N_19958,N_19655);
nor U20326 (N_20326,N_19760,N_19979);
and U20327 (N_20327,N_19600,N_19597);
xor U20328 (N_20328,N_19631,N_19701);
or U20329 (N_20329,N_19581,N_19826);
nand U20330 (N_20330,N_19768,N_19656);
xnor U20331 (N_20331,N_19769,N_19709);
nand U20332 (N_20332,N_19870,N_19826);
or U20333 (N_20333,N_19600,N_19721);
and U20334 (N_20334,N_19665,N_19691);
or U20335 (N_20335,N_19895,N_19671);
or U20336 (N_20336,N_19755,N_19698);
xnor U20337 (N_20337,N_19978,N_19632);
xor U20338 (N_20338,N_19771,N_19838);
xor U20339 (N_20339,N_19776,N_19540);
xnor U20340 (N_20340,N_19729,N_19597);
nand U20341 (N_20341,N_19998,N_19975);
nand U20342 (N_20342,N_19824,N_19771);
or U20343 (N_20343,N_19768,N_19592);
nor U20344 (N_20344,N_19597,N_19827);
nor U20345 (N_20345,N_19777,N_19617);
and U20346 (N_20346,N_19770,N_19895);
nand U20347 (N_20347,N_19748,N_19871);
and U20348 (N_20348,N_19912,N_19582);
or U20349 (N_20349,N_19945,N_19631);
and U20350 (N_20350,N_19712,N_19530);
or U20351 (N_20351,N_19814,N_19541);
nor U20352 (N_20352,N_19545,N_19678);
nand U20353 (N_20353,N_19583,N_19717);
nor U20354 (N_20354,N_19509,N_19782);
and U20355 (N_20355,N_19597,N_19519);
nand U20356 (N_20356,N_19943,N_19501);
xor U20357 (N_20357,N_19888,N_19603);
nand U20358 (N_20358,N_19970,N_19997);
nor U20359 (N_20359,N_19565,N_19700);
nor U20360 (N_20360,N_19551,N_19809);
nor U20361 (N_20361,N_19559,N_19843);
xor U20362 (N_20362,N_19791,N_19522);
and U20363 (N_20363,N_19878,N_19785);
nor U20364 (N_20364,N_19510,N_19689);
nand U20365 (N_20365,N_19887,N_19832);
nor U20366 (N_20366,N_19736,N_19647);
nand U20367 (N_20367,N_19985,N_19895);
or U20368 (N_20368,N_19958,N_19847);
or U20369 (N_20369,N_19637,N_19800);
and U20370 (N_20370,N_19742,N_19501);
or U20371 (N_20371,N_19600,N_19964);
or U20372 (N_20372,N_19556,N_19610);
nand U20373 (N_20373,N_19938,N_19638);
or U20374 (N_20374,N_19623,N_19996);
and U20375 (N_20375,N_19969,N_19598);
and U20376 (N_20376,N_19973,N_19600);
nand U20377 (N_20377,N_19614,N_19968);
and U20378 (N_20378,N_19583,N_19973);
xor U20379 (N_20379,N_19946,N_19998);
or U20380 (N_20380,N_19672,N_19990);
nor U20381 (N_20381,N_19583,N_19565);
nand U20382 (N_20382,N_19570,N_19945);
nor U20383 (N_20383,N_19611,N_19724);
or U20384 (N_20384,N_19518,N_19535);
and U20385 (N_20385,N_19551,N_19531);
nor U20386 (N_20386,N_19977,N_19831);
and U20387 (N_20387,N_19785,N_19594);
nor U20388 (N_20388,N_19864,N_19917);
or U20389 (N_20389,N_19560,N_19991);
xnor U20390 (N_20390,N_19758,N_19506);
xnor U20391 (N_20391,N_19711,N_19791);
xnor U20392 (N_20392,N_19838,N_19610);
nor U20393 (N_20393,N_19979,N_19871);
nand U20394 (N_20394,N_19817,N_19590);
and U20395 (N_20395,N_19614,N_19831);
or U20396 (N_20396,N_19510,N_19616);
and U20397 (N_20397,N_19711,N_19652);
and U20398 (N_20398,N_19818,N_19623);
xor U20399 (N_20399,N_19750,N_19892);
xor U20400 (N_20400,N_19900,N_19561);
nor U20401 (N_20401,N_19995,N_19603);
nand U20402 (N_20402,N_19551,N_19588);
nand U20403 (N_20403,N_19564,N_19649);
nand U20404 (N_20404,N_19645,N_19845);
nand U20405 (N_20405,N_19858,N_19878);
xnor U20406 (N_20406,N_19570,N_19652);
xor U20407 (N_20407,N_19925,N_19621);
and U20408 (N_20408,N_19831,N_19860);
xnor U20409 (N_20409,N_19527,N_19893);
nand U20410 (N_20410,N_19547,N_19840);
nand U20411 (N_20411,N_19653,N_19644);
nor U20412 (N_20412,N_19929,N_19708);
nor U20413 (N_20413,N_19506,N_19606);
xor U20414 (N_20414,N_19720,N_19977);
nor U20415 (N_20415,N_19984,N_19946);
xor U20416 (N_20416,N_19767,N_19920);
xnor U20417 (N_20417,N_19707,N_19555);
nor U20418 (N_20418,N_19800,N_19654);
nor U20419 (N_20419,N_19779,N_19815);
nor U20420 (N_20420,N_19681,N_19827);
nand U20421 (N_20421,N_19934,N_19788);
nand U20422 (N_20422,N_19816,N_19830);
and U20423 (N_20423,N_19564,N_19733);
nand U20424 (N_20424,N_19701,N_19981);
nand U20425 (N_20425,N_19768,N_19751);
nor U20426 (N_20426,N_19915,N_19559);
and U20427 (N_20427,N_19619,N_19783);
and U20428 (N_20428,N_19536,N_19898);
nor U20429 (N_20429,N_19733,N_19662);
or U20430 (N_20430,N_19833,N_19834);
nor U20431 (N_20431,N_19730,N_19500);
nor U20432 (N_20432,N_19533,N_19506);
xor U20433 (N_20433,N_19744,N_19962);
xnor U20434 (N_20434,N_19700,N_19621);
nor U20435 (N_20435,N_19855,N_19754);
and U20436 (N_20436,N_19607,N_19996);
and U20437 (N_20437,N_19570,N_19891);
or U20438 (N_20438,N_19924,N_19978);
nand U20439 (N_20439,N_19763,N_19687);
or U20440 (N_20440,N_19915,N_19837);
nor U20441 (N_20441,N_19507,N_19585);
xor U20442 (N_20442,N_19892,N_19642);
xor U20443 (N_20443,N_19754,N_19910);
and U20444 (N_20444,N_19866,N_19618);
or U20445 (N_20445,N_19863,N_19643);
nand U20446 (N_20446,N_19631,N_19978);
nor U20447 (N_20447,N_19597,N_19863);
and U20448 (N_20448,N_19871,N_19603);
nand U20449 (N_20449,N_19701,N_19751);
and U20450 (N_20450,N_19716,N_19847);
nor U20451 (N_20451,N_19706,N_19771);
and U20452 (N_20452,N_19669,N_19959);
nand U20453 (N_20453,N_19563,N_19564);
nand U20454 (N_20454,N_19892,N_19579);
nor U20455 (N_20455,N_19702,N_19580);
nor U20456 (N_20456,N_19848,N_19767);
nor U20457 (N_20457,N_19508,N_19717);
and U20458 (N_20458,N_19598,N_19625);
xor U20459 (N_20459,N_19617,N_19519);
or U20460 (N_20460,N_19581,N_19865);
nor U20461 (N_20461,N_19798,N_19838);
nor U20462 (N_20462,N_19665,N_19697);
xor U20463 (N_20463,N_19999,N_19930);
nor U20464 (N_20464,N_19903,N_19680);
or U20465 (N_20465,N_19858,N_19754);
nor U20466 (N_20466,N_19768,N_19644);
xor U20467 (N_20467,N_19704,N_19665);
nand U20468 (N_20468,N_19841,N_19899);
or U20469 (N_20469,N_19637,N_19777);
or U20470 (N_20470,N_19541,N_19701);
and U20471 (N_20471,N_19540,N_19546);
xnor U20472 (N_20472,N_19738,N_19654);
xor U20473 (N_20473,N_19958,N_19721);
nor U20474 (N_20474,N_19500,N_19660);
or U20475 (N_20475,N_19962,N_19578);
and U20476 (N_20476,N_19942,N_19590);
nand U20477 (N_20477,N_19546,N_19606);
or U20478 (N_20478,N_19659,N_19764);
nor U20479 (N_20479,N_19684,N_19886);
xnor U20480 (N_20480,N_19914,N_19994);
xnor U20481 (N_20481,N_19578,N_19581);
nor U20482 (N_20482,N_19802,N_19551);
xnor U20483 (N_20483,N_19803,N_19796);
nand U20484 (N_20484,N_19697,N_19763);
nor U20485 (N_20485,N_19605,N_19815);
or U20486 (N_20486,N_19700,N_19774);
nor U20487 (N_20487,N_19855,N_19584);
nand U20488 (N_20488,N_19770,N_19690);
xor U20489 (N_20489,N_19752,N_19568);
nor U20490 (N_20490,N_19630,N_19889);
nand U20491 (N_20491,N_19927,N_19964);
nor U20492 (N_20492,N_19802,N_19691);
nand U20493 (N_20493,N_19870,N_19714);
xnor U20494 (N_20494,N_19678,N_19585);
nor U20495 (N_20495,N_19973,N_19532);
nand U20496 (N_20496,N_19686,N_19990);
or U20497 (N_20497,N_19789,N_19635);
xor U20498 (N_20498,N_19982,N_19896);
or U20499 (N_20499,N_19837,N_19865);
nor U20500 (N_20500,N_20062,N_20300);
or U20501 (N_20501,N_20343,N_20056);
nand U20502 (N_20502,N_20184,N_20455);
and U20503 (N_20503,N_20412,N_20360);
and U20504 (N_20504,N_20094,N_20376);
xor U20505 (N_20505,N_20108,N_20086);
nor U20506 (N_20506,N_20043,N_20245);
xnor U20507 (N_20507,N_20117,N_20379);
xor U20508 (N_20508,N_20282,N_20123);
nand U20509 (N_20509,N_20393,N_20491);
nor U20510 (N_20510,N_20220,N_20075);
xnor U20511 (N_20511,N_20232,N_20302);
nor U20512 (N_20512,N_20027,N_20244);
nand U20513 (N_20513,N_20292,N_20210);
nand U20514 (N_20514,N_20110,N_20095);
or U20515 (N_20515,N_20299,N_20364);
and U20516 (N_20516,N_20164,N_20191);
nand U20517 (N_20517,N_20338,N_20207);
and U20518 (N_20518,N_20145,N_20327);
xnor U20519 (N_20519,N_20285,N_20240);
or U20520 (N_20520,N_20028,N_20443);
and U20521 (N_20521,N_20187,N_20355);
or U20522 (N_20522,N_20135,N_20332);
nor U20523 (N_20523,N_20142,N_20259);
xor U20524 (N_20524,N_20146,N_20369);
or U20525 (N_20525,N_20228,N_20406);
nor U20526 (N_20526,N_20494,N_20440);
and U20527 (N_20527,N_20174,N_20474);
nand U20528 (N_20528,N_20417,N_20324);
or U20529 (N_20529,N_20462,N_20144);
nand U20530 (N_20530,N_20169,N_20435);
nor U20531 (N_20531,N_20185,N_20383);
nor U20532 (N_20532,N_20446,N_20141);
or U20533 (N_20533,N_20005,N_20218);
nand U20534 (N_20534,N_20444,N_20290);
nor U20535 (N_20535,N_20463,N_20154);
xor U20536 (N_20536,N_20353,N_20118);
and U20537 (N_20537,N_20140,N_20002);
or U20538 (N_20538,N_20429,N_20033);
nor U20539 (N_20539,N_20466,N_20167);
nor U20540 (N_20540,N_20223,N_20350);
xor U20541 (N_20541,N_20403,N_20480);
and U20542 (N_20542,N_20205,N_20241);
nand U20543 (N_20543,N_20490,N_20298);
nor U20544 (N_20544,N_20226,N_20131);
nand U20545 (N_20545,N_20041,N_20323);
nor U20546 (N_20546,N_20365,N_20199);
and U20547 (N_20547,N_20022,N_20073);
nor U20548 (N_20548,N_20288,N_20105);
xnor U20549 (N_20549,N_20243,N_20196);
nor U20550 (N_20550,N_20030,N_20126);
and U20551 (N_20551,N_20212,N_20251);
or U20552 (N_20552,N_20348,N_20473);
nor U20553 (N_20553,N_20394,N_20032);
xnor U20554 (N_20554,N_20268,N_20049);
xor U20555 (N_20555,N_20470,N_20242);
xnor U20556 (N_20556,N_20414,N_20458);
nor U20557 (N_20557,N_20180,N_20349);
xnor U20558 (N_20558,N_20465,N_20333);
nand U20559 (N_20559,N_20283,N_20279);
nor U20560 (N_20560,N_20267,N_20203);
xor U20561 (N_20561,N_20287,N_20488);
or U20562 (N_20562,N_20224,N_20341);
nand U20563 (N_20563,N_20193,N_20426);
nand U20564 (N_20564,N_20297,N_20265);
or U20565 (N_20565,N_20399,N_20451);
xnor U20566 (N_20566,N_20000,N_20020);
xnor U20567 (N_20567,N_20478,N_20115);
and U20568 (N_20568,N_20270,N_20031);
xor U20569 (N_20569,N_20420,N_20404);
nor U20570 (N_20570,N_20217,N_20254);
and U20571 (N_20571,N_20104,N_20206);
nand U20572 (N_20572,N_20070,N_20239);
or U20573 (N_20573,N_20124,N_20281);
nor U20574 (N_20574,N_20029,N_20371);
and U20575 (N_20575,N_20266,N_20066);
and U20576 (N_20576,N_20401,N_20137);
nor U20577 (N_20577,N_20319,N_20321);
nand U20578 (N_20578,N_20172,N_20485);
or U20579 (N_20579,N_20296,N_20111);
xor U20580 (N_20580,N_20234,N_20256);
nor U20581 (N_20581,N_20192,N_20475);
nand U20582 (N_20582,N_20158,N_20088);
and U20583 (N_20583,N_20069,N_20122);
or U20584 (N_20584,N_20074,N_20246);
nor U20585 (N_20585,N_20015,N_20334);
xor U20586 (N_20586,N_20467,N_20021);
nor U20587 (N_20587,N_20219,N_20114);
nand U20588 (N_20588,N_20099,N_20395);
and U20589 (N_20589,N_20405,N_20004);
or U20590 (N_20590,N_20410,N_20082);
xor U20591 (N_20591,N_20186,N_20389);
xor U20592 (N_20592,N_20061,N_20106);
and U20593 (N_20593,N_20397,N_20222);
xnor U20594 (N_20594,N_20120,N_20042);
and U20595 (N_20595,N_20328,N_20036);
nor U20596 (N_20596,N_20472,N_20498);
nand U20597 (N_20597,N_20316,N_20024);
and U20598 (N_20598,N_20459,N_20358);
nand U20599 (N_20599,N_20482,N_20311);
nand U20600 (N_20600,N_20447,N_20037);
and U20601 (N_20601,N_20149,N_20409);
nand U20602 (N_20602,N_20121,N_20214);
or U20603 (N_20603,N_20047,N_20318);
or U20604 (N_20604,N_20017,N_20384);
and U20605 (N_20605,N_20044,N_20125);
xnor U20606 (N_20606,N_20305,N_20163);
and U20607 (N_20607,N_20059,N_20434);
and U20608 (N_20608,N_20176,N_20381);
and U20609 (N_20609,N_20424,N_20452);
nand U20610 (N_20610,N_20456,N_20178);
and U20611 (N_20611,N_20419,N_20089);
and U20612 (N_20612,N_20018,N_20454);
or U20613 (N_20613,N_20127,N_20077);
or U20614 (N_20614,N_20391,N_20257);
xnor U20615 (N_20615,N_20198,N_20188);
nand U20616 (N_20616,N_20377,N_20116);
and U20617 (N_20617,N_20335,N_20177);
xor U20618 (N_20618,N_20481,N_20008);
or U20619 (N_20619,N_20392,N_20190);
nand U20620 (N_20620,N_20170,N_20157);
nor U20621 (N_20621,N_20211,N_20057);
and U20622 (N_20622,N_20469,N_20293);
and U20623 (N_20623,N_20312,N_20495);
or U20624 (N_20624,N_20003,N_20402);
nor U20625 (N_20625,N_20130,N_20413);
xor U20626 (N_20626,N_20045,N_20442);
or U20627 (N_20627,N_20342,N_20489);
xnor U20628 (N_20628,N_20295,N_20247);
nand U20629 (N_20629,N_20171,N_20215);
nor U20630 (N_20630,N_20119,N_20252);
or U20631 (N_20631,N_20040,N_20237);
and U20632 (N_20632,N_20152,N_20441);
xnor U20633 (N_20633,N_20189,N_20289);
or U20634 (N_20634,N_20109,N_20150);
or U20635 (N_20635,N_20432,N_20079);
nand U20636 (N_20636,N_20204,N_20098);
nand U20637 (N_20637,N_20398,N_20138);
and U20638 (N_20638,N_20453,N_20275);
nor U20639 (N_20639,N_20202,N_20357);
and U20640 (N_20640,N_20320,N_20476);
and U20641 (N_20641,N_20085,N_20361);
nor U20642 (N_20642,N_20197,N_20340);
nor U20643 (N_20643,N_20132,N_20304);
and U20644 (N_20644,N_20483,N_20009);
xnor U20645 (N_20645,N_20097,N_20326);
nand U20646 (N_20646,N_20368,N_20229);
nand U20647 (N_20647,N_20236,N_20448);
nor U20648 (N_20648,N_20183,N_20407);
xor U20649 (N_20649,N_20081,N_20136);
or U20650 (N_20650,N_20133,N_20148);
or U20651 (N_20651,N_20486,N_20165);
xnor U20652 (N_20652,N_20162,N_20306);
or U20653 (N_20653,N_20225,N_20103);
or U20654 (N_20654,N_20011,N_20055);
xnor U20655 (N_20655,N_20034,N_20194);
or U20656 (N_20656,N_20060,N_20261);
nand U20657 (N_20657,N_20416,N_20280);
or U20658 (N_20658,N_20012,N_20050);
xor U20659 (N_20659,N_20013,N_20255);
and U20660 (N_20660,N_20068,N_20449);
and U20661 (N_20661,N_20415,N_20421);
or U20662 (N_20662,N_20496,N_20272);
nand U20663 (N_20663,N_20039,N_20390);
nand U20664 (N_20664,N_20129,N_20425);
or U20665 (N_20665,N_20388,N_20271);
and U20666 (N_20666,N_20273,N_20307);
or U20667 (N_20667,N_20195,N_20262);
and U20668 (N_20668,N_20484,N_20301);
nor U20669 (N_20669,N_20336,N_20385);
or U20670 (N_20670,N_20227,N_20291);
nand U20671 (N_20671,N_20209,N_20064);
and U20672 (N_20672,N_20235,N_20303);
nor U20673 (N_20673,N_20433,N_20208);
and U20674 (N_20674,N_20309,N_20411);
nor U20675 (N_20675,N_20260,N_20200);
nand U20676 (N_20676,N_20084,N_20160);
or U20677 (N_20677,N_20352,N_20370);
xor U20678 (N_20678,N_20155,N_20052);
or U20679 (N_20679,N_20372,N_20366);
nor U20680 (N_20680,N_20418,N_20233);
xor U20681 (N_20681,N_20181,N_20007);
nor U20682 (N_20682,N_20436,N_20354);
and U20683 (N_20683,N_20038,N_20010);
and U20684 (N_20684,N_20487,N_20026);
or U20685 (N_20685,N_20048,N_20249);
or U20686 (N_20686,N_20499,N_20035);
xnor U20687 (N_20687,N_20173,N_20100);
and U20688 (N_20688,N_20386,N_20083);
xnor U20689 (N_20689,N_20310,N_20294);
nor U20690 (N_20690,N_20445,N_20263);
or U20691 (N_20691,N_20277,N_20367);
nor U20692 (N_20692,N_20065,N_20380);
and U20693 (N_20693,N_20213,N_20479);
nand U20694 (N_20694,N_20096,N_20438);
or U20695 (N_20695,N_20450,N_20317);
and U20696 (N_20696,N_20166,N_20477);
xnor U20697 (N_20697,N_20468,N_20063);
nor U20698 (N_20698,N_20457,N_20153);
xnor U20699 (N_20699,N_20087,N_20308);
and U20700 (N_20700,N_20238,N_20019);
nor U20701 (N_20701,N_20359,N_20216);
or U20702 (N_20702,N_20351,N_20253);
nor U20703 (N_20703,N_20315,N_20387);
or U20704 (N_20704,N_20101,N_20014);
nand U20705 (N_20705,N_20072,N_20471);
or U20706 (N_20706,N_20400,N_20378);
xor U20707 (N_20707,N_20461,N_20313);
and U20708 (N_20708,N_20071,N_20314);
nor U20709 (N_20709,N_20330,N_20025);
or U20710 (N_20710,N_20113,N_20179);
nor U20711 (N_20711,N_20151,N_20058);
nor U20712 (N_20712,N_20016,N_20076);
and U20713 (N_20713,N_20382,N_20339);
xnor U20714 (N_20714,N_20182,N_20363);
xor U20715 (N_20715,N_20344,N_20258);
xor U20716 (N_20716,N_20346,N_20437);
or U20717 (N_20717,N_20428,N_20345);
nor U20718 (N_20718,N_20337,N_20001);
and U20719 (N_20719,N_20067,N_20046);
or U20720 (N_20720,N_20325,N_20373);
or U20721 (N_20721,N_20143,N_20147);
nand U20722 (N_20722,N_20134,N_20139);
xnor U20723 (N_20723,N_20269,N_20053);
nor U20724 (N_20724,N_20460,N_20286);
and U20725 (N_20725,N_20156,N_20090);
nor U20726 (N_20726,N_20248,N_20102);
or U20727 (N_20727,N_20493,N_20284);
nor U20728 (N_20728,N_20175,N_20159);
nor U20729 (N_20729,N_20128,N_20006);
nand U20730 (N_20730,N_20264,N_20408);
nand U20731 (N_20731,N_20464,N_20331);
nand U20732 (N_20732,N_20168,N_20497);
nand U20733 (N_20733,N_20051,N_20250);
nand U20734 (N_20734,N_20107,N_20430);
or U20735 (N_20735,N_20439,N_20278);
nor U20736 (N_20736,N_20322,N_20092);
nor U20737 (N_20737,N_20080,N_20422);
xor U20738 (N_20738,N_20274,N_20201);
xnor U20739 (N_20739,N_20362,N_20374);
or U20740 (N_20740,N_20054,N_20091);
and U20741 (N_20741,N_20347,N_20276);
nor U20742 (N_20742,N_20221,N_20023);
and U20743 (N_20743,N_20396,N_20161);
nor U20744 (N_20744,N_20356,N_20231);
nor U20745 (N_20745,N_20423,N_20427);
xnor U20746 (N_20746,N_20112,N_20375);
nand U20747 (N_20747,N_20492,N_20431);
nor U20748 (N_20748,N_20078,N_20230);
nand U20749 (N_20749,N_20093,N_20329);
nor U20750 (N_20750,N_20117,N_20235);
and U20751 (N_20751,N_20156,N_20327);
nor U20752 (N_20752,N_20150,N_20265);
nand U20753 (N_20753,N_20401,N_20419);
nor U20754 (N_20754,N_20499,N_20406);
and U20755 (N_20755,N_20051,N_20392);
nand U20756 (N_20756,N_20307,N_20209);
xnor U20757 (N_20757,N_20474,N_20300);
xnor U20758 (N_20758,N_20334,N_20499);
xnor U20759 (N_20759,N_20000,N_20230);
xor U20760 (N_20760,N_20098,N_20062);
nand U20761 (N_20761,N_20157,N_20478);
or U20762 (N_20762,N_20003,N_20008);
or U20763 (N_20763,N_20137,N_20490);
or U20764 (N_20764,N_20124,N_20399);
and U20765 (N_20765,N_20240,N_20210);
nand U20766 (N_20766,N_20050,N_20299);
xnor U20767 (N_20767,N_20418,N_20253);
nor U20768 (N_20768,N_20485,N_20400);
and U20769 (N_20769,N_20469,N_20004);
and U20770 (N_20770,N_20296,N_20090);
and U20771 (N_20771,N_20359,N_20349);
or U20772 (N_20772,N_20000,N_20067);
or U20773 (N_20773,N_20408,N_20020);
xnor U20774 (N_20774,N_20359,N_20345);
xnor U20775 (N_20775,N_20005,N_20205);
nand U20776 (N_20776,N_20458,N_20473);
xor U20777 (N_20777,N_20472,N_20257);
nand U20778 (N_20778,N_20132,N_20038);
xor U20779 (N_20779,N_20108,N_20065);
nor U20780 (N_20780,N_20300,N_20448);
xor U20781 (N_20781,N_20183,N_20456);
nor U20782 (N_20782,N_20475,N_20265);
nand U20783 (N_20783,N_20349,N_20287);
and U20784 (N_20784,N_20227,N_20238);
and U20785 (N_20785,N_20235,N_20484);
xor U20786 (N_20786,N_20184,N_20284);
nand U20787 (N_20787,N_20201,N_20378);
or U20788 (N_20788,N_20215,N_20404);
nand U20789 (N_20789,N_20001,N_20053);
nand U20790 (N_20790,N_20469,N_20384);
or U20791 (N_20791,N_20134,N_20319);
and U20792 (N_20792,N_20251,N_20196);
or U20793 (N_20793,N_20411,N_20174);
xor U20794 (N_20794,N_20166,N_20258);
or U20795 (N_20795,N_20333,N_20267);
or U20796 (N_20796,N_20442,N_20203);
nor U20797 (N_20797,N_20382,N_20350);
xnor U20798 (N_20798,N_20487,N_20099);
and U20799 (N_20799,N_20280,N_20312);
and U20800 (N_20800,N_20493,N_20422);
nor U20801 (N_20801,N_20437,N_20355);
nand U20802 (N_20802,N_20031,N_20084);
or U20803 (N_20803,N_20404,N_20103);
and U20804 (N_20804,N_20491,N_20010);
xor U20805 (N_20805,N_20317,N_20300);
and U20806 (N_20806,N_20217,N_20224);
or U20807 (N_20807,N_20367,N_20279);
nand U20808 (N_20808,N_20233,N_20309);
nor U20809 (N_20809,N_20183,N_20486);
nand U20810 (N_20810,N_20011,N_20102);
xnor U20811 (N_20811,N_20467,N_20290);
nand U20812 (N_20812,N_20016,N_20273);
nor U20813 (N_20813,N_20002,N_20032);
and U20814 (N_20814,N_20110,N_20216);
nand U20815 (N_20815,N_20487,N_20335);
nor U20816 (N_20816,N_20070,N_20476);
or U20817 (N_20817,N_20464,N_20061);
nand U20818 (N_20818,N_20021,N_20346);
or U20819 (N_20819,N_20405,N_20062);
xnor U20820 (N_20820,N_20098,N_20358);
xor U20821 (N_20821,N_20228,N_20399);
nor U20822 (N_20822,N_20351,N_20270);
nor U20823 (N_20823,N_20210,N_20023);
or U20824 (N_20824,N_20125,N_20370);
or U20825 (N_20825,N_20366,N_20085);
nand U20826 (N_20826,N_20304,N_20103);
xor U20827 (N_20827,N_20237,N_20112);
nand U20828 (N_20828,N_20011,N_20156);
and U20829 (N_20829,N_20119,N_20175);
xnor U20830 (N_20830,N_20229,N_20461);
or U20831 (N_20831,N_20044,N_20472);
and U20832 (N_20832,N_20459,N_20247);
nor U20833 (N_20833,N_20149,N_20290);
nand U20834 (N_20834,N_20134,N_20349);
nand U20835 (N_20835,N_20426,N_20162);
nor U20836 (N_20836,N_20368,N_20079);
nand U20837 (N_20837,N_20394,N_20010);
or U20838 (N_20838,N_20423,N_20394);
xor U20839 (N_20839,N_20216,N_20149);
nor U20840 (N_20840,N_20479,N_20391);
nand U20841 (N_20841,N_20100,N_20176);
and U20842 (N_20842,N_20015,N_20133);
nand U20843 (N_20843,N_20421,N_20408);
xor U20844 (N_20844,N_20221,N_20109);
nor U20845 (N_20845,N_20246,N_20101);
nor U20846 (N_20846,N_20411,N_20216);
or U20847 (N_20847,N_20240,N_20374);
xor U20848 (N_20848,N_20203,N_20126);
and U20849 (N_20849,N_20397,N_20059);
or U20850 (N_20850,N_20330,N_20351);
or U20851 (N_20851,N_20046,N_20038);
xnor U20852 (N_20852,N_20094,N_20385);
nor U20853 (N_20853,N_20447,N_20141);
nand U20854 (N_20854,N_20310,N_20089);
nor U20855 (N_20855,N_20225,N_20300);
nand U20856 (N_20856,N_20130,N_20208);
xnor U20857 (N_20857,N_20426,N_20424);
nand U20858 (N_20858,N_20413,N_20007);
nand U20859 (N_20859,N_20160,N_20478);
xnor U20860 (N_20860,N_20263,N_20024);
nor U20861 (N_20861,N_20485,N_20071);
or U20862 (N_20862,N_20174,N_20245);
xor U20863 (N_20863,N_20356,N_20379);
nand U20864 (N_20864,N_20485,N_20022);
xor U20865 (N_20865,N_20176,N_20236);
and U20866 (N_20866,N_20212,N_20482);
xnor U20867 (N_20867,N_20412,N_20210);
and U20868 (N_20868,N_20222,N_20171);
nand U20869 (N_20869,N_20402,N_20322);
nor U20870 (N_20870,N_20199,N_20137);
nor U20871 (N_20871,N_20034,N_20010);
xor U20872 (N_20872,N_20044,N_20387);
or U20873 (N_20873,N_20101,N_20028);
or U20874 (N_20874,N_20101,N_20031);
or U20875 (N_20875,N_20446,N_20186);
xnor U20876 (N_20876,N_20349,N_20209);
or U20877 (N_20877,N_20288,N_20085);
and U20878 (N_20878,N_20377,N_20162);
nand U20879 (N_20879,N_20127,N_20160);
nor U20880 (N_20880,N_20103,N_20167);
or U20881 (N_20881,N_20295,N_20042);
xnor U20882 (N_20882,N_20118,N_20263);
xor U20883 (N_20883,N_20486,N_20356);
and U20884 (N_20884,N_20330,N_20188);
nand U20885 (N_20885,N_20351,N_20288);
or U20886 (N_20886,N_20195,N_20145);
nor U20887 (N_20887,N_20398,N_20048);
and U20888 (N_20888,N_20443,N_20452);
or U20889 (N_20889,N_20255,N_20306);
nor U20890 (N_20890,N_20143,N_20005);
and U20891 (N_20891,N_20165,N_20441);
xnor U20892 (N_20892,N_20100,N_20429);
nand U20893 (N_20893,N_20395,N_20306);
or U20894 (N_20894,N_20268,N_20255);
or U20895 (N_20895,N_20250,N_20391);
nor U20896 (N_20896,N_20402,N_20397);
and U20897 (N_20897,N_20230,N_20142);
and U20898 (N_20898,N_20399,N_20179);
xor U20899 (N_20899,N_20211,N_20447);
and U20900 (N_20900,N_20123,N_20483);
nand U20901 (N_20901,N_20474,N_20211);
nor U20902 (N_20902,N_20153,N_20005);
nand U20903 (N_20903,N_20017,N_20471);
nand U20904 (N_20904,N_20487,N_20361);
or U20905 (N_20905,N_20310,N_20109);
and U20906 (N_20906,N_20388,N_20134);
nand U20907 (N_20907,N_20257,N_20445);
and U20908 (N_20908,N_20212,N_20492);
xnor U20909 (N_20909,N_20101,N_20382);
and U20910 (N_20910,N_20257,N_20166);
or U20911 (N_20911,N_20260,N_20373);
nand U20912 (N_20912,N_20051,N_20076);
or U20913 (N_20913,N_20349,N_20272);
or U20914 (N_20914,N_20332,N_20492);
or U20915 (N_20915,N_20475,N_20198);
nor U20916 (N_20916,N_20381,N_20067);
xnor U20917 (N_20917,N_20442,N_20087);
and U20918 (N_20918,N_20337,N_20487);
and U20919 (N_20919,N_20350,N_20369);
nand U20920 (N_20920,N_20184,N_20012);
and U20921 (N_20921,N_20436,N_20384);
nor U20922 (N_20922,N_20154,N_20281);
or U20923 (N_20923,N_20128,N_20330);
nand U20924 (N_20924,N_20464,N_20242);
xnor U20925 (N_20925,N_20073,N_20160);
and U20926 (N_20926,N_20410,N_20313);
nand U20927 (N_20927,N_20376,N_20059);
nand U20928 (N_20928,N_20151,N_20251);
and U20929 (N_20929,N_20097,N_20005);
xor U20930 (N_20930,N_20044,N_20460);
xnor U20931 (N_20931,N_20172,N_20255);
and U20932 (N_20932,N_20203,N_20288);
xnor U20933 (N_20933,N_20491,N_20215);
and U20934 (N_20934,N_20053,N_20228);
xnor U20935 (N_20935,N_20282,N_20140);
and U20936 (N_20936,N_20172,N_20446);
nor U20937 (N_20937,N_20145,N_20258);
and U20938 (N_20938,N_20088,N_20199);
xor U20939 (N_20939,N_20364,N_20212);
nor U20940 (N_20940,N_20112,N_20055);
nor U20941 (N_20941,N_20079,N_20033);
or U20942 (N_20942,N_20154,N_20058);
nand U20943 (N_20943,N_20475,N_20006);
nor U20944 (N_20944,N_20394,N_20338);
nor U20945 (N_20945,N_20139,N_20316);
nor U20946 (N_20946,N_20392,N_20450);
nor U20947 (N_20947,N_20116,N_20130);
and U20948 (N_20948,N_20473,N_20387);
nor U20949 (N_20949,N_20106,N_20022);
xnor U20950 (N_20950,N_20420,N_20479);
nor U20951 (N_20951,N_20152,N_20151);
or U20952 (N_20952,N_20438,N_20281);
nor U20953 (N_20953,N_20128,N_20197);
nand U20954 (N_20954,N_20482,N_20131);
xor U20955 (N_20955,N_20073,N_20067);
nand U20956 (N_20956,N_20261,N_20292);
and U20957 (N_20957,N_20220,N_20479);
nor U20958 (N_20958,N_20104,N_20258);
or U20959 (N_20959,N_20235,N_20126);
or U20960 (N_20960,N_20274,N_20437);
nor U20961 (N_20961,N_20403,N_20088);
or U20962 (N_20962,N_20336,N_20018);
nand U20963 (N_20963,N_20176,N_20459);
and U20964 (N_20964,N_20434,N_20370);
or U20965 (N_20965,N_20243,N_20427);
or U20966 (N_20966,N_20012,N_20212);
xor U20967 (N_20967,N_20140,N_20042);
nand U20968 (N_20968,N_20380,N_20283);
nor U20969 (N_20969,N_20233,N_20166);
nand U20970 (N_20970,N_20095,N_20254);
nand U20971 (N_20971,N_20431,N_20225);
or U20972 (N_20972,N_20096,N_20481);
xnor U20973 (N_20973,N_20071,N_20045);
xor U20974 (N_20974,N_20150,N_20374);
nand U20975 (N_20975,N_20464,N_20179);
and U20976 (N_20976,N_20137,N_20449);
xor U20977 (N_20977,N_20183,N_20312);
nor U20978 (N_20978,N_20188,N_20116);
and U20979 (N_20979,N_20057,N_20466);
and U20980 (N_20980,N_20315,N_20076);
nand U20981 (N_20981,N_20464,N_20334);
or U20982 (N_20982,N_20207,N_20356);
nand U20983 (N_20983,N_20047,N_20210);
xnor U20984 (N_20984,N_20282,N_20409);
nor U20985 (N_20985,N_20133,N_20489);
xor U20986 (N_20986,N_20467,N_20454);
xnor U20987 (N_20987,N_20222,N_20201);
nor U20988 (N_20988,N_20078,N_20131);
nand U20989 (N_20989,N_20100,N_20023);
and U20990 (N_20990,N_20202,N_20377);
and U20991 (N_20991,N_20375,N_20377);
xor U20992 (N_20992,N_20361,N_20175);
or U20993 (N_20993,N_20026,N_20019);
xnor U20994 (N_20994,N_20395,N_20105);
or U20995 (N_20995,N_20299,N_20097);
nand U20996 (N_20996,N_20224,N_20293);
nor U20997 (N_20997,N_20373,N_20181);
nor U20998 (N_20998,N_20296,N_20285);
or U20999 (N_20999,N_20224,N_20455);
or U21000 (N_21000,N_20612,N_20790);
or U21001 (N_21001,N_20582,N_20560);
and U21002 (N_21002,N_20845,N_20822);
xnor U21003 (N_21003,N_20562,N_20633);
and U21004 (N_21004,N_20974,N_20975);
or U21005 (N_21005,N_20777,N_20594);
nor U21006 (N_21006,N_20662,N_20933);
nor U21007 (N_21007,N_20892,N_20963);
xor U21008 (N_21008,N_20574,N_20957);
xor U21009 (N_21009,N_20593,N_20720);
or U21010 (N_21010,N_20508,N_20919);
nor U21011 (N_21011,N_20638,N_20561);
and U21012 (N_21012,N_20616,N_20819);
and U21013 (N_21013,N_20799,N_20710);
nand U21014 (N_21014,N_20903,N_20642);
and U21015 (N_21015,N_20726,N_20770);
and U21016 (N_21016,N_20967,N_20526);
nor U21017 (N_21017,N_20838,N_20865);
and U21018 (N_21018,N_20929,N_20745);
and U21019 (N_21019,N_20983,N_20960);
xnor U21020 (N_21020,N_20917,N_20698);
nand U21021 (N_21021,N_20961,N_20940);
nand U21022 (N_21022,N_20518,N_20944);
and U21023 (N_21023,N_20655,N_20935);
xor U21024 (N_21024,N_20922,N_20876);
nand U21025 (N_21025,N_20839,N_20849);
or U21026 (N_21026,N_20636,N_20817);
xnor U21027 (N_21027,N_20846,N_20816);
xnor U21028 (N_21028,N_20718,N_20524);
or U21029 (N_21029,N_20614,N_20528);
xor U21030 (N_21030,N_20567,N_20559);
nand U21031 (N_21031,N_20910,N_20990);
nor U21032 (N_21032,N_20600,N_20856);
nor U21033 (N_21033,N_20527,N_20908);
xor U21034 (N_21034,N_20690,N_20580);
xor U21035 (N_21035,N_20533,N_20679);
xnor U21036 (N_21036,N_20926,N_20753);
nand U21037 (N_21037,N_20982,N_20999);
nor U21038 (N_21038,N_20854,N_20813);
nor U21039 (N_21039,N_20937,N_20557);
and U21040 (N_21040,N_20714,N_20936);
nand U21041 (N_21041,N_20664,N_20667);
xor U21042 (N_21042,N_20723,N_20644);
nand U21043 (N_21043,N_20500,N_20599);
or U21044 (N_21044,N_20611,N_20871);
or U21045 (N_21045,N_20847,N_20850);
nand U21046 (N_21046,N_20551,N_20877);
nand U21047 (N_21047,N_20881,N_20731);
nand U21048 (N_21048,N_20860,N_20661);
nand U21049 (N_21049,N_20716,N_20568);
nor U21050 (N_21050,N_20652,N_20949);
xor U21051 (N_21051,N_20989,N_20758);
xnor U21052 (N_21052,N_20907,N_20658);
nor U21053 (N_21053,N_20870,N_20793);
xnor U21054 (N_21054,N_20747,N_20890);
and U21055 (N_21055,N_20992,N_20824);
nand U21056 (N_21056,N_20730,N_20520);
and U21057 (N_21057,N_20738,N_20687);
and U21058 (N_21058,N_20986,N_20680);
nor U21059 (N_21059,N_20515,N_20646);
or U21060 (N_21060,N_20981,N_20853);
or U21061 (N_21061,N_20739,N_20634);
nand U21062 (N_21062,N_20618,N_20809);
xnor U21063 (N_21063,N_20620,N_20621);
xor U21064 (N_21064,N_20529,N_20884);
and U21065 (N_21065,N_20828,N_20615);
or U21066 (N_21066,N_20588,N_20746);
nor U21067 (N_21067,N_20796,N_20898);
nand U21068 (N_21068,N_20915,N_20744);
nand U21069 (N_21069,N_20886,N_20894);
or U21070 (N_21070,N_20976,N_20649);
nand U21071 (N_21071,N_20872,N_20647);
nand U21072 (N_21072,N_20566,N_20706);
nor U21073 (N_21073,N_20888,N_20656);
nand U21074 (N_21074,N_20752,N_20810);
xor U21075 (N_21075,N_20959,N_20887);
xnor U21076 (N_21076,N_20665,N_20504);
xor U21077 (N_21077,N_20998,N_20815);
and U21078 (N_21078,N_20630,N_20556);
xor U21079 (N_21079,N_20546,N_20639);
xor U21080 (N_21080,N_20604,N_20765);
nand U21081 (N_21081,N_20727,N_20626);
xnor U21082 (N_21082,N_20991,N_20570);
or U21083 (N_21083,N_20812,N_20941);
and U21084 (N_21084,N_20757,N_20781);
and U21085 (N_21085,N_20945,N_20558);
xor U21086 (N_21086,N_20724,N_20563);
and U21087 (N_21087,N_20993,N_20525);
nand U21088 (N_21088,N_20632,N_20767);
nand U21089 (N_21089,N_20843,N_20754);
nand U21090 (N_21090,N_20509,N_20764);
nand U21091 (N_21091,N_20923,N_20831);
or U21092 (N_21092,N_20885,N_20947);
and U21093 (N_21093,N_20789,N_20514);
nor U21094 (N_21094,N_20977,N_20841);
or U21095 (N_21095,N_20659,N_20713);
xnor U21096 (N_21096,N_20925,N_20891);
or U21097 (N_21097,N_20674,N_20958);
nand U21098 (N_21098,N_20511,N_20997);
nand U21099 (N_21099,N_20503,N_20741);
xnor U21100 (N_21100,N_20984,N_20603);
and U21101 (N_21101,N_20875,N_20700);
nand U21102 (N_21102,N_20994,N_20802);
and U21103 (N_21103,N_20932,N_20590);
nor U21104 (N_21104,N_20797,N_20507);
and U21105 (N_21105,N_20717,N_20712);
nor U21106 (N_21106,N_20804,N_20857);
xor U21107 (N_21107,N_20607,N_20651);
or U21108 (N_21108,N_20787,N_20948);
and U21109 (N_21109,N_20609,N_20592);
or U21110 (N_21110,N_20707,N_20627);
nor U21111 (N_21111,N_20668,N_20800);
nor U21112 (N_21112,N_20595,N_20697);
nand U21113 (N_21113,N_20985,N_20641);
nor U21114 (N_21114,N_20534,N_20942);
xnor U21115 (N_21115,N_20517,N_20904);
or U21116 (N_21116,N_20541,N_20808);
nand U21117 (N_21117,N_20805,N_20766);
nand U21118 (N_21118,N_20788,N_20965);
and U21119 (N_21119,N_20951,N_20749);
or U21120 (N_21120,N_20869,N_20598);
nand U21121 (N_21121,N_20553,N_20863);
nand U21122 (N_21122,N_20597,N_20729);
nand U21123 (N_21123,N_20859,N_20848);
or U21124 (N_21124,N_20814,N_20768);
nor U21125 (N_21125,N_20613,N_20708);
xor U21126 (N_21126,N_20535,N_20775);
nor U21127 (N_21127,N_20950,N_20868);
and U21128 (N_21128,N_20791,N_20979);
and U21129 (N_21129,N_20513,N_20676);
xnor U21130 (N_21130,N_20905,N_20643);
or U21131 (N_21131,N_20601,N_20693);
xnor U21132 (N_21132,N_20801,N_20873);
nor U21133 (N_21133,N_20778,N_20893);
nand U21134 (N_21134,N_20895,N_20677);
nand U21135 (N_21135,N_20798,N_20773);
nor U21136 (N_21136,N_20913,N_20931);
nor U21137 (N_21137,N_20896,N_20874);
nand U21138 (N_21138,N_20722,N_20970);
or U21139 (N_21139,N_20930,N_20579);
nor U21140 (N_21140,N_20692,N_20617);
nor U21141 (N_21141,N_20521,N_20995);
nor U21142 (N_21142,N_20756,N_20540);
xor U21143 (N_21143,N_20988,N_20996);
nor U21144 (N_21144,N_20519,N_20537);
xnor U21145 (N_21145,N_20751,N_20939);
or U21146 (N_21146,N_20653,N_20637);
and U21147 (N_21147,N_20571,N_20512);
and U21148 (N_21148,N_20682,N_20625);
xnor U21149 (N_21149,N_20699,N_20840);
xnor U21150 (N_21150,N_20530,N_20762);
nand U21151 (N_21151,N_20502,N_20946);
xnor U21152 (N_21152,N_20704,N_20811);
nor U21153 (N_21153,N_20901,N_20830);
xnor U21154 (N_21154,N_20702,N_20596);
or U21155 (N_21155,N_20532,N_20782);
nand U21156 (N_21156,N_20629,N_20681);
nand U21157 (N_21157,N_20779,N_20971);
xor U21158 (N_21158,N_20759,N_20536);
nor U21159 (N_21159,N_20867,N_20964);
or U21160 (N_21160,N_20921,N_20861);
nand U21161 (N_21161,N_20862,N_20721);
or U21162 (N_21162,N_20835,N_20978);
or U21163 (N_21163,N_20924,N_20663);
nand U21164 (N_21164,N_20539,N_20882);
and U21165 (N_21165,N_20866,N_20624);
nand U21166 (N_21166,N_20550,N_20962);
nor U21167 (N_21167,N_20672,N_20750);
xor U21168 (N_21168,N_20542,N_20523);
nor U21169 (N_21169,N_20780,N_20623);
xnor U21170 (N_21170,N_20719,N_20736);
xor U21171 (N_21171,N_20705,N_20578);
and U21172 (N_21172,N_20934,N_20807);
and U21173 (N_21173,N_20826,N_20569);
and U21174 (N_21174,N_20734,N_20952);
and U21175 (N_21175,N_20538,N_20585);
nor U21176 (N_21176,N_20640,N_20825);
or U21177 (N_21177,N_20784,N_20694);
and U21178 (N_21178,N_20654,N_20968);
xor U21179 (N_21179,N_20920,N_20956);
or U21180 (N_21180,N_20648,N_20555);
or U21181 (N_21181,N_20545,N_20575);
and U21182 (N_21182,N_20696,N_20883);
nand U21183 (N_21183,N_20688,N_20691);
and U21184 (N_21184,N_20549,N_20842);
or U21185 (N_21185,N_20733,N_20880);
nand U21186 (N_21186,N_20827,N_20670);
nand U21187 (N_21187,N_20878,N_20619);
and U21188 (N_21188,N_20836,N_20683);
xor U21189 (N_21189,N_20685,N_20743);
and U21190 (N_21190,N_20973,N_20844);
nor U21191 (N_21191,N_20610,N_20628);
and U21192 (N_21192,N_20581,N_20548);
xnor U21193 (N_21193,N_20760,N_20954);
or U21194 (N_21194,N_20605,N_20879);
nand U21195 (N_21195,N_20927,N_20742);
xnor U21196 (N_21196,N_20669,N_20889);
nand U21197 (N_21197,N_20689,N_20980);
nor U21198 (N_21198,N_20715,N_20510);
xor U21199 (N_21199,N_20833,N_20916);
or U21200 (N_21200,N_20602,N_20820);
nand U21201 (N_21201,N_20666,N_20506);
nand U21202 (N_21202,N_20587,N_20684);
xor U21203 (N_21203,N_20650,N_20783);
nand U21204 (N_21204,N_20928,N_20823);
nand U21205 (N_21205,N_20899,N_20645);
nand U21206 (N_21206,N_20591,N_20606);
nand U21207 (N_21207,N_20794,N_20740);
nand U21208 (N_21208,N_20858,N_20755);
nor U21209 (N_21209,N_20725,N_20852);
xnor U21210 (N_21210,N_20748,N_20586);
nand U21211 (N_21211,N_20786,N_20912);
nand U21212 (N_21212,N_20732,N_20834);
and U21213 (N_21213,N_20911,N_20675);
xor U21214 (N_21214,N_20806,N_20953);
nand U21215 (N_21215,N_20564,N_20505);
xor U21216 (N_21216,N_20583,N_20552);
and U21217 (N_21217,N_20671,N_20776);
xnor U21218 (N_21218,N_20686,N_20774);
xnor U21219 (N_21219,N_20711,N_20544);
and U21220 (N_21220,N_20703,N_20829);
nor U21221 (N_21221,N_20821,N_20897);
nor U21222 (N_21222,N_20554,N_20772);
or U21223 (N_21223,N_20673,N_20622);
nor U21224 (N_21224,N_20966,N_20576);
nand U21225 (N_21225,N_20516,N_20631);
xnor U21226 (N_21226,N_20635,N_20577);
and U21227 (N_21227,N_20972,N_20589);
xnor U21228 (N_21228,N_20660,N_20761);
and U21229 (N_21229,N_20573,N_20501);
or U21230 (N_21230,N_20769,N_20522);
nor U21231 (N_21231,N_20864,N_20695);
nand U21232 (N_21232,N_20906,N_20735);
nor U21233 (N_21233,N_20531,N_20572);
nor U21234 (N_21234,N_20771,N_20543);
nand U21235 (N_21235,N_20678,N_20837);
xnor U21236 (N_21236,N_20584,N_20608);
xnor U21237 (N_21237,N_20938,N_20737);
nor U21238 (N_21238,N_20763,N_20900);
nand U21239 (N_21239,N_20728,N_20943);
or U21240 (N_21240,N_20709,N_20795);
xor U21241 (N_21241,N_20701,N_20855);
nor U21242 (N_21242,N_20792,N_20832);
nand U21243 (N_21243,N_20565,N_20987);
nor U21244 (N_21244,N_20803,N_20914);
and U21245 (N_21245,N_20851,N_20955);
or U21246 (N_21246,N_20547,N_20969);
nor U21247 (N_21247,N_20818,N_20909);
xnor U21248 (N_21248,N_20785,N_20902);
xor U21249 (N_21249,N_20657,N_20918);
or U21250 (N_21250,N_20759,N_20535);
xnor U21251 (N_21251,N_20901,N_20788);
xor U21252 (N_21252,N_20990,N_20844);
and U21253 (N_21253,N_20936,N_20713);
or U21254 (N_21254,N_20951,N_20935);
and U21255 (N_21255,N_20949,N_20809);
xnor U21256 (N_21256,N_20989,N_20994);
nor U21257 (N_21257,N_20845,N_20745);
and U21258 (N_21258,N_20806,N_20848);
or U21259 (N_21259,N_20757,N_20811);
xor U21260 (N_21260,N_20571,N_20681);
nand U21261 (N_21261,N_20922,N_20869);
or U21262 (N_21262,N_20749,N_20636);
and U21263 (N_21263,N_20881,N_20598);
and U21264 (N_21264,N_20873,N_20655);
nor U21265 (N_21265,N_20983,N_20921);
xnor U21266 (N_21266,N_20749,N_20799);
and U21267 (N_21267,N_20728,N_20964);
or U21268 (N_21268,N_20945,N_20798);
and U21269 (N_21269,N_20694,N_20873);
or U21270 (N_21270,N_20946,N_20741);
or U21271 (N_21271,N_20936,N_20938);
nand U21272 (N_21272,N_20840,N_20737);
or U21273 (N_21273,N_20968,N_20922);
xnor U21274 (N_21274,N_20888,N_20646);
nor U21275 (N_21275,N_20769,N_20630);
nand U21276 (N_21276,N_20538,N_20586);
xor U21277 (N_21277,N_20825,N_20633);
xnor U21278 (N_21278,N_20862,N_20516);
nand U21279 (N_21279,N_20877,N_20893);
or U21280 (N_21280,N_20930,N_20578);
xnor U21281 (N_21281,N_20979,N_20881);
nor U21282 (N_21282,N_20848,N_20964);
xor U21283 (N_21283,N_20705,N_20783);
xor U21284 (N_21284,N_20657,N_20835);
and U21285 (N_21285,N_20599,N_20756);
nor U21286 (N_21286,N_20988,N_20937);
nor U21287 (N_21287,N_20610,N_20869);
nor U21288 (N_21288,N_20642,N_20913);
and U21289 (N_21289,N_20896,N_20891);
or U21290 (N_21290,N_20862,N_20822);
or U21291 (N_21291,N_20942,N_20889);
or U21292 (N_21292,N_20614,N_20604);
nand U21293 (N_21293,N_20727,N_20565);
xor U21294 (N_21294,N_20864,N_20947);
or U21295 (N_21295,N_20936,N_20799);
nor U21296 (N_21296,N_20682,N_20911);
or U21297 (N_21297,N_20599,N_20921);
or U21298 (N_21298,N_20735,N_20956);
or U21299 (N_21299,N_20505,N_20622);
or U21300 (N_21300,N_20587,N_20995);
and U21301 (N_21301,N_20813,N_20845);
or U21302 (N_21302,N_20665,N_20687);
nand U21303 (N_21303,N_20685,N_20581);
xor U21304 (N_21304,N_20825,N_20947);
nor U21305 (N_21305,N_20818,N_20788);
nor U21306 (N_21306,N_20577,N_20721);
or U21307 (N_21307,N_20805,N_20901);
or U21308 (N_21308,N_20764,N_20506);
nor U21309 (N_21309,N_20749,N_20507);
or U21310 (N_21310,N_20569,N_20783);
nand U21311 (N_21311,N_20880,N_20526);
nor U21312 (N_21312,N_20844,N_20619);
or U21313 (N_21313,N_20681,N_20646);
xnor U21314 (N_21314,N_20677,N_20891);
nand U21315 (N_21315,N_20554,N_20882);
nor U21316 (N_21316,N_20749,N_20940);
and U21317 (N_21317,N_20500,N_20671);
or U21318 (N_21318,N_20587,N_20827);
or U21319 (N_21319,N_20525,N_20606);
nand U21320 (N_21320,N_20736,N_20548);
and U21321 (N_21321,N_20515,N_20845);
nand U21322 (N_21322,N_20614,N_20616);
nand U21323 (N_21323,N_20538,N_20799);
or U21324 (N_21324,N_20629,N_20730);
and U21325 (N_21325,N_20693,N_20699);
nor U21326 (N_21326,N_20993,N_20602);
xnor U21327 (N_21327,N_20676,N_20930);
nor U21328 (N_21328,N_20918,N_20577);
or U21329 (N_21329,N_20971,N_20703);
xnor U21330 (N_21330,N_20678,N_20967);
and U21331 (N_21331,N_20761,N_20945);
xor U21332 (N_21332,N_20965,N_20943);
and U21333 (N_21333,N_20887,N_20705);
and U21334 (N_21334,N_20992,N_20709);
xor U21335 (N_21335,N_20790,N_20510);
or U21336 (N_21336,N_20531,N_20578);
and U21337 (N_21337,N_20985,N_20963);
nand U21338 (N_21338,N_20616,N_20579);
nand U21339 (N_21339,N_20720,N_20841);
or U21340 (N_21340,N_20563,N_20675);
nor U21341 (N_21341,N_20791,N_20803);
and U21342 (N_21342,N_20973,N_20871);
or U21343 (N_21343,N_20719,N_20543);
nor U21344 (N_21344,N_20634,N_20662);
xor U21345 (N_21345,N_20946,N_20593);
and U21346 (N_21346,N_20976,N_20746);
xnor U21347 (N_21347,N_20623,N_20841);
nor U21348 (N_21348,N_20820,N_20707);
nor U21349 (N_21349,N_20548,N_20743);
or U21350 (N_21350,N_20909,N_20975);
xnor U21351 (N_21351,N_20920,N_20576);
nor U21352 (N_21352,N_20508,N_20529);
and U21353 (N_21353,N_20773,N_20968);
and U21354 (N_21354,N_20552,N_20896);
or U21355 (N_21355,N_20824,N_20630);
and U21356 (N_21356,N_20672,N_20674);
or U21357 (N_21357,N_20534,N_20594);
xor U21358 (N_21358,N_20540,N_20736);
xor U21359 (N_21359,N_20604,N_20946);
nand U21360 (N_21360,N_20529,N_20984);
xor U21361 (N_21361,N_20710,N_20707);
nand U21362 (N_21362,N_20615,N_20590);
xnor U21363 (N_21363,N_20883,N_20649);
and U21364 (N_21364,N_20903,N_20665);
xnor U21365 (N_21365,N_20562,N_20802);
nor U21366 (N_21366,N_20662,N_20950);
and U21367 (N_21367,N_20754,N_20656);
and U21368 (N_21368,N_20820,N_20811);
and U21369 (N_21369,N_20691,N_20631);
or U21370 (N_21370,N_20870,N_20852);
xor U21371 (N_21371,N_20862,N_20750);
nand U21372 (N_21372,N_20802,N_20933);
nor U21373 (N_21373,N_20965,N_20772);
or U21374 (N_21374,N_20993,N_20601);
xor U21375 (N_21375,N_20916,N_20879);
nor U21376 (N_21376,N_20795,N_20697);
and U21377 (N_21377,N_20632,N_20786);
nor U21378 (N_21378,N_20566,N_20733);
nand U21379 (N_21379,N_20910,N_20883);
nor U21380 (N_21380,N_20809,N_20987);
xnor U21381 (N_21381,N_20843,N_20991);
xnor U21382 (N_21382,N_20937,N_20676);
xor U21383 (N_21383,N_20669,N_20778);
nor U21384 (N_21384,N_20528,N_20981);
or U21385 (N_21385,N_20532,N_20767);
nor U21386 (N_21386,N_20886,N_20750);
xor U21387 (N_21387,N_20699,N_20843);
or U21388 (N_21388,N_20648,N_20774);
or U21389 (N_21389,N_20998,N_20979);
nand U21390 (N_21390,N_20924,N_20675);
nand U21391 (N_21391,N_20532,N_20734);
nand U21392 (N_21392,N_20757,N_20645);
xnor U21393 (N_21393,N_20700,N_20879);
nor U21394 (N_21394,N_20927,N_20626);
xnor U21395 (N_21395,N_20786,N_20587);
nand U21396 (N_21396,N_20953,N_20982);
and U21397 (N_21397,N_20677,N_20816);
nand U21398 (N_21398,N_20809,N_20696);
or U21399 (N_21399,N_20578,N_20821);
or U21400 (N_21400,N_20985,N_20883);
xnor U21401 (N_21401,N_20739,N_20650);
nor U21402 (N_21402,N_20850,N_20774);
or U21403 (N_21403,N_20930,N_20783);
and U21404 (N_21404,N_20957,N_20515);
and U21405 (N_21405,N_20979,N_20788);
nand U21406 (N_21406,N_20836,N_20842);
or U21407 (N_21407,N_20838,N_20762);
or U21408 (N_21408,N_20753,N_20804);
and U21409 (N_21409,N_20807,N_20741);
nand U21410 (N_21410,N_20687,N_20789);
and U21411 (N_21411,N_20853,N_20993);
and U21412 (N_21412,N_20681,N_20673);
nand U21413 (N_21413,N_20630,N_20898);
and U21414 (N_21414,N_20584,N_20598);
nor U21415 (N_21415,N_20828,N_20839);
nand U21416 (N_21416,N_20725,N_20987);
nand U21417 (N_21417,N_20863,N_20728);
or U21418 (N_21418,N_20664,N_20723);
and U21419 (N_21419,N_20559,N_20865);
or U21420 (N_21420,N_20991,N_20768);
nand U21421 (N_21421,N_20952,N_20603);
or U21422 (N_21422,N_20903,N_20781);
nand U21423 (N_21423,N_20954,N_20728);
nor U21424 (N_21424,N_20560,N_20541);
nor U21425 (N_21425,N_20735,N_20746);
nor U21426 (N_21426,N_20709,N_20659);
xor U21427 (N_21427,N_20810,N_20587);
and U21428 (N_21428,N_20927,N_20694);
nand U21429 (N_21429,N_20624,N_20609);
nor U21430 (N_21430,N_20569,N_20834);
or U21431 (N_21431,N_20771,N_20984);
xnor U21432 (N_21432,N_20780,N_20662);
xnor U21433 (N_21433,N_20961,N_20948);
xnor U21434 (N_21434,N_20843,N_20503);
xnor U21435 (N_21435,N_20788,N_20609);
and U21436 (N_21436,N_20895,N_20976);
nand U21437 (N_21437,N_20735,N_20916);
xnor U21438 (N_21438,N_20733,N_20993);
nor U21439 (N_21439,N_20788,N_20678);
or U21440 (N_21440,N_20758,N_20926);
xnor U21441 (N_21441,N_20622,N_20862);
nor U21442 (N_21442,N_20640,N_20848);
and U21443 (N_21443,N_20637,N_20544);
and U21444 (N_21444,N_20740,N_20672);
nand U21445 (N_21445,N_20755,N_20964);
nand U21446 (N_21446,N_20656,N_20958);
nand U21447 (N_21447,N_20799,N_20958);
or U21448 (N_21448,N_20580,N_20713);
nand U21449 (N_21449,N_20800,N_20860);
xnor U21450 (N_21450,N_20570,N_20676);
and U21451 (N_21451,N_20665,N_20901);
or U21452 (N_21452,N_20889,N_20788);
xnor U21453 (N_21453,N_20560,N_20856);
nor U21454 (N_21454,N_20910,N_20610);
nand U21455 (N_21455,N_20758,N_20946);
xor U21456 (N_21456,N_20540,N_20944);
or U21457 (N_21457,N_20924,N_20542);
nor U21458 (N_21458,N_20500,N_20630);
nor U21459 (N_21459,N_20970,N_20765);
nor U21460 (N_21460,N_20966,N_20997);
and U21461 (N_21461,N_20926,N_20749);
and U21462 (N_21462,N_20906,N_20573);
and U21463 (N_21463,N_20537,N_20761);
or U21464 (N_21464,N_20596,N_20508);
nor U21465 (N_21465,N_20608,N_20815);
xor U21466 (N_21466,N_20963,N_20718);
nand U21467 (N_21467,N_20943,N_20839);
xnor U21468 (N_21468,N_20944,N_20579);
nand U21469 (N_21469,N_20694,N_20992);
or U21470 (N_21470,N_20927,N_20780);
and U21471 (N_21471,N_20999,N_20623);
nand U21472 (N_21472,N_20814,N_20836);
or U21473 (N_21473,N_20824,N_20537);
nand U21474 (N_21474,N_20672,N_20715);
and U21475 (N_21475,N_20829,N_20517);
xor U21476 (N_21476,N_20592,N_20624);
nor U21477 (N_21477,N_20544,N_20721);
and U21478 (N_21478,N_20671,N_20638);
xnor U21479 (N_21479,N_20571,N_20730);
nand U21480 (N_21480,N_20607,N_20904);
and U21481 (N_21481,N_20830,N_20819);
or U21482 (N_21482,N_20868,N_20581);
xnor U21483 (N_21483,N_20610,N_20607);
nor U21484 (N_21484,N_20518,N_20956);
or U21485 (N_21485,N_20712,N_20749);
xor U21486 (N_21486,N_20631,N_20561);
nor U21487 (N_21487,N_20620,N_20535);
or U21488 (N_21488,N_20952,N_20766);
or U21489 (N_21489,N_20723,N_20831);
xnor U21490 (N_21490,N_20616,N_20610);
or U21491 (N_21491,N_20588,N_20735);
or U21492 (N_21492,N_20754,N_20584);
nor U21493 (N_21493,N_20605,N_20885);
nand U21494 (N_21494,N_20504,N_20738);
and U21495 (N_21495,N_20837,N_20872);
xor U21496 (N_21496,N_20964,N_20586);
nand U21497 (N_21497,N_20972,N_20790);
or U21498 (N_21498,N_20887,N_20934);
nand U21499 (N_21499,N_20796,N_20816);
xor U21500 (N_21500,N_21338,N_21107);
and U21501 (N_21501,N_21317,N_21253);
xor U21502 (N_21502,N_21115,N_21116);
or U21503 (N_21503,N_21148,N_21449);
nand U21504 (N_21504,N_21096,N_21040);
and U21505 (N_21505,N_21427,N_21225);
and U21506 (N_21506,N_21254,N_21266);
xnor U21507 (N_21507,N_21187,N_21043);
nor U21508 (N_21508,N_21357,N_21000);
nand U21509 (N_21509,N_21349,N_21101);
or U21510 (N_21510,N_21197,N_21273);
nor U21511 (N_21511,N_21214,N_21471);
and U21512 (N_21512,N_21161,N_21049);
and U21513 (N_21513,N_21026,N_21469);
nand U21514 (N_21514,N_21193,N_21324);
nor U21515 (N_21515,N_21461,N_21231);
or U21516 (N_21516,N_21439,N_21311);
nand U21517 (N_21517,N_21344,N_21270);
or U21518 (N_21518,N_21218,N_21323);
or U21519 (N_21519,N_21068,N_21285);
xor U21520 (N_21520,N_21013,N_21297);
nand U21521 (N_21521,N_21367,N_21292);
xor U21522 (N_21522,N_21054,N_21089);
and U21523 (N_21523,N_21224,N_21412);
and U21524 (N_21524,N_21408,N_21024);
or U21525 (N_21525,N_21183,N_21376);
nand U21526 (N_21526,N_21372,N_21246);
and U21527 (N_21527,N_21097,N_21150);
and U21528 (N_21528,N_21245,N_21361);
and U21529 (N_21529,N_21064,N_21299);
or U21530 (N_21530,N_21258,N_21459);
or U21531 (N_21531,N_21241,N_21496);
or U21532 (N_21532,N_21446,N_21379);
nand U21533 (N_21533,N_21256,N_21399);
or U21534 (N_21534,N_21313,N_21030);
or U21535 (N_21535,N_21125,N_21133);
or U21536 (N_21536,N_21084,N_21380);
nand U21537 (N_21537,N_21059,N_21221);
and U21538 (N_21538,N_21127,N_21473);
nand U21539 (N_21539,N_21450,N_21422);
nor U21540 (N_21540,N_21041,N_21001);
nand U21541 (N_21541,N_21111,N_21342);
xnor U21542 (N_21542,N_21331,N_21397);
xnor U21543 (N_21543,N_21110,N_21077);
xor U21544 (N_21544,N_21400,N_21444);
and U21545 (N_21545,N_21011,N_21199);
nand U21546 (N_21546,N_21472,N_21136);
or U21547 (N_21547,N_21207,N_21491);
xor U21548 (N_21548,N_21384,N_21147);
or U21549 (N_21549,N_21365,N_21120);
xnor U21550 (N_21550,N_21490,N_21060);
and U21551 (N_21551,N_21424,N_21360);
or U21552 (N_21552,N_21442,N_21179);
nor U21553 (N_21553,N_21015,N_21204);
nand U21554 (N_21554,N_21401,N_21158);
and U21555 (N_21555,N_21188,N_21033);
and U21556 (N_21556,N_21137,N_21353);
nor U21557 (N_21557,N_21304,N_21470);
nor U21558 (N_21558,N_21182,N_21028);
nor U21559 (N_21559,N_21435,N_21250);
or U21560 (N_21560,N_21319,N_21257);
or U21561 (N_21561,N_21070,N_21190);
nor U21562 (N_21562,N_21144,N_21093);
nor U21563 (N_21563,N_21140,N_21209);
and U21564 (N_21564,N_21240,N_21483);
xor U21565 (N_21565,N_21226,N_21301);
nor U21566 (N_21566,N_21099,N_21385);
xnor U21567 (N_21567,N_21466,N_21062);
nand U21568 (N_21568,N_21235,N_21355);
xor U21569 (N_21569,N_21335,N_21264);
and U21570 (N_21570,N_21429,N_21244);
nand U21571 (N_21571,N_21251,N_21481);
or U21572 (N_21572,N_21411,N_21282);
nor U21573 (N_21573,N_21016,N_21298);
and U21574 (N_21574,N_21328,N_21498);
nor U21575 (N_21575,N_21407,N_21104);
xor U21576 (N_21576,N_21008,N_21362);
nor U21577 (N_21577,N_21057,N_21234);
or U21578 (N_21578,N_21039,N_21050);
and U21579 (N_21579,N_21325,N_21051);
or U21580 (N_21580,N_21172,N_21153);
nand U21581 (N_21581,N_21102,N_21237);
nor U21582 (N_21582,N_21392,N_21262);
and U21583 (N_21583,N_21388,N_21306);
nand U21584 (N_21584,N_21090,N_21086);
and U21585 (N_21585,N_21129,N_21118);
xnor U21586 (N_21586,N_21404,N_21072);
xor U21587 (N_21587,N_21109,N_21479);
nor U21588 (N_21588,N_21315,N_21027);
xor U21589 (N_21589,N_21437,N_21322);
or U21590 (N_21590,N_21268,N_21484);
nand U21591 (N_21591,N_21433,N_21042);
nand U21592 (N_21592,N_21351,N_21291);
and U21593 (N_21593,N_21417,N_21163);
xnor U21594 (N_21594,N_21112,N_21123);
xnor U21595 (N_21595,N_21100,N_21196);
and U21596 (N_21596,N_21073,N_21205);
nor U21597 (N_21597,N_21094,N_21443);
nor U21598 (N_21598,N_21395,N_21434);
or U21599 (N_21599,N_21006,N_21326);
and U21600 (N_21600,N_21467,N_21159);
nor U21601 (N_21601,N_21398,N_21267);
xnor U21602 (N_21602,N_21162,N_21296);
and U21603 (N_21603,N_21402,N_21465);
nand U21604 (N_21604,N_21122,N_21287);
xnor U21605 (N_21605,N_21451,N_21284);
or U21606 (N_21606,N_21430,N_21076);
and U21607 (N_21607,N_21255,N_21352);
and U21608 (N_21608,N_21113,N_21242);
or U21609 (N_21609,N_21020,N_21208);
or U21610 (N_21610,N_21095,N_21048);
and U21611 (N_21611,N_21075,N_21438);
and U21612 (N_21612,N_21281,N_21277);
xor U21613 (N_21613,N_21171,N_21189);
and U21614 (N_21614,N_21203,N_21363);
and U21615 (N_21615,N_21098,N_21421);
nand U21616 (N_21616,N_21170,N_21428);
nand U21617 (N_21617,N_21103,N_21494);
or U21618 (N_21618,N_21227,N_21348);
xor U21619 (N_21619,N_21202,N_21175);
or U21620 (N_21620,N_21327,N_21493);
xor U21621 (N_21621,N_21217,N_21124);
xor U21622 (N_21622,N_21164,N_21128);
xnor U21623 (N_21623,N_21414,N_21154);
nand U21624 (N_21624,N_21452,N_21002);
nand U21625 (N_21625,N_21061,N_21091);
and U21626 (N_21626,N_21354,N_21261);
and U21627 (N_21627,N_21047,N_21044);
nand U21628 (N_21628,N_21377,N_21106);
or U21629 (N_21629,N_21152,N_21223);
or U21630 (N_21630,N_21393,N_21337);
xor U21631 (N_21631,N_21478,N_21195);
or U21632 (N_21632,N_21213,N_21166);
nand U21633 (N_21633,N_21046,N_21426);
and U21634 (N_21634,N_21482,N_21343);
nor U21635 (N_21635,N_21206,N_21371);
xnor U21636 (N_21636,N_21456,N_21014);
and U21637 (N_21637,N_21463,N_21280);
nand U21638 (N_21638,N_21278,N_21228);
nor U21639 (N_21639,N_21283,N_21383);
and U21640 (N_21640,N_21276,N_21074);
xor U21641 (N_21641,N_21167,N_21249);
nand U21642 (N_21642,N_21032,N_21143);
nand U21643 (N_21643,N_21269,N_21263);
xor U21644 (N_21644,N_21010,N_21366);
or U21645 (N_21645,N_21378,N_21055);
nand U21646 (N_21646,N_21037,N_21198);
and U21647 (N_21647,N_21274,N_21488);
or U21648 (N_21648,N_21271,N_21364);
xor U21649 (N_21649,N_21087,N_21121);
nor U21650 (N_21650,N_21448,N_21031);
or U21651 (N_21651,N_21294,N_21447);
and U21652 (N_21652,N_21295,N_21440);
nor U21653 (N_21653,N_21425,N_21080);
or U21654 (N_21654,N_21194,N_21441);
nand U21655 (N_21655,N_21165,N_21088);
nand U21656 (N_21656,N_21489,N_21069);
or U21657 (N_21657,N_21025,N_21035);
and U21658 (N_21658,N_21219,N_21374);
and U21659 (N_21659,N_21334,N_21081);
or U21660 (N_21660,N_21012,N_21078);
nand U21661 (N_21661,N_21370,N_21248);
and U21662 (N_21662,N_21457,N_21359);
xor U21663 (N_21663,N_21117,N_21339);
xor U21664 (N_21664,N_21114,N_21038);
or U21665 (N_21665,N_21460,N_21174);
or U21666 (N_21666,N_21105,N_21135);
or U21667 (N_21667,N_21168,N_21177);
nor U21668 (N_21668,N_21476,N_21492);
nor U21669 (N_21669,N_21141,N_21132);
and U21670 (N_21670,N_21021,N_21350);
nor U21671 (N_21671,N_21329,N_21119);
xor U21672 (N_21672,N_21022,N_21369);
nor U21673 (N_21673,N_21394,N_21139);
nand U21674 (N_21674,N_21239,N_21464);
and U21675 (N_21675,N_21368,N_21056);
xnor U21676 (N_21676,N_21176,N_21346);
or U21677 (N_21677,N_21238,N_21149);
or U21678 (N_21678,N_21432,N_21308);
nor U21679 (N_21679,N_21215,N_21382);
nand U21680 (N_21680,N_21211,N_21279);
nor U21681 (N_21681,N_21300,N_21316);
or U21682 (N_21682,N_21336,N_21222);
xor U21683 (N_21683,N_21455,N_21318);
or U21684 (N_21684,N_21232,N_21418);
or U21685 (N_21685,N_21083,N_21007);
nand U21686 (N_21686,N_21052,N_21431);
or U21687 (N_21687,N_21063,N_21458);
or U21688 (N_21688,N_21333,N_21216);
nor U21689 (N_21689,N_21330,N_21307);
xnor U21690 (N_21690,N_21480,N_21071);
and U21691 (N_21691,N_21423,N_21477);
or U21692 (N_21692,N_21468,N_21356);
and U21693 (N_21693,N_21390,N_21293);
and U21694 (N_21694,N_21169,N_21082);
xor U21695 (N_21695,N_21260,N_21058);
or U21696 (N_21696,N_21286,N_21288);
nor U21697 (N_21697,N_21066,N_21358);
or U21698 (N_21698,N_21184,N_21445);
and U21699 (N_21699,N_21375,N_21151);
or U21700 (N_21700,N_21005,N_21029);
nand U21701 (N_21701,N_21185,N_21065);
nand U21702 (N_21702,N_21036,N_21067);
nor U21703 (N_21703,N_21178,N_21192);
nor U21704 (N_21704,N_21034,N_21310);
nand U21705 (N_21705,N_21079,N_21134);
nand U21706 (N_21706,N_21309,N_21145);
xnor U21707 (N_21707,N_21314,N_21138);
or U21708 (N_21708,N_21220,N_21289);
nand U21709 (N_21709,N_21181,N_21045);
nor U21710 (N_21710,N_21160,N_21415);
nand U21711 (N_21711,N_21436,N_21212);
or U21712 (N_21712,N_21389,N_21462);
nand U21713 (N_21713,N_21230,N_21092);
or U21714 (N_21714,N_21236,N_21191);
nand U21715 (N_21715,N_21180,N_21108);
or U21716 (N_21716,N_21131,N_21453);
or U21717 (N_21717,N_21416,N_21396);
nand U21718 (N_21718,N_21053,N_21386);
xor U21719 (N_21719,N_21004,N_21275);
or U21720 (N_21720,N_21243,N_21173);
and U21721 (N_21721,N_21341,N_21247);
nand U21722 (N_21722,N_21146,N_21387);
and U21723 (N_21723,N_21321,N_21320);
or U21724 (N_21724,N_21487,N_21003);
xnor U21725 (N_21725,N_21312,N_21486);
nor U21726 (N_21726,N_21233,N_21157);
nand U21727 (N_21727,N_21085,N_21485);
nor U21728 (N_21728,N_21410,N_21475);
nand U21729 (N_21729,N_21403,N_21405);
xnor U21730 (N_21730,N_21017,N_21406);
xnor U21731 (N_21731,N_21413,N_21419);
and U21732 (N_21732,N_21126,N_21272);
and U21733 (N_21733,N_21229,N_21019);
and U21734 (N_21734,N_21023,N_21259);
xor U21735 (N_21735,N_21474,N_21142);
nand U21736 (N_21736,N_21252,N_21155);
xor U21737 (N_21737,N_21290,N_21373);
nor U21738 (N_21738,N_21391,N_21200);
or U21739 (N_21739,N_21332,N_21340);
nor U21740 (N_21740,N_21499,N_21201);
nor U21741 (N_21741,N_21302,N_21009);
and U21742 (N_21742,N_21497,N_21381);
xor U21743 (N_21743,N_21345,N_21409);
nand U21744 (N_21744,N_21420,N_21495);
nand U21745 (N_21745,N_21265,N_21018);
nand U21746 (N_21746,N_21156,N_21130);
nor U21747 (N_21747,N_21303,N_21454);
nand U21748 (N_21748,N_21305,N_21186);
nor U21749 (N_21749,N_21347,N_21210);
xnor U21750 (N_21750,N_21216,N_21236);
xor U21751 (N_21751,N_21144,N_21046);
or U21752 (N_21752,N_21052,N_21112);
xor U21753 (N_21753,N_21043,N_21127);
xor U21754 (N_21754,N_21212,N_21131);
xnor U21755 (N_21755,N_21283,N_21408);
xnor U21756 (N_21756,N_21009,N_21132);
or U21757 (N_21757,N_21147,N_21495);
nand U21758 (N_21758,N_21183,N_21047);
or U21759 (N_21759,N_21017,N_21225);
and U21760 (N_21760,N_21336,N_21083);
nand U21761 (N_21761,N_21380,N_21457);
and U21762 (N_21762,N_21270,N_21405);
nor U21763 (N_21763,N_21266,N_21272);
xor U21764 (N_21764,N_21048,N_21213);
nor U21765 (N_21765,N_21082,N_21464);
and U21766 (N_21766,N_21415,N_21044);
nor U21767 (N_21767,N_21087,N_21071);
xnor U21768 (N_21768,N_21092,N_21304);
or U21769 (N_21769,N_21341,N_21198);
xnor U21770 (N_21770,N_21161,N_21284);
nor U21771 (N_21771,N_21480,N_21155);
xnor U21772 (N_21772,N_21469,N_21441);
and U21773 (N_21773,N_21307,N_21426);
and U21774 (N_21774,N_21488,N_21370);
nor U21775 (N_21775,N_21484,N_21014);
and U21776 (N_21776,N_21104,N_21470);
or U21777 (N_21777,N_21370,N_21123);
or U21778 (N_21778,N_21441,N_21000);
or U21779 (N_21779,N_21206,N_21104);
xnor U21780 (N_21780,N_21295,N_21152);
or U21781 (N_21781,N_21348,N_21017);
nor U21782 (N_21782,N_21286,N_21112);
nand U21783 (N_21783,N_21130,N_21067);
nand U21784 (N_21784,N_21344,N_21313);
and U21785 (N_21785,N_21434,N_21176);
or U21786 (N_21786,N_21074,N_21183);
or U21787 (N_21787,N_21375,N_21207);
and U21788 (N_21788,N_21176,N_21100);
and U21789 (N_21789,N_21398,N_21130);
or U21790 (N_21790,N_21347,N_21277);
nand U21791 (N_21791,N_21399,N_21387);
xnor U21792 (N_21792,N_21256,N_21231);
and U21793 (N_21793,N_21026,N_21370);
nor U21794 (N_21794,N_21289,N_21394);
xnor U21795 (N_21795,N_21280,N_21216);
or U21796 (N_21796,N_21418,N_21024);
nand U21797 (N_21797,N_21072,N_21158);
nor U21798 (N_21798,N_21311,N_21222);
nand U21799 (N_21799,N_21029,N_21341);
nor U21800 (N_21800,N_21243,N_21190);
xor U21801 (N_21801,N_21448,N_21237);
or U21802 (N_21802,N_21281,N_21165);
or U21803 (N_21803,N_21264,N_21373);
nor U21804 (N_21804,N_21318,N_21089);
or U21805 (N_21805,N_21329,N_21147);
and U21806 (N_21806,N_21368,N_21198);
nand U21807 (N_21807,N_21136,N_21438);
or U21808 (N_21808,N_21269,N_21375);
and U21809 (N_21809,N_21053,N_21381);
and U21810 (N_21810,N_21207,N_21373);
xnor U21811 (N_21811,N_21166,N_21359);
xnor U21812 (N_21812,N_21070,N_21178);
and U21813 (N_21813,N_21021,N_21105);
and U21814 (N_21814,N_21472,N_21105);
or U21815 (N_21815,N_21384,N_21367);
nand U21816 (N_21816,N_21060,N_21233);
xor U21817 (N_21817,N_21319,N_21150);
nor U21818 (N_21818,N_21243,N_21196);
nor U21819 (N_21819,N_21077,N_21390);
or U21820 (N_21820,N_21364,N_21092);
nor U21821 (N_21821,N_21445,N_21124);
nor U21822 (N_21822,N_21286,N_21317);
and U21823 (N_21823,N_21415,N_21266);
nor U21824 (N_21824,N_21447,N_21217);
and U21825 (N_21825,N_21333,N_21411);
nand U21826 (N_21826,N_21427,N_21155);
nand U21827 (N_21827,N_21091,N_21195);
or U21828 (N_21828,N_21432,N_21137);
nand U21829 (N_21829,N_21393,N_21289);
and U21830 (N_21830,N_21256,N_21274);
nand U21831 (N_21831,N_21324,N_21115);
xor U21832 (N_21832,N_21311,N_21156);
xor U21833 (N_21833,N_21107,N_21397);
or U21834 (N_21834,N_21394,N_21380);
nor U21835 (N_21835,N_21251,N_21241);
xor U21836 (N_21836,N_21348,N_21073);
and U21837 (N_21837,N_21189,N_21311);
nand U21838 (N_21838,N_21293,N_21380);
nand U21839 (N_21839,N_21118,N_21157);
or U21840 (N_21840,N_21219,N_21284);
nor U21841 (N_21841,N_21094,N_21419);
and U21842 (N_21842,N_21215,N_21243);
nor U21843 (N_21843,N_21334,N_21379);
or U21844 (N_21844,N_21394,N_21143);
or U21845 (N_21845,N_21255,N_21302);
and U21846 (N_21846,N_21185,N_21276);
nor U21847 (N_21847,N_21173,N_21264);
or U21848 (N_21848,N_21404,N_21281);
or U21849 (N_21849,N_21349,N_21110);
xor U21850 (N_21850,N_21307,N_21129);
nor U21851 (N_21851,N_21444,N_21333);
xor U21852 (N_21852,N_21180,N_21416);
nand U21853 (N_21853,N_21486,N_21135);
nor U21854 (N_21854,N_21265,N_21427);
nor U21855 (N_21855,N_21132,N_21392);
nor U21856 (N_21856,N_21414,N_21136);
or U21857 (N_21857,N_21289,N_21097);
nand U21858 (N_21858,N_21103,N_21472);
nand U21859 (N_21859,N_21304,N_21452);
nand U21860 (N_21860,N_21018,N_21315);
xor U21861 (N_21861,N_21404,N_21090);
and U21862 (N_21862,N_21420,N_21172);
nor U21863 (N_21863,N_21413,N_21085);
and U21864 (N_21864,N_21069,N_21251);
nor U21865 (N_21865,N_21215,N_21011);
xnor U21866 (N_21866,N_21395,N_21279);
nor U21867 (N_21867,N_21247,N_21407);
and U21868 (N_21868,N_21140,N_21498);
nor U21869 (N_21869,N_21326,N_21364);
and U21870 (N_21870,N_21040,N_21216);
xor U21871 (N_21871,N_21432,N_21387);
nand U21872 (N_21872,N_21385,N_21264);
or U21873 (N_21873,N_21237,N_21003);
nand U21874 (N_21874,N_21316,N_21138);
nand U21875 (N_21875,N_21258,N_21380);
nand U21876 (N_21876,N_21184,N_21440);
xnor U21877 (N_21877,N_21279,N_21212);
xor U21878 (N_21878,N_21431,N_21313);
xnor U21879 (N_21879,N_21441,N_21222);
or U21880 (N_21880,N_21197,N_21179);
nor U21881 (N_21881,N_21098,N_21344);
nor U21882 (N_21882,N_21260,N_21137);
nand U21883 (N_21883,N_21155,N_21050);
or U21884 (N_21884,N_21390,N_21289);
and U21885 (N_21885,N_21163,N_21034);
nand U21886 (N_21886,N_21430,N_21369);
and U21887 (N_21887,N_21477,N_21289);
nor U21888 (N_21888,N_21289,N_21364);
nand U21889 (N_21889,N_21459,N_21158);
nand U21890 (N_21890,N_21349,N_21084);
nand U21891 (N_21891,N_21123,N_21025);
nor U21892 (N_21892,N_21104,N_21055);
and U21893 (N_21893,N_21443,N_21341);
nand U21894 (N_21894,N_21090,N_21257);
or U21895 (N_21895,N_21440,N_21357);
nor U21896 (N_21896,N_21114,N_21166);
xnor U21897 (N_21897,N_21223,N_21326);
nor U21898 (N_21898,N_21320,N_21124);
and U21899 (N_21899,N_21410,N_21290);
or U21900 (N_21900,N_21079,N_21435);
nor U21901 (N_21901,N_21001,N_21148);
nand U21902 (N_21902,N_21252,N_21362);
nand U21903 (N_21903,N_21391,N_21082);
xnor U21904 (N_21904,N_21344,N_21332);
and U21905 (N_21905,N_21418,N_21179);
xnor U21906 (N_21906,N_21367,N_21245);
and U21907 (N_21907,N_21011,N_21499);
and U21908 (N_21908,N_21211,N_21266);
and U21909 (N_21909,N_21399,N_21264);
nand U21910 (N_21910,N_21240,N_21226);
xor U21911 (N_21911,N_21383,N_21265);
and U21912 (N_21912,N_21193,N_21123);
and U21913 (N_21913,N_21022,N_21404);
nand U21914 (N_21914,N_21435,N_21187);
and U21915 (N_21915,N_21254,N_21471);
or U21916 (N_21916,N_21192,N_21484);
xor U21917 (N_21917,N_21410,N_21270);
nand U21918 (N_21918,N_21130,N_21289);
xnor U21919 (N_21919,N_21285,N_21159);
and U21920 (N_21920,N_21164,N_21011);
or U21921 (N_21921,N_21073,N_21448);
nor U21922 (N_21922,N_21275,N_21157);
nand U21923 (N_21923,N_21473,N_21451);
or U21924 (N_21924,N_21058,N_21004);
or U21925 (N_21925,N_21030,N_21011);
or U21926 (N_21926,N_21041,N_21259);
or U21927 (N_21927,N_21446,N_21061);
and U21928 (N_21928,N_21106,N_21269);
xor U21929 (N_21929,N_21161,N_21369);
or U21930 (N_21930,N_21239,N_21386);
and U21931 (N_21931,N_21472,N_21077);
nor U21932 (N_21932,N_21028,N_21203);
and U21933 (N_21933,N_21030,N_21280);
xor U21934 (N_21934,N_21311,N_21098);
and U21935 (N_21935,N_21303,N_21446);
nand U21936 (N_21936,N_21394,N_21295);
and U21937 (N_21937,N_21201,N_21037);
or U21938 (N_21938,N_21119,N_21319);
xnor U21939 (N_21939,N_21102,N_21273);
nand U21940 (N_21940,N_21239,N_21307);
xnor U21941 (N_21941,N_21041,N_21046);
nand U21942 (N_21942,N_21420,N_21381);
nor U21943 (N_21943,N_21393,N_21403);
nor U21944 (N_21944,N_21160,N_21377);
nand U21945 (N_21945,N_21350,N_21236);
nand U21946 (N_21946,N_21112,N_21342);
nor U21947 (N_21947,N_21308,N_21198);
nor U21948 (N_21948,N_21195,N_21387);
or U21949 (N_21949,N_21275,N_21229);
or U21950 (N_21950,N_21486,N_21439);
nand U21951 (N_21951,N_21009,N_21107);
or U21952 (N_21952,N_21105,N_21383);
or U21953 (N_21953,N_21380,N_21302);
xor U21954 (N_21954,N_21370,N_21282);
nor U21955 (N_21955,N_21329,N_21048);
and U21956 (N_21956,N_21125,N_21389);
xor U21957 (N_21957,N_21278,N_21304);
xnor U21958 (N_21958,N_21417,N_21328);
or U21959 (N_21959,N_21203,N_21457);
and U21960 (N_21960,N_21246,N_21139);
nand U21961 (N_21961,N_21305,N_21167);
nor U21962 (N_21962,N_21113,N_21164);
or U21963 (N_21963,N_21033,N_21472);
nand U21964 (N_21964,N_21123,N_21068);
or U21965 (N_21965,N_21404,N_21214);
xor U21966 (N_21966,N_21285,N_21383);
and U21967 (N_21967,N_21495,N_21197);
and U21968 (N_21968,N_21355,N_21109);
nand U21969 (N_21969,N_21006,N_21088);
xor U21970 (N_21970,N_21011,N_21455);
or U21971 (N_21971,N_21236,N_21242);
nand U21972 (N_21972,N_21480,N_21163);
or U21973 (N_21973,N_21434,N_21113);
nor U21974 (N_21974,N_21414,N_21071);
nand U21975 (N_21975,N_21385,N_21298);
xor U21976 (N_21976,N_21280,N_21047);
nand U21977 (N_21977,N_21042,N_21149);
nand U21978 (N_21978,N_21163,N_21232);
nor U21979 (N_21979,N_21073,N_21350);
or U21980 (N_21980,N_21217,N_21087);
and U21981 (N_21981,N_21002,N_21485);
or U21982 (N_21982,N_21015,N_21154);
or U21983 (N_21983,N_21469,N_21154);
xor U21984 (N_21984,N_21423,N_21042);
nor U21985 (N_21985,N_21407,N_21386);
xnor U21986 (N_21986,N_21122,N_21435);
or U21987 (N_21987,N_21056,N_21391);
nor U21988 (N_21988,N_21022,N_21300);
xor U21989 (N_21989,N_21420,N_21491);
nor U21990 (N_21990,N_21172,N_21457);
nand U21991 (N_21991,N_21158,N_21290);
nand U21992 (N_21992,N_21236,N_21363);
and U21993 (N_21993,N_21001,N_21484);
nand U21994 (N_21994,N_21324,N_21054);
nand U21995 (N_21995,N_21091,N_21249);
or U21996 (N_21996,N_21363,N_21436);
nand U21997 (N_21997,N_21243,N_21288);
nor U21998 (N_21998,N_21143,N_21260);
or U21999 (N_21999,N_21163,N_21103);
xnor U22000 (N_22000,N_21926,N_21817);
or U22001 (N_22001,N_21626,N_21580);
and U22002 (N_22002,N_21864,N_21677);
or U22003 (N_22003,N_21916,N_21886);
nand U22004 (N_22004,N_21813,N_21610);
nand U22005 (N_22005,N_21850,N_21814);
or U22006 (N_22006,N_21912,N_21902);
xnor U22007 (N_22007,N_21984,N_21785);
and U22008 (N_22008,N_21568,N_21944);
nor U22009 (N_22009,N_21666,N_21865);
xor U22010 (N_22010,N_21546,N_21513);
and U22011 (N_22011,N_21507,N_21908);
nor U22012 (N_22012,N_21711,N_21592);
nand U22013 (N_22013,N_21995,N_21958);
xor U22014 (N_22014,N_21528,N_21824);
nor U22015 (N_22015,N_21974,N_21803);
xor U22016 (N_22016,N_21981,N_21617);
and U22017 (N_22017,N_21828,N_21838);
and U22018 (N_22018,N_21538,N_21520);
xnor U22019 (N_22019,N_21705,N_21728);
xor U22020 (N_22020,N_21591,N_21941);
or U22021 (N_22021,N_21953,N_21578);
xor U22022 (N_22022,N_21972,N_21544);
xor U22023 (N_22023,N_21554,N_21766);
nand U22024 (N_22024,N_21964,N_21920);
nand U22025 (N_22025,N_21852,N_21631);
xor U22026 (N_22026,N_21843,N_21527);
xnor U22027 (N_22027,N_21980,N_21834);
and U22028 (N_22028,N_21907,N_21888);
nand U22029 (N_22029,N_21909,N_21581);
or U22030 (N_22030,N_21519,N_21690);
nor U22031 (N_22031,N_21783,N_21982);
nor U22032 (N_22032,N_21654,N_21812);
xor U22033 (N_22033,N_21988,N_21603);
or U22034 (N_22034,N_21949,N_21582);
nand U22035 (N_22035,N_21618,N_21717);
nor U22036 (N_22036,N_21773,N_21868);
nand U22037 (N_22037,N_21771,N_21628);
or U22038 (N_22038,N_21742,N_21891);
xor U22039 (N_22039,N_21877,N_21967);
and U22040 (N_22040,N_21727,N_21752);
nor U22041 (N_22041,N_21526,N_21685);
xor U22042 (N_22042,N_21811,N_21575);
or U22043 (N_22043,N_21691,N_21657);
nor U22044 (N_22044,N_21589,N_21833);
and U22045 (N_22045,N_21930,N_21741);
xnor U22046 (N_22046,N_21790,N_21639);
xor U22047 (N_22047,N_21969,N_21718);
nor U22048 (N_22048,N_21855,N_21579);
and U22049 (N_22049,N_21616,N_21897);
nor U22050 (N_22050,N_21956,N_21830);
or U22051 (N_22051,N_21846,N_21750);
xnor U22052 (N_22052,N_21861,N_21583);
and U22053 (N_22053,N_21665,N_21681);
or U22054 (N_22054,N_21904,N_21775);
xnor U22055 (N_22055,N_21608,N_21553);
or U22056 (N_22056,N_21720,N_21703);
and U22057 (N_22057,N_21649,N_21643);
nor U22058 (N_22058,N_21596,N_21551);
nand U22059 (N_22059,N_21895,N_21735);
nor U22060 (N_22060,N_21726,N_21801);
and U22061 (N_22061,N_21802,N_21925);
and U22062 (N_22062,N_21731,N_21598);
xor U22063 (N_22063,N_21706,N_21947);
xnor U22064 (N_22064,N_21531,N_21970);
xnor U22065 (N_22065,N_21655,N_21839);
nand U22066 (N_22066,N_21857,N_21585);
or U22067 (N_22067,N_21670,N_21522);
and U22068 (N_22068,N_21822,N_21879);
xnor U22069 (N_22069,N_21683,N_21662);
nand U22070 (N_22070,N_21695,N_21632);
xor U22071 (N_22071,N_21653,N_21863);
xor U22072 (N_22072,N_21704,N_21832);
and U22073 (N_22073,N_21876,N_21723);
nand U22074 (N_22074,N_21621,N_21883);
or U22075 (N_22075,N_21799,N_21523);
xnor U22076 (N_22076,N_21928,N_21664);
and U22077 (N_22077,N_21829,N_21569);
or U22078 (N_22078,N_21633,N_21744);
nor U22079 (N_22079,N_21772,N_21881);
and U22080 (N_22080,N_21743,N_21647);
nand U22081 (N_22081,N_21699,N_21692);
nor U22082 (N_22082,N_21784,N_21660);
nor U22083 (N_22083,N_21746,N_21989);
nor U22084 (N_22084,N_21763,N_21619);
xor U22085 (N_22085,N_21797,N_21511);
xnor U22086 (N_22086,N_21714,N_21640);
nand U22087 (N_22087,N_21567,N_21851);
and U22088 (N_22088,N_21937,N_21795);
and U22089 (N_22089,N_21805,N_21506);
xnor U22090 (N_22090,N_21867,N_21914);
nand U22091 (N_22091,N_21565,N_21793);
and U22092 (N_22092,N_21900,N_21827);
and U22093 (N_22093,N_21870,N_21976);
xnor U22094 (N_22094,N_21777,N_21906);
nor U22095 (N_22095,N_21586,N_21635);
and U22096 (N_22096,N_21738,N_21588);
and U22097 (N_22097,N_21757,N_21869);
and U22098 (N_22098,N_21796,N_21505);
and U22099 (N_22099,N_21792,N_21535);
nand U22100 (N_22100,N_21678,N_21558);
nor U22101 (N_22101,N_21627,N_21963);
nand U22102 (N_22102,N_21740,N_21878);
nor U22103 (N_22103,N_21543,N_21753);
nor U22104 (N_22104,N_21570,N_21894);
and U22105 (N_22105,N_21954,N_21917);
xnor U22106 (N_22106,N_21629,N_21840);
xor U22107 (N_22107,N_21547,N_21638);
nand U22108 (N_22108,N_21957,N_21856);
nor U22109 (N_22109,N_21573,N_21890);
and U22110 (N_22110,N_21826,N_21605);
xor U22111 (N_22111,N_21787,N_21921);
xnor U22112 (N_22112,N_21593,N_21502);
xnor U22113 (N_22113,N_21701,N_21836);
nor U22114 (N_22114,N_21842,N_21689);
and U22115 (N_22115,N_21550,N_21774);
xnor U22116 (N_22116,N_21676,N_21599);
or U22117 (N_22117,N_21584,N_21533);
nand U22118 (N_22118,N_21809,N_21860);
and U22119 (N_22119,N_21945,N_21871);
nor U22120 (N_22120,N_21806,N_21698);
or U22121 (N_22121,N_21684,N_21913);
nor U22122 (N_22122,N_21854,N_21675);
nand U22123 (N_22123,N_21896,N_21776);
nand U22124 (N_22124,N_21667,N_21786);
nand U22125 (N_22125,N_21931,N_21899);
xnor U22126 (N_22126,N_21755,N_21874);
xor U22127 (N_22127,N_21898,N_21503);
nor U22128 (N_22128,N_21566,N_21724);
and U22129 (N_22129,N_21509,N_21892);
nor U22130 (N_22130,N_21782,N_21905);
xor U22131 (N_22131,N_21821,N_21911);
and U22132 (N_22132,N_21759,N_21745);
and U22133 (N_22133,N_21923,N_21500);
and U22134 (N_22134,N_21819,N_21656);
or U22135 (N_22135,N_21534,N_21977);
xor U22136 (N_22136,N_21985,N_21901);
nor U22137 (N_22137,N_21997,N_21614);
and U22138 (N_22138,N_21688,N_21780);
or U22139 (N_22139,N_21501,N_21548);
nand U22140 (N_22140,N_21996,N_21722);
nor U22141 (N_22141,N_21791,N_21968);
nand U22142 (N_22142,N_21760,N_21927);
nand U22143 (N_22143,N_21915,N_21674);
xor U22144 (N_22144,N_21672,N_21708);
nor U22145 (N_22145,N_21934,N_21630);
nand U22146 (N_22146,N_21889,N_21983);
nor U22147 (N_22147,N_21719,N_21707);
and U22148 (N_22148,N_21936,N_21542);
xor U22149 (N_22149,N_21929,N_21693);
nand U22150 (N_22150,N_21948,N_21768);
xnor U22151 (N_22151,N_21994,N_21918);
or U22152 (N_22152,N_21966,N_21645);
and U22153 (N_22153,N_21823,N_21794);
nand U22154 (N_22154,N_21650,N_21517);
nand U22155 (N_22155,N_21940,N_21648);
xnor U22156 (N_22156,N_21807,N_21748);
and U22157 (N_22157,N_21739,N_21725);
xor U22158 (N_22158,N_21611,N_21564);
nor U22159 (N_22159,N_21761,N_21576);
xor U22160 (N_22160,N_21978,N_21571);
nor U22161 (N_22161,N_21525,N_21991);
nand U22162 (N_22162,N_21789,N_21710);
xnor U22163 (N_22163,N_21998,N_21646);
and U22164 (N_22164,N_21788,N_21975);
and U22165 (N_22165,N_21607,N_21623);
xnor U22166 (N_22166,N_21552,N_21721);
nor U22167 (N_22167,N_21993,N_21514);
or U22168 (N_22168,N_21734,N_21634);
xnor U22169 (N_22169,N_21778,N_21600);
nand U22170 (N_22170,N_21700,N_21938);
nor U22171 (N_22171,N_21999,N_21518);
or U22172 (N_22172,N_21504,N_21668);
nand U22173 (N_22173,N_21922,N_21979);
and U22174 (N_22174,N_21767,N_21873);
or U22175 (N_22175,N_21884,N_21971);
and U22176 (N_22176,N_21804,N_21624);
or U22177 (N_22177,N_21754,N_21820);
nand U22178 (N_22178,N_21713,N_21539);
and U22179 (N_22179,N_21651,N_21955);
and U22180 (N_22180,N_21959,N_21781);
nand U22181 (N_22181,N_21555,N_21559);
nor U22182 (N_22182,N_21549,N_21560);
and U22183 (N_22183,N_21663,N_21682);
nand U22184 (N_22184,N_21730,N_21951);
nand U22185 (N_22185,N_21530,N_21545);
and U22186 (N_22186,N_21694,N_21620);
and U22187 (N_22187,N_21875,N_21841);
and U22188 (N_22188,N_21715,N_21960);
and U22189 (N_22189,N_21800,N_21816);
and U22190 (N_22190,N_21764,N_21636);
nand U22191 (N_22191,N_21686,N_21882);
xor U22192 (N_22192,N_21933,N_21537);
and U22193 (N_22193,N_21987,N_21758);
nor U22194 (N_22194,N_21587,N_21529);
or U22195 (N_22195,N_21737,N_21765);
nor U22196 (N_22196,N_21815,N_21961);
nor U22197 (N_22197,N_21818,N_21601);
nand U22198 (N_22198,N_21973,N_21524);
xor U22199 (N_22199,N_21946,N_21798);
nand U22200 (N_22200,N_21512,N_21613);
or U22201 (N_22201,N_21862,N_21604);
nor U22202 (N_22202,N_21844,N_21680);
and U22203 (N_22203,N_21561,N_21669);
nor U22204 (N_22204,N_21712,N_21590);
nand U22205 (N_22205,N_21943,N_21595);
or U22206 (N_22206,N_21562,N_21556);
or U22207 (N_22207,N_21986,N_21942);
nor U22208 (N_22208,N_21779,N_21848);
or U22209 (N_22209,N_21965,N_21853);
nor U22210 (N_22210,N_21516,N_21935);
and U22211 (N_22211,N_21687,N_21697);
nand U22212 (N_22212,N_21950,N_21924);
xnor U22213 (N_22213,N_21858,N_21887);
nor U22214 (N_22214,N_21609,N_21992);
and U22215 (N_22215,N_21729,N_21732);
nand U22216 (N_22216,N_21859,N_21845);
nand U22217 (N_22217,N_21749,N_21835);
nand U22218 (N_22218,N_21747,N_21849);
nor U22219 (N_22219,N_21637,N_21661);
and U22220 (N_22220,N_21919,N_21837);
xor U22221 (N_22221,N_21885,N_21541);
nand U22222 (N_22222,N_21536,N_21733);
or U22223 (N_22223,N_21532,N_21577);
nor U22224 (N_22224,N_21903,N_21810);
xor U22225 (N_22225,N_21510,N_21910);
and U22226 (N_22226,N_21866,N_21594);
xnor U22227 (N_22227,N_21880,N_21825);
or U22228 (N_22228,N_21831,N_21642);
xnor U22229 (N_22229,N_21612,N_21508);
nor U22230 (N_22230,N_21671,N_21658);
nor U22231 (N_22231,N_21625,N_21872);
or U22232 (N_22232,N_21709,N_21990);
nor U22233 (N_22233,N_21597,N_21808);
and U22234 (N_22234,N_21602,N_21932);
xnor U22235 (N_22235,N_21644,N_21659);
or U22236 (N_22236,N_21736,N_21641);
or U22237 (N_22237,N_21673,N_21847);
and U22238 (N_22238,N_21893,N_21952);
xnor U22239 (N_22239,N_21572,N_21939);
or U22240 (N_22240,N_21679,N_21615);
nand U22241 (N_22241,N_21606,N_21716);
nand U22242 (N_22242,N_21762,N_21769);
and U22243 (N_22243,N_21557,N_21770);
nand U22244 (N_22244,N_21652,N_21751);
and U22245 (N_22245,N_21622,N_21540);
xor U22246 (N_22246,N_21756,N_21515);
nand U22247 (N_22247,N_21563,N_21521);
or U22248 (N_22248,N_21962,N_21696);
nand U22249 (N_22249,N_21702,N_21574);
and U22250 (N_22250,N_21742,N_21621);
nor U22251 (N_22251,N_21831,N_21867);
or U22252 (N_22252,N_21761,N_21832);
xnor U22253 (N_22253,N_21778,N_21591);
or U22254 (N_22254,N_21811,N_21930);
or U22255 (N_22255,N_21733,N_21825);
xnor U22256 (N_22256,N_21655,N_21650);
nand U22257 (N_22257,N_21615,N_21752);
nor U22258 (N_22258,N_21884,N_21968);
nor U22259 (N_22259,N_21699,N_21591);
nor U22260 (N_22260,N_21690,N_21590);
nand U22261 (N_22261,N_21618,N_21567);
and U22262 (N_22262,N_21694,N_21579);
xor U22263 (N_22263,N_21850,N_21946);
nor U22264 (N_22264,N_21736,N_21964);
xor U22265 (N_22265,N_21607,N_21714);
or U22266 (N_22266,N_21516,N_21926);
xor U22267 (N_22267,N_21860,N_21823);
and U22268 (N_22268,N_21711,N_21891);
or U22269 (N_22269,N_21975,N_21759);
xnor U22270 (N_22270,N_21984,N_21650);
xor U22271 (N_22271,N_21549,N_21568);
nor U22272 (N_22272,N_21906,N_21530);
xor U22273 (N_22273,N_21763,N_21960);
or U22274 (N_22274,N_21922,N_21682);
or U22275 (N_22275,N_21833,N_21959);
and U22276 (N_22276,N_21915,N_21970);
or U22277 (N_22277,N_21805,N_21684);
nand U22278 (N_22278,N_21686,N_21552);
nor U22279 (N_22279,N_21935,N_21561);
or U22280 (N_22280,N_21502,N_21519);
xor U22281 (N_22281,N_21724,N_21830);
nor U22282 (N_22282,N_21866,N_21857);
and U22283 (N_22283,N_21537,N_21567);
nor U22284 (N_22284,N_21558,N_21773);
xor U22285 (N_22285,N_21901,N_21813);
and U22286 (N_22286,N_21863,N_21946);
and U22287 (N_22287,N_21893,N_21517);
and U22288 (N_22288,N_21533,N_21793);
xor U22289 (N_22289,N_21703,N_21746);
nand U22290 (N_22290,N_21701,N_21774);
xor U22291 (N_22291,N_21752,N_21888);
and U22292 (N_22292,N_21775,N_21886);
xor U22293 (N_22293,N_21810,N_21547);
xnor U22294 (N_22294,N_21592,N_21602);
xnor U22295 (N_22295,N_21913,N_21765);
nor U22296 (N_22296,N_21849,N_21757);
xor U22297 (N_22297,N_21774,N_21589);
and U22298 (N_22298,N_21620,N_21825);
nor U22299 (N_22299,N_21659,N_21741);
and U22300 (N_22300,N_21699,N_21889);
and U22301 (N_22301,N_21914,N_21509);
xnor U22302 (N_22302,N_21895,N_21780);
nor U22303 (N_22303,N_21749,N_21802);
and U22304 (N_22304,N_21880,N_21903);
nor U22305 (N_22305,N_21767,N_21900);
xor U22306 (N_22306,N_21994,N_21596);
nor U22307 (N_22307,N_21537,N_21942);
xnor U22308 (N_22308,N_21839,N_21789);
nor U22309 (N_22309,N_21547,N_21933);
and U22310 (N_22310,N_21594,N_21774);
xor U22311 (N_22311,N_21535,N_21914);
or U22312 (N_22312,N_21811,N_21882);
xor U22313 (N_22313,N_21890,N_21707);
or U22314 (N_22314,N_21528,N_21635);
nor U22315 (N_22315,N_21958,N_21949);
nor U22316 (N_22316,N_21942,N_21949);
nor U22317 (N_22317,N_21821,N_21577);
and U22318 (N_22318,N_21961,N_21811);
nor U22319 (N_22319,N_21553,N_21807);
and U22320 (N_22320,N_21914,N_21769);
and U22321 (N_22321,N_21573,N_21633);
or U22322 (N_22322,N_21586,N_21850);
xor U22323 (N_22323,N_21828,N_21750);
nand U22324 (N_22324,N_21968,N_21504);
nor U22325 (N_22325,N_21602,N_21525);
nand U22326 (N_22326,N_21763,N_21698);
and U22327 (N_22327,N_21572,N_21511);
or U22328 (N_22328,N_21654,N_21818);
and U22329 (N_22329,N_21800,N_21863);
nand U22330 (N_22330,N_21583,N_21969);
and U22331 (N_22331,N_21722,N_21824);
nand U22332 (N_22332,N_21874,N_21676);
xor U22333 (N_22333,N_21548,N_21734);
or U22334 (N_22334,N_21569,N_21726);
and U22335 (N_22335,N_21737,N_21714);
xor U22336 (N_22336,N_21917,N_21866);
nand U22337 (N_22337,N_21662,N_21963);
or U22338 (N_22338,N_21705,N_21805);
or U22339 (N_22339,N_21597,N_21883);
nand U22340 (N_22340,N_21600,N_21665);
nor U22341 (N_22341,N_21832,N_21792);
xor U22342 (N_22342,N_21828,N_21955);
and U22343 (N_22343,N_21979,N_21563);
xor U22344 (N_22344,N_21889,N_21582);
nor U22345 (N_22345,N_21523,N_21681);
xor U22346 (N_22346,N_21992,N_21790);
nor U22347 (N_22347,N_21705,N_21685);
or U22348 (N_22348,N_21721,N_21720);
xnor U22349 (N_22349,N_21739,N_21581);
and U22350 (N_22350,N_21850,N_21994);
nor U22351 (N_22351,N_21856,N_21552);
nand U22352 (N_22352,N_21816,N_21521);
nand U22353 (N_22353,N_21579,N_21727);
or U22354 (N_22354,N_21684,N_21977);
xor U22355 (N_22355,N_21796,N_21651);
xnor U22356 (N_22356,N_21740,N_21770);
and U22357 (N_22357,N_21977,N_21939);
nand U22358 (N_22358,N_21878,N_21589);
xor U22359 (N_22359,N_21795,N_21737);
nand U22360 (N_22360,N_21763,N_21500);
nor U22361 (N_22361,N_21628,N_21572);
nand U22362 (N_22362,N_21975,N_21633);
nand U22363 (N_22363,N_21730,N_21586);
nand U22364 (N_22364,N_21870,N_21722);
nor U22365 (N_22365,N_21814,N_21692);
xor U22366 (N_22366,N_21817,N_21722);
nor U22367 (N_22367,N_21824,N_21907);
nand U22368 (N_22368,N_21681,N_21624);
xnor U22369 (N_22369,N_21781,N_21988);
xor U22370 (N_22370,N_21901,N_21863);
xor U22371 (N_22371,N_21590,N_21941);
or U22372 (N_22372,N_21952,N_21780);
or U22373 (N_22373,N_21679,N_21916);
nand U22374 (N_22374,N_21797,N_21801);
xnor U22375 (N_22375,N_21563,N_21514);
nor U22376 (N_22376,N_21717,N_21847);
and U22377 (N_22377,N_21535,N_21882);
nor U22378 (N_22378,N_21580,N_21864);
xnor U22379 (N_22379,N_21631,N_21809);
xnor U22380 (N_22380,N_21903,N_21660);
xor U22381 (N_22381,N_21673,N_21775);
xnor U22382 (N_22382,N_21767,N_21985);
xor U22383 (N_22383,N_21733,N_21642);
nand U22384 (N_22384,N_21923,N_21784);
or U22385 (N_22385,N_21804,N_21538);
xor U22386 (N_22386,N_21746,N_21507);
and U22387 (N_22387,N_21568,N_21841);
and U22388 (N_22388,N_21777,N_21991);
and U22389 (N_22389,N_21941,N_21887);
and U22390 (N_22390,N_21892,N_21623);
or U22391 (N_22391,N_21508,N_21940);
nor U22392 (N_22392,N_21653,N_21944);
xnor U22393 (N_22393,N_21709,N_21867);
xor U22394 (N_22394,N_21661,N_21837);
nor U22395 (N_22395,N_21864,N_21644);
nor U22396 (N_22396,N_21854,N_21914);
nand U22397 (N_22397,N_21813,N_21997);
or U22398 (N_22398,N_21510,N_21727);
nor U22399 (N_22399,N_21551,N_21762);
nor U22400 (N_22400,N_21836,N_21938);
nand U22401 (N_22401,N_21983,N_21852);
or U22402 (N_22402,N_21766,N_21514);
nand U22403 (N_22403,N_21819,N_21916);
or U22404 (N_22404,N_21711,N_21714);
and U22405 (N_22405,N_21788,N_21644);
nand U22406 (N_22406,N_21905,N_21813);
nor U22407 (N_22407,N_21545,N_21958);
nor U22408 (N_22408,N_21551,N_21547);
or U22409 (N_22409,N_21939,N_21644);
xnor U22410 (N_22410,N_21934,N_21542);
nor U22411 (N_22411,N_21646,N_21944);
and U22412 (N_22412,N_21838,N_21931);
or U22413 (N_22413,N_21907,N_21926);
nor U22414 (N_22414,N_21534,N_21558);
nand U22415 (N_22415,N_21568,N_21832);
nand U22416 (N_22416,N_21672,N_21633);
and U22417 (N_22417,N_21699,N_21863);
nand U22418 (N_22418,N_21589,N_21634);
xnor U22419 (N_22419,N_21753,N_21769);
and U22420 (N_22420,N_21835,N_21615);
nor U22421 (N_22421,N_21625,N_21829);
or U22422 (N_22422,N_21607,N_21682);
nor U22423 (N_22423,N_21894,N_21883);
or U22424 (N_22424,N_21522,N_21701);
nor U22425 (N_22425,N_21574,N_21844);
and U22426 (N_22426,N_21996,N_21849);
and U22427 (N_22427,N_21894,N_21533);
nand U22428 (N_22428,N_21578,N_21554);
or U22429 (N_22429,N_21550,N_21799);
nor U22430 (N_22430,N_21855,N_21791);
xor U22431 (N_22431,N_21711,N_21915);
nor U22432 (N_22432,N_21762,N_21600);
or U22433 (N_22433,N_21784,N_21901);
or U22434 (N_22434,N_21871,N_21690);
and U22435 (N_22435,N_21812,N_21672);
nand U22436 (N_22436,N_21527,N_21892);
nor U22437 (N_22437,N_21578,N_21847);
nor U22438 (N_22438,N_21525,N_21584);
xnor U22439 (N_22439,N_21899,N_21804);
or U22440 (N_22440,N_21961,N_21638);
or U22441 (N_22441,N_21776,N_21569);
xor U22442 (N_22442,N_21811,N_21589);
xor U22443 (N_22443,N_21757,N_21903);
and U22444 (N_22444,N_21924,N_21974);
nand U22445 (N_22445,N_21734,N_21912);
nand U22446 (N_22446,N_21874,N_21888);
or U22447 (N_22447,N_21556,N_21573);
nor U22448 (N_22448,N_21605,N_21626);
nor U22449 (N_22449,N_21552,N_21674);
nor U22450 (N_22450,N_21561,N_21588);
xor U22451 (N_22451,N_21552,N_21970);
nand U22452 (N_22452,N_21687,N_21926);
xor U22453 (N_22453,N_21596,N_21928);
or U22454 (N_22454,N_21665,N_21624);
or U22455 (N_22455,N_21735,N_21966);
and U22456 (N_22456,N_21531,N_21590);
xnor U22457 (N_22457,N_21721,N_21620);
or U22458 (N_22458,N_21951,N_21846);
and U22459 (N_22459,N_21619,N_21572);
and U22460 (N_22460,N_21974,N_21513);
or U22461 (N_22461,N_21866,N_21610);
or U22462 (N_22462,N_21501,N_21640);
or U22463 (N_22463,N_21578,N_21506);
xor U22464 (N_22464,N_21993,N_21941);
or U22465 (N_22465,N_21884,N_21505);
nand U22466 (N_22466,N_21715,N_21968);
or U22467 (N_22467,N_21825,N_21994);
nand U22468 (N_22468,N_21796,N_21589);
or U22469 (N_22469,N_21672,N_21651);
xnor U22470 (N_22470,N_21964,N_21746);
nor U22471 (N_22471,N_21607,N_21689);
nor U22472 (N_22472,N_21541,N_21946);
nand U22473 (N_22473,N_21839,N_21765);
xnor U22474 (N_22474,N_21999,N_21990);
xor U22475 (N_22475,N_21615,N_21928);
nor U22476 (N_22476,N_21736,N_21879);
nand U22477 (N_22477,N_21719,N_21512);
or U22478 (N_22478,N_21715,N_21669);
xnor U22479 (N_22479,N_21869,N_21957);
nor U22480 (N_22480,N_21593,N_21952);
and U22481 (N_22481,N_21774,N_21924);
xor U22482 (N_22482,N_21824,N_21970);
nor U22483 (N_22483,N_21861,N_21515);
or U22484 (N_22484,N_21639,N_21612);
nand U22485 (N_22485,N_21719,N_21623);
and U22486 (N_22486,N_21647,N_21630);
xor U22487 (N_22487,N_21945,N_21539);
or U22488 (N_22488,N_21816,N_21569);
xor U22489 (N_22489,N_21897,N_21751);
nor U22490 (N_22490,N_21892,N_21538);
nand U22491 (N_22491,N_21829,N_21841);
or U22492 (N_22492,N_21669,N_21834);
and U22493 (N_22493,N_21870,N_21712);
and U22494 (N_22494,N_21782,N_21823);
and U22495 (N_22495,N_21598,N_21569);
xor U22496 (N_22496,N_21767,N_21573);
and U22497 (N_22497,N_21665,N_21992);
and U22498 (N_22498,N_21625,N_21847);
xor U22499 (N_22499,N_21901,N_21690);
or U22500 (N_22500,N_22084,N_22124);
or U22501 (N_22501,N_22202,N_22417);
xor U22502 (N_22502,N_22366,N_22476);
nand U22503 (N_22503,N_22160,N_22112);
nand U22504 (N_22504,N_22182,N_22425);
or U22505 (N_22505,N_22135,N_22304);
xnor U22506 (N_22506,N_22376,N_22231);
and U22507 (N_22507,N_22164,N_22411);
and U22508 (N_22508,N_22488,N_22079);
nand U22509 (N_22509,N_22009,N_22424);
or U22510 (N_22510,N_22186,N_22350);
nor U22511 (N_22511,N_22318,N_22441);
or U22512 (N_22512,N_22222,N_22352);
xnor U22513 (N_22513,N_22220,N_22263);
or U22514 (N_22514,N_22052,N_22058);
nand U22515 (N_22515,N_22308,N_22224);
nor U22516 (N_22516,N_22282,N_22130);
and U22517 (N_22517,N_22322,N_22024);
nand U22518 (N_22518,N_22319,N_22167);
nor U22519 (N_22519,N_22148,N_22074);
xor U22520 (N_22520,N_22384,N_22383);
nor U22521 (N_22521,N_22152,N_22485);
xor U22522 (N_22522,N_22387,N_22083);
xnor U22523 (N_22523,N_22109,N_22474);
and U22524 (N_22524,N_22397,N_22420);
nand U22525 (N_22525,N_22405,N_22492);
or U22526 (N_22526,N_22293,N_22195);
and U22527 (N_22527,N_22310,N_22363);
xor U22528 (N_22528,N_22144,N_22131);
and U22529 (N_22529,N_22015,N_22280);
nor U22530 (N_22530,N_22257,N_22359);
nor U22531 (N_22531,N_22415,N_22315);
nand U22532 (N_22532,N_22029,N_22400);
or U22533 (N_22533,N_22106,N_22171);
nand U22534 (N_22534,N_22028,N_22126);
nand U22535 (N_22535,N_22031,N_22380);
nor U22536 (N_22536,N_22334,N_22023);
or U22537 (N_22537,N_22372,N_22409);
nor U22538 (N_22538,N_22462,N_22139);
xor U22539 (N_22539,N_22272,N_22165);
nor U22540 (N_22540,N_22404,N_22001);
nor U22541 (N_22541,N_22197,N_22393);
or U22542 (N_22542,N_22456,N_22064);
and U22543 (N_22543,N_22453,N_22207);
and U22544 (N_22544,N_22180,N_22209);
xnor U22545 (N_22545,N_22091,N_22089);
xor U22546 (N_22546,N_22045,N_22273);
nor U22547 (N_22547,N_22275,N_22175);
xor U22548 (N_22548,N_22078,N_22427);
or U22549 (N_22549,N_22337,N_22090);
or U22550 (N_22550,N_22094,N_22082);
and U22551 (N_22551,N_22295,N_22373);
xor U22552 (N_22552,N_22204,N_22184);
xnor U22553 (N_22553,N_22253,N_22431);
xnor U22554 (N_22554,N_22020,N_22391);
nand U22555 (N_22555,N_22348,N_22287);
nor U22556 (N_22556,N_22369,N_22395);
nor U22557 (N_22557,N_22357,N_22223);
nor U22558 (N_22558,N_22101,N_22098);
and U22559 (N_22559,N_22166,N_22149);
nand U22560 (N_22560,N_22245,N_22459);
nor U22561 (N_22561,N_22193,N_22057);
xnor U22562 (N_22562,N_22191,N_22181);
and U22563 (N_22563,N_22004,N_22185);
or U22564 (N_22564,N_22085,N_22070);
xor U22565 (N_22565,N_22413,N_22136);
or U22566 (N_22566,N_22343,N_22030);
xor U22567 (N_22567,N_22340,N_22241);
or U22568 (N_22568,N_22143,N_22068);
or U22569 (N_22569,N_22303,N_22258);
xnor U22570 (N_22570,N_22483,N_22328);
xor U22571 (N_22571,N_22033,N_22339);
xnor U22572 (N_22572,N_22086,N_22433);
nand U22573 (N_22573,N_22443,N_22429);
nand U22574 (N_22574,N_22019,N_22403);
nand U22575 (N_22575,N_22076,N_22386);
nor U22576 (N_22576,N_22438,N_22205);
nand U22577 (N_22577,N_22290,N_22196);
nor U22578 (N_22578,N_22103,N_22330);
nand U22579 (N_22579,N_22016,N_22137);
nor U22580 (N_22580,N_22497,N_22450);
nor U22581 (N_22581,N_22134,N_22174);
or U22582 (N_22582,N_22219,N_22478);
and U22583 (N_22583,N_22296,N_22027);
nor U22584 (N_22584,N_22236,N_22466);
or U22585 (N_22585,N_22270,N_22495);
or U22586 (N_22586,N_22260,N_22121);
and U22587 (N_22587,N_22323,N_22440);
nor U22588 (N_22588,N_22163,N_22013);
or U22589 (N_22589,N_22277,N_22235);
xor U22590 (N_22590,N_22201,N_22170);
or U22591 (N_22591,N_22423,N_22344);
nand U22592 (N_22592,N_22324,N_22002);
or U22593 (N_22593,N_22189,N_22056);
and U22594 (N_22594,N_22188,N_22269);
or U22595 (N_22595,N_22436,N_22102);
nor U22596 (N_22596,N_22448,N_22421);
and U22597 (N_22597,N_22177,N_22128);
xnor U22598 (N_22598,N_22161,N_22491);
nand U22599 (N_22599,N_22410,N_22454);
and U22600 (N_22600,N_22368,N_22381);
nand U22601 (N_22601,N_22012,N_22317);
nor U22602 (N_22602,N_22370,N_22138);
and U22603 (N_22603,N_22120,N_22242);
nor U22604 (N_22604,N_22355,N_22298);
xnor U22605 (N_22605,N_22375,N_22458);
xor U22606 (N_22606,N_22008,N_22168);
and U22607 (N_22607,N_22218,N_22301);
nor U22608 (N_22608,N_22244,N_22468);
nand U22609 (N_22609,N_22125,N_22479);
or U22610 (N_22610,N_22155,N_22416);
or U22611 (N_22611,N_22435,N_22210);
xnor U22612 (N_22612,N_22158,N_22095);
nor U22613 (N_22613,N_22108,N_22407);
xnor U22614 (N_22614,N_22477,N_22461);
nand U22615 (N_22615,N_22358,N_22087);
xor U22616 (N_22616,N_22104,N_22025);
or U22617 (N_22617,N_22046,N_22036);
and U22618 (N_22618,N_22005,N_22329);
or U22619 (N_22619,N_22014,N_22034);
and U22620 (N_22620,N_22011,N_22499);
nand U22621 (N_22621,N_22316,N_22153);
nor U22622 (N_22622,N_22059,N_22053);
nand U22623 (N_22623,N_22469,N_22447);
xnor U22624 (N_22624,N_22035,N_22299);
nor U22625 (N_22625,N_22238,N_22365);
nor U22626 (N_22626,N_22183,N_22455);
nand U22627 (N_22627,N_22229,N_22412);
nor U22628 (N_22628,N_22278,N_22345);
nand U22629 (N_22629,N_22051,N_22038);
and U22630 (N_22630,N_22162,N_22142);
nor U22631 (N_22631,N_22156,N_22394);
or U22632 (N_22632,N_22347,N_22279);
xnor U22633 (N_22633,N_22115,N_22065);
or U22634 (N_22634,N_22093,N_22389);
and U22635 (N_22635,N_22467,N_22401);
and U22636 (N_22636,N_22026,N_22061);
nor U22637 (N_22637,N_22037,N_22498);
xor U22638 (N_22638,N_22234,N_22221);
or U22639 (N_22639,N_22157,N_22073);
xor U22640 (N_22640,N_22044,N_22276);
nor U22641 (N_22641,N_22226,N_22463);
or U22642 (N_22642,N_22169,N_22040);
xor U22643 (N_22643,N_22364,N_22192);
nor U22644 (N_22644,N_22489,N_22105);
or U22645 (N_22645,N_22398,N_22042);
or U22646 (N_22646,N_22041,N_22388);
nor U22647 (N_22647,N_22261,N_22252);
nand U22648 (N_22648,N_22378,N_22274);
nor U22649 (N_22649,N_22206,N_22419);
nand U22650 (N_22650,N_22396,N_22346);
or U22651 (N_22651,N_22406,N_22333);
nor U22652 (N_22652,N_22217,N_22362);
nand U22653 (N_22653,N_22232,N_22018);
or U22654 (N_22654,N_22190,N_22493);
and U22655 (N_22655,N_22471,N_22060);
xnor U22656 (N_22656,N_22147,N_22306);
nor U22657 (N_22657,N_22043,N_22000);
nor U22658 (N_22658,N_22281,N_22356);
nand U22659 (N_22659,N_22114,N_22486);
or U22660 (N_22660,N_22338,N_22266);
nor U22661 (N_22661,N_22141,N_22017);
xor U22662 (N_22662,N_22311,N_22211);
and U22663 (N_22663,N_22256,N_22048);
nand U22664 (N_22664,N_22063,N_22097);
nor U22665 (N_22665,N_22198,N_22006);
or U22666 (N_22666,N_22426,N_22442);
and U22667 (N_22667,N_22075,N_22484);
or U22668 (N_22668,N_22314,N_22003);
nand U22669 (N_22669,N_22176,N_22255);
and U22670 (N_22670,N_22110,N_22203);
nor U22671 (N_22671,N_22129,N_22250);
nor U22672 (N_22672,N_22451,N_22259);
nor U22673 (N_22673,N_22422,N_22151);
xnor U22674 (N_22674,N_22313,N_22213);
or U22675 (N_22675,N_22123,N_22360);
and U22676 (N_22676,N_22305,N_22268);
nor U22677 (N_22677,N_22122,N_22418);
and U22678 (N_22678,N_22445,N_22371);
or U22679 (N_22679,N_22228,N_22374);
nor U22680 (N_22680,N_22145,N_22237);
or U22681 (N_22681,N_22199,N_22490);
nor U22682 (N_22682,N_22481,N_22119);
nor U22683 (N_22683,N_22464,N_22351);
and U22684 (N_22684,N_22286,N_22353);
or U22685 (N_22685,N_22361,N_22178);
nand U22686 (N_22686,N_22284,N_22179);
nor U22687 (N_22687,N_22039,N_22062);
or U22688 (N_22688,N_22377,N_22473);
or U22689 (N_22689,N_22312,N_22309);
nand U22690 (N_22690,N_22050,N_22265);
nor U22691 (N_22691,N_22264,N_22099);
nand U22692 (N_22692,N_22444,N_22283);
and U22693 (N_22693,N_22172,N_22254);
nor U22694 (N_22694,N_22327,N_22480);
nand U22695 (N_22695,N_22227,N_22225);
and U22696 (N_22696,N_22320,N_22392);
nor U22697 (N_22697,N_22249,N_22132);
and U22698 (N_22698,N_22247,N_22472);
and U22699 (N_22699,N_22146,N_22288);
nor U22700 (N_22700,N_22096,N_22494);
nand U22701 (N_22701,N_22470,N_22187);
or U22702 (N_22702,N_22460,N_22430);
and U22703 (N_22703,N_22292,N_22321);
or U22704 (N_22704,N_22248,N_22331);
xor U22705 (N_22705,N_22437,N_22335);
nor U22706 (N_22706,N_22414,N_22294);
or U22707 (N_22707,N_22496,N_22066);
and U22708 (N_22708,N_22118,N_22173);
and U22709 (N_22709,N_22341,N_22326);
and U22710 (N_22710,N_22246,N_22072);
nor U22711 (N_22711,N_22200,N_22214);
nand U22712 (N_22712,N_22285,N_22081);
or U22713 (N_22713,N_22251,N_22216);
nor U22714 (N_22714,N_22054,N_22067);
nand U22715 (N_22715,N_22159,N_22194);
xnor U22716 (N_22716,N_22239,N_22071);
nand U22717 (N_22717,N_22069,N_22007);
xor U22718 (N_22718,N_22336,N_22342);
xor U22719 (N_22719,N_22077,N_22262);
nand U22720 (N_22720,N_22439,N_22230);
xnor U22721 (N_22721,N_22297,N_22302);
and U22722 (N_22722,N_22116,N_22271);
xnor U22723 (N_22723,N_22332,N_22399);
nor U22724 (N_22724,N_22212,N_22113);
nor U22725 (N_22725,N_22408,N_22289);
nor U22726 (N_22726,N_22117,N_22055);
nand U22727 (N_22727,N_22010,N_22291);
or U22728 (N_22728,N_22154,N_22475);
nand U22729 (N_22729,N_22449,N_22402);
xnor U22730 (N_22730,N_22100,N_22452);
nor U22731 (N_22731,N_22307,N_22107);
and U22732 (N_22732,N_22133,N_22208);
nor U22733 (N_22733,N_22487,N_22127);
or U22734 (N_22734,N_22482,N_22385);
nand U22735 (N_22735,N_22092,N_22446);
or U22736 (N_22736,N_22432,N_22267);
xor U22737 (N_22737,N_22465,N_22367);
or U22738 (N_22738,N_22080,N_22022);
nand U22739 (N_22739,N_22049,N_22150);
or U22740 (N_22740,N_22243,N_22088);
xnor U22741 (N_22741,N_22140,N_22111);
xor U22742 (N_22742,N_22215,N_22047);
or U22743 (N_22743,N_22354,N_22434);
and U22744 (N_22744,N_22032,N_22233);
nand U22745 (N_22745,N_22300,N_22382);
nand U22746 (N_22746,N_22390,N_22428);
nand U22747 (N_22747,N_22349,N_22240);
and U22748 (N_22748,N_22457,N_22325);
nand U22749 (N_22749,N_22021,N_22379);
and U22750 (N_22750,N_22395,N_22009);
and U22751 (N_22751,N_22037,N_22088);
or U22752 (N_22752,N_22351,N_22016);
xor U22753 (N_22753,N_22069,N_22225);
or U22754 (N_22754,N_22324,N_22422);
nor U22755 (N_22755,N_22381,N_22203);
nand U22756 (N_22756,N_22429,N_22174);
or U22757 (N_22757,N_22175,N_22307);
nor U22758 (N_22758,N_22079,N_22331);
nor U22759 (N_22759,N_22108,N_22375);
or U22760 (N_22760,N_22327,N_22216);
and U22761 (N_22761,N_22004,N_22033);
xor U22762 (N_22762,N_22390,N_22446);
nor U22763 (N_22763,N_22341,N_22459);
nand U22764 (N_22764,N_22337,N_22421);
or U22765 (N_22765,N_22383,N_22492);
or U22766 (N_22766,N_22000,N_22067);
nor U22767 (N_22767,N_22094,N_22370);
nand U22768 (N_22768,N_22383,N_22457);
nor U22769 (N_22769,N_22270,N_22211);
nor U22770 (N_22770,N_22013,N_22434);
and U22771 (N_22771,N_22250,N_22033);
or U22772 (N_22772,N_22211,N_22100);
nor U22773 (N_22773,N_22403,N_22008);
or U22774 (N_22774,N_22057,N_22419);
xnor U22775 (N_22775,N_22140,N_22160);
or U22776 (N_22776,N_22277,N_22384);
or U22777 (N_22777,N_22436,N_22190);
xnor U22778 (N_22778,N_22297,N_22330);
xnor U22779 (N_22779,N_22369,N_22078);
nand U22780 (N_22780,N_22092,N_22422);
nor U22781 (N_22781,N_22246,N_22462);
xor U22782 (N_22782,N_22459,N_22286);
nand U22783 (N_22783,N_22276,N_22367);
and U22784 (N_22784,N_22458,N_22283);
nor U22785 (N_22785,N_22331,N_22406);
and U22786 (N_22786,N_22249,N_22317);
nor U22787 (N_22787,N_22317,N_22489);
and U22788 (N_22788,N_22030,N_22373);
and U22789 (N_22789,N_22402,N_22201);
xor U22790 (N_22790,N_22298,N_22378);
and U22791 (N_22791,N_22192,N_22235);
nor U22792 (N_22792,N_22032,N_22243);
xor U22793 (N_22793,N_22030,N_22344);
or U22794 (N_22794,N_22235,N_22248);
nor U22795 (N_22795,N_22183,N_22052);
xor U22796 (N_22796,N_22390,N_22133);
or U22797 (N_22797,N_22195,N_22401);
nand U22798 (N_22798,N_22405,N_22427);
xor U22799 (N_22799,N_22091,N_22376);
and U22800 (N_22800,N_22098,N_22488);
nor U22801 (N_22801,N_22270,N_22057);
nand U22802 (N_22802,N_22448,N_22288);
nor U22803 (N_22803,N_22322,N_22277);
nor U22804 (N_22804,N_22488,N_22082);
or U22805 (N_22805,N_22007,N_22190);
or U22806 (N_22806,N_22211,N_22358);
nand U22807 (N_22807,N_22046,N_22177);
nor U22808 (N_22808,N_22254,N_22038);
nand U22809 (N_22809,N_22450,N_22479);
xnor U22810 (N_22810,N_22013,N_22311);
and U22811 (N_22811,N_22360,N_22076);
nor U22812 (N_22812,N_22413,N_22277);
nand U22813 (N_22813,N_22156,N_22220);
nor U22814 (N_22814,N_22369,N_22430);
xnor U22815 (N_22815,N_22217,N_22147);
or U22816 (N_22816,N_22249,N_22074);
and U22817 (N_22817,N_22201,N_22416);
nor U22818 (N_22818,N_22305,N_22007);
nand U22819 (N_22819,N_22384,N_22060);
nand U22820 (N_22820,N_22100,N_22360);
and U22821 (N_22821,N_22031,N_22268);
nor U22822 (N_22822,N_22140,N_22123);
nand U22823 (N_22823,N_22230,N_22047);
nand U22824 (N_22824,N_22421,N_22237);
nor U22825 (N_22825,N_22258,N_22357);
nand U22826 (N_22826,N_22153,N_22126);
xor U22827 (N_22827,N_22173,N_22075);
xor U22828 (N_22828,N_22345,N_22188);
xnor U22829 (N_22829,N_22316,N_22221);
nand U22830 (N_22830,N_22471,N_22141);
and U22831 (N_22831,N_22348,N_22364);
nand U22832 (N_22832,N_22236,N_22069);
and U22833 (N_22833,N_22318,N_22392);
or U22834 (N_22834,N_22156,N_22463);
nor U22835 (N_22835,N_22223,N_22189);
and U22836 (N_22836,N_22057,N_22228);
or U22837 (N_22837,N_22401,N_22321);
and U22838 (N_22838,N_22058,N_22184);
and U22839 (N_22839,N_22168,N_22243);
or U22840 (N_22840,N_22164,N_22424);
and U22841 (N_22841,N_22192,N_22158);
nand U22842 (N_22842,N_22050,N_22467);
nand U22843 (N_22843,N_22241,N_22332);
nand U22844 (N_22844,N_22154,N_22171);
xnor U22845 (N_22845,N_22353,N_22023);
nand U22846 (N_22846,N_22301,N_22098);
nor U22847 (N_22847,N_22354,N_22045);
xnor U22848 (N_22848,N_22102,N_22101);
or U22849 (N_22849,N_22226,N_22092);
and U22850 (N_22850,N_22126,N_22352);
nor U22851 (N_22851,N_22406,N_22499);
or U22852 (N_22852,N_22172,N_22280);
and U22853 (N_22853,N_22498,N_22305);
nand U22854 (N_22854,N_22056,N_22016);
xnor U22855 (N_22855,N_22144,N_22325);
or U22856 (N_22856,N_22059,N_22184);
xnor U22857 (N_22857,N_22078,N_22269);
xor U22858 (N_22858,N_22142,N_22268);
xnor U22859 (N_22859,N_22364,N_22494);
or U22860 (N_22860,N_22460,N_22199);
and U22861 (N_22861,N_22297,N_22388);
and U22862 (N_22862,N_22043,N_22344);
nand U22863 (N_22863,N_22318,N_22365);
or U22864 (N_22864,N_22339,N_22060);
nor U22865 (N_22865,N_22425,N_22326);
and U22866 (N_22866,N_22368,N_22337);
and U22867 (N_22867,N_22316,N_22238);
or U22868 (N_22868,N_22121,N_22231);
nand U22869 (N_22869,N_22174,N_22474);
nor U22870 (N_22870,N_22409,N_22010);
and U22871 (N_22871,N_22120,N_22060);
nand U22872 (N_22872,N_22390,N_22489);
xor U22873 (N_22873,N_22224,N_22352);
or U22874 (N_22874,N_22112,N_22299);
xnor U22875 (N_22875,N_22493,N_22027);
and U22876 (N_22876,N_22236,N_22134);
nor U22877 (N_22877,N_22447,N_22083);
and U22878 (N_22878,N_22114,N_22171);
and U22879 (N_22879,N_22263,N_22193);
or U22880 (N_22880,N_22086,N_22291);
nor U22881 (N_22881,N_22057,N_22015);
nor U22882 (N_22882,N_22022,N_22335);
xor U22883 (N_22883,N_22008,N_22499);
xor U22884 (N_22884,N_22388,N_22214);
nand U22885 (N_22885,N_22058,N_22144);
or U22886 (N_22886,N_22341,N_22485);
nor U22887 (N_22887,N_22192,N_22191);
nand U22888 (N_22888,N_22438,N_22390);
xnor U22889 (N_22889,N_22229,N_22126);
xnor U22890 (N_22890,N_22206,N_22173);
xor U22891 (N_22891,N_22092,N_22038);
nand U22892 (N_22892,N_22445,N_22125);
nand U22893 (N_22893,N_22026,N_22485);
nor U22894 (N_22894,N_22282,N_22188);
and U22895 (N_22895,N_22476,N_22054);
nand U22896 (N_22896,N_22127,N_22412);
nand U22897 (N_22897,N_22059,N_22121);
or U22898 (N_22898,N_22498,N_22219);
nand U22899 (N_22899,N_22161,N_22065);
and U22900 (N_22900,N_22116,N_22382);
or U22901 (N_22901,N_22143,N_22233);
nor U22902 (N_22902,N_22006,N_22287);
nand U22903 (N_22903,N_22036,N_22221);
nand U22904 (N_22904,N_22376,N_22291);
nand U22905 (N_22905,N_22049,N_22328);
or U22906 (N_22906,N_22381,N_22017);
or U22907 (N_22907,N_22483,N_22058);
xnor U22908 (N_22908,N_22013,N_22068);
xor U22909 (N_22909,N_22165,N_22121);
or U22910 (N_22910,N_22344,N_22128);
or U22911 (N_22911,N_22393,N_22192);
xor U22912 (N_22912,N_22089,N_22044);
nand U22913 (N_22913,N_22221,N_22004);
xor U22914 (N_22914,N_22496,N_22214);
nand U22915 (N_22915,N_22149,N_22376);
and U22916 (N_22916,N_22115,N_22449);
and U22917 (N_22917,N_22385,N_22040);
or U22918 (N_22918,N_22201,N_22394);
xnor U22919 (N_22919,N_22377,N_22498);
nand U22920 (N_22920,N_22482,N_22408);
nand U22921 (N_22921,N_22461,N_22428);
nand U22922 (N_22922,N_22412,N_22346);
nand U22923 (N_22923,N_22076,N_22303);
and U22924 (N_22924,N_22310,N_22216);
xnor U22925 (N_22925,N_22452,N_22476);
nand U22926 (N_22926,N_22324,N_22346);
and U22927 (N_22927,N_22467,N_22436);
nand U22928 (N_22928,N_22437,N_22461);
or U22929 (N_22929,N_22139,N_22195);
nor U22930 (N_22930,N_22016,N_22404);
and U22931 (N_22931,N_22153,N_22331);
nand U22932 (N_22932,N_22173,N_22308);
or U22933 (N_22933,N_22066,N_22259);
or U22934 (N_22934,N_22322,N_22466);
xor U22935 (N_22935,N_22168,N_22055);
nand U22936 (N_22936,N_22085,N_22014);
nor U22937 (N_22937,N_22299,N_22072);
or U22938 (N_22938,N_22447,N_22488);
nor U22939 (N_22939,N_22436,N_22087);
nor U22940 (N_22940,N_22498,N_22308);
and U22941 (N_22941,N_22063,N_22190);
and U22942 (N_22942,N_22019,N_22175);
xnor U22943 (N_22943,N_22455,N_22133);
nand U22944 (N_22944,N_22466,N_22428);
nand U22945 (N_22945,N_22483,N_22197);
or U22946 (N_22946,N_22023,N_22096);
nand U22947 (N_22947,N_22346,N_22129);
nand U22948 (N_22948,N_22213,N_22101);
xnor U22949 (N_22949,N_22379,N_22414);
nand U22950 (N_22950,N_22378,N_22261);
nor U22951 (N_22951,N_22164,N_22431);
and U22952 (N_22952,N_22181,N_22434);
nand U22953 (N_22953,N_22277,N_22159);
xor U22954 (N_22954,N_22404,N_22236);
and U22955 (N_22955,N_22159,N_22383);
nor U22956 (N_22956,N_22433,N_22455);
and U22957 (N_22957,N_22126,N_22270);
or U22958 (N_22958,N_22241,N_22008);
or U22959 (N_22959,N_22046,N_22038);
and U22960 (N_22960,N_22169,N_22081);
nand U22961 (N_22961,N_22286,N_22412);
or U22962 (N_22962,N_22054,N_22316);
nand U22963 (N_22963,N_22386,N_22098);
nand U22964 (N_22964,N_22298,N_22381);
nor U22965 (N_22965,N_22488,N_22478);
nor U22966 (N_22966,N_22011,N_22091);
nand U22967 (N_22967,N_22407,N_22462);
xor U22968 (N_22968,N_22114,N_22248);
nor U22969 (N_22969,N_22167,N_22081);
and U22970 (N_22970,N_22087,N_22086);
nand U22971 (N_22971,N_22306,N_22290);
or U22972 (N_22972,N_22224,N_22345);
and U22973 (N_22973,N_22165,N_22085);
nand U22974 (N_22974,N_22285,N_22301);
nand U22975 (N_22975,N_22065,N_22314);
nor U22976 (N_22976,N_22238,N_22144);
or U22977 (N_22977,N_22474,N_22281);
xnor U22978 (N_22978,N_22146,N_22090);
or U22979 (N_22979,N_22292,N_22096);
and U22980 (N_22980,N_22359,N_22006);
xnor U22981 (N_22981,N_22445,N_22259);
nand U22982 (N_22982,N_22198,N_22440);
or U22983 (N_22983,N_22153,N_22052);
nor U22984 (N_22984,N_22112,N_22458);
nor U22985 (N_22985,N_22065,N_22308);
nor U22986 (N_22986,N_22220,N_22288);
or U22987 (N_22987,N_22256,N_22367);
nor U22988 (N_22988,N_22216,N_22479);
and U22989 (N_22989,N_22390,N_22185);
nand U22990 (N_22990,N_22433,N_22176);
and U22991 (N_22991,N_22498,N_22323);
nand U22992 (N_22992,N_22434,N_22462);
xnor U22993 (N_22993,N_22457,N_22254);
or U22994 (N_22994,N_22193,N_22484);
xnor U22995 (N_22995,N_22110,N_22187);
xor U22996 (N_22996,N_22472,N_22300);
nor U22997 (N_22997,N_22462,N_22089);
xnor U22998 (N_22998,N_22052,N_22348);
and U22999 (N_22999,N_22258,N_22229);
and U23000 (N_23000,N_22858,N_22921);
or U23001 (N_23001,N_22922,N_22866);
xor U23002 (N_23002,N_22729,N_22935);
nand U23003 (N_23003,N_22779,N_22513);
nand U23004 (N_23004,N_22524,N_22792);
nor U23005 (N_23005,N_22506,N_22931);
nor U23006 (N_23006,N_22679,N_22548);
or U23007 (N_23007,N_22791,N_22592);
or U23008 (N_23008,N_22528,N_22938);
and U23009 (N_23009,N_22706,N_22811);
nand U23010 (N_23010,N_22633,N_22560);
nand U23011 (N_23011,N_22957,N_22596);
nand U23012 (N_23012,N_22700,N_22508);
nand U23013 (N_23013,N_22683,N_22650);
and U23014 (N_23014,N_22972,N_22542);
nand U23015 (N_23015,N_22517,N_22704);
nor U23016 (N_23016,N_22607,N_22887);
or U23017 (N_23017,N_22876,N_22603);
nand U23018 (N_23018,N_22881,N_22762);
and U23019 (N_23019,N_22557,N_22971);
or U23020 (N_23020,N_22622,N_22813);
nor U23021 (N_23021,N_22702,N_22979);
or U23022 (N_23022,N_22997,N_22719);
xor U23023 (N_23023,N_22527,N_22711);
xor U23024 (N_23024,N_22894,N_22849);
or U23025 (N_23025,N_22657,N_22751);
and U23026 (N_23026,N_22944,N_22757);
or U23027 (N_23027,N_22746,N_22594);
nor U23028 (N_23028,N_22768,N_22648);
nand U23029 (N_23029,N_22776,N_22816);
nor U23030 (N_23030,N_22896,N_22807);
xor U23031 (N_23031,N_22755,N_22786);
nand U23032 (N_23032,N_22736,N_22758);
nand U23033 (N_23033,N_22580,N_22684);
xnor U23034 (N_23034,N_22628,N_22617);
and U23035 (N_23035,N_22664,N_22604);
nor U23036 (N_23036,N_22649,N_22593);
xnor U23037 (N_23037,N_22843,N_22629);
and U23038 (N_23038,N_22999,N_22728);
or U23039 (N_23039,N_22698,N_22837);
nor U23040 (N_23040,N_22828,N_22605);
xor U23041 (N_23041,N_22609,N_22988);
and U23042 (N_23042,N_22942,N_22774);
nand U23043 (N_23043,N_22533,N_22920);
nor U23044 (N_23044,N_22611,N_22620);
nor U23045 (N_23045,N_22785,N_22500);
or U23046 (N_23046,N_22985,N_22818);
and U23047 (N_23047,N_22636,N_22632);
or U23048 (N_23048,N_22602,N_22903);
and U23049 (N_23049,N_22529,N_22968);
nand U23050 (N_23050,N_22678,N_22518);
and U23051 (N_23051,N_22685,N_22502);
nand U23052 (N_23052,N_22720,N_22731);
or U23053 (N_23053,N_22770,N_22898);
nor U23054 (N_23054,N_22950,N_22760);
nor U23055 (N_23055,N_22616,N_22914);
nor U23056 (N_23056,N_22676,N_22745);
nor U23057 (N_23057,N_22638,N_22544);
nor U23058 (N_23058,N_22927,N_22627);
xnor U23059 (N_23059,N_22515,N_22589);
nor U23060 (N_23060,N_22565,N_22850);
or U23061 (N_23061,N_22802,N_22952);
and U23062 (N_23062,N_22724,N_22530);
and U23063 (N_23063,N_22918,N_22913);
nor U23064 (N_23064,N_22998,N_22710);
xor U23065 (N_23065,N_22939,N_22868);
or U23066 (N_23066,N_22709,N_22695);
nor U23067 (N_23067,N_22672,N_22897);
nand U23068 (N_23068,N_22582,N_22579);
nand U23069 (N_23069,N_22608,N_22925);
xor U23070 (N_23070,N_22847,N_22715);
nand U23071 (N_23071,N_22996,N_22919);
nand U23072 (N_23072,N_22688,N_22916);
xnor U23073 (N_23073,N_22839,N_22960);
nand U23074 (N_23074,N_22738,N_22783);
and U23075 (N_23075,N_22795,N_22781);
nor U23076 (N_23076,N_22835,N_22651);
xnor U23077 (N_23077,N_22808,N_22780);
nor U23078 (N_23078,N_22778,N_22521);
nor U23079 (N_23079,N_22965,N_22567);
nand U23080 (N_23080,N_22964,N_22930);
nand U23081 (N_23081,N_22507,N_22976);
or U23082 (N_23082,N_22810,N_22573);
xor U23083 (N_23083,N_22665,N_22687);
or U23084 (N_23084,N_22949,N_22547);
xnor U23085 (N_23085,N_22559,N_22578);
or U23086 (N_23086,N_22563,N_22987);
nand U23087 (N_23087,N_22519,N_22825);
xnor U23088 (N_23088,N_22819,N_22618);
nand U23089 (N_23089,N_22993,N_22644);
nor U23090 (N_23090,N_22884,N_22569);
nand U23091 (N_23091,N_22872,N_22955);
or U23092 (N_23092,N_22788,N_22861);
xnor U23093 (N_23093,N_22973,N_22697);
xnor U23094 (N_23094,N_22851,N_22984);
and U23095 (N_23095,N_22641,N_22734);
or U23096 (N_23096,N_22646,N_22862);
nand U23097 (N_23097,N_22540,N_22550);
nor U23098 (N_23098,N_22994,N_22765);
xnor U23099 (N_23099,N_22782,N_22653);
xor U23100 (N_23100,N_22800,N_22798);
nor U23101 (N_23101,N_22926,N_22889);
xnor U23102 (N_23102,N_22552,N_22553);
xor U23103 (N_23103,N_22662,N_22936);
nor U23104 (N_23104,N_22891,N_22566);
nand U23105 (N_23105,N_22686,N_22789);
nand U23106 (N_23106,N_22990,N_22943);
or U23107 (N_23107,N_22630,N_22784);
or U23108 (N_23108,N_22883,N_22947);
nor U23109 (N_23109,N_22621,N_22701);
nand U23110 (N_23110,N_22767,N_22848);
or U23111 (N_23111,N_22805,N_22829);
nor U23112 (N_23112,N_22820,N_22631);
and U23113 (N_23113,N_22860,N_22836);
and U23114 (N_23114,N_22655,N_22771);
nor U23115 (N_23115,N_22725,N_22674);
nor U23116 (N_23116,N_22723,N_22708);
and U23117 (N_23117,N_22536,N_22954);
xnor U23118 (N_23118,N_22908,N_22714);
nand U23119 (N_23119,N_22525,N_22899);
or U23120 (N_23120,N_22904,N_22977);
nor U23121 (N_23121,N_22945,N_22556);
xnor U23122 (N_23122,N_22934,N_22777);
nand U23123 (N_23123,N_22859,N_22703);
nand U23124 (N_23124,N_22880,N_22895);
and U23125 (N_23125,N_22743,N_22871);
nor U23126 (N_23126,N_22575,N_22591);
nor U23127 (N_23127,N_22598,N_22753);
nor U23128 (N_23128,N_22915,N_22982);
and U23129 (N_23129,N_22970,N_22614);
xnor U23130 (N_23130,N_22824,N_22523);
and U23131 (N_23131,N_22727,N_22772);
nand U23132 (N_23132,N_22796,N_22750);
or U23133 (N_23133,N_22863,N_22948);
nor U23134 (N_23134,N_22585,N_22561);
nand U23135 (N_23135,N_22804,N_22832);
or U23136 (N_23136,N_22877,N_22551);
and U23137 (N_23137,N_22509,N_22534);
or U23138 (N_23138,N_22873,N_22831);
nor U23139 (N_23139,N_22726,N_22597);
nand U23140 (N_23140,N_22639,N_22992);
nor U23141 (N_23141,N_22692,N_22554);
nor U23142 (N_23142,N_22748,N_22989);
or U23143 (N_23143,N_22787,N_22577);
nor U23144 (N_23144,N_22923,N_22867);
or U23145 (N_23145,N_22924,N_22546);
and U23146 (N_23146,N_22713,N_22969);
nand U23147 (N_23147,N_22503,N_22911);
xor U23148 (N_23148,N_22857,N_22535);
nor U23149 (N_23149,N_22574,N_22600);
nor U23150 (N_23150,N_22537,N_22512);
nand U23151 (N_23151,N_22716,N_22652);
xnor U23152 (N_23152,N_22610,N_22742);
xnor U23153 (N_23153,N_22599,N_22681);
xor U23154 (N_23154,N_22689,N_22531);
xor U23155 (N_23155,N_22659,N_22673);
and U23156 (N_23156,N_22626,N_22658);
or U23157 (N_23157,N_22888,N_22510);
nand U23158 (N_23158,N_22606,N_22739);
xnor U23159 (N_23159,N_22654,N_22830);
and U23160 (N_23160,N_22730,N_22959);
nand U23161 (N_23161,N_22583,N_22613);
and U23162 (N_23162,N_22669,N_22840);
nand U23163 (N_23163,N_22951,N_22846);
nand U23164 (N_23164,N_22761,N_22937);
nor U23165 (N_23165,N_22826,N_22907);
and U23166 (N_23166,N_22838,N_22623);
or U23167 (N_23167,N_22526,N_22568);
nand U23168 (N_23168,N_22667,N_22775);
and U23169 (N_23169,N_22961,N_22893);
nand U23170 (N_23170,N_22680,N_22735);
nand U23171 (N_23171,N_22545,N_22834);
xnor U23172 (N_23172,N_22815,N_22752);
and U23173 (N_23173,N_22797,N_22675);
or U23174 (N_23174,N_22699,N_22995);
and U23175 (N_23175,N_22974,N_22590);
nor U23176 (N_23176,N_22615,N_22940);
xor U23177 (N_23177,N_22640,N_22928);
or U23178 (N_23178,N_22690,N_22754);
or U23179 (N_23179,N_22549,N_22647);
nor U23180 (N_23180,N_22890,N_22522);
nand U23181 (N_23181,N_22801,N_22817);
or U23182 (N_23182,N_22759,N_22842);
and U23183 (N_23183,N_22747,N_22929);
and U23184 (N_23184,N_22538,N_22769);
xnor U23185 (N_23185,N_22696,N_22744);
nor U23186 (N_23186,N_22886,N_22809);
and U23187 (N_23187,N_22666,N_22645);
and U23188 (N_23188,N_22763,N_22885);
or U23189 (N_23189,N_22571,N_22793);
xnor U23190 (N_23190,N_22511,N_22933);
nand U23191 (N_23191,N_22790,N_22584);
nand U23192 (N_23192,N_22705,N_22981);
and U23193 (N_23193,N_22588,N_22514);
nand U23194 (N_23194,N_22878,N_22660);
nor U23195 (N_23195,N_22543,N_22587);
and U23196 (N_23196,N_22682,N_22991);
or U23197 (N_23197,N_22501,N_22879);
and U23198 (N_23198,N_22677,N_22827);
xnor U23199 (N_23199,N_22595,N_22721);
nor U23200 (N_23200,N_22656,N_22794);
xnor U23201 (N_23201,N_22741,N_22882);
and U23202 (N_23202,N_22975,N_22668);
or U23203 (N_23203,N_22856,N_22956);
or U23204 (N_23204,N_22740,N_22852);
xor U23205 (N_23205,N_22912,N_22845);
or U23206 (N_23206,N_22901,N_22986);
nand U23207 (N_23207,N_22576,N_22821);
xnor U23208 (N_23208,N_22624,N_22691);
nor U23209 (N_23209,N_22865,N_22516);
or U23210 (N_23210,N_22764,N_22844);
and U23211 (N_23211,N_22558,N_22718);
or U23212 (N_23212,N_22661,N_22637);
nand U23213 (N_23213,N_22539,N_22833);
nand U23214 (N_23214,N_22505,N_22823);
nand U23215 (N_23215,N_22962,N_22773);
nor U23216 (N_23216,N_22946,N_22642);
nand U23217 (N_23217,N_22814,N_22841);
nor U23218 (N_23218,N_22555,N_22900);
nor U23219 (N_23219,N_22853,N_22693);
or U23220 (N_23220,N_22932,N_22733);
or U23221 (N_23221,N_22581,N_22917);
or U23222 (N_23222,N_22619,N_22756);
or U23223 (N_23223,N_22803,N_22905);
nor U23224 (N_23224,N_22707,N_22906);
nor U23225 (N_23225,N_22564,N_22874);
xnor U23226 (N_23226,N_22967,N_22966);
nor U23227 (N_23227,N_22570,N_22799);
nand U23228 (N_23228,N_22712,N_22812);
nor U23229 (N_23229,N_22562,N_22963);
xor U23230 (N_23230,N_22635,N_22854);
nor U23231 (N_23231,N_22806,N_22910);
nor U23232 (N_23232,N_22902,N_22612);
nor U23233 (N_23233,N_22541,N_22983);
and U23234 (N_23234,N_22855,N_22663);
and U23235 (N_23235,N_22892,N_22601);
or U23236 (N_23236,N_22980,N_22941);
or U23237 (N_23237,N_22520,N_22766);
nor U23238 (N_23238,N_22953,N_22749);
xnor U23239 (N_23239,N_22870,N_22909);
nor U23240 (N_23240,N_22978,N_22732);
and U23241 (N_23241,N_22625,N_22694);
nand U23242 (N_23242,N_22717,N_22958);
or U23243 (N_23243,N_22586,N_22671);
xor U23244 (N_23244,N_22875,N_22822);
xnor U23245 (N_23245,N_22504,N_22864);
nand U23246 (N_23246,N_22634,N_22643);
xor U23247 (N_23247,N_22737,N_22722);
or U23248 (N_23248,N_22532,N_22670);
or U23249 (N_23249,N_22869,N_22572);
nand U23250 (N_23250,N_22922,N_22892);
nand U23251 (N_23251,N_22691,N_22829);
nand U23252 (N_23252,N_22572,N_22633);
xor U23253 (N_23253,N_22968,N_22763);
or U23254 (N_23254,N_22698,N_22802);
or U23255 (N_23255,N_22622,N_22822);
nor U23256 (N_23256,N_22703,N_22727);
xor U23257 (N_23257,N_22553,N_22905);
or U23258 (N_23258,N_22964,N_22572);
nand U23259 (N_23259,N_22840,N_22771);
nand U23260 (N_23260,N_22631,N_22648);
or U23261 (N_23261,N_22712,N_22918);
or U23262 (N_23262,N_22667,N_22539);
xor U23263 (N_23263,N_22843,N_22657);
xnor U23264 (N_23264,N_22746,N_22710);
and U23265 (N_23265,N_22810,N_22621);
and U23266 (N_23266,N_22638,N_22915);
xor U23267 (N_23267,N_22795,N_22906);
nand U23268 (N_23268,N_22909,N_22825);
nor U23269 (N_23269,N_22853,N_22941);
or U23270 (N_23270,N_22762,N_22896);
and U23271 (N_23271,N_22679,N_22610);
and U23272 (N_23272,N_22740,N_22769);
and U23273 (N_23273,N_22923,N_22918);
nor U23274 (N_23274,N_22640,N_22566);
nor U23275 (N_23275,N_22651,N_22518);
nand U23276 (N_23276,N_22901,N_22979);
nand U23277 (N_23277,N_22643,N_22895);
or U23278 (N_23278,N_22817,N_22536);
or U23279 (N_23279,N_22502,N_22944);
and U23280 (N_23280,N_22662,N_22733);
xnor U23281 (N_23281,N_22985,N_22988);
nor U23282 (N_23282,N_22514,N_22811);
and U23283 (N_23283,N_22635,N_22542);
nor U23284 (N_23284,N_22951,N_22699);
nand U23285 (N_23285,N_22545,N_22989);
and U23286 (N_23286,N_22857,N_22673);
xor U23287 (N_23287,N_22705,N_22956);
nand U23288 (N_23288,N_22987,N_22564);
nand U23289 (N_23289,N_22508,N_22948);
nor U23290 (N_23290,N_22784,N_22918);
or U23291 (N_23291,N_22511,N_22642);
nor U23292 (N_23292,N_22805,N_22791);
or U23293 (N_23293,N_22689,N_22982);
nand U23294 (N_23294,N_22860,N_22905);
xor U23295 (N_23295,N_22537,N_22737);
xnor U23296 (N_23296,N_22598,N_22749);
nand U23297 (N_23297,N_22704,N_22726);
nor U23298 (N_23298,N_22994,N_22881);
or U23299 (N_23299,N_22774,N_22550);
xor U23300 (N_23300,N_22553,N_22977);
nand U23301 (N_23301,N_22973,N_22946);
and U23302 (N_23302,N_22620,N_22742);
nand U23303 (N_23303,N_22687,N_22965);
xor U23304 (N_23304,N_22747,N_22902);
nand U23305 (N_23305,N_22811,N_22789);
nand U23306 (N_23306,N_22543,N_22879);
xnor U23307 (N_23307,N_22882,N_22994);
nand U23308 (N_23308,N_22528,N_22569);
and U23309 (N_23309,N_22642,N_22542);
nand U23310 (N_23310,N_22592,N_22608);
nor U23311 (N_23311,N_22752,N_22952);
or U23312 (N_23312,N_22925,N_22529);
and U23313 (N_23313,N_22552,N_22516);
xor U23314 (N_23314,N_22979,N_22545);
xnor U23315 (N_23315,N_22563,N_22510);
or U23316 (N_23316,N_22836,N_22650);
nand U23317 (N_23317,N_22912,N_22947);
nand U23318 (N_23318,N_22970,N_22597);
or U23319 (N_23319,N_22547,N_22944);
nor U23320 (N_23320,N_22689,N_22734);
nor U23321 (N_23321,N_22882,N_22677);
or U23322 (N_23322,N_22633,N_22797);
nor U23323 (N_23323,N_22787,N_22667);
or U23324 (N_23324,N_22578,N_22871);
or U23325 (N_23325,N_22808,N_22965);
and U23326 (N_23326,N_22818,N_22535);
and U23327 (N_23327,N_22610,N_22654);
and U23328 (N_23328,N_22991,N_22671);
or U23329 (N_23329,N_22573,N_22556);
and U23330 (N_23330,N_22944,N_22932);
or U23331 (N_23331,N_22938,N_22761);
nor U23332 (N_23332,N_22872,N_22656);
nand U23333 (N_23333,N_22627,N_22716);
or U23334 (N_23334,N_22615,N_22601);
nand U23335 (N_23335,N_22529,N_22565);
nor U23336 (N_23336,N_22746,N_22657);
nor U23337 (N_23337,N_22842,N_22764);
or U23338 (N_23338,N_22818,N_22872);
xnor U23339 (N_23339,N_22817,N_22986);
xor U23340 (N_23340,N_22576,N_22809);
nor U23341 (N_23341,N_22689,N_22695);
nand U23342 (N_23342,N_22894,N_22679);
nand U23343 (N_23343,N_22525,N_22682);
nor U23344 (N_23344,N_22856,N_22518);
or U23345 (N_23345,N_22905,N_22571);
xor U23346 (N_23346,N_22528,N_22745);
and U23347 (N_23347,N_22922,N_22862);
and U23348 (N_23348,N_22900,N_22757);
nor U23349 (N_23349,N_22804,N_22624);
xor U23350 (N_23350,N_22930,N_22560);
and U23351 (N_23351,N_22562,N_22546);
xor U23352 (N_23352,N_22755,N_22734);
nand U23353 (N_23353,N_22953,N_22965);
or U23354 (N_23354,N_22649,N_22500);
nor U23355 (N_23355,N_22940,N_22922);
and U23356 (N_23356,N_22948,N_22820);
xnor U23357 (N_23357,N_22995,N_22624);
or U23358 (N_23358,N_22816,N_22630);
and U23359 (N_23359,N_22958,N_22779);
or U23360 (N_23360,N_22923,N_22745);
or U23361 (N_23361,N_22789,N_22631);
and U23362 (N_23362,N_22590,N_22768);
nand U23363 (N_23363,N_22623,N_22616);
and U23364 (N_23364,N_22849,N_22955);
xor U23365 (N_23365,N_22845,N_22595);
xor U23366 (N_23366,N_22716,N_22759);
and U23367 (N_23367,N_22722,N_22538);
or U23368 (N_23368,N_22673,N_22950);
nor U23369 (N_23369,N_22601,N_22747);
nor U23370 (N_23370,N_22660,N_22681);
nor U23371 (N_23371,N_22801,N_22559);
or U23372 (N_23372,N_22713,N_22843);
and U23373 (N_23373,N_22836,N_22977);
xnor U23374 (N_23374,N_22744,N_22848);
and U23375 (N_23375,N_22749,N_22675);
nand U23376 (N_23376,N_22528,N_22509);
xnor U23377 (N_23377,N_22964,N_22980);
or U23378 (N_23378,N_22782,N_22596);
nor U23379 (N_23379,N_22931,N_22987);
nor U23380 (N_23380,N_22538,N_22830);
nor U23381 (N_23381,N_22805,N_22848);
xor U23382 (N_23382,N_22831,N_22580);
nor U23383 (N_23383,N_22877,N_22845);
nor U23384 (N_23384,N_22768,N_22938);
or U23385 (N_23385,N_22797,N_22783);
or U23386 (N_23386,N_22529,N_22864);
nand U23387 (N_23387,N_22595,N_22522);
and U23388 (N_23388,N_22500,N_22745);
nand U23389 (N_23389,N_22891,N_22676);
xnor U23390 (N_23390,N_22548,N_22798);
nand U23391 (N_23391,N_22956,N_22758);
or U23392 (N_23392,N_22817,N_22505);
or U23393 (N_23393,N_22533,N_22586);
xor U23394 (N_23394,N_22738,N_22676);
nand U23395 (N_23395,N_22687,N_22931);
nand U23396 (N_23396,N_22608,N_22947);
xnor U23397 (N_23397,N_22851,N_22980);
or U23398 (N_23398,N_22595,N_22558);
xnor U23399 (N_23399,N_22606,N_22930);
nor U23400 (N_23400,N_22827,N_22623);
nand U23401 (N_23401,N_22913,N_22827);
nor U23402 (N_23402,N_22902,N_22734);
xnor U23403 (N_23403,N_22783,N_22548);
nand U23404 (N_23404,N_22949,N_22763);
nand U23405 (N_23405,N_22577,N_22865);
nand U23406 (N_23406,N_22648,N_22500);
xor U23407 (N_23407,N_22526,N_22963);
or U23408 (N_23408,N_22816,N_22612);
and U23409 (N_23409,N_22625,N_22904);
nand U23410 (N_23410,N_22729,N_22777);
xor U23411 (N_23411,N_22870,N_22762);
nand U23412 (N_23412,N_22519,N_22718);
nand U23413 (N_23413,N_22540,N_22996);
and U23414 (N_23414,N_22536,N_22782);
nor U23415 (N_23415,N_22555,N_22948);
xor U23416 (N_23416,N_22691,N_22904);
nor U23417 (N_23417,N_22727,N_22650);
or U23418 (N_23418,N_22663,N_22659);
nand U23419 (N_23419,N_22819,N_22799);
and U23420 (N_23420,N_22958,N_22553);
or U23421 (N_23421,N_22721,N_22776);
or U23422 (N_23422,N_22590,N_22975);
nor U23423 (N_23423,N_22830,N_22999);
or U23424 (N_23424,N_22767,N_22917);
nor U23425 (N_23425,N_22884,N_22959);
xnor U23426 (N_23426,N_22955,N_22589);
xor U23427 (N_23427,N_22898,N_22570);
or U23428 (N_23428,N_22807,N_22960);
nor U23429 (N_23429,N_22938,N_22529);
and U23430 (N_23430,N_22892,N_22501);
or U23431 (N_23431,N_22764,N_22685);
or U23432 (N_23432,N_22832,N_22656);
or U23433 (N_23433,N_22886,N_22595);
nor U23434 (N_23434,N_22861,N_22627);
nor U23435 (N_23435,N_22824,N_22886);
nand U23436 (N_23436,N_22618,N_22811);
or U23437 (N_23437,N_22547,N_22728);
xnor U23438 (N_23438,N_22838,N_22682);
xor U23439 (N_23439,N_22603,N_22901);
xnor U23440 (N_23440,N_22744,N_22752);
nand U23441 (N_23441,N_22720,N_22967);
and U23442 (N_23442,N_22855,N_22727);
and U23443 (N_23443,N_22968,N_22701);
or U23444 (N_23444,N_22819,N_22717);
nand U23445 (N_23445,N_22978,N_22532);
nor U23446 (N_23446,N_22984,N_22798);
and U23447 (N_23447,N_22768,N_22610);
nand U23448 (N_23448,N_22699,N_22615);
xnor U23449 (N_23449,N_22546,N_22680);
and U23450 (N_23450,N_22834,N_22956);
xor U23451 (N_23451,N_22834,N_22532);
nand U23452 (N_23452,N_22892,N_22957);
xor U23453 (N_23453,N_22821,N_22726);
xor U23454 (N_23454,N_22763,N_22981);
nor U23455 (N_23455,N_22557,N_22961);
nand U23456 (N_23456,N_22709,N_22542);
nand U23457 (N_23457,N_22896,N_22624);
or U23458 (N_23458,N_22714,N_22506);
and U23459 (N_23459,N_22770,N_22792);
and U23460 (N_23460,N_22677,N_22777);
and U23461 (N_23461,N_22774,N_22599);
or U23462 (N_23462,N_22989,N_22578);
xor U23463 (N_23463,N_22695,N_22818);
or U23464 (N_23464,N_22546,N_22826);
nor U23465 (N_23465,N_22532,N_22869);
and U23466 (N_23466,N_22751,N_22628);
or U23467 (N_23467,N_22546,N_22660);
nand U23468 (N_23468,N_22549,N_22925);
xnor U23469 (N_23469,N_22919,N_22619);
nand U23470 (N_23470,N_22612,N_22652);
or U23471 (N_23471,N_22685,N_22969);
xor U23472 (N_23472,N_22593,N_22962);
xor U23473 (N_23473,N_22806,N_22580);
and U23474 (N_23474,N_22913,N_22886);
xnor U23475 (N_23475,N_22802,N_22870);
or U23476 (N_23476,N_22604,N_22854);
nor U23477 (N_23477,N_22589,N_22648);
and U23478 (N_23478,N_22582,N_22920);
and U23479 (N_23479,N_22928,N_22681);
nor U23480 (N_23480,N_22708,N_22948);
or U23481 (N_23481,N_22527,N_22851);
nand U23482 (N_23482,N_22570,N_22546);
or U23483 (N_23483,N_22517,N_22508);
xor U23484 (N_23484,N_22579,N_22910);
nand U23485 (N_23485,N_22599,N_22953);
xor U23486 (N_23486,N_22765,N_22561);
and U23487 (N_23487,N_22565,N_22537);
xnor U23488 (N_23488,N_22701,N_22535);
or U23489 (N_23489,N_22866,N_22782);
or U23490 (N_23490,N_22593,N_22752);
nand U23491 (N_23491,N_22668,N_22764);
nor U23492 (N_23492,N_22663,N_22846);
nor U23493 (N_23493,N_22615,N_22686);
xnor U23494 (N_23494,N_22870,N_22960);
xor U23495 (N_23495,N_22897,N_22809);
xor U23496 (N_23496,N_22682,N_22677);
nand U23497 (N_23497,N_22781,N_22747);
or U23498 (N_23498,N_22687,N_22752);
or U23499 (N_23499,N_22969,N_22634);
or U23500 (N_23500,N_23129,N_23392);
nand U23501 (N_23501,N_23202,N_23370);
xor U23502 (N_23502,N_23314,N_23347);
or U23503 (N_23503,N_23003,N_23442);
xnor U23504 (N_23504,N_23371,N_23061);
nand U23505 (N_23505,N_23119,N_23391);
and U23506 (N_23506,N_23486,N_23215);
xor U23507 (N_23507,N_23039,N_23007);
or U23508 (N_23508,N_23141,N_23151);
nor U23509 (N_23509,N_23170,N_23335);
and U23510 (N_23510,N_23208,N_23341);
nor U23511 (N_23511,N_23269,N_23225);
or U23512 (N_23512,N_23136,N_23477);
xor U23513 (N_23513,N_23374,N_23142);
or U23514 (N_23514,N_23196,N_23465);
and U23515 (N_23515,N_23248,N_23333);
nand U23516 (N_23516,N_23143,N_23016);
or U23517 (N_23517,N_23033,N_23308);
nand U23518 (N_23518,N_23412,N_23020);
xor U23519 (N_23519,N_23177,N_23176);
or U23520 (N_23520,N_23309,N_23073);
nor U23521 (N_23521,N_23031,N_23226);
xnor U23522 (N_23522,N_23022,N_23419);
or U23523 (N_23523,N_23153,N_23005);
or U23524 (N_23524,N_23305,N_23366);
nor U23525 (N_23525,N_23490,N_23461);
xor U23526 (N_23526,N_23244,N_23476);
and U23527 (N_23527,N_23279,N_23071);
xor U23528 (N_23528,N_23012,N_23349);
xnor U23529 (N_23529,N_23014,N_23250);
and U23530 (N_23530,N_23032,N_23369);
and U23531 (N_23531,N_23413,N_23043);
or U23532 (N_23532,N_23154,N_23418);
nand U23533 (N_23533,N_23066,N_23409);
nor U23534 (N_23534,N_23259,N_23346);
xnor U23535 (N_23535,N_23009,N_23132);
nand U23536 (N_23536,N_23275,N_23240);
or U23537 (N_23537,N_23090,N_23284);
xor U23538 (N_23538,N_23239,N_23188);
or U23539 (N_23539,N_23040,N_23258);
or U23540 (N_23540,N_23048,N_23357);
nand U23541 (N_23541,N_23289,N_23420);
xor U23542 (N_23542,N_23292,N_23303);
or U23543 (N_23543,N_23446,N_23311);
and U23544 (N_23544,N_23382,N_23107);
nand U23545 (N_23545,N_23232,N_23015);
or U23546 (N_23546,N_23011,N_23381);
or U23547 (N_23547,N_23192,N_23120);
and U23548 (N_23548,N_23281,N_23114);
nor U23549 (N_23549,N_23000,N_23029);
nand U23550 (N_23550,N_23023,N_23220);
nand U23551 (N_23551,N_23463,N_23488);
nor U23552 (N_23552,N_23448,N_23222);
or U23553 (N_23553,N_23408,N_23415);
nor U23554 (N_23554,N_23169,N_23312);
and U23555 (N_23555,N_23199,N_23326);
or U23556 (N_23556,N_23484,N_23320);
xnor U23557 (N_23557,N_23152,N_23037);
or U23558 (N_23558,N_23173,N_23083);
nor U23559 (N_23559,N_23236,N_23495);
xor U23560 (N_23560,N_23057,N_23283);
nand U23561 (N_23561,N_23301,N_23254);
or U23562 (N_23562,N_23462,N_23110);
nor U23563 (N_23563,N_23439,N_23430);
and U23564 (N_23564,N_23055,N_23316);
nand U23565 (N_23565,N_23195,N_23358);
xor U23566 (N_23566,N_23267,N_23424);
xor U23567 (N_23567,N_23051,N_23416);
nor U23568 (N_23568,N_23296,N_23332);
xnor U23569 (N_23569,N_23046,N_23181);
or U23570 (N_23570,N_23001,N_23218);
nand U23571 (N_23571,N_23214,N_23013);
or U23572 (N_23572,N_23386,N_23148);
nand U23573 (N_23573,N_23004,N_23124);
or U23574 (N_23574,N_23323,N_23200);
xor U23575 (N_23575,N_23111,N_23094);
and U23576 (N_23576,N_23479,N_23102);
nand U23577 (N_23577,N_23487,N_23231);
nor U23578 (N_23578,N_23384,N_23451);
nand U23579 (N_23579,N_23079,N_23454);
nor U23580 (N_23580,N_23118,N_23441);
nor U23581 (N_23581,N_23262,N_23298);
nand U23582 (N_23582,N_23393,N_23185);
nor U23583 (N_23583,N_23489,N_23466);
or U23584 (N_23584,N_23134,N_23460);
nor U23585 (N_23585,N_23087,N_23198);
or U23586 (N_23586,N_23457,N_23359);
and U23587 (N_23587,N_23445,N_23427);
nor U23588 (N_23588,N_23189,N_23274);
nand U23589 (N_23589,N_23131,N_23163);
and U23590 (N_23590,N_23184,N_23045);
xnor U23591 (N_23591,N_23260,N_23078);
xnor U23592 (N_23592,N_23186,N_23036);
nand U23593 (N_23593,N_23315,N_23276);
xor U23594 (N_23594,N_23426,N_23191);
nand U23595 (N_23595,N_23336,N_23287);
nor U23596 (N_23596,N_23054,N_23130);
or U23597 (N_23597,N_23128,N_23104);
nand U23598 (N_23598,N_23331,N_23383);
xnor U23599 (N_23599,N_23449,N_23273);
nor U23600 (N_23600,N_23174,N_23085);
or U23601 (N_23601,N_23389,N_23237);
xor U23602 (N_23602,N_23021,N_23318);
and U23603 (N_23603,N_23024,N_23277);
nor U23604 (N_23604,N_23150,N_23388);
nand U23605 (N_23605,N_23362,N_23084);
and U23606 (N_23606,N_23027,N_23076);
and U23607 (N_23607,N_23405,N_23182);
nand U23608 (N_23608,N_23069,N_23330);
or U23609 (N_23609,N_23035,N_23140);
or U23610 (N_23610,N_23178,N_23355);
or U23611 (N_23611,N_23253,N_23172);
nand U23612 (N_23612,N_23478,N_23086);
nor U23613 (N_23613,N_23068,N_23394);
or U23614 (N_23614,N_23437,N_23300);
nand U23615 (N_23615,N_23204,N_23497);
and U23616 (N_23616,N_23286,N_23146);
xnor U23617 (N_23617,N_23459,N_23443);
and U23618 (N_23618,N_23180,N_23127);
nand U23619 (N_23619,N_23411,N_23351);
nand U23620 (N_23620,N_23288,N_23241);
nor U23621 (N_23621,N_23377,N_23455);
and U23622 (N_23622,N_23428,N_23444);
and U23623 (N_23623,N_23352,N_23155);
xnor U23624 (N_23624,N_23203,N_23100);
or U23625 (N_23625,N_23266,N_23270);
or U23626 (N_23626,N_23268,N_23211);
or U23627 (N_23627,N_23414,N_23160);
nor U23628 (N_23628,N_23390,N_23157);
nor U23629 (N_23629,N_23089,N_23207);
nor U23630 (N_23630,N_23356,N_23217);
xnor U23631 (N_23631,N_23480,N_23285);
and U23632 (N_23632,N_23025,N_23280);
nor U23633 (N_23633,N_23229,N_23201);
xor U23634 (N_23634,N_23272,N_23345);
nand U23635 (N_23635,N_23363,N_23247);
nand U23636 (N_23636,N_23385,N_23395);
nor U23637 (N_23637,N_23145,N_23434);
nand U23638 (N_23638,N_23194,N_23494);
nand U23639 (N_23639,N_23167,N_23026);
and U23640 (N_23640,N_23321,N_23492);
xnor U23641 (N_23641,N_23493,N_23337);
or U23642 (N_23642,N_23242,N_23469);
xnor U23643 (N_23643,N_23334,N_23233);
nand U23644 (N_23644,N_23103,N_23081);
nor U23645 (N_23645,N_23325,N_23041);
or U23646 (N_23646,N_23062,N_23473);
nor U23647 (N_23647,N_23075,N_23179);
or U23648 (N_23648,N_23397,N_23246);
nor U23649 (N_23649,N_23396,N_23453);
or U23650 (N_23650,N_23158,N_23126);
nand U23651 (N_23651,N_23482,N_23149);
nand U23652 (N_23652,N_23210,N_23113);
xor U23653 (N_23653,N_23044,N_23243);
nor U23654 (N_23654,N_23091,N_23304);
nand U23655 (N_23655,N_23498,N_23452);
xor U23656 (N_23656,N_23265,N_23125);
and U23657 (N_23657,N_23074,N_23400);
xor U23658 (N_23658,N_23249,N_23019);
nor U23659 (N_23659,N_23168,N_23431);
nand U23660 (N_23660,N_23213,N_23343);
nor U23661 (N_23661,N_23018,N_23438);
xor U23662 (N_23662,N_23219,N_23373);
nor U23663 (N_23663,N_23139,N_23212);
nor U23664 (N_23664,N_23399,N_23109);
nand U23665 (N_23665,N_23474,N_23067);
nand U23666 (N_23666,N_23450,N_23034);
nand U23667 (N_23667,N_23360,N_23008);
or U23668 (N_23668,N_23447,N_23324);
xor U23669 (N_23669,N_23053,N_23380);
and U23670 (N_23670,N_23271,N_23293);
or U23671 (N_23671,N_23458,N_23227);
and U23672 (N_23672,N_23425,N_23310);
xor U23673 (N_23673,N_23354,N_23407);
and U23674 (N_23674,N_23423,N_23010);
nand U23675 (N_23675,N_23297,N_23307);
or U23676 (N_23676,N_23106,N_23187);
and U23677 (N_23677,N_23166,N_23299);
nand U23678 (N_23678,N_23436,N_23230);
and U23679 (N_23679,N_23294,N_23093);
nand U23680 (N_23680,N_23162,N_23095);
nand U23681 (N_23681,N_23038,N_23077);
or U23682 (N_23682,N_23047,N_23133);
xnor U23683 (N_23683,N_23491,N_23108);
nor U23684 (N_23684,N_23499,N_23161);
xnor U23685 (N_23685,N_23209,N_23175);
xnor U23686 (N_23686,N_23368,N_23421);
or U23687 (N_23687,N_23485,N_23123);
nand U23688 (N_23688,N_23261,N_23080);
xor U23689 (N_23689,N_23252,N_23156);
or U23690 (N_23690,N_23440,N_23468);
and U23691 (N_23691,N_23238,N_23379);
nand U23692 (N_23692,N_23410,N_23295);
and U23693 (N_23693,N_23002,N_23375);
xor U23694 (N_23694,N_23245,N_23056);
xor U23695 (N_23695,N_23101,N_23344);
xor U23696 (N_23696,N_23350,N_23403);
nand U23697 (N_23697,N_23464,N_23072);
and U23698 (N_23698,N_23483,N_23313);
nor U23699 (N_23699,N_23302,N_23329);
xor U23700 (N_23700,N_23467,N_23402);
nor U23701 (N_23701,N_23098,N_23116);
or U23702 (N_23702,N_23322,N_23147);
and U23703 (N_23703,N_23205,N_23082);
or U23704 (N_23704,N_23121,N_23190);
nand U23705 (N_23705,N_23291,N_23006);
xnor U23706 (N_23706,N_23429,N_23122);
and U23707 (N_23707,N_23105,N_23052);
xor U23708 (N_23708,N_23496,N_23342);
nor U23709 (N_23709,N_23234,N_23092);
or U23710 (N_23710,N_23028,N_23099);
nor U23711 (N_23711,N_23376,N_23058);
or U23712 (N_23712,N_23137,N_23235);
nand U23713 (N_23713,N_23117,N_23481);
or U23714 (N_23714,N_23353,N_23417);
nor U23715 (N_23715,N_23206,N_23340);
or U23716 (N_23716,N_23306,N_23263);
and U23717 (N_23717,N_23197,N_23327);
nand U23718 (N_23718,N_23338,N_23317);
and U23719 (N_23719,N_23367,N_23216);
or U23720 (N_23720,N_23097,N_23435);
nor U23721 (N_23721,N_23159,N_23063);
and U23722 (N_23722,N_23433,N_23387);
nor U23723 (N_23723,N_23406,N_23183);
and U23724 (N_23724,N_23144,N_23456);
nor U23725 (N_23725,N_23088,N_23372);
and U23726 (N_23726,N_23255,N_23290);
xor U23727 (N_23727,N_23042,N_23112);
nor U23728 (N_23728,N_23165,N_23348);
and U23729 (N_23729,N_23404,N_23470);
nor U23730 (N_23730,N_23223,N_23070);
nand U23731 (N_23731,N_23050,N_23224);
or U23732 (N_23732,N_23319,N_23228);
nand U23733 (N_23733,N_23096,N_23030);
nor U23734 (N_23734,N_23115,N_23064);
xor U23735 (N_23735,N_23361,N_23065);
nand U23736 (N_23736,N_23059,N_23472);
nand U23737 (N_23737,N_23060,N_23135);
nor U23738 (N_23738,N_23339,N_23278);
nand U23739 (N_23739,N_23164,N_23398);
and U23740 (N_23740,N_23432,N_23401);
nor U23741 (N_23741,N_23471,N_23256);
or U23742 (N_23742,N_23017,N_23257);
or U23743 (N_23743,N_23365,N_23364);
nor U23744 (N_23744,N_23171,N_23193);
xnor U23745 (N_23745,N_23221,N_23138);
and U23746 (N_23746,N_23282,N_23422);
and U23747 (N_23747,N_23251,N_23264);
xnor U23748 (N_23748,N_23378,N_23475);
xnor U23749 (N_23749,N_23328,N_23049);
or U23750 (N_23750,N_23324,N_23251);
and U23751 (N_23751,N_23047,N_23382);
nor U23752 (N_23752,N_23372,N_23142);
nor U23753 (N_23753,N_23473,N_23309);
nor U23754 (N_23754,N_23479,N_23028);
xnor U23755 (N_23755,N_23196,N_23352);
nor U23756 (N_23756,N_23277,N_23336);
nand U23757 (N_23757,N_23234,N_23425);
xnor U23758 (N_23758,N_23269,N_23428);
nor U23759 (N_23759,N_23473,N_23035);
nand U23760 (N_23760,N_23174,N_23343);
or U23761 (N_23761,N_23494,N_23047);
xnor U23762 (N_23762,N_23013,N_23347);
nand U23763 (N_23763,N_23198,N_23493);
and U23764 (N_23764,N_23373,N_23254);
or U23765 (N_23765,N_23114,N_23075);
xnor U23766 (N_23766,N_23291,N_23176);
nand U23767 (N_23767,N_23000,N_23414);
or U23768 (N_23768,N_23199,N_23213);
and U23769 (N_23769,N_23258,N_23314);
nor U23770 (N_23770,N_23318,N_23218);
and U23771 (N_23771,N_23478,N_23356);
or U23772 (N_23772,N_23173,N_23020);
nor U23773 (N_23773,N_23478,N_23112);
xnor U23774 (N_23774,N_23222,N_23088);
and U23775 (N_23775,N_23374,N_23041);
and U23776 (N_23776,N_23243,N_23374);
or U23777 (N_23777,N_23154,N_23328);
or U23778 (N_23778,N_23019,N_23042);
or U23779 (N_23779,N_23379,N_23409);
and U23780 (N_23780,N_23237,N_23201);
and U23781 (N_23781,N_23087,N_23492);
xor U23782 (N_23782,N_23009,N_23030);
nor U23783 (N_23783,N_23144,N_23343);
xor U23784 (N_23784,N_23125,N_23181);
xnor U23785 (N_23785,N_23245,N_23194);
xor U23786 (N_23786,N_23069,N_23351);
and U23787 (N_23787,N_23448,N_23053);
xnor U23788 (N_23788,N_23101,N_23333);
and U23789 (N_23789,N_23325,N_23308);
or U23790 (N_23790,N_23311,N_23489);
or U23791 (N_23791,N_23190,N_23225);
xor U23792 (N_23792,N_23479,N_23191);
nand U23793 (N_23793,N_23148,N_23258);
nand U23794 (N_23794,N_23445,N_23492);
and U23795 (N_23795,N_23305,N_23187);
nor U23796 (N_23796,N_23323,N_23338);
or U23797 (N_23797,N_23031,N_23253);
nand U23798 (N_23798,N_23022,N_23012);
or U23799 (N_23799,N_23235,N_23249);
and U23800 (N_23800,N_23391,N_23229);
or U23801 (N_23801,N_23384,N_23177);
xnor U23802 (N_23802,N_23013,N_23126);
or U23803 (N_23803,N_23000,N_23217);
or U23804 (N_23804,N_23051,N_23386);
nor U23805 (N_23805,N_23224,N_23420);
nand U23806 (N_23806,N_23300,N_23097);
nand U23807 (N_23807,N_23262,N_23038);
nor U23808 (N_23808,N_23428,N_23124);
nor U23809 (N_23809,N_23426,N_23468);
and U23810 (N_23810,N_23314,N_23193);
or U23811 (N_23811,N_23045,N_23386);
xnor U23812 (N_23812,N_23275,N_23157);
nor U23813 (N_23813,N_23373,N_23479);
nor U23814 (N_23814,N_23325,N_23261);
or U23815 (N_23815,N_23319,N_23487);
and U23816 (N_23816,N_23330,N_23453);
nor U23817 (N_23817,N_23205,N_23017);
or U23818 (N_23818,N_23293,N_23422);
nor U23819 (N_23819,N_23057,N_23211);
xnor U23820 (N_23820,N_23435,N_23259);
xnor U23821 (N_23821,N_23105,N_23324);
xnor U23822 (N_23822,N_23084,N_23292);
xnor U23823 (N_23823,N_23137,N_23095);
nor U23824 (N_23824,N_23475,N_23357);
xnor U23825 (N_23825,N_23349,N_23305);
xnor U23826 (N_23826,N_23248,N_23423);
xnor U23827 (N_23827,N_23019,N_23178);
nor U23828 (N_23828,N_23025,N_23100);
nand U23829 (N_23829,N_23042,N_23194);
nor U23830 (N_23830,N_23148,N_23170);
nor U23831 (N_23831,N_23467,N_23105);
nand U23832 (N_23832,N_23259,N_23306);
nand U23833 (N_23833,N_23336,N_23224);
and U23834 (N_23834,N_23266,N_23268);
or U23835 (N_23835,N_23331,N_23435);
xor U23836 (N_23836,N_23292,N_23325);
nand U23837 (N_23837,N_23407,N_23151);
and U23838 (N_23838,N_23310,N_23156);
or U23839 (N_23839,N_23345,N_23072);
nand U23840 (N_23840,N_23494,N_23248);
xor U23841 (N_23841,N_23032,N_23008);
or U23842 (N_23842,N_23238,N_23412);
and U23843 (N_23843,N_23101,N_23493);
or U23844 (N_23844,N_23353,N_23176);
and U23845 (N_23845,N_23199,N_23483);
nor U23846 (N_23846,N_23363,N_23491);
or U23847 (N_23847,N_23440,N_23421);
and U23848 (N_23848,N_23290,N_23399);
or U23849 (N_23849,N_23325,N_23342);
and U23850 (N_23850,N_23455,N_23052);
xnor U23851 (N_23851,N_23409,N_23219);
nand U23852 (N_23852,N_23299,N_23479);
nor U23853 (N_23853,N_23268,N_23421);
xor U23854 (N_23854,N_23360,N_23091);
nand U23855 (N_23855,N_23189,N_23418);
and U23856 (N_23856,N_23459,N_23029);
or U23857 (N_23857,N_23282,N_23475);
and U23858 (N_23858,N_23133,N_23409);
and U23859 (N_23859,N_23232,N_23065);
and U23860 (N_23860,N_23203,N_23326);
nand U23861 (N_23861,N_23341,N_23081);
nand U23862 (N_23862,N_23062,N_23059);
xor U23863 (N_23863,N_23060,N_23178);
or U23864 (N_23864,N_23246,N_23139);
or U23865 (N_23865,N_23454,N_23053);
or U23866 (N_23866,N_23267,N_23191);
nand U23867 (N_23867,N_23040,N_23077);
nor U23868 (N_23868,N_23188,N_23482);
and U23869 (N_23869,N_23272,N_23112);
nand U23870 (N_23870,N_23222,N_23193);
or U23871 (N_23871,N_23340,N_23341);
nor U23872 (N_23872,N_23378,N_23481);
and U23873 (N_23873,N_23441,N_23122);
nand U23874 (N_23874,N_23453,N_23403);
and U23875 (N_23875,N_23396,N_23269);
nor U23876 (N_23876,N_23064,N_23063);
nand U23877 (N_23877,N_23317,N_23275);
and U23878 (N_23878,N_23111,N_23419);
xor U23879 (N_23879,N_23103,N_23145);
xor U23880 (N_23880,N_23072,N_23330);
or U23881 (N_23881,N_23210,N_23246);
nor U23882 (N_23882,N_23001,N_23188);
nand U23883 (N_23883,N_23169,N_23194);
xor U23884 (N_23884,N_23013,N_23368);
nor U23885 (N_23885,N_23451,N_23047);
and U23886 (N_23886,N_23438,N_23094);
nor U23887 (N_23887,N_23001,N_23226);
xnor U23888 (N_23888,N_23208,N_23494);
nand U23889 (N_23889,N_23219,N_23136);
xnor U23890 (N_23890,N_23093,N_23155);
nand U23891 (N_23891,N_23145,N_23266);
nand U23892 (N_23892,N_23342,N_23301);
xnor U23893 (N_23893,N_23457,N_23388);
and U23894 (N_23894,N_23403,N_23095);
nor U23895 (N_23895,N_23194,N_23358);
or U23896 (N_23896,N_23162,N_23265);
xnor U23897 (N_23897,N_23264,N_23217);
nor U23898 (N_23898,N_23000,N_23344);
nand U23899 (N_23899,N_23419,N_23279);
or U23900 (N_23900,N_23297,N_23322);
and U23901 (N_23901,N_23001,N_23435);
and U23902 (N_23902,N_23231,N_23229);
nor U23903 (N_23903,N_23352,N_23041);
nand U23904 (N_23904,N_23477,N_23253);
nand U23905 (N_23905,N_23357,N_23145);
or U23906 (N_23906,N_23112,N_23055);
nand U23907 (N_23907,N_23280,N_23362);
nor U23908 (N_23908,N_23292,N_23026);
xnor U23909 (N_23909,N_23036,N_23394);
and U23910 (N_23910,N_23411,N_23037);
or U23911 (N_23911,N_23026,N_23047);
nor U23912 (N_23912,N_23340,N_23324);
xor U23913 (N_23913,N_23023,N_23170);
nand U23914 (N_23914,N_23159,N_23156);
nand U23915 (N_23915,N_23312,N_23471);
nor U23916 (N_23916,N_23034,N_23196);
xor U23917 (N_23917,N_23095,N_23400);
or U23918 (N_23918,N_23381,N_23009);
and U23919 (N_23919,N_23454,N_23423);
or U23920 (N_23920,N_23125,N_23398);
and U23921 (N_23921,N_23258,N_23238);
xnor U23922 (N_23922,N_23341,N_23041);
nand U23923 (N_23923,N_23363,N_23475);
xnor U23924 (N_23924,N_23069,N_23325);
and U23925 (N_23925,N_23394,N_23447);
nor U23926 (N_23926,N_23071,N_23123);
xor U23927 (N_23927,N_23008,N_23314);
xnor U23928 (N_23928,N_23450,N_23385);
and U23929 (N_23929,N_23393,N_23319);
and U23930 (N_23930,N_23319,N_23021);
nand U23931 (N_23931,N_23419,N_23214);
xnor U23932 (N_23932,N_23373,N_23450);
and U23933 (N_23933,N_23085,N_23227);
or U23934 (N_23934,N_23174,N_23345);
nand U23935 (N_23935,N_23114,N_23137);
or U23936 (N_23936,N_23202,N_23121);
nand U23937 (N_23937,N_23173,N_23164);
or U23938 (N_23938,N_23475,N_23097);
xnor U23939 (N_23939,N_23402,N_23355);
and U23940 (N_23940,N_23258,N_23325);
and U23941 (N_23941,N_23118,N_23019);
xor U23942 (N_23942,N_23089,N_23035);
or U23943 (N_23943,N_23193,N_23443);
or U23944 (N_23944,N_23460,N_23412);
nor U23945 (N_23945,N_23257,N_23028);
and U23946 (N_23946,N_23370,N_23243);
and U23947 (N_23947,N_23247,N_23263);
or U23948 (N_23948,N_23374,N_23232);
or U23949 (N_23949,N_23349,N_23133);
nor U23950 (N_23950,N_23277,N_23449);
nand U23951 (N_23951,N_23483,N_23281);
and U23952 (N_23952,N_23255,N_23175);
nor U23953 (N_23953,N_23200,N_23185);
nand U23954 (N_23954,N_23219,N_23101);
nand U23955 (N_23955,N_23133,N_23070);
nand U23956 (N_23956,N_23039,N_23182);
nand U23957 (N_23957,N_23285,N_23313);
and U23958 (N_23958,N_23049,N_23262);
and U23959 (N_23959,N_23131,N_23053);
and U23960 (N_23960,N_23403,N_23299);
or U23961 (N_23961,N_23134,N_23088);
xnor U23962 (N_23962,N_23010,N_23324);
nand U23963 (N_23963,N_23142,N_23109);
nand U23964 (N_23964,N_23204,N_23259);
or U23965 (N_23965,N_23428,N_23229);
nand U23966 (N_23966,N_23280,N_23359);
nand U23967 (N_23967,N_23288,N_23482);
or U23968 (N_23968,N_23177,N_23096);
xor U23969 (N_23969,N_23411,N_23364);
and U23970 (N_23970,N_23460,N_23024);
nor U23971 (N_23971,N_23498,N_23391);
xnor U23972 (N_23972,N_23382,N_23044);
nor U23973 (N_23973,N_23222,N_23467);
nor U23974 (N_23974,N_23112,N_23222);
xor U23975 (N_23975,N_23109,N_23181);
or U23976 (N_23976,N_23253,N_23204);
nor U23977 (N_23977,N_23469,N_23086);
and U23978 (N_23978,N_23234,N_23492);
nor U23979 (N_23979,N_23133,N_23498);
nand U23980 (N_23980,N_23113,N_23432);
xnor U23981 (N_23981,N_23354,N_23064);
nor U23982 (N_23982,N_23377,N_23102);
nor U23983 (N_23983,N_23373,N_23058);
or U23984 (N_23984,N_23490,N_23179);
nand U23985 (N_23985,N_23174,N_23290);
nand U23986 (N_23986,N_23206,N_23043);
or U23987 (N_23987,N_23462,N_23146);
or U23988 (N_23988,N_23332,N_23234);
xnor U23989 (N_23989,N_23265,N_23432);
xnor U23990 (N_23990,N_23295,N_23383);
and U23991 (N_23991,N_23119,N_23055);
nor U23992 (N_23992,N_23489,N_23394);
xor U23993 (N_23993,N_23328,N_23000);
and U23994 (N_23994,N_23393,N_23311);
nand U23995 (N_23995,N_23455,N_23206);
nor U23996 (N_23996,N_23038,N_23355);
nor U23997 (N_23997,N_23094,N_23074);
xor U23998 (N_23998,N_23354,N_23347);
or U23999 (N_23999,N_23154,N_23246);
or U24000 (N_24000,N_23982,N_23593);
xnor U24001 (N_24001,N_23512,N_23776);
xnor U24002 (N_24002,N_23906,N_23703);
and U24003 (N_24003,N_23643,N_23855);
xor U24004 (N_24004,N_23939,N_23661);
nand U24005 (N_24005,N_23699,N_23790);
nor U24006 (N_24006,N_23969,N_23917);
and U24007 (N_24007,N_23730,N_23875);
nand U24008 (N_24008,N_23582,N_23524);
xor U24009 (N_24009,N_23992,N_23731);
and U24010 (N_24010,N_23907,N_23911);
and U24011 (N_24011,N_23801,N_23710);
xor U24012 (N_24012,N_23720,N_23686);
xnor U24013 (N_24013,N_23774,N_23778);
nor U24014 (N_24014,N_23599,N_23928);
or U24015 (N_24015,N_23962,N_23974);
and U24016 (N_24016,N_23777,N_23878);
nor U24017 (N_24017,N_23530,N_23850);
nand U24018 (N_24018,N_23747,N_23708);
nor U24019 (N_24019,N_23542,N_23967);
and U24020 (N_24020,N_23973,N_23722);
nor U24021 (N_24021,N_23990,N_23684);
nand U24022 (N_24022,N_23632,N_23539);
and U24023 (N_24023,N_23667,N_23834);
or U24024 (N_24024,N_23729,N_23680);
or U24025 (N_24025,N_23619,N_23757);
nand U24026 (N_24026,N_23791,N_23972);
nor U24027 (N_24027,N_23980,N_23944);
xor U24028 (N_24028,N_23798,N_23578);
nand U24029 (N_24029,N_23700,N_23821);
and U24030 (N_24030,N_23615,N_23891);
xnor U24031 (N_24031,N_23500,N_23690);
xnor U24032 (N_24032,N_23693,N_23601);
and U24033 (N_24033,N_23859,N_23544);
and U24034 (N_24034,N_23871,N_23828);
or U24035 (N_24035,N_23697,N_23943);
nand U24036 (N_24036,N_23689,N_23754);
or U24037 (N_24037,N_23677,N_23585);
xor U24038 (N_24038,N_23614,N_23823);
nand U24039 (N_24039,N_23957,N_23502);
nor U24040 (N_24040,N_23675,N_23549);
nand U24041 (N_24041,N_23711,N_23607);
or U24042 (N_24042,N_23641,N_23999);
nor U24043 (N_24043,N_23885,N_23877);
and U24044 (N_24044,N_23818,N_23958);
or U24045 (N_24045,N_23636,N_23597);
and U24046 (N_24046,N_23649,N_23545);
nand U24047 (N_24047,N_23803,N_23836);
nor U24048 (N_24048,N_23587,N_23576);
and U24049 (N_24049,N_23892,N_23648);
and U24050 (N_24050,N_23640,N_23922);
or U24051 (N_24051,N_23504,N_23868);
xor U24052 (N_24052,N_23620,N_23724);
xnor U24053 (N_24053,N_23751,N_23725);
xnor U24054 (N_24054,N_23808,N_23795);
or U24055 (N_24055,N_23880,N_23752);
nor U24056 (N_24056,N_23896,N_23901);
and U24057 (N_24057,N_23625,N_23514);
or U24058 (N_24058,N_23874,N_23904);
or U24059 (N_24059,N_23537,N_23920);
xor U24060 (N_24060,N_23695,N_23622);
nand U24061 (N_24061,N_23737,N_23705);
nor U24062 (N_24062,N_23735,N_23561);
xnor U24063 (N_24063,N_23520,N_23959);
nor U24064 (N_24064,N_23817,N_23704);
nor U24065 (N_24065,N_23580,N_23989);
xor U24066 (N_24066,N_23937,N_23764);
xnor U24067 (N_24067,N_23867,N_23598);
nor U24068 (N_24068,N_23851,N_23794);
nor U24069 (N_24069,N_23954,N_23914);
xor U24070 (N_24070,N_23952,N_23555);
nor U24071 (N_24071,N_23694,N_23845);
and U24072 (N_24072,N_23673,N_23941);
nand U24073 (N_24073,N_23556,N_23883);
and U24074 (N_24074,N_23560,N_23986);
nor U24075 (N_24075,N_23984,N_23709);
nand U24076 (N_24076,N_23988,N_23857);
nand U24077 (N_24077,N_23733,N_23740);
nand U24078 (N_24078,N_23863,N_23756);
xnor U24079 (N_24079,N_23628,N_23876);
or U24080 (N_24080,N_23548,N_23603);
nand U24081 (N_24081,N_23565,N_23832);
nor U24082 (N_24082,N_23951,N_23706);
xnor U24083 (N_24083,N_23559,N_23976);
or U24084 (N_24084,N_23780,N_23616);
nand U24085 (N_24085,N_23717,N_23698);
nand U24086 (N_24086,N_23932,N_23543);
nand U24087 (N_24087,N_23511,N_23748);
xnor U24088 (N_24088,N_23535,N_23668);
nand U24089 (N_24089,N_23602,N_23547);
nand U24090 (N_24090,N_23617,N_23910);
or U24091 (N_24091,N_23788,N_23792);
xor U24092 (N_24092,N_23749,N_23590);
and U24093 (N_24093,N_23770,N_23767);
and U24094 (N_24094,N_23899,N_23666);
nand U24095 (N_24095,N_23866,N_23925);
nor U24096 (N_24096,N_23806,N_23786);
nor U24097 (N_24097,N_23771,N_23738);
nor U24098 (N_24098,N_23660,N_23835);
or U24099 (N_24099,N_23965,N_23936);
nor U24100 (N_24100,N_23948,N_23807);
xor U24101 (N_24101,N_23827,N_23997);
nor U24102 (N_24102,N_23853,N_23696);
nand U24103 (N_24103,N_23926,N_23744);
or U24104 (N_24104,N_23996,N_23844);
nand U24105 (N_24105,N_23812,N_23831);
xor U24106 (N_24106,N_23721,N_23956);
xor U24107 (N_24107,N_23626,N_23682);
xor U24108 (N_24108,N_23970,N_23513);
nand U24109 (N_24109,N_23650,N_23782);
xor U24110 (N_24110,N_23657,N_23830);
xnor U24111 (N_24111,N_23769,N_23852);
and U24112 (N_24112,N_23995,N_23586);
nor U24113 (N_24113,N_23915,N_23654);
nand U24114 (N_24114,N_23631,N_23604);
nor U24115 (N_24115,N_23509,N_23858);
xor U24116 (N_24116,N_23663,N_23618);
nand U24117 (N_24117,N_23713,N_23589);
nor U24118 (N_24118,N_23946,N_23856);
xnor U24119 (N_24119,N_23676,N_23692);
nand U24120 (N_24120,N_23762,N_23532);
nand U24121 (N_24121,N_23758,N_23913);
nand U24122 (N_24122,N_23805,N_23505);
nor U24123 (N_24123,N_23779,N_23701);
nand U24124 (N_24124,N_23864,N_23596);
or U24125 (N_24125,N_23557,N_23687);
xor U24126 (N_24126,N_23799,N_23960);
or U24127 (N_24127,N_23865,N_23889);
or U24128 (N_24128,N_23563,N_23552);
or U24129 (N_24129,N_23612,N_23564);
nand U24130 (N_24130,N_23633,N_23723);
and U24131 (N_24131,N_23789,N_23678);
or U24132 (N_24132,N_23567,N_23683);
or U24133 (N_24133,N_23569,N_23536);
nor U24134 (N_24134,N_23670,N_23881);
xor U24135 (N_24135,N_23674,N_23726);
and U24136 (N_24136,N_23785,N_23662);
and U24137 (N_24137,N_23558,N_23966);
xor U24138 (N_24138,N_23783,N_23518);
or U24139 (N_24139,N_23506,N_23921);
nand U24140 (N_24140,N_23727,N_23934);
and U24141 (N_24141,N_23888,N_23655);
nand U24142 (N_24142,N_23659,N_23507);
nand U24143 (N_24143,N_23810,N_23861);
nor U24144 (N_24144,N_23645,N_23908);
and U24145 (N_24145,N_23642,N_23873);
and U24146 (N_24146,N_23572,N_23734);
nor U24147 (N_24147,N_23950,N_23826);
nand U24148 (N_24148,N_23897,N_23784);
xnor U24149 (N_24149,N_23947,N_23765);
or U24150 (N_24150,N_23577,N_23975);
xor U24151 (N_24151,N_23775,N_23630);
and U24152 (N_24152,N_23594,N_23571);
xor U24153 (N_24153,N_23574,N_23613);
nand U24154 (N_24154,N_23581,N_23849);
nor U24155 (N_24155,N_23610,N_23608);
nor U24156 (N_24156,N_23815,N_23820);
and U24157 (N_24157,N_23813,N_23681);
nor U24158 (N_24158,N_23998,N_23755);
and U24159 (N_24159,N_23522,N_23651);
nand U24160 (N_24160,N_23766,N_23869);
and U24161 (N_24161,N_23846,N_23517);
nand U24162 (N_24162,N_23860,N_23551);
xor U24163 (N_24163,N_23847,N_23665);
xnor U24164 (N_24164,N_23637,N_23554);
or U24165 (N_24165,N_23890,N_23924);
and U24166 (N_24166,N_23819,N_23745);
nor U24167 (N_24167,N_23624,N_23742);
or U24168 (N_24168,N_23743,N_23994);
or U24169 (N_24169,N_23584,N_23829);
or U24170 (N_24170,N_23900,N_23718);
and U24171 (N_24171,N_23629,N_23912);
nand U24172 (N_24172,N_23987,N_23719);
and U24173 (N_24173,N_23595,N_23716);
or U24174 (N_24174,N_23712,N_23971);
or U24175 (N_24175,N_23949,N_23644);
nand U24176 (N_24176,N_23882,N_23872);
nand U24177 (N_24177,N_23903,N_23942);
or U24178 (N_24178,N_23728,N_23905);
xnor U24179 (N_24179,N_23526,N_23739);
xnor U24180 (N_24180,N_23916,N_23592);
xor U24181 (N_24181,N_23679,N_23991);
and U24182 (N_24182,N_23553,N_23816);
xnor U24183 (N_24183,N_23508,N_23627);
xor U24184 (N_24184,N_23879,N_23886);
or U24185 (N_24185,N_23575,N_23541);
or U24186 (N_24186,N_23732,N_23750);
nor U24187 (N_24187,N_23570,N_23741);
and U24188 (N_24188,N_23707,N_23521);
and U24189 (N_24189,N_23893,N_23528);
xor U24190 (N_24190,N_23773,N_23605);
xor U24191 (N_24191,N_23837,N_23533);
and U24192 (N_24192,N_23688,N_23927);
and U24193 (N_24193,N_23895,N_23652);
nor U24194 (N_24194,N_23919,N_23977);
nor U24195 (N_24195,N_23804,N_23656);
or U24196 (N_24196,N_23838,N_23550);
nor U24197 (N_24197,N_23525,N_23887);
nor U24198 (N_24198,N_23638,N_23979);
nand U24199 (N_24199,N_23515,N_23968);
or U24200 (N_24200,N_23940,N_23894);
nand U24201 (N_24201,N_23796,N_23978);
nor U24202 (N_24202,N_23923,N_23839);
and U24203 (N_24203,N_23546,N_23902);
nor U24204 (N_24204,N_23993,N_23811);
nand U24205 (N_24205,N_23573,N_23843);
nor U24206 (N_24206,N_23898,N_23983);
xor U24207 (N_24207,N_23753,N_23583);
xnor U24208 (N_24208,N_23702,N_23600);
and U24209 (N_24209,N_23963,N_23929);
nor U24210 (N_24210,N_23822,N_23964);
or U24211 (N_24211,N_23534,N_23621);
xor U24212 (N_24212,N_23579,N_23930);
xnor U24213 (N_24213,N_23588,N_23763);
xor U24214 (N_24214,N_23529,N_23945);
or U24215 (N_24215,N_23800,N_23523);
xnor U24216 (N_24216,N_23519,N_23814);
and U24217 (N_24217,N_23772,N_23761);
xor U24218 (N_24218,N_23609,N_23635);
nand U24219 (N_24219,N_23797,N_23759);
xnor U24220 (N_24220,N_23848,N_23691);
nor U24221 (N_24221,N_23562,N_23664);
xnor U24222 (N_24222,N_23736,N_23931);
nor U24223 (N_24223,N_23685,N_23503);
nor U24224 (N_24224,N_23606,N_23909);
or U24225 (N_24225,N_23809,N_23714);
or U24226 (N_24226,N_23842,N_23933);
xnor U24227 (N_24227,N_23802,N_23623);
nand U24228 (N_24228,N_23672,N_23611);
xnor U24229 (N_24229,N_23824,N_23981);
nor U24230 (N_24230,N_23985,N_23639);
and U24231 (N_24231,N_23501,N_23793);
nand U24232 (N_24232,N_23787,N_23653);
nor U24233 (N_24233,N_23955,N_23669);
or U24234 (N_24234,N_23540,N_23531);
xnor U24235 (N_24235,N_23961,N_23870);
and U24236 (N_24236,N_23768,N_23833);
and U24237 (N_24237,N_23516,N_23634);
nand U24238 (N_24238,N_23760,N_23862);
and U24239 (N_24239,N_23746,N_23854);
xnor U24240 (N_24240,N_23781,N_23918);
nor U24241 (N_24241,N_23566,N_23510);
nand U24242 (N_24242,N_23591,N_23884);
xor U24243 (N_24243,N_23647,N_23840);
nor U24244 (N_24244,N_23646,N_23538);
xor U24245 (N_24245,N_23953,N_23715);
xnor U24246 (N_24246,N_23671,N_23568);
xnor U24247 (N_24247,N_23825,N_23658);
nor U24248 (N_24248,N_23527,N_23841);
nand U24249 (N_24249,N_23938,N_23935);
and U24250 (N_24250,N_23943,N_23992);
nor U24251 (N_24251,N_23527,N_23626);
xor U24252 (N_24252,N_23841,N_23953);
nor U24253 (N_24253,N_23935,N_23660);
nor U24254 (N_24254,N_23771,N_23691);
or U24255 (N_24255,N_23612,N_23592);
xor U24256 (N_24256,N_23624,N_23759);
xor U24257 (N_24257,N_23954,N_23952);
and U24258 (N_24258,N_23846,N_23926);
nand U24259 (N_24259,N_23605,N_23982);
nand U24260 (N_24260,N_23771,N_23608);
nor U24261 (N_24261,N_23849,N_23986);
or U24262 (N_24262,N_23619,N_23523);
nor U24263 (N_24263,N_23747,N_23549);
and U24264 (N_24264,N_23601,N_23695);
or U24265 (N_24265,N_23626,N_23756);
xor U24266 (N_24266,N_23576,N_23828);
or U24267 (N_24267,N_23744,N_23526);
xnor U24268 (N_24268,N_23862,N_23947);
or U24269 (N_24269,N_23505,N_23948);
xnor U24270 (N_24270,N_23640,N_23758);
nand U24271 (N_24271,N_23842,N_23970);
or U24272 (N_24272,N_23809,N_23557);
xnor U24273 (N_24273,N_23729,N_23956);
nor U24274 (N_24274,N_23731,N_23759);
xnor U24275 (N_24275,N_23793,N_23987);
nor U24276 (N_24276,N_23746,N_23918);
nor U24277 (N_24277,N_23949,N_23888);
nand U24278 (N_24278,N_23903,N_23827);
or U24279 (N_24279,N_23664,N_23704);
or U24280 (N_24280,N_23724,N_23804);
or U24281 (N_24281,N_23665,N_23840);
nor U24282 (N_24282,N_23574,N_23804);
nor U24283 (N_24283,N_23854,N_23865);
nand U24284 (N_24284,N_23738,N_23974);
nand U24285 (N_24285,N_23762,N_23830);
nor U24286 (N_24286,N_23552,N_23650);
and U24287 (N_24287,N_23538,N_23709);
or U24288 (N_24288,N_23699,N_23748);
nor U24289 (N_24289,N_23565,N_23828);
or U24290 (N_24290,N_23878,N_23991);
or U24291 (N_24291,N_23910,N_23892);
nand U24292 (N_24292,N_23894,N_23561);
xor U24293 (N_24293,N_23507,N_23946);
xor U24294 (N_24294,N_23572,N_23725);
or U24295 (N_24295,N_23670,N_23785);
nand U24296 (N_24296,N_23545,N_23740);
or U24297 (N_24297,N_23522,N_23731);
nor U24298 (N_24298,N_23772,N_23621);
nor U24299 (N_24299,N_23764,N_23649);
nand U24300 (N_24300,N_23911,N_23948);
nor U24301 (N_24301,N_23677,N_23847);
nand U24302 (N_24302,N_23771,N_23636);
nor U24303 (N_24303,N_23920,N_23999);
nand U24304 (N_24304,N_23756,N_23711);
or U24305 (N_24305,N_23965,N_23963);
nand U24306 (N_24306,N_23817,N_23867);
or U24307 (N_24307,N_23870,N_23737);
and U24308 (N_24308,N_23595,N_23718);
nor U24309 (N_24309,N_23761,N_23815);
or U24310 (N_24310,N_23629,N_23813);
and U24311 (N_24311,N_23825,N_23596);
nand U24312 (N_24312,N_23879,N_23779);
nor U24313 (N_24313,N_23802,N_23811);
and U24314 (N_24314,N_23950,N_23629);
and U24315 (N_24315,N_23661,N_23772);
nor U24316 (N_24316,N_23849,N_23743);
nor U24317 (N_24317,N_23592,N_23548);
nand U24318 (N_24318,N_23827,N_23593);
and U24319 (N_24319,N_23909,N_23553);
nor U24320 (N_24320,N_23505,N_23707);
nor U24321 (N_24321,N_23553,N_23536);
or U24322 (N_24322,N_23808,N_23618);
nand U24323 (N_24323,N_23970,N_23839);
xor U24324 (N_24324,N_23547,N_23561);
and U24325 (N_24325,N_23644,N_23980);
and U24326 (N_24326,N_23808,N_23723);
or U24327 (N_24327,N_23942,N_23863);
nor U24328 (N_24328,N_23697,N_23758);
or U24329 (N_24329,N_23945,N_23619);
xor U24330 (N_24330,N_23820,N_23854);
xor U24331 (N_24331,N_23887,N_23775);
and U24332 (N_24332,N_23562,N_23558);
xor U24333 (N_24333,N_23609,N_23893);
or U24334 (N_24334,N_23968,N_23956);
xnor U24335 (N_24335,N_23679,N_23777);
nor U24336 (N_24336,N_23889,N_23991);
xnor U24337 (N_24337,N_23651,N_23813);
and U24338 (N_24338,N_23562,N_23809);
nand U24339 (N_24339,N_23832,N_23944);
and U24340 (N_24340,N_23899,N_23878);
nor U24341 (N_24341,N_23981,N_23980);
xnor U24342 (N_24342,N_23995,N_23985);
nor U24343 (N_24343,N_23602,N_23568);
nand U24344 (N_24344,N_23544,N_23712);
and U24345 (N_24345,N_23671,N_23904);
xnor U24346 (N_24346,N_23805,N_23647);
and U24347 (N_24347,N_23953,N_23606);
xnor U24348 (N_24348,N_23873,N_23766);
or U24349 (N_24349,N_23608,N_23605);
nor U24350 (N_24350,N_23737,N_23848);
nor U24351 (N_24351,N_23512,N_23619);
and U24352 (N_24352,N_23564,N_23776);
nor U24353 (N_24353,N_23641,N_23904);
nor U24354 (N_24354,N_23909,N_23802);
or U24355 (N_24355,N_23639,N_23931);
and U24356 (N_24356,N_23890,N_23560);
nand U24357 (N_24357,N_23869,N_23666);
nor U24358 (N_24358,N_23932,N_23770);
xor U24359 (N_24359,N_23668,N_23989);
and U24360 (N_24360,N_23546,N_23872);
nor U24361 (N_24361,N_23570,N_23806);
nor U24362 (N_24362,N_23747,N_23556);
xor U24363 (N_24363,N_23879,N_23620);
nand U24364 (N_24364,N_23543,N_23884);
nor U24365 (N_24365,N_23889,N_23505);
or U24366 (N_24366,N_23655,N_23759);
nor U24367 (N_24367,N_23885,N_23655);
and U24368 (N_24368,N_23586,N_23923);
and U24369 (N_24369,N_23580,N_23634);
or U24370 (N_24370,N_23661,N_23762);
and U24371 (N_24371,N_23500,N_23814);
and U24372 (N_24372,N_23937,N_23968);
nor U24373 (N_24373,N_23667,N_23767);
nor U24374 (N_24374,N_23508,N_23637);
and U24375 (N_24375,N_23656,N_23980);
or U24376 (N_24376,N_23526,N_23960);
xor U24377 (N_24377,N_23954,N_23958);
nor U24378 (N_24378,N_23605,N_23940);
nor U24379 (N_24379,N_23793,N_23954);
nor U24380 (N_24380,N_23573,N_23665);
xnor U24381 (N_24381,N_23743,N_23538);
and U24382 (N_24382,N_23544,N_23531);
nor U24383 (N_24383,N_23983,N_23834);
or U24384 (N_24384,N_23839,N_23925);
and U24385 (N_24385,N_23716,N_23696);
or U24386 (N_24386,N_23674,N_23893);
xnor U24387 (N_24387,N_23522,N_23818);
and U24388 (N_24388,N_23923,N_23696);
and U24389 (N_24389,N_23581,N_23547);
and U24390 (N_24390,N_23507,N_23738);
nand U24391 (N_24391,N_23601,N_23707);
nor U24392 (N_24392,N_23567,N_23596);
and U24393 (N_24393,N_23941,N_23899);
nor U24394 (N_24394,N_23605,N_23775);
nand U24395 (N_24395,N_23609,N_23810);
xnor U24396 (N_24396,N_23586,N_23623);
or U24397 (N_24397,N_23649,N_23915);
nor U24398 (N_24398,N_23777,N_23971);
and U24399 (N_24399,N_23542,N_23984);
nand U24400 (N_24400,N_23830,N_23995);
xnor U24401 (N_24401,N_23750,N_23705);
nand U24402 (N_24402,N_23922,N_23777);
xor U24403 (N_24403,N_23611,N_23816);
and U24404 (N_24404,N_23955,N_23655);
xnor U24405 (N_24405,N_23872,N_23549);
and U24406 (N_24406,N_23602,N_23988);
or U24407 (N_24407,N_23860,N_23517);
and U24408 (N_24408,N_23957,N_23688);
or U24409 (N_24409,N_23528,N_23918);
nor U24410 (N_24410,N_23800,N_23716);
nand U24411 (N_24411,N_23943,N_23668);
and U24412 (N_24412,N_23787,N_23517);
nand U24413 (N_24413,N_23739,N_23709);
nand U24414 (N_24414,N_23762,N_23925);
and U24415 (N_24415,N_23545,N_23546);
xnor U24416 (N_24416,N_23998,N_23896);
and U24417 (N_24417,N_23898,N_23793);
and U24418 (N_24418,N_23839,N_23852);
or U24419 (N_24419,N_23647,N_23733);
nand U24420 (N_24420,N_23812,N_23967);
or U24421 (N_24421,N_23718,N_23622);
nor U24422 (N_24422,N_23567,N_23765);
nand U24423 (N_24423,N_23789,N_23973);
nor U24424 (N_24424,N_23940,N_23885);
nand U24425 (N_24425,N_23783,N_23872);
xnor U24426 (N_24426,N_23774,N_23857);
and U24427 (N_24427,N_23992,N_23935);
nand U24428 (N_24428,N_23808,N_23502);
and U24429 (N_24429,N_23782,N_23818);
nor U24430 (N_24430,N_23623,N_23524);
xnor U24431 (N_24431,N_23518,N_23553);
or U24432 (N_24432,N_23963,N_23737);
xor U24433 (N_24433,N_23516,N_23950);
and U24434 (N_24434,N_23903,N_23549);
xor U24435 (N_24435,N_23701,N_23869);
nor U24436 (N_24436,N_23532,N_23821);
nand U24437 (N_24437,N_23623,N_23652);
and U24438 (N_24438,N_23896,N_23914);
and U24439 (N_24439,N_23538,N_23944);
xor U24440 (N_24440,N_23654,N_23696);
xnor U24441 (N_24441,N_23829,N_23695);
or U24442 (N_24442,N_23821,N_23902);
nor U24443 (N_24443,N_23597,N_23970);
and U24444 (N_24444,N_23775,N_23729);
nand U24445 (N_24445,N_23901,N_23779);
or U24446 (N_24446,N_23908,N_23854);
or U24447 (N_24447,N_23638,N_23550);
nand U24448 (N_24448,N_23552,N_23816);
nand U24449 (N_24449,N_23725,N_23857);
nor U24450 (N_24450,N_23518,N_23652);
nand U24451 (N_24451,N_23834,N_23805);
xor U24452 (N_24452,N_23862,N_23945);
and U24453 (N_24453,N_23797,N_23765);
xor U24454 (N_24454,N_23611,N_23830);
xor U24455 (N_24455,N_23575,N_23905);
xor U24456 (N_24456,N_23664,N_23918);
or U24457 (N_24457,N_23694,N_23626);
nor U24458 (N_24458,N_23991,N_23854);
or U24459 (N_24459,N_23611,N_23551);
and U24460 (N_24460,N_23938,N_23798);
xor U24461 (N_24461,N_23623,N_23873);
nand U24462 (N_24462,N_23818,N_23545);
xor U24463 (N_24463,N_23833,N_23615);
and U24464 (N_24464,N_23646,N_23667);
or U24465 (N_24465,N_23718,N_23767);
nand U24466 (N_24466,N_23658,N_23889);
or U24467 (N_24467,N_23624,N_23888);
nand U24468 (N_24468,N_23526,N_23946);
xnor U24469 (N_24469,N_23772,N_23693);
xnor U24470 (N_24470,N_23743,N_23662);
or U24471 (N_24471,N_23622,N_23726);
nor U24472 (N_24472,N_23547,N_23536);
nand U24473 (N_24473,N_23985,N_23843);
xor U24474 (N_24474,N_23785,N_23860);
or U24475 (N_24475,N_23975,N_23995);
nand U24476 (N_24476,N_23834,N_23769);
or U24477 (N_24477,N_23828,N_23503);
or U24478 (N_24478,N_23570,N_23980);
or U24479 (N_24479,N_23750,N_23939);
nor U24480 (N_24480,N_23600,N_23809);
xnor U24481 (N_24481,N_23831,N_23745);
and U24482 (N_24482,N_23518,N_23965);
nand U24483 (N_24483,N_23800,N_23612);
and U24484 (N_24484,N_23518,N_23511);
nand U24485 (N_24485,N_23995,N_23799);
nand U24486 (N_24486,N_23606,N_23727);
and U24487 (N_24487,N_23640,N_23590);
xor U24488 (N_24488,N_23525,N_23567);
xnor U24489 (N_24489,N_23539,N_23535);
nor U24490 (N_24490,N_23781,N_23819);
and U24491 (N_24491,N_23880,N_23808);
nor U24492 (N_24492,N_23719,N_23686);
nand U24493 (N_24493,N_23675,N_23606);
and U24494 (N_24494,N_23515,N_23779);
xnor U24495 (N_24495,N_23672,N_23640);
and U24496 (N_24496,N_23582,N_23748);
xor U24497 (N_24497,N_23529,N_23944);
and U24498 (N_24498,N_23876,N_23974);
and U24499 (N_24499,N_23654,N_23746);
or U24500 (N_24500,N_24275,N_24000);
xnor U24501 (N_24501,N_24208,N_24036);
nand U24502 (N_24502,N_24379,N_24322);
and U24503 (N_24503,N_24062,N_24189);
or U24504 (N_24504,N_24236,N_24212);
nand U24505 (N_24505,N_24076,N_24056);
and U24506 (N_24506,N_24040,N_24021);
xor U24507 (N_24507,N_24432,N_24271);
or U24508 (N_24508,N_24319,N_24240);
xor U24509 (N_24509,N_24103,N_24371);
xor U24510 (N_24510,N_24199,N_24229);
nor U24511 (N_24511,N_24362,N_24377);
nor U24512 (N_24512,N_24116,N_24260);
nand U24513 (N_24513,N_24344,N_24442);
nor U24514 (N_24514,N_24012,N_24176);
nand U24515 (N_24515,N_24304,N_24462);
or U24516 (N_24516,N_24065,N_24293);
nand U24517 (N_24517,N_24493,N_24218);
xor U24518 (N_24518,N_24487,N_24484);
nand U24519 (N_24519,N_24324,N_24339);
nor U24520 (N_24520,N_24064,N_24035);
and U24521 (N_24521,N_24367,N_24125);
nor U24522 (N_24522,N_24210,N_24426);
or U24523 (N_24523,N_24029,N_24238);
xor U24524 (N_24524,N_24084,N_24004);
xnor U24525 (N_24525,N_24131,N_24245);
nor U24526 (N_24526,N_24494,N_24204);
xor U24527 (N_24527,N_24030,N_24312);
or U24528 (N_24528,N_24300,N_24305);
and U24529 (N_24529,N_24412,N_24042);
xnor U24530 (N_24530,N_24227,N_24273);
xor U24531 (N_24531,N_24150,N_24429);
or U24532 (N_24532,N_24460,N_24058);
nand U24533 (N_24533,N_24311,N_24485);
nand U24534 (N_24534,N_24378,N_24153);
nand U24535 (N_24535,N_24255,N_24482);
xnor U24536 (N_24536,N_24451,N_24157);
or U24537 (N_24537,N_24336,N_24111);
nand U24538 (N_24538,N_24025,N_24100);
xnor U24539 (N_24539,N_24235,N_24452);
and U24540 (N_24540,N_24207,N_24028);
or U24541 (N_24541,N_24106,N_24239);
xnor U24542 (N_24542,N_24201,N_24225);
nor U24543 (N_24543,N_24213,N_24327);
and U24544 (N_24544,N_24047,N_24481);
and U24545 (N_24545,N_24135,N_24385);
nand U24546 (N_24546,N_24140,N_24003);
nor U24547 (N_24547,N_24123,N_24474);
nor U24548 (N_24548,N_24489,N_24326);
or U24549 (N_24549,N_24441,N_24161);
xor U24550 (N_24550,N_24110,N_24053);
or U24551 (N_24551,N_24285,N_24133);
nand U24552 (N_24552,N_24470,N_24366);
nand U24553 (N_24553,N_24302,N_24043);
xor U24554 (N_24554,N_24099,N_24018);
and U24555 (N_24555,N_24461,N_24050);
or U24556 (N_24556,N_24403,N_24347);
and U24557 (N_24557,N_24093,N_24194);
nor U24558 (N_24558,N_24145,N_24231);
or U24559 (N_24559,N_24364,N_24016);
nand U24560 (N_24560,N_24413,N_24148);
nor U24561 (N_24561,N_24097,N_24181);
xnor U24562 (N_24562,N_24015,N_24120);
or U24563 (N_24563,N_24078,N_24288);
nor U24564 (N_24564,N_24262,N_24320);
and U24565 (N_24565,N_24142,N_24007);
xnor U24566 (N_24566,N_24284,N_24417);
nand U24567 (N_24567,N_24323,N_24476);
nor U24568 (N_24568,N_24349,N_24276);
nor U24569 (N_24569,N_24159,N_24292);
xor U24570 (N_24570,N_24248,N_24444);
and U24571 (N_24571,N_24196,N_24317);
nor U24572 (N_24572,N_24496,N_24002);
and U24573 (N_24573,N_24400,N_24269);
nand U24574 (N_24574,N_24373,N_24254);
nor U24575 (N_24575,N_24290,N_24465);
nor U24576 (N_24576,N_24039,N_24114);
nor U24577 (N_24577,N_24399,N_24149);
nand U24578 (N_24578,N_24202,N_24329);
xnor U24579 (N_24579,N_24232,N_24085);
xnor U24580 (N_24580,N_24249,N_24282);
and U24581 (N_24581,N_24203,N_24309);
or U24582 (N_24582,N_24080,N_24321);
nand U24583 (N_24583,N_24431,N_24361);
nand U24584 (N_24584,N_24092,N_24328);
xnor U24585 (N_24585,N_24343,N_24448);
or U24586 (N_24586,N_24155,N_24310);
xor U24587 (N_24587,N_24277,N_24386);
and U24588 (N_24588,N_24384,N_24340);
xor U24589 (N_24589,N_24104,N_24486);
nor U24590 (N_24590,N_24251,N_24172);
and U24591 (N_24591,N_24105,N_24478);
xor U24592 (N_24592,N_24077,N_24205);
nor U24593 (N_24593,N_24393,N_24224);
or U24594 (N_24594,N_24352,N_24475);
nor U24595 (N_24595,N_24453,N_24391);
or U24596 (N_24596,N_24160,N_24253);
and U24597 (N_24597,N_24087,N_24169);
xnor U24598 (N_24598,N_24139,N_24298);
and U24599 (N_24599,N_24415,N_24073);
xor U24600 (N_24600,N_24468,N_24112);
xnor U24601 (N_24601,N_24369,N_24198);
nand U24602 (N_24602,N_24286,N_24197);
nand U24603 (N_24603,N_24033,N_24355);
and U24604 (N_24604,N_24049,N_24045);
or U24605 (N_24605,N_24348,N_24443);
nand U24606 (N_24606,N_24283,N_24353);
nor U24607 (N_24607,N_24418,N_24265);
and U24608 (N_24608,N_24409,N_24346);
nor U24609 (N_24609,N_24458,N_24422);
nand U24610 (N_24610,N_24261,N_24214);
nand U24611 (N_24611,N_24301,N_24094);
xor U24612 (N_24612,N_24318,N_24368);
nor U24613 (N_24613,N_24044,N_24427);
nor U24614 (N_24614,N_24250,N_24419);
xnor U24615 (N_24615,N_24308,N_24438);
xor U24616 (N_24616,N_24022,N_24136);
nor U24617 (N_24617,N_24332,N_24156);
and U24618 (N_24618,N_24166,N_24287);
xor U24619 (N_24619,N_24168,N_24178);
and U24620 (N_24620,N_24020,N_24134);
nor U24621 (N_24621,N_24257,N_24471);
nand U24622 (N_24622,N_24380,N_24041);
nand U24623 (N_24623,N_24370,N_24387);
nand U24624 (N_24624,N_24101,N_24278);
xor U24625 (N_24625,N_24061,N_24375);
and U24626 (N_24626,N_24054,N_24372);
and U24627 (N_24627,N_24404,N_24463);
and U24628 (N_24628,N_24147,N_24469);
and U24629 (N_24629,N_24401,N_24006);
xor U24630 (N_24630,N_24488,N_24128);
xor U24631 (N_24631,N_24389,N_24209);
or U24632 (N_24632,N_24289,N_24244);
and U24633 (N_24633,N_24267,N_24024);
and U24634 (N_24634,N_24032,N_24026);
nor U24635 (N_24635,N_24407,N_24472);
and U24636 (N_24636,N_24437,N_24118);
or U24637 (N_24637,N_24129,N_24408);
or U24638 (N_24638,N_24424,N_24206);
xor U24639 (N_24639,N_24005,N_24423);
xnor U24640 (N_24640,N_24001,N_24241);
nand U24641 (N_24641,N_24009,N_24215);
nand U24642 (N_24642,N_24190,N_24013);
xnor U24643 (N_24643,N_24060,N_24174);
or U24644 (N_24644,N_24428,N_24495);
and U24645 (N_24645,N_24138,N_24052);
or U24646 (N_24646,N_24182,N_24263);
nor U24647 (N_24647,N_24046,N_24011);
and U24648 (N_24648,N_24497,N_24363);
nor U24649 (N_24649,N_24337,N_24086);
nor U24650 (N_24650,N_24242,N_24115);
xnor U24651 (N_24651,N_24274,N_24295);
and U24652 (N_24652,N_24102,N_24083);
and U24653 (N_24653,N_24457,N_24158);
nand U24654 (N_24654,N_24167,N_24165);
or U24655 (N_24655,N_24081,N_24068);
or U24656 (N_24656,N_24019,N_24233);
nor U24657 (N_24657,N_24491,N_24072);
and U24658 (N_24658,N_24330,N_24358);
or U24659 (N_24659,N_24063,N_24070);
and U24660 (N_24660,N_24108,N_24057);
nand U24661 (N_24661,N_24243,N_24055);
and U24662 (N_24662,N_24187,N_24141);
and U24663 (N_24663,N_24354,N_24272);
nand U24664 (N_24664,N_24416,N_24221);
nand U24665 (N_24665,N_24027,N_24307);
or U24666 (N_24666,N_24395,N_24430);
nor U24667 (N_24667,N_24294,N_24455);
nor U24668 (N_24668,N_24193,N_24096);
and U24669 (N_24669,N_24188,N_24479);
or U24670 (N_24670,N_24192,N_24306);
nand U24671 (N_24671,N_24048,N_24051);
nor U24672 (N_24672,N_24171,N_24477);
nand U24673 (N_24673,N_24303,N_24331);
xor U24674 (N_24674,N_24420,N_24398);
or U24675 (N_24675,N_24126,N_24091);
or U24676 (N_24676,N_24466,N_24392);
nand U24677 (N_24677,N_24490,N_24154);
nand U24678 (N_24678,N_24071,N_24335);
or U24679 (N_24679,N_24338,N_24410);
xor U24680 (N_24680,N_24449,N_24281);
xor U24681 (N_24681,N_24264,N_24492);
or U24682 (N_24682,N_24359,N_24183);
nor U24683 (N_24683,N_24217,N_24360);
nand U24684 (N_24684,N_24402,N_24414);
nand U24685 (N_24685,N_24334,N_24010);
xor U24686 (N_24686,N_24195,N_24216);
nand U24687 (N_24687,N_24237,N_24014);
nor U24688 (N_24688,N_24185,N_24177);
xnor U24689 (N_24689,N_24483,N_24146);
xnor U24690 (N_24690,N_24023,N_24314);
or U24691 (N_24691,N_24256,N_24383);
and U24692 (N_24692,N_24357,N_24088);
or U24693 (N_24693,N_24067,N_24456);
or U24694 (N_24694,N_24162,N_24152);
nor U24695 (N_24695,N_24333,N_24222);
or U24696 (N_24696,N_24299,N_24075);
nand U24697 (N_24697,N_24396,N_24137);
nand U24698 (N_24698,N_24069,N_24315);
and U24699 (N_24699,N_24200,N_24350);
or U24700 (N_24700,N_24252,N_24220);
nand U24701 (N_24701,N_24388,N_24079);
xor U24702 (N_24702,N_24436,N_24464);
xor U24703 (N_24703,N_24226,N_24342);
xnor U24704 (N_24704,N_24127,N_24280);
nand U24705 (N_24705,N_24098,N_24341);
nor U24706 (N_24706,N_24117,N_24297);
and U24707 (N_24707,N_24163,N_24119);
or U24708 (N_24708,N_24038,N_24439);
nand U24709 (N_24709,N_24121,N_24059);
and U24710 (N_24710,N_24107,N_24445);
nor U24711 (N_24711,N_24143,N_24008);
xnor U24712 (N_24712,N_24089,N_24180);
or U24713 (N_24713,N_24406,N_24175);
or U24714 (N_24714,N_24219,N_24405);
nand U24715 (N_24715,N_24130,N_24473);
nor U24716 (N_24716,N_24132,N_24382);
xor U24717 (N_24717,N_24296,N_24109);
nand U24718 (N_24718,N_24031,N_24365);
or U24719 (N_24719,N_24316,N_24228);
xor U24720 (N_24720,N_24440,N_24268);
nor U24721 (N_24721,N_24186,N_24381);
xor U24722 (N_24722,N_24173,N_24184);
or U24723 (N_24723,N_24390,N_24313);
xnor U24724 (N_24724,N_24179,N_24113);
or U24725 (N_24725,N_24234,N_24291);
nor U24726 (N_24726,N_24425,N_24266);
xnor U24727 (N_24727,N_24223,N_24394);
xor U24728 (N_24728,N_24279,N_24258);
xnor U24729 (N_24729,N_24450,N_24480);
nand U24730 (N_24730,N_24246,N_24435);
and U24731 (N_24731,N_24230,N_24374);
nor U24732 (N_24732,N_24211,N_24434);
and U24733 (N_24733,N_24164,N_24325);
and U24734 (N_24734,N_24170,N_24454);
nor U24735 (N_24735,N_24090,N_24259);
xnor U24736 (N_24736,N_24270,N_24247);
and U24737 (N_24737,N_24191,N_24037);
and U24738 (N_24738,N_24151,N_24459);
or U24739 (N_24739,N_24345,N_24467);
or U24740 (N_24740,N_24074,N_24144);
nand U24741 (N_24741,N_24122,N_24066);
and U24742 (N_24742,N_24411,N_24421);
and U24743 (N_24743,N_24433,N_24447);
xor U24744 (N_24744,N_24124,N_24034);
nand U24745 (N_24745,N_24397,N_24095);
xor U24746 (N_24746,N_24356,N_24376);
nor U24747 (N_24747,N_24082,N_24351);
nand U24748 (N_24748,N_24017,N_24446);
nand U24749 (N_24749,N_24499,N_24498);
xnor U24750 (N_24750,N_24477,N_24084);
or U24751 (N_24751,N_24040,N_24195);
or U24752 (N_24752,N_24371,N_24204);
xnor U24753 (N_24753,N_24370,N_24298);
xor U24754 (N_24754,N_24140,N_24271);
nor U24755 (N_24755,N_24384,N_24180);
or U24756 (N_24756,N_24119,N_24258);
nor U24757 (N_24757,N_24165,N_24295);
nand U24758 (N_24758,N_24235,N_24252);
nor U24759 (N_24759,N_24443,N_24420);
nand U24760 (N_24760,N_24034,N_24055);
nand U24761 (N_24761,N_24159,N_24498);
nor U24762 (N_24762,N_24186,N_24145);
or U24763 (N_24763,N_24077,N_24455);
nand U24764 (N_24764,N_24216,N_24175);
or U24765 (N_24765,N_24026,N_24237);
or U24766 (N_24766,N_24483,N_24273);
nand U24767 (N_24767,N_24092,N_24071);
and U24768 (N_24768,N_24293,N_24382);
nand U24769 (N_24769,N_24131,N_24063);
or U24770 (N_24770,N_24025,N_24252);
nor U24771 (N_24771,N_24344,N_24057);
nand U24772 (N_24772,N_24156,N_24106);
or U24773 (N_24773,N_24327,N_24385);
nor U24774 (N_24774,N_24449,N_24258);
and U24775 (N_24775,N_24138,N_24085);
nand U24776 (N_24776,N_24364,N_24362);
xnor U24777 (N_24777,N_24307,N_24430);
and U24778 (N_24778,N_24428,N_24340);
xor U24779 (N_24779,N_24078,N_24306);
and U24780 (N_24780,N_24303,N_24460);
and U24781 (N_24781,N_24462,N_24157);
and U24782 (N_24782,N_24141,N_24112);
nor U24783 (N_24783,N_24113,N_24456);
or U24784 (N_24784,N_24444,N_24389);
nor U24785 (N_24785,N_24419,N_24073);
or U24786 (N_24786,N_24384,N_24189);
or U24787 (N_24787,N_24011,N_24499);
nand U24788 (N_24788,N_24324,N_24005);
nand U24789 (N_24789,N_24135,N_24497);
and U24790 (N_24790,N_24046,N_24039);
xnor U24791 (N_24791,N_24492,N_24200);
and U24792 (N_24792,N_24309,N_24305);
xor U24793 (N_24793,N_24390,N_24112);
or U24794 (N_24794,N_24465,N_24041);
and U24795 (N_24795,N_24316,N_24137);
xnor U24796 (N_24796,N_24031,N_24125);
nand U24797 (N_24797,N_24270,N_24044);
xor U24798 (N_24798,N_24428,N_24004);
nand U24799 (N_24799,N_24081,N_24464);
xnor U24800 (N_24800,N_24061,N_24481);
nor U24801 (N_24801,N_24072,N_24068);
and U24802 (N_24802,N_24465,N_24456);
xor U24803 (N_24803,N_24465,N_24418);
or U24804 (N_24804,N_24085,N_24132);
and U24805 (N_24805,N_24423,N_24006);
nand U24806 (N_24806,N_24246,N_24306);
nor U24807 (N_24807,N_24454,N_24254);
xor U24808 (N_24808,N_24481,N_24287);
nand U24809 (N_24809,N_24342,N_24157);
xor U24810 (N_24810,N_24127,N_24162);
xnor U24811 (N_24811,N_24172,N_24480);
nand U24812 (N_24812,N_24432,N_24376);
or U24813 (N_24813,N_24123,N_24471);
xnor U24814 (N_24814,N_24075,N_24303);
nand U24815 (N_24815,N_24216,N_24344);
and U24816 (N_24816,N_24439,N_24002);
and U24817 (N_24817,N_24309,N_24114);
and U24818 (N_24818,N_24369,N_24301);
nand U24819 (N_24819,N_24284,N_24203);
and U24820 (N_24820,N_24206,N_24091);
or U24821 (N_24821,N_24168,N_24002);
nor U24822 (N_24822,N_24486,N_24373);
and U24823 (N_24823,N_24360,N_24253);
nor U24824 (N_24824,N_24198,N_24329);
nand U24825 (N_24825,N_24277,N_24353);
xor U24826 (N_24826,N_24277,N_24419);
nand U24827 (N_24827,N_24478,N_24073);
and U24828 (N_24828,N_24091,N_24067);
nand U24829 (N_24829,N_24304,N_24007);
xnor U24830 (N_24830,N_24007,N_24251);
or U24831 (N_24831,N_24053,N_24037);
or U24832 (N_24832,N_24008,N_24162);
nor U24833 (N_24833,N_24311,N_24382);
nor U24834 (N_24834,N_24261,N_24190);
or U24835 (N_24835,N_24385,N_24073);
nand U24836 (N_24836,N_24303,N_24232);
nor U24837 (N_24837,N_24239,N_24037);
nor U24838 (N_24838,N_24026,N_24364);
nor U24839 (N_24839,N_24068,N_24243);
and U24840 (N_24840,N_24289,N_24029);
nand U24841 (N_24841,N_24277,N_24178);
or U24842 (N_24842,N_24075,N_24016);
xnor U24843 (N_24843,N_24108,N_24081);
or U24844 (N_24844,N_24117,N_24486);
and U24845 (N_24845,N_24381,N_24044);
xnor U24846 (N_24846,N_24326,N_24223);
nand U24847 (N_24847,N_24146,N_24372);
xor U24848 (N_24848,N_24093,N_24373);
or U24849 (N_24849,N_24396,N_24013);
nor U24850 (N_24850,N_24349,N_24100);
or U24851 (N_24851,N_24458,N_24468);
xnor U24852 (N_24852,N_24136,N_24402);
or U24853 (N_24853,N_24431,N_24258);
xor U24854 (N_24854,N_24491,N_24031);
and U24855 (N_24855,N_24008,N_24130);
nand U24856 (N_24856,N_24491,N_24246);
and U24857 (N_24857,N_24464,N_24383);
xnor U24858 (N_24858,N_24292,N_24390);
nand U24859 (N_24859,N_24027,N_24254);
nor U24860 (N_24860,N_24266,N_24335);
and U24861 (N_24861,N_24325,N_24329);
nand U24862 (N_24862,N_24053,N_24315);
xnor U24863 (N_24863,N_24057,N_24310);
or U24864 (N_24864,N_24132,N_24181);
nand U24865 (N_24865,N_24080,N_24340);
nand U24866 (N_24866,N_24407,N_24161);
nand U24867 (N_24867,N_24155,N_24498);
nand U24868 (N_24868,N_24366,N_24410);
nor U24869 (N_24869,N_24057,N_24167);
or U24870 (N_24870,N_24098,N_24137);
nor U24871 (N_24871,N_24016,N_24121);
or U24872 (N_24872,N_24132,N_24274);
xnor U24873 (N_24873,N_24413,N_24337);
or U24874 (N_24874,N_24306,N_24310);
nand U24875 (N_24875,N_24341,N_24113);
nor U24876 (N_24876,N_24211,N_24251);
nand U24877 (N_24877,N_24365,N_24126);
xor U24878 (N_24878,N_24129,N_24273);
and U24879 (N_24879,N_24205,N_24351);
and U24880 (N_24880,N_24049,N_24221);
and U24881 (N_24881,N_24238,N_24042);
xor U24882 (N_24882,N_24153,N_24059);
and U24883 (N_24883,N_24260,N_24096);
and U24884 (N_24884,N_24346,N_24324);
xnor U24885 (N_24885,N_24379,N_24275);
nor U24886 (N_24886,N_24253,N_24281);
or U24887 (N_24887,N_24075,N_24373);
xnor U24888 (N_24888,N_24062,N_24228);
xor U24889 (N_24889,N_24069,N_24028);
nor U24890 (N_24890,N_24243,N_24417);
and U24891 (N_24891,N_24259,N_24004);
and U24892 (N_24892,N_24017,N_24250);
or U24893 (N_24893,N_24152,N_24445);
nand U24894 (N_24894,N_24175,N_24277);
or U24895 (N_24895,N_24184,N_24468);
or U24896 (N_24896,N_24227,N_24313);
nand U24897 (N_24897,N_24276,N_24478);
nand U24898 (N_24898,N_24376,N_24024);
xnor U24899 (N_24899,N_24415,N_24264);
and U24900 (N_24900,N_24264,N_24113);
and U24901 (N_24901,N_24136,N_24007);
nand U24902 (N_24902,N_24148,N_24108);
and U24903 (N_24903,N_24201,N_24118);
or U24904 (N_24904,N_24128,N_24419);
or U24905 (N_24905,N_24072,N_24085);
nor U24906 (N_24906,N_24067,N_24295);
nor U24907 (N_24907,N_24211,N_24316);
xnor U24908 (N_24908,N_24404,N_24173);
or U24909 (N_24909,N_24072,N_24437);
xor U24910 (N_24910,N_24382,N_24242);
nand U24911 (N_24911,N_24170,N_24191);
nor U24912 (N_24912,N_24458,N_24298);
or U24913 (N_24913,N_24345,N_24293);
nand U24914 (N_24914,N_24165,N_24281);
and U24915 (N_24915,N_24239,N_24303);
xor U24916 (N_24916,N_24129,N_24124);
nor U24917 (N_24917,N_24236,N_24206);
xor U24918 (N_24918,N_24162,N_24331);
nor U24919 (N_24919,N_24183,N_24129);
and U24920 (N_24920,N_24350,N_24392);
nor U24921 (N_24921,N_24476,N_24489);
nor U24922 (N_24922,N_24390,N_24339);
or U24923 (N_24923,N_24155,N_24314);
nand U24924 (N_24924,N_24280,N_24185);
nor U24925 (N_24925,N_24174,N_24065);
nand U24926 (N_24926,N_24042,N_24235);
xnor U24927 (N_24927,N_24300,N_24085);
nand U24928 (N_24928,N_24068,N_24419);
and U24929 (N_24929,N_24138,N_24329);
or U24930 (N_24930,N_24129,N_24145);
and U24931 (N_24931,N_24498,N_24455);
and U24932 (N_24932,N_24330,N_24172);
or U24933 (N_24933,N_24179,N_24372);
nor U24934 (N_24934,N_24215,N_24442);
xor U24935 (N_24935,N_24047,N_24339);
nor U24936 (N_24936,N_24353,N_24409);
nand U24937 (N_24937,N_24189,N_24368);
xor U24938 (N_24938,N_24208,N_24493);
xnor U24939 (N_24939,N_24275,N_24483);
nor U24940 (N_24940,N_24453,N_24449);
and U24941 (N_24941,N_24379,N_24204);
xnor U24942 (N_24942,N_24447,N_24378);
nor U24943 (N_24943,N_24295,N_24424);
or U24944 (N_24944,N_24254,N_24078);
nor U24945 (N_24945,N_24116,N_24086);
nor U24946 (N_24946,N_24150,N_24256);
nor U24947 (N_24947,N_24247,N_24456);
xor U24948 (N_24948,N_24117,N_24475);
nand U24949 (N_24949,N_24302,N_24478);
or U24950 (N_24950,N_24202,N_24231);
nand U24951 (N_24951,N_24186,N_24322);
or U24952 (N_24952,N_24142,N_24426);
or U24953 (N_24953,N_24426,N_24187);
xnor U24954 (N_24954,N_24170,N_24429);
nand U24955 (N_24955,N_24190,N_24207);
nand U24956 (N_24956,N_24433,N_24318);
and U24957 (N_24957,N_24125,N_24091);
nor U24958 (N_24958,N_24077,N_24468);
xnor U24959 (N_24959,N_24030,N_24159);
xor U24960 (N_24960,N_24138,N_24498);
and U24961 (N_24961,N_24053,N_24082);
or U24962 (N_24962,N_24485,N_24224);
and U24963 (N_24963,N_24200,N_24411);
nor U24964 (N_24964,N_24252,N_24376);
or U24965 (N_24965,N_24049,N_24329);
nor U24966 (N_24966,N_24010,N_24230);
nor U24967 (N_24967,N_24156,N_24155);
or U24968 (N_24968,N_24434,N_24361);
or U24969 (N_24969,N_24228,N_24224);
xnor U24970 (N_24970,N_24251,N_24443);
and U24971 (N_24971,N_24453,N_24373);
or U24972 (N_24972,N_24274,N_24232);
and U24973 (N_24973,N_24054,N_24364);
xor U24974 (N_24974,N_24150,N_24201);
and U24975 (N_24975,N_24031,N_24317);
xor U24976 (N_24976,N_24182,N_24249);
nor U24977 (N_24977,N_24271,N_24424);
nor U24978 (N_24978,N_24261,N_24085);
nor U24979 (N_24979,N_24413,N_24074);
nand U24980 (N_24980,N_24216,N_24163);
and U24981 (N_24981,N_24185,N_24437);
nand U24982 (N_24982,N_24188,N_24109);
nand U24983 (N_24983,N_24305,N_24013);
and U24984 (N_24984,N_24328,N_24262);
and U24985 (N_24985,N_24437,N_24353);
nor U24986 (N_24986,N_24305,N_24104);
nand U24987 (N_24987,N_24044,N_24117);
or U24988 (N_24988,N_24307,N_24331);
or U24989 (N_24989,N_24131,N_24075);
or U24990 (N_24990,N_24436,N_24247);
nor U24991 (N_24991,N_24250,N_24203);
nand U24992 (N_24992,N_24105,N_24294);
nand U24993 (N_24993,N_24092,N_24195);
nand U24994 (N_24994,N_24254,N_24116);
nand U24995 (N_24995,N_24136,N_24040);
and U24996 (N_24996,N_24495,N_24085);
xnor U24997 (N_24997,N_24018,N_24428);
nor U24998 (N_24998,N_24390,N_24355);
and U24999 (N_24999,N_24297,N_24222);
nand U25000 (N_25000,N_24885,N_24533);
xnor U25001 (N_25001,N_24626,N_24792);
xnor U25002 (N_25002,N_24699,N_24754);
nor U25003 (N_25003,N_24982,N_24538);
and U25004 (N_25004,N_24740,N_24537);
or U25005 (N_25005,N_24513,N_24834);
nand U25006 (N_25006,N_24749,N_24735);
nor U25007 (N_25007,N_24852,N_24633);
nand U25008 (N_25008,N_24644,N_24684);
xnor U25009 (N_25009,N_24935,N_24845);
xnor U25010 (N_25010,N_24587,N_24772);
and U25011 (N_25011,N_24958,N_24655);
xor U25012 (N_25012,N_24803,N_24500);
and U25013 (N_25013,N_24777,N_24704);
nor U25014 (N_25014,N_24534,N_24857);
or U25015 (N_25015,N_24530,N_24584);
and U25016 (N_25016,N_24940,N_24952);
nand U25017 (N_25017,N_24739,N_24931);
nor U25018 (N_25018,N_24599,N_24720);
nor U25019 (N_25019,N_24631,N_24971);
and U25020 (N_25020,N_24868,N_24645);
nand U25021 (N_25021,N_24515,N_24997);
or U25022 (N_25022,N_24681,N_24510);
and U25023 (N_25023,N_24966,N_24719);
and U25024 (N_25024,N_24815,N_24901);
nor U25025 (N_25025,N_24891,N_24934);
nor U25026 (N_25026,N_24668,N_24665);
nand U25027 (N_25027,N_24718,N_24562);
xor U25028 (N_25028,N_24503,N_24814);
nor U25029 (N_25029,N_24551,N_24524);
nor U25030 (N_25030,N_24862,N_24799);
or U25031 (N_25031,N_24957,N_24567);
xnor U25032 (N_25032,N_24673,N_24566);
and U25033 (N_25033,N_24948,N_24913);
nor U25034 (N_25034,N_24775,N_24748);
xor U25035 (N_25035,N_24701,N_24653);
and U25036 (N_25036,N_24797,N_24585);
xor U25037 (N_25037,N_24568,N_24927);
nor U25038 (N_25038,N_24519,N_24962);
xor U25039 (N_25039,N_24604,N_24542);
and U25040 (N_25040,N_24933,N_24677);
xnor U25041 (N_25041,N_24564,N_24911);
xor U25042 (N_25042,N_24511,N_24759);
and U25043 (N_25043,N_24916,N_24922);
nand U25044 (N_25044,N_24976,N_24611);
and U25045 (N_25045,N_24540,N_24967);
nor U25046 (N_25046,N_24992,N_24643);
and U25047 (N_25047,N_24581,N_24921);
and U25048 (N_25048,N_24732,N_24810);
nor U25049 (N_25049,N_24809,N_24918);
or U25050 (N_25050,N_24696,N_24595);
xor U25051 (N_25051,N_24906,N_24629);
nor U25052 (N_25052,N_24963,N_24956);
or U25053 (N_25053,N_24794,N_24782);
and U25054 (N_25054,N_24742,N_24915);
or U25055 (N_25055,N_24985,N_24787);
xnor U25056 (N_25056,N_24640,N_24838);
xor U25057 (N_25057,N_24709,N_24688);
xor U25058 (N_25058,N_24725,N_24898);
nand U25059 (N_25059,N_24778,N_24945);
nand U25060 (N_25060,N_24618,N_24726);
and U25061 (N_25061,N_24846,N_24817);
xnor U25062 (N_25062,N_24751,N_24964);
or U25063 (N_25063,N_24990,N_24711);
nor U25064 (N_25064,N_24907,N_24569);
and U25065 (N_25065,N_24526,N_24950);
or U25066 (N_25066,N_24892,N_24578);
or U25067 (N_25067,N_24986,N_24924);
nor U25068 (N_25068,N_24975,N_24501);
and U25069 (N_25069,N_24822,N_24682);
xor U25070 (N_25070,N_24779,N_24687);
or U25071 (N_25071,N_24756,N_24965);
or U25072 (N_25072,N_24660,N_24552);
xor U25073 (N_25073,N_24840,N_24606);
xnor U25074 (N_25074,N_24766,N_24555);
xnor U25075 (N_25075,N_24616,N_24580);
and U25076 (N_25076,N_24662,N_24747);
xor U25077 (N_25077,N_24991,N_24758);
xor U25078 (N_25078,N_24657,N_24883);
or U25079 (N_25079,N_24661,N_24713);
or U25080 (N_25080,N_24832,N_24805);
nand U25081 (N_25081,N_24752,N_24613);
nor U25082 (N_25082,N_24977,N_24521);
nand U25083 (N_25083,N_24853,N_24692);
and U25084 (N_25084,N_24548,N_24903);
or U25085 (N_25085,N_24955,N_24667);
xnor U25086 (N_25086,N_24850,N_24535);
or U25087 (N_25087,N_24763,N_24638);
nand U25088 (N_25088,N_24532,N_24553);
nor U25089 (N_25089,N_24917,N_24848);
xor U25090 (N_25090,N_24813,N_24539);
xnor U25091 (N_25091,N_24762,N_24820);
nor U25092 (N_25092,N_24972,N_24531);
and U25093 (N_25093,N_24855,N_24802);
nand U25094 (N_25094,N_24959,N_24690);
and U25095 (N_25095,N_24887,N_24973);
or U25096 (N_25096,N_24801,N_24741);
xor U25097 (N_25097,N_24880,N_24789);
or U25098 (N_25098,N_24761,N_24560);
nor U25099 (N_25099,N_24517,N_24575);
or U25100 (N_25100,N_24561,N_24942);
nor U25101 (N_25101,N_24625,N_24523);
nor U25102 (N_25102,N_24632,N_24926);
xor U25103 (N_25103,N_24755,N_24938);
and U25104 (N_25104,N_24571,N_24818);
or U25105 (N_25105,N_24793,N_24819);
nor U25106 (N_25106,N_24894,N_24858);
and U25107 (N_25107,N_24508,N_24574);
nor U25108 (N_25108,N_24823,N_24708);
xnor U25109 (N_25109,N_24695,N_24603);
and U25110 (N_25110,N_24981,N_24659);
and U25111 (N_25111,N_24577,N_24786);
nand U25112 (N_25112,N_24974,N_24544);
and U25113 (N_25113,N_24920,N_24860);
nand U25114 (N_25114,N_24863,N_24723);
nor U25115 (N_25115,N_24602,N_24827);
nor U25116 (N_25116,N_24745,N_24543);
or U25117 (N_25117,N_24825,N_24694);
or U25118 (N_25118,N_24506,N_24698);
nor U25119 (N_25119,N_24522,N_24944);
nand U25120 (N_25120,N_24769,N_24502);
nand U25121 (N_25121,N_24843,N_24930);
and U25122 (N_25122,N_24656,N_24686);
xor U25123 (N_25123,N_24649,N_24685);
or U25124 (N_25124,N_24984,N_24689);
xnor U25125 (N_25125,N_24791,N_24664);
xnor U25126 (N_25126,N_24619,N_24676);
or U25127 (N_25127,N_24856,N_24788);
xor U25128 (N_25128,N_24703,N_24837);
or U25129 (N_25129,N_24893,N_24909);
and U25130 (N_25130,N_24724,N_24760);
and U25131 (N_25131,N_24648,N_24528);
and U25132 (N_25132,N_24881,N_24637);
nand U25133 (N_25133,N_24798,N_24650);
nor U25134 (N_25134,N_24878,N_24890);
and U25135 (N_25135,N_24558,N_24936);
nor U25136 (N_25136,N_24851,N_24888);
nor U25137 (N_25137,N_24663,N_24615);
xnor U25138 (N_25138,N_24705,N_24919);
and U25139 (N_25139,N_24872,N_24570);
and U25140 (N_25140,N_24614,N_24721);
nor U25141 (N_25141,N_24716,N_24807);
nor U25142 (N_25142,N_24597,N_24849);
and U25143 (N_25143,N_24784,N_24678);
nor U25144 (N_25144,N_24764,N_24557);
nand U25145 (N_25145,N_24646,N_24623);
xnor U25146 (N_25146,N_24527,N_24790);
or U25147 (N_25147,N_24999,N_24712);
xor U25148 (N_25148,N_24811,N_24556);
nand U25149 (N_25149,N_24546,N_24854);
and U25150 (N_25150,N_24715,N_24969);
and U25151 (N_25151,N_24842,N_24579);
nand U25152 (N_25152,N_24620,N_24744);
nor U25153 (N_25153,N_24925,N_24714);
nand U25154 (N_25154,N_24536,N_24844);
xnor U25155 (N_25155,N_24598,N_24871);
or U25156 (N_25156,N_24547,N_24841);
or U25157 (N_25157,N_24554,N_24774);
or U25158 (N_25158,N_24833,N_24796);
xor U25159 (N_25159,N_24882,N_24672);
nand U25160 (N_25160,N_24954,N_24781);
nand U25161 (N_25161,N_24884,N_24504);
xnor U25162 (N_25162,N_24905,N_24586);
and U25163 (N_25163,N_24867,N_24812);
nor U25164 (N_25164,N_24675,N_24970);
nor U25165 (N_25165,N_24874,N_24624);
or U25166 (N_25166,N_24590,N_24647);
nor U25167 (N_25167,N_24943,N_24785);
xnor U25168 (N_25168,N_24601,N_24979);
xnor U25169 (N_25169,N_24549,N_24953);
nor U25170 (N_25170,N_24988,N_24731);
or U25171 (N_25171,N_24592,N_24859);
nand U25172 (N_25172,N_24671,N_24768);
nand U25173 (N_25173,N_24877,N_24697);
nand U25174 (N_25174,N_24621,N_24666);
nand U25175 (N_25175,N_24847,N_24896);
and U25176 (N_25176,N_24565,N_24995);
nand U25177 (N_25177,N_24563,N_24706);
nand U25178 (N_25178,N_24545,N_24722);
and U25179 (N_25179,N_24669,N_24989);
xor U25180 (N_25180,N_24912,N_24873);
nor U25181 (N_25181,N_24937,N_24830);
nor U25182 (N_25182,N_24652,N_24869);
and U25183 (N_25183,N_24609,N_24826);
or U25184 (N_25184,N_24861,N_24900);
nor U25185 (N_25185,N_24776,N_24836);
nand U25186 (N_25186,N_24824,N_24939);
and U25187 (N_25187,N_24910,N_24505);
xnor U25188 (N_25188,N_24983,N_24780);
and U25189 (N_25189,N_24866,N_24512);
nor U25190 (N_25190,N_24757,N_24765);
xor U25191 (N_25191,N_24717,N_24738);
or U25192 (N_25192,N_24641,N_24808);
and U25193 (N_25193,N_24914,N_24516);
or U25194 (N_25194,N_24951,N_24541);
nand U25195 (N_25195,N_24583,N_24899);
nand U25196 (N_25196,N_24897,N_24932);
or U25197 (N_25197,N_24870,N_24691);
nand U25198 (N_25198,N_24902,N_24771);
nor U25199 (N_25199,N_24831,N_24642);
xor U25200 (N_25200,N_24929,N_24821);
nor U25201 (N_25201,N_24593,N_24617);
or U25202 (N_25202,N_24839,N_24507);
xor U25203 (N_25203,N_24730,N_24634);
and U25204 (N_25204,N_24978,N_24835);
nand U25205 (N_25205,N_24576,N_24743);
nand U25206 (N_25206,N_24514,N_24700);
and U25207 (N_25207,N_24996,N_24795);
nand U25208 (N_25208,N_24736,N_24733);
nand U25209 (N_25209,N_24600,N_24591);
nand U25210 (N_25210,N_24947,N_24949);
xor U25211 (N_25211,N_24800,N_24594);
nand U25212 (N_25212,N_24816,N_24679);
or U25213 (N_25213,N_24734,N_24550);
nand U25214 (N_25214,N_24589,N_24980);
xor U25215 (N_25215,N_24773,N_24895);
xor U25216 (N_25216,N_24630,N_24710);
and U25217 (N_25217,N_24509,N_24702);
xnor U25218 (N_25218,N_24559,N_24889);
and U25219 (N_25219,N_24573,N_24728);
nor U25220 (N_25220,N_24828,N_24683);
and U25221 (N_25221,N_24960,N_24804);
nor U25222 (N_25222,N_24612,N_24968);
or U25223 (N_25223,N_24904,N_24572);
nor U25224 (N_25224,N_24635,N_24865);
and U25225 (N_25225,N_24627,N_24670);
or U25226 (N_25226,N_24987,N_24622);
nand U25227 (N_25227,N_24727,N_24993);
xor U25228 (N_25228,N_24636,N_24886);
nor U25229 (N_25229,N_24876,N_24783);
or U25230 (N_25230,N_24767,N_24607);
nand U25231 (N_25231,N_24529,N_24525);
nor U25232 (N_25232,N_24864,N_24753);
and U25233 (N_25233,N_24707,N_24605);
or U25234 (N_25234,N_24674,N_24651);
nand U25235 (N_25235,N_24941,N_24829);
or U25236 (N_25236,N_24770,N_24596);
xnor U25237 (N_25237,N_24654,N_24875);
or U25238 (N_25238,N_24658,N_24908);
nand U25239 (N_25239,N_24923,N_24750);
or U25240 (N_25240,N_24518,N_24994);
nor U25241 (N_25241,N_24610,N_24928);
xnor U25242 (N_25242,N_24806,N_24737);
nand U25243 (N_25243,N_24520,N_24729);
nor U25244 (N_25244,N_24582,N_24639);
nor U25245 (N_25245,N_24588,N_24693);
and U25246 (N_25246,N_24879,N_24628);
nor U25247 (N_25247,N_24680,N_24608);
nand U25248 (N_25248,N_24946,N_24746);
nor U25249 (N_25249,N_24961,N_24998);
or U25250 (N_25250,N_24657,N_24827);
or U25251 (N_25251,N_24592,N_24551);
xor U25252 (N_25252,N_24868,N_24658);
xnor U25253 (N_25253,N_24607,N_24940);
nand U25254 (N_25254,N_24924,N_24964);
xnor U25255 (N_25255,N_24993,N_24617);
or U25256 (N_25256,N_24513,N_24882);
or U25257 (N_25257,N_24851,N_24702);
nand U25258 (N_25258,N_24970,N_24876);
or U25259 (N_25259,N_24846,N_24535);
nor U25260 (N_25260,N_24888,N_24798);
nand U25261 (N_25261,N_24667,N_24562);
and U25262 (N_25262,N_24505,N_24611);
nand U25263 (N_25263,N_24614,N_24727);
and U25264 (N_25264,N_24962,N_24740);
nand U25265 (N_25265,N_24820,N_24617);
or U25266 (N_25266,N_24735,N_24620);
and U25267 (N_25267,N_24994,N_24937);
nor U25268 (N_25268,N_24747,N_24502);
nor U25269 (N_25269,N_24919,N_24864);
nor U25270 (N_25270,N_24725,N_24678);
nor U25271 (N_25271,N_24653,N_24752);
xor U25272 (N_25272,N_24829,N_24532);
xor U25273 (N_25273,N_24796,N_24884);
nor U25274 (N_25274,N_24835,N_24617);
or U25275 (N_25275,N_24773,N_24687);
xor U25276 (N_25276,N_24885,N_24940);
or U25277 (N_25277,N_24847,N_24664);
xor U25278 (N_25278,N_24992,N_24618);
or U25279 (N_25279,N_24729,N_24773);
nand U25280 (N_25280,N_24645,N_24526);
nor U25281 (N_25281,N_24698,N_24558);
or U25282 (N_25282,N_24792,N_24627);
xnor U25283 (N_25283,N_24868,N_24527);
xor U25284 (N_25284,N_24668,N_24885);
or U25285 (N_25285,N_24851,N_24709);
and U25286 (N_25286,N_24834,N_24739);
xor U25287 (N_25287,N_24877,N_24716);
or U25288 (N_25288,N_24953,N_24943);
nand U25289 (N_25289,N_24515,N_24645);
xor U25290 (N_25290,N_24922,N_24810);
or U25291 (N_25291,N_24718,N_24845);
xor U25292 (N_25292,N_24547,N_24964);
nor U25293 (N_25293,N_24782,N_24545);
nor U25294 (N_25294,N_24872,N_24915);
xnor U25295 (N_25295,N_24559,N_24652);
and U25296 (N_25296,N_24665,N_24707);
nor U25297 (N_25297,N_24601,N_24603);
xnor U25298 (N_25298,N_24875,N_24928);
and U25299 (N_25299,N_24932,N_24801);
xnor U25300 (N_25300,N_24610,N_24861);
xnor U25301 (N_25301,N_24601,N_24559);
and U25302 (N_25302,N_24982,N_24689);
or U25303 (N_25303,N_24525,N_24558);
xnor U25304 (N_25304,N_24559,N_24756);
or U25305 (N_25305,N_24621,N_24955);
or U25306 (N_25306,N_24862,N_24820);
nor U25307 (N_25307,N_24555,N_24700);
nor U25308 (N_25308,N_24573,N_24730);
xor U25309 (N_25309,N_24714,N_24526);
xor U25310 (N_25310,N_24847,N_24841);
nand U25311 (N_25311,N_24691,N_24506);
and U25312 (N_25312,N_24944,N_24733);
xnor U25313 (N_25313,N_24843,N_24711);
xor U25314 (N_25314,N_24525,N_24747);
nand U25315 (N_25315,N_24713,N_24897);
nor U25316 (N_25316,N_24964,N_24775);
nor U25317 (N_25317,N_24700,N_24546);
nor U25318 (N_25318,N_24722,N_24694);
xnor U25319 (N_25319,N_24722,N_24639);
and U25320 (N_25320,N_24588,N_24572);
nand U25321 (N_25321,N_24590,N_24996);
xnor U25322 (N_25322,N_24794,N_24752);
and U25323 (N_25323,N_24818,N_24804);
xnor U25324 (N_25324,N_24669,N_24611);
xnor U25325 (N_25325,N_24709,N_24588);
nor U25326 (N_25326,N_24832,N_24621);
nor U25327 (N_25327,N_24916,N_24789);
or U25328 (N_25328,N_24946,N_24535);
or U25329 (N_25329,N_24908,N_24845);
nor U25330 (N_25330,N_24740,N_24817);
or U25331 (N_25331,N_24822,N_24913);
and U25332 (N_25332,N_24862,N_24564);
nor U25333 (N_25333,N_24794,N_24883);
and U25334 (N_25334,N_24917,N_24518);
and U25335 (N_25335,N_24651,N_24628);
xnor U25336 (N_25336,N_24819,N_24761);
and U25337 (N_25337,N_24815,N_24526);
nor U25338 (N_25338,N_24524,N_24821);
nor U25339 (N_25339,N_24609,N_24539);
nand U25340 (N_25340,N_24890,N_24545);
xor U25341 (N_25341,N_24744,N_24577);
xnor U25342 (N_25342,N_24985,N_24684);
nand U25343 (N_25343,N_24861,N_24836);
or U25344 (N_25344,N_24847,N_24812);
nand U25345 (N_25345,N_24945,N_24843);
nor U25346 (N_25346,N_24789,N_24941);
and U25347 (N_25347,N_24827,N_24704);
or U25348 (N_25348,N_24879,N_24546);
xor U25349 (N_25349,N_24677,N_24654);
or U25350 (N_25350,N_24673,N_24546);
xor U25351 (N_25351,N_24594,N_24587);
nand U25352 (N_25352,N_24674,N_24891);
and U25353 (N_25353,N_24579,N_24944);
xnor U25354 (N_25354,N_24984,N_24843);
or U25355 (N_25355,N_24851,N_24651);
nor U25356 (N_25356,N_24971,N_24584);
and U25357 (N_25357,N_24877,N_24876);
and U25358 (N_25358,N_24769,N_24999);
or U25359 (N_25359,N_24826,N_24610);
xor U25360 (N_25360,N_24934,N_24788);
or U25361 (N_25361,N_24830,N_24942);
xor U25362 (N_25362,N_24520,N_24727);
or U25363 (N_25363,N_24561,N_24598);
and U25364 (N_25364,N_24966,N_24515);
nor U25365 (N_25365,N_24871,N_24535);
and U25366 (N_25366,N_24663,N_24761);
nand U25367 (N_25367,N_24716,N_24960);
or U25368 (N_25368,N_24615,N_24948);
nand U25369 (N_25369,N_24547,N_24721);
or U25370 (N_25370,N_24994,N_24740);
or U25371 (N_25371,N_24795,N_24824);
nor U25372 (N_25372,N_24913,N_24532);
nor U25373 (N_25373,N_24560,N_24882);
and U25374 (N_25374,N_24944,N_24595);
nand U25375 (N_25375,N_24606,N_24728);
nand U25376 (N_25376,N_24973,N_24858);
xor U25377 (N_25377,N_24607,N_24861);
nor U25378 (N_25378,N_24953,N_24759);
xnor U25379 (N_25379,N_24556,N_24807);
or U25380 (N_25380,N_24533,N_24654);
nor U25381 (N_25381,N_24828,N_24982);
nand U25382 (N_25382,N_24775,N_24850);
xnor U25383 (N_25383,N_24711,N_24691);
or U25384 (N_25384,N_24792,N_24523);
nand U25385 (N_25385,N_24568,N_24995);
and U25386 (N_25386,N_24531,N_24746);
xor U25387 (N_25387,N_24885,N_24563);
and U25388 (N_25388,N_24937,N_24807);
xor U25389 (N_25389,N_24578,N_24644);
nand U25390 (N_25390,N_24726,N_24774);
or U25391 (N_25391,N_24841,N_24512);
nand U25392 (N_25392,N_24948,N_24733);
and U25393 (N_25393,N_24648,N_24862);
or U25394 (N_25394,N_24660,N_24511);
nor U25395 (N_25395,N_24640,N_24944);
xnor U25396 (N_25396,N_24847,N_24733);
xnor U25397 (N_25397,N_24733,N_24951);
or U25398 (N_25398,N_24769,N_24747);
nand U25399 (N_25399,N_24991,N_24725);
or U25400 (N_25400,N_24829,N_24503);
or U25401 (N_25401,N_24616,N_24766);
nand U25402 (N_25402,N_24881,N_24821);
xnor U25403 (N_25403,N_24591,N_24554);
or U25404 (N_25404,N_24867,N_24965);
and U25405 (N_25405,N_24537,N_24948);
and U25406 (N_25406,N_24863,N_24757);
nand U25407 (N_25407,N_24830,N_24505);
xor U25408 (N_25408,N_24770,N_24814);
or U25409 (N_25409,N_24636,N_24581);
and U25410 (N_25410,N_24948,N_24981);
nand U25411 (N_25411,N_24956,N_24874);
nand U25412 (N_25412,N_24837,N_24638);
or U25413 (N_25413,N_24962,N_24969);
and U25414 (N_25414,N_24514,N_24550);
xor U25415 (N_25415,N_24804,N_24512);
nor U25416 (N_25416,N_24530,N_24585);
nand U25417 (N_25417,N_24619,N_24991);
nand U25418 (N_25418,N_24761,N_24576);
and U25419 (N_25419,N_24663,N_24774);
or U25420 (N_25420,N_24657,N_24547);
or U25421 (N_25421,N_24613,N_24962);
nand U25422 (N_25422,N_24870,N_24935);
or U25423 (N_25423,N_24802,N_24660);
or U25424 (N_25424,N_24690,N_24732);
or U25425 (N_25425,N_24907,N_24600);
nand U25426 (N_25426,N_24820,N_24831);
nor U25427 (N_25427,N_24934,N_24899);
nor U25428 (N_25428,N_24991,N_24990);
nand U25429 (N_25429,N_24739,N_24895);
nand U25430 (N_25430,N_24637,N_24519);
nand U25431 (N_25431,N_24653,N_24793);
and U25432 (N_25432,N_24549,N_24720);
and U25433 (N_25433,N_24821,N_24728);
and U25434 (N_25434,N_24777,N_24745);
or U25435 (N_25435,N_24720,N_24647);
nor U25436 (N_25436,N_24949,N_24911);
xor U25437 (N_25437,N_24677,N_24928);
xnor U25438 (N_25438,N_24886,N_24907);
or U25439 (N_25439,N_24691,N_24576);
nor U25440 (N_25440,N_24505,N_24583);
or U25441 (N_25441,N_24699,N_24501);
nand U25442 (N_25442,N_24703,N_24933);
xor U25443 (N_25443,N_24893,N_24980);
and U25444 (N_25444,N_24557,N_24827);
nand U25445 (N_25445,N_24670,N_24589);
and U25446 (N_25446,N_24963,N_24882);
xnor U25447 (N_25447,N_24874,N_24751);
or U25448 (N_25448,N_24708,N_24535);
nand U25449 (N_25449,N_24989,N_24837);
or U25450 (N_25450,N_24916,N_24943);
nand U25451 (N_25451,N_24725,N_24964);
nand U25452 (N_25452,N_24864,N_24763);
xnor U25453 (N_25453,N_24649,N_24723);
xor U25454 (N_25454,N_24724,N_24755);
xnor U25455 (N_25455,N_24822,N_24686);
or U25456 (N_25456,N_24736,N_24712);
xor U25457 (N_25457,N_24980,N_24812);
nor U25458 (N_25458,N_24592,N_24986);
nor U25459 (N_25459,N_24854,N_24809);
nor U25460 (N_25460,N_24856,N_24655);
nand U25461 (N_25461,N_24590,N_24709);
nand U25462 (N_25462,N_24925,N_24507);
nand U25463 (N_25463,N_24752,N_24711);
xnor U25464 (N_25464,N_24626,N_24714);
or U25465 (N_25465,N_24685,N_24678);
xnor U25466 (N_25466,N_24619,N_24869);
and U25467 (N_25467,N_24513,N_24830);
xnor U25468 (N_25468,N_24698,N_24938);
xnor U25469 (N_25469,N_24778,N_24510);
nand U25470 (N_25470,N_24672,N_24579);
nor U25471 (N_25471,N_24962,N_24676);
nand U25472 (N_25472,N_24553,N_24520);
or U25473 (N_25473,N_24607,N_24776);
xnor U25474 (N_25474,N_24731,N_24823);
xnor U25475 (N_25475,N_24667,N_24748);
nor U25476 (N_25476,N_24886,N_24667);
and U25477 (N_25477,N_24987,N_24802);
and U25478 (N_25478,N_24947,N_24556);
nor U25479 (N_25479,N_24543,N_24802);
and U25480 (N_25480,N_24939,N_24868);
nand U25481 (N_25481,N_24644,N_24742);
nor U25482 (N_25482,N_24506,N_24897);
or U25483 (N_25483,N_24539,N_24633);
xnor U25484 (N_25484,N_24977,N_24985);
and U25485 (N_25485,N_24976,N_24561);
xor U25486 (N_25486,N_24628,N_24781);
or U25487 (N_25487,N_24686,N_24636);
nor U25488 (N_25488,N_24553,N_24723);
and U25489 (N_25489,N_24603,N_24723);
nand U25490 (N_25490,N_24821,N_24825);
and U25491 (N_25491,N_24710,N_24712);
xnor U25492 (N_25492,N_24959,N_24937);
xnor U25493 (N_25493,N_24702,N_24986);
nor U25494 (N_25494,N_24615,N_24507);
and U25495 (N_25495,N_24995,N_24893);
xnor U25496 (N_25496,N_24562,N_24757);
and U25497 (N_25497,N_24637,N_24682);
xnor U25498 (N_25498,N_24872,N_24826);
nor U25499 (N_25499,N_24546,N_24667);
nand U25500 (N_25500,N_25364,N_25420);
or U25501 (N_25501,N_25133,N_25129);
nand U25502 (N_25502,N_25235,N_25011);
nor U25503 (N_25503,N_25348,N_25093);
nand U25504 (N_25504,N_25338,N_25095);
or U25505 (N_25505,N_25271,N_25044);
nand U25506 (N_25506,N_25322,N_25302);
and U25507 (N_25507,N_25466,N_25134);
nand U25508 (N_25508,N_25279,N_25376);
and U25509 (N_25509,N_25113,N_25075);
nor U25510 (N_25510,N_25243,N_25265);
nand U25511 (N_25511,N_25051,N_25112);
nand U25512 (N_25512,N_25216,N_25189);
and U25513 (N_25513,N_25452,N_25146);
or U25514 (N_25514,N_25124,N_25144);
nand U25515 (N_25515,N_25008,N_25222);
xnor U25516 (N_25516,N_25223,N_25212);
nand U25517 (N_25517,N_25491,N_25142);
or U25518 (N_25518,N_25307,N_25204);
nand U25519 (N_25519,N_25382,N_25337);
xor U25520 (N_25520,N_25476,N_25018);
nand U25521 (N_25521,N_25464,N_25050);
xor U25522 (N_25522,N_25237,N_25393);
nor U25523 (N_25523,N_25045,N_25236);
nor U25524 (N_25524,N_25082,N_25114);
xnor U25525 (N_25525,N_25149,N_25024);
or U25526 (N_25526,N_25168,N_25202);
nor U25527 (N_25527,N_25078,N_25296);
nand U25528 (N_25528,N_25274,N_25319);
nor U25529 (N_25529,N_25176,N_25010);
xnor U25530 (N_25530,N_25059,N_25211);
and U25531 (N_25531,N_25346,N_25173);
and U25532 (N_25532,N_25115,N_25229);
and U25533 (N_25533,N_25012,N_25039);
nand U25534 (N_25534,N_25109,N_25436);
or U25535 (N_25535,N_25431,N_25259);
nor U25536 (N_25536,N_25118,N_25401);
nor U25537 (N_25537,N_25290,N_25323);
nor U25538 (N_25538,N_25298,N_25384);
and U25539 (N_25539,N_25282,N_25254);
xnor U25540 (N_25540,N_25398,N_25230);
and U25541 (N_25541,N_25154,N_25281);
nand U25542 (N_25542,N_25448,N_25005);
xor U25543 (N_25543,N_25092,N_25485);
nand U25544 (N_25544,N_25200,N_25349);
nor U25545 (N_25545,N_25233,N_25308);
or U25546 (N_25546,N_25358,N_25463);
and U25547 (N_25547,N_25170,N_25494);
or U25548 (N_25548,N_25457,N_25096);
nand U25549 (N_25549,N_25462,N_25294);
xnor U25550 (N_25550,N_25369,N_25194);
and U25551 (N_25551,N_25185,N_25107);
and U25552 (N_25552,N_25057,N_25079);
nand U25553 (N_25553,N_25140,N_25496);
or U25554 (N_25554,N_25071,N_25207);
nor U25555 (N_25555,N_25120,N_25110);
or U25556 (N_25556,N_25231,N_25397);
xnor U25557 (N_25557,N_25460,N_25101);
xnor U25558 (N_25558,N_25312,N_25257);
nand U25559 (N_25559,N_25385,N_25210);
nor U25560 (N_25560,N_25374,N_25127);
nand U25561 (N_25561,N_25013,N_25316);
or U25562 (N_25562,N_25378,N_25326);
nor U25563 (N_25563,N_25089,N_25042);
nor U25564 (N_25564,N_25002,N_25126);
nor U25565 (N_25565,N_25329,N_25111);
and U25566 (N_25566,N_25219,N_25062);
xnor U25567 (N_25567,N_25411,N_25108);
nor U25568 (N_25568,N_25291,N_25400);
or U25569 (N_25569,N_25106,N_25284);
xnor U25570 (N_25570,N_25440,N_25234);
xnor U25571 (N_25571,N_25285,N_25371);
nand U25572 (N_25572,N_25052,N_25297);
and U25573 (N_25573,N_25341,N_25033);
xnor U25574 (N_25574,N_25343,N_25069);
and U25575 (N_25575,N_25418,N_25487);
or U25576 (N_25576,N_25060,N_25488);
nor U25577 (N_25577,N_25416,N_25152);
xnor U25578 (N_25578,N_25232,N_25255);
xnor U25579 (N_25579,N_25034,N_25193);
nand U25580 (N_25580,N_25131,N_25245);
or U25581 (N_25581,N_25339,N_25186);
xnor U25582 (N_25582,N_25141,N_25276);
and U25583 (N_25583,N_25305,N_25187);
nor U25584 (N_25584,N_25153,N_25399);
xnor U25585 (N_25585,N_25188,N_25482);
nand U25586 (N_25586,N_25102,N_25434);
or U25587 (N_25587,N_25354,N_25270);
nor U25588 (N_25588,N_25099,N_25077);
nand U25589 (N_25589,N_25480,N_25438);
nand U25590 (N_25590,N_25150,N_25098);
and U25591 (N_25591,N_25227,N_25492);
nor U25592 (N_25592,N_25481,N_25461);
or U25593 (N_25593,N_25250,N_25363);
xnor U25594 (N_25594,N_25471,N_25321);
xnor U25595 (N_25595,N_25449,N_25361);
and U25596 (N_25596,N_25201,N_25238);
nor U25597 (N_25597,N_25064,N_25084);
or U25598 (N_25598,N_25428,N_25320);
nand U25599 (N_25599,N_25286,N_25396);
nor U25600 (N_25600,N_25088,N_25309);
nand U25601 (N_25601,N_25182,N_25006);
nand U25602 (N_25602,N_25100,N_25003);
and U25603 (N_25603,N_25375,N_25038);
nor U25604 (N_25604,N_25067,N_25446);
nor U25605 (N_25605,N_25221,N_25454);
nor U25606 (N_25606,N_25184,N_25432);
nor U25607 (N_25607,N_25001,N_25162);
nand U25608 (N_25608,N_25347,N_25292);
xnor U25609 (N_25609,N_25402,N_25391);
xnor U25610 (N_25610,N_25181,N_25264);
xor U25611 (N_25611,N_25097,N_25036);
and U25612 (N_25612,N_25273,N_25444);
xnor U25613 (N_25613,N_25157,N_25335);
xor U25614 (N_25614,N_25239,N_25055);
and U25615 (N_25615,N_25394,N_25000);
nor U25616 (N_25616,N_25165,N_25248);
or U25617 (N_25617,N_25087,N_25315);
and U25618 (N_25618,N_25499,N_25479);
or U25619 (N_25619,N_25373,N_25260);
nand U25620 (N_25620,N_25137,N_25179);
or U25621 (N_25621,N_25405,N_25327);
xor U25622 (N_25622,N_25083,N_25415);
or U25623 (N_25623,N_25081,N_25442);
xnor U25624 (N_25624,N_25392,N_25379);
xnor U25625 (N_25625,N_25228,N_25156);
xnor U25626 (N_25626,N_25249,N_25105);
xor U25627 (N_25627,N_25037,N_25130);
and U25628 (N_25628,N_25443,N_25015);
xnor U25629 (N_25629,N_25251,N_25409);
and U25630 (N_25630,N_25041,N_25388);
nand U25631 (N_25631,N_25117,N_25277);
xnor U25632 (N_25632,N_25342,N_25301);
and U25633 (N_25633,N_25299,N_25498);
nor U25634 (N_25634,N_25021,N_25331);
nor U25635 (N_25635,N_25303,N_25068);
or U25636 (N_25636,N_25429,N_25390);
or U25637 (N_25637,N_25351,N_25287);
nand U25638 (N_25638,N_25203,N_25404);
nor U25639 (N_25639,N_25020,N_25355);
and U25640 (N_25640,N_25340,N_25004);
and U25641 (N_25641,N_25439,N_25225);
nand U25642 (N_25642,N_25447,N_25074);
and U25643 (N_25643,N_25226,N_25258);
and U25644 (N_25644,N_25218,N_25007);
and U25645 (N_25645,N_25043,N_25387);
nor U25646 (N_25646,N_25383,N_25493);
and U25647 (N_25647,N_25275,N_25483);
and U25648 (N_25648,N_25190,N_25160);
and U25649 (N_25649,N_25070,N_25362);
or U25650 (N_25650,N_25336,N_25121);
xnor U25651 (N_25651,N_25430,N_25224);
nand U25652 (N_25652,N_25330,N_25016);
nand U25653 (N_25653,N_25048,N_25198);
and U25654 (N_25654,N_25313,N_25090);
or U25655 (N_25655,N_25054,N_25425);
nor U25656 (N_25656,N_25353,N_25380);
nand U25657 (N_25657,N_25125,N_25453);
or U25658 (N_25658,N_25241,N_25423);
and U25659 (N_25659,N_25386,N_25172);
and U25660 (N_25660,N_25408,N_25132);
nor U25661 (N_25661,N_25459,N_25143);
nor U25662 (N_25662,N_25389,N_25094);
or U25663 (N_25663,N_25147,N_25473);
or U25664 (N_25664,N_25091,N_25197);
nand U25665 (N_25665,N_25161,N_25360);
or U25666 (N_25666,N_25433,N_25441);
nor U25667 (N_25667,N_25325,N_25047);
nor U25668 (N_25668,N_25310,N_25407);
xnor U25669 (N_25669,N_25080,N_25304);
nor U25670 (N_25670,N_25269,N_25475);
nand U25671 (N_25671,N_25497,N_25470);
and U25672 (N_25672,N_25220,N_25177);
nand U25673 (N_25673,N_25300,N_25138);
or U25674 (N_25674,N_25208,N_25159);
nand U25675 (N_25675,N_25023,N_25029);
xor U25676 (N_25676,N_25451,N_25283);
and U25677 (N_25677,N_25246,N_25306);
or U25678 (N_25678,N_25073,N_25116);
nor U25679 (N_25679,N_25345,N_25357);
xnor U25680 (N_25680,N_25410,N_25334);
or U25681 (N_25681,N_25213,N_25065);
and U25682 (N_25682,N_25242,N_25403);
nor U25683 (N_25683,N_25195,N_25318);
or U25684 (N_25684,N_25031,N_25009);
or U25685 (N_25685,N_25040,N_25465);
nand U25686 (N_25686,N_25086,N_25486);
and U25687 (N_25687,N_25427,N_25247);
nor U25688 (N_25688,N_25217,N_25368);
or U25689 (N_25689,N_25139,N_25085);
and U25690 (N_25690,N_25214,N_25046);
nand U25691 (N_25691,N_25215,N_25104);
xnor U25692 (N_25692,N_25458,N_25135);
nand U25693 (N_25693,N_25289,N_25352);
or U25694 (N_25694,N_25350,N_25426);
and U25695 (N_25695,N_25183,N_25295);
nor U25696 (N_25696,N_25252,N_25017);
xnor U25697 (N_25697,N_25474,N_25419);
xor U25698 (N_25698,N_25435,N_25365);
nand U25699 (N_25699,N_25311,N_25063);
nand U25700 (N_25700,N_25490,N_25122);
or U25701 (N_25701,N_25123,N_25367);
nor U25702 (N_25702,N_25026,N_25032);
xnor U25703 (N_25703,N_25192,N_25406);
and U25704 (N_25704,N_25049,N_25167);
xnor U25705 (N_25705,N_25456,N_25293);
xnor U25706 (N_25706,N_25199,N_25035);
and U25707 (N_25707,N_25145,N_25025);
and U25708 (N_25708,N_25437,N_25478);
or U25709 (N_25709,N_25366,N_25395);
or U25710 (N_25710,N_25412,N_25058);
and U25711 (N_25711,N_25477,N_25267);
xnor U25712 (N_25712,N_25261,N_25163);
nor U25713 (N_25713,N_25467,N_25278);
nand U25714 (N_25714,N_25484,N_25148);
xor U25715 (N_25715,N_25030,N_25022);
nor U25716 (N_25716,N_25280,N_25061);
xor U25717 (N_25717,N_25455,N_25171);
nand U25718 (N_25718,N_25332,N_25076);
or U25719 (N_25719,N_25272,N_25468);
and U25720 (N_25720,N_25053,N_25450);
nor U25721 (N_25721,N_25266,N_25469);
xor U25722 (N_25722,N_25262,N_25174);
nor U25723 (N_25723,N_25495,N_25317);
and U25724 (N_25724,N_25263,N_25424);
nor U25725 (N_25725,N_25158,N_25205);
nor U25726 (N_25726,N_25240,N_25019);
xnor U25727 (N_25727,N_25413,N_25253);
nand U25728 (N_25728,N_25119,N_25372);
nor U25729 (N_25729,N_25472,N_25256);
nor U25730 (N_25730,N_25377,N_25066);
nor U25731 (N_25731,N_25206,N_25196);
nor U25732 (N_25732,N_25489,N_25414);
xnor U25733 (N_25733,N_25151,N_25244);
nand U25734 (N_25734,N_25333,N_25136);
nand U25735 (N_25735,N_25370,N_25381);
nand U25736 (N_25736,N_25191,N_25324);
or U25737 (N_25737,N_25209,N_25028);
xor U25738 (N_25738,N_25356,N_25166);
or U25739 (N_25739,N_25178,N_25169);
or U25740 (N_25740,N_25314,N_25445);
nor U25741 (N_25741,N_25359,N_25422);
and U25742 (N_25742,N_25175,N_25072);
nor U25743 (N_25743,N_25128,N_25164);
and U25744 (N_25744,N_25014,N_25103);
and U25745 (N_25745,N_25288,N_25155);
and U25746 (N_25746,N_25027,N_25180);
xor U25747 (N_25747,N_25344,N_25417);
xnor U25748 (N_25748,N_25268,N_25056);
and U25749 (N_25749,N_25328,N_25421);
and U25750 (N_25750,N_25259,N_25401);
nand U25751 (N_25751,N_25466,N_25318);
nand U25752 (N_25752,N_25323,N_25085);
and U25753 (N_25753,N_25211,N_25032);
nand U25754 (N_25754,N_25344,N_25371);
nand U25755 (N_25755,N_25017,N_25105);
nand U25756 (N_25756,N_25270,N_25451);
xor U25757 (N_25757,N_25111,N_25388);
nor U25758 (N_25758,N_25482,N_25474);
nand U25759 (N_25759,N_25138,N_25271);
nand U25760 (N_25760,N_25232,N_25070);
nor U25761 (N_25761,N_25184,N_25219);
xor U25762 (N_25762,N_25395,N_25181);
nand U25763 (N_25763,N_25018,N_25161);
nor U25764 (N_25764,N_25152,N_25144);
xnor U25765 (N_25765,N_25120,N_25454);
and U25766 (N_25766,N_25001,N_25074);
and U25767 (N_25767,N_25303,N_25066);
nor U25768 (N_25768,N_25343,N_25094);
nand U25769 (N_25769,N_25420,N_25431);
or U25770 (N_25770,N_25018,N_25185);
and U25771 (N_25771,N_25124,N_25280);
xor U25772 (N_25772,N_25396,N_25388);
or U25773 (N_25773,N_25278,N_25117);
and U25774 (N_25774,N_25184,N_25409);
nand U25775 (N_25775,N_25260,N_25350);
nor U25776 (N_25776,N_25449,N_25186);
and U25777 (N_25777,N_25237,N_25445);
or U25778 (N_25778,N_25060,N_25203);
or U25779 (N_25779,N_25010,N_25249);
and U25780 (N_25780,N_25187,N_25497);
or U25781 (N_25781,N_25451,N_25000);
or U25782 (N_25782,N_25391,N_25431);
xnor U25783 (N_25783,N_25296,N_25248);
and U25784 (N_25784,N_25479,N_25483);
nor U25785 (N_25785,N_25433,N_25448);
and U25786 (N_25786,N_25096,N_25011);
nor U25787 (N_25787,N_25312,N_25360);
xor U25788 (N_25788,N_25179,N_25497);
xor U25789 (N_25789,N_25224,N_25024);
nor U25790 (N_25790,N_25443,N_25394);
nand U25791 (N_25791,N_25202,N_25171);
nand U25792 (N_25792,N_25370,N_25142);
nor U25793 (N_25793,N_25332,N_25473);
nand U25794 (N_25794,N_25379,N_25015);
nor U25795 (N_25795,N_25363,N_25439);
nand U25796 (N_25796,N_25186,N_25266);
nand U25797 (N_25797,N_25050,N_25385);
nand U25798 (N_25798,N_25310,N_25213);
and U25799 (N_25799,N_25200,N_25159);
nand U25800 (N_25800,N_25275,N_25210);
or U25801 (N_25801,N_25456,N_25351);
or U25802 (N_25802,N_25401,N_25174);
or U25803 (N_25803,N_25254,N_25105);
or U25804 (N_25804,N_25156,N_25418);
or U25805 (N_25805,N_25291,N_25265);
and U25806 (N_25806,N_25075,N_25124);
and U25807 (N_25807,N_25472,N_25387);
nor U25808 (N_25808,N_25122,N_25331);
xor U25809 (N_25809,N_25128,N_25389);
nand U25810 (N_25810,N_25380,N_25219);
nor U25811 (N_25811,N_25340,N_25437);
or U25812 (N_25812,N_25249,N_25357);
nor U25813 (N_25813,N_25085,N_25130);
and U25814 (N_25814,N_25351,N_25088);
or U25815 (N_25815,N_25377,N_25201);
nor U25816 (N_25816,N_25085,N_25496);
nand U25817 (N_25817,N_25089,N_25186);
xnor U25818 (N_25818,N_25334,N_25235);
and U25819 (N_25819,N_25273,N_25233);
or U25820 (N_25820,N_25069,N_25036);
and U25821 (N_25821,N_25450,N_25158);
and U25822 (N_25822,N_25177,N_25459);
or U25823 (N_25823,N_25187,N_25024);
or U25824 (N_25824,N_25474,N_25059);
and U25825 (N_25825,N_25404,N_25077);
nor U25826 (N_25826,N_25452,N_25331);
nand U25827 (N_25827,N_25330,N_25451);
and U25828 (N_25828,N_25269,N_25352);
or U25829 (N_25829,N_25231,N_25230);
xor U25830 (N_25830,N_25476,N_25210);
or U25831 (N_25831,N_25113,N_25068);
xnor U25832 (N_25832,N_25063,N_25409);
nor U25833 (N_25833,N_25453,N_25314);
nor U25834 (N_25834,N_25069,N_25291);
nand U25835 (N_25835,N_25271,N_25389);
or U25836 (N_25836,N_25305,N_25081);
and U25837 (N_25837,N_25014,N_25071);
nand U25838 (N_25838,N_25146,N_25428);
and U25839 (N_25839,N_25317,N_25103);
and U25840 (N_25840,N_25031,N_25178);
or U25841 (N_25841,N_25064,N_25374);
or U25842 (N_25842,N_25301,N_25451);
or U25843 (N_25843,N_25020,N_25164);
nor U25844 (N_25844,N_25112,N_25137);
nand U25845 (N_25845,N_25352,N_25146);
nor U25846 (N_25846,N_25225,N_25277);
nand U25847 (N_25847,N_25349,N_25016);
or U25848 (N_25848,N_25406,N_25321);
or U25849 (N_25849,N_25451,N_25236);
xnor U25850 (N_25850,N_25152,N_25260);
nor U25851 (N_25851,N_25215,N_25364);
and U25852 (N_25852,N_25020,N_25498);
or U25853 (N_25853,N_25495,N_25298);
nand U25854 (N_25854,N_25280,N_25456);
and U25855 (N_25855,N_25489,N_25495);
xnor U25856 (N_25856,N_25378,N_25123);
and U25857 (N_25857,N_25194,N_25253);
xor U25858 (N_25858,N_25308,N_25132);
nor U25859 (N_25859,N_25283,N_25148);
and U25860 (N_25860,N_25368,N_25467);
or U25861 (N_25861,N_25032,N_25130);
or U25862 (N_25862,N_25462,N_25098);
xor U25863 (N_25863,N_25349,N_25155);
nor U25864 (N_25864,N_25266,N_25095);
or U25865 (N_25865,N_25070,N_25137);
xor U25866 (N_25866,N_25275,N_25045);
nor U25867 (N_25867,N_25140,N_25272);
and U25868 (N_25868,N_25131,N_25368);
xnor U25869 (N_25869,N_25156,N_25020);
nor U25870 (N_25870,N_25075,N_25395);
and U25871 (N_25871,N_25188,N_25324);
or U25872 (N_25872,N_25378,N_25026);
and U25873 (N_25873,N_25273,N_25454);
xor U25874 (N_25874,N_25315,N_25122);
nand U25875 (N_25875,N_25441,N_25484);
xor U25876 (N_25876,N_25035,N_25228);
or U25877 (N_25877,N_25395,N_25153);
nor U25878 (N_25878,N_25206,N_25088);
xnor U25879 (N_25879,N_25402,N_25313);
nor U25880 (N_25880,N_25141,N_25401);
nor U25881 (N_25881,N_25106,N_25336);
and U25882 (N_25882,N_25339,N_25368);
nand U25883 (N_25883,N_25389,N_25054);
xnor U25884 (N_25884,N_25473,N_25069);
and U25885 (N_25885,N_25113,N_25258);
and U25886 (N_25886,N_25384,N_25209);
xnor U25887 (N_25887,N_25466,N_25267);
and U25888 (N_25888,N_25233,N_25011);
nand U25889 (N_25889,N_25029,N_25135);
xnor U25890 (N_25890,N_25194,N_25212);
nor U25891 (N_25891,N_25448,N_25007);
or U25892 (N_25892,N_25436,N_25246);
nor U25893 (N_25893,N_25321,N_25102);
nand U25894 (N_25894,N_25498,N_25281);
or U25895 (N_25895,N_25280,N_25033);
nor U25896 (N_25896,N_25174,N_25072);
xor U25897 (N_25897,N_25061,N_25337);
or U25898 (N_25898,N_25285,N_25268);
xnor U25899 (N_25899,N_25056,N_25139);
or U25900 (N_25900,N_25341,N_25231);
and U25901 (N_25901,N_25271,N_25127);
or U25902 (N_25902,N_25132,N_25466);
and U25903 (N_25903,N_25049,N_25289);
xor U25904 (N_25904,N_25224,N_25370);
nor U25905 (N_25905,N_25313,N_25077);
nand U25906 (N_25906,N_25101,N_25302);
or U25907 (N_25907,N_25449,N_25395);
or U25908 (N_25908,N_25248,N_25334);
nand U25909 (N_25909,N_25241,N_25337);
nand U25910 (N_25910,N_25056,N_25390);
xor U25911 (N_25911,N_25210,N_25055);
nand U25912 (N_25912,N_25314,N_25072);
nand U25913 (N_25913,N_25251,N_25154);
or U25914 (N_25914,N_25041,N_25094);
nand U25915 (N_25915,N_25128,N_25283);
or U25916 (N_25916,N_25220,N_25019);
nand U25917 (N_25917,N_25213,N_25159);
and U25918 (N_25918,N_25384,N_25319);
nand U25919 (N_25919,N_25342,N_25243);
and U25920 (N_25920,N_25104,N_25319);
nor U25921 (N_25921,N_25249,N_25175);
or U25922 (N_25922,N_25079,N_25026);
and U25923 (N_25923,N_25313,N_25099);
xor U25924 (N_25924,N_25258,N_25270);
and U25925 (N_25925,N_25452,N_25224);
or U25926 (N_25926,N_25084,N_25145);
xor U25927 (N_25927,N_25499,N_25281);
and U25928 (N_25928,N_25442,N_25152);
or U25929 (N_25929,N_25247,N_25275);
nand U25930 (N_25930,N_25492,N_25146);
or U25931 (N_25931,N_25300,N_25337);
or U25932 (N_25932,N_25321,N_25487);
nand U25933 (N_25933,N_25340,N_25337);
nor U25934 (N_25934,N_25003,N_25128);
and U25935 (N_25935,N_25430,N_25445);
nor U25936 (N_25936,N_25309,N_25390);
nand U25937 (N_25937,N_25167,N_25235);
xor U25938 (N_25938,N_25294,N_25269);
xnor U25939 (N_25939,N_25094,N_25434);
or U25940 (N_25940,N_25032,N_25298);
or U25941 (N_25941,N_25360,N_25019);
nand U25942 (N_25942,N_25463,N_25343);
or U25943 (N_25943,N_25096,N_25328);
nor U25944 (N_25944,N_25439,N_25021);
or U25945 (N_25945,N_25011,N_25494);
and U25946 (N_25946,N_25422,N_25079);
nor U25947 (N_25947,N_25498,N_25043);
and U25948 (N_25948,N_25001,N_25121);
and U25949 (N_25949,N_25066,N_25029);
nor U25950 (N_25950,N_25131,N_25296);
xnor U25951 (N_25951,N_25326,N_25127);
or U25952 (N_25952,N_25191,N_25030);
nand U25953 (N_25953,N_25324,N_25338);
xnor U25954 (N_25954,N_25384,N_25375);
or U25955 (N_25955,N_25409,N_25154);
and U25956 (N_25956,N_25064,N_25153);
or U25957 (N_25957,N_25273,N_25326);
nand U25958 (N_25958,N_25389,N_25286);
and U25959 (N_25959,N_25260,N_25406);
nand U25960 (N_25960,N_25226,N_25046);
xor U25961 (N_25961,N_25326,N_25113);
and U25962 (N_25962,N_25483,N_25302);
nor U25963 (N_25963,N_25465,N_25036);
and U25964 (N_25964,N_25323,N_25301);
xnor U25965 (N_25965,N_25206,N_25219);
nor U25966 (N_25966,N_25440,N_25349);
xor U25967 (N_25967,N_25109,N_25128);
nand U25968 (N_25968,N_25028,N_25041);
or U25969 (N_25969,N_25372,N_25425);
and U25970 (N_25970,N_25426,N_25017);
nand U25971 (N_25971,N_25411,N_25236);
xnor U25972 (N_25972,N_25332,N_25399);
nor U25973 (N_25973,N_25267,N_25231);
xnor U25974 (N_25974,N_25457,N_25283);
or U25975 (N_25975,N_25398,N_25025);
nor U25976 (N_25976,N_25257,N_25321);
or U25977 (N_25977,N_25237,N_25463);
xnor U25978 (N_25978,N_25384,N_25222);
xnor U25979 (N_25979,N_25099,N_25295);
or U25980 (N_25980,N_25453,N_25048);
or U25981 (N_25981,N_25223,N_25079);
and U25982 (N_25982,N_25194,N_25488);
or U25983 (N_25983,N_25171,N_25427);
xnor U25984 (N_25984,N_25253,N_25048);
or U25985 (N_25985,N_25406,N_25019);
or U25986 (N_25986,N_25313,N_25331);
or U25987 (N_25987,N_25145,N_25174);
or U25988 (N_25988,N_25065,N_25132);
nand U25989 (N_25989,N_25209,N_25177);
and U25990 (N_25990,N_25154,N_25377);
nand U25991 (N_25991,N_25001,N_25146);
xor U25992 (N_25992,N_25209,N_25127);
nand U25993 (N_25993,N_25331,N_25453);
or U25994 (N_25994,N_25058,N_25145);
xnor U25995 (N_25995,N_25462,N_25101);
nor U25996 (N_25996,N_25251,N_25439);
xnor U25997 (N_25997,N_25034,N_25417);
nand U25998 (N_25998,N_25338,N_25258);
nor U25999 (N_25999,N_25425,N_25375);
xor U26000 (N_26000,N_25798,N_25644);
nor U26001 (N_26001,N_25926,N_25646);
nor U26002 (N_26002,N_25595,N_25839);
xnor U26003 (N_26003,N_25596,N_25529);
and U26004 (N_26004,N_25904,N_25675);
or U26005 (N_26005,N_25815,N_25650);
xnor U26006 (N_26006,N_25516,N_25505);
or U26007 (N_26007,N_25671,N_25912);
nand U26008 (N_26008,N_25584,N_25860);
xor U26009 (N_26009,N_25531,N_25514);
and U26010 (N_26010,N_25820,N_25694);
or U26011 (N_26011,N_25852,N_25717);
nand U26012 (N_26012,N_25978,N_25826);
nand U26013 (N_26013,N_25939,N_25603);
xor U26014 (N_26014,N_25913,N_25897);
nand U26015 (N_26015,N_25631,N_25903);
nand U26016 (N_26016,N_25754,N_25512);
and U26017 (N_26017,N_25676,N_25742);
nand U26018 (N_26018,N_25550,N_25682);
nor U26019 (N_26019,N_25848,N_25506);
and U26020 (N_26020,N_25801,N_25991);
xnor U26021 (N_26021,N_25953,N_25870);
xor U26022 (N_26022,N_25916,N_25971);
or U26023 (N_26023,N_25645,N_25735);
or U26024 (N_26024,N_25950,N_25804);
xor U26025 (N_26025,N_25859,N_25936);
nand U26026 (N_26026,N_25655,N_25948);
nor U26027 (N_26027,N_25575,N_25522);
and U26028 (N_26028,N_25614,N_25768);
xor U26029 (N_26029,N_25715,N_25758);
or U26030 (N_26030,N_25841,N_25803);
and U26031 (N_26031,N_25554,N_25532);
nand U26032 (N_26032,N_25877,N_25980);
or U26033 (N_26033,N_25802,N_25538);
and U26034 (N_26034,N_25875,N_25564);
xor U26035 (N_26035,N_25502,N_25769);
or U26036 (N_26036,N_25995,N_25500);
nand U26037 (N_26037,N_25880,N_25785);
nand U26038 (N_26038,N_25581,N_25790);
nand U26039 (N_26039,N_25600,N_25610);
or U26040 (N_26040,N_25873,N_25965);
nand U26041 (N_26041,N_25632,N_25621);
or U26042 (N_26042,N_25606,N_25961);
nand U26043 (N_26043,N_25780,N_25837);
and U26044 (N_26044,N_25602,N_25823);
or U26045 (N_26045,N_25756,N_25917);
and U26046 (N_26046,N_25541,N_25836);
nor U26047 (N_26047,N_25952,N_25762);
nor U26048 (N_26048,N_25734,N_25871);
and U26049 (N_26049,N_25716,N_25844);
xor U26050 (N_26050,N_25507,N_25892);
nand U26051 (N_26051,N_25623,N_25583);
and U26052 (N_26052,N_25821,N_25570);
xnor U26053 (N_26053,N_25729,N_25993);
nor U26054 (N_26054,N_25558,N_25647);
or U26055 (N_26055,N_25775,N_25774);
nor U26056 (N_26056,N_25789,N_25966);
xnor U26057 (N_26057,N_25984,N_25910);
nand U26058 (N_26058,N_25914,N_25868);
nand U26059 (N_26059,N_25518,N_25555);
nand U26060 (N_26060,N_25767,N_25686);
and U26061 (N_26061,N_25963,N_25891);
xnor U26062 (N_26062,N_25760,N_25510);
and U26063 (N_26063,N_25743,N_25695);
and U26064 (N_26064,N_25799,N_25628);
nor U26065 (N_26065,N_25778,N_25863);
nor U26066 (N_26066,N_25572,N_25582);
or U26067 (N_26067,N_25562,N_25976);
and U26068 (N_26068,N_25761,N_25730);
nand U26069 (N_26069,N_25755,N_25824);
xnor U26070 (N_26070,N_25657,N_25659);
nand U26071 (N_26071,N_25784,N_25713);
and U26072 (N_26072,N_25559,N_25683);
and U26073 (N_26073,N_25578,N_25690);
nor U26074 (N_26074,N_25940,N_25818);
nand U26075 (N_26075,N_25704,N_25827);
nor U26076 (N_26076,N_25731,N_25857);
nand U26077 (N_26077,N_25988,N_25751);
nand U26078 (N_26078,N_25997,N_25604);
and U26079 (N_26079,N_25535,N_25864);
nor U26080 (N_26080,N_25893,N_25673);
and U26081 (N_26081,N_25783,N_25526);
or U26082 (N_26082,N_25616,N_25981);
xnor U26083 (N_26083,N_25739,N_25782);
xor U26084 (N_26084,N_25560,N_25662);
xor U26085 (N_26085,N_25781,N_25901);
or U26086 (N_26086,N_25688,N_25908);
and U26087 (N_26087,N_25511,N_25585);
and U26088 (N_26088,N_25525,N_25958);
or U26089 (N_26089,N_25915,N_25771);
nand U26090 (N_26090,N_25987,N_25850);
nor U26091 (N_26091,N_25548,N_25626);
and U26092 (N_26092,N_25501,N_25816);
nor U26093 (N_26093,N_25598,N_25708);
xnor U26094 (N_26094,N_25979,N_25990);
and U26095 (N_26095,N_25625,N_25931);
and U26096 (N_26096,N_25527,N_25546);
xnor U26097 (N_26097,N_25609,N_25925);
nand U26098 (N_26098,N_25842,N_25504);
xnor U26099 (N_26099,N_25545,N_25797);
nand U26100 (N_26100,N_25949,N_25831);
nand U26101 (N_26101,N_25668,N_25664);
nor U26102 (N_26102,N_25744,N_25918);
or U26103 (N_26103,N_25720,N_25938);
xnor U26104 (N_26104,N_25854,N_25661);
or U26105 (N_26105,N_25772,N_25919);
nor U26106 (N_26106,N_25969,N_25568);
or U26107 (N_26107,N_25763,N_25648);
nor U26108 (N_26108,N_25843,N_25725);
and U26109 (N_26109,N_25660,N_25951);
and U26110 (N_26110,N_25773,N_25736);
xor U26111 (N_26111,N_25537,N_25569);
and U26112 (N_26112,N_25520,N_25999);
nor U26113 (N_26113,N_25796,N_25653);
nor U26114 (N_26114,N_25835,N_25513);
and U26115 (N_26115,N_25874,N_25989);
and U26116 (N_26116,N_25779,N_25574);
xor U26117 (N_26117,N_25576,N_25975);
and U26118 (N_26118,N_25639,N_25866);
or U26119 (N_26119,N_25884,N_25807);
or U26120 (N_26120,N_25861,N_25776);
nor U26121 (N_26121,N_25705,N_25737);
nand U26122 (N_26122,N_25895,N_25882);
nand U26123 (N_26123,N_25642,N_25964);
nand U26124 (N_26124,N_25552,N_25654);
xor U26125 (N_26125,N_25928,N_25613);
nor U26126 (N_26126,N_25937,N_25753);
or U26127 (N_26127,N_25996,N_25846);
and U26128 (N_26128,N_25845,N_25832);
and U26129 (N_26129,N_25956,N_25945);
nand U26130 (N_26130,N_25898,N_25929);
nand U26131 (N_26131,N_25721,N_25765);
and U26132 (N_26132,N_25921,N_25643);
xor U26133 (N_26133,N_25542,N_25651);
or U26134 (N_26134,N_25543,N_25817);
nand U26135 (N_26135,N_25573,N_25687);
or U26136 (N_26136,N_25508,N_25791);
or U26137 (N_26137,N_25896,N_25795);
and U26138 (N_26138,N_25732,N_25786);
nand U26139 (N_26139,N_25906,N_25800);
nand U26140 (N_26140,N_25698,N_25867);
nand U26141 (N_26141,N_25833,N_25923);
or U26142 (N_26142,N_25813,N_25794);
xnor U26143 (N_26143,N_25515,N_25630);
and U26144 (N_26144,N_25986,N_25567);
nand U26145 (N_26145,N_25615,N_25766);
nor U26146 (N_26146,N_25959,N_25770);
nand U26147 (N_26147,N_25930,N_25649);
or U26148 (N_26148,N_25551,N_25556);
and U26149 (N_26149,N_25530,N_25656);
nor U26150 (N_26150,N_25828,N_25983);
and U26151 (N_26151,N_25962,N_25876);
and U26152 (N_26152,N_25968,N_25670);
nor U26153 (N_26153,N_25722,N_25883);
nor U26154 (N_26154,N_25738,N_25911);
and U26155 (N_26155,N_25881,N_25580);
or U26156 (N_26156,N_25973,N_25565);
and U26157 (N_26157,N_25579,N_25701);
and U26158 (N_26158,N_25932,N_25809);
nor U26159 (N_26159,N_25679,N_25922);
and U26160 (N_26160,N_25849,N_25719);
nor U26161 (N_26161,N_25669,N_25697);
and U26162 (N_26162,N_25622,N_25985);
and U26163 (N_26163,N_25703,N_25748);
xnor U26164 (N_26164,N_25752,N_25637);
xor U26165 (N_26165,N_25955,N_25636);
or U26166 (N_26166,N_25710,N_25706);
or U26167 (N_26167,N_25992,N_25601);
nor U26168 (N_26168,N_25718,N_25788);
nor U26169 (N_26169,N_25693,N_25692);
nand U26170 (N_26170,N_25733,N_25812);
nand U26171 (N_26171,N_25757,N_25792);
and U26172 (N_26172,N_25519,N_25685);
or U26173 (N_26173,N_25829,N_25900);
or U26174 (N_26174,N_25960,N_25635);
nor U26175 (N_26175,N_25509,N_25633);
nor U26176 (N_26176,N_25855,N_25547);
nor U26177 (N_26177,N_25764,N_25561);
and U26178 (N_26178,N_25957,N_25699);
xor U26179 (N_26179,N_25994,N_25618);
nor U26180 (N_26180,N_25889,N_25702);
and U26181 (N_26181,N_25521,N_25640);
and U26182 (N_26182,N_25907,N_25599);
xor U26183 (N_26183,N_25680,N_25593);
xor U26184 (N_26184,N_25941,N_25566);
or U26185 (N_26185,N_25712,N_25681);
or U26186 (N_26186,N_25641,N_25726);
nor U26187 (N_26187,N_25665,N_25629);
nand U26188 (N_26188,N_25549,N_25970);
or U26189 (N_26189,N_25819,N_25747);
and U26190 (N_26190,N_25862,N_25577);
nand U26191 (N_26191,N_25607,N_25878);
or U26192 (N_26192,N_25974,N_25724);
or U26193 (N_26193,N_25793,N_25856);
xor U26194 (N_26194,N_25700,N_25838);
xnor U26195 (N_26195,N_25967,N_25617);
nor U26196 (N_26196,N_25759,N_25777);
xnor U26197 (N_26197,N_25749,N_25811);
or U26198 (N_26198,N_25840,N_25553);
nor U26199 (N_26199,N_25540,N_25887);
nand U26200 (N_26200,N_25740,N_25954);
nor U26201 (N_26201,N_25587,N_25658);
nand U26202 (N_26202,N_25944,N_25707);
nand U26203 (N_26203,N_25746,N_25528);
nor U26204 (N_26204,N_25689,N_25638);
xnor U26205 (N_26205,N_25869,N_25533);
or U26206 (N_26206,N_25709,N_25851);
and U26207 (N_26207,N_25674,N_25691);
xor U26208 (N_26208,N_25666,N_25608);
nand U26209 (N_26209,N_25563,N_25590);
nor U26210 (N_26210,N_25594,N_25998);
or U26211 (N_26211,N_25899,N_25909);
nor U26212 (N_26212,N_25741,N_25684);
xor U26213 (N_26213,N_25524,N_25627);
nor U26214 (N_26214,N_25830,N_25787);
and U26215 (N_26215,N_25677,N_25539);
and U26216 (N_26216,N_25678,N_25597);
nor U26217 (N_26217,N_25853,N_25591);
nor U26218 (N_26218,N_25605,N_25806);
xnor U26219 (N_26219,N_25624,N_25972);
or U26220 (N_26220,N_25544,N_25750);
nand U26221 (N_26221,N_25652,N_25611);
or U26222 (N_26222,N_25696,N_25727);
or U26223 (N_26223,N_25589,N_25942);
xnor U26224 (N_26224,N_25503,N_25586);
xnor U26225 (N_26225,N_25612,N_25517);
nand U26226 (N_26226,N_25920,N_25805);
and U26227 (N_26227,N_25934,N_25534);
nor U26228 (N_26228,N_25933,N_25865);
xnor U26229 (N_26229,N_25523,N_25847);
and U26230 (N_26230,N_25634,N_25834);
nand U26231 (N_26231,N_25822,N_25808);
nor U26232 (N_26232,N_25888,N_25714);
and U26233 (N_26233,N_25723,N_25943);
or U26234 (N_26234,N_25872,N_25745);
nor U26235 (N_26235,N_25588,N_25894);
or U26236 (N_26236,N_25902,N_25924);
or U26237 (N_26237,N_25890,N_25982);
or U26238 (N_26238,N_25879,N_25571);
nor U26239 (N_26239,N_25927,N_25592);
xor U26240 (N_26240,N_25886,N_25667);
and U26241 (N_26241,N_25935,N_25728);
nand U26242 (N_26242,N_25557,N_25858);
xnor U26243 (N_26243,N_25977,N_25672);
nand U26244 (N_26244,N_25885,N_25536);
or U26245 (N_26245,N_25825,N_25620);
nor U26246 (N_26246,N_25905,N_25810);
nor U26247 (N_26247,N_25619,N_25663);
and U26248 (N_26248,N_25946,N_25947);
and U26249 (N_26249,N_25814,N_25711);
nand U26250 (N_26250,N_25923,N_25609);
and U26251 (N_26251,N_25844,N_25929);
nor U26252 (N_26252,N_25971,N_25813);
nand U26253 (N_26253,N_25697,N_25549);
nor U26254 (N_26254,N_25513,N_25788);
xor U26255 (N_26255,N_25642,N_25532);
and U26256 (N_26256,N_25860,N_25835);
nor U26257 (N_26257,N_25791,N_25586);
or U26258 (N_26258,N_25548,N_25722);
nand U26259 (N_26259,N_25650,N_25691);
xnor U26260 (N_26260,N_25863,N_25880);
and U26261 (N_26261,N_25988,N_25506);
xnor U26262 (N_26262,N_25963,N_25974);
nor U26263 (N_26263,N_25740,N_25794);
nor U26264 (N_26264,N_25747,N_25504);
and U26265 (N_26265,N_25766,N_25812);
xnor U26266 (N_26266,N_25987,N_25513);
nand U26267 (N_26267,N_25879,N_25659);
and U26268 (N_26268,N_25977,N_25945);
or U26269 (N_26269,N_25503,N_25950);
nor U26270 (N_26270,N_25696,N_25818);
xnor U26271 (N_26271,N_25881,N_25699);
and U26272 (N_26272,N_25839,N_25721);
nor U26273 (N_26273,N_25882,N_25845);
or U26274 (N_26274,N_25712,N_25579);
xor U26275 (N_26275,N_25618,N_25563);
and U26276 (N_26276,N_25708,N_25691);
nor U26277 (N_26277,N_25712,N_25853);
nor U26278 (N_26278,N_25936,N_25955);
or U26279 (N_26279,N_25648,N_25754);
or U26280 (N_26280,N_25532,N_25557);
or U26281 (N_26281,N_25561,N_25822);
nand U26282 (N_26282,N_25952,N_25677);
and U26283 (N_26283,N_25564,N_25578);
nor U26284 (N_26284,N_25710,N_25889);
or U26285 (N_26285,N_25616,N_25733);
and U26286 (N_26286,N_25609,N_25533);
xor U26287 (N_26287,N_25637,N_25516);
or U26288 (N_26288,N_25819,N_25840);
nand U26289 (N_26289,N_25881,N_25563);
and U26290 (N_26290,N_25618,N_25650);
xnor U26291 (N_26291,N_25671,N_25945);
and U26292 (N_26292,N_25903,N_25699);
xor U26293 (N_26293,N_25623,N_25807);
xnor U26294 (N_26294,N_25789,N_25588);
nor U26295 (N_26295,N_25580,N_25672);
nand U26296 (N_26296,N_25954,N_25854);
and U26297 (N_26297,N_25880,N_25653);
or U26298 (N_26298,N_25960,N_25850);
nor U26299 (N_26299,N_25997,N_25627);
nor U26300 (N_26300,N_25734,N_25528);
or U26301 (N_26301,N_25914,N_25880);
nand U26302 (N_26302,N_25838,N_25745);
nand U26303 (N_26303,N_25805,N_25574);
or U26304 (N_26304,N_25602,N_25582);
xor U26305 (N_26305,N_25814,N_25532);
xor U26306 (N_26306,N_25885,N_25916);
nand U26307 (N_26307,N_25673,N_25628);
nor U26308 (N_26308,N_25858,N_25914);
nand U26309 (N_26309,N_25522,N_25946);
or U26310 (N_26310,N_25984,N_25827);
and U26311 (N_26311,N_25545,N_25896);
xnor U26312 (N_26312,N_25916,N_25636);
or U26313 (N_26313,N_25814,N_25713);
and U26314 (N_26314,N_25808,N_25512);
nor U26315 (N_26315,N_25880,N_25576);
and U26316 (N_26316,N_25875,N_25924);
and U26317 (N_26317,N_25658,N_25991);
and U26318 (N_26318,N_25698,N_25838);
and U26319 (N_26319,N_25917,N_25531);
or U26320 (N_26320,N_25839,N_25803);
xnor U26321 (N_26321,N_25920,N_25636);
nand U26322 (N_26322,N_25964,N_25593);
or U26323 (N_26323,N_25675,N_25526);
and U26324 (N_26324,N_25532,N_25759);
nor U26325 (N_26325,N_25960,N_25697);
or U26326 (N_26326,N_25908,N_25965);
nand U26327 (N_26327,N_25529,N_25569);
xor U26328 (N_26328,N_25819,N_25760);
nor U26329 (N_26329,N_25816,N_25857);
nand U26330 (N_26330,N_25871,N_25830);
or U26331 (N_26331,N_25718,N_25853);
and U26332 (N_26332,N_25787,N_25568);
and U26333 (N_26333,N_25710,N_25829);
nand U26334 (N_26334,N_25527,N_25522);
nand U26335 (N_26335,N_25612,N_25645);
xnor U26336 (N_26336,N_25950,N_25852);
xor U26337 (N_26337,N_25644,N_25675);
and U26338 (N_26338,N_25555,N_25661);
nand U26339 (N_26339,N_25913,N_25579);
nor U26340 (N_26340,N_25843,N_25560);
nor U26341 (N_26341,N_25956,N_25768);
xor U26342 (N_26342,N_25807,N_25600);
xnor U26343 (N_26343,N_25635,N_25592);
nand U26344 (N_26344,N_25519,N_25892);
xnor U26345 (N_26345,N_25560,N_25654);
nand U26346 (N_26346,N_25613,N_25883);
nand U26347 (N_26347,N_25965,N_25713);
and U26348 (N_26348,N_25985,N_25884);
and U26349 (N_26349,N_25525,N_25821);
nor U26350 (N_26350,N_25989,N_25793);
xor U26351 (N_26351,N_25670,N_25938);
nand U26352 (N_26352,N_25929,N_25749);
or U26353 (N_26353,N_25689,N_25634);
or U26354 (N_26354,N_25680,N_25932);
xor U26355 (N_26355,N_25849,N_25571);
nor U26356 (N_26356,N_25729,N_25574);
nand U26357 (N_26357,N_25552,N_25517);
and U26358 (N_26358,N_25570,N_25689);
nand U26359 (N_26359,N_25606,N_25747);
nor U26360 (N_26360,N_25572,N_25875);
nand U26361 (N_26361,N_25681,N_25984);
or U26362 (N_26362,N_25869,N_25722);
or U26363 (N_26363,N_25516,N_25924);
or U26364 (N_26364,N_25645,N_25861);
xnor U26365 (N_26365,N_25583,N_25541);
nand U26366 (N_26366,N_25551,N_25717);
xor U26367 (N_26367,N_25995,N_25988);
and U26368 (N_26368,N_25860,N_25768);
nor U26369 (N_26369,N_25595,N_25867);
nand U26370 (N_26370,N_25667,N_25757);
nand U26371 (N_26371,N_25907,N_25673);
xor U26372 (N_26372,N_25664,N_25737);
nand U26373 (N_26373,N_25766,N_25664);
nand U26374 (N_26374,N_25679,N_25645);
and U26375 (N_26375,N_25690,N_25943);
nand U26376 (N_26376,N_25772,N_25899);
nand U26377 (N_26377,N_25790,N_25511);
nor U26378 (N_26378,N_25972,N_25833);
and U26379 (N_26379,N_25564,N_25607);
xnor U26380 (N_26380,N_25642,N_25999);
and U26381 (N_26381,N_25811,N_25724);
xnor U26382 (N_26382,N_25689,N_25900);
and U26383 (N_26383,N_25708,N_25819);
nor U26384 (N_26384,N_25770,N_25877);
nor U26385 (N_26385,N_25643,N_25905);
nor U26386 (N_26386,N_25639,N_25992);
nand U26387 (N_26387,N_25907,N_25672);
or U26388 (N_26388,N_25531,N_25869);
nand U26389 (N_26389,N_25958,N_25770);
or U26390 (N_26390,N_25915,N_25504);
and U26391 (N_26391,N_25758,N_25683);
and U26392 (N_26392,N_25944,N_25718);
nor U26393 (N_26393,N_25865,N_25925);
nand U26394 (N_26394,N_25515,N_25703);
nand U26395 (N_26395,N_25928,N_25547);
xnor U26396 (N_26396,N_25771,N_25769);
xor U26397 (N_26397,N_25886,N_25706);
or U26398 (N_26398,N_25841,N_25901);
nand U26399 (N_26399,N_25630,N_25876);
nand U26400 (N_26400,N_25722,N_25601);
nand U26401 (N_26401,N_25778,N_25966);
or U26402 (N_26402,N_25523,N_25774);
nand U26403 (N_26403,N_25766,N_25833);
xor U26404 (N_26404,N_25772,N_25924);
nor U26405 (N_26405,N_25899,N_25643);
xnor U26406 (N_26406,N_25745,N_25821);
and U26407 (N_26407,N_25915,N_25847);
and U26408 (N_26408,N_25956,N_25767);
and U26409 (N_26409,N_25593,N_25951);
nor U26410 (N_26410,N_25668,N_25595);
or U26411 (N_26411,N_25955,N_25767);
xnor U26412 (N_26412,N_25887,N_25781);
xor U26413 (N_26413,N_25931,N_25520);
and U26414 (N_26414,N_25565,N_25531);
xor U26415 (N_26415,N_25594,N_25673);
or U26416 (N_26416,N_25896,N_25603);
xor U26417 (N_26417,N_25673,N_25993);
nor U26418 (N_26418,N_25756,N_25786);
xor U26419 (N_26419,N_25570,N_25682);
nand U26420 (N_26420,N_25962,N_25709);
nand U26421 (N_26421,N_25938,N_25936);
or U26422 (N_26422,N_25716,N_25561);
nand U26423 (N_26423,N_25691,N_25509);
xor U26424 (N_26424,N_25802,N_25693);
or U26425 (N_26425,N_25974,N_25981);
and U26426 (N_26426,N_25814,N_25561);
nor U26427 (N_26427,N_25589,N_25654);
or U26428 (N_26428,N_25710,N_25678);
xor U26429 (N_26429,N_25610,N_25915);
or U26430 (N_26430,N_25536,N_25687);
nor U26431 (N_26431,N_25946,N_25909);
nand U26432 (N_26432,N_25976,N_25928);
and U26433 (N_26433,N_25959,N_25697);
nor U26434 (N_26434,N_25531,N_25606);
nor U26435 (N_26435,N_25571,N_25585);
xor U26436 (N_26436,N_25689,N_25844);
nor U26437 (N_26437,N_25897,N_25628);
or U26438 (N_26438,N_25681,N_25512);
or U26439 (N_26439,N_25885,N_25713);
xor U26440 (N_26440,N_25910,N_25666);
or U26441 (N_26441,N_25754,N_25681);
or U26442 (N_26442,N_25915,N_25816);
nor U26443 (N_26443,N_25524,N_25992);
nor U26444 (N_26444,N_25907,N_25975);
or U26445 (N_26445,N_25746,N_25520);
nand U26446 (N_26446,N_25938,N_25859);
nor U26447 (N_26447,N_25765,N_25972);
and U26448 (N_26448,N_25669,N_25915);
or U26449 (N_26449,N_25929,N_25916);
or U26450 (N_26450,N_25523,N_25865);
or U26451 (N_26451,N_25762,N_25916);
or U26452 (N_26452,N_25610,N_25980);
nand U26453 (N_26453,N_25881,N_25833);
xnor U26454 (N_26454,N_25838,N_25515);
nor U26455 (N_26455,N_25813,N_25809);
nor U26456 (N_26456,N_25610,N_25602);
or U26457 (N_26457,N_25969,N_25664);
or U26458 (N_26458,N_25811,N_25785);
nand U26459 (N_26459,N_25759,N_25853);
xnor U26460 (N_26460,N_25725,N_25962);
and U26461 (N_26461,N_25510,N_25556);
xor U26462 (N_26462,N_25651,N_25532);
xnor U26463 (N_26463,N_25619,N_25873);
nor U26464 (N_26464,N_25904,N_25687);
nor U26465 (N_26465,N_25949,N_25879);
nor U26466 (N_26466,N_25983,N_25934);
and U26467 (N_26467,N_25822,N_25547);
and U26468 (N_26468,N_25753,N_25903);
nand U26469 (N_26469,N_25581,N_25799);
nand U26470 (N_26470,N_25816,N_25656);
and U26471 (N_26471,N_25724,N_25503);
and U26472 (N_26472,N_25800,N_25805);
and U26473 (N_26473,N_25635,N_25937);
or U26474 (N_26474,N_25514,N_25846);
nand U26475 (N_26475,N_25812,N_25856);
nand U26476 (N_26476,N_25581,N_25849);
nor U26477 (N_26477,N_25805,N_25615);
or U26478 (N_26478,N_25817,N_25902);
nor U26479 (N_26479,N_25590,N_25649);
or U26480 (N_26480,N_25800,N_25680);
and U26481 (N_26481,N_25519,N_25840);
or U26482 (N_26482,N_25986,N_25886);
and U26483 (N_26483,N_25789,N_25660);
nand U26484 (N_26484,N_25637,N_25717);
nand U26485 (N_26485,N_25614,N_25833);
nand U26486 (N_26486,N_25888,N_25661);
nor U26487 (N_26487,N_25928,N_25610);
or U26488 (N_26488,N_25984,N_25518);
xnor U26489 (N_26489,N_25729,N_25504);
and U26490 (N_26490,N_25966,N_25611);
xor U26491 (N_26491,N_25725,N_25923);
or U26492 (N_26492,N_25913,N_25862);
nor U26493 (N_26493,N_25588,N_25767);
xor U26494 (N_26494,N_25766,N_25986);
xor U26495 (N_26495,N_25561,N_25808);
nor U26496 (N_26496,N_25760,N_25752);
or U26497 (N_26497,N_25545,N_25565);
nor U26498 (N_26498,N_25963,N_25576);
nand U26499 (N_26499,N_25629,N_25810);
nor U26500 (N_26500,N_26388,N_26441);
and U26501 (N_26501,N_26078,N_26019);
nand U26502 (N_26502,N_26090,N_26207);
xnor U26503 (N_26503,N_26270,N_26381);
nor U26504 (N_26504,N_26389,N_26427);
and U26505 (N_26505,N_26179,N_26260);
xnor U26506 (N_26506,N_26176,N_26481);
nand U26507 (N_26507,N_26408,N_26340);
nand U26508 (N_26508,N_26014,N_26295);
and U26509 (N_26509,N_26470,N_26405);
nand U26510 (N_26510,N_26048,N_26466);
or U26511 (N_26511,N_26069,N_26232);
or U26512 (N_26512,N_26430,N_26010);
nand U26513 (N_26513,N_26290,N_26031);
and U26514 (N_26514,N_26462,N_26171);
xor U26515 (N_26515,N_26442,N_26224);
or U26516 (N_26516,N_26001,N_26355);
nand U26517 (N_26517,N_26140,N_26184);
nand U26518 (N_26518,N_26280,N_26017);
nand U26519 (N_26519,N_26312,N_26372);
and U26520 (N_26520,N_26066,N_26020);
nor U26521 (N_26521,N_26465,N_26170);
xor U26522 (N_26522,N_26160,N_26122);
xnor U26523 (N_26523,N_26114,N_26229);
xor U26524 (N_26524,N_26238,N_26094);
nor U26525 (N_26525,N_26086,N_26198);
nand U26526 (N_26526,N_26040,N_26366);
and U26527 (N_26527,N_26080,N_26436);
or U26528 (N_26528,N_26460,N_26100);
nor U26529 (N_26529,N_26396,N_26415);
and U26530 (N_26530,N_26189,N_26126);
xor U26531 (N_26531,N_26474,N_26104);
nand U26532 (N_26532,N_26488,N_26044);
nand U26533 (N_26533,N_26392,N_26226);
nand U26534 (N_26534,N_26306,N_26116);
and U26535 (N_26535,N_26391,N_26130);
or U26536 (N_26536,N_26360,N_26275);
xor U26537 (N_26537,N_26028,N_26320);
and U26538 (N_26538,N_26431,N_26233);
nor U26539 (N_26539,N_26099,N_26012);
and U26540 (N_26540,N_26065,N_26083);
or U26541 (N_26541,N_26487,N_26315);
nor U26542 (N_26542,N_26254,N_26305);
nor U26543 (N_26543,N_26288,N_26060);
or U26544 (N_26544,N_26006,N_26303);
and U26545 (N_26545,N_26287,N_26241);
xnor U26546 (N_26546,N_26084,N_26380);
xor U26547 (N_26547,N_26110,N_26141);
xnor U26548 (N_26548,N_26301,N_26369);
nand U26549 (N_26549,N_26145,N_26429);
nand U26550 (N_26550,N_26418,N_26218);
nor U26551 (N_26551,N_26188,N_26491);
nor U26552 (N_26552,N_26117,N_26333);
nand U26553 (N_26553,N_26399,N_26349);
xnor U26554 (N_26554,N_26225,N_26223);
and U26555 (N_26555,N_26367,N_26265);
and U26556 (N_26556,N_26385,N_26482);
nor U26557 (N_26557,N_26216,N_26063);
xnor U26558 (N_26558,N_26456,N_26345);
xor U26559 (N_26559,N_26322,N_26486);
nor U26560 (N_26560,N_26298,N_26330);
nor U26561 (N_26561,N_26492,N_26029);
or U26562 (N_26562,N_26213,N_26237);
xnor U26563 (N_26563,N_26095,N_26251);
and U26564 (N_26564,N_26489,N_26119);
or U26565 (N_26565,N_26464,N_26495);
and U26566 (N_26566,N_26473,N_26284);
xor U26567 (N_26567,N_26037,N_26416);
and U26568 (N_26568,N_26304,N_26432);
xnor U26569 (N_26569,N_26476,N_26445);
and U26570 (N_26570,N_26199,N_26309);
nor U26571 (N_26571,N_26267,N_26478);
or U26572 (N_26572,N_26249,N_26153);
xnor U26573 (N_26573,N_26087,N_26068);
nor U26574 (N_26574,N_26274,N_26386);
nor U26575 (N_26575,N_26376,N_26371);
nand U26576 (N_26576,N_26440,N_26053);
and U26577 (N_26577,N_26258,N_26294);
and U26578 (N_26578,N_26455,N_26361);
or U26579 (N_26579,N_26246,N_26434);
xnor U26580 (N_26580,N_26424,N_26142);
nand U26581 (N_26581,N_26348,N_26013);
or U26582 (N_26582,N_26394,N_26051);
nand U26583 (N_26583,N_26273,N_26124);
or U26584 (N_26584,N_26458,N_26278);
and U26585 (N_26585,N_26190,N_26056);
and U26586 (N_26586,N_26036,N_26477);
or U26587 (N_26587,N_26469,N_26209);
xnor U26588 (N_26588,N_26039,N_26230);
nand U26589 (N_26589,N_26005,N_26148);
and U26590 (N_26590,N_26067,N_26313);
and U26591 (N_26591,N_26096,N_26475);
or U26592 (N_26592,N_26335,N_26490);
and U26593 (N_26593,N_26472,N_26336);
nand U26594 (N_26594,N_26215,N_26368);
and U26595 (N_26595,N_26195,N_26422);
nor U26596 (N_26596,N_26410,N_26387);
nor U26597 (N_26597,N_26158,N_26159);
xor U26598 (N_26598,N_26334,N_26297);
and U26599 (N_26599,N_26054,N_26314);
nand U26600 (N_26600,N_26281,N_26098);
nor U26601 (N_26601,N_26057,N_26454);
nor U26602 (N_26602,N_26205,N_26425);
nor U26603 (N_26603,N_26459,N_26292);
or U26604 (N_26604,N_26191,N_26093);
nand U26605 (N_26605,N_26018,N_26131);
and U26606 (N_26606,N_26463,N_26296);
nor U26607 (N_26607,N_26112,N_26026);
or U26608 (N_26608,N_26252,N_26354);
and U26609 (N_26609,N_26062,N_26497);
and U26610 (N_26610,N_26344,N_26253);
and U26611 (N_26611,N_26185,N_26438);
xor U26612 (N_26612,N_26412,N_26151);
nand U26613 (N_26613,N_26339,N_26433);
nor U26614 (N_26614,N_26435,N_26332);
or U26615 (N_26615,N_26496,N_26137);
nand U26616 (N_26616,N_26164,N_26206);
and U26617 (N_26617,N_26318,N_26033);
xnor U26618 (N_26618,N_26042,N_26419);
and U26619 (N_26619,N_26310,N_26045);
and U26620 (N_26620,N_26308,N_26139);
and U26621 (N_26621,N_26214,N_26004);
nand U26622 (N_26622,N_26453,N_26446);
xor U26623 (N_26623,N_26328,N_26220);
or U26624 (N_26624,N_26072,N_26420);
nand U26625 (N_26625,N_26135,N_26269);
xnor U26626 (N_26626,N_26437,N_26245);
or U26627 (N_26627,N_26201,N_26228);
or U26628 (N_26628,N_26406,N_26485);
xnor U26629 (N_26629,N_26319,N_26413);
nor U26630 (N_26630,N_26421,N_26426);
xor U26631 (N_26631,N_26043,N_26082);
nand U26632 (N_26632,N_26146,N_26250);
xor U26633 (N_26633,N_26293,N_26107);
nor U26634 (N_26634,N_26374,N_26091);
or U26635 (N_26635,N_26038,N_26011);
or U26636 (N_26636,N_26341,N_26167);
or U26637 (N_26637,N_26248,N_26147);
or U26638 (N_26638,N_26353,N_26144);
or U26639 (N_26639,N_26452,N_26257);
or U26640 (N_26640,N_26120,N_26172);
and U26641 (N_26641,N_26217,N_26326);
nor U26642 (N_26642,N_26134,N_26236);
or U26643 (N_26643,N_26390,N_26003);
or U26644 (N_26644,N_26202,N_26261);
nand U26645 (N_26645,N_26168,N_26000);
or U26646 (N_26646,N_26115,N_26423);
xnor U26647 (N_26647,N_26210,N_26102);
xnor U26648 (N_26648,N_26041,N_26384);
xor U26649 (N_26649,N_26174,N_26483);
xnor U26650 (N_26650,N_26383,N_26109);
and U26651 (N_26651,N_26443,N_26157);
xor U26652 (N_26652,N_26307,N_26331);
nand U26653 (N_26653,N_26279,N_26365);
nor U26654 (N_26654,N_26357,N_26049);
or U26655 (N_26655,N_26125,N_26363);
and U26656 (N_26656,N_26276,N_26402);
nor U26657 (N_26657,N_26343,N_26370);
nor U26658 (N_26658,N_26149,N_26272);
xnor U26659 (N_26659,N_26092,N_26059);
and U26660 (N_26660,N_26193,N_26359);
or U26661 (N_26661,N_26074,N_26030);
xnor U26662 (N_26662,N_26085,N_26187);
nand U26663 (N_26663,N_26327,N_26259);
xor U26664 (N_26664,N_26009,N_26398);
nand U26665 (N_26665,N_26178,N_26373);
nand U26666 (N_26666,N_26375,N_26052);
nor U26667 (N_26667,N_26282,N_26152);
and U26668 (N_26668,N_26173,N_26351);
nand U26669 (N_26669,N_26311,N_26242);
xnor U26670 (N_26670,N_26212,N_26493);
nor U26671 (N_26671,N_26499,N_26071);
nand U26672 (N_26672,N_26032,N_26204);
and U26673 (N_26673,N_26123,N_26024);
xnor U26674 (N_26674,N_26034,N_26263);
and U26675 (N_26675,N_26317,N_26008);
and U26676 (N_26676,N_26227,N_26047);
and U26677 (N_26677,N_26108,N_26113);
and U26678 (N_26678,N_26180,N_26448);
nand U26679 (N_26679,N_26409,N_26457);
nand U26680 (N_26680,N_26155,N_26286);
and U26681 (N_26681,N_26471,N_26182);
nand U26682 (N_26682,N_26444,N_26132);
xor U26683 (N_26683,N_26285,N_26136);
xnor U26684 (N_26684,N_26244,N_26055);
and U26685 (N_26685,N_26329,N_26480);
and U26686 (N_26686,N_26479,N_26362);
or U26687 (N_26687,N_26299,N_26404);
nor U26688 (N_26688,N_26400,N_26411);
nand U26689 (N_26689,N_26243,N_26169);
and U26690 (N_26690,N_26323,N_26161);
nor U26691 (N_26691,N_26395,N_26143);
xor U26692 (N_26692,N_26118,N_26023);
or U26693 (N_26693,N_26358,N_26035);
nor U26694 (N_26694,N_26247,N_26468);
nor U26695 (N_26695,N_26088,N_26077);
xor U26696 (N_26696,N_26186,N_26264);
nand U26697 (N_26697,N_26061,N_26291);
xnor U26698 (N_26698,N_26181,N_26221);
nor U26699 (N_26699,N_26447,N_26200);
nor U26700 (N_26700,N_26165,N_26467);
nor U26701 (N_26701,N_26283,N_26075);
or U26702 (N_26702,N_26203,N_26002);
nor U26703 (N_26703,N_26271,N_26064);
nor U26704 (N_26704,N_26127,N_26166);
or U26705 (N_26705,N_26162,N_26154);
and U26706 (N_26706,N_26316,N_26106);
and U26707 (N_26707,N_26428,N_26050);
nor U26708 (N_26708,N_26255,N_26342);
and U26709 (N_26709,N_26407,N_26377);
nor U26710 (N_26710,N_26128,N_26121);
nor U26711 (N_26711,N_26081,N_26403);
or U26712 (N_26712,N_26133,N_26022);
nor U26713 (N_26713,N_26222,N_26058);
nor U26714 (N_26714,N_26234,N_26382);
and U26715 (N_26715,N_26484,N_26240);
xnor U26716 (N_26716,N_26194,N_26076);
nand U26717 (N_26717,N_26239,N_26007);
xnor U26718 (N_26718,N_26070,N_26150);
nor U26719 (N_26719,N_26211,N_26325);
nor U26720 (N_26720,N_26256,N_26197);
xor U26721 (N_26721,N_26138,N_26111);
nor U26722 (N_26722,N_26262,N_26235);
or U26723 (N_26723,N_26101,N_26027);
or U26724 (N_26724,N_26208,N_26025);
nor U26725 (N_26725,N_26364,N_26451);
nor U26726 (N_26726,N_26089,N_26494);
or U26727 (N_26727,N_26417,N_26352);
and U26728 (N_26728,N_26129,N_26461);
or U26729 (N_26729,N_26175,N_26401);
nand U26730 (N_26730,N_26338,N_26397);
and U26731 (N_26731,N_26450,N_26156);
and U26732 (N_26732,N_26393,N_26219);
and U26733 (N_26733,N_26277,N_26015);
and U26734 (N_26734,N_26414,N_26346);
and U26735 (N_26735,N_26449,N_26300);
and U26736 (N_26736,N_26302,N_26021);
xnor U26737 (N_26737,N_26498,N_26289);
xnor U26738 (N_26738,N_26097,N_26073);
xnor U26739 (N_26739,N_26347,N_26016);
xnor U26740 (N_26740,N_26183,N_26105);
nor U26741 (N_26741,N_26356,N_26268);
and U26742 (N_26742,N_26163,N_26439);
xor U26743 (N_26743,N_26379,N_26192);
or U26744 (N_26744,N_26231,N_26046);
nand U26745 (N_26745,N_26079,N_26103);
xor U26746 (N_26746,N_26378,N_26266);
and U26747 (N_26747,N_26177,N_26196);
xor U26748 (N_26748,N_26324,N_26337);
nor U26749 (N_26749,N_26350,N_26321);
or U26750 (N_26750,N_26451,N_26461);
nand U26751 (N_26751,N_26186,N_26319);
nand U26752 (N_26752,N_26486,N_26379);
nor U26753 (N_26753,N_26229,N_26013);
or U26754 (N_26754,N_26050,N_26005);
and U26755 (N_26755,N_26409,N_26247);
or U26756 (N_26756,N_26125,N_26236);
xor U26757 (N_26757,N_26303,N_26008);
and U26758 (N_26758,N_26348,N_26392);
and U26759 (N_26759,N_26312,N_26269);
or U26760 (N_26760,N_26173,N_26320);
nor U26761 (N_26761,N_26307,N_26277);
xor U26762 (N_26762,N_26131,N_26102);
nand U26763 (N_26763,N_26219,N_26377);
or U26764 (N_26764,N_26007,N_26123);
or U26765 (N_26765,N_26324,N_26025);
nor U26766 (N_26766,N_26481,N_26490);
nor U26767 (N_26767,N_26210,N_26364);
nor U26768 (N_26768,N_26184,N_26143);
and U26769 (N_26769,N_26300,N_26325);
nand U26770 (N_26770,N_26200,N_26390);
nor U26771 (N_26771,N_26308,N_26047);
and U26772 (N_26772,N_26308,N_26210);
nand U26773 (N_26773,N_26430,N_26480);
and U26774 (N_26774,N_26483,N_26358);
xor U26775 (N_26775,N_26335,N_26095);
nand U26776 (N_26776,N_26144,N_26027);
xor U26777 (N_26777,N_26327,N_26028);
or U26778 (N_26778,N_26061,N_26060);
nand U26779 (N_26779,N_26396,N_26259);
nor U26780 (N_26780,N_26425,N_26363);
and U26781 (N_26781,N_26484,N_26353);
and U26782 (N_26782,N_26386,N_26264);
and U26783 (N_26783,N_26349,N_26430);
or U26784 (N_26784,N_26224,N_26227);
nor U26785 (N_26785,N_26383,N_26445);
nor U26786 (N_26786,N_26443,N_26357);
or U26787 (N_26787,N_26206,N_26352);
nand U26788 (N_26788,N_26440,N_26286);
xor U26789 (N_26789,N_26409,N_26086);
or U26790 (N_26790,N_26271,N_26262);
and U26791 (N_26791,N_26326,N_26122);
and U26792 (N_26792,N_26211,N_26083);
or U26793 (N_26793,N_26337,N_26344);
nand U26794 (N_26794,N_26126,N_26441);
xor U26795 (N_26795,N_26039,N_26369);
xor U26796 (N_26796,N_26015,N_26118);
and U26797 (N_26797,N_26045,N_26166);
xor U26798 (N_26798,N_26283,N_26114);
nand U26799 (N_26799,N_26229,N_26422);
or U26800 (N_26800,N_26105,N_26061);
and U26801 (N_26801,N_26312,N_26366);
xnor U26802 (N_26802,N_26076,N_26269);
nor U26803 (N_26803,N_26498,N_26450);
nand U26804 (N_26804,N_26140,N_26239);
and U26805 (N_26805,N_26039,N_26101);
nor U26806 (N_26806,N_26478,N_26147);
and U26807 (N_26807,N_26349,N_26355);
and U26808 (N_26808,N_26080,N_26005);
or U26809 (N_26809,N_26092,N_26097);
xnor U26810 (N_26810,N_26324,N_26144);
and U26811 (N_26811,N_26273,N_26172);
and U26812 (N_26812,N_26200,N_26378);
nor U26813 (N_26813,N_26198,N_26480);
and U26814 (N_26814,N_26326,N_26230);
nand U26815 (N_26815,N_26453,N_26067);
xnor U26816 (N_26816,N_26393,N_26066);
nor U26817 (N_26817,N_26453,N_26046);
or U26818 (N_26818,N_26473,N_26427);
or U26819 (N_26819,N_26075,N_26272);
or U26820 (N_26820,N_26044,N_26226);
nor U26821 (N_26821,N_26469,N_26014);
nor U26822 (N_26822,N_26106,N_26232);
xor U26823 (N_26823,N_26225,N_26389);
or U26824 (N_26824,N_26193,N_26055);
nor U26825 (N_26825,N_26499,N_26448);
nor U26826 (N_26826,N_26153,N_26486);
xor U26827 (N_26827,N_26181,N_26003);
and U26828 (N_26828,N_26310,N_26293);
xnor U26829 (N_26829,N_26245,N_26061);
nand U26830 (N_26830,N_26465,N_26422);
or U26831 (N_26831,N_26411,N_26309);
xnor U26832 (N_26832,N_26321,N_26025);
xor U26833 (N_26833,N_26123,N_26053);
nor U26834 (N_26834,N_26397,N_26258);
nor U26835 (N_26835,N_26303,N_26388);
and U26836 (N_26836,N_26320,N_26125);
nor U26837 (N_26837,N_26344,N_26356);
or U26838 (N_26838,N_26406,N_26253);
and U26839 (N_26839,N_26213,N_26219);
nand U26840 (N_26840,N_26235,N_26014);
or U26841 (N_26841,N_26452,N_26264);
xor U26842 (N_26842,N_26050,N_26306);
xnor U26843 (N_26843,N_26363,N_26489);
xnor U26844 (N_26844,N_26494,N_26021);
or U26845 (N_26845,N_26422,N_26042);
and U26846 (N_26846,N_26490,N_26497);
nor U26847 (N_26847,N_26048,N_26288);
or U26848 (N_26848,N_26339,N_26370);
xor U26849 (N_26849,N_26009,N_26497);
or U26850 (N_26850,N_26294,N_26281);
nor U26851 (N_26851,N_26190,N_26243);
nor U26852 (N_26852,N_26244,N_26313);
xnor U26853 (N_26853,N_26251,N_26339);
and U26854 (N_26854,N_26300,N_26197);
or U26855 (N_26855,N_26226,N_26239);
or U26856 (N_26856,N_26212,N_26360);
and U26857 (N_26857,N_26337,N_26094);
or U26858 (N_26858,N_26447,N_26330);
xor U26859 (N_26859,N_26023,N_26379);
or U26860 (N_26860,N_26453,N_26172);
or U26861 (N_26861,N_26168,N_26274);
nand U26862 (N_26862,N_26483,N_26114);
or U26863 (N_26863,N_26280,N_26182);
and U26864 (N_26864,N_26139,N_26009);
nand U26865 (N_26865,N_26136,N_26483);
or U26866 (N_26866,N_26231,N_26317);
nor U26867 (N_26867,N_26093,N_26374);
or U26868 (N_26868,N_26468,N_26441);
nor U26869 (N_26869,N_26404,N_26088);
nor U26870 (N_26870,N_26093,N_26358);
nand U26871 (N_26871,N_26187,N_26229);
nand U26872 (N_26872,N_26325,N_26126);
xnor U26873 (N_26873,N_26149,N_26238);
nor U26874 (N_26874,N_26441,N_26171);
nor U26875 (N_26875,N_26493,N_26088);
nand U26876 (N_26876,N_26113,N_26206);
nor U26877 (N_26877,N_26447,N_26148);
nor U26878 (N_26878,N_26291,N_26318);
or U26879 (N_26879,N_26434,N_26216);
nand U26880 (N_26880,N_26132,N_26435);
xor U26881 (N_26881,N_26194,N_26446);
nand U26882 (N_26882,N_26170,N_26292);
and U26883 (N_26883,N_26107,N_26008);
and U26884 (N_26884,N_26432,N_26340);
xnor U26885 (N_26885,N_26358,N_26432);
nand U26886 (N_26886,N_26390,N_26074);
or U26887 (N_26887,N_26402,N_26400);
or U26888 (N_26888,N_26436,N_26284);
and U26889 (N_26889,N_26103,N_26323);
and U26890 (N_26890,N_26105,N_26200);
and U26891 (N_26891,N_26275,N_26470);
or U26892 (N_26892,N_26145,N_26017);
nand U26893 (N_26893,N_26202,N_26093);
xor U26894 (N_26894,N_26326,N_26014);
xnor U26895 (N_26895,N_26263,N_26442);
xnor U26896 (N_26896,N_26102,N_26337);
or U26897 (N_26897,N_26397,N_26011);
nand U26898 (N_26898,N_26451,N_26091);
or U26899 (N_26899,N_26350,N_26317);
xor U26900 (N_26900,N_26345,N_26354);
xor U26901 (N_26901,N_26125,N_26210);
nor U26902 (N_26902,N_26146,N_26061);
and U26903 (N_26903,N_26426,N_26101);
or U26904 (N_26904,N_26034,N_26205);
nand U26905 (N_26905,N_26183,N_26072);
nand U26906 (N_26906,N_26403,N_26282);
xor U26907 (N_26907,N_26109,N_26244);
nor U26908 (N_26908,N_26065,N_26365);
or U26909 (N_26909,N_26167,N_26112);
nand U26910 (N_26910,N_26410,N_26214);
or U26911 (N_26911,N_26362,N_26276);
and U26912 (N_26912,N_26268,N_26012);
nand U26913 (N_26913,N_26179,N_26340);
or U26914 (N_26914,N_26309,N_26124);
nor U26915 (N_26915,N_26350,N_26245);
nand U26916 (N_26916,N_26429,N_26490);
and U26917 (N_26917,N_26264,N_26248);
or U26918 (N_26918,N_26203,N_26106);
or U26919 (N_26919,N_26124,N_26255);
or U26920 (N_26920,N_26387,N_26028);
nand U26921 (N_26921,N_26149,N_26211);
nand U26922 (N_26922,N_26081,N_26250);
or U26923 (N_26923,N_26121,N_26473);
nor U26924 (N_26924,N_26196,N_26002);
nand U26925 (N_26925,N_26116,N_26436);
and U26926 (N_26926,N_26276,N_26400);
and U26927 (N_26927,N_26008,N_26342);
or U26928 (N_26928,N_26168,N_26394);
or U26929 (N_26929,N_26384,N_26448);
nand U26930 (N_26930,N_26096,N_26430);
nor U26931 (N_26931,N_26252,N_26385);
nand U26932 (N_26932,N_26300,N_26042);
nand U26933 (N_26933,N_26321,N_26472);
and U26934 (N_26934,N_26433,N_26086);
nor U26935 (N_26935,N_26047,N_26008);
and U26936 (N_26936,N_26207,N_26482);
xor U26937 (N_26937,N_26455,N_26011);
and U26938 (N_26938,N_26180,N_26298);
nor U26939 (N_26939,N_26315,N_26498);
or U26940 (N_26940,N_26080,N_26383);
and U26941 (N_26941,N_26487,N_26264);
nand U26942 (N_26942,N_26101,N_26324);
nand U26943 (N_26943,N_26079,N_26277);
and U26944 (N_26944,N_26238,N_26438);
nand U26945 (N_26945,N_26381,N_26234);
xor U26946 (N_26946,N_26461,N_26252);
and U26947 (N_26947,N_26326,N_26358);
or U26948 (N_26948,N_26152,N_26309);
xnor U26949 (N_26949,N_26281,N_26196);
nand U26950 (N_26950,N_26006,N_26254);
nor U26951 (N_26951,N_26324,N_26124);
nor U26952 (N_26952,N_26266,N_26383);
nor U26953 (N_26953,N_26304,N_26468);
and U26954 (N_26954,N_26237,N_26048);
nor U26955 (N_26955,N_26164,N_26093);
xor U26956 (N_26956,N_26045,N_26248);
and U26957 (N_26957,N_26276,N_26184);
nor U26958 (N_26958,N_26480,N_26482);
and U26959 (N_26959,N_26227,N_26461);
xnor U26960 (N_26960,N_26376,N_26348);
nor U26961 (N_26961,N_26207,N_26001);
and U26962 (N_26962,N_26152,N_26412);
xor U26963 (N_26963,N_26249,N_26386);
nand U26964 (N_26964,N_26211,N_26282);
nand U26965 (N_26965,N_26329,N_26359);
xnor U26966 (N_26966,N_26361,N_26443);
nand U26967 (N_26967,N_26257,N_26360);
nand U26968 (N_26968,N_26262,N_26137);
or U26969 (N_26969,N_26213,N_26464);
and U26970 (N_26970,N_26382,N_26438);
nor U26971 (N_26971,N_26474,N_26447);
xor U26972 (N_26972,N_26138,N_26074);
or U26973 (N_26973,N_26447,N_26498);
or U26974 (N_26974,N_26295,N_26084);
nand U26975 (N_26975,N_26426,N_26053);
xor U26976 (N_26976,N_26322,N_26008);
or U26977 (N_26977,N_26369,N_26126);
xor U26978 (N_26978,N_26435,N_26339);
nor U26979 (N_26979,N_26489,N_26005);
nor U26980 (N_26980,N_26494,N_26108);
and U26981 (N_26981,N_26152,N_26015);
nor U26982 (N_26982,N_26154,N_26048);
and U26983 (N_26983,N_26324,N_26082);
and U26984 (N_26984,N_26376,N_26393);
nor U26985 (N_26985,N_26379,N_26355);
nand U26986 (N_26986,N_26467,N_26423);
or U26987 (N_26987,N_26380,N_26149);
nand U26988 (N_26988,N_26088,N_26217);
nor U26989 (N_26989,N_26071,N_26368);
nor U26990 (N_26990,N_26290,N_26107);
nor U26991 (N_26991,N_26342,N_26134);
nor U26992 (N_26992,N_26392,N_26373);
xnor U26993 (N_26993,N_26171,N_26466);
nor U26994 (N_26994,N_26353,N_26245);
xnor U26995 (N_26995,N_26044,N_26087);
xnor U26996 (N_26996,N_26317,N_26144);
or U26997 (N_26997,N_26345,N_26328);
nand U26998 (N_26998,N_26053,N_26344);
and U26999 (N_26999,N_26005,N_26363);
nor U27000 (N_27000,N_26658,N_26602);
nand U27001 (N_27001,N_26846,N_26760);
nor U27002 (N_27002,N_26519,N_26879);
nand U27003 (N_27003,N_26682,N_26515);
xnor U27004 (N_27004,N_26777,N_26980);
nor U27005 (N_27005,N_26954,N_26797);
nand U27006 (N_27006,N_26664,N_26925);
xnor U27007 (N_27007,N_26520,N_26801);
xor U27008 (N_27008,N_26819,N_26653);
nor U27009 (N_27009,N_26942,N_26640);
xnor U27010 (N_27010,N_26953,N_26633);
nor U27011 (N_27011,N_26986,N_26768);
nor U27012 (N_27012,N_26997,N_26504);
nor U27013 (N_27013,N_26606,N_26669);
nand U27014 (N_27014,N_26680,N_26533);
and U27015 (N_27015,N_26648,N_26730);
xor U27016 (N_27016,N_26800,N_26710);
nor U27017 (N_27017,N_26556,N_26848);
nor U27018 (N_27018,N_26774,N_26950);
xor U27019 (N_27019,N_26558,N_26501);
nand U27020 (N_27020,N_26759,N_26857);
xnor U27021 (N_27021,N_26655,N_26629);
nand U27022 (N_27022,N_26766,N_26994);
and U27023 (N_27023,N_26502,N_26827);
or U27024 (N_27024,N_26749,N_26559);
xor U27025 (N_27025,N_26951,N_26686);
and U27026 (N_27026,N_26940,N_26674);
or U27027 (N_27027,N_26804,N_26647);
and U27028 (N_27028,N_26784,N_26833);
nand U27029 (N_27029,N_26775,N_26931);
nor U27030 (N_27030,N_26756,N_26945);
nor U27031 (N_27031,N_26522,N_26660);
or U27032 (N_27032,N_26729,N_26896);
and U27033 (N_27033,N_26864,N_26512);
xnor U27034 (N_27034,N_26972,N_26707);
nor U27035 (N_27035,N_26910,N_26700);
xnor U27036 (N_27036,N_26635,N_26875);
nor U27037 (N_27037,N_26921,N_26706);
or U27038 (N_27038,N_26928,N_26685);
nor U27039 (N_27039,N_26897,N_26981);
nor U27040 (N_27040,N_26553,N_26575);
xor U27041 (N_27041,N_26528,N_26592);
and U27042 (N_27042,N_26870,N_26702);
and U27043 (N_27043,N_26531,N_26639);
xor U27044 (N_27044,N_26943,N_26649);
and U27045 (N_27045,N_26672,N_26899);
xor U27046 (N_27046,N_26565,N_26969);
nand U27047 (N_27047,N_26826,N_26934);
or U27048 (N_27048,N_26740,N_26936);
nand U27049 (N_27049,N_26718,N_26576);
nand U27050 (N_27050,N_26891,N_26693);
xnor U27051 (N_27051,N_26789,N_26738);
nand U27052 (N_27052,N_26927,N_26643);
nand U27053 (N_27053,N_26714,N_26871);
and U27054 (N_27054,N_26569,N_26703);
nand U27055 (N_27055,N_26816,N_26652);
or U27056 (N_27056,N_26673,N_26621);
and U27057 (N_27057,N_26930,N_26709);
or U27058 (N_27058,N_26546,N_26688);
xor U27059 (N_27059,N_26771,N_26717);
and U27060 (N_27060,N_26661,N_26666);
or U27061 (N_27061,N_26701,N_26572);
or U27062 (N_27062,N_26723,N_26765);
or U27063 (N_27063,N_26787,N_26825);
or U27064 (N_27064,N_26868,N_26617);
xor U27065 (N_27065,N_26841,N_26835);
xor U27066 (N_27066,N_26935,N_26968);
nor U27067 (N_27067,N_26625,N_26914);
or U27068 (N_27068,N_26615,N_26806);
nor U27069 (N_27069,N_26975,N_26788);
xnor U27070 (N_27070,N_26743,N_26588);
nor U27071 (N_27071,N_26690,N_26890);
nand U27072 (N_27072,N_26607,N_26585);
xor U27073 (N_27073,N_26911,N_26903);
and U27074 (N_27074,N_26810,N_26503);
xnor U27075 (N_27075,N_26527,N_26798);
nand U27076 (N_27076,N_26555,N_26694);
nor U27077 (N_27077,N_26644,N_26795);
and U27078 (N_27078,N_26962,N_26862);
and U27079 (N_27079,N_26605,N_26614);
or U27080 (N_27080,N_26873,N_26638);
xor U27081 (N_27081,N_26529,N_26889);
or U27082 (N_27082,N_26594,N_26601);
and U27083 (N_27083,N_26739,N_26654);
or U27084 (N_27084,N_26755,N_26513);
or U27085 (N_27085,N_26853,N_26637);
xnor U27086 (N_27086,N_26807,N_26947);
and U27087 (N_27087,N_26987,N_26850);
and U27088 (N_27088,N_26630,N_26915);
nand U27089 (N_27089,N_26802,N_26562);
or U27090 (N_27090,N_26741,N_26623);
or U27091 (N_27091,N_26544,N_26860);
and U27092 (N_27092,N_26995,N_26612);
or U27093 (N_27093,N_26970,N_26832);
and U27094 (N_27094,N_26855,N_26811);
and U27095 (N_27095,N_26874,N_26699);
or U27096 (N_27096,N_26747,N_26753);
and U27097 (N_27097,N_26821,N_26627);
and U27098 (N_27098,N_26563,N_26634);
or U27099 (N_27099,N_26878,N_26781);
or U27100 (N_27100,N_26847,N_26941);
or U27101 (N_27101,N_26772,N_26955);
nor U27102 (N_27102,N_26780,N_26996);
xor U27103 (N_27103,N_26737,N_26902);
or U27104 (N_27104,N_26919,N_26991);
nand U27105 (N_27105,N_26603,N_26507);
or U27106 (N_27106,N_26577,N_26523);
nand U27107 (N_27107,N_26920,N_26861);
xor U27108 (N_27108,N_26731,N_26641);
and U27109 (N_27109,N_26887,N_26877);
nor U27110 (N_27110,N_26564,N_26793);
or U27111 (N_27111,N_26837,N_26537);
and U27112 (N_27112,N_26786,N_26525);
nor U27113 (N_27113,N_26814,N_26657);
or U27114 (N_27114,N_26608,N_26521);
nor U27115 (N_27115,N_26586,N_26626);
xor U27116 (N_27116,N_26982,N_26705);
or U27117 (N_27117,N_26509,N_26882);
and U27118 (N_27118,N_26526,N_26551);
nor U27119 (N_27119,N_26552,N_26582);
xnor U27120 (N_27120,N_26984,N_26778);
xor U27121 (N_27121,N_26557,N_26611);
nor U27122 (N_27122,N_26510,N_26845);
nor U27123 (N_27123,N_26895,N_26662);
xor U27124 (N_27124,N_26754,N_26763);
nor U27125 (N_27125,N_26712,N_26720);
xnor U27126 (N_27126,N_26906,N_26550);
xor U27127 (N_27127,N_26888,N_26578);
nand U27128 (N_27128,N_26842,N_26764);
xnor U27129 (N_27129,N_26719,N_26727);
and U27130 (N_27130,N_26813,N_26618);
nand U27131 (N_27131,N_26628,N_26535);
xor U27132 (N_27132,N_26536,N_26990);
or U27133 (N_27133,N_26574,N_26993);
xor U27134 (N_27134,N_26966,N_26622);
and U27135 (N_27135,N_26865,N_26584);
nor U27136 (N_27136,N_26532,N_26783);
or U27137 (N_27137,N_26632,N_26758);
nand U27138 (N_27138,N_26595,N_26677);
or U27139 (N_27139,N_26851,N_26604);
nor U27140 (N_27140,N_26790,N_26583);
or U27141 (N_27141,N_26866,N_26971);
and U27142 (N_27142,N_26561,N_26988);
nand U27143 (N_27143,N_26883,N_26500);
nand U27144 (N_27144,N_26518,N_26734);
and U27145 (N_27145,N_26824,N_26828);
xor U27146 (N_27146,N_26668,N_26681);
nor U27147 (N_27147,N_26963,N_26684);
or U27148 (N_27148,N_26964,N_26867);
or U27149 (N_27149,N_26769,N_26676);
nand U27150 (N_27150,N_26696,N_26506);
xnor U27151 (N_27151,N_26619,N_26530);
xnor U27152 (N_27152,N_26683,N_26748);
nor U27153 (N_27153,N_26908,N_26616);
and U27154 (N_27154,N_26838,N_26610);
nor U27155 (N_27155,N_26998,N_26913);
nor U27156 (N_27156,N_26923,N_26894);
nor U27157 (N_27157,N_26695,N_26983);
or U27158 (N_27158,N_26762,N_26593);
nand U27159 (N_27159,N_26679,N_26960);
xor U27160 (N_27160,N_26542,N_26967);
xor U27161 (N_27161,N_26568,N_26820);
or U27162 (N_27162,N_26973,N_26534);
nand U27163 (N_27163,N_26721,N_26692);
nor U27164 (N_27164,N_26933,N_26733);
nand U27165 (N_27165,N_26961,N_26805);
nor U27166 (N_27166,N_26946,N_26932);
or U27167 (N_27167,N_26566,N_26830);
and U27168 (N_27168,N_26948,N_26886);
or U27169 (N_27169,N_26571,N_26803);
nor U27170 (N_27170,N_26881,N_26916);
nand U27171 (N_27171,N_26650,N_26905);
and U27172 (N_27172,N_26907,N_26773);
and U27173 (N_27173,N_26691,N_26989);
nor U27174 (N_27174,N_26959,N_26976);
nor U27175 (N_27175,N_26651,N_26596);
nand U27176 (N_27176,N_26770,N_26573);
or U27177 (N_27177,N_26722,N_26876);
and U27178 (N_27178,N_26761,N_26540);
nand U27179 (N_27179,N_26999,N_26587);
xnor U27180 (N_27180,N_26517,N_26904);
and U27181 (N_27181,N_26646,N_26742);
and U27182 (N_27182,N_26547,N_26809);
and U27183 (N_27183,N_26977,N_26645);
nor U27184 (N_27184,N_26598,N_26929);
or U27185 (N_27185,N_26843,N_26918);
nor U27186 (N_27186,N_26538,N_26831);
and U27187 (N_27187,N_26901,N_26750);
nor U27188 (N_27188,N_26687,N_26815);
xnor U27189 (N_27189,N_26579,N_26689);
nand U27190 (N_27190,N_26785,N_26880);
xor U27191 (N_27191,N_26757,N_26708);
or U27192 (N_27192,N_26799,N_26898);
nand U27193 (N_27193,N_26746,N_26840);
or U27194 (N_27194,N_26985,N_26613);
nor U27195 (N_27195,N_26726,N_26590);
xor U27196 (N_27196,N_26979,N_26912);
xnor U27197 (N_27197,N_26567,N_26505);
nand U27198 (N_27198,N_26745,N_26670);
nand U27199 (N_27199,N_26600,N_26711);
xor U27200 (N_27200,N_26965,N_26675);
or U27201 (N_27201,N_26570,N_26872);
and U27202 (N_27202,N_26952,N_26885);
and U27203 (N_27203,N_26944,N_26663);
nand U27204 (N_27204,N_26597,N_26808);
and U27205 (N_27205,N_26716,N_26508);
nand U27206 (N_27206,N_26839,N_26822);
and U27207 (N_27207,N_26949,N_26698);
xnor U27208 (N_27208,N_26704,N_26580);
nor U27209 (N_27209,N_26869,N_26665);
xnor U27210 (N_27210,N_26958,N_26697);
nor U27211 (N_27211,N_26836,N_26554);
and U27212 (N_27212,N_26844,N_26856);
xnor U27213 (N_27213,N_26854,N_26909);
and U27214 (N_27214,N_26591,N_26581);
xor U27215 (N_27215,N_26794,N_26782);
nand U27216 (N_27216,N_26642,N_26725);
xnor U27217 (N_27217,N_26545,N_26543);
and U27218 (N_27218,N_26884,N_26818);
nand U27219 (N_27219,N_26956,N_26541);
nor U27220 (N_27220,N_26767,N_26924);
and U27221 (N_27221,N_26852,N_26812);
xnor U27222 (N_27222,N_26631,N_26549);
and U27223 (N_27223,N_26667,N_26744);
nor U27224 (N_27224,N_26609,N_26957);
xor U27225 (N_27225,N_26776,N_26978);
xnor U27226 (N_27226,N_26751,N_26516);
nor U27227 (N_27227,N_26834,N_26589);
and U27228 (N_27228,N_26829,N_26659);
nor U27229 (N_27229,N_26937,N_26859);
xor U27230 (N_27230,N_26791,N_26539);
nand U27231 (N_27231,N_26779,N_26863);
or U27232 (N_27232,N_26636,N_26713);
and U27233 (N_27233,N_26715,N_26678);
or U27234 (N_27234,N_26671,N_26858);
and U27235 (N_27235,N_26735,N_26992);
and U27236 (N_27236,N_26893,N_26926);
nand U27237 (N_27237,N_26599,N_26939);
or U27238 (N_27238,N_26736,N_26823);
xor U27239 (N_27239,N_26624,N_26548);
xnor U27240 (N_27240,N_26922,N_26892);
nand U27241 (N_27241,N_26560,N_26724);
nand U27242 (N_27242,N_26728,N_26514);
xor U27243 (N_27243,N_26849,N_26511);
xor U27244 (N_27244,N_26524,N_26900);
and U27245 (N_27245,N_26792,N_26796);
xor U27246 (N_27246,N_26917,N_26620);
nor U27247 (N_27247,N_26817,N_26732);
nor U27248 (N_27248,N_26656,N_26938);
nor U27249 (N_27249,N_26752,N_26974);
xor U27250 (N_27250,N_26927,N_26695);
xnor U27251 (N_27251,N_26774,N_26905);
nand U27252 (N_27252,N_26907,N_26739);
and U27253 (N_27253,N_26616,N_26873);
and U27254 (N_27254,N_26683,N_26878);
and U27255 (N_27255,N_26572,N_26649);
and U27256 (N_27256,N_26640,N_26631);
xnor U27257 (N_27257,N_26620,N_26715);
nor U27258 (N_27258,N_26528,N_26750);
nor U27259 (N_27259,N_26576,N_26804);
xor U27260 (N_27260,N_26609,N_26907);
nand U27261 (N_27261,N_26691,N_26881);
or U27262 (N_27262,N_26568,N_26778);
or U27263 (N_27263,N_26754,N_26791);
xnor U27264 (N_27264,N_26533,N_26975);
nand U27265 (N_27265,N_26802,N_26512);
nor U27266 (N_27266,N_26852,N_26882);
xnor U27267 (N_27267,N_26766,N_26571);
xnor U27268 (N_27268,N_26551,N_26510);
nor U27269 (N_27269,N_26709,N_26518);
nand U27270 (N_27270,N_26664,N_26634);
or U27271 (N_27271,N_26630,N_26796);
nor U27272 (N_27272,N_26542,N_26877);
or U27273 (N_27273,N_26816,N_26654);
and U27274 (N_27274,N_26656,N_26769);
nand U27275 (N_27275,N_26769,N_26909);
or U27276 (N_27276,N_26833,N_26575);
and U27277 (N_27277,N_26696,N_26800);
nor U27278 (N_27278,N_26792,N_26774);
nor U27279 (N_27279,N_26961,N_26630);
nor U27280 (N_27280,N_26529,N_26535);
nor U27281 (N_27281,N_26943,N_26988);
nor U27282 (N_27282,N_26892,N_26843);
and U27283 (N_27283,N_26886,N_26577);
nand U27284 (N_27284,N_26577,N_26891);
nand U27285 (N_27285,N_26663,N_26740);
nor U27286 (N_27286,N_26594,N_26537);
xnor U27287 (N_27287,N_26712,N_26936);
nor U27288 (N_27288,N_26646,N_26712);
xnor U27289 (N_27289,N_26725,N_26711);
or U27290 (N_27290,N_26503,N_26568);
and U27291 (N_27291,N_26676,N_26934);
and U27292 (N_27292,N_26966,N_26664);
nor U27293 (N_27293,N_26936,N_26850);
and U27294 (N_27294,N_26506,N_26957);
and U27295 (N_27295,N_26944,N_26978);
or U27296 (N_27296,N_26833,N_26512);
nand U27297 (N_27297,N_26630,N_26974);
nand U27298 (N_27298,N_26712,N_26861);
and U27299 (N_27299,N_26947,N_26940);
nand U27300 (N_27300,N_26949,N_26587);
nand U27301 (N_27301,N_26948,N_26578);
nor U27302 (N_27302,N_26789,N_26881);
xnor U27303 (N_27303,N_26941,N_26533);
and U27304 (N_27304,N_26586,N_26944);
and U27305 (N_27305,N_26564,N_26517);
and U27306 (N_27306,N_26545,N_26726);
xnor U27307 (N_27307,N_26738,N_26990);
xor U27308 (N_27308,N_26999,N_26903);
xor U27309 (N_27309,N_26723,N_26519);
xor U27310 (N_27310,N_26634,N_26717);
nor U27311 (N_27311,N_26764,N_26994);
xnor U27312 (N_27312,N_26519,N_26855);
nor U27313 (N_27313,N_26884,N_26770);
and U27314 (N_27314,N_26539,N_26804);
and U27315 (N_27315,N_26967,N_26887);
nand U27316 (N_27316,N_26644,N_26549);
or U27317 (N_27317,N_26626,N_26565);
or U27318 (N_27318,N_26738,N_26528);
xor U27319 (N_27319,N_26760,N_26795);
xor U27320 (N_27320,N_26743,N_26629);
and U27321 (N_27321,N_26649,N_26597);
nor U27322 (N_27322,N_26921,N_26918);
or U27323 (N_27323,N_26874,N_26581);
nor U27324 (N_27324,N_26640,N_26954);
and U27325 (N_27325,N_26869,N_26672);
nor U27326 (N_27326,N_26711,N_26956);
nor U27327 (N_27327,N_26539,N_26574);
xor U27328 (N_27328,N_26677,N_26912);
and U27329 (N_27329,N_26645,N_26585);
nand U27330 (N_27330,N_26856,N_26921);
nor U27331 (N_27331,N_26695,N_26599);
and U27332 (N_27332,N_26585,N_26812);
or U27333 (N_27333,N_26671,N_26832);
or U27334 (N_27334,N_26779,N_26510);
nand U27335 (N_27335,N_26731,N_26873);
nand U27336 (N_27336,N_26563,N_26819);
nor U27337 (N_27337,N_26565,N_26539);
or U27338 (N_27338,N_26647,N_26572);
nand U27339 (N_27339,N_26925,N_26604);
and U27340 (N_27340,N_26838,N_26830);
or U27341 (N_27341,N_26533,N_26678);
nor U27342 (N_27342,N_26675,N_26787);
and U27343 (N_27343,N_26819,N_26722);
nand U27344 (N_27344,N_26707,N_26852);
nand U27345 (N_27345,N_26706,N_26998);
nor U27346 (N_27346,N_26974,N_26688);
nand U27347 (N_27347,N_26951,N_26792);
nand U27348 (N_27348,N_26573,N_26763);
xor U27349 (N_27349,N_26659,N_26528);
or U27350 (N_27350,N_26997,N_26913);
nand U27351 (N_27351,N_26870,N_26902);
xnor U27352 (N_27352,N_26747,N_26861);
xor U27353 (N_27353,N_26910,N_26939);
and U27354 (N_27354,N_26775,N_26972);
nor U27355 (N_27355,N_26894,N_26935);
and U27356 (N_27356,N_26601,N_26522);
nor U27357 (N_27357,N_26993,N_26518);
xnor U27358 (N_27358,N_26978,N_26703);
and U27359 (N_27359,N_26509,N_26507);
or U27360 (N_27360,N_26825,N_26814);
xnor U27361 (N_27361,N_26621,N_26759);
or U27362 (N_27362,N_26859,N_26783);
or U27363 (N_27363,N_26620,N_26900);
nand U27364 (N_27364,N_26578,N_26913);
xor U27365 (N_27365,N_26582,N_26578);
nor U27366 (N_27366,N_26866,N_26677);
or U27367 (N_27367,N_26627,N_26823);
nor U27368 (N_27368,N_26736,N_26528);
xnor U27369 (N_27369,N_26604,N_26663);
or U27370 (N_27370,N_26953,N_26657);
nor U27371 (N_27371,N_26519,N_26730);
xnor U27372 (N_27372,N_26534,N_26734);
nand U27373 (N_27373,N_26981,N_26603);
xnor U27374 (N_27374,N_26963,N_26508);
or U27375 (N_27375,N_26631,N_26619);
xor U27376 (N_27376,N_26632,N_26962);
nand U27377 (N_27377,N_26941,N_26797);
nor U27378 (N_27378,N_26679,N_26821);
xor U27379 (N_27379,N_26975,N_26622);
and U27380 (N_27380,N_26727,N_26629);
and U27381 (N_27381,N_26619,N_26606);
and U27382 (N_27382,N_26707,N_26956);
or U27383 (N_27383,N_26603,N_26620);
or U27384 (N_27384,N_26577,N_26612);
nand U27385 (N_27385,N_26658,N_26997);
nor U27386 (N_27386,N_26502,N_26598);
xnor U27387 (N_27387,N_26638,N_26780);
xor U27388 (N_27388,N_26787,N_26881);
and U27389 (N_27389,N_26806,N_26927);
or U27390 (N_27390,N_26839,N_26656);
nor U27391 (N_27391,N_26527,N_26713);
or U27392 (N_27392,N_26519,N_26577);
or U27393 (N_27393,N_26885,N_26673);
nand U27394 (N_27394,N_26693,N_26890);
nor U27395 (N_27395,N_26599,N_26991);
nand U27396 (N_27396,N_26788,N_26681);
and U27397 (N_27397,N_26813,N_26664);
nand U27398 (N_27398,N_26562,N_26602);
nand U27399 (N_27399,N_26827,N_26708);
nor U27400 (N_27400,N_26507,N_26659);
or U27401 (N_27401,N_26856,N_26538);
nand U27402 (N_27402,N_26827,N_26518);
xor U27403 (N_27403,N_26530,N_26766);
and U27404 (N_27404,N_26506,N_26679);
xor U27405 (N_27405,N_26561,N_26593);
xnor U27406 (N_27406,N_26865,N_26589);
xnor U27407 (N_27407,N_26708,N_26855);
nor U27408 (N_27408,N_26718,N_26719);
xnor U27409 (N_27409,N_26819,N_26759);
xor U27410 (N_27410,N_26943,N_26623);
nand U27411 (N_27411,N_26944,N_26837);
or U27412 (N_27412,N_26839,N_26977);
nor U27413 (N_27413,N_26810,N_26671);
nand U27414 (N_27414,N_26690,N_26961);
xnor U27415 (N_27415,N_26694,N_26955);
or U27416 (N_27416,N_26802,N_26549);
xor U27417 (N_27417,N_26511,N_26684);
and U27418 (N_27418,N_26529,N_26678);
nand U27419 (N_27419,N_26885,N_26613);
nor U27420 (N_27420,N_26912,N_26639);
xor U27421 (N_27421,N_26622,N_26594);
and U27422 (N_27422,N_26958,N_26670);
and U27423 (N_27423,N_26938,N_26600);
nor U27424 (N_27424,N_26968,N_26612);
xor U27425 (N_27425,N_26900,N_26974);
xnor U27426 (N_27426,N_26806,N_26703);
and U27427 (N_27427,N_26773,N_26828);
and U27428 (N_27428,N_26582,N_26678);
or U27429 (N_27429,N_26905,N_26880);
nor U27430 (N_27430,N_26964,N_26887);
and U27431 (N_27431,N_26859,N_26851);
nor U27432 (N_27432,N_26825,N_26777);
and U27433 (N_27433,N_26843,N_26640);
nor U27434 (N_27434,N_26994,N_26776);
and U27435 (N_27435,N_26939,N_26797);
and U27436 (N_27436,N_26538,N_26510);
nand U27437 (N_27437,N_26929,N_26512);
or U27438 (N_27438,N_26776,N_26709);
or U27439 (N_27439,N_26612,N_26510);
nor U27440 (N_27440,N_26653,N_26853);
nor U27441 (N_27441,N_26519,N_26866);
and U27442 (N_27442,N_26592,N_26529);
nor U27443 (N_27443,N_26673,N_26989);
nor U27444 (N_27444,N_26709,N_26607);
nor U27445 (N_27445,N_26938,N_26955);
or U27446 (N_27446,N_26838,N_26674);
xor U27447 (N_27447,N_26868,N_26669);
nand U27448 (N_27448,N_26774,N_26864);
nand U27449 (N_27449,N_26824,N_26592);
nand U27450 (N_27450,N_26763,N_26602);
or U27451 (N_27451,N_26826,N_26976);
or U27452 (N_27452,N_26691,N_26973);
xor U27453 (N_27453,N_26572,N_26803);
nand U27454 (N_27454,N_26840,N_26994);
nand U27455 (N_27455,N_26916,N_26876);
nor U27456 (N_27456,N_26663,N_26967);
and U27457 (N_27457,N_26665,N_26514);
nor U27458 (N_27458,N_26865,N_26960);
and U27459 (N_27459,N_26757,N_26627);
xnor U27460 (N_27460,N_26749,N_26539);
nand U27461 (N_27461,N_26946,N_26909);
or U27462 (N_27462,N_26614,N_26807);
and U27463 (N_27463,N_26831,N_26566);
xnor U27464 (N_27464,N_26564,N_26668);
nor U27465 (N_27465,N_26666,N_26952);
and U27466 (N_27466,N_26987,N_26725);
nor U27467 (N_27467,N_26739,N_26894);
nor U27468 (N_27468,N_26947,N_26851);
nor U27469 (N_27469,N_26668,N_26964);
nor U27470 (N_27470,N_26898,N_26557);
or U27471 (N_27471,N_26667,N_26519);
nand U27472 (N_27472,N_26954,N_26594);
nor U27473 (N_27473,N_26987,N_26780);
nor U27474 (N_27474,N_26507,N_26915);
nand U27475 (N_27475,N_26798,N_26723);
or U27476 (N_27476,N_26810,N_26560);
or U27477 (N_27477,N_26989,N_26928);
nor U27478 (N_27478,N_26957,N_26501);
or U27479 (N_27479,N_26714,N_26722);
nor U27480 (N_27480,N_26947,N_26768);
nor U27481 (N_27481,N_26585,N_26912);
xnor U27482 (N_27482,N_26790,N_26665);
or U27483 (N_27483,N_26994,N_26957);
xnor U27484 (N_27484,N_26657,N_26786);
nand U27485 (N_27485,N_26828,N_26541);
and U27486 (N_27486,N_26691,N_26660);
nor U27487 (N_27487,N_26519,N_26542);
nor U27488 (N_27488,N_26536,N_26507);
and U27489 (N_27489,N_26934,N_26514);
and U27490 (N_27490,N_26960,N_26665);
xnor U27491 (N_27491,N_26678,N_26953);
nand U27492 (N_27492,N_26640,N_26988);
nor U27493 (N_27493,N_26749,N_26884);
or U27494 (N_27494,N_26891,N_26654);
nor U27495 (N_27495,N_26810,N_26911);
nor U27496 (N_27496,N_26641,N_26524);
nand U27497 (N_27497,N_26769,N_26535);
nand U27498 (N_27498,N_26890,N_26601);
nand U27499 (N_27499,N_26930,N_26735);
xnor U27500 (N_27500,N_27022,N_27199);
and U27501 (N_27501,N_27190,N_27215);
and U27502 (N_27502,N_27276,N_27440);
nor U27503 (N_27503,N_27493,N_27149);
or U27504 (N_27504,N_27317,N_27391);
nand U27505 (N_27505,N_27231,N_27067);
xnor U27506 (N_27506,N_27275,N_27363);
or U27507 (N_27507,N_27433,N_27125);
and U27508 (N_27508,N_27047,N_27128);
nor U27509 (N_27509,N_27112,N_27158);
nand U27510 (N_27510,N_27250,N_27238);
nor U27511 (N_27511,N_27348,N_27173);
xor U27512 (N_27512,N_27123,N_27080);
and U27513 (N_27513,N_27419,N_27027);
nand U27514 (N_27514,N_27380,N_27443);
xor U27515 (N_27515,N_27362,N_27464);
nand U27516 (N_27516,N_27011,N_27498);
nand U27517 (N_27517,N_27437,N_27249);
or U27518 (N_27518,N_27478,N_27079);
and U27519 (N_27519,N_27203,N_27313);
and U27520 (N_27520,N_27485,N_27000);
and U27521 (N_27521,N_27164,N_27182);
nor U27522 (N_27522,N_27188,N_27127);
or U27523 (N_27523,N_27356,N_27017);
and U27524 (N_27524,N_27014,N_27365);
nand U27525 (N_27525,N_27183,N_27427);
nor U27526 (N_27526,N_27179,N_27075);
and U27527 (N_27527,N_27048,N_27445);
and U27528 (N_27528,N_27358,N_27103);
xor U27529 (N_27529,N_27269,N_27018);
or U27530 (N_27530,N_27359,N_27434);
xor U27531 (N_27531,N_27194,N_27052);
nor U27532 (N_27532,N_27056,N_27405);
nor U27533 (N_27533,N_27133,N_27422);
nor U27534 (N_27534,N_27366,N_27452);
nor U27535 (N_27535,N_27344,N_27216);
nor U27536 (N_27536,N_27286,N_27144);
nor U27537 (N_27537,N_27161,N_27071);
nor U27538 (N_27538,N_27432,N_27104);
and U27539 (N_27539,N_27303,N_27092);
and U27540 (N_27540,N_27336,N_27408);
or U27541 (N_27541,N_27007,N_27069);
or U27542 (N_27542,N_27016,N_27438);
and U27543 (N_27543,N_27145,N_27245);
or U27544 (N_27544,N_27113,N_27414);
or U27545 (N_27545,N_27316,N_27187);
nand U27546 (N_27546,N_27480,N_27138);
and U27547 (N_27547,N_27054,N_27415);
nor U27548 (N_27548,N_27255,N_27383);
nor U27549 (N_27549,N_27346,N_27244);
or U27550 (N_27550,N_27428,N_27093);
nor U27551 (N_27551,N_27479,N_27084);
nor U27552 (N_27552,N_27417,N_27451);
xnor U27553 (N_27553,N_27001,N_27390);
nand U27554 (N_27554,N_27354,N_27262);
xor U27555 (N_27555,N_27297,N_27494);
xor U27556 (N_27556,N_27239,N_27219);
nand U27557 (N_27557,N_27483,N_27040);
xnor U27558 (N_27558,N_27287,N_27002);
and U27559 (N_27559,N_27253,N_27025);
xnor U27560 (N_27560,N_27137,N_27270);
and U27561 (N_27561,N_27213,N_27361);
xnor U27562 (N_27562,N_27453,N_27281);
nor U27563 (N_27563,N_27241,N_27473);
and U27564 (N_27564,N_27030,N_27139);
or U27565 (N_27565,N_27311,N_27257);
xnor U27566 (N_27566,N_27264,N_27205);
or U27567 (N_27567,N_27298,N_27246);
nor U27568 (N_27568,N_27094,N_27220);
xor U27569 (N_27569,N_27381,N_27301);
nor U27570 (N_27570,N_27406,N_27459);
and U27571 (N_27571,N_27395,N_27147);
nor U27572 (N_27572,N_27413,N_27468);
or U27573 (N_27573,N_27386,N_27212);
nand U27574 (N_27574,N_27260,N_27055);
xnor U27575 (N_27575,N_27283,N_27095);
nor U27576 (N_27576,N_27321,N_27058);
or U27577 (N_27577,N_27122,N_27057);
or U27578 (N_27578,N_27261,N_27292);
nor U27579 (N_27579,N_27240,N_27198);
and U27580 (N_27580,N_27285,N_27463);
xor U27581 (N_27581,N_27338,N_27349);
and U27582 (N_27582,N_27121,N_27439);
nand U27583 (N_27583,N_27465,N_27259);
xor U27584 (N_27584,N_27117,N_27174);
nand U27585 (N_27585,N_27471,N_27430);
and U27586 (N_27586,N_27177,N_27461);
and U27587 (N_27587,N_27387,N_27475);
and U27588 (N_27588,N_27331,N_27300);
nor U27589 (N_27589,N_27114,N_27252);
nor U27590 (N_27590,N_27063,N_27305);
or U27591 (N_27591,N_27091,N_27169);
nor U27592 (N_27592,N_27446,N_27330);
nor U27593 (N_27593,N_27053,N_27242);
and U27594 (N_27594,N_27120,N_27407);
or U27595 (N_27595,N_27416,N_27102);
nand U27596 (N_27596,N_27211,N_27332);
xor U27597 (N_27597,N_27266,N_27481);
and U27598 (N_27598,N_27009,N_27106);
and U27599 (N_27599,N_27090,N_27491);
or U27600 (N_27600,N_27237,N_27426);
nor U27601 (N_27601,N_27265,N_27150);
nor U27602 (N_27602,N_27031,N_27282);
nand U27603 (N_27603,N_27083,N_27005);
nor U27604 (N_27604,N_27107,N_27455);
and U27605 (N_27605,N_27396,N_27026);
and U27606 (N_27606,N_27312,N_27377);
and U27607 (N_27607,N_27142,N_27327);
or U27608 (N_27608,N_27061,N_27111);
or U27609 (N_27609,N_27289,N_27364);
xor U27610 (N_27610,N_27315,N_27006);
and U27611 (N_27611,N_27319,N_27410);
and U27612 (N_27612,N_27224,N_27490);
nand U27613 (N_27613,N_27448,N_27098);
or U27614 (N_27614,N_27482,N_27489);
xnor U27615 (N_27615,N_27012,N_27256);
and U27616 (N_27616,N_27214,N_27195);
or U27617 (N_27617,N_27068,N_27230);
and U27618 (N_27618,N_27488,N_27207);
or U27619 (N_27619,N_27166,N_27404);
nand U27620 (N_27620,N_27352,N_27134);
xnor U27621 (N_27621,N_27148,N_27372);
nand U27622 (N_27622,N_27236,N_27487);
nor U27623 (N_27623,N_27400,N_27227);
and U27624 (N_27624,N_27254,N_27039);
or U27625 (N_27625,N_27497,N_27099);
and U27626 (N_27626,N_27221,N_27467);
or U27627 (N_27627,N_27288,N_27401);
xor U27628 (N_27628,N_27096,N_27496);
or U27629 (N_27629,N_27458,N_27184);
xnor U27630 (N_27630,N_27167,N_27170);
xor U27631 (N_27631,N_27435,N_27192);
xnor U27632 (N_27632,N_27196,N_27228);
nor U27633 (N_27633,N_27323,N_27029);
or U27634 (N_27634,N_27193,N_27329);
or U27635 (N_27635,N_27476,N_27035);
nand U27636 (N_27636,N_27337,N_27340);
or U27637 (N_27637,N_27100,N_27278);
nor U27638 (N_27638,N_27367,N_27304);
nand U27639 (N_27639,N_27412,N_27004);
nand U27640 (N_27640,N_27146,N_27105);
nand U27641 (N_27641,N_27036,N_27399);
nor U27642 (N_27642,N_27424,N_27389);
nand U27643 (N_27643,N_27347,N_27333);
xor U27644 (N_27644,N_27339,N_27234);
nor U27645 (N_27645,N_27020,N_27232);
nor U27646 (N_27646,N_27155,N_27351);
or U27647 (N_27647,N_27308,N_27322);
nand U27648 (N_27648,N_27402,N_27457);
nor U27649 (N_27649,N_27073,N_27101);
and U27650 (N_27650,N_27124,N_27420);
xor U27651 (N_27651,N_27041,N_27126);
or U27652 (N_27652,N_27157,N_27248);
and U27653 (N_27653,N_27397,N_27225);
or U27654 (N_27654,N_27046,N_27409);
or U27655 (N_27655,N_27411,N_27165);
or U27656 (N_27656,N_27119,N_27484);
nor U27657 (N_27657,N_27388,N_27328);
nand U27658 (N_27658,N_27447,N_27129);
nand U27659 (N_27659,N_27038,N_27431);
or U27660 (N_27660,N_27243,N_27015);
or U27661 (N_27661,N_27066,N_27291);
and U27662 (N_27662,N_27076,N_27325);
xor U27663 (N_27663,N_27210,N_27206);
xor U27664 (N_27664,N_27293,N_27175);
or U27665 (N_27665,N_27176,N_27049);
nand U27666 (N_27666,N_27044,N_27074);
xor U27667 (N_27667,N_27217,N_27403);
nand U27668 (N_27668,N_27136,N_27070);
xnor U27669 (N_27669,N_27109,N_27191);
xor U27670 (N_27670,N_27472,N_27263);
nand U27671 (N_27671,N_27394,N_27486);
or U27672 (N_27672,N_27460,N_27097);
xnor U27673 (N_27673,N_27385,N_27171);
xor U27674 (N_27674,N_27296,N_27318);
and U27675 (N_27675,N_27274,N_27115);
nand U27676 (N_27676,N_27462,N_27421);
and U27677 (N_27677,N_27280,N_27172);
nor U27678 (N_27678,N_27268,N_27130);
xnor U27679 (N_27679,N_27226,N_27392);
nor U27680 (N_27680,N_27143,N_27131);
nand U27681 (N_27681,N_27369,N_27309);
and U27682 (N_27682,N_27118,N_27449);
and U27683 (N_27683,N_27202,N_27425);
and U27684 (N_27684,N_27051,N_27334);
nor U27685 (N_27685,N_27023,N_27222);
or U27686 (N_27686,N_27087,N_27272);
and U27687 (N_27687,N_27082,N_27444);
nor U27688 (N_27688,N_27477,N_27470);
or U27689 (N_27689,N_27186,N_27258);
nand U27690 (N_27690,N_27441,N_27353);
and U27691 (N_27691,N_27163,N_27132);
or U27692 (N_27692,N_27078,N_27034);
and U27693 (N_27693,N_27373,N_27060);
nor U27694 (N_27694,N_27368,N_27469);
nand U27695 (N_27695,N_27350,N_27159);
and U27696 (N_27696,N_27492,N_27277);
and U27697 (N_27697,N_27156,N_27357);
xor U27698 (N_27698,N_27065,N_27279);
xnor U27699 (N_27699,N_27466,N_27162);
xor U27700 (N_27700,N_27152,N_27062);
nand U27701 (N_27701,N_27375,N_27178);
nand U27702 (N_27702,N_27393,N_27341);
or U27703 (N_27703,N_27181,N_27335);
xor U27704 (N_27704,N_27233,N_27379);
and U27705 (N_27705,N_27010,N_27085);
and U27706 (N_27706,N_27324,N_27450);
or U27707 (N_27707,N_27037,N_27108);
nand U27708 (N_27708,N_27294,N_27306);
or U27709 (N_27709,N_27495,N_27442);
and U27710 (N_27710,N_27271,N_27081);
or U27711 (N_27711,N_27345,N_27343);
nor U27712 (N_27712,N_27140,N_27429);
and U27713 (N_27713,N_27474,N_27045);
nor U27714 (N_27714,N_27378,N_27021);
and U27715 (N_27715,N_27185,N_27355);
xor U27716 (N_27716,N_27374,N_27032);
xnor U27717 (N_27717,N_27326,N_27423);
and U27718 (N_27718,N_27135,N_27003);
and U27719 (N_27719,N_27314,N_27376);
and U27720 (N_27720,N_27043,N_27189);
or U27721 (N_27721,N_27295,N_27008);
nor U27722 (N_27722,N_27360,N_27310);
or U27723 (N_27723,N_27072,N_27371);
nor U27724 (N_27724,N_27168,N_27382);
nor U27725 (N_27725,N_27370,N_27418);
nor U27726 (N_27726,N_27064,N_27086);
xnor U27727 (N_27727,N_27019,N_27251);
nor U27728 (N_27728,N_27160,N_27208);
xnor U27729 (N_27729,N_27436,N_27267);
nand U27730 (N_27730,N_27059,N_27110);
nor U27731 (N_27731,N_27307,N_27151);
or U27732 (N_27732,N_27384,N_27499);
nand U27733 (N_27733,N_27398,N_27223);
nor U27734 (N_27734,N_27302,N_27284);
xor U27735 (N_27735,N_27273,N_27229);
or U27736 (N_27736,N_27042,N_27200);
nand U27737 (N_27737,N_27201,N_27320);
and U27738 (N_27738,N_27050,N_27141);
nand U27739 (N_27739,N_27013,N_27089);
and U27740 (N_27740,N_27456,N_27290);
or U27741 (N_27741,N_27454,N_27204);
xnor U27742 (N_27742,N_27028,N_27299);
and U27743 (N_27743,N_27209,N_27218);
xnor U27744 (N_27744,N_27180,N_27154);
and U27745 (N_27745,N_27235,N_27197);
nand U27746 (N_27746,N_27088,N_27033);
nand U27747 (N_27747,N_27077,N_27153);
xor U27748 (N_27748,N_27342,N_27024);
or U27749 (N_27749,N_27116,N_27247);
nor U27750 (N_27750,N_27028,N_27174);
xor U27751 (N_27751,N_27300,N_27178);
nor U27752 (N_27752,N_27331,N_27384);
or U27753 (N_27753,N_27447,N_27444);
nor U27754 (N_27754,N_27086,N_27486);
or U27755 (N_27755,N_27479,N_27073);
nand U27756 (N_27756,N_27315,N_27090);
xor U27757 (N_27757,N_27108,N_27130);
and U27758 (N_27758,N_27412,N_27041);
and U27759 (N_27759,N_27149,N_27204);
or U27760 (N_27760,N_27176,N_27263);
or U27761 (N_27761,N_27422,N_27401);
xnor U27762 (N_27762,N_27080,N_27345);
nor U27763 (N_27763,N_27148,N_27397);
nand U27764 (N_27764,N_27362,N_27432);
and U27765 (N_27765,N_27218,N_27034);
nor U27766 (N_27766,N_27028,N_27340);
and U27767 (N_27767,N_27182,N_27244);
and U27768 (N_27768,N_27017,N_27364);
or U27769 (N_27769,N_27039,N_27317);
and U27770 (N_27770,N_27369,N_27045);
nor U27771 (N_27771,N_27042,N_27243);
and U27772 (N_27772,N_27133,N_27185);
and U27773 (N_27773,N_27221,N_27139);
nand U27774 (N_27774,N_27197,N_27404);
and U27775 (N_27775,N_27236,N_27141);
and U27776 (N_27776,N_27170,N_27107);
and U27777 (N_27777,N_27308,N_27459);
or U27778 (N_27778,N_27433,N_27348);
and U27779 (N_27779,N_27466,N_27251);
nand U27780 (N_27780,N_27039,N_27306);
and U27781 (N_27781,N_27194,N_27406);
and U27782 (N_27782,N_27428,N_27094);
or U27783 (N_27783,N_27342,N_27015);
nand U27784 (N_27784,N_27079,N_27440);
xnor U27785 (N_27785,N_27169,N_27485);
nor U27786 (N_27786,N_27151,N_27273);
or U27787 (N_27787,N_27351,N_27160);
or U27788 (N_27788,N_27254,N_27107);
xnor U27789 (N_27789,N_27144,N_27250);
nand U27790 (N_27790,N_27168,N_27357);
nand U27791 (N_27791,N_27076,N_27128);
or U27792 (N_27792,N_27317,N_27427);
nor U27793 (N_27793,N_27142,N_27216);
nor U27794 (N_27794,N_27177,N_27334);
and U27795 (N_27795,N_27498,N_27229);
xor U27796 (N_27796,N_27286,N_27352);
and U27797 (N_27797,N_27273,N_27042);
nand U27798 (N_27798,N_27239,N_27399);
or U27799 (N_27799,N_27006,N_27488);
nor U27800 (N_27800,N_27316,N_27158);
or U27801 (N_27801,N_27304,N_27462);
nor U27802 (N_27802,N_27211,N_27033);
or U27803 (N_27803,N_27110,N_27115);
nand U27804 (N_27804,N_27194,N_27150);
or U27805 (N_27805,N_27010,N_27443);
xnor U27806 (N_27806,N_27353,N_27132);
nand U27807 (N_27807,N_27474,N_27264);
xnor U27808 (N_27808,N_27042,N_27210);
and U27809 (N_27809,N_27288,N_27045);
nand U27810 (N_27810,N_27087,N_27292);
nor U27811 (N_27811,N_27117,N_27027);
nand U27812 (N_27812,N_27475,N_27252);
nor U27813 (N_27813,N_27000,N_27295);
or U27814 (N_27814,N_27354,N_27353);
xor U27815 (N_27815,N_27006,N_27358);
xor U27816 (N_27816,N_27354,N_27438);
nand U27817 (N_27817,N_27112,N_27200);
nand U27818 (N_27818,N_27010,N_27226);
or U27819 (N_27819,N_27140,N_27043);
or U27820 (N_27820,N_27385,N_27437);
nor U27821 (N_27821,N_27171,N_27429);
nor U27822 (N_27822,N_27095,N_27042);
xnor U27823 (N_27823,N_27449,N_27366);
nor U27824 (N_27824,N_27308,N_27001);
nand U27825 (N_27825,N_27139,N_27201);
xor U27826 (N_27826,N_27295,N_27298);
and U27827 (N_27827,N_27042,N_27110);
nor U27828 (N_27828,N_27284,N_27013);
xor U27829 (N_27829,N_27467,N_27110);
or U27830 (N_27830,N_27482,N_27466);
or U27831 (N_27831,N_27445,N_27243);
and U27832 (N_27832,N_27097,N_27360);
or U27833 (N_27833,N_27309,N_27354);
or U27834 (N_27834,N_27106,N_27121);
and U27835 (N_27835,N_27324,N_27048);
xor U27836 (N_27836,N_27494,N_27187);
xor U27837 (N_27837,N_27348,N_27331);
nor U27838 (N_27838,N_27084,N_27346);
xor U27839 (N_27839,N_27480,N_27043);
and U27840 (N_27840,N_27324,N_27396);
and U27841 (N_27841,N_27282,N_27106);
and U27842 (N_27842,N_27404,N_27002);
and U27843 (N_27843,N_27065,N_27293);
nand U27844 (N_27844,N_27437,N_27271);
xor U27845 (N_27845,N_27215,N_27245);
or U27846 (N_27846,N_27018,N_27412);
or U27847 (N_27847,N_27396,N_27241);
or U27848 (N_27848,N_27293,N_27130);
xor U27849 (N_27849,N_27017,N_27319);
nor U27850 (N_27850,N_27228,N_27244);
or U27851 (N_27851,N_27488,N_27003);
nor U27852 (N_27852,N_27490,N_27269);
nand U27853 (N_27853,N_27490,N_27201);
xor U27854 (N_27854,N_27428,N_27037);
nand U27855 (N_27855,N_27252,N_27016);
xor U27856 (N_27856,N_27314,N_27013);
or U27857 (N_27857,N_27283,N_27202);
or U27858 (N_27858,N_27395,N_27193);
or U27859 (N_27859,N_27122,N_27475);
or U27860 (N_27860,N_27238,N_27099);
nor U27861 (N_27861,N_27284,N_27419);
nor U27862 (N_27862,N_27116,N_27314);
xor U27863 (N_27863,N_27084,N_27014);
and U27864 (N_27864,N_27261,N_27056);
xor U27865 (N_27865,N_27246,N_27487);
xnor U27866 (N_27866,N_27196,N_27494);
xor U27867 (N_27867,N_27091,N_27402);
nand U27868 (N_27868,N_27177,N_27048);
or U27869 (N_27869,N_27385,N_27458);
nand U27870 (N_27870,N_27054,N_27371);
xor U27871 (N_27871,N_27414,N_27260);
nand U27872 (N_27872,N_27011,N_27374);
nor U27873 (N_27873,N_27126,N_27455);
xnor U27874 (N_27874,N_27206,N_27240);
nor U27875 (N_27875,N_27401,N_27113);
nor U27876 (N_27876,N_27088,N_27454);
and U27877 (N_27877,N_27291,N_27426);
nand U27878 (N_27878,N_27165,N_27121);
nor U27879 (N_27879,N_27364,N_27408);
or U27880 (N_27880,N_27472,N_27180);
or U27881 (N_27881,N_27134,N_27496);
nor U27882 (N_27882,N_27058,N_27193);
and U27883 (N_27883,N_27173,N_27460);
nand U27884 (N_27884,N_27075,N_27443);
and U27885 (N_27885,N_27032,N_27294);
or U27886 (N_27886,N_27300,N_27160);
nor U27887 (N_27887,N_27137,N_27240);
nand U27888 (N_27888,N_27426,N_27008);
or U27889 (N_27889,N_27245,N_27129);
nor U27890 (N_27890,N_27413,N_27145);
nor U27891 (N_27891,N_27248,N_27116);
and U27892 (N_27892,N_27009,N_27304);
or U27893 (N_27893,N_27381,N_27163);
nand U27894 (N_27894,N_27337,N_27169);
nor U27895 (N_27895,N_27037,N_27459);
nor U27896 (N_27896,N_27062,N_27090);
and U27897 (N_27897,N_27404,N_27265);
xor U27898 (N_27898,N_27157,N_27017);
and U27899 (N_27899,N_27035,N_27382);
nand U27900 (N_27900,N_27186,N_27115);
nor U27901 (N_27901,N_27086,N_27495);
or U27902 (N_27902,N_27260,N_27353);
and U27903 (N_27903,N_27191,N_27272);
xnor U27904 (N_27904,N_27129,N_27088);
nand U27905 (N_27905,N_27305,N_27024);
nand U27906 (N_27906,N_27201,N_27138);
or U27907 (N_27907,N_27106,N_27460);
nor U27908 (N_27908,N_27486,N_27234);
nand U27909 (N_27909,N_27051,N_27018);
nand U27910 (N_27910,N_27164,N_27462);
nand U27911 (N_27911,N_27288,N_27213);
nor U27912 (N_27912,N_27262,N_27135);
xnor U27913 (N_27913,N_27060,N_27087);
and U27914 (N_27914,N_27263,N_27108);
and U27915 (N_27915,N_27156,N_27064);
xnor U27916 (N_27916,N_27002,N_27073);
and U27917 (N_27917,N_27373,N_27009);
nand U27918 (N_27918,N_27167,N_27438);
nand U27919 (N_27919,N_27167,N_27078);
xnor U27920 (N_27920,N_27037,N_27383);
nor U27921 (N_27921,N_27166,N_27476);
xor U27922 (N_27922,N_27190,N_27007);
and U27923 (N_27923,N_27357,N_27166);
nor U27924 (N_27924,N_27161,N_27285);
nor U27925 (N_27925,N_27485,N_27492);
xnor U27926 (N_27926,N_27323,N_27119);
xor U27927 (N_27927,N_27212,N_27220);
xor U27928 (N_27928,N_27220,N_27354);
or U27929 (N_27929,N_27465,N_27338);
xor U27930 (N_27930,N_27444,N_27440);
xnor U27931 (N_27931,N_27380,N_27058);
and U27932 (N_27932,N_27087,N_27099);
xnor U27933 (N_27933,N_27067,N_27140);
nor U27934 (N_27934,N_27485,N_27105);
nand U27935 (N_27935,N_27286,N_27479);
nor U27936 (N_27936,N_27090,N_27197);
or U27937 (N_27937,N_27172,N_27259);
xnor U27938 (N_27938,N_27208,N_27415);
xor U27939 (N_27939,N_27465,N_27360);
xnor U27940 (N_27940,N_27418,N_27207);
and U27941 (N_27941,N_27421,N_27410);
xnor U27942 (N_27942,N_27271,N_27204);
nand U27943 (N_27943,N_27062,N_27142);
and U27944 (N_27944,N_27053,N_27481);
xor U27945 (N_27945,N_27313,N_27151);
xor U27946 (N_27946,N_27426,N_27231);
nor U27947 (N_27947,N_27086,N_27179);
xor U27948 (N_27948,N_27399,N_27269);
nor U27949 (N_27949,N_27122,N_27300);
xor U27950 (N_27950,N_27480,N_27159);
and U27951 (N_27951,N_27353,N_27430);
nor U27952 (N_27952,N_27331,N_27204);
xor U27953 (N_27953,N_27112,N_27264);
or U27954 (N_27954,N_27285,N_27223);
nor U27955 (N_27955,N_27417,N_27360);
nand U27956 (N_27956,N_27041,N_27136);
nor U27957 (N_27957,N_27019,N_27344);
nor U27958 (N_27958,N_27070,N_27486);
nand U27959 (N_27959,N_27410,N_27067);
and U27960 (N_27960,N_27227,N_27106);
or U27961 (N_27961,N_27242,N_27240);
and U27962 (N_27962,N_27118,N_27493);
and U27963 (N_27963,N_27004,N_27276);
nand U27964 (N_27964,N_27194,N_27408);
or U27965 (N_27965,N_27106,N_27425);
nand U27966 (N_27966,N_27301,N_27484);
and U27967 (N_27967,N_27295,N_27285);
xor U27968 (N_27968,N_27445,N_27375);
xnor U27969 (N_27969,N_27182,N_27480);
nand U27970 (N_27970,N_27469,N_27463);
xnor U27971 (N_27971,N_27076,N_27021);
and U27972 (N_27972,N_27107,N_27410);
xnor U27973 (N_27973,N_27222,N_27455);
xor U27974 (N_27974,N_27081,N_27372);
and U27975 (N_27975,N_27098,N_27126);
nand U27976 (N_27976,N_27002,N_27133);
nor U27977 (N_27977,N_27114,N_27393);
or U27978 (N_27978,N_27169,N_27181);
or U27979 (N_27979,N_27348,N_27349);
nor U27980 (N_27980,N_27219,N_27193);
and U27981 (N_27981,N_27003,N_27078);
xnor U27982 (N_27982,N_27049,N_27328);
and U27983 (N_27983,N_27468,N_27081);
or U27984 (N_27984,N_27415,N_27487);
nand U27985 (N_27985,N_27141,N_27403);
nor U27986 (N_27986,N_27162,N_27457);
xnor U27987 (N_27987,N_27127,N_27176);
nor U27988 (N_27988,N_27116,N_27305);
or U27989 (N_27989,N_27286,N_27194);
nor U27990 (N_27990,N_27358,N_27059);
xnor U27991 (N_27991,N_27485,N_27402);
xor U27992 (N_27992,N_27132,N_27198);
or U27993 (N_27993,N_27018,N_27182);
and U27994 (N_27994,N_27382,N_27449);
xnor U27995 (N_27995,N_27102,N_27267);
nor U27996 (N_27996,N_27411,N_27005);
nor U27997 (N_27997,N_27411,N_27447);
or U27998 (N_27998,N_27288,N_27462);
nand U27999 (N_27999,N_27147,N_27266);
nor U28000 (N_28000,N_27894,N_27580);
nor U28001 (N_28001,N_27596,N_27540);
and U28002 (N_28002,N_27880,N_27778);
and U28003 (N_28003,N_27742,N_27845);
or U28004 (N_28004,N_27825,N_27747);
or U28005 (N_28005,N_27775,N_27895);
and U28006 (N_28006,N_27565,N_27854);
and U28007 (N_28007,N_27952,N_27502);
nand U28008 (N_28008,N_27641,N_27792);
and U28009 (N_28009,N_27759,N_27917);
nor U28010 (N_28010,N_27713,N_27719);
xnor U28011 (N_28011,N_27616,N_27663);
xor U28012 (N_28012,N_27909,N_27798);
or U28013 (N_28013,N_27509,N_27701);
and U28014 (N_28014,N_27762,N_27769);
xor U28015 (N_28015,N_27715,N_27910);
and U28016 (N_28016,N_27939,N_27964);
nand U28017 (N_28017,N_27853,N_27805);
and U28018 (N_28018,N_27730,N_27693);
nor U28019 (N_28019,N_27623,N_27525);
or U28020 (N_28020,N_27878,N_27501);
nand U28021 (N_28021,N_27500,N_27735);
or U28022 (N_28022,N_27632,N_27832);
xnor U28023 (N_28023,N_27947,N_27538);
and U28024 (N_28024,N_27506,N_27593);
nor U28025 (N_28025,N_27619,N_27757);
nand U28026 (N_28026,N_27599,N_27592);
nor U28027 (N_28027,N_27691,N_27667);
xnor U28028 (N_28028,N_27652,N_27557);
and U28029 (N_28029,N_27718,N_27709);
or U28030 (N_28030,N_27626,N_27521);
nor U28031 (N_28031,N_27914,N_27886);
and U28032 (N_28032,N_27546,N_27885);
or U28033 (N_28033,N_27806,N_27802);
nand U28034 (N_28034,N_27508,N_27631);
xnor U28035 (N_28035,N_27793,N_27949);
nand U28036 (N_28036,N_27927,N_27651);
nor U28037 (N_28037,N_27916,N_27660);
xnor U28038 (N_28038,N_27512,N_27669);
nand U28039 (N_28039,N_27714,N_27530);
and U28040 (N_28040,N_27789,N_27563);
nand U28041 (N_28041,N_27955,N_27847);
nand U28042 (N_28042,N_27956,N_27542);
nand U28043 (N_28043,N_27911,N_27970);
or U28044 (N_28044,N_27884,N_27865);
or U28045 (N_28045,N_27566,N_27581);
nand U28046 (N_28046,N_27639,N_27923);
nand U28047 (N_28047,N_27570,N_27782);
nor U28048 (N_28048,N_27823,N_27680);
and U28049 (N_28049,N_27649,N_27737);
nand U28050 (N_28050,N_27932,N_27594);
or U28051 (N_28051,N_27934,N_27564);
and U28052 (N_28052,N_27533,N_27888);
nor U28053 (N_28053,N_27846,N_27803);
and U28054 (N_28054,N_27905,N_27582);
xnor U28055 (N_28055,N_27658,N_27867);
nor U28056 (N_28056,N_27527,N_27951);
xor U28057 (N_28057,N_27962,N_27813);
nand U28058 (N_28058,N_27796,N_27568);
or U28059 (N_28059,N_27705,N_27583);
xnor U28060 (N_28060,N_27943,N_27835);
or U28061 (N_28061,N_27824,N_27598);
xor U28062 (N_28062,N_27958,N_27627);
and U28063 (N_28063,N_27859,N_27842);
nor U28064 (N_28064,N_27768,N_27694);
and U28065 (N_28065,N_27586,N_27706);
nand U28066 (N_28066,N_27812,N_27901);
nand U28067 (N_28067,N_27689,N_27942);
and U28068 (N_28068,N_27703,N_27666);
xnor U28069 (N_28069,N_27961,N_27863);
nor U28070 (N_28070,N_27595,N_27821);
or U28071 (N_28071,N_27673,N_27638);
nand U28072 (N_28072,N_27571,N_27869);
xor U28073 (N_28073,N_27969,N_27868);
and U28074 (N_28074,N_27553,N_27558);
and U28075 (N_28075,N_27817,N_27839);
nor U28076 (N_28076,N_27556,N_27918);
nand U28077 (N_28077,N_27588,N_27975);
nor U28078 (N_28078,N_27562,N_27881);
or U28079 (N_28079,N_27618,N_27681);
nand U28080 (N_28080,N_27721,N_27576);
or U28081 (N_28081,N_27851,N_27785);
xnor U28082 (N_28082,N_27944,N_27702);
nor U28083 (N_28083,N_27860,N_27953);
and U28084 (N_28084,N_27931,N_27620);
nor U28085 (N_28085,N_27629,N_27797);
or U28086 (N_28086,N_27840,N_27763);
or U28087 (N_28087,N_27892,N_27528);
and U28088 (N_28088,N_27809,N_27552);
or U28089 (N_28089,N_27799,N_27532);
nor U28090 (N_28090,N_27684,N_27606);
nand U28091 (N_28091,N_27993,N_27904);
nor U28092 (N_28092,N_27624,N_27529);
nor U28093 (N_28093,N_27725,N_27536);
nand U28094 (N_28094,N_27539,N_27643);
and U28095 (N_28095,N_27991,N_27729);
xor U28096 (N_28096,N_27661,N_27779);
xnor U28097 (N_28097,N_27848,N_27692);
nor U28098 (N_28098,N_27541,N_27994);
nor U28099 (N_28099,N_27511,N_27555);
xor U28100 (N_28100,N_27781,N_27928);
nand U28101 (N_28101,N_27731,N_27844);
or U28102 (N_28102,N_27996,N_27740);
xnor U28103 (N_28103,N_27516,N_27647);
xor U28104 (N_28104,N_27985,N_27526);
xor U28105 (N_28105,N_27834,N_27548);
xnor U28106 (N_28106,N_27872,N_27518);
or U28107 (N_28107,N_27941,N_27987);
nor U28108 (N_28108,N_27976,N_27788);
xnor U28109 (N_28109,N_27707,N_27800);
nor U28110 (N_28110,N_27773,N_27831);
nor U28111 (N_28111,N_27610,N_27889);
nor U28112 (N_28112,N_27621,N_27977);
nor U28113 (N_28113,N_27810,N_27611);
or U28114 (N_28114,N_27640,N_27561);
and U28115 (N_28115,N_27790,N_27559);
xnor U28116 (N_28116,N_27929,N_27676);
and U28117 (N_28117,N_27843,N_27664);
nor U28118 (N_28118,N_27816,N_27672);
nand U28119 (N_28119,N_27601,N_27791);
nand U28120 (N_28120,N_27613,N_27567);
xor U28121 (N_28121,N_27732,N_27874);
xnor U28122 (N_28122,N_27883,N_27890);
nor U28123 (N_28123,N_27551,N_27711);
or U28124 (N_28124,N_27671,N_27897);
nor U28125 (N_28125,N_27899,N_27836);
nor U28126 (N_28126,N_27614,N_27534);
nor U28127 (N_28127,N_27877,N_27830);
nand U28128 (N_28128,N_27630,N_27745);
or U28129 (N_28129,N_27900,N_27907);
and U28130 (N_28130,N_27504,N_27645);
xor U28131 (N_28131,N_27723,N_27537);
and U28132 (N_28132,N_27891,N_27515);
nand U28133 (N_28133,N_27544,N_27770);
or U28134 (N_28134,N_27764,N_27675);
nor U28135 (N_28135,N_27695,N_27980);
nand U28136 (N_28136,N_27841,N_27677);
and U28137 (N_28137,N_27655,N_27815);
xnor U28138 (N_28138,N_27690,N_27688);
or U28139 (N_28139,N_27925,N_27820);
nor U28140 (N_28140,N_27653,N_27746);
xnor U28141 (N_28141,N_27879,N_27963);
nand U28142 (N_28142,N_27849,N_27524);
xnor U28143 (N_28143,N_27995,N_27650);
and U28144 (N_28144,N_27654,N_27972);
nor U28145 (N_28145,N_27744,N_27600);
xor U28146 (N_28146,N_27968,N_27887);
nor U28147 (N_28147,N_27876,N_27992);
xnor U28148 (N_28148,N_27716,N_27607);
nand U28149 (N_28149,N_27545,N_27922);
xnor U28150 (N_28150,N_27870,N_27862);
nor U28151 (N_28151,N_27808,N_27999);
nor U28152 (N_28152,N_27998,N_27902);
xor U28153 (N_28153,N_27728,N_27549);
or U28154 (N_28154,N_27828,N_27678);
nand U28155 (N_28155,N_27748,N_27893);
xor U28156 (N_28156,N_27578,N_27979);
or U28157 (N_28157,N_27665,N_27915);
xor U28158 (N_28158,N_27615,N_27531);
nor U28159 (N_28159,N_27698,N_27628);
nor U28160 (N_28160,N_27858,N_27741);
and U28161 (N_28161,N_27726,N_27818);
xnor U28162 (N_28162,N_27967,N_27605);
nand U28163 (N_28163,N_27777,N_27749);
nor U28164 (N_28164,N_27736,N_27882);
nand U28165 (N_28165,N_27560,N_27924);
or U28166 (N_28166,N_27520,N_27717);
nand U28167 (N_28167,N_27722,N_27896);
nand U28168 (N_28168,N_27786,N_27753);
nor U28169 (N_28169,N_27503,N_27523);
nor U28170 (N_28170,N_27783,N_27751);
and U28171 (N_28171,N_27871,N_27829);
or U28172 (N_28172,N_27683,N_27966);
or U28173 (N_28173,N_27569,N_27597);
nand U28174 (N_28174,N_27724,N_27921);
or U28175 (N_28175,N_27866,N_27855);
and U28176 (N_28176,N_27982,N_27852);
nor U28177 (N_28177,N_27959,N_27700);
xnor U28178 (N_28178,N_27765,N_27756);
and U28179 (N_28179,N_27513,N_27838);
nor U28180 (N_28180,N_27644,N_27755);
and U28181 (N_28181,N_27981,N_27873);
nor U28182 (N_28182,N_27656,N_27648);
xor U28183 (N_28183,N_27794,N_27760);
nor U28184 (N_28184,N_27990,N_27609);
nor U28185 (N_28185,N_27575,N_27752);
nor U28186 (N_28186,N_27633,N_27602);
or U28187 (N_28187,N_27795,N_27585);
nor U28188 (N_28188,N_27517,N_27819);
or U28189 (N_28189,N_27584,N_27804);
or U28190 (N_28190,N_27727,N_27510);
xor U28191 (N_28191,N_27543,N_27739);
nand U28192 (N_28192,N_27974,N_27761);
nor U28193 (N_28193,N_27950,N_27612);
nor U28194 (N_28194,N_27634,N_27903);
xor U28195 (N_28195,N_27906,N_27772);
nor U28196 (N_28196,N_27674,N_27668);
nand U28197 (N_28197,N_27784,N_27935);
and U28198 (N_28198,N_27590,N_27547);
xor U28199 (N_28199,N_27938,N_27919);
nand U28200 (N_28200,N_27734,N_27573);
nor U28201 (N_28201,N_27637,N_27807);
nor U28202 (N_28202,N_27965,N_27774);
or U28203 (N_28203,N_27926,N_27603);
nor U28204 (N_28204,N_27940,N_27697);
nor U28205 (N_28205,N_27948,N_27933);
and U28206 (N_28206,N_27720,N_27591);
nor U28207 (N_28207,N_27936,N_27913);
and U28208 (N_28208,N_27930,N_27507);
nand U28209 (N_28209,N_27758,N_27780);
nand U28210 (N_28210,N_27687,N_27635);
or U28211 (N_28211,N_27801,N_27642);
or U28212 (N_28212,N_27577,N_27657);
xor U28213 (N_28213,N_27646,N_27945);
xor U28214 (N_28214,N_27814,N_27861);
nand U28215 (N_28215,N_27754,N_27875);
xor U28216 (N_28216,N_27946,N_27983);
or U28217 (N_28217,N_27986,N_27898);
xnor U28218 (N_28218,N_27771,N_27957);
or U28219 (N_28219,N_27554,N_27522);
and U28220 (N_28220,N_27954,N_27750);
nor U28221 (N_28221,N_27685,N_27837);
nor U28222 (N_28222,N_27589,N_27579);
and U28223 (N_28223,N_27997,N_27514);
or U28224 (N_28224,N_27574,N_27710);
xnor U28225 (N_28225,N_27960,N_27822);
nor U28226 (N_28226,N_27827,N_27622);
and U28227 (N_28227,N_27587,N_27712);
nor U28228 (N_28228,N_27662,N_27519);
or U28229 (N_28229,N_27978,N_27696);
or U28230 (N_28230,N_27686,N_27550);
and U28231 (N_28231,N_27973,N_27833);
or U28232 (N_28232,N_27811,N_27787);
nor U28233 (N_28233,N_27708,N_27733);
and U28234 (N_28234,N_27617,N_27670);
or U28235 (N_28235,N_27738,N_27776);
nand U28236 (N_28236,N_27984,N_27767);
xnor U28237 (N_28237,N_27625,N_27608);
nor U28238 (N_28238,N_27912,N_27699);
nand U28239 (N_28239,N_27857,N_27971);
or U28240 (N_28240,N_27850,N_27766);
nand U28241 (N_28241,N_27679,N_27920);
xnor U28242 (N_28242,N_27989,N_27743);
nand U28243 (N_28243,N_27659,N_27604);
xnor U28244 (N_28244,N_27682,N_27704);
nor U28245 (N_28245,N_27572,N_27908);
or U28246 (N_28246,N_27826,N_27937);
or U28247 (N_28247,N_27864,N_27535);
and U28248 (N_28248,N_27988,N_27856);
xor U28249 (N_28249,N_27505,N_27636);
nand U28250 (N_28250,N_27806,N_27912);
or U28251 (N_28251,N_27876,N_27677);
nand U28252 (N_28252,N_27564,N_27843);
or U28253 (N_28253,N_27677,N_27962);
or U28254 (N_28254,N_27802,N_27914);
or U28255 (N_28255,N_27703,N_27969);
or U28256 (N_28256,N_27773,N_27500);
and U28257 (N_28257,N_27581,N_27954);
and U28258 (N_28258,N_27995,N_27652);
nand U28259 (N_28259,N_27729,N_27606);
or U28260 (N_28260,N_27712,N_27870);
nand U28261 (N_28261,N_27834,N_27636);
nand U28262 (N_28262,N_27982,N_27722);
and U28263 (N_28263,N_27794,N_27652);
nand U28264 (N_28264,N_27934,N_27704);
xnor U28265 (N_28265,N_27666,N_27717);
or U28266 (N_28266,N_27558,N_27939);
nor U28267 (N_28267,N_27616,N_27597);
nor U28268 (N_28268,N_27569,N_27826);
xnor U28269 (N_28269,N_27747,N_27751);
xor U28270 (N_28270,N_27613,N_27820);
nand U28271 (N_28271,N_27661,N_27763);
nand U28272 (N_28272,N_27733,N_27513);
xnor U28273 (N_28273,N_27776,N_27797);
nand U28274 (N_28274,N_27539,N_27633);
and U28275 (N_28275,N_27566,N_27649);
nand U28276 (N_28276,N_27594,N_27993);
nor U28277 (N_28277,N_27942,N_27877);
xnor U28278 (N_28278,N_27982,N_27931);
nand U28279 (N_28279,N_27963,N_27628);
nor U28280 (N_28280,N_27907,N_27722);
nor U28281 (N_28281,N_27704,N_27526);
xor U28282 (N_28282,N_27721,N_27619);
or U28283 (N_28283,N_27990,N_27867);
xor U28284 (N_28284,N_27738,N_27868);
xnor U28285 (N_28285,N_27953,N_27586);
nor U28286 (N_28286,N_27687,N_27797);
nand U28287 (N_28287,N_27808,N_27939);
and U28288 (N_28288,N_27841,N_27600);
or U28289 (N_28289,N_27943,N_27649);
nor U28290 (N_28290,N_27539,N_27937);
nor U28291 (N_28291,N_27972,N_27537);
or U28292 (N_28292,N_27811,N_27674);
nor U28293 (N_28293,N_27905,N_27725);
and U28294 (N_28294,N_27885,N_27810);
nor U28295 (N_28295,N_27844,N_27918);
or U28296 (N_28296,N_27935,N_27778);
xor U28297 (N_28297,N_27550,N_27871);
xnor U28298 (N_28298,N_27690,N_27680);
nand U28299 (N_28299,N_27887,N_27639);
nor U28300 (N_28300,N_27777,N_27506);
nand U28301 (N_28301,N_27859,N_27907);
nand U28302 (N_28302,N_27584,N_27614);
xor U28303 (N_28303,N_27620,N_27782);
and U28304 (N_28304,N_27554,N_27747);
nor U28305 (N_28305,N_27759,N_27536);
nand U28306 (N_28306,N_27685,N_27663);
nand U28307 (N_28307,N_27905,N_27871);
and U28308 (N_28308,N_27640,N_27990);
or U28309 (N_28309,N_27587,N_27669);
xor U28310 (N_28310,N_27632,N_27741);
nand U28311 (N_28311,N_27958,N_27969);
nor U28312 (N_28312,N_27746,N_27517);
nand U28313 (N_28313,N_27763,N_27714);
xnor U28314 (N_28314,N_27909,N_27808);
xnor U28315 (N_28315,N_27845,N_27771);
or U28316 (N_28316,N_27780,N_27565);
or U28317 (N_28317,N_27634,N_27875);
nand U28318 (N_28318,N_27904,N_27891);
nor U28319 (N_28319,N_27722,N_27991);
xnor U28320 (N_28320,N_27640,N_27519);
and U28321 (N_28321,N_27725,N_27745);
xnor U28322 (N_28322,N_27622,N_27929);
and U28323 (N_28323,N_27597,N_27629);
and U28324 (N_28324,N_27597,N_27879);
nor U28325 (N_28325,N_27710,N_27649);
or U28326 (N_28326,N_27999,N_27893);
nor U28327 (N_28327,N_27908,N_27737);
nor U28328 (N_28328,N_27545,N_27772);
nand U28329 (N_28329,N_27825,N_27794);
nor U28330 (N_28330,N_27598,N_27819);
or U28331 (N_28331,N_27909,N_27816);
xnor U28332 (N_28332,N_27959,N_27912);
xor U28333 (N_28333,N_27559,N_27899);
nor U28334 (N_28334,N_27548,N_27600);
xor U28335 (N_28335,N_27666,N_27587);
xnor U28336 (N_28336,N_27646,N_27502);
xor U28337 (N_28337,N_27518,N_27751);
or U28338 (N_28338,N_27769,N_27960);
nor U28339 (N_28339,N_27881,N_27580);
or U28340 (N_28340,N_27614,N_27990);
and U28341 (N_28341,N_27745,N_27583);
xor U28342 (N_28342,N_27976,N_27692);
xor U28343 (N_28343,N_27978,N_27827);
xnor U28344 (N_28344,N_27749,N_27960);
or U28345 (N_28345,N_27851,N_27674);
xnor U28346 (N_28346,N_27537,N_27912);
or U28347 (N_28347,N_27720,N_27877);
or U28348 (N_28348,N_27947,N_27640);
nor U28349 (N_28349,N_27503,N_27644);
or U28350 (N_28350,N_27835,N_27746);
or U28351 (N_28351,N_27693,N_27506);
and U28352 (N_28352,N_27883,N_27548);
nand U28353 (N_28353,N_27547,N_27902);
or U28354 (N_28354,N_27661,N_27884);
xnor U28355 (N_28355,N_27817,N_27621);
xnor U28356 (N_28356,N_27533,N_27856);
or U28357 (N_28357,N_27637,N_27665);
or U28358 (N_28358,N_27729,N_27709);
nand U28359 (N_28359,N_27770,N_27933);
and U28360 (N_28360,N_27819,N_27633);
and U28361 (N_28361,N_27850,N_27573);
nand U28362 (N_28362,N_27608,N_27563);
xor U28363 (N_28363,N_27702,N_27657);
xnor U28364 (N_28364,N_27981,N_27588);
and U28365 (N_28365,N_27952,N_27608);
and U28366 (N_28366,N_27658,N_27605);
nand U28367 (N_28367,N_27793,N_27857);
nand U28368 (N_28368,N_27777,N_27926);
or U28369 (N_28369,N_27942,N_27578);
and U28370 (N_28370,N_27508,N_27583);
nand U28371 (N_28371,N_27666,N_27828);
xor U28372 (N_28372,N_27928,N_27677);
xor U28373 (N_28373,N_27694,N_27935);
nand U28374 (N_28374,N_27549,N_27526);
or U28375 (N_28375,N_27912,N_27546);
or U28376 (N_28376,N_27708,N_27956);
nand U28377 (N_28377,N_27591,N_27830);
nor U28378 (N_28378,N_27672,N_27555);
nor U28379 (N_28379,N_27925,N_27963);
nor U28380 (N_28380,N_27768,N_27515);
or U28381 (N_28381,N_27579,N_27640);
xor U28382 (N_28382,N_27787,N_27795);
or U28383 (N_28383,N_27954,N_27828);
nor U28384 (N_28384,N_27700,N_27806);
and U28385 (N_28385,N_27782,N_27538);
and U28386 (N_28386,N_27906,N_27540);
and U28387 (N_28387,N_27799,N_27631);
or U28388 (N_28388,N_27622,N_27995);
and U28389 (N_28389,N_27927,N_27758);
xor U28390 (N_28390,N_27834,N_27615);
and U28391 (N_28391,N_27622,N_27872);
or U28392 (N_28392,N_27933,N_27816);
xnor U28393 (N_28393,N_27775,N_27999);
nor U28394 (N_28394,N_27634,N_27602);
nor U28395 (N_28395,N_27617,N_27708);
or U28396 (N_28396,N_27941,N_27750);
nand U28397 (N_28397,N_27502,N_27734);
xor U28398 (N_28398,N_27756,N_27593);
xnor U28399 (N_28399,N_27767,N_27776);
and U28400 (N_28400,N_27588,N_27693);
nand U28401 (N_28401,N_27610,N_27609);
nand U28402 (N_28402,N_27949,N_27792);
or U28403 (N_28403,N_27941,N_27741);
and U28404 (N_28404,N_27628,N_27568);
nor U28405 (N_28405,N_27746,N_27885);
nor U28406 (N_28406,N_27949,N_27691);
nand U28407 (N_28407,N_27612,N_27896);
or U28408 (N_28408,N_27566,N_27940);
and U28409 (N_28409,N_27778,N_27731);
nand U28410 (N_28410,N_27941,N_27564);
nor U28411 (N_28411,N_27644,N_27759);
nor U28412 (N_28412,N_27503,N_27802);
xnor U28413 (N_28413,N_27773,N_27987);
or U28414 (N_28414,N_27632,N_27700);
nand U28415 (N_28415,N_27601,N_27885);
xor U28416 (N_28416,N_27748,N_27882);
xnor U28417 (N_28417,N_27891,N_27965);
or U28418 (N_28418,N_27760,N_27714);
and U28419 (N_28419,N_27928,N_27807);
nor U28420 (N_28420,N_27813,N_27670);
nor U28421 (N_28421,N_27831,N_27969);
xor U28422 (N_28422,N_27600,N_27799);
nand U28423 (N_28423,N_27718,N_27508);
or U28424 (N_28424,N_27967,N_27582);
and U28425 (N_28425,N_27704,N_27699);
nor U28426 (N_28426,N_27888,N_27819);
nand U28427 (N_28427,N_27511,N_27771);
nor U28428 (N_28428,N_27793,N_27743);
xnor U28429 (N_28429,N_27711,N_27655);
nor U28430 (N_28430,N_27540,N_27744);
or U28431 (N_28431,N_27796,N_27944);
and U28432 (N_28432,N_27945,N_27934);
or U28433 (N_28433,N_27594,N_27598);
xnor U28434 (N_28434,N_27910,N_27638);
or U28435 (N_28435,N_27564,N_27755);
and U28436 (N_28436,N_27518,N_27635);
xor U28437 (N_28437,N_27872,N_27799);
nand U28438 (N_28438,N_27524,N_27994);
or U28439 (N_28439,N_27722,N_27604);
nor U28440 (N_28440,N_27700,N_27525);
or U28441 (N_28441,N_27767,N_27620);
nand U28442 (N_28442,N_27567,N_27950);
xnor U28443 (N_28443,N_27580,N_27649);
nor U28444 (N_28444,N_27904,N_27728);
and U28445 (N_28445,N_27600,N_27856);
nor U28446 (N_28446,N_27617,N_27795);
and U28447 (N_28447,N_27864,N_27792);
or U28448 (N_28448,N_27612,N_27751);
nand U28449 (N_28449,N_27963,N_27589);
nor U28450 (N_28450,N_27681,N_27623);
nand U28451 (N_28451,N_27893,N_27730);
and U28452 (N_28452,N_27960,N_27939);
nor U28453 (N_28453,N_27925,N_27686);
and U28454 (N_28454,N_27689,N_27810);
nor U28455 (N_28455,N_27890,N_27545);
nor U28456 (N_28456,N_27589,N_27516);
or U28457 (N_28457,N_27906,N_27695);
nand U28458 (N_28458,N_27514,N_27942);
or U28459 (N_28459,N_27676,N_27579);
and U28460 (N_28460,N_27691,N_27851);
or U28461 (N_28461,N_27961,N_27991);
and U28462 (N_28462,N_27943,N_27961);
nand U28463 (N_28463,N_27842,N_27535);
nand U28464 (N_28464,N_27946,N_27764);
and U28465 (N_28465,N_27903,N_27980);
nand U28466 (N_28466,N_27966,N_27553);
and U28467 (N_28467,N_27669,N_27693);
and U28468 (N_28468,N_27712,N_27656);
or U28469 (N_28469,N_27645,N_27933);
and U28470 (N_28470,N_27701,N_27625);
and U28471 (N_28471,N_27695,N_27583);
nor U28472 (N_28472,N_27862,N_27868);
nor U28473 (N_28473,N_27930,N_27608);
nand U28474 (N_28474,N_27946,N_27712);
xor U28475 (N_28475,N_27792,N_27505);
nand U28476 (N_28476,N_27584,N_27705);
nand U28477 (N_28477,N_27925,N_27680);
or U28478 (N_28478,N_27662,N_27768);
or U28479 (N_28479,N_27840,N_27762);
nor U28480 (N_28480,N_27560,N_27658);
nand U28481 (N_28481,N_27749,N_27898);
xnor U28482 (N_28482,N_27777,N_27866);
nand U28483 (N_28483,N_27805,N_27877);
nand U28484 (N_28484,N_27634,N_27534);
or U28485 (N_28485,N_27541,N_27672);
and U28486 (N_28486,N_27588,N_27554);
or U28487 (N_28487,N_27835,N_27571);
or U28488 (N_28488,N_27977,N_27647);
and U28489 (N_28489,N_27538,N_27774);
xor U28490 (N_28490,N_27505,N_27816);
xnor U28491 (N_28491,N_27827,N_27722);
and U28492 (N_28492,N_27983,N_27858);
xor U28493 (N_28493,N_27887,N_27807);
nand U28494 (N_28494,N_27914,N_27955);
xnor U28495 (N_28495,N_27692,N_27525);
nand U28496 (N_28496,N_27975,N_27679);
or U28497 (N_28497,N_27969,N_27737);
xnor U28498 (N_28498,N_27516,N_27788);
nand U28499 (N_28499,N_27600,N_27894);
and U28500 (N_28500,N_28266,N_28460);
and U28501 (N_28501,N_28434,N_28011);
nor U28502 (N_28502,N_28202,N_28335);
nand U28503 (N_28503,N_28171,N_28096);
nand U28504 (N_28504,N_28341,N_28254);
nor U28505 (N_28505,N_28264,N_28483);
or U28506 (N_28506,N_28403,N_28122);
and U28507 (N_28507,N_28091,N_28253);
or U28508 (N_28508,N_28380,N_28466);
nand U28509 (N_28509,N_28092,N_28265);
and U28510 (N_28510,N_28182,N_28411);
xnor U28511 (N_28511,N_28159,N_28248);
nand U28512 (N_28512,N_28414,N_28377);
xnor U28513 (N_28513,N_28062,N_28222);
or U28514 (N_28514,N_28018,N_28493);
or U28515 (N_28515,N_28427,N_28256);
and U28516 (N_28516,N_28196,N_28086);
nand U28517 (N_28517,N_28119,N_28170);
or U28518 (N_28518,N_28418,N_28213);
nand U28519 (N_28519,N_28234,N_28140);
nand U28520 (N_28520,N_28218,N_28349);
or U28521 (N_28521,N_28481,N_28039);
or U28522 (N_28522,N_28142,N_28429);
xor U28523 (N_28523,N_28157,N_28004);
nor U28524 (N_28524,N_28195,N_28278);
and U28525 (N_28525,N_28371,N_28391);
and U28526 (N_28526,N_28022,N_28121);
nand U28527 (N_28527,N_28058,N_28310);
nor U28528 (N_28528,N_28276,N_28442);
and U28529 (N_28529,N_28361,N_28387);
nand U28530 (N_28530,N_28488,N_28379);
and U28531 (N_28531,N_28472,N_28072);
and U28532 (N_28532,N_28482,N_28409);
and U28533 (N_28533,N_28107,N_28273);
and U28534 (N_28534,N_28238,N_28325);
nand U28535 (N_28535,N_28315,N_28005);
nand U28536 (N_28536,N_28372,N_28324);
xnor U28537 (N_28537,N_28164,N_28223);
nor U28538 (N_28538,N_28211,N_28279);
and U28539 (N_28539,N_28158,N_28436);
xnor U28540 (N_28540,N_28048,N_28024);
nand U28541 (N_28541,N_28282,N_28149);
nor U28542 (N_28542,N_28113,N_28464);
and U28543 (N_28543,N_28413,N_28351);
nand U28544 (N_28544,N_28255,N_28165);
nor U28545 (N_28545,N_28305,N_28304);
or U28546 (N_28546,N_28449,N_28212);
nor U28547 (N_28547,N_28428,N_28098);
xor U28548 (N_28548,N_28071,N_28032);
nor U28549 (N_28549,N_28154,N_28246);
or U28550 (N_28550,N_28152,N_28221);
and U28551 (N_28551,N_28043,N_28247);
nand U28552 (N_28552,N_28283,N_28134);
or U28553 (N_28553,N_28061,N_28399);
and U28554 (N_28554,N_28344,N_28003);
or U28555 (N_28555,N_28240,N_28068);
nand U28556 (N_28556,N_28063,N_28451);
nand U28557 (N_28557,N_28366,N_28210);
xnor U28558 (N_28558,N_28095,N_28023);
and U28559 (N_28559,N_28016,N_28345);
nand U28560 (N_28560,N_28186,N_28079);
nor U28561 (N_28561,N_28307,N_28026);
nor U28562 (N_28562,N_28469,N_28497);
xnor U28563 (N_28563,N_28178,N_28357);
xor U28564 (N_28564,N_28360,N_28020);
or U28565 (N_28565,N_28089,N_28342);
xnor U28566 (N_28566,N_28476,N_28373);
or U28567 (N_28567,N_28130,N_28285);
and U28568 (N_28568,N_28350,N_28495);
nand U28569 (N_28569,N_28271,N_28115);
nand U28570 (N_28570,N_28274,N_28289);
nand U28571 (N_28571,N_28475,N_28419);
or U28572 (N_28572,N_28425,N_28463);
or U28573 (N_28573,N_28309,N_28124);
xnor U28574 (N_28574,N_28067,N_28146);
nand U28575 (N_28575,N_28394,N_28204);
nand U28576 (N_28576,N_28287,N_28090);
nor U28577 (N_28577,N_28284,N_28433);
nand U28578 (N_28578,N_28006,N_28027);
nor U28579 (N_28579,N_28487,N_28021);
or U28580 (N_28580,N_28491,N_28192);
or U28581 (N_28581,N_28249,N_28454);
and U28582 (N_28582,N_28462,N_28015);
and U28583 (N_28583,N_28423,N_28199);
or U28584 (N_28584,N_28311,N_28225);
xnor U28585 (N_28585,N_28384,N_28161);
nand U28586 (N_28586,N_28480,N_28106);
and U28587 (N_28587,N_28431,N_28314);
and U28588 (N_28588,N_28336,N_28382);
nor U28589 (N_28589,N_28406,N_28236);
and U28590 (N_28590,N_28037,N_28343);
and U28591 (N_28591,N_28308,N_28293);
or U28592 (N_28592,N_28331,N_28147);
nand U28593 (N_28593,N_28070,N_28041);
xnor U28594 (N_28594,N_28185,N_28028);
and U28595 (N_28595,N_28370,N_28458);
nor U28596 (N_28596,N_28494,N_28328);
or U28597 (N_28597,N_28174,N_28395);
xor U28598 (N_28598,N_28286,N_28390);
xor U28599 (N_28599,N_28132,N_28054);
nand U28600 (N_28600,N_28378,N_28139);
nor U28601 (N_28601,N_28337,N_28323);
nand U28602 (N_28602,N_28381,N_28258);
or U28603 (N_28603,N_28486,N_28045);
xnor U28604 (N_28604,N_28228,N_28319);
and U28605 (N_28605,N_28208,N_28322);
nand U28606 (N_28606,N_28239,N_28127);
xor U28607 (N_28607,N_28321,N_28422);
xor U28608 (N_28608,N_28330,N_28261);
xor U28609 (N_28609,N_28153,N_28402);
and U28610 (N_28610,N_28160,N_28053);
nor U28611 (N_28611,N_28137,N_28009);
and U28612 (N_28612,N_28117,N_28346);
xnor U28613 (N_28613,N_28201,N_28272);
nor U28614 (N_28614,N_28415,N_28112);
nand U28615 (N_28615,N_28155,N_28465);
and U28616 (N_28616,N_28232,N_28446);
nor U28617 (N_28617,N_28299,N_28468);
nor U28618 (N_28618,N_28224,N_28320);
nand U28619 (N_28619,N_28099,N_28440);
nand U28620 (N_28620,N_28268,N_28038);
nand U28621 (N_28621,N_28363,N_28455);
or U28622 (N_28622,N_28163,N_28338);
nor U28623 (N_28623,N_28367,N_28435);
nor U28624 (N_28624,N_28209,N_28181);
nand U28625 (N_28625,N_28456,N_28355);
or U28626 (N_28626,N_28243,N_28241);
nand U28627 (N_28627,N_28097,N_28025);
nand U28628 (N_28628,N_28252,N_28471);
xor U28629 (N_28629,N_28417,N_28128);
nor U28630 (N_28630,N_28148,N_28441);
and U28631 (N_28631,N_28369,N_28110);
nand U28632 (N_28632,N_28162,N_28051);
and U28633 (N_28633,N_28376,N_28049);
nor U28634 (N_28634,N_28180,N_28206);
xnor U28635 (N_28635,N_28275,N_28059);
nor U28636 (N_28636,N_28060,N_28075);
xor U28637 (N_28637,N_28042,N_28150);
or U28638 (N_28638,N_28116,N_28100);
nand U28639 (N_28639,N_28453,N_28281);
and U28640 (N_28640,N_28074,N_28136);
or U28641 (N_28641,N_28479,N_28392);
and U28642 (N_28642,N_28297,N_28034);
xor U28643 (N_28643,N_28359,N_28404);
xor U28644 (N_28644,N_28292,N_28229);
and U28645 (N_28645,N_28069,N_28470);
xnor U28646 (N_28646,N_28104,N_28296);
nand U28647 (N_28647,N_28242,N_28401);
and U28648 (N_28648,N_28093,N_28010);
nand U28649 (N_28649,N_28172,N_28105);
and U28650 (N_28650,N_28416,N_28393);
nor U28651 (N_28651,N_28030,N_28179);
xnor U28652 (N_28652,N_28076,N_28078);
and U28653 (N_28653,N_28151,N_28033);
and U28654 (N_28654,N_28250,N_28303);
nand U28655 (N_28655,N_28013,N_28398);
or U28656 (N_28656,N_28467,N_28012);
or U28657 (N_28657,N_28088,N_28101);
or U28658 (N_28658,N_28044,N_28126);
nor U28659 (N_28659,N_28187,N_28114);
or U28660 (N_28660,N_28167,N_28014);
nor U28661 (N_28661,N_28191,N_28216);
nand U28662 (N_28662,N_28207,N_28365);
nor U28663 (N_28663,N_28189,N_28430);
nor U28664 (N_28664,N_28019,N_28008);
xnor U28665 (N_28665,N_28348,N_28040);
nand U28666 (N_28666,N_28329,N_28368);
xnor U28667 (N_28667,N_28485,N_28347);
xor U28668 (N_28668,N_28017,N_28235);
and U28669 (N_28669,N_28461,N_28318);
or U28670 (N_28670,N_28144,N_28388);
or U28671 (N_28671,N_28439,N_28103);
xor U28672 (N_28672,N_28452,N_28400);
nor U28673 (N_28673,N_28002,N_28490);
nor U28674 (N_28674,N_28405,N_28197);
xor U28675 (N_28675,N_28169,N_28364);
nor U28676 (N_28676,N_28007,N_28385);
and U28677 (N_28677,N_28001,N_28190);
or U28678 (N_28678,N_28220,N_28295);
nor U28679 (N_28679,N_28410,N_28362);
xor U28680 (N_28680,N_28291,N_28496);
and U28681 (N_28681,N_28300,N_28492);
nand U28682 (N_28682,N_28407,N_28141);
and U28683 (N_28683,N_28437,N_28358);
nor U28684 (N_28684,N_28133,N_28447);
or U28685 (N_28685,N_28035,N_28432);
or U28686 (N_28686,N_28166,N_28082);
nor U28687 (N_28687,N_28031,N_28029);
and U28688 (N_28688,N_28156,N_28135);
nor U28689 (N_28689,N_28257,N_28176);
xnor U28690 (N_28690,N_28263,N_28484);
and U28691 (N_28691,N_28109,N_28374);
or U28692 (N_28692,N_28226,N_28056);
nand U28693 (N_28693,N_28237,N_28052);
and U28694 (N_28694,N_28177,N_28397);
and U28695 (N_28695,N_28094,N_28084);
nand U28696 (N_28696,N_28233,N_28129);
and U28697 (N_28697,N_28443,N_28474);
or U28698 (N_28698,N_28267,N_28260);
or U28699 (N_28699,N_28064,N_28057);
nand U28700 (N_28700,N_28083,N_28298);
and U28701 (N_28701,N_28420,N_28175);
xnor U28702 (N_28702,N_28389,N_28200);
xor U28703 (N_28703,N_28230,N_28294);
nand U28704 (N_28704,N_28473,N_28426);
or U28705 (N_28705,N_28312,N_28073);
nand U28706 (N_28706,N_28087,N_28219);
xnor U28707 (N_28707,N_28280,N_28339);
nor U28708 (N_28708,N_28316,N_28332);
nand U28709 (N_28709,N_28194,N_28408);
nand U28710 (N_28710,N_28356,N_28244);
and U28711 (N_28711,N_28077,N_28111);
xnor U28712 (N_28712,N_28173,N_28055);
and U28713 (N_28713,N_28340,N_28489);
xnor U28714 (N_28714,N_28424,N_28326);
and U28715 (N_28715,N_28448,N_28459);
xnor U28716 (N_28716,N_28193,N_28145);
and U28717 (N_28717,N_28386,N_28270);
xnor U28718 (N_28718,N_28217,N_28198);
and U28719 (N_28719,N_28333,N_28450);
xnor U28720 (N_28720,N_28102,N_28353);
xor U28721 (N_28721,N_28066,N_28231);
or U28722 (N_28722,N_28203,N_28445);
nor U28723 (N_28723,N_28036,N_28050);
nor U28724 (N_28724,N_28227,N_28131);
and U28725 (N_28725,N_28215,N_28138);
nand U28726 (N_28726,N_28000,N_28245);
xnor U28727 (N_28727,N_28205,N_28269);
nor U28728 (N_28728,N_28498,N_28184);
and U28729 (N_28729,N_28188,N_28444);
nor U28730 (N_28730,N_28327,N_28065);
xnor U28731 (N_28731,N_28125,N_28168);
nand U28732 (N_28732,N_28047,N_28457);
nor U28733 (N_28733,N_28302,N_28499);
nand U28734 (N_28734,N_28313,N_28108);
xor U28735 (N_28735,N_28046,N_28354);
and U28736 (N_28736,N_28334,N_28396);
nor U28737 (N_28737,N_28214,N_28383);
xor U28738 (N_28738,N_28478,N_28120);
nor U28739 (N_28739,N_28123,N_28262);
nand U28740 (N_28740,N_28080,N_28412);
nand U28741 (N_28741,N_28375,N_28143);
xor U28742 (N_28742,N_28352,N_28290);
xnor U28743 (N_28743,N_28301,N_28251);
xor U28744 (N_28744,N_28081,N_28438);
xnor U28745 (N_28745,N_28288,N_28085);
nand U28746 (N_28746,N_28259,N_28277);
and U28747 (N_28747,N_28317,N_28306);
and U28748 (N_28748,N_28118,N_28421);
or U28749 (N_28749,N_28183,N_28477);
or U28750 (N_28750,N_28484,N_28186);
nand U28751 (N_28751,N_28210,N_28420);
nand U28752 (N_28752,N_28070,N_28272);
and U28753 (N_28753,N_28363,N_28094);
nand U28754 (N_28754,N_28029,N_28439);
or U28755 (N_28755,N_28096,N_28154);
and U28756 (N_28756,N_28388,N_28357);
and U28757 (N_28757,N_28372,N_28472);
nor U28758 (N_28758,N_28365,N_28265);
xnor U28759 (N_28759,N_28463,N_28138);
and U28760 (N_28760,N_28162,N_28387);
nand U28761 (N_28761,N_28459,N_28455);
xor U28762 (N_28762,N_28032,N_28368);
nand U28763 (N_28763,N_28423,N_28036);
or U28764 (N_28764,N_28477,N_28310);
xnor U28765 (N_28765,N_28196,N_28191);
or U28766 (N_28766,N_28196,N_28484);
nand U28767 (N_28767,N_28067,N_28312);
or U28768 (N_28768,N_28446,N_28135);
or U28769 (N_28769,N_28040,N_28086);
xnor U28770 (N_28770,N_28218,N_28364);
and U28771 (N_28771,N_28220,N_28406);
nor U28772 (N_28772,N_28498,N_28347);
nand U28773 (N_28773,N_28034,N_28011);
or U28774 (N_28774,N_28438,N_28128);
nand U28775 (N_28775,N_28056,N_28469);
and U28776 (N_28776,N_28377,N_28141);
and U28777 (N_28777,N_28179,N_28320);
nor U28778 (N_28778,N_28312,N_28392);
xnor U28779 (N_28779,N_28293,N_28412);
nor U28780 (N_28780,N_28498,N_28181);
or U28781 (N_28781,N_28084,N_28397);
nand U28782 (N_28782,N_28329,N_28104);
nand U28783 (N_28783,N_28163,N_28006);
nand U28784 (N_28784,N_28339,N_28229);
and U28785 (N_28785,N_28391,N_28049);
and U28786 (N_28786,N_28352,N_28348);
or U28787 (N_28787,N_28419,N_28449);
nor U28788 (N_28788,N_28361,N_28277);
and U28789 (N_28789,N_28246,N_28212);
or U28790 (N_28790,N_28424,N_28139);
nor U28791 (N_28791,N_28312,N_28352);
and U28792 (N_28792,N_28352,N_28116);
xor U28793 (N_28793,N_28221,N_28399);
nor U28794 (N_28794,N_28306,N_28496);
nand U28795 (N_28795,N_28118,N_28432);
xnor U28796 (N_28796,N_28428,N_28492);
or U28797 (N_28797,N_28251,N_28077);
nor U28798 (N_28798,N_28057,N_28424);
and U28799 (N_28799,N_28283,N_28070);
or U28800 (N_28800,N_28414,N_28265);
nor U28801 (N_28801,N_28010,N_28487);
or U28802 (N_28802,N_28100,N_28165);
nand U28803 (N_28803,N_28296,N_28279);
nor U28804 (N_28804,N_28042,N_28304);
or U28805 (N_28805,N_28014,N_28020);
nor U28806 (N_28806,N_28243,N_28365);
nand U28807 (N_28807,N_28032,N_28272);
nor U28808 (N_28808,N_28350,N_28147);
nand U28809 (N_28809,N_28263,N_28360);
nor U28810 (N_28810,N_28119,N_28123);
nor U28811 (N_28811,N_28119,N_28143);
and U28812 (N_28812,N_28188,N_28238);
nand U28813 (N_28813,N_28046,N_28251);
and U28814 (N_28814,N_28185,N_28361);
xnor U28815 (N_28815,N_28340,N_28320);
or U28816 (N_28816,N_28404,N_28169);
nand U28817 (N_28817,N_28331,N_28192);
nor U28818 (N_28818,N_28110,N_28416);
and U28819 (N_28819,N_28393,N_28491);
and U28820 (N_28820,N_28332,N_28386);
xor U28821 (N_28821,N_28121,N_28228);
nor U28822 (N_28822,N_28407,N_28294);
and U28823 (N_28823,N_28464,N_28268);
and U28824 (N_28824,N_28294,N_28034);
nor U28825 (N_28825,N_28011,N_28026);
and U28826 (N_28826,N_28477,N_28387);
nand U28827 (N_28827,N_28251,N_28461);
nor U28828 (N_28828,N_28342,N_28087);
nor U28829 (N_28829,N_28236,N_28409);
and U28830 (N_28830,N_28154,N_28296);
or U28831 (N_28831,N_28434,N_28424);
and U28832 (N_28832,N_28188,N_28001);
nand U28833 (N_28833,N_28076,N_28061);
and U28834 (N_28834,N_28429,N_28091);
nor U28835 (N_28835,N_28029,N_28075);
or U28836 (N_28836,N_28110,N_28083);
nor U28837 (N_28837,N_28202,N_28201);
and U28838 (N_28838,N_28103,N_28461);
nand U28839 (N_28839,N_28076,N_28454);
nor U28840 (N_28840,N_28473,N_28498);
or U28841 (N_28841,N_28133,N_28370);
nand U28842 (N_28842,N_28270,N_28496);
or U28843 (N_28843,N_28440,N_28489);
or U28844 (N_28844,N_28323,N_28099);
or U28845 (N_28845,N_28119,N_28067);
nor U28846 (N_28846,N_28125,N_28050);
nand U28847 (N_28847,N_28468,N_28087);
nand U28848 (N_28848,N_28075,N_28492);
or U28849 (N_28849,N_28320,N_28140);
nor U28850 (N_28850,N_28088,N_28295);
nor U28851 (N_28851,N_28265,N_28089);
nor U28852 (N_28852,N_28089,N_28199);
and U28853 (N_28853,N_28121,N_28434);
nor U28854 (N_28854,N_28374,N_28193);
xor U28855 (N_28855,N_28342,N_28361);
xor U28856 (N_28856,N_28314,N_28126);
or U28857 (N_28857,N_28496,N_28185);
xnor U28858 (N_28858,N_28426,N_28394);
and U28859 (N_28859,N_28191,N_28385);
xor U28860 (N_28860,N_28212,N_28026);
and U28861 (N_28861,N_28023,N_28479);
or U28862 (N_28862,N_28285,N_28004);
and U28863 (N_28863,N_28365,N_28126);
or U28864 (N_28864,N_28350,N_28202);
or U28865 (N_28865,N_28380,N_28177);
nand U28866 (N_28866,N_28392,N_28481);
nor U28867 (N_28867,N_28371,N_28007);
or U28868 (N_28868,N_28160,N_28245);
nor U28869 (N_28869,N_28053,N_28263);
xnor U28870 (N_28870,N_28487,N_28262);
xnor U28871 (N_28871,N_28304,N_28054);
nor U28872 (N_28872,N_28489,N_28039);
xor U28873 (N_28873,N_28467,N_28124);
nor U28874 (N_28874,N_28234,N_28472);
and U28875 (N_28875,N_28441,N_28422);
nand U28876 (N_28876,N_28433,N_28145);
xnor U28877 (N_28877,N_28264,N_28271);
or U28878 (N_28878,N_28344,N_28396);
or U28879 (N_28879,N_28069,N_28317);
nand U28880 (N_28880,N_28149,N_28269);
and U28881 (N_28881,N_28360,N_28066);
xor U28882 (N_28882,N_28174,N_28350);
xor U28883 (N_28883,N_28096,N_28366);
nor U28884 (N_28884,N_28353,N_28143);
or U28885 (N_28885,N_28308,N_28135);
and U28886 (N_28886,N_28386,N_28357);
nand U28887 (N_28887,N_28283,N_28191);
nand U28888 (N_28888,N_28207,N_28385);
nor U28889 (N_28889,N_28025,N_28103);
nor U28890 (N_28890,N_28168,N_28163);
nand U28891 (N_28891,N_28233,N_28423);
nand U28892 (N_28892,N_28468,N_28446);
nor U28893 (N_28893,N_28283,N_28417);
nor U28894 (N_28894,N_28470,N_28400);
xnor U28895 (N_28895,N_28294,N_28080);
xor U28896 (N_28896,N_28294,N_28495);
nor U28897 (N_28897,N_28364,N_28459);
xnor U28898 (N_28898,N_28262,N_28117);
and U28899 (N_28899,N_28151,N_28416);
nor U28900 (N_28900,N_28011,N_28390);
or U28901 (N_28901,N_28290,N_28415);
xor U28902 (N_28902,N_28140,N_28278);
and U28903 (N_28903,N_28374,N_28322);
nand U28904 (N_28904,N_28197,N_28441);
and U28905 (N_28905,N_28137,N_28388);
xnor U28906 (N_28906,N_28430,N_28376);
or U28907 (N_28907,N_28058,N_28065);
nand U28908 (N_28908,N_28064,N_28153);
nand U28909 (N_28909,N_28261,N_28361);
nor U28910 (N_28910,N_28251,N_28303);
nor U28911 (N_28911,N_28030,N_28053);
or U28912 (N_28912,N_28124,N_28115);
nor U28913 (N_28913,N_28419,N_28457);
xor U28914 (N_28914,N_28383,N_28426);
or U28915 (N_28915,N_28043,N_28116);
and U28916 (N_28916,N_28445,N_28095);
and U28917 (N_28917,N_28232,N_28340);
nor U28918 (N_28918,N_28141,N_28165);
and U28919 (N_28919,N_28477,N_28320);
xnor U28920 (N_28920,N_28303,N_28307);
or U28921 (N_28921,N_28364,N_28481);
nor U28922 (N_28922,N_28468,N_28099);
nor U28923 (N_28923,N_28389,N_28490);
or U28924 (N_28924,N_28147,N_28165);
and U28925 (N_28925,N_28158,N_28070);
and U28926 (N_28926,N_28376,N_28042);
xnor U28927 (N_28927,N_28132,N_28333);
or U28928 (N_28928,N_28203,N_28266);
or U28929 (N_28929,N_28292,N_28107);
xnor U28930 (N_28930,N_28283,N_28463);
or U28931 (N_28931,N_28302,N_28133);
and U28932 (N_28932,N_28289,N_28043);
nor U28933 (N_28933,N_28236,N_28390);
and U28934 (N_28934,N_28263,N_28167);
nand U28935 (N_28935,N_28080,N_28263);
nor U28936 (N_28936,N_28242,N_28186);
nand U28937 (N_28937,N_28209,N_28289);
or U28938 (N_28938,N_28114,N_28242);
nand U28939 (N_28939,N_28086,N_28463);
nor U28940 (N_28940,N_28243,N_28162);
xor U28941 (N_28941,N_28103,N_28435);
and U28942 (N_28942,N_28169,N_28379);
nor U28943 (N_28943,N_28317,N_28360);
or U28944 (N_28944,N_28092,N_28138);
and U28945 (N_28945,N_28292,N_28363);
and U28946 (N_28946,N_28033,N_28325);
and U28947 (N_28947,N_28469,N_28365);
nor U28948 (N_28948,N_28274,N_28187);
or U28949 (N_28949,N_28241,N_28292);
xnor U28950 (N_28950,N_28142,N_28159);
nor U28951 (N_28951,N_28245,N_28357);
nand U28952 (N_28952,N_28480,N_28152);
and U28953 (N_28953,N_28179,N_28250);
nand U28954 (N_28954,N_28427,N_28109);
nand U28955 (N_28955,N_28123,N_28453);
nor U28956 (N_28956,N_28036,N_28086);
nand U28957 (N_28957,N_28073,N_28108);
and U28958 (N_28958,N_28397,N_28440);
nor U28959 (N_28959,N_28435,N_28473);
and U28960 (N_28960,N_28022,N_28357);
nand U28961 (N_28961,N_28117,N_28111);
xnor U28962 (N_28962,N_28093,N_28267);
xor U28963 (N_28963,N_28241,N_28165);
xor U28964 (N_28964,N_28322,N_28350);
nor U28965 (N_28965,N_28475,N_28152);
xnor U28966 (N_28966,N_28018,N_28420);
nand U28967 (N_28967,N_28082,N_28473);
nor U28968 (N_28968,N_28351,N_28320);
nor U28969 (N_28969,N_28356,N_28450);
nor U28970 (N_28970,N_28174,N_28457);
xnor U28971 (N_28971,N_28304,N_28410);
and U28972 (N_28972,N_28450,N_28019);
nor U28973 (N_28973,N_28436,N_28287);
xnor U28974 (N_28974,N_28066,N_28344);
and U28975 (N_28975,N_28461,N_28396);
or U28976 (N_28976,N_28197,N_28416);
or U28977 (N_28977,N_28183,N_28153);
nand U28978 (N_28978,N_28241,N_28426);
nor U28979 (N_28979,N_28171,N_28015);
xor U28980 (N_28980,N_28133,N_28162);
nand U28981 (N_28981,N_28281,N_28031);
and U28982 (N_28982,N_28396,N_28127);
and U28983 (N_28983,N_28252,N_28288);
nor U28984 (N_28984,N_28316,N_28302);
or U28985 (N_28985,N_28264,N_28002);
xor U28986 (N_28986,N_28410,N_28490);
and U28987 (N_28987,N_28220,N_28262);
nor U28988 (N_28988,N_28135,N_28492);
xnor U28989 (N_28989,N_28363,N_28214);
or U28990 (N_28990,N_28232,N_28017);
or U28991 (N_28991,N_28118,N_28368);
and U28992 (N_28992,N_28405,N_28121);
xor U28993 (N_28993,N_28454,N_28321);
and U28994 (N_28994,N_28140,N_28391);
xor U28995 (N_28995,N_28048,N_28300);
nand U28996 (N_28996,N_28237,N_28169);
nor U28997 (N_28997,N_28443,N_28012);
xor U28998 (N_28998,N_28304,N_28148);
nand U28999 (N_28999,N_28455,N_28208);
nor U29000 (N_29000,N_28545,N_28745);
nor U29001 (N_29001,N_28721,N_28844);
xnor U29002 (N_29002,N_28589,N_28794);
nand U29003 (N_29003,N_28725,N_28920);
nor U29004 (N_29004,N_28879,N_28703);
or U29005 (N_29005,N_28840,N_28740);
nand U29006 (N_29006,N_28551,N_28549);
xnor U29007 (N_29007,N_28859,N_28623);
and U29008 (N_29008,N_28510,N_28702);
or U29009 (N_29009,N_28601,N_28747);
xor U29010 (N_29010,N_28641,N_28704);
nand U29011 (N_29011,N_28916,N_28946);
nand U29012 (N_29012,N_28961,N_28507);
nand U29013 (N_29013,N_28887,N_28811);
and U29014 (N_29014,N_28959,N_28850);
nor U29015 (N_29015,N_28791,N_28627);
and U29016 (N_29016,N_28554,N_28588);
or U29017 (N_29017,N_28636,N_28829);
or U29018 (N_29018,N_28754,N_28683);
nor U29019 (N_29019,N_28854,N_28712);
and U29020 (N_29020,N_28790,N_28518);
xor U29021 (N_29021,N_28918,N_28985);
nand U29022 (N_29022,N_28528,N_28841);
nor U29023 (N_29023,N_28722,N_28967);
or U29024 (N_29024,N_28734,N_28547);
nand U29025 (N_29025,N_28557,N_28668);
or U29026 (N_29026,N_28759,N_28559);
xor U29027 (N_29027,N_28569,N_28585);
and U29028 (N_29028,N_28860,N_28945);
nand U29029 (N_29029,N_28966,N_28981);
and U29030 (N_29030,N_28730,N_28755);
xnor U29031 (N_29031,N_28731,N_28670);
and U29032 (N_29032,N_28911,N_28933);
and U29033 (N_29033,N_28766,N_28746);
and U29034 (N_29034,N_28855,N_28960);
xor U29035 (N_29035,N_28706,N_28656);
xor U29036 (N_29036,N_28948,N_28931);
or U29037 (N_29037,N_28564,N_28815);
or U29038 (N_29038,N_28870,N_28897);
and U29039 (N_29039,N_28613,N_28503);
nand U29040 (N_29040,N_28999,N_28552);
xor U29041 (N_29041,N_28816,N_28509);
xnor U29042 (N_29042,N_28572,N_28753);
nor U29043 (N_29043,N_28717,N_28789);
nand U29044 (N_29044,N_28581,N_28957);
or U29045 (N_29045,N_28672,N_28727);
or U29046 (N_29046,N_28531,N_28906);
nand U29047 (N_29047,N_28535,N_28534);
nor U29048 (N_29048,N_28775,N_28874);
nor U29049 (N_29049,N_28849,N_28788);
nand U29050 (N_29050,N_28776,N_28863);
and U29051 (N_29051,N_28778,N_28714);
or U29052 (N_29052,N_28500,N_28939);
xnor U29053 (N_29053,N_28763,N_28780);
xnor U29054 (N_29054,N_28839,N_28521);
nand U29055 (N_29055,N_28944,N_28963);
and U29056 (N_29056,N_28680,N_28977);
nor U29057 (N_29057,N_28560,N_28996);
nor U29058 (N_29058,N_28513,N_28825);
and U29059 (N_29059,N_28846,N_28857);
nor U29060 (N_29060,N_28867,N_28701);
or U29061 (N_29061,N_28677,N_28881);
and U29062 (N_29062,N_28741,N_28861);
nand U29063 (N_29063,N_28678,N_28919);
and U29064 (N_29064,N_28760,N_28597);
or U29065 (N_29065,N_28884,N_28526);
nor U29066 (N_29066,N_28893,N_28616);
and U29067 (N_29067,N_28512,N_28882);
and U29068 (N_29068,N_28573,N_28566);
xor U29069 (N_29069,N_28538,N_28992);
or U29070 (N_29070,N_28797,N_28617);
nor U29071 (N_29071,N_28924,N_28889);
or U29072 (N_29072,N_28749,N_28579);
or U29073 (N_29073,N_28932,N_28669);
and U29074 (N_29074,N_28748,N_28762);
nor U29075 (N_29075,N_28649,N_28671);
nor U29076 (N_29076,N_28805,N_28876);
or U29077 (N_29077,N_28691,N_28516);
or U29078 (N_29078,N_28699,N_28506);
nand U29079 (N_29079,N_28980,N_28765);
xor U29080 (N_29080,N_28847,N_28655);
and U29081 (N_29081,N_28978,N_28718);
and U29082 (N_29082,N_28705,N_28527);
and U29083 (N_29083,N_28508,N_28761);
and U29084 (N_29084,N_28925,N_28688);
and U29085 (N_29085,N_28729,N_28833);
or U29086 (N_29086,N_28772,N_28519);
nand U29087 (N_29087,N_28594,N_28515);
or U29088 (N_29088,N_28983,N_28986);
and U29089 (N_29089,N_28645,N_28611);
and U29090 (N_29090,N_28837,N_28993);
xnor U29091 (N_29091,N_28796,N_28709);
or U29092 (N_29092,N_28836,N_28886);
and U29093 (N_29093,N_28696,N_28767);
and U29094 (N_29094,N_28615,N_28896);
xnor U29095 (N_29095,N_28888,N_28635);
nor U29096 (N_29096,N_28715,N_28553);
or U29097 (N_29097,N_28739,N_28812);
or U29098 (N_29098,N_28998,N_28523);
and U29099 (N_29099,N_28923,N_28899);
nor U29100 (N_29100,N_28631,N_28593);
xor U29101 (N_29101,N_28824,N_28972);
xnor U29102 (N_29102,N_28629,N_28851);
xnor U29103 (N_29103,N_28938,N_28726);
and U29104 (N_29104,N_28908,N_28758);
nand U29105 (N_29105,N_28864,N_28591);
and U29106 (N_29106,N_28880,N_28885);
nand U29107 (N_29107,N_28757,N_28813);
and U29108 (N_29108,N_28638,N_28912);
or U29109 (N_29109,N_28673,N_28647);
xor U29110 (N_29110,N_28803,N_28943);
and U29111 (N_29111,N_28930,N_28546);
and U29112 (N_29112,N_28785,N_28533);
xor U29113 (N_29113,N_28976,N_28556);
nand U29114 (N_29114,N_28643,N_28894);
xor U29115 (N_29115,N_28536,N_28743);
nand U29116 (N_29116,N_28660,N_28633);
nor U29117 (N_29117,N_28865,N_28604);
nor U29118 (N_29118,N_28792,N_28603);
nand U29119 (N_29119,N_28768,N_28926);
xnor U29120 (N_29120,N_28587,N_28653);
and U29121 (N_29121,N_28558,N_28822);
and U29122 (N_29122,N_28922,N_28806);
or U29123 (N_29123,N_28630,N_28781);
nand U29124 (N_29124,N_28567,N_28644);
and U29125 (N_29125,N_28878,N_28583);
nand U29126 (N_29126,N_28774,N_28783);
nor U29127 (N_29127,N_28862,N_28662);
xnor U29128 (N_29128,N_28586,N_28654);
nand U29129 (N_29129,N_28804,N_28901);
or U29130 (N_29130,N_28646,N_28651);
or U29131 (N_29131,N_28949,N_28777);
nor U29132 (N_29132,N_28707,N_28689);
or U29133 (N_29133,N_28842,N_28802);
or U29134 (N_29134,N_28929,N_28698);
nand U29135 (N_29135,N_28543,N_28735);
and U29136 (N_29136,N_28530,N_28845);
or U29137 (N_29137,N_28711,N_28544);
xnor U29138 (N_29138,N_28900,N_28808);
or U29139 (N_29139,N_28708,N_28562);
nor U29140 (N_29140,N_28625,N_28756);
xnor U29141 (N_29141,N_28661,N_28628);
nor U29142 (N_29142,N_28541,N_28724);
xor U29143 (N_29143,N_28801,N_28575);
nor U29144 (N_29144,N_28610,N_28764);
or U29145 (N_29145,N_28773,N_28770);
and U29146 (N_29146,N_28728,N_28624);
and U29147 (N_29147,N_28873,N_28947);
nor U29148 (N_29148,N_28952,N_28550);
or U29149 (N_29149,N_28955,N_28958);
nand U29150 (N_29150,N_28737,N_28875);
and U29151 (N_29151,N_28525,N_28866);
and U29152 (N_29152,N_28663,N_28692);
and U29153 (N_29153,N_28973,N_28834);
or U29154 (N_29154,N_28713,N_28561);
or U29155 (N_29155,N_28710,N_28674);
or U29156 (N_29156,N_28969,N_28814);
nor U29157 (N_29157,N_28719,N_28975);
and U29158 (N_29158,N_28990,N_28511);
and U29159 (N_29159,N_28612,N_28577);
or U29160 (N_29160,N_28852,N_28989);
or U29161 (N_29161,N_28891,N_28571);
nor U29162 (N_29162,N_28809,N_28823);
nor U29163 (N_29163,N_28830,N_28807);
and U29164 (N_29164,N_28954,N_28532);
nand U29165 (N_29165,N_28574,N_28838);
nand U29166 (N_29166,N_28898,N_28858);
or U29167 (N_29167,N_28994,N_28940);
nand U29168 (N_29168,N_28652,N_28658);
and U29169 (N_29169,N_28520,N_28871);
and U29170 (N_29170,N_28582,N_28974);
nand U29171 (N_29171,N_28921,N_28584);
xnor U29172 (N_29172,N_28695,N_28892);
xnor U29173 (N_29173,N_28716,N_28693);
xnor U29174 (N_29174,N_28872,N_28514);
or U29175 (N_29175,N_28956,N_28987);
xor U29176 (N_29176,N_28848,N_28694);
xor U29177 (N_29177,N_28979,N_28602);
xnor U29178 (N_29178,N_28659,N_28843);
nor U29179 (N_29179,N_28936,N_28608);
nor U29180 (N_29180,N_28917,N_28793);
and U29181 (N_29181,N_28626,N_28614);
nand U29182 (N_29182,N_28964,N_28667);
xnor U29183 (N_29183,N_28596,N_28622);
xnor U29184 (N_29184,N_28568,N_28982);
nand U29185 (N_29185,N_28817,N_28738);
nor U29186 (N_29186,N_28732,N_28524);
or U29187 (N_29187,N_28675,N_28934);
or U29188 (N_29188,N_28600,N_28609);
nor U29189 (N_29189,N_28942,N_28913);
nor U29190 (N_29190,N_28909,N_28539);
nand U29191 (N_29191,N_28697,N_28517);
or U29192 (N_29192,N_28657,N_28914);
and U29193 (N_29193,N_28779,N_28501);
or U29194 (N_29194,N_28800,N_28769);
nand U29195 (N_29195,N_28666,N_28869);
nor U29196 (N_29196,N_28927,N_28682);
and U29197 (N_29197,N_28787,N_28821);
or U29198 (N_29198,N_28690,N_28819);
and U29199 (N_29199,N_28799,N_28832);
or U29200 (N_29200,N_28895,N_28971);
or U29201 (N_29201,N_28782,N_28650);
xor U29202 (N_29202,N_28563,N_28742);
nor U29203 (N_29203,N_28634,N_28522);
xor U29204 (N_29204,N_28723,N_28818);
xnor U29205 (N_29205,N_28950,N_28798);
nor U29206 (N_29206,N_28590,N_28720);
nand U29207 (N_29207,N_28771,N_28620);
nand U29208 (N_29208,N_28605,N_28548);
or U29209 (N_29209,N_28915,N_28984);
nor U29210 (N_29210,N_28570,N_28700);
and U29211 (N_29211,N_28679,N_28676);
or U29212 (N_29212,N_28580,N_28595);
and U29213 (N_29213,N_28937,N_28744);
or U29214 (N_29214,N_28751,N_28820);
xor U29215 (N_29215,N_28951,N_28907);
or U29216 (N_29216,N_28621,N_28997);
nor U29217 (N_29217,N_28618,N_28505);
nand U29218 (N_29218,N_28685,N_28965);
nor U29219 (N_29219,N_28928,N_28890);
and U29220 (N_29220,N_28736,N_28504);
nor U29221 (N_29221,N_28752,N_28540);
or U29222 (N_29222,N_28642,N_28868);
nand U29223 (N_29223,N_28598,N_28665);
nand U29224 (N_29224,N_28795,N_28565);
nor U29225 (N_29225,N_28877,N_28592);
and U29226 (N_29226,N_28640,N_28606);
nand U29227 (N_29227,N_28750,N_28684);
nor U29228 (N_29228,N_28687,N_28786);
and U29229 (N_29229,N_28542,N_28995);
or U29230 (N_29230,N_28970,N_28828);
or U29231 (N_29231,N_28883,N_28537);
nand U29232 (N_29232,N_28856,N_28953);
and U29233 (N_29233,N_28988,N_28733);
xnor U29234 (N_29234,N_28941,N_28681);
nand U29235 (N_29235,N_28648,N_28599);
or U29236 (N_29236,N_28831,N_28827);
nand U29237 (N_29237,N_28904,N_28619);
xnor U29238 (N_29238,N_28607,N_28991);
or U29239 (N_29239,N_28502,N_28902);
nor U29240 (N_29240,N_28968,N_28664);
xor U29241 (N_29241,N_28555,N_28784);
or U29242 (N_29242,N_28962,N_28826);
or U29243 (N_29243,N_28686,N_28810);
or U29244 (N_29244,N_28903,N_28910);
nand U29245 (N_29245,N_28935,N_28835);
nor U29246 (N_29246,N_28529,N_28576);
nand U29247 (N_29247,N_28632,N_28853);
nand U29248 (N_29248,N_28637,N_28578);
nor U29249 (N_29249,N_28905,N_28639);
nor U29250 (N_29250,N_28598,N_28565);
xnor U29251 (N_29251,N_28827,N_28913);
or U29252 (N_29252,N_28572,N_28809);
xor U29253 (N_29253,N_28864,N_28873);
xnor U29254 (N_29254,N_28560,N_28801);
and U29255 (N_29255,N_28708,N_28936);
nor U29256 (N_29256,N_28700,N_28885);
and U29257 (N_29257,N_28504,N_28901);
and U29258 (N_29258,N_28753,N_28954);
and U29259 (N_29259,N_28967,N_28720);
or U29260 (N_29260,N_28733,N_28514);
or U29261 (N_29261,N_28944,N_28997);
nor U29262 (N_29262,N_28771,N_28915);
nor U29263 (N_29263,N_28977,N_28822);
and U29264 (N_29264,N_28730,N_28696);
nand U29265 (N_29265,N_28868,N_28843);
or U29266 (N_29266,N_28968,N_28826);
and U29267 (N_29267,N_28763,N_28535);
or U29268 (N_29268,N_28571,N_28895);
or U29269 (N_29269,N_28812,N_28996);
xnor U29270 (N_29270,N_28917,N_28892);
or U29271 (N_29271,N_28931,N_28713);
nor U29272 (N_29272,N_28742,N_28809);
xnor U29273 (N_29273,N_28948,N_28514);
or U29274 (N_29274,N_28846,N_28974);
xor U29275 (N_29275,N_28865,N_28631);
and U29276 (N_29276,N_28907,N_28679);
or U29277 (N_29277,N_28860,N_28736);
nand U29278 (N_29278,N_28648,N_28987);
and U29279 (N_29279,N_28906,N_28804);
and U29280 (N_29280,N_28769,N_28939);
or U29281 (N_29281,N_28602,N_28762);
nor U29282 (N_29282,N_28535,N_28943);
nand U29283 (N_29283,N_28646,N_28669);
and U29284 (N_29284,N_28770,N_28761);
nand U29285 (N_29285,N_28808,N_28558);
nor U29286 (N_29286,N_28756,N_28798);
nand U29287 (N_29287,N_28742,N_28514);
or U29288 (N_29288,N_28508,N_28987);
nor U29289 (N_29289,N_28940,N_28684);
or U29290 (N_29290,N_28529,N_28526);
and U29291 (N_29291,N_28831,N_28721);
or U29292 (N_29292,N_28617,N_28514);
nor U29293 (N_29293,N_28825,N_28870);
and U29294 (N_29294,N_28560,N_28932);
xor U29295 (N_29295,N_28571,N_28694);
or U29296 (N_29296,N_28527,N_28788);
and U29297 (N_29297,N_28784,N_28950);
xor U29298 (N_29298,N_28709,N_28922);
xor U29299 (N_29299,N_28987,N_28725);
xnor U29300 (N_29300,N_28738,N_28987);
or U29301 (N_29301,N_28738,N_28914);
and U29302 (N_29302,N_28675,N_28759);
or U29303 (N_29303,N_28968,N_28592);
nor U29304 (N_29304,N_28575,N_28730);
xnor U29305 (N_29305,N_28784,N_28916);
nor U29306 (N_29306,N_28616,N_28907);
or U29307 (N_29307,N_28582,N_28898);
nand U29308 (N_29308,N_28737,N_28892);
nor U29309 (N_29309,N_28884,N_28597);
and U29310 (N_29310,N_28593,N_28926);
xor U29311 (N_29311,N_28924,N_28565);
xor U29312 (N_29312,N_28986,N_28504);
nor U29313 (N_29313,N_28891,N_28947);
xnor U29314 (N_29314,N_28729,N_28511);
and U29315 (N_29315,N_28655,N_28916);
nor U29316 (N_29316,N_28571,N_28940);
nand U29317 (N_29317,N_28585,N_28523);
xor U29318 (N_29318,N_28669,N_28790);
or U29319 (N_29319,N_28690,N_28834);
or U29320 (N_29320,N_28692,N_28753);
xor U29321 (N_29321,N_28957,N_28891);
nor U29322 (N_29322,N_28973,N_28784);
nor U29323 (N_29323,N_28694,N_28959);
or U29324 (N_29324,N_28542,N_28715);
and U29325 (N_29325,N_28558,N_28783);
or U29326 (N_29326,N_28955,N_28673);
and U29327 (N_29327,N_28574,N_28585);
nand U29328 (N_29328,N_28817,N_28604);
xnor U29329 (N_29329,N_28603,N_28861);
nor U29330 (N_29330,N_28810,N_28806);
and U29331 (N_29331,N_28797,N_28834);
xnor U29332 (N_29332,N_28899,N_28538);
xnor U29333 (N_29333,N_28803,N_28940);
or U29334 (N_29334,N_28598,N_28827);
and U29335 (N_29335,N_28515,N_28822);
xor U29336 (N_29336,N_28966,N_28557);
xor U29337 (N_29337,N_28990,N_28807);
xnor U29338 (N_29338,N_28760,N_28596);
nor U29339 (N_29339,N_28638,N_28633);
nand U29340 (N_29340,N_28834,N_28560);
or U29341 (N_29341,N_28981,N_28917);
nor U29342 (N_29342,N_28776,N_28689);
and U29343 (N_29343,N_28709,N_28975);
nor U29344 (N_29344,N_28732,N_28905);
nand U29345 (N_29345,N_28615,N_28680);
nor U29346 (N_29346,N_28936,N_28937);
or U29347 (N_29347,N_28936,N_28531);
xnor U29348 (N_29348,N_28687,N_28599);
xnor U29349 (N_29349,N_28645,N_28630);
nand U29350 (N_29350,N_28895,N_28573);
or U29351 (N_29351,N_28586,N_28913);
nor U29352 (N_29352,N_28715,N_28779);
nand U29353 (N_29353,N_28833,N_28865);
xor U29354 (N_29354,N_28885,N_28951);
xor U29355 (N_29355,N_28783,N_28747);
xor U29356 (N_29356,N_28892,N_28734);
nand U29357 (N_29357,N_28736,N_28990);
nor U29358 (N_29358,N_28772,N_28534);
and U29359 (N_29359,N_28993,N_28596);
or U29360 (N_29360,N_28859,N_28833);
nand U29361 (N_29361,N_28943,N_28538);
or U29362 (N_29362,N_28555,N_28989);
nor U29363 (N_29363,N_28817,N_28812);
or U29364 (N_29364,N_28589,N_28524);
or U29365 (N_29365,N_28982,N_28826);
and U29366 (N_29366,N_28759,N_28789);
and U29367 (N_29367,N_28661,N_28768);
or U29368 (N_29368,N_28694,N_28676);
nor U29369 (N_29369,N_28924,N_28632);
nor U29370 (N_29370,N_28785,N_28903);
nand U29371 (N_29371,N_28725,N_28804);
or U29372 (N_29372,N_28535,N_28997);
or U29373 (N_29373,N_28521,N_28941);
nand U29374 (N_29374,N_28962,N_28799);
xnor U29375 (N_29375,N_28677,N_28782);
xor U29376 (N_29376,N_28514,N_28905);
nand U29377 (N_29377,N_28574,N_28658);
nor U29378 (N_29378,N_28615,N_28658);
nand U29379 (N_29379,N_28912,N_28541);
or U29380 (N_29380,N_28789,N_28839);
nand U29381 (N_29381,N_28661,N_28524);
or U29382 (N_29382,N_28834,N_28552);
and U29383 (N_29383,N_28804,N_28957);
or U29384 (N_29384,N_28557,N_28864);
xnor U29385 (N_29385,N_28703,N_28627);
xor U29386 (N_29386,N_28735,N_28821);
nand U29387 (N_29387,N_28777,N_28899);
and U29388 (N_29388,N_28999,N_28882);
and U29389 (N_29389,N_28815,N_28728);
and U29390 (N_29390,N_28686,N_28730);
nor U29391 (N_29391,N_28762,N_28712);
nor U29392 (N_29392,N_28503,N_28502);
or U29393 (N_29393,N_28896,N_28756);
and U29394 (N_29394,N_28501,N_28642);
or U29395 (N_29395,N_28897,N_28996);
and U29396 (N_29396,N_28806,N_28824);
nor U29397 (N_29397,N_28956,N_28843);
and U29398 (N_29398,N_28521,N_28905);
xor U29399 (N_29399,N_28717,N_28909);
and U29400 (N_29400,N_28777,N_28906);
or U29401 (N_29401,N_28682,N_28591);
nor U29402 (N_29402,N_28551,N_28884);
or U29403 (N_29403,N_28578,N_28702);
nand U29404 (N_29404,N_28508,N_28653);
and U29405 (N_29405,N_28608,N_28838);
and U29406 (N_29406,N_28663,N_28970);
or U29407 (N_29407,N_28900,N_28892);
nand U29408 (N_29408,N_28799,N_28975);
nor U29409 (N_29409,N_28635,N_28652);
nand U29410 (N_29410,N_28907,N_28868);
xor U29411 (N_29411,N_28625,N_28521);
nor U29412 (N_29412,N_28653,N_28635);
or U29413 (N_29413,N_28738,N_28964);
or U29414 (N_29414,N_28523,N_28872);
xor U29415 (N_29415,N_28697,N_28776);
xnor U29416 (N_29416,N_28503,N_28507);
nand U29417 (N_29417,N_28971,N_28945);
and U29418 (N_29418,N_28662,N_28634);
nor U29419 (N_29419,N_28953,N_28590);
or U29420 (N_29420,N_28870,N_28508);
and U29421 (N_29421,N_28680,N_28743);
and U29422 (N_29422,N_28879,N_28933);
and U29423 (N_29423,N_28941,N_28792);
xor U29424 (N_29424,N_28826,N_28764);
and U29425 (N_29425,N_28673,N_28638);
nand U29426 (N_29426,N_28646,N_28535);
nand U29427 (N_29427,N_28523,N_28569);
or U29428 (N_29428,N_28954,N_28647);
nand U29429 (N_29429,N_28916,N_28633);
or U29430 (N_29430,N_28595,N_28555);
xnor U29431 (N_29431,N_28539,N_28935);
xnor U29432 (N_29432,N_28649,N_28742);
nand U29433 (N_29433,N_28725,N_28670);
or U29434 (N_29434,N_28735,N_28759);
nand U29435 (N_29435,N_28593,N_28923);
xnor U29436 (N_29436,N_28588,N_28659);
nand U29437 (N_29437,N_28675,N_28892);
nand U29438 (N_29438,N_28831,N_28650);
or U29439 (N_29439,N_28988,N_28868);
nand U29440 (N_29440,N_28827,N_28560);
nand U29441 (N_29441,N_28955,N_28903);
nand U29442 (N_29442,N_28639,N_28682);
nand U29443 (N_29443,N_28904,N_28865);
nor U29444 (N_29444,N_28828,N_28577);
nand U29445 (N_29445,N_28752,N_28988);
nand U29446 (N_29446,N_28992,N_28986);
nand U29447 (N_29447,N_28802,N_28952);
and U29448 (N_29448,N_28824,N_28654);
nor U29449 (N_29449,N_28675,N_28804);
or U29450 (N_29450,N_28972,N_28876);
and U29451 (N_29451,N_28612,N_28676);
and U29452 (N_29452,N_28872,N_28691);
nor U29453 (N_29453,N_28750,N_28957);
nor U29454 (N_29454,N_28671,N_28923);
nand U29455 (N_29455,N_28970,N_28784);
or U29456 (N_29456,N_28926,N_28911);
or U29457 (N_29457,N_28947,N_28704);
nor U29458 (N_29458,N_28983,N_28858);
or U29459 (N_29459,N_28857,N_28507);
nand U29460 (N_29460,N_28986,N_28813);
xnor U29461 (N_29461,N_28595,N_28985);
nand U29462 (N_29462,N_28706,N_28722);
and U29463 (N_29463,N_28726,N_28740);
xor U29464 (N_29464,N_28747,N_28977);
xor U29465 (N_29465,N_28994,N_28951);
nor U29466 (N_29466,N_28976,N_28989);
and U29467 (N_29467,N_28595,N_28510);
xor U29468 (N_29468,N_28942,N_28507);
and U29469 (N_29469,N_28705,N_28532);
nand U29470 (N_29470,N_28777,N_28647);
and U29471 (N_29471,N_28774,N_28801);
nand U29472 (N_29472,N_28866,N_28804);
or U29473 (N_29473,N_28789,N_28567);
xor U29474 (N_29474,N_28757,N_28863);
nor U29475 (N_29475,N_28818,N_28560);
xnor U29476 (N_29476,N_28745,N_28652);
nor U29477 (N_29477,N_28967,N_28705);
or U29478 (N_29478,N_28615,N_28829);
nor U29479 (N_29479,N_28779,N_28911);
xnor U29480 (N_29480,N_28791,N_28577);
nor U29481 (N_29481,N_28795,N_28846);
xor U29482 (N_29482,N_28899,N_28836);
nor U29483 (N_29483,N_28590,N_28987);
nand U29484 (N_29484,N_28967,N_28862);
and U29485 (N_29485,N_28834,N_28566);
xnor U29486 (N_29486,N_28527,N_28683);
and U29487 (N_29487,N_28533,N_28607);
or U29488 (N_29488,N_28650,N_28612);
or U29489 (N_29489,N_28598,N_28527);
nand U29490 (N_29490,N_28519,N_28567);
nand U29491 (N_29491,N_28966,N_28827);
nor U29492 (N_29492,N_28746,N_28564);
and U29493 (N_29493,N_28747,N_28996);
nor U29494 (N_29494,N_28728,N_28756);
or U29495 (N_29495,N_28827,N_28821);
and U29496 (N_29496,N_28683,N_28786);
or U29497 (N_29497,N_28900,N_28982);
xor U29498 (N_29498,N_28694,N_28649);
or U29499 (N_29499,N_28726,N_28587);
nor U29500 (N_29500,N_29045,N_29188);
or U29501 (N_29501,N_29404,N_29490);
nor U29502 (N_29502,N_29467,N_29100);
nand U29503 (N_29503,N_29290,N_29259);
nor U29504 (N_29504,N_29406,N_29476);
nand U29505 (N_29505,N_29136,N_29277);
nor U29506 (N_29506,N_29401,N_29203);
nand U29507 (N_29507,N_29382,N_29035);
and U29508 (N_29508,N_29305,N_29037);
or U29509 (N_29509,N_29351,N_29071);
and U29510 (N_29510,N_29472,N_29286);
nand U29511 (N_29511,N_29260,N_29226);
nand U29512 (N_29512,N_29345,N_29448);
nand U29513 (N_29513,N_29067,N_29279);
xor U29514 (N_29514,N_29094,N_29042);
or U29515 (N_29515,N_29184,N_29295);
nand U29516 (N_29516,N_29074,N_29271);
nand U29517 (N_29517,N_29106,N_29254);
or U29518 (N_29518,N_29311,N_29170);
or U29519 (N_29519,N_29114,N_29312);
nor U29520 (N_29520,N_29486,N_29264);
nor U29521 (N_29521,N_29245,N_29430);
and U29522 (N_29522,N_29176,N_29428);
and U29523 (N_29523,N_29481,N_29052);
nor U29524 (N_29524,N_29319,N_29174);
xnor U29525 (N_29525,N_29473,N_29381);
xor U29526 (N_29526,N_29018,N_29200);
xnor U29527 (N_29527,N_29364,N_29123);
or U29528 (N_29528,N_29454,N_29463);
nor U29529 (N_29529,N_29040,N_29474);
xor U29530 (N_29530,N_29014,N_29142);
and U29531 (N_29531,N_29355,N_29113);
or U29532 (N_29532,N_29433,N_29363);
nor U29533 (N_29533,N_29118,N_29144);
nor U29534 (N_29534,N_29165,N_29220);
nor U29535 (N_29535,N_29301,N_29039);
or U29536 (N_29536,N_29055,N_29267);
nor U29537 (N_29537,N_29047,N_29438);
nor U29538 (N_29538,N_29346,N_29069);
xor U29539 (N_29539,N_29198,N_29225);
nand U29540 (N_29540,N_29053,N_29031);
nand U29541 (N_29541,N_29131,N_29120);
or U29542 (N_29542,N_29297,N_29041);
or U29543 (N_29543,N_29491,N_29426);
and U29544 (N_29544,N_29325,N_29195);
and U29545 (N_29545,N_29166,N_29077);
and U29546 (N_29546,N_29076,N_29348);
or U29547 (N_29547,N_29101,N_29026);
or U29548 (N_29548,N_29344,N_29365);
and U29549 (N_29549,N_29459,N_29098);
nand U29550 (N_29550,N_29202,N_29065);
nor U29551 (N_29551,N_29180,N_29419);
xnor U29552 (N_29552,N_29300,N_29462);
nor U29553 (N_29553,N_29493,N_29289);
or U29554 (N_29554,N_29083,N_29232);
xor U29555 (N_29555,N_29058,N_29450);
xnor U29556 (N_29556,N_29262,N_29334);
xor U29557 (N_29557,N_29273,N_29028);
xor U29558 (N_29558,N_29337,N_29299);
or U29559 (N_29559,N_29284,N_29499);
and U29560 (N_29560,N_29379,N_29274);
nor U29561 (N_29561,N_29377,N_29024);
or U29562 (N_29562,N_29358,N_29051);
xor U29563 (N_29563,N_29475,N_29070);
xnor U29564 (N_29564,N_29244,N_29078);
nor U29565 (N_29565,N_29164,N_29169);
or U29566 (N_29566,N_29292,N_29460);
xnor U29567 (N_29567,N_29457,N_29089);
xor U29568 (N_29568,N_29294,N_29362);
and U29569 (N_29569,N_29064,N_29395);
nand U29570 (N_29570,N_29167,N_29233);
nand U29571 (N_29571,N_29372,N_29272);
xnor U29572 (N_29572,N_29258,N_29335);
and U29573 (N_29573,N_29062,N_29234);
or U29574 (N_29574,N_29445,N_29405);
and U29575 (N_29575,N_29376,N_29352);
nor U29576 (N_29576,N_29353,N_29321);
nor U29577 (N_29577,N_29266,N_29011);
nand U29578 (N_29578,N_29086,N_29153);
or U29579 (N_29579,N_29084,N_29402);
xnor U29580 (N_29580,N_29310,N_29020);
xnor U29581 (N_29581,N_29398,N_29073);
xnor U29582 (N_29582,N_29343,N_29477);
or U29583 (N_29583,N_29196,N_29326);
or U29584 (N_29584,N_29239,N_29126);
and U29585 (N_29585,N_29434,N_29494);
nand U29586 (N_29586,N_29096,N_29141);
xor U29587 (N_29587,N_29480,N_29392);
and U29588 (N_29588,N_29022,N_29417);
xnor U29589 (N_29589,N_29054,N_29361);
and U29590 (N_29590,N_29149,N_29440);
nand U29591 (N_29591,N_29161,N_29383);
or U29592 (N_29592,N_29420,N_29479);
nor U29593 (N_29593,N_29158,N_29338);
nand U29594 (N_29594,N_29498,N_29139);
nor U29595 (N_29595,N_29129,N_29190);
or U29596 (N_29596,N_29241,N_29132);
xor U29597 (N_29597,N_29119,N_29194);
nor U29598 (N_29598,N_29308,N_29108);
and U29599 (N_29599,N_29110,N_29323);
xor U29600 (N_29600,N_29210,N_29302);
nand U29601 (N_29601,N_29303,N_29025);
xor U29602 (N_29602,N_29093,N_29044);
nor U29603 (N_29603,N_29324,N_29207);
nor U29604 (N_29604,N_29464,N_29341);
xor U29605 (N_29605,N_29327,N_29103);
xor U29606 (N_29606,N_29489,N_29214);
nand U29607 (N_29607,N_29437,N_29060);
or U29608 (N_29608,N_29012,N_29121);
and U29609 (N_29609,N_29436,N_29191);
nand U29610 (N_29610,N_29015,N_29206);
or U29611 (N_29611,N_29322,N_29487);
or U29612 (N_29612,N_29332,N_29399);
xnor U29613 (N_29613,N_29005,N_29143);
nand U29614 (N_29614,N_29160,N_29138);
xnor U29615 (N_29615,N_29342,N_29116);
and U29616 (N_29616,N_29411,N_29228);
xnor U29617 (N_29617,N_29270,N_29168);
xor U29618 (N_29618,N_29293,N_29000);
xnor U29619 (N_29619,N_29019,N_29181);
and U29620 (N_29620,N_29368,N_29304);
nor U29621 (N_29621,N_29049,N_29235);
xnor U29622 (N_29622,N_29378,N_29127);
nor U29623 (N_29623,N_29407,N_29213);
and U29624 (N_29624,N_29124,N_29246);
or U29625 (N_29625,N_29389,N_29291);
and U29626 (N_29626,N_29257,N_29097);
nor U29627 (N_29627,N_29238,N_29066);
nor U29628 (N_29628,N_29380,N_29313);
nor U29629 (N_29629,N_29135,N_29057);
nor U29630 (N_29630,N_29115,N_29090);
xnor U29631 (N_29631,N_29468,N_29151);
nor U29632 (N_29632,N_29409,N_29027);
nand U29633 (N_29633,N_29029,N_29186);
or U29634 (N_29634,N_29488,N_29004);
nand U29635 (N_29635,N_29092,N_29256);
xnor U29636 (N_29636,N_29485,N_29229);
nor U29637 (N_29637,N_29133,N_29340);
or U29638 (N_29638,N_29208,N_29243);
or U29639 (N_29639,N_29209,N_29163);
xor U29640 (N_29640,N_29424,N_29449);
xor U29641 (N_29641,N_29223,N_29001);
or U29642 (N_29642,N_29105,N_29285);
and U29643 (N_29643,N_29193,N_29393);
nor U29644 (N_29644,N_29287,N_29387);
xnor U29645 (N_29645,N_29384,N_29217);
or U29646 (N_29646,N_29453,N_29043);
nand U29647 (N_29647,N_29492,N_29231);
nor U29648 (N_29648,N_29038,N_29173);
and U29649 (N_29649,N_29212,N_29400);
nor U29650 (N_29650,N_29439,N_29320);
nand U29651 (N_29651,N_29375,N_29386);
or U29652 (N_29652,N_29183,N_29242);
and U29653 (N_29653,N_29427,N_29403);
nand U29654 (N_29654,N_29162,N_29224);
and U29655 (N_29655,N_29339,N_29109);
and U29656 (N_29656,N_29391,N_29081);
or U29657 (N_29657,N_29354,N_29315);
nand U29658 (N_29658,N_29429,N_29046);
or U29659 (N_29659,N_29478,N_29061);
xnor U29660 (N_29660,N_29248,N_29349);
and U29661 (N_29661,N_29178,N_29413);
or U29662 (N_29662,N_29140,N_29150);
nor U29663 (N_29663,N_29314,N_29425);
and U29664 (N_29664,N_29441,N_29280);
nand U29665 (N_29665,N_29189,N_29227);
nor U29666 (N_29666,N_29360,N_29152);
or U29667 (N_29667,N_29282,N_29099);
xnor U29668 (N_29668,N_29374,N_29444);
nand U29669 (N_29669,N_29385,N_29397);
nor U29670 (N_29670,N_29048,N_29009);
or U29671 (N_29671,N_29456,N_29471);
nor U29672 (N_29672,N_29204,N_29175);
xnor U29673 (N_29673,N_29495,N_29415);
xor U29674 (N_29674,N_29388,N_29033);
nor U29675 (N_29675,N_29366,N_29298);
and U29676 (N_29676,N_29091,N_29145);
xor U29677 (N_29677,N_29222,N_29316);
xor U29678 (N_29678,N_29010,N_29112);
nor U29679 (N_29679,N_29177,N_29357);
and U29680 (N_29680,N_29269,N_29156);
nand U29681 (N_29681,N_29102,N_29185);
xnor U29682 (N_29682,N_29215,N_29159);
and U29683 (N_29683,N_29182,N_29367);
xnor U29684 (N_29684,N_29331,N_29416);
and U29685 (N_29685,N_29219,N_29036);
nand U29686 (N_29686,N_29137,N_29087);
nor U29687 (N_29687,N_29251,N_29455);
or U29688 (N_29688,N_29032,N_29470);
and U29689 (N_29689,N_29216,N_29482);
or U29690 (N_29690,N_29157,N_29171);
nor U29691 (N_29691,N_29082,N_29201);
and U29692 (N_29692,N_29068,N_29147);
xor U29693 (N_29693,N_29281,N_29007);
or U29694 (N_29694,N_29394,N_29063);
xnor U29695 (N_29695,N_29418,N_29469);
nand U29696 (N_29696,N_29423,N_29451);
and U29697 (N_29697,N_29017,N_29432);
or U29698 (N_29698,N_29261,N_29431);
and U29699 (N_29699,N_29333,N_29421);
and U29700 (N_29700,N_29023,N_29104);
or U29701 (N_29701,N_29288,N_29329);
xor U29702 (N_29702,N_29088,N_29249);
nand U29703 (N_29703,N_29317,N_29197);
xnor U29704 (N_29704,N_29075,N_29111);
nand U29705 (N_29705,N_29034,N_29107);
and U29706 (N_29706,N_29496,N_29148);
xor U29707 (N_29707,N_29013,N_29199);
nand U29708 (N_29708,N_29452,N_29296);
xnor U29709 (N_29709,N_29336,N_29172);
nor U29710 (N_29710,N_29056,N_29356);
and U29711 (N_29711,N_29347,N_29465);
or U29712 (N_29712,N_29179,N_29359);
and U29713 (N_29713,N_29371,N_29390);
nor U29714 (N_29714,N_29373,N_29059);
xor U29715 (N_29715,N_29252,N_29205);
nand U29716 (N_29716,N_29085,N_29484);
nand U29717 (N_29717,N_29412,N_29122);
or U29718 (N_29718,N_29117,N_29370);
and U29719 (N_29719,N_29250,N_29350);
nand U29720 (N_29720,N_29237,N_29247);
nand U29721 (N_29721,N_29461,N_29442);
or U29722 (N_29722,N_29283,N_29211);
nor U29723 (N_29723,N_29240,N_29307);
and U29724 (N_29724,N_29080,N_29276);
nand U29725 (N_29725,N_29072,N_29435);
xnor U29726 (N_29726,N_29408,N_29497);
and U29727 (N_29727,N_29446,N_29002);
xnor U29728 (N_29728,N_29230,N_29134);
nor U29729 (N_29729,N_29447,N_29253);
nand U29730 (N_29730,N_29218,N_29410);
nand U29731 (N_29731,N_29146,N_29130);
or U29732 (N_29732,N_29330,N_29050);
xnor U29733 (N_29733,N_29306,N_29221);
and U29734 (N_29734,N_29396,N_29030);
and U29735 (N_29735,N_29255,N_29155);
or U29736 (N_29736,N_29275,N_29263);
xor U29737 (N_29737,N_29422,N_29008);
nor U29738 (N_29738,N_29466,N_29318);
or U29739 (N_29739,N_29125,N_29187);
xor U29740 (N_29740,N_29016,N_29192);
nor U29741 (N_29741,N_29483,N_29021);
nand U29742 (N_29742,N_29128,N_29095);
xor U29743 (N_29743,N_29369,N_29154);
nor U29744 (N_29744,N_29278,N_29265);
nand U29745 (N_29745,N_29328,N_29268);
nand U29746 (N_29746,N_29414,N_29443);
nand U29747 (N_29747,N_29309,N_29236);
or U29748 (N_29748,N_29003,N_29006);
xor U29749 (N_29749,N_29079,N_29458);
and U29750 (N_29750,N_29169,N_29493);
or U29751 (N_29751,N_29477,N_29476);
xnor U29752 (N_29752,N_29205,N_29188);
nor U29753 (N_29753,N_29053,N_29440);
xnor U29754 (N_29754,N_29128,N_29105);
nand U29755 (N_29755,N_29009,N_29234);
or U29756 (N_29756,N_29073,N_29177);
xnor U29757 (N_29757,N_29119,N_29279);
and U29758 (N_29758,N_29483,N_29068);
nand U29759 (N_29759,N_29415,N_29268);
or U29760 (N_29760,N_29099,N_29268);
and U29761 (N_29761,N_29388,N_29165);
xnor U29762 (N_29762,N_29330,N_29403);
and U29763 (N_29763,N_29191,N_29074);
nand U29764 (N_29764,N_29122,N_29254);
or U29765 (N_29765,N_29326,N_29156);
and U29766 (N_29766,N_29096,N_29458);
or U29767 (N_29767,N_29350,N_29331);
or U29768 (N_29768,N_29380,N_29376);
nor U29769 (N_29769,N_29087,N_29428);
and U29770 (N_29770,N_29491,N_29425);
or U29771 (N_29771,N_29270,N_29054);
nand U29772 (N_29772,N_29166,N_29229);
nand U29773 (N_29773,N_29306,N_29132);
nand U29774 (N_29774,N_29095,N_29201);
xor U29775 (N_29775,N_29134,N_29008);
xor U29776 (N_29776,N_29040,N_29081);
or U29777 (N_29777,N_29023,N_29231);
and U29778 (N_29778,N_29139,N_29440);
nor U29779 (N_29779,N_29287,N_29239);
nand U29780 (N_29780,N_29352,N_29033);
and U29781 (N_29781,N_29027,N_29184);
and U29782 (N_29782,N_29155,N_29217);
nand U29783 (N_29783,N_29133,N_29406);
nor U29784 (N_29784,N_29038,N_29054);
nor U29785 (N_29785,N_29413,N_29053);
and U29786 (N_29786,N_29133,N_29375);
or U29787 (N_29787,N_29032,N_29221);
or U29788 (N_29788,N_29076,N_29084);
xnor U29789 (N_29789,N_29359,N_29007);
or U29790 (N_29790,N_29328,N_29471);
or U29791 (N_29791,N_29015,N_29047);
nor U29792 (N_29792,N_29393,N_29048);
and U29793 (N_29793,N_29051,N_29211);
xnor U29794 (N_29794,N_29236,N_29266);
or U29795 (N_29795,N_29312,N_29241);
or U29796 (N_29796,N_29338,N_29172);
xnor U29797 (N_29797,N_29149,N_29271);
and U29798 (N_29798,N_29086,N_29163);
or U29799 (N_29799,N_29186,N_29185);
or U29800 (N_29800,N_29009,N_29171);
nor U29801 (N_29801,N_29019,N_29434);
nor U29802 (N_29802,N_29052,N_29199);
nor U29803 (N_29803,N_29305,N_29023);
or U29804 (N_29804,N_29378,N_29062);
or U29805 (N_29805,N_29007,N_29318);
nand U29806 (N_29806,N_29433,N_29349);
xor U29807 (N_29807,N_29481,N_29163);
nor U29808 (N_29808,N_29484,N_29084);
or U29809 (N_29809,N_29057,N_29344);
and U29810 (N_29810,N_29191,N_29343);
nand U29811 (N_29811,N_29149,N_29338);
or U29812 (N_29812,N_29447,N_29071);
xnor U29813 (N_29813,N_29313,N_29456);
nor U29814 (N_29814,N_29474,N_29084);
xor U29815 (N_29815,N_29061,N_29324);
and U29816 (N_29816,N_29064,N_29397);
and U29817 (N_29817,N_29020,N_29302);
xor U29818 (N_29818,N_29420,N_29104);
nand U29819 (N_29819,N_29024,N_29497);
or U29820 (N_29820,N_29289,N_29096);
xnor U29821 (N_29821,N_29350,N_29383);
nor U29822 (N_29822,N_29419,N_29323);
nand U29823 (N_29823,N_29099,N_29283);
xnor U29824 (N_29824,N_29390,N_29323);
nor U29825 (N_29825,N_29351,N_29014);
xor U29826 (N_29826,N_29296,N_29078);
nor U29827 (N_29827,N_29442,N_29098);
and U29828 (N_29828,N_29145,N_29497);
nand U29829 (N_29829,N_29014,N_29388);
nand U29830 (N_29830,N_29010,N_29156);
and U29831 (N_29831,N_29378,N_29398);
and U29832 (N_29832,N_29094,N_29481);
and U29833 (N_29833,N_29235,N_29289);
or U29834 (N_29834,N_29454,N_29222);
nand U29835 (N_29835,N_29045,N_29152);
nor U29836 (N_29836,N_29316,N_29330);
nand U29837 (N_29837,N_29096,N_29238);
and U29838 (N_29838,N_29378,N_29459);
nand U29839 (N_29839,N_29381,N_29291);
xnor U29840 (N_29840,N_29061,N_29309);
nor U29841 (N_29841,N_29347,N_29080);
or U29842 (N_29842,N_29007,N_29206);
and U29843 (N_29843,N_29162,N_29491);
or U29844 (N_29844,N_29450,N_29053);
nor U29845 (N_29845,N_29041,N_29261);
nor U29846 (N_29846,N_29020,N_29300);
xnor U29847 (N_29847,N_29082,N_29319);
or U29848 (N_29848,N_29352,N_29408);
xnor U29849 (N_29849,N_29158,N_29295);
nor U29850 (N_29850,N_29499,N_29291);
nor U29851 (N_29851,N_29359,N_29483);
nor U29852 (N_29852,N_29086,N_29387);
and U29853 (N_29853,N_29274,N_29195);
nand U29854 (N_29854,N_29242,N_29422);
nor U29855 (N_29855,N_29071,N_29481);
nand U29856 (N_29856,N_29307,N_29416);
and U29857 (N_29857,N_29026,N_29453);
xor U29858 (N_29858,N_29166,N_29218);
nand U29859 (N_29859,N_29014,N_29373);
nor U29860 (N_29860,N_29284,N_29048);
nor U29861 (N_29861,N_29051,N_29483);
nand U29862 (N_29862,N_29159,N_29258);
and U29863 (N_29863,N_29260,N_29073);
xor U29864 (N_29864,N_29195,N_29387);
nor U29865 (N_29865,N_29085,N_29297);
nor U29866 (N_29866,N_29344,N_29287);
nand U29867 (N_29867,N_29251,N_29038);
xnor U29868 (N_29868,N_29035,N_29038);
or U29869 (N_29869,N_29450,N_29247);
nor U29870 (N_29870,N_29072,N_29156);
and U29871 (N_29871,N_29018,N_29368);
or U29872 (N_29872,N_29339,N_29056);
and U29873 (N_29873,N_29058,N_29018);
nor U29874 (N_29874,N_29228,N_29034);
nand U29875 (N_29875,N_29317,N_29378);
nand U29876 (N_29876,N_29447,N_29426);
nand U29877 (N_29877,N_29170,N_29268);
nand U29878 (N_29878,N_29480,N_29236);
and U29879 (N_29879,N_29234,N_29008);
and U29880 (N_29880,N_29450,N_29212);
nand U29881 (N_29881,N_29313,N_29133);
xnor U29882 (N_29882,N_29268,N_29116);
or U29883 (N_29883,N_29254,N_29449);
xnor U29884 (N_29884,N_29098,N_29316);
or U29885 (N_29885,N_29213,N_29185);
nor U29886 (N_29886,N_29049,N_29330);
nor U29887 (N_29887,N_29137,N_29016);
nor U29888 (N_29888,N_29176,N_29244);
nand U29889 (N_29889,N_29176,N_29154);
and U29890 (N_29890,N_29197,N_29111);
nand U29891 (N_29891,N_29340,N_29348);
nor U29892 (N_29892,N_29395,N_29436);
or U29893 (N_29893,N_29094,N_29195);
or U29894 (N_29894,N_29128,N_29319);
nor U29895 (N_29895,N_29440,N_29207);
and U29896 (N_29896,N_29031,N_29373);
or U29897 (N_29897,N_29187,N_29257);
and U29898 (N_29898,N_29077,N_29300);
nor U29899 (N_29899,N_29443,N_29209);
nor U29900 (N_29900,N_29132,N_29364);
nor U29901 (N_29901,N_29079,N_29118);
nor U29902 (N_29902,N_29089,N_29394);
nand U29903 (N_29903,N_29205,N_29174);
xnor U29904 (N_29904,N_29469,N_29133);
or U29905 (N_29905,N_29152,N_29448);
nand U29906 (N_29906,N_29022,N_29049);
and U29907 (N_29907,N_29134,N_29085);
nor U29908 (N_29908,N_29296,N_29170);
or U29909 (N_29909,N_29412,N_29047);
nand U29910 (N_29910,N_29072,N_29307);
and U29911 (N_29911,N_29457,N_29098);
xor U29912 (N_29912,N_29472,N_29419);
nor U29913 (N_29913,N_29408,N_29023);
or U29914 (N_29914,N_29496,N_29481);
and U29915 (N_29915,N_29457,N_29375);
nor U29916 (N_29916,N_29018,N_29103);
and U29917 (N_29917,N_29064,N_29099);
and U29918 (N_29918,N_29064,N_29151);
and U29919 (N_29919,N_29424,N_29151);
nor U29920 (N_29920,N_29027,N_29262);
or U29921 (N_29921,N_29273,N_29357);
nand U29922 (N_29922,N_29083,N_29058);
nand U29923 (N_29923,N_29037,N_29107);
and U29924 (N_29924,N_29267,N_29391);
xor U29925 (N_29925,N_29163,N_29287);
or U29926 (N_29926,N_29182,N_29402);
nor U29927 (N_29927,N_29108,N_29276);
xor U29928 (N_29928,N_29355,N_29024);
nor U29929 (N_29929,N_29306,N_29493);
or U29930 (N_29930,N_29300,N_29152);
nor U29931 (N_29931,N_29359,N_29047);
nand U29932 (N_29932,N_29077,N_29087);
xor U29933 (N_29933,N_29155,N_29326);
xor U29934 (N_29934,N_29457,N_29231);
nor U29935 (N_29935,N_29440,N_29275);
xnor U29936 (N_29936,N_29057,N_29224);
nor U29937 (N_29937,N_29080,N_29238);
or U29938 (N_29938,N_29013,N_29377);
or U29939 (N_29939,N_29148,N_29047);
nand U29940 (N_29940,N_29229,N_29168);
nand U29941 (N_29941,N_29257,N_29076);
or U29942 (N_29942,N_29474,N_29203);
and U29943 (N_29943,N_29069,N_29049);
nand U29944 (N_29944,N_29438,N_29024);
nor U29945 (N_29945,N_29276,N_29177);
nor U29946 (N_29946,N_29456,N_29079);
nor U29947 (N_29947,N_29212,N_29062);
xor U29948 (N_29948,N_29198,N_29143);
nor U29949 (N_29949,N_29065,N_29066);
or U29950 (N_29950,N_29480,N_29267);
nand U29951 (N_29951,N_29045,N_29064);
and U29952 (N_29952,N_29429,N_29217);
nand U29953 (N_29953,N_29043,N_29402);
nor U29954 (N_29954,N_29219,N_29040);
and U29955 (N_29955,N_29143,N_29241);
or U29956 (N_29956,N_29021,N_29226);
or U29957 (N_29957,N_29199,N_29404);
and U29958 (N_29958,N_29484,N_29193);
or U29959 (N_29959,N_29282,N_29362);
nand U29960 (N_29960,N_29191,N_29082);
nor U29961 (N_29961,N_29047,N_29184);
xor U29962 (N_29962,N_29153,N_29095);
or U29963 (N_29963,N_29366,N_29444);
nand U29964 (N_29964,N_29466,N_29002);
or U29965 (N_29965,N_29284,N_29229);
xnor U29966 (N_29966,N_29172,N_29044);
and U29967 (N_29967,N_29092,N_29082);
nor U29968 (N_29968,N_29399,N_29463);
xnor U29969 (N_29969,N_29062,N_29166);
and U29970 (N_29970,N_29051,N_29325);
xnor U29971 (N_29971,N_29013,N_29479);
xor U29972 (N_29972,N_29225,N_29090);
nand U29973 (N_29973,N_29186,N_29427);
xor U29974 (N_29974,N_29418,N_29305);
nor U29975 (N_29975,N_29070,N_29128);
nand U29976 (N_29976,N_29233,N_29324);
xor U29977 (N_29977,N_29188,N_29094);
nor U29978 (N_29978,N_29460,N_29003);
or U29979 (N_29979,N_29173,N_29223);
and U29980 (N_29980,N_29301,N_29266);
and U29981 (N_29981,N_29036,N_29162);
and U29982 (N_29982,N_29103,N_29371);
and U29983 (N_29983,N_29072,N_29083);
xor U29984 (N_29984,N_29291,N_29153);
nor U29985 (N_29985,N_29315,N_29475);
nand U29986 (N_29986,N_29321,N_29267);
nor U29987 (N_29987,N_29028,N_29201);
or U29988 (N_29988,N_29017,N_29170);
and U29989 (N_29989,N_29190,N_29320);
nor U29990 (N_29990,N_29198,N_29322);
or U29991 (N_29991,N_29323,N_29172);
and U29992 (N_29992,N_29258,N_29239);
and U29993 (N_29993,N_29137,N_29388);
or U29994 (N_29994,N_29306,N_29374);
nand U29995 (N_29995,N_29082,N_29424);
and U29996 (N_29996,N_29028,N_29332);
nand U29997 (N_29997,N_29275,N_29322);
nand U29998 (N_29998,N_29261,N_29254);
and U29999 (N_29999,N_29488,N_29324);
or UO_0 (O_0,N_29518,N_29925);
nand UO_1 (O_1,N_29665,N_29607);
xnor UO_2 (O_2,N_29877,N_29967);
nand UO_3 (O_3,N_29619,N_29782);
and UO_4 (O_4,N_29680,N_29610);
or UO_5 (O_5,N_29966,N_29831);
or UO_6 (O_6,N_29906,N_29540);
nor UO_7 (O_7,N_29555,N_29760);
nor UO_8 (O_8,N_29813,N_29505);
nand UO_9 (O_9,N_29626,N_29734);
nand UO_10 (O_10,N_29705,N_29554);
or UO_11 (O_11,N_29566,N_29524);
xnor UO_12 (O_12,N_29930,N_29561);
nor UO_13 (O_13,N_29787,N_29748);
or UO_14 (O_14,N_29886,N_29798);
nor UO_15 (O_15,N_29909,N_29501);
xnor UO_16 (O_16,N_29857,N_29799);
xnor UO_17 (O_17,N_29975,N_29692);
and UO_18 (O_18,N_29821,N_29574);
and UO_19 (O_19,N_29573,N_29990);
nand UO_20 (O_20,N_29685,N_29859);
nor UO_21 (O_21,N_29987,N_29582);
and UO_22 (O_22,N_29522,N_29593);
and UO_23 (O_23,N_29598,N_29550);
or UO_24 (O_24,N_29735,N_29669);
or UO_25 (O_25,N_29919,N_29750);
or UO_26 (O_26,N_29972,N_29914);
or UO_27 (O_27,N_29786,N_29584);
xor UO_28 (O_28,N_29768,N_29892);
nor UO_29 (O_29,N_29700,N_29648);
and UO_30 (O_30,N_29915,N_29929);
xor UO_31 (O_31,N_29873,N_29643);
or UO_32 (O_32,N_29537,N_29592);
nand UO_33 (O_33,N_29704,N_29994);
and UO_34 (O_34,N_29870,N_29809);
xnor UO_35 (O_35,N_29781,N_29846);
or UO_36 (O_36,N_29536,N_29594);
or UO_37 (O_37,N_29698,N_29960);
or UO_38 (O_38,N_29689,N_29562);
or UO_39 (O_39,N_29503,N_29568);
nor UO_40 (O_40,N_29931,N_29741);
or UO_41 (O_41,N_29844,N_29955);
nor UO_42 (O_42,N_29595,N_29811);
xnor UO_43 (O_43,N_29634,N_29625);
nand UO_44 (O_44,N_29645,N_29507);
xor UO_45 (O_45,N_29693,N_29564);
nor UO_46 (O_46,N_29519,N_29928);
nor UO_47 (O_47,N_29812,N_29856);
nor UO_48 (O_48,N_29826,N_29765);
or UO_49 (O_49,N_29899,N_29606);
nand UO_50 (O_50,N_29957,N_29604);
and UO_51 (O_51,N_29728,N_29618);
or UO_52 (O_52,N_29862,N_29706);
nand UO_53 (O_53,N_29726,N_29684);
and UO_54 (O_54,N_29679,N_29800);
xor UO_55 (O_55,N_29942,N_29926);
nand UO_56 (O_56,N_29767,N_29512);
and UO_57 (O_57,N_29657,N_29622);
nor UO_58 (O_58,N_29916,N_29756);
or UO_59 (O_59,N_29934,N_29514);
xnor UO_60 (O_60,N_29631,N_29515);
nor UO_61 (O_61,N_29690,N_29729);
and UO_62 (O_62,N_29526,N_29713);
xnor UO_63 (O_63,N_29790,N_29829);
or UO_64 (O_64,N_29753,N_29673);
or UO_65 (O_65,N_29570,N_29939);
nor UO_66 (O_66,N_29907,N_29981);
xnor UO_67 (O_67,N_29985,N_29810);
xor UO_68 (O_68,N_29553,N_29817);
or UO_69 (O_69,N_29612,N_29749);
nand UO_70 (O_70,N_29897,N_29794);
nand UO_71 (O_71,N_29961,N_29746);
or UO_72 (O_72,N_29864,N_29656);
nor UO_73 (O_73,N_29983,N_29991);
and UO_74 (O_74,N_29950,N_29971);
nand UO_75 (O_75,N_29855,N_29941);
and UO_76 (O_76,N_29544,N_29615);
nand UO_77 (O_77,N_29658,N_29703);
nand UO_78 (O_78,N_29517,N_29903);
or UO_79 (O_79,N_29774,N_29633);
nand UO_80 (O_80,N_29640,N_29761);
or UO_81 (O_81,N_29986,N_29823);
and UO_82 (O_82,N_29565,N_29725);
xnor UO_83 (O_83,N_29576,N_29718);
or UO_84 (O_84,N_29874,N_29940);
nor UO_85 (O_85,N_29865,N_29629);
and UO_86 (O_86,N_29552,N_29732);
nand UO_87 (O_87,N_29752,N_29827);
and UO_88 (O_88,N_29954,N_29947);
xnor UO_89 (O_89,N_29951,N_29912);
nand UO_90 (O_90,N_29569,N_29647);
or UO_91 (O_91,N_29599,N_29624);
nor UO_92 (O_92,N_29807,N_29816);
or UO_93 (O_93,N_29567,N_29614);
and UO_94 (O_94,N_29714,N_29575);
and UO_95 (O_95,N_29683,N_29970);
and UO_96 (O_96,N_29720,N_29998);
nor UO_97 (O_97,N_29688,N_29742);
nor UO_98 (O_98,N_29850,N_29922);
nor UO_99 (O_99,N_29952,N_29836);
or UO_100 (O_100,N_29762,N_29992);
nand UO_101 (O_101,N_29989,N_29893);
nor UO_102 (O_102,N_29905,N_29508);
nand UO_103 (O_103,N_29521,N_29910);
nand UO_104 (O_104,N_29997,N_29891);
nand UO_105 (O_105,N_29597,N_29695);
nand UO_106 (O_106,N_29847,N_29852);
or UO_107 (O_107,N_29697,N_29819);
and UO_108 (O_108,N_29721,N_29801);
nand UO_109 (O_109,N_29835,N_29825);
and UO_110 (O_110,N_29506,N_29660);
xor UO_111 (O_111,N_29666,N_29712);
nand UO_112 (O_112,N_29995,N_29853);
or UO_113 (O_113,N_29839,N_29655);
nand UO_114 (O_114,N_29775,N_29830);
nand UO_115 (O_115,N_29636,N_29982);
nand UO_116 (O_116,N_29806,N_29523);
and UO_117 (O_117,N_29535,N_29722);
nor UO_118 (O_118,N_29945,N_29671);
xor UO_119 (O_119,N_29984,N_29956);
or UO_120 (O_120,N_29791,N_29937);
nand UO_121 (O_121,N_29757,N_29737);
and UO_122 (O_122,N_29820,N_29818);
and UO_123 (O_123,N_29670,N_29642);
or UO_124 (O_124,N_29878,N_29557);
nor UO_125 (O_125,N_29858,N_29938);
or UO_126 (O_126,N_29845,N_29571);
and UO_127 (O_127,N_29534,N_29682);
or UO_128 (O_128,N_29964,N_29920);
and UO_129 (O_129,N_29841,N_29911);
nand UO_130 (O_130,N_29978,N_29663);
and UO_131 (O_131,N_29860,N_29867);
nand UO_132 (O_132,N_29927,N_29711);
nand UO_133 (O_133,N_29667,N_29556);
xor UO_134 (O_134,N_29677,N_29848);
nand UO_135 (O_135,N_29805,N_29739);
xor UO_136 (O_136,N_29751,N_29918);
nor UO_137 (O_137,N_29585,N_29933);
nor UO_138 (O_138,N_29963,N_29861);
nand UO_139 (O_139,N_29516,N_29548);
nand UO_140 (O_140,N_29935,N_29600);
xnor UO_141 (O_141,N_29894,N_29745);
or UO_142 (O_142,N_29500,N_29730);
or UO_143 (O_143,N_29646,N_29771);
and UO_144 (O_144,N_29763,N_29780);
xnor UO_145 (O_145,N_29590,N_29976);
nand UO_146 (O_146,N_29546,N_29959);
or UO_147 (O_147,N_29779,N_29551);
nor UO_148 (O_148,N_29943,N_29587);
and UO_149 (O_149,N_29898,N_29999);
nor UO_150 (O_150,N_29843,N_29889);
xnor UO_151 (O_151,N_29502,N_29731);
xor UO_152 (O_152,N_29627,N_29702);
and UO_153 (O_153,N_29803,N_29686);
nor UO_154 (O_154,N_29504,N_29542);
and UO_155 (O_155,N_29630,N_29789);
nand UO_156 (O_156,N_29532,N_29513);
and UO_157 (O_157,N_29871,N_29738);
xor UO_158 (O_158,N_29883,N_29724);
and UO_159 (O_159,N_29900,N_29896);
xor UO_160 (O_160,N_29773,N_29675);
and UO_161 (O_161,N_29511,N_29733);
and UO_162 (O_162,N_29795,N_29545);
xnor UO_163 (O_163,N_29815,N_29530);
xnor UO_164 (O_164,N_29838,N_29525);
xor UO_165 (O_165,N_29736,N_29635);
nand UO_166 (O_166,N_29908,N_29895);
or UO_167 (O_167,N_29958,N_29709);
nor UO_168 (O_168,N_29681,N_29904);
nand UO_169 (O_169,N_29837,N_29876);
nand UO_170 (O_170,N_29993,N_29572);
xor UO_171 (O_171,N_29601,N_29701);
nand UO_172 (O_172,N_29694,N_29814);
nand UO_173 (O_173,N_29988,N_29560);
or UO_174 (O_174,N_29887,N_29699);
nand UO_175 (O_175,N_29849,N_29792);
or UO_176 (O_176,N_29832,N_29758);
xor UO_177 (O_177,N_29890,N_29868);
xnor UO_178 (O_178,N_29659,N_29788);
nor UO_179 (O_179,N_29558,N_29880);
nor UO_180 (O_180,N_29885,N_29577);
nand UO_181 (O_181,N_29901,N_29678);
nand UO_182 (O_182,N_29609,N_29539);
and UO_183 (O_183,N_29651,N_29628);
nor UO_184 (O_184,N_29676,N_29632);
nand UO_185 (O_185,N_29769,N_29638);
nor UO_186 (O_186,N_29527,N_29840);
xor UO_187 (O_187,N_29654,N_29872);
xnor UO_188 (O_188,N_29596,N_29533);
or UO_189 (O_189,N_29962,N_29580);
nand UO_190 (O_190,N_29608,N_29854);
xor UO_191 (O_191,N_29793,N_29969);
or UO_192 (O_192,N_29649,N_29979);
or UO_193 (O_193,N_29672,N_29974);
xor UO_194 (O_194,N_29824,N_29644);
nand UO_195 (O_195,N_29591,N_29586);
xnor UO_196 (O_196,N_29509,N_29917);
or UO_197 (O_197,N_29833,N_29716);
and UO_198 (O_198,N_29881,N_29973);
xnor UO_199 (O_199,N_29538,N_29804);
nand UO_200 (O_200,N_29747,N_29932);
nor UO_201 (O_201,N_29796,N_29579);
nand UO_202 (O_202,N_29866,N_29547);
nor UO_203 (O_203,N_29875,N_29921);
nand UO_204 (O_204,N_29639,N_29802);
xor UO_205 (O_205,N_29664,N_29652);
and UO_206 (O_206,N_29616,N_29842);
nand UO_207 (O_207,N_29863,N_29581);
nand UO_208 (O_208,N_29783,N_29583);
nand UO_209 (O_209,N_29770,N_29784);
and UO_210 (O_210,N_29902,N_29661);
or UO_211 (O_211,N_29529,N_29520);
xnor UO_212 (O_212,N_29611,N_29674);
xor UO_213 (O_213,N_29882,N_29717);
nand UO_214 (O_214,N_29888,N_29707);
xor UO_215 (O_215,N_29563,N_29923);
nor UO_216 (O_216,N_29528,N_29764);
nor UO_217 (O_217,N_29936,N_29549);
nand UO_218 (O_218,N_29723,N_29641);
xnor UO_219 (O_219,N_29662,N_29965);
nor UO_220 (O_220,N_29543,N_29778);
or UO_221 (O_221,N_29879,N_29602);
and UO_222 (O_222,N_29589,N_29605);
nand UO_223 (O_223,N_29623,N_29588);
xnor UO_224 (O_224,N_29617,N_29869);
xor UO_225 (O_225,N_29559,N_29668);
xor UO_226 (O_226,N_29996,N_29653);
nor UO_227 (O_227,N_29766,N_29743);
or UO_228 (O_228,N_29777,N_29719);
or UO_229 (O_229,N_29687,N_29696);
or UO_230 (O_230,N_29946,N_29740);
nor UO_231 (O_231,N_29822,N_29620);
or UO_232 (O_232,N_29968,N_29755);
and UO_233 (O_233,N_29754,N_29744);
xnor UO_234 (O_234,N_29948,N_29785);
xnor UO_235 (O_235,N_29797,N_29828);
xnor UO_236 (O_236,N_29977,N_29650);
xnor UO_237 (O_237,N_29710,N_29851);
xor UO_238 (O_238,N_29834,N_29510);
or UO_239 (O_239,N_29808,N_29531);
and UO_240 (O_240,N_29759,N_29913);
or UO_241 (O_241,N_29949,N_29924);
or UO_242 (O_242,N_29578,N_29621);
nor UO_243 (O_243,N_29637,N_29727);
nor UO_244 (O_244,N_29603,N_29715);
xor UO_245 (O_245,N_29944,N_29772);
and UO_246 (O_246,N_29541,N_29953);
and UO_247 (O_247,N_29980,N_29613);
nor UO_248 (O_248,N_29691,N_29776);
and UO_249 (O_249,N_29708,N_29884);
xnor UO_250 (O_250,N_29865,N_29592);
nor UO_251 (O_251,N_29928,N_29951);
nand UO_252 (O_252,N_29837,N_29525);
or UO_253 (O_253,N_29663,N_29602);
or UO_254 (O_254,N_29679,N_29845);
and UO_255 (O_255,N_29986,N_29942);
and UO_256 (O_256,N_29891,N_29533);
nor UO_257 (O_257,N_29533,N_29768);
or UO_258 (O_258,N_29984,N_29660);
or UO_259 (O_259,N_29787,N_29705);
nand UO_260 (O_260,N_29981,N_29821);
and UO_261 (O_261,N_29994,N_29505);
nand UO_262 (O_262,N_29739,N_29554);
nand UO_263 (O_263,N_29841,N_29940);
and UO_264 (O_264,N_29774,N_29506);
nand UO_265 (O_265,N_29664,N_29820);
nand UO_266 (O_266,N_29986,N_29598);
and UO_267 (O_267,N_29953,N_29986);
and UO_268 (O_268,N_29546,N_29596);
nor UO_269 (O_269,N_29957,N_29528);
nand UO_270 (O_270,N_29638,N_29743);
nor UO_271 (O_271,N_29913,N_29944);
nor UO_272 (O_272,N_29579,N_29662);
xnor UO_273 (O_273,N_29922,N_29762);
xnor UO_274 (O_274,N_29532,N_29621);
nor UO_275 (O_275,N_29876,N_29784);
nand UO_276 (O_276,N_29704,N_29978);
nand UO_277 (O_277,N_29636,N_29658);
nand UO_278 (O_278,N_29882,N_29854);
nor UO_279 (O_279,N_29824,N_29878);
nand UO_280 (O_280,N_29587,N_29739);
xor UO_281 (O_281,N_29643,N_29668);
xor UO_282 (O_282,N_29962,N_29608);
nand UO_283 (O_283,N_29592,N_29788);
xnor UO_284 (O_284,N_29979,N_29624);
or UO_285 (O_285,N_29979,N_29673);
and UO_286 (O_286,N_29546,N_29572);
or UO_287 (O_287,N_29508,N_29845);
or UO_288 (O_288,N_29934,N_29624);
nor UO_289 (O_289,N_29969,N_29710);
nand UO_290 (O_290,N_29993,N_29577);
and UO_291 (O_291,N_29957,N_29845);
nor UO_292 (O_292,N_29848,N_29702);
nand UO_293 (O_293,N_29541,N_29956);
or UO_294 (O_294,N_29678,N_29950);
or UO_295 (O_295,N_29560,N_29971);
nand UO_296 (O_296,N_29512,N_29516);
or UO_297 (O_297,N_29828,N_29981);
and UO_298 (O_298,N_29840,N_29756);
nand UO_299 (O_299,N_29554,N_29654);
and UO_300 (O_300,N_29791,N_29892);
nor UO_301 (O_301,N_29534,N_29925);
nand UO_302 (O_302,N_29730,N_29822);
nand UO_303 (O_303,N_29726,N_29825);
xnor UO_304 (O_304,N_29805,N_29761);
or UO_305 (O_305,N_29648,N_29827);
xnor UO_306 (O_306,N_29572,N_29976);
and UO_307 (O_307,N_29507,N_29748);
nand UO_308 (O_308,N_29682,N_29513);
xnor UO_309 (O_309,N_29790,N_29955);
nor UO_310 (O_310,N_29665,N_29958);
and UO_311 (O_311,N_29565,N_29677);
nand UO_312 (O_312,N_29791,N_29687);
nand UO_313 (O_313,N_29727,N_29996);
xor UO_314 (O_314,N_29592,N_29535);
nand UO_315 (O_315,N_29942,N_29742);
nor UO_316 (O_316,N_29957,N_29623);
nor UO_317 (O_317,N_29914,N_29947);
nand UO_318 (O_318,N_29665,N_29587);
or UO_319 (O_319,N_29596,N_29863);
or UO_320 (O_320,N_29941,N_29659);
xnor UO_321 (O_321,N_29581,N_29807);
or UO_322 (O_322,N_29913,N_29752);
and UO_323 (O_323,N_29857,N_29806);
or UO_324 (O_324,N_29711,N_29632);
nand UO_325 (O_325,N_29560,N_29642);
nor UO_326 (O_326,N_29568,N_29540);
xor UO_327 (O_327,N_29774,N_29977);
or UO_328 (O_328,N_29590,N_29598);
xnor UO_329 (O_329,N_29636,N_29518);
xor UO_330 (O_330,N_29626,N_29961);
or UO_331 (O_331,N_29953,N_29835);
and UO_332 (O_332,N_29589,N_29672);
or UO_333 (O_333,N_29562,N_29840);
xor UO_334 (O_334,N_29859,N_29548);
xnor UO_335 (O_335,N_29702,N_29793);
xnor UO_336 (O_336,N_29864,N_29765);
and UO_337 (O_337,N_29753,N_29823);
nor UO_338 (O_338,N_29508,N_29858);
nor UO_339 (O_339,N_29943,N_29534);
xor UO_340 (O_340,N_29693,N_29815);
xor UO_341 (O_341,N_29785,N_29725);
or UO_342 (O_342,N_29950,N_29765);
nor UO_343 (O_343,N_29838,N_29901);
nor UO_344 (O_344,N_29678,N_29709);
nor UO_345 (O_345,N_29676,N_29612);
and UO_346 (O_346,N_29595,N_29583);
and UO_347 (O_347,N_29519,N_29834);
nor UO_348 (O_348,N_29522,N_29603);
nor UO_349 (O_349,N_29580,N_29764);
and UO_350 (O_350,N_29792,N_29566);
xnor UO_351 (O_351,N_29503,N_29997);
nor UO_352 (O_352,N_29684,N_29981);
and UO_353 (O_353,N_29979,N_29984);
nand UO_354 (O_354,N_29734,N_29514);
nor UO_355 (O_355,N_29767,N_29866);
nor UO_356 (O_356,N_29952,N_29828);
xor UO_357 (O_357,N_29965,N_29617);
or UO_358 (O_358,N_29658,N_29971);
xnor UO_359 (O_359,N_29519,N_29830);
nor UO_360 (O_360,N_29990,N_29731);
xnor UO_361 (O_361,N_29954,N_29545);
or UO_362 (O_362,N_29846,N_29854);
nor UO_363 (O_363,N_29686,N_29547);
and UO_364 (O_364,N_29588,N_29770);
nand UO_365 (O_365,N_29916,N_29904);
nor UO_366 (O_366,N_29560,N_29703);
nand UO_367 (O_367,N_29516,N_29635);
nor UO_368 (O_368,N_29702,N_29976);
or UO_369 (O_369,N_29792,N_29514);
xor UO_370 (O_370,N_29851,N_29731);
nor UO_371 (O_371,N_29798,N_29860);
nand UO_372 (O_372,N_29817,N_29688);
nor UO_373 (O_373,N_29978,N_29944);
nand UO_374 (O_374,N_29828,N_29768);
xor UO_375 (O_375,N_29653,N_29854);
nand UO_376 (O_376,N_29816,N_29743);
xnor UO_377 (O_377,N_29578,N_29952);
and UO_378 (O_378,N_29743,N_29998);
xor UO_379 (O_379,N_29956,N_29818);
nor UO_380 (O_380,N_29727,N_29522);
nor UO_381 (O_381,N_29508,N_29585);
nor UO_382 (O_382,N_29660,N_29781);
nor UO_383 (O_383,N_29911,N_29715);
or UO_384 (O_384,N_29875,N_29763);
or UO_385 (O_385,N_29736,N_29803);
and UO_386 (O_386,N_29818,N_29753);
nand UO_387 (O_387,N_29866,N_29724);
nor UO_388 (O_388,N_29869,N_29939);
and UO_389 (O_389,N_29924,N_29663);
and UO_390 (O_390,N_29875,N_29854);
nand UO_391 (O_391,N_29779,N_29757);
nor UO_392 (O_392,N_29964,N_29899);
nand UO_393 (O_393,N_29667,N_29749);
or UO_394 (O_394,N_29953,N_29748);
nor UO_395 (O_395,N_29505,N_29680);
nand UO_396 (O_396,N_29692,N_29958);
or UO_397 (O_397,N_29912,N_29504);
xnor UO_398 (O_398,N_29845,N_29706);
and UO_399 (O_399,N_29798,N_29981);
nor UO_400 (O_400,N_29758,N_29780);
xnor UO_401 (O_401,N_29934,N_29832);
or UO_402 (O_402,N_29630,N_29586);
xor UO_403 (O_403,N_29786,N_29672);
xnor UO_404 (O_404,N_29785,N_29586);
or UO_405 (O_405,N_29748,N_29983);
or UO_406 (O_406,N_29728,N_29547);
nand UO_407 (O_407,N_29567,N_29584);
and UO_408 (O_408,N_29980,N_29500);
nor UO_409 (O_409,N_29602,N_29604);
nand UO_410 (O_410,N_29859,N_29504);
or UO_411 (O_411,N_29784,N_29963);
nand UO_412 (O_412,N_29814,N_29926);
xnor UO_413 (O_413,N_29749,N_29584);
or UO_414 (O_414,N_29622,N_29828);
nand UO_415 (O_415,N_29502,N_29735);
and UO_416 (O_416,N_29972,N_29558);
xor UO_417 (O_417,N_29568,N_29797);
or UO_418 (O_418,N_29641,N_29816);
and UO_419 (O_419,N_29713,N_29747);
nor UO_420 (O_420,N_29584,N_29948);
nor UO_421 (O_421,N_29797,N_29827);
or UO_422 (O_422,N_29932,N_29912);
or UO_423 (O_423,N_29632,N_29733);
xnor UO_424 (O_424,N_29846,N_29957);
and UO_425 (O_425,N_29678,N_29636);
or UO_426 (O_426,N_29646,N_29668);
nand UO_427 (O_427,N_29718,N_29602);
xnor UO_428 (O_428,N_29679,N_29954);
and UO_429 (O_429,N_29856,N_29704);
nor UO_430 (O_430,N_29827,N_29765);
xnor UO_431 (O_431,N_29603,N_29625);
nor UO_432 (O_432,N_29758,N_29528);
nor UO_433 (O_433,N_29789,N_29957);
xor UO_434 (O_434,N_29982,N_29686);
or UO_435 (O_435,N_29844,N_29868);
nand UO_436 (O_436,N_29678,N_29509);
and UO_437 (O_437,N_29665,N_29544);
or UO_438 (O_438,N_29715,N_29843);
and UO_439 (O_439,N_29915,N_29543);
and UO_440 (O_440,N_29644,N_29533);
nor UO_441 (O_441,N_29725,N_29603);
xnor UO_442 (O_442,N_29701,N_29766);
and UO_443 (O_443,N_29657,N_29534);
nand UO_444 (O_444,N_29771,N_29698);
and UO_445 (O_445,N_29615,N_29652);
nand UO_446 (O_446,N_29833,N_29794);
nor UO_447 (O_447,N_29877,N_29529);
xnor UO_448 (O_448,N_29945,N_29787);
and UO_449 (O_449,N_29894,N_29608);
nor UO_450 (O_450,N_29961,N_29868);
nand UO_451 (O_451,N_29556,N_29665);
and UO_452 (O_452,N_29989,N_29799);
nand UO_453 (O_453,N_29900,N_29529);
xnor UO_454 (O_454,N_29921,N_29526);
nand UO_455 (O_455,N_29553,N_29978);
nor UO_456 (O_456,N_29550,N_29962);
or UO_457 (O_457,N_29507,N_29835);
and UO_458 (O_458,N_29840,N_29806);
nor UO_459 (O_459,N_29748,N_29724);
or UO_460 (O_460,N_29664,N_29536);
xor UO_461 (O_461,N_29858,N_29999);
or UO_462 (O_462,N_29635,N_29514);
xnor UO_463 (O_463,N_29677,N_29958);
xor UO_464 (O_464,N_29952,N_29547);
nand UO_465 (O_465,N_29666,N_29581);
nand UO_466 (O_466,N_29670,N_29729);
nor UO_467 (O_467,N_29672,N_29870);
nor UO_468 (O_468,N_29753,N_29674);
nor UO_469 (O_469,N_29639,N_29587);
and UO_470 (O_470,N_29802,N_29641);
nand UO_471 (O_471,N_29850,N_29689);
nor UO_472 (O_472,N_29671,N_29750);
xor UO_473 (O_473,N_29991,N_29509);
nor UO_474 (O_474,N_29705,N_29808);
xor UO_475 (O_475,N_29641,N_29662);
and UO_476 (O_476,N_29623,N_29956);
nor UO_477 (O_477,N_29726,N_29573);
xnor UO_478 (O_478,N_29743,N_29857);
nor UO_479 (O_479,N_29929,N_29536);
xnor UO_480 (O_480,N_29630,N_29607);
or UO_481 (O_481,N_29891,N_29563);
xor UO_482 (O_482,N_29716,N_29576);
xnor UO_483 (O_483,N_29642,N_29982);
or UO_484 (O_484,N_29521,N_29659);
and UO_485 (O_485,N_29783,N_29814);
or UO_486 (O_486,N_29903,N_29834);
and UO_487 (O_487,N_29779,N_29663);
or UO_488 (O_488,N_29521,N_29985);
or UO_489 (O_489,N_29700,N_29726);
xor UO_490 (O_490,N_29912,N_29603);
nand UO_491 (O_491,N_29880,N_29834);
xor UO_492 (O_492,N_29735,N_29729);
nor UO_493 (O_493,N_29766,N_29585);
or UO_494 (O_494,N_29947,N_29513);
or UO_495 (O_495,N_29567,N_29652);
nor UO_496 (O_496,N_29631,N_29815);
nand UO_497 (O_497,N_29957,N_29588);
xor UO_498 (O_498,N_29506,N_29809);
xor UO_499 (O_499,N_29844,N_29985);
xor UO_500 (O_500,N_29902,N_29743);
or UO_501 (O_501,N_29563,N_29875);
nand UO_502 (O_502,N_29936,N_29777);
nand UO_503 (O_503,N_29941,N_29859);
nor UO_504 (O_504,N_29510,N_29644);
nor UO_505 (O_505,N_29891,N_29896);
nor UO_506 (O_506,N_29681,N_29935);
nand UO_507 (O_507,N_29861,N_29633);
or UO_508 (O_508,N_29933,N_29720);
nor UO_509 (O_509,N_29685,N_29884);
nor UO_510 (O_510,N_29755,N_29773);
and UO_511 (O_511,N_29701,N_29579);
nand UO_512 (O_512,N_29736,N_29926);
or UO_513 (O_513,N_29865,N_29893);
nand UO_514 (O_514,N_29714,N_29681);
nor UO_515 (O_515,N_29525,N_29518);
xor UO_516 (O_516,N_29684,N_29913);
and UO_517 (O_517,N_29812,N_29818);
nor UO_518 (O_518,N_29912,N_29685);
nor UO_519 (O_519,N_29821,N_29774);
and UO_520 (O_520,N_29947,N_29748);
and UO_521 (O_521,N_29705,N_29805);
nand UO_522 (O_522,N_29896,N_29849);
nand UO_523 (O_523,N_29674,N_29720);
nor UO_524 (O_524,N_29950,N_29520);
xor UO_525 (O_525,N_29813,N_29847);
nand UO_526 (O_526,N_29842,N_29586);
nor UO_527 (O_527,N_29633,N_29545);
nand UO_528 (O_528,N_29802,N_29710);
or UO_529 (O_529,N_29631,N_29911);
or UO_530 (O_530,N_29715,N_29879);
xnor UO_531 (O_531,N_29953,N_29561);
nor UO_532 (O_532,N_29581,N_29995);
nand UO_533 (O_533,N_29776,N_29975);
nand UO_534 (O_534,N_29852,N_29707);
or UO_535 (O_535,N_29714,N_29667);
nor UO_536 (O_536,N_29832,N_29625);
nor UO_537 (O_537,N_29853,N_29814);
or UO_538 (O_538,N_29843,N_29926);
xor UO_539 (O_539,N_29516,N_29952);
nor UO_540 (O_540,N_29943,N_29869);
and UO_541 (O_541,N_29573,N_29603);
or UO_542 (O_542,N_29735,N_29734);
nand UO_543 (O_543,N_29573,N_29548);
nor UO_544 (O_544,N_29740,N_29701);
and UO_545 (O_545,N_29514,N_29888);
and UO_546 (O_546,N_29827,N_29555);
and UO_547 (O_547,N_29626,N_29801);
nand UO_548 (O_548,N_29560,N_29621);
nor UO_549 (O_549,N_29513,N_29652);
nand UO_550 (O_550,N_29879,N_29562);
and UO_551 (O_551,N_29782,N_29626);
nand UO_552 (O_552,N_29603,N_29572);
xnor UO_553 (O_553,N_29507,N_29539);
nand UO_554 (O_554,N_29909,N_29913);
nand UO_555 (O_555,N_29984,N_29722);
or UO_556 (O_556,N_29573,N_29595);
nand UO_557 (O_557,N_29632,N_29859);
nand UO_558 (O_558,N_29638,N_29709);
nand UO_559 (O_559,N_29515,N_29684);
or UO_560 (O_560,N_29840,N_29990);
nand UO_561 (O_561,N_29566,N_29760);
nand UO_562 (O_562,N_29622,N_29762);
and UO_563 (O_563,N_29641,N_29973);
xor UO_564 (O_564,N_29997,N_29570);
xor UO_565 (O_565,N_29831,N_29703);
nor UO_566 (O_566,N_29542,N_29743);
or UO_567 (O_567,N_29871,N_29824);
nor UO_568 (O_568,N_29667,N_29763);
nand UO_569 (O_569,N_29801,N_29882);
nand UO_570 (O_570,N_29807,N_29788);
or UO_571 (O_571,N_29662,N_29766);
xor UO_572 (O_572,N_29534,N_29931);
nand UO_573 (O_573,N_29910,N_29726);
nand UO_574 (O_574,N_29888,N_29630);
nand UO_575 (O_575,N_29689,N_29888);
or UO_576 (O_576,N_29582,N_29587);
and UO_577 (O_577,N_29817,N_29896);
and UO_578 (O_578,N_29594,N_29895);
or UO_579 (O_579,N_29623,N_29931);
xor UO_580 (O_580,N_29571,N_29670);
xnor UO_581 (O_581,N_29594,N_29797);
or UO_582 (O_582,N_29720,N_29716);
and UO_583 (O_583,N_29675,N_29897);
and UO_584 (O_584,N_29925,N_29883);
xor UO_585 (O_585,N_29776,N_29596);
xor UO_586 (O_586,N_29863,N_29764);
or UO_587 (O_587,N_29998,N_29591);
or UO_588 (O_588,N_29958,N_29809);
and UO_589 (O_589,N_29801,N_29565);
xnor UO_590 (O_590,N_29958,N_29706);
or UO_591 (O_591,N_29944,N_29961);
or UO_592 (O_592,N_29713,N_29889);
and UO_593 (O_593,N_29731,N_29939);
or UO_594 (O_594,N_29865,N_29963);
xnor UO_595 (O_595,N_29770,N_29746);
or UO_596 (O_596,N_29546,N_29979);
xnor UO_597 (O_597,N_29600,N_29704);
xnor UO_598 (O_598,N_29836,N_29941);
or UO_599 (O_599,N_29593,N_29934);
nand UO_600 (O_600,N_29597,N_29786);
nor UO_601 (O_601,N_29548,N_29923);
nor UO_602 (O_602,N_29991,N_29953);
or UO_603 (O_603,N_29535,N_29795);
and UO_604 (O_604,N_29987,N_29992);
nand UO_605 (O_605,N_29754,N_29527);
nand UO_606 (O_606,N_29691,N_29803);
xor UO_607 (O_607,N_29756,N_29779);
nand UO_608 (O_608,N_29673,N_29931);
xor UO_609 (O_609,N_29607,N_29713);
xor UO_610 (O_610,N_29681,N_29721);
xor UO_611 (O_611,N_29748,N_29622);
nor UO_612 (O_612,N_29906,N_29513);
nor UO_613 (O_613,N_29819,N_29741);
or UO_614 (O_614,N_29626,N_29748);
or UO_615 (O_615,N_29506,N_29643);
xnor UO_616 (O_616,N_29687,N_29686);
nor UO_617 (O_617,N_29578,N_29634);
xor UO_618 (O_618,N_29884,N_29741);
nor UO_619 (O_619,N_29790,N_29755);
or UO_620 (O_620,N_29831,N_29694);
nor UO_621 (O_621,N_29796,N_29757);
or UO_622 (O_622,N_29520,N_29599);
xor UO_623 (O_623,N_29724,N_29936);
xor UO_624 (O_624,N_29507,N_29747);
nor UO_625 (O_625,N_29950,N_29781);
or UO_626 (O_626,N_29645,N_29608);
xnor UO_627 (O_627,N_29581,N_29503);
xor UO_628 (O_628,N_29632,N_29509);
xor UO_629 (O_629,N_29664,N_29934);
xnor UO_630 (O_630,N_29528,N_29752);
nor UO_631 (O_631,N_29700,N_29886);
nand UO_632 (O_632,N_29878,N_29526);
xnor UO_633 (O_633,N_29886,N_29610);
nor UO_634 (O_634,N_29526,N_29630);
or UO_635 (O_635,N_29724,N_29514);
or UO_636 (O_636,N_29675,N_29978);
nand UO_637 (O_637,N_29925,N_29828);
nor UO_638 (O_638,N_29720,N_29578);
xnor UO_639 (O_639,N_29599,N_29566);
and UO_640 (O_640,N_29767,N_29553);
nor UO_641 (O_641,N_29575,N_29987);
nor UO_642 (O_642,N_29704,N_29640);
xor UO_643 (O_643,N_29941,N_29605);
nand UO_644 (O_644,N_29647,N_29523);
nand UO_645 (O_645,N_29519,N_29819);
and UO_646 (O_646,N_29954,N_29721);
and UO_647 (O_647,N_29661,N_29726);
and UO_648 (O_648,N_29951,N_29966);
nand UO_649 (O_649,N_29645,N_29681);
xor UO_650 (O_650,N_29616,N_29868);
xor UO_651 (O_651,N_29775,N_29851);
xor UO_652 (O_652,N_29909,N_29612);
nand UO_653 (O_653,N_29718,N_29882);
nand UO_654 (O_654,N_29560,N_29672);
nor UO_655 (O_655,N_29874,N_29991);
nand UO_656 (O_656,N_29519,N_29849);
and UO_657 (O_657,N_29997,N_29602);
nand UO_658 (O_658,N_29694,N_29844);
nand UO_659 (O_659,N_29791,N_29977);
xnor UO_660 (O_660,N_29526,N_29539);
nand UO_661 (O_661,N_29650,N_29906);
nand UO_662 (O_662,N_29549,N_29509);
xor UO_663 (O_663,N_29872,N_29677);
xnor UO_664 (O_664,N_29680,N_29630);
and UO_665 (O_665,N_29714,N_29699);
and UO_666 (O_666,N_29927,N_29818);
nand UO_667 (O_667,N_29768,N_29711);
nand UO_668 (O_668,N_29656,N_29584);
and UO_669 (O_669,N_29930,N_29922);
xnor UO_670 (O_670,N_29622,N_29566);
or UO_671 (O_671,N_29800,N_29674);
nor UO_672 (O_672,N_29519,N_29821);
nor UO_673 (O_673,N_29860,N_29671);
xnor UO_674 (O_674,N_29507,N_29846);
nor UO_675 (O_675,N_29510,N_29642);
and UO_676 (O_676,N_29871,N_29680);
xnor UO_677 (O_677,N_29635,N_29605);
and UO_678 (O_678,N_29756,N_29530);
and UO_679 (O_679,N_29561,N_29960);
and UO_680 (O_680,N_29741,N_29929);
xnor UO_681 (O_681,N_29931,N_29923);
or UO_682 (O_682,N_29703,N_29791);
xnor UO_683 (O_683,N_29528,N_29538);
or UO_684 (O_684,N_29864,N_29583);
xnor UO_685 (O_685,N_29608,N_29574);
and UO_686 (O_686,N_29659,N_29601);
or UO_687 (O_687,N_29531,N_29648);
and UO_688 (O_688,N_29948,N_29743);
nand UO_689 (O_689,N_29997,N_29514);
or UO_690 (O_690,N_29555,N_29901);
or UO_691 (O_691,N_29948,N_29651);
or UO_692 (O_692,N_29605,N_29593);
xor UO_693 (O_693,N_29861,N_29847);
nor UO_694 (O_694,N_29788,N_29608);
nand UO_695 (O_695,N_29981,N_29897);
or UO_696 (O_696,N_29548,N_29630);
nor UO_697 (O_697,N_29896,N_29836);
or UO_698 (O_698,N_29752,N_29575);
or UO_699 (O_699,N_29710,N_29901);
nand UO_700 (O_700,N_29856,N_29731);
nor UO_701 (O_701,N_29897,N_29861);
xnor UO_702 (O_702,N_29719,N_29650);
xnor UO_703 (O_703,N_29503,N_29710);
or UO_704 (O_704,N_29926,N_29755);
nor UO_705 (O_705,N_29645,N_29881);
nand UO_706 (O_706,N_29949,N_29922);
and UO_707 (O_707,N_29573,N_29985);
xor UO_708 (O_708,N_29601,N_29942);
nand UO_709 (O_709,N_29916,N_29655);
xor UO_710 (O_710,N_29874,N_29823);
nand UO_711 (O_711,N_29876,N_29952);
or UO_712 (O_712,N_29685,N_29767);
and UO_713 (O_713,N_29815,N_29765);
xor UO_714 (O_714,N_29525,N_29917);
nand UO_715 (O_715,N_29759,N_29540);
nor UO_716 (O_716,N_29588,N_29643);
nand UO_717 (O_717,N_29697,N_29809);
xnor UO_718 (O_718,N_29988,N_29855);
xnor UO_719 (O_719,N_29589,N_29775);
and UO_720 (O_720,N_29816,N_29574);
nor UO_721 (O_721,N_29618,N_29819);
nand UO_722 (O_722,N_29654,N_29717);
nand UO_723 (O_723,N_29517,N_29541);
xnor UO_724 (O_724,N_29666,N_29769);
or UO_725 (O_725,N_29731,N_29547);
and UO_726 (O_726,N_29993,N_29717);
nand UO_727 (O_727,N_29773,N_29726);
xnor UO_728 (O_728,N_29907,N_29681);
nor UO_729 (O_729,N_29761,N_29753);
nor UO_730 (O_730,N_29564,N_29680);
nand UO_731 (O_731,N_29912,N_29943);
or UO_732 (O_732,N_29967,N_29602);
nand UO_733 (O_733,N_29574,N_29708);
or UO_734 (O_734,N_29626,N_29543);
nand UO_735 (O_735,N_29574,N_29796);
nand UO_736 (O_736,N_29962,N_29518);
or UO_737 (O_737,N_29600,N_29852);
nor UO_738 (O_738,N_29520,N_29852);
nor UO_739 (O_739,N_29919,N_29630);
nand UO_740 (O_740,N_29504,N_29993);
nor UO_741 (O_741,N_29735,N_29866);
nand UO_742 (O_742,N_29686,N_29821);
nor UO_743 (O_743,N_29776,N_29558);
xnor UO_744 (O_744,N_29763,N_29607);
and UO_745 (O_745,N_29746,N_29501);
xor UO_746 (O_746,N_29671,N_29932);
and UO_747 (O_747,N_29565,N_29861);
nor UO_748 (O_748,N_29980,N_29581);
or UO_749 (O_749,N_29812,N_29560);
nand UO_750 (O_750,N_29921,N_29514);
xor UO_751 (O_751,N_29591,N_29736);
nor UO_752 (O_752,N_29551,N_29586);
or UO_753 (O_753,N_29730,N_29550);
and UO_754 (O_754,N_29682,N_29658);
xnor UO_755 (O_755,N_29924,N_29583);
nor UO_756 (O_756,N_29535,N_29692);
nand UO_757 (O_757,N_29834,N_29720);
nand UO_758 (O_758,N_29581,N_29734);
or UO_759 (O_759,N_29680,N_29952);
xnor UO_760 (O_760,N_29865,N_29688);
nand UO_761 (O_761,N_29937,N_29736);
and UO_762 (O_762,N_29613,N_29704);
or UO_763 (O_763,N_29618,N_29620);
and UO_764 (O_764,N_29745,N_29523);
and UO_765 (O_765,N_29811,N_29660);
xor UO_766 (O_766,N_29541,N_29742);
nor UO_767 (O_767,N_29863,N_29931);
and UO_768 (O_768,N_29629,N_29930);
and UO_769 (O_769,N_29748,N_29540);
nand UO_770 (O_770,N_29972,N_29900);
xnor UO_771 (O_771,N_29824,N_29993);
nand UO_772 (O_772,N_29651,N_29632);
nand UO_773 (O_773,N_29758,N_29581);
and UO_774 (O_774,N_29524,N_29898);
and UO_775 (O_775,N_29612,N_29670);
xor UO_776 (O_776,N_29528,N_29788);
xnor UO_777 (O_777,N_29540,N_29698);
or UO_778 (O_778,N_29952,N_29660);
nor UO_779 (O_779,N_29964,N_29642);
and UO_780 (O_780,N_29595,N_29728);
nand UO_781 (O_781,N_29506,N_29746);
nor UO_782 (O_782,N_29993,N_29700);
nand UO_783 (O_783,N_29858,N_29948);
xor UO_784 (O_784,N_29632,N_29506);
xor UO_785 (O_785,N_29703,N_29661);
xor UO_786 (O_786,N_29983,N_29704);
nor UO_787 (O_787,N_29769,N_29529);
or UO_788 (O_788,N_29586,N_29709);
or UO_789 (O_789,N_29778,N_29895);
nand UO_790 (O_790,N_29774,N_29658);
nor UO_791 (O_791,N_29932,N_29805);
nand UO_792 (O_792,N_29805,N_29813);
xor UO_793 (O_793,N_29947,N_29687);
nand UO_794 (O_794,N_29697,N_29611);
nand UO_795 (O_795,N_29810,N_29935);
nand UO_796 (O_796,N_29529,N_29999);
nand UO_797 (O_797,N_29595,N_29544);
and UO_798 (O_798,N_29528,N_29854);
xor UO_799 (O_799,N_29746,N_29792);
and UO_800 (O_800,N_29828,N_29675);
or UO_801 (O_801,N_29829,N_29977);
or UO_802 (O_802,N_29679,N_29521);
nand UO_803 (O_803,N_29855,N_29935);
xnor UO_804 (O_804,N_29527,N_29551);
or UO_805 (O_805,N_29600,N_29516);
xor UO_806 (O_806,N_29716,N_29879);
and UO_807 (O_807,N_29878,N_29977);
xor UO_808 (O_808,N_29733,N_29967);
nand UO_809 (O_809,N_29550,N_29715);
nor UO_810 (O_810,N_29792,N_29945);
nor UO_811 (O_811,N_29948,N_29918);
xor UO_812 (O_812,N_29527,N_29932);
nand UO_813 (O_813,N_29526,N_29548);
and UO_814 (O_814,N_29793,N_29921);
or UO_815 (O_815,N_29927,N_29985);
or UO_816 (O_816,N_29933,N_29890);
nand UO_817 (O_817,N_29548,N_29722);
nor UO_818 (O_818,N_29894,N_29878);
nand UO_819 (O_819,N_29897,N_29954);
or UO_820 (O_820,N_29978,N_29575);
xnor UO_821 (O_821,N_29914,N_29594);
or UO_822 (O_822,N_29848,N_29938);
and UO_823 (O_823,N_29997,N_29670);
nor UO_824 (O_824,N_29625,N_29718);
xor UO_825 (O_825,N_29685,N_29670);
nor UO_826 (O_826,N_29613,N_29739);
and UO_827 (O_827,N_29943,N_29761);
or UO_828 (O_828,N_29902,N_29769);
xor UO_829 (O_829,N_29567,N_29739);
xor UO_830 (O_830,N_29742,N_29945);
nor UO_831 (O_831,N_29556,N_29579);
or UO_832 (O_832,N_29747,N_29889);
xnor UO_833 (O_833,N_29536,N_29528);
and UO_834 (O_834,N_29787,N_29641);
or UO_835 (O_835,N_29981,N_29819);
nor UO_836 (O_836,N_29758,N_29791);
or UO_837 (O_837,N_29618,N_29637);
xor UO_838 (O_838,N_29801,N_29794);
xnor UO_839 (O_839,N_29796,N_29907);
and UO_840 (O_840,N_29624,N_29609);
xnor UO_841 (O_841,N_29520,N_29632);
nor UO_842 (O_842,N_29915,N_29998);
or UO_843 (O_843,N_29839,N_29889);
xor UO_844 (O_844,N_29980,N_29583);
and UO_845 (O_845,N_29712,N_29700);
nor UO_846 (O_846,N_29846,N_29548);
and UO_847 (O_847,N_29912,N_29781);
nor UO_848 (O_848,N_29602,N_29514);
or UO_849 (O_849,N_29979,N_29584);
xnor UO_850 (O_850,N_29972,N_29769);
nor UO_851 (O_851,N_29887,N_29778);
nand UO_852 (O_852,N_29599,N_29715);
xor UO_853 (O_853,N_29589,N_29673);
and UO_854 (O_854,N_29714,N_29687);
xnor UO_855 (O_855,N_29939,N_29619);
nand UO_856 (O_856,N_29918,N_29814);
xnor UO_857 (O_857,N_29847,N_29620);
xnor UO_858 (O_858,N_29985,N_29881);
nand UO_859 (O_859,N_29613,N_29571);
xnor UO_860 (O_860,N_29760,N_29946);
or UO_861 (O_861,N_29894,N_29829);
nand UO_862 (O_862,N_29532,N_29782);
nor UO_863 (O_863,N_29578,N_29853);
xor UO_864 (O_864,N_29833,N_29662);
and UO_865 (O_865,N_29644,N_29592);
nand UO_866 (O_866,N_29784,N_29839);
nor UO_867 (O_867,N_29946,N_29691);
or UO_868 (O_868,N_29521,N_29966);
and UO_869 (O_869,N_29560,N_29922);
xnor UO_870 (O_870,N_29810,N_29629);
and UO_871 (O_871,N_29511,N_29603);
nor UO_872 (O_872,N_29641,N_29849);
xnor UO_873 (O_873,N_29997,N_29626);
xor UO_874 (O_874,N_29998,N_29625);
nor UO_875 (O_875,N_29820,N_29671);
nand UO_876 (O_876,N_29685,N_29755);
and UO_877 (O_877,N_29536,N_29551);
xnor UO_878 (O_878,N_29986,N_29925);
or UO_879 (O_879,N_29609,N_29679);
nand UO_880 (O_880,N_29869,N_29581);
nand UO_881 (O_881,N_29875,N_29972);
or UO_882 (O_882,N_29852,N_29726);
or UO_883 (O_883,N_29862,N_29580);
or UO_884 (O_884,N_29861,N_29803);
and UO_885 (O_885,N_29562,N_29927);
nand UO_886 (O_886,N_29666,N_29941);
xor UO_887 (O_887,N_29813,N_29725);
or UO_888 (O_888,N_29964,N_29753);
nand UO_889 (O_889,N_29719,N_29591);
or UO_890 (O_890,N_29867,N_29726);
or UO_891 (O_891,N_29964,N_29519);
nand UO_892 (O_892,N_29657,N_29721);
xnor UO_893 (O_893,N_29664,N_29706);
nand UO_894 (O_894,N_29524,N_29579);
xnor UO_895 (O_895,N_29786,N_29652);
or UO_896 (O_896,N_29918,N_29806);
nor UO_897 (O_897,N_29780,N_29726);
nor UO_898 (O_898,N_29609,N_29929);
and UO_899 (O_899,N_29705,N_29967);
nand UO_900 (O_900,N_29725,N_29598);
nor UO_901 (O_901,N_29601,N_29736);
nor UO_902 (O_902,N_29987,N_29549);
nand UO_903 (O_903,N_29566,N_29748);
and UO_904 (O_904,N_29558,N_29890);
and UO_905 (O_905,N_29975,N_29922);
nand UO_906 (O_906,N_29653,N_29783);
xnor UO_907 (O_907,N_29566,N_29618);
nor UO_908 (O_908,N_29598,N_29521);
or UO_909 (O_909,N_29605,N_29572);
or UO_910 (O_910,N_29825,N_29549);
or UO_911 (O_911,N_29962,N_29897);
nand UO_912 (O_912,N_29568,N_29585);
or UO_913 (O_913,N_29540,N_29824);
and UO_914 (O_914,N_29889,N_29934);
nor UO_915 (O_915,N_29851,N_29674);
or UO_916 (O_916,N_29637,N_29651);
xnor UO_917 (O_917,N_29665,N_29993);
or UO_918 (O_918,N_29501,N_29717);
and UO_919 (O_919,N_29623,N_29596);
nor UO_920 (O_920,N_29974,N_29977);
nand UO_921 (O_921,N_29935,N_29952);
nand UO_922 (O_922,N_29988,N_29940);
nor UO_923 (O_923,N_29886,N_29952);
or UO_924 (O_924,N_29877,N_29902);
nor UO_925 (O_925,N_29975,N_29996);
xor UO_926 (O_926,N_29692,N_29785);
nand UO_927 (O_927,N_29944,N_29814);
or UO_928 (O_928,N_29670,N_29875);
nand UO_929 (O_929,N_29520,N_29890);
and UO_930 (O_930,N_29915,N_29683);
or UO_931 (O_931,N_29615,N_29676);
or UO_932 (O_932,N_29682,N_29930);
nor UO_933 (O_933,N_29886,N_29778);
nand UO_934 (O_934,N_29593,N_29971);
nor UO_935 (O_935,N_29704,N_29853);
xnor UO_936 (O_936,N_29773,N_29982);
nor UO_937 (O_937,N_29613,N_29649);
and UO_938 (O_938,N_29576,N_29595);
nand UO_939 (O_939,N_29576,N_29996);
nand UO_940 (O_940,N_29956,N_29697);
and UO_941 (O_941,N_29593,N_29929);
or UO_942 (O_942,N_29832,N_29857);
xnor UO_943 (O_943,N_29985,N_29600);
nand UO_944 (O_944,N_29593,N_29573);
xnor UO_945 (O_945,N_29802,N_29994);
xor UO_946 (O_946,N_29683,N_29933);
xnor UO_947 (O_947,N_29540,N_29589);
and UO_948 (O_948,N_29600,N_29707);
nand UO_949 (O_949,N_29917,N_29578);
nor UO_950 (O_950,N_29941,N_29928);
nor UO_951 (O_951,N_29847,N_29751);
nand UO_952 (O_952,N_29713,N_29965);
and UO_953 (O_953,N_29713,N_29754);
and UO_954 (O_954,N_29991,N_29651);
xor UO_955 (O_955,N_29529,N_29770);
or UO_956 (O_956,N_29916,N_29987);
nand UO_957 (O_957,N_29821,N_29623);
nor UO_958 (O_958,N_29590,N_29670);
nand UO_959 (O_959,N_29607,N_29856);
xor UO_960 (O_960,N_29679,N_29802);
xor UO_961 (O_961,N_29683,N_29744);
nor UO_962 (O_962,N_29616,N_29836);
and UO_963 (O_963,N_29556,N_29847);
nor UO_964 (O_964,N_29558,N_29806);
nand UO_965 (O_965,N_29983,N_29680);
nand UO_966 (O_966,N_29667,N_29878);
nand UO_967 (O_967,N_29894,N_29590);
xor UO_968 (O_968,N_29910,N_29985);
nand UO_969 (O_969,N_29593,N_29746);
and UO_970 (O_970,N_29704,N_29751);
and UO_971 (O_971,N_29812,N_29820);
nand UO_972 (O_972,N_29998,N_29910);
or UO_973 (O_973,N_29854,N_29759);
and UO_974 (O_974,N_29757,N_29602);
or UO_975 (O_975,N_29790,N_29855);
nor UO_976 (O_976,N_29711,N_29664);
and UO_977 (O_977,N_29733,N_29553);
or UO_978 (O_978,N_29885,N_29948);
nor UO_979 (O_979,N_29891,N_29681);
or UO_980 (O_980,N_29753,N_29631);
or UO_981 (O_981,N_29753,N_29954);
nor UO_982 (O_982,N_29599,N_29678);
nand UO_983 (O_983,N_29715,N_29695);
nand UO_984 (O_984,N_29705,N_29948);
xor UO_985 (O_985,N_29507,N_29697);
xor UO_986 (O_986,N_29939,N_29936);
or UO_987 (O_987,N_29920,N_29597);
xor UO_988 (O_988,N_29842,N_29615);
nand UO_989 (O_989,N_29980,N_29719);
nand UO_990 (O_990,N_29577,N_29668);
nand UO_991 (O_991,N_29704,N_29975);
xnor UO_992 (O_992,N_29525,N_29828);
nor UO_993 (O_993,N_29708,N_29500);
or UO_994 (O_994,N_29952,N_29668);
nand UO_995 (O_995,N_29724,N_29878);
nand UO_996 (O_996,N_29867,N_29542);
or UO_997 (O_997,N_29693,N_29563);
nand UO_998 (O_998,N_29511,N_29716);
xor UO_999 (O_999,N_29593,N_29764);
nor UO_1000 (O_1000,N_29668,N_29839);
nor UO_1001 (O_1001,N_29687,N_29567);
nor UO_1002 (O_1002,N_29890,N_29812);
or UO_1003 (O_1003,N_29609,N_29513);
nand UO_1004 (O_1004,N_29836,N_29653);
xnor UO_1005 (O_1005,N_29994,N_29854);
xor UO_1006 (O_1006,N_29949,N_29624);
and UO_1007 (O_1007,N_29988,N_29633);
nor UO_1008 (O_1008,N_29757,N_29517);
xnor UO_1009 (O_1009,N_29521,N_29719);
and UO_1010 (O_1010,N_29516,N_29886);
nand UO_1011 (O_1011,N_29553,N_29918);
nor UO_1012 (O_1012,N_29897,N_29836);
nor UO_1013 (O_1013,N_29610,N_29948);
nor UO_1014 (O_1014,N_29546,N_29757);
and UO_1015 (O_1015,N_29912,N_29732);
xor UO_1016 (O_1016,N_29765,N_29744);
nand UO_1017 (O_1017,N_29988,N_29806);
xor UO_1018 (O_1018,N_29550,N_29795);
or UO_1019 (O_1019,N_29625,N_29643);
and UO_1020 (O_1020,N_29924,N_29986);
nor UO_1021 (O_1021,N_29858,N_29562);
or UO_1022 (O_1022,N_29763,N_29702);
nor UO_1023 (O_1023,N_29963,N_29973);
xnor UO_1024 (O_1024,N_29971,N_29961);
and UO_1025 (O_1025,N_29832,N_29736);
nor UO_1026 (O_1026,N_29576,N_29665);
or UO_1027 (O_1027,N_29591,N_29621);
nand UO_1028 (O_1028,N_29520,N_29779);
nand UO_1029 (O_1029,N_29954,N_29811);
and UO_1030 (O_1030,N_29968,N_29692);
xor UO_1031 (O_1031,N_29786,N_29851);
xnor UO_1032 (O_1032,N_29979,N_29619);
xor UO_1033 (O_1033,N_29816,N_29651);
nor UO_1034 (O_1034,N_29617,N_29937);
or UO_1035 (O_1035,N_29886,N_29709);
xor UO_1036 (O_1036,N_29510,N_29930);
and UO_1037 (O_1037,N_29513,N_29619);
xor UO_1038 (O_1038,N_29552,N_29769);
nor UO_1039 (O_1039,N_29961,N_29692);
and UO_1040 (O_1040,N_29973,N_29874);
and UO_1041 (O_1041,N_29641,N_29892);
or UO_1042 (O_1042,N_29763,N_29826);
and UO_1043 (O_1043,N_29762,N_29842);
nand UO_1044 (O_1044,N_29702,N_29817);
or UO_1045 (O_1045,N_29944,N_29599);
xnor UO_1046 (O_1046,N_29539,N_29629);
nand UO_1047 (O_1047,N_29602,N_29788);
or UO_1048 (O_1048,N_29999,N_29873);
xor UO_1049 (O_1049,N_29716,N_29960);
and UO_1050 (O_1050,N_29578,N_29751);
and UO_1051 (O_1051,N_29517,N_29660);
nand UO_1052 (O_1052,N_29515,N_29966);
and UO_1053 (O_1053,N_29855,N_29607);
xnor UO_1054 (O_1054,N_29884,N_29644);
or UO_1055 (O_1055,N_29938,N_29924);
xor UO_1056 (O_1056,N_29507,N_29752);
nor UO_1057 (O_1057,N_29862,N_29581);
and UO_1058 (O_1058,N_29884,N_29557);
xor UO_1059 (O_1059,N_29671,N_29957);
xnor UO_1060 (O_1060,N_29757,N_29983);
or UO_1061 (O_1061,N_29590,N_29887);
and UO_1062 (O_1062,N_29832,N_29920);
xor UO_1063 (O_1063,N_29582,N_29656);
nor UO_1064 (O_1064,N_29600,N_29614);
or UO_1065 (O_1065,N_29890,N_29631);
nor UO_1066 (O_1066,N_29687,N_29950);
nand UO_1067 (O_1067,N_29969,N_29783);
nand UO_1068 (O_1068,N_29541,N_29703);
xor UO_1069 (O_1069,N_29574,N_29570);
xnor UO_1070 (O_1070,N_29794,N_29861);
nand UO_1071 (O_1071,N_29837,N_29755);
and UO_1072 (O_1072,N_29532,N_29734);
and UO_1073 (O_1073,N_29824,N_29602);
and UO_1074 (O_1074,N_29853,N_29802);
and UO_1075 (O_1075,N_29514,N_29563);
nor UO_1076 (O_1076,N_29537,N_29924);
xor UO_1077 (O_1077,N_29688,N_29972);
xor UO_1078 (O_1078,N_29686,N_29655);
nand UO_1079 (O_1079,N_29600,N_29929);
nand UO_1080 (O_1080,N_29889,N_29544);
nor UO_1081 (O_1081,N_29521,N_29531);
xnor UO_1082 (O_1082,N_29636,N_29573);
or UO_1083 (O_1083,N_29812,N_29874);
nor UO_1084 (O_1084,N_29879,N_29712);
or UO_1085 (O_1085,N_29781,N_29648);
nand UO_1086 (O_1086,N_29685,N_29608);
nor UO_1087 (O_1087,N_29639,N_29980);
nand UO_1088 (O_1088,N_29956,N_29547);
nand UO_1089 (O_1089,N_29574,N_29715);
or UO_1090 (O_1090,N_29532,N_29825);
xor UO_1091 (O_1091,N_29754,N_29818);
and UO_1092 (O_1092,N_29644,N_29776);
nor UO_1093 (O_1093,N_29525,N_29744);
or UO_1094 (O_1094,N_29813,N_29966);
nor UO_1095 (O_1095,N_29514,N_29889);
xnor UO_1096 (O_1096,N_29665,N_29640);
xnor UO_1097 (O_1097,N_29696,N_29782);
or UO_1098 (O_1098,N_29878,N_29829);
or UO_1099 (O_1099,N_29999,N_29978);
and UO_1100 (O_1100,N_29976,N_29806);
or UO_1101 (O_1101,N_29725,N_29766);
xnor UO_1102 (O_1102,N_29558,N_29824);
and UO_1103 (O_1103,N_29953,N_29984);
xnor UO_1104 (O_1104,N_29931,N_29928);
nand UO_1105 (O_1105,N_29899,N_29944);
xnor UO_1106 (O_1106,N_29729,N_29763);
and UO_1107 (O_1107,N_29569,N_29961);
xor UO_1108 (O_1108,N_29907,N_29914);
xnor UO_1109 (O_1109,N_29875,N_29678);
xor UO_1110 (O_1110,N_29849,N_29891);
nor UO_1111 (O_1111,N_29776,N_29774);
nand UO_1112 (O_1112,N_29972,N_29684);
nand UO_1113 (O_1113,N_29673,N_29553);
xor UO_1114 (O_1114,N_29696,N_29595);
nand UO_1115 (O_1115,N_29554,N_29571);
nor UO_1116 (O_1116,N_29639,N_29806);
nor UO_1117 (O_1117,N_29504,N_29714);
nand UO_1118 (O_1118,N_29716,N_29655);
and UO_1119 (O_1119,N_29757,N_29866);
xor UO_1120 (O_1120,N_29563,N_29616);
or UO_1121 (O_1121,N_29516,N_29723);
xnor UO_1122 (O_1122,N_29997,N_29815);
nand UO_1123 (O_1123,N_29879,N_29885);
xor UO_1124 (O_1124,N_29805,N_29627);
xor UO_1125 (O_1125,N_29709,N_29735);
nor UO_1126 (O_1126,N_29605,N_29690);
or UO_1127 (O_1127,N_29688,N_29870);
and UO_1128 (O_1128,N_29860,N_29537);
nor UO_1129 (O_1129,N_29913,N_29586);
xor UO_1130 (O_1130,N_29563,N_29900);
and UO_1131 (O_1131,N_29828,N_29610);
xor UO_1132 (O_1132,N_29801,N_29841);
nor UO_1133 (O_1133,N_29850,N_29549);
nor UO_1134 (O_1134,N_29812,N_29919);
nor UO_1135 (O_1135,N_29731,N_29535);
and UO_1136 (O_1136,N_29768,N_29732);
xor UO_1137 (O_1137,N_29981,N_29552);
nand UO_1138 (O_1138,N_29669,N_29688);
and UO_1139 (O_1139,N_29715,N_29725);
or UO_1140 (O_1140,N_29723,N_29540);
xnor UO_1141 (O_1141,N_29761,N_29788);
nand UO_1142 (O_1142,N_29746,N_29788);
nor UO_1143 (O_1143,N_29504,N_29755);
or UO_1144 (O_1144,N_29849,N_29898);
xnor UO_1145 (O_1145,N_29743,N_29858);
and UO_1146 (O_1146,N_29773,N_29888);
nor UO_1147 (O_1147,N_29517,N_29537);
nand UO_1148 (O_1148,N_29946,N_29950);
xnor UO_1149 (O_1149,N_29798,N_29530);
and UO_1150 (O_1150,N_29829,N_29732);
nand UO_1151 (O_1151,N_29640,N_29834);
or UO_1152 (O_1152,N_29764,N_29823);
nor UO_1153 (O_1153,N_29857,N_29813);
and UO_1154 (O_1154,N_29836,N_29955);
xnor UO_1155 (O_1155,N_29717,N_29545);
xnor UO_1156 (O_1156,N_29691,N_29880);
and UO_1157 (O_1157,N_29628,N_29742);
nand UO_1158 (O_1158,N_29667,N_29703);
or UO_1159 (O_1159,N_29622,N_29609);
nor UO_1160 (O_1160,N_29555,N_29869);
or UO_1161 (O_1161,N_29992,N_29674);
and UO_1162 (O_1162,N_29563,N_29691);
or UO_1163 (O_1163,N_29621,N_29695);
or UO_1164 (O_1164,N_29594,N_29738);
nand UO_1165 (O_1165,N_29696,N_29599);
or UO_1166 (O_1166,N_29762,N_29834);
or UO_1167 (O_1167,N_29722,N_29824);
xnor UO_1168 (O_1168,N_29980,N_29654);
and UO_1169 (O_1169,N_29691,N_29647);
and UO_1170 (O_1170,N_29754,N_29542);
nor UO_1171 (O_1171,N_29537,N_29908);
nor UO_1172 (O_1172,N_29884,N_29953);
nand UO_1173 (O_1173,N_29929,N_29967);
and UO_1174 (O_1174,N_29640,N_29839);
xnor UO_1175 (O_1175,N_29744,N_29672);
xnor UO_1176 (O_1176,N_29920,N_29676);
nor UO_1177 (O_1177,N_29778,N_29647);
nand UO_1178 (O_1178,N_29663,N_29533);
or UO_1179 (O_1179,N_29565,N_29866);
and UO_1180 (O_1180,N_29782,N_29590);
xnor UO_1181 (O_1181,N_29765,N_29809);
nand UO_1182 (O_1182,N_29543,N_29822);
xnor UO_1183 (O_1183,N_29866,N_29589);
and UO_1184 (O_1184,N_29846,N_29570);
nand UO_1185 (O_1185,N_29556,N_29587);
nand UO_1186 (O_1186,N_29774,N_29963);
or UO_1187 (O_1187,N_29870,N_29593);
and UO_1188 (O_1188,N_29603,N_29503);
and UO_1189 (O_1189,N_29549,N_29578);
xnor UO_1190 (O_1190,N_29563,N_29821);
nor UO_1191 (O_1191,N_29795,N_29615);
nor UO_1192 (O_1192,N_29885,N_29524);
and UO_1193 (O_1193,N_29682,N_29607);
xnor UO_1194 (O_1194,N_29714,N_29999);
xor UO_1195 (O_1195,N_29606,N_29977);
and UO_1196 (O_1196,N_29590,N_29634);
xnor UO_1197 (O_1197,N_29509,N_29599);
nand UO_1198 (O_1198,N_29731,N_29740);
xor UO_1199 (O_1199,N_29565,N_29849);
or UO_1200 (O_1200,N_29837,N_29517);
xor UO_1201 (O_1201,N_29627,N_29991);
xnor UO_1202 (O_1202,N_29547,N_29530);
and UO_1203 (O_1203,N_29995,N_29580);
xor UO_1204 (O_1204,N_29943,N_29967);
xnor UO_1205 (O_1205,N_29621,N_29875);
xnor UO_1206 (O_1206,N_29944,N_29551);
and UO_1207 (O_1207,N_29701,N_29739);
or UO_1208 (O_1208,N_29667,N_29730);
and UO_1209 (O_1209,N_29614,N_29748);
nor UO_1210 (O_1210,N_29535,N_29732);
and UO_1211 (O_1211,N_29509,N_29803);
nand UO_1212 (O_1212,N_29891,N_29569);
and UO_1213 (O_1213,N_29680,N_29985);
nor UO_1214 (O_1214,N_29662,N_29813);
and UO_1215 (O_1215,N_29729,N_29775);
and UO_1216 (O_1216,N_29923,N_29579);
and UO_1217 (O_1217,N_29899,N_29880);
xor UO_1218 (O_1218,N_29745,N_29730);
xnor UO_1219 (O_1219,N_29807,N_29550);
xor UO_1220 (O_1220,N_29966,N_29987);
or UO_1221 (O_1221,N_29646,N_29658);
nor UO_1222 (O_1222,N_29807,N_29932);
and UO_1223 (O_1223,N_29942,N_29642);
or UO_1224 (O_1224,N_29544,N_29763);
or UO_1225 (O_1225,N_29942,N_29834);
and UO_1226 (O_1226,N_29505,N_29696);
or UO_1227 (O_1227,N_29909,N_29989);
or UO_1228 (O_1228,N_29754,N_29533);
or UO_1229 (O_1229,N_29699,N_29848);
nor UO_1230 (O_1230,N_29797,N_29915);
nand UO_1231 (O_1231,N_29559,N_29933);
and UO_1232 (O_1232,N_29665,N_29926);
nor UO_1233 (O_1233,N_29882,N_29911);
xor UO_1234 (O_1234,N_29784,N_29516);
or UO_1235 (O_1235,N_29811,N_29593);
nand UO_1236 (O_1236,N_29973,N_29837);
and UO_1237 (O_1237,N_29655,N_29781);
nor UO_1238 (O_1238,N_29980,N_29548);
and UO_1239 (O_1239,N_29694,N_29944);
or UO_1240 (O_1240,N_29901,N_29657);
xnor UO_1241 (O_1241,N_29527,N_29903);
or UO_1242 (O_1242,N_29879,N_29516);
and UO_1243 (O_1243,N_29882,N_29682);
nor UO_1244 (O_1244,N_29731,N_29914);
xnor UO_1245 (O_1245,N_29787,N_29926);
nor UO_1246 (O_1246,N_29742,N_29748);
or UO_1247 (O_1247,N_29772,N_29980);
xor UO_1248 (O_1248,N_29980,N_29536);
xnor UO_1249 (O_1249,N_29616,N_29818);
nand UO_1250 (O_1250,N_29706,N_29871);
or UO_1251 (O_1251,N_29650,N_29798);
and UO_1252 (O_1252,N_29952,N_29725);
nand UO_1253 (O_1253,N_29642,N_29855);
xnor UO_1254 (O_1254,N_29733,N_29530);
nand UO_1255 (O_1255,N_29637,N_29579);
xnor UO_1256 (O_1256,N_29879,N_29624);
xnor UO_1257 (O_1257,N_29656,N_29774);
or UO_1258 (O_1258,N_29779,N_29595);
and UO_1259 (O_1259,N_29657,N_29999);
xnor UO_1260 (O_1260,N_29955,N_29885);
nor UO_1261 (O_1261,N_29951,N_29990);
or UO_1262 (O_1262,N_29627,N_29517);
nor UO_1263 (O_1263,N_29598,N_29657);
xnor UO_1264 (O_1264,N_29756,N_29852);
and UO_1265 (O_1265,N_29887,N_29507);
or UO_1266 (O_1266,N_29963,N_29552);
and UO_1267 (O_1267,N_29790,N_29803);
xnor UO_1268 (O_1268,N_29979,N_29634);
nand UO_1269 (O_1269,N_29705,N_29696);
or UO_1270 (O_1270,N_29919,N_29751);
xnor UO_1271 (O_1271,N_29770,N_29817);
nand UO_1272 (O_1272,N_29874,N_29981);
or UO_1273 (O_1273,N_29885,N_29818);
nor UO_1274 (O_1274,N_29531,N_29787);
or UO_1275 (O_1275,N_29955,N_29586);
nand UO_1276 (O_1276,N_29523,N_29851);
nor UO_1277 (O_1277,N_29889,N_29875);
nand UO_1278 (O_1278,N_29677,N_29642);
nand UO_1279 (O_1279,N_29602,N_29530);
or UO_1280 (O_1280,N_29902,N_29517);
xor UO_1281 (O_1281,N_29696,N_29896);
and UO_1282 (O_1282,N_29996,N_29570);
or UO_1283 (O_1283,N_29909,N_29895);
nand UO_1284 (O_1284,N_29664,N_29895);
or UO_1285 (O_1285,N_29562,N_29924);
nor UO_1286 (O_1286,N_29960,N_29686);
and UO_1287 (O_1287,N_29631,N_29614);
and UO_1288 (O_1288,N_29806,N_29933);
xor UO_1289 (O_1289,N_29547,N_29912);
or UO_1290 (O_1290,N_29991,N_29727);
or UO_1291 (O_1291,N_29947,N_29728);
or UO_1292 (O_1292,N_29597,N_29534);
and UO_1293 (O_1293,N_29740,N_29778);
or UO_1294 (O_1294,N_29882,N_29647);
or UO_1295 (O_1295,N_29638,N_29949);
xnor UO_1296 (O_1296,N_29860,N_29788);
xor UO_1297 (O_1297,N_29711,N_29961);
and UO_1298 (O_1298,N_29834,N_29653);
and UO_1299 (O_1299,N_29872,N_29761);
nand UO_1300 (O_1300,N_29843,N_29535);
or UO_1301 (O_1301,N_29708,N_29634);
xor UO_1302 (O_1302,N_29832,N_29883);
nand UO_1303 (O_1303,N_29596,N_29632);
or UO_1304 (O_1304,N_29535,N_29831);
and UO_1305 (O_1305,N_29920,N_29547);
and UO_1306 (O_1306,N_29696,N_29706);
nor UO_1307 (O_1307,N_29790,N_29757);
or UO_1308 (O_1308,N_29585,N_29573);
nor UO_1309 (O_1309,N_29537,N_29890);
nand UO_1310 (O_1310,N_29535,N_29869);
nor UO_1311 (O_1311,N_29643,N_29912);
and UO_1312 (O_1312,N_29593,N_29950);
and UO_1313 (O_1313,N_29547,N_29736);
and UO_1314 (O_1314,N_29686,N_29818);
nand UO_1315 (O_1315,N_29721,N_29606);
and UO_1316 (O_1316,N_29941,N_29522);
nor UO_1317 (O_1317,N_29989,N_29927);
xor UO_1318 (O_1318,N_29936,N_29852);
nand UO_1319 (O_1319,N_29696,N_29707);
and UO_1320 (O_1320,N_29752,N_29894);
or UO_1321 (O_1321,N_29577,N_29992);
or UO_1322 (O_1322,N_29516,N_29685);
nor UO_1323 (O_1323,N_29591,N_29559);
xor UO_1324 (O_1324,N_29836,N_29610);
nor UO_1325 (O_1325,N_29877,N_29853);
nand UO_1326 (O_1326,N_29894,N_29665);
xor UO_1327 (O_1327,N_29873,N_29938);
and UO_1328 (O_1328,N_29772,N_29729);
and UO_1329 (O_1329,N_29792,N_29978);
nor UO_1330 (O_1330,N_29644,N_29979);
nor UO_1331 (O_1331,N_29641,N_29778);
xnor UO_1332 (O_1332,N_29613,N_29714);
or UO_1333 (O_1333,N_29520,N_29826);
and UO_1334 (O_1334,N_29598,N_29936);
nor UO_1335 (O_1335,N_29503,N_29812);
and UO_1336 (O_1336,N_29831,N_29715);
or UO_1337 (O_1337,N_29832,N_29992);
nand UO_1338 (O_1338,N_29859,N_29652);
or UO_1339 (O_1339,N_29908,N_29730);
or UO_1340 (O_1340,N_29801,N_29653);
or UO_1341 (O_1341,N_29691,N_29657);
and UO_1342 (O_1342,N_29879,N_29749);
nand UO_1343 (O_1343,N_29787,N_29789);
xnor UO_1344 (O_1344,N_29538,N_29944);
xor UO_1345 (O_1345,N_29984,N_29773);
nand UO_1346 (O_1346,N_29587,N_29628);
and UO_1347 (O_1347,N_29580,N_29871);
nand UO_1348 (O_1348,N_29633,N_29972);
xnor UO_1349 (O_1349,N_29845,N_29766);
or UO_1350 (O_1350,N_29856,N_29825);
and UO_1351 (O_1351,N_29659,N_29731);
xnor UO_1352 (O_1352,N_29932,N_29739);
nand UO_1353 (O_1353,N_29524,N_29735);
xnor UO_1354 (O_1354,N_29835,N_29963);
nand UO_1355 (O_1355,N_29575,N_29660);
xnor UO_1356 (O_1356,N_29619,N_29707);
nand UO_1357 (O_1357,N_29563,N_29739);
nor UO_1358 (O_1358,N_29675,N_29950);
nor UO_1359 (O_1359,N_29804,N_29598);
or UO_1360 (O_1360,N_29547,N_29584);
or UO_1361 (O_1361,N_29907,N_29791);
nand UO_1362 (O_1362,N_29761,N_29531);
and UO_1363 (O_1363,N_29915,N_29888);
nor UO_1364 (O_1364,N_29773,N_29562);
and UO_1365 (O_1365,N_29694,N_29914);
xnor UO_1366 (O_1366,N_29883,N_29785);
nor UO_1367 (O_1367,N_29739,N_29561);
or UO_1368 (O_1368,N_29861,N_29759);
and UO_1369 (O_1369,N_29729,N_29986);
xor UO_1370 (O_1370,N_29582,N_29806);
nand UO_1371 (O_1371,N_29544,N_29836);
and UO_1372 (O_1372,N_29695,N_29750);
or UO_1373 (O_1373,N_29636,N_29835);
nor UO_1374 (O_1374,N_29875,N_29636);
nor UO_1375 (O_1375,N_29899,N_29600);
nand UO_1376 (O_1376,N_29811,N_29903);
nand UO_1377 (O_1377,N_29753,N_29819);
or UO_1378 (O_1378,N_29835,N_29943);
nor UO_1379 (O_1379,N_29821,N_29518);
xnor UO_1380 (O_1380,N_29893,N_29872);
and UO_1381 (O_1381,N_29786,N_29519);
xnor UO_1382 (O_1382,N_29693,N_29902);
xnor UO_1383 (O_1383,N_29639,N_29995);
or UO_1384 (O_1384,N_29810,N_29865);
nand UO_1385 (O_1385,N_29933,N_29957);
nand UO_1386 (O_1386,N_29758,N_29775);
nand UO_1387 (O_1387,N_29935,N_29638);
and UO_1388 (O_1388,N_29803,N_29852);
or UO_1389 (O_1389,N_29762,N_29881);
nand UO_1390 (O_1390,N_29501,N_29623);
xnor UO_1391 (O_1391,N_29723,N_29952);
or UO_1392 (O_1392,N_29970,N_29624);
nor UO_1393 (O_1393,N_29669,N_29744);
and UO_1394 (O_1394,N_29839,N_29521);
and UO_1395 (O_1395,N_29975,N_29563);
nand UO_1396 (O_1396,N_29563,N_29832);
nor UO_1397 (O_1397,N_29676,N_29927);
or UO_1398 (O_1398,N_29651,N_29621);
nand UO_1399 (O_1399,N_29746,N_29969);
nand UO_1400 (O_1400,N_29590,N_29772);
nand UO_1401 (O_1401,N_29805,N_29735);
nor UO_1402 (O_1402,N_29974,N_29702);
xor UO_1403 (O_1403,N_29730,N_29964);
and UO_1404 (O_1404,N_29980,N_29786);
or UO_1405 (O_1405,N_29572,N_29868);
and UO_1406 (O_1406,N_29525,N_29965);
or UO_1407 (O_1407,N_29893,N_29524);
xnor UO_1408 (O_1408,N_29926,N_29714);
and UO_1409 (O_1409,N_29692,N_29715);
nand UO_1410 (O_1410,N_29807,N_29824);
and UO_1411 (O_1411,N_29673,N_29892);
and UO_1412 (O_1412,N_29896,N_29641);
and UO_1413 (O_1413,N_29887,N_29571);
nor UO_1414 (O_1414,N_29912,N_29545);
nand UO_1415 (O_1415,N_29866,N_29750);
xor UO_1416 (O_1416,N_29670,N_29825);
and UO_1417 (O_1417,N_29710,N_29772);
xnor UO_1418 (O_1418,N_29967,N_29891);
nand UO_1419 (O_1419,N_29879,N_29619);
and UO_1420 (O_1420,N_29943,N_29872);
nand UO_1421 (O_1421,N_29885,N_29639);
nand UO_1422 (O_1422,N_29956,N_29962);
and UO_1423 (O_1423,N_29571,N_29992);
nor UO_1424 (O_1424,N_29993,N_29885);
nor UO_1425 (O_1425,N_29835,N_29939);
nand UO_1426 (O_1426,N_29967,N_29725);
or UO_1427 (O_1427,N_29511,N_29780);
or UO_1428 (O_1428,N_29881,N_29543);
xnor UO_1429 (O_1429,N_29664,N_29645);
or UO_1430 (O_1430,N_29630,N_29865);
nor UO_1431 (O_1431,N_29915,N_29552);
nor UO_1432 (O_1432,N_29549,N_29792);
or UO_1433 (O_1433,N_29701,N_29860);
nand UO_1434 (O_1434,N_29872,N_29635);
xnor UO_1435 (O_1435,N_29531,N_29509);
nor UO_1436 (O_1436,N_29912,N_29852);
nor UO_1437 (O_1437,N_29726,N_29568);
and UO_1438 (O_1438,N_29825,N_29643);
xor UO_1439 (O_1439,N_29629,N_29741);
nand UO_1440 (O_1440,N_29620,N_29664);
or UO_1441 (O_1441,N_29903,N_29882);
nor UO_1442 (O_1442,N_29660,N_29591);
nand UO_1443 (O_1443,N_29579,N_29508);
xor UO_1444 (O_1444,N_29610,N_29947);
and UO_1445 (O_1445,N_29523,N_29583);
nand UO_1446 (O_1446,N_29902,N_29534);
nor UO_1447 (O_1447,N_29742,N_29640);
nand UO_1448 (O_1448,N_29685,N_29915);
nor UO_1449 (O_1449,N_29918,N_29914);
xnor UO_1450 (O_1450,N_29512,N_29607);
nor UO_1451 (O_1451,N_29923,N_29805);
nor UO_1452 (O_1452,N_29625,N_29839);
xor UO_1453 (O_1453,N_29828,N_29561);
xnor UO_1454 (O_1454,N_29830,N_29711);
or UO_1455 (O_1455,N_29649,N_29880);
xor UO_1456 (O_1456,N_29818,N_29762);
nand UO_1457 (O_1457,N_29878,N_29712);
and UO_1458 (O_1458,N_29946,N_29558);
nand UO_1459 (O_1459,N_29530,N_29557);
nor UO_1460 (O_1460,N_29631,N_29685);
or UO_1461 (O_1461,N_29512,N_29565);
and UO_1462 (O_1462,N_29983,N_29875);
and UO_1463 (O_1463,N_29777,N_29675);
nor UO_1464 (O_1464,N_29938,N_29944);
and UO_1465 (O_1465,N_29605,N_29956);
and UO_1466 (O_1466,N_29897,N_29638);
and UO_1467 (O_1467,N_29888,N_29605);
nor UO_1468 (O_1468,N_29571,N_29544);
nand UO_1469 (O_1469,N_29870,N_29632);
and UO_1470 (O_1470,N_29518,N_29571);
xor UO_1471 (O_1471,N_29873,N_29758);
nor UO_1472 (O_1472,N_29758,N_29589);
or UO_1473 (O_1473,N_29552,N_29930);
nand UO_1474 (O_1474,N_29545,N_29629);
and UO_1475 (O_1475,N_29816,N_29599);
and UO_1476 (O_1476,N_29849,N_29862);
and UO_1477 (O_1477,N_29786,N_29753);
or UO_1478 (O_1478,N_29575,N_29560);
or UO_1479 (O_1479,N_29794,N_29559);
and UO_1480 (O_1480,N_29505,N_29748);
and UO_1481 (O_1481,N_29636,N_29532);
and UO_1482 (O_1482,N_29714,N_29763);
nand UO_1483 (O_1483,N_29643,N_29561);
and UO_1484 (O_1484,N_29995,N_29594);
and UO_1485 (O_1485,N_29824,N_29821);
nor UO_1486 (O_1486,N_29644,N_29848);
xor UO_1487 (O_1487,N_29616,N_29644);
nand UO_1488 (O_1488,N_29605,N_29529);
or UO_1489 (O_1489,N_29617,N_29712);
or UO_1490 (O_1490,N_29551,N_29992);
xor UO_1491 (O_1491,N_29628,N_29760);
and UO_1492 (O_1492,N_29598,N_29558);
and UO_1493 (O_1493,N_29679,N_29674);
or UO_1494 (O_1494,N_29820,N_29976);
and UO_1495 (O_1495,N_29634,N_29978);
and UO_1496 (O_1496,N_29897,N_29888);
nand UO_1497 (O_1497,N_29789,N_29597);
and UO_1498 (O_1498,N_29996,N_29696);
xnor UO_1499 (O_1499,N_29937,N_29946);
or UO_1500 (O_1500,N_29743,N_29541);
and UO_1501 (O_1501,N_29736,N_29986);
xnor UO_1502 (O_1502,N_29533,N_29511);
or UO_1503 (O_1503,N_29545,N_29989);
or UO_1504 (O_1504,N_29942,N_29770);
nor UO_1505 (O_1505,N_29768,N_29934);
nand UO_1506 (O_1506,N_29693,N_29509);
and UO_1507 (O_1507,N_29766,N_29746);
nor UO_1508 (O_1508,N_29746,N_29537);
nor UO_1509 (O_1509,N_29733,N_29584);
xnor UO_1510 (O_1510,N_29800,N_29719);
or UO_1511 (O_1511,N_29694,N_29751);
xnor UO_1512 (O_1512,N_29897,N_29931);
and UO_1513 (O_1513,N_29595,N_29963);
or UO_1514 (O_1514,N_29986,N_29666);
or UO_1515 (O_1515,N_29825,N_29978);
nor UO_1516 (O_1516,N_29627,N_29607);
and UO_1517 (O_1517,N_29546,N_29782);
nand UO_1518 (O_1518,N_29758,N_29949);
and UO_1519 (O_1519,N_29553,N_29902);
xnor UO_1520 (O_1520,N_29529,N_29984);
xnor UO_1521 (O_1521,N_29594,N_29814);
xor UO_1522 (O_1522,N_29714,N_29846);
or UO_1523 (O_1523,N_29956,N_29764);
xnor UO_1524 (O_1524,N_29655,N_29668);
and UO_1525 (O_1525,N_29537,N_29715);
nand UO_1526 (O_1526,N_29911,N_29603);
nor UO_1527 (O_1527,N_29703,N_29569);
nand UO_1528 (O_1528,N_29625,N_29620);
nand UO_1529 (O_1529,N_29628,N_29540);
and UO_1530 (O_1530,N_29834,N_29965);
and UO_1531 (O_1531,N_29911,N_29877);
xnor UO_1532 (O_1532,N_29581,N_29733);
nor UO_1533 (O_1533,N_29733,N_29835);
xnor UO_1534 (O_1534,N_29968,N_29961);
and UO_1535 (O_1535,N_29765,N_29570);
or UO_1536 (O_1536,N_29533,N_29698);
and UO_1537 (O_1537,N_29547,N_29911);
and UO_1538 (O_1538,N_29988,N_29963);
or UO_1539 (O_1539,N_29626,N_29631);
nand UO_1540 (O_1540,N_29726,N_29829);
nand UO_1541 (O_1541,N_29711,N_29877);
or UO_1542 (O_1542,N_29981,N_29641);
nand UO_1543 (O_1543,N_29563,N_29998);
xnor UO_1544 (O_1544,N_29539,N_29506);
xnor UO_1545 (O_1545,N_29684,N_29990);
nor UO_1546 (O_1546,N_29794,N_29931);
nor UO_1547 (O_1547,N_29651,N_29780);
or UO_1548 (O_1548,N_29919,N_29931);
xnor UO_1549 (O_1549,N_29836,N_29841);
or UO_1550 (O_1550,N_29998,N_29786);
nand UO_1551 (O_1551,N_29752,N_29978);
and UO_1552 (O_1552,N_29786,N_29971);
and UO_1553 (O_1553,N_29960,N_29573);
nand UO_1554 (O_1554,N_29569,N_29816);
xnor UO_1555 (O_1555,N_29673,N_29672);
nor UO_1556 (O_1556,N_29696,N_29625);
xor UO_1557 (O_1557,N_29681,N_29768);
or UO_1558 (O_1558,N_29707,N_29934);
or UO_1559 (O_1559,N_29727,N_29889);
and UO_1560 (O_1560,N_29597,N_29523);
or UO_1561 (O_1561,N_29748,N_29808);
or UO_1562 (O_1562,N_29899,N_29589);
or UO_1563 (O_1563,N_29505,N_29633);
nand UO_1564 (O_1564,N_29828,N_29728);
or UO_1565 (O_1565,N_29579,N_29603);
or UO_1566 (O_1566,N_29509,N_29504);
nand UO_1567 (O_1567,N_29841,N_29741);
nor UO_1568 (O_1568,N_29688,N_29645);
xor UO_1569 (O_1569,N_29857,N_29685);
nand UO_1570 (O_1570,N_29647,N_29923);
and UO_1571 (O_1571,N_29878,N_29769);
nand UO_1572 (O_1572,N_29942,N_29567);
xor UO_1573 (O_1573,N_29914,N_29616);
nand UO_1574 (O_1574,N_29754,N_29832);
nor UO_1575 (O_1575,N_29520,N_29712);
xor UO_1576 (O_1576,N_29720,N_29897);
and UO_1577 (O_1577,N_29593,N_29562);
and UO_1578 (O_1578,N_29678,N_29600);
xor UO_1579 (O_1579,N_29717,N_29837);
and UO_1580 (O_1580,N_29761,N_29517);
or UO_1581 (O_1581,N_29578,N_29815);
nand UO_1582 (O_1582,N_29837,N_29803);
xnor UO_1583 (O_1583,N_29874,N_29796);
nand UO_1584 (O_1584,N_29929,N_29679);
nand UO_1585 (O_1585,N_29876,N_29877);
xnor UO_1586 (O_1586,N_29994,N_29654);
or UO_1587 (O_1587,N_29980,N_29589);
xnor UO_1588 (O_1588,N_29677,N_29632);
nand UO_1589 (O_1589,N_29614,N_29569);
nor UO_1590 (O_1590,N_29818,N_29746);
or UO_1591 (O_1591,N_29971,N_29679);
nand UO_1592 (O_1592,N_29542,N_29590);
nand UO_1593 (O_1593,N_29927,N_29621);
or UO_1594 (O_1594,N_29572,N_29949);
and UO_1595 (O_1595,N_29545,N_29919);
or UO_1596 (O_1596,N_29828,N_29836);
xnor UO_1597 (O_1597,N_29501,N_29579);
nand UO_1598 (O_1598,N_29662,N_29769);
nand UO_1599 (O_1599,N_29594,N_29745);
and UO_1600 (O_1600,N_29647,N_29625);
or UO_1601 (O_1601,N_29813,N_29668);
nor UO_1602 (O_1602,N_29697,N_29508);
xor UO_1603 (O_1603,N_29783,N_29629);
nor UO_1604 (O_1604,N_29645,N_29977);
nor UO_1605 (O_1605,N_29716,N_29747);
or UO_1606 (O_1606,N_29925,N_29654);
or UO_1607 (O_1607,N_29941,N_29596);
xor UO_1608 (O_1608,N_29899,N_29649);
nand UO_1609 (O_1609,N_29550,N_29862);
nand UO_1610 (O_1610,N_29702,N_29561);
xnor UO_1611 (O_1611,N_29629,N_29679);
nand UO_1612 (O_1612,N_29527,N_29873);
xnor UO_1613 (O_1613,N_29509,N_29935);
or UO_1614 (O_1614,N_29951,N_29710);
or UO_1615 (O_1615,N_29957,N_29512);
nor UO_1616 (O_1616,N_29782,N_29582);
nand UO_1617 (O_1617,N_29640,N_29950);
and UO_1618 (O_1618,N_29742,N_29774);
nand UO_1619 (O_1619,N_29647,N_29524);
nor UO_1620 (O_1620,N_29610,N_29742);
and UO_1621 (O_1621,N_29867,N_29951);
xor UO_1622 (O_1622,N_29882,N_29678);
nand UO_1623 (O_1623,N_29621,N_29596);
and UO_1624 (O_1624,N_29672,N_29509);
nor UO_1625 (O_1625,N_29856,N_29997);
xor UO_1626 (O_1626,N_29671,N_29514);
and UO_1627 (O_1627,N_29935,N_29713);
and UO_1628 (O_1628,N_29523,N_29502);
xor UO_1629 (O_1629,N_29580,N_29791);
nor UO_1630 (O_1630,N_29799,N_29999);
nor UO_1631 (O_1631,N_29558,N_29527);
nor UO_1632 (O_1632,N_29827,N_29673);
nor UO_1633 (O_1633,N_29632,N_29565);
xnor UO_1634 (O_1634,N_29514,N_29935);
and UO_1635 (O_1635,N_29982,N_29908);
nand UO_1636 (O_1636,N_29826,N_29554);
or UO_1637 (O_1637,N_29518,N_29953);
or UO_1638 (O_1638,N_29852,N_29979);
and UO_1639 (O_1639,N_29608,N_29667);
or UO_1640 (O_1640,N_29594,N_29795);
and UO_1641 (O_1641,N_29550,N_29887);
nand UO_1642 (O_1642,N_29665,N_29836);
or UO_1643 (O_1643,N_29993,N_29950);
nor UO_1644 (O_1644,N_29730,N_29891);
nand UO_1645 (O_1645,N_29991,N_29632);
xor UO_1646 (O_1646,N_29952,N_29894);
xnor UO_1647 (O_1647,N_29841,N_29708);
and UO_1648 (O_1648,N_29949,N_29665);
nor UO_1649 (O_1649,N_29840,N_29620);
or UO_1650 (O_1650,N_29877,N_29884);
xnor UO_1651 (O_1651,N_29520,N_29923);
nor UO_1652 (O_1652,N_29803,N_29590);
nor UO_1653 (O_1653,N_29975,N_29907);
nor UO_1654 (O_1654,N_29842,N_29838);
and UO_1655 (O_1655,N_29700,N_29654);
nand UO_1656 (O_1656,N_29764,N_29657);
nand UO_1657 (O_1657,N_29634,N_29648);
nor UO_1658 (O_1658,N_29894,N_29706);
nor UO_1659 (O_1659,N_29604,N_29924);
nor UO_1660 (O_1660,N_29531,N_29564);
nor UO_1661 (O_1661,N_29619,N_29877);
nand UO_1662 (O_1662,N_29764,N_29647);
xnor UO_1663 (O_1663,N_29634,N_29616);
xor UO_1664 (O_1664,N_29885,N_29797);
or UO_1665 (O_1665,N_29698,N_29883);
xor UO_1666 (O_1666,N_29580,N_29940);
xnor UO_1667 (O_1667,N_29624,N_29773);
nand UO_1668 (O_1668,N_29964,N_29966);
and UO_1669 (O_1669,N_29892,N_29549);
and UO_1670 (O_1670,N_29782,N_29598);
nand UO_1671 (O_1671,N_29642,N_29983);
nor UO_1672 (O_1672,N_29536,N_29630);
and UO_1673 (O_1673,N_29926,N_29606);
and UO_1674 (O_1674,N_29635,N_29973);
xnor UO_1675 (O_1675,N_29532,N_29757);
nand UO_1676 (O_1676,N_29847,N_29579);
nand UO_1677 (O_1677,N_29575,N_29739);
or UO_1678 (O_1678,N_29813,N_29825);
or UO_1679 (O_1679,N_29506,N_29665);
nand UO_1680 (O_1680,N_29898,N_29948);
or UO_1681 (O_1681,N_29951,N_29606);
nand UO_1682 (O_1682,N_29888,N_29775);
or UO_1683 (O_1683,N_29524,N_29664);
or UO_1684 (O_1684,N_29884,N_29782);
nand UO_1685 (O_1685,N_29974,N_29557);
or UO_1686 (O_1686,N_29560,N_29648);
or UO_1687 (O_1687,N_29738,N_29930);
nor UO_1688 (O_1688,N_29673,N_29973);
or UO_1689 (O_1689,N_29778,N_29541);
nand UO_1690 (O_1690,N_29735,N_29527);
xnor UO_1691 (O_1691,N_29865,N_29983);
nand UO_1692 (O_1692,N_29759,N_29692);
or UO_1693 (O_1693,N_29605,N_29687);
and UO_1694 (O_1694,N_29502,N_29944);
and UO_1695 (O_1695,N_29928,N_29994);
or UO_1696 (O_1696,N_29834,N_29752);
nor UO_1697 (O_1697,N_29840,N_29791);
or UO_1698 (O_1698,N_29905,N_29934);
or UO_1699 (O_1699,N_29930,N_29726);
or UO_1700 (O_1700,N_29825,N_29758);
xor UO_1701 (O_1701,N_29714,N_29951);
and UO_1702 (O_1702,N_29613,N_29703);
nand UO_1703 (O_1703,N_29860,N_29742);
and UO_1704 (O_1704,N_29534,N_29686);
and UO_1705 (O_1705,N_29927,N_29508);
xor UO_1706 (O_1706,N_29738,N_29612);
nand UO_1707 (O_1707,N_29840,N_29685);
xnor UO_1708 (O_1708,N_29903,N_29576);
xnor UO_1709 (O_1709,N_29566,N_29877);
nor UO_1710 (O_1710,N_29776,N_29522);
and UO_1711 (O_1711,N_29965,N_29633);
or UO_1712 (O_1712,N_29774,N_29806);
xor UO_1713 (O_1713,N_29884,N_29755);
xnor UO_1714 (O_1714,N_29612,N_29779);
nand UO_1715 (O_1715,N_29795,N_29624);
nor UO_1716 (O_1716,N_29756,N_29742);
nor UO_1717 (O_1717,N_29876,N_29825);
and UO_1718 (O_1718,N_29839,N_29523);
or UO_1719 (O_1719,N_29991,N_29765);
or UO_1720 (O_1720,N_29809,N_29846);
or UO_1721 (O_1721,N_29731,N_29963);
nand UO_1722 (O_1722,N_29861,N_29636);
and UO_1723 (O_1723,N_29817,N_29736);
or UO_1724 (O_1724,N_29896,N_29821);
nor UO_1725 (O_1725,N_29715,N_29679);
xnor UO_1726 (O_1726,N_29909,N_29654);
nor UO_1727 (O_1727,N_29982,N_29535);
or UO_1728 (O_1728,N_29655,N_29576);
nor UO_1729 (O_1729,N_29869,N_29715);
and UO_1730 (O_1730,N_29692,N_29548);
or UO_1731 (O_1731,N_29606,N_29551);
and UO_1732 (O_1732,N_29543,N_29841);
xor UO_1733 (O_1733,N_29741,N_29916);
xnor UO_1734 (O_1734,N_29656,N_29580);
and UO_1735 (O_1735,N_29507,N_29812);
and UO_1736 (O_1736,N_29814,N_29907);
and UO_1737 (O_1737,N_29537,N_29967);
xor UO_1738 (O_1738,N_29573,N_29895);
or UO_1739 (O_1739,N_29837,N_29555);
and UO_1740 (O_1740,N_29636,N_29677);
xor UO_1741 (O_1741,N_29643,N_29563);
and UO_1742 (O_1742,N_29720,N_29995);
xnor UO_1743 (O_1743,N_29542,N_29630);
nand UO_1744 (O_1744,N_29949,N_29639);
nor UO_1745 (O_1745,N_29678,N_29652);
or UO_1746 (O_1746,N_29989,N_29925);
nor UO_1747 (O_1747,N_29690,N_29929);
or UO_1748 (O_1748,N_29528,N_29965);
xnor UO_1749 (O_1749,N_29526,N_29669);
nand UO_1750 (O_1750,N_29677,N_29838);
and UO_1751 (O_1751,N_29911,N_29839);
xnor UO_1752 (O_1752,N_29729,N_29798);
or UO_1753 (O_1753,N_29518,N_29723);
nor UO_1754 (O_1754,N_29506,N_29851);
nand UO_1755 (O_1755,N_29967,N_29656);
or UO_1756 (O_1756,N_29915,N_29842);
nand UO_1757 (O_1757,N_29761,N_29567);
nand UO_1758 (O_1758,N_29679,N_29993);
xor UO_1759 (O_1759,N_29996,N_29788);
nand UO_1760 (O_1760,N_29628,N_29969);
xor UO_1761 (O_1761,N_29716,N_29757);
nand UO_1762 (O_1762,N_29812,N_29668);
nand UO_1763 (O_1763,N_29630,N_29987);
and UO_1764 (O_1764,N_29645,N_29560);
and UO_1765 (O_1765,N_29534,N_29811);
nor UO_1766 (O_1766,N_29973,N_29807);
xor UO_1767 (O_1767,N_29543,N_29686);
and UO_1768 (O_1768,N_29873,N_29982);
or UO_1769 (O_1769,N_29892,N_29929);
nor UO_1770 (O_1770,N_29639,N_29948);
xor UO_1771 (O_1771,N_29833,N_29983);
xnor UO_1772 (O_1772,N_29916,N_29673);
and UO_1773 (O_1773,N_29586,N_29627);
xnor UO_1774 (O_1774,N_29645,N_29870);
nand UO_1775 (O_1775,N_29707,N_29679);
and UO_1776 (O_1776,N_29807,N_29969);
nand UO_1777 (O_1777,N_29661,N_29616);
and UO_1778 (O_1778,N_29893,N_29909);
or UO_1779 (O_1779,N_29657,N_29624);
and UO_1780 (O_1780,N_29577,N_29698);
and UO_1781 (O_1781,N_29555,N_29521);
or UO_1782 (O_1782,N_29706,N_29713);
xor UO_1783 (O_1783,N_29527,N_29553);
and UO_1784 (O_1784,N_29982,N_29582);
xor UO_1785 (O_1785,N_29772,N_29815);
and UO_1786 (O_1786,N_29619,N_29671);
nor UO_1787 (O_1787,N_29976,N_29569);
nor UO_1788 (O_1788,N_29713,N_29517);
xor UO_1789 (O_1789,N_29975,N_29968);
or UO_1790 (O_1790,N_29802,N_29747);
xnor UO_1791 (O_1791,N_29681,N_29964);
nor UO_1792 (O_1792,N_29987,N_29839);
and UO_1793 (O_1793,N_29767,N_29728);
nor UO_1794 (O_1794,N_29675,N_29569);
and UO_1795 (O_1795,N_29956,N_29503);
and UO_1796 (O_1796,N_29732,N_29580);
nor UO_1797 (O_1797,N_29535,N_29636);
or UO_1798 (O_1798,N_29857,N_29811);
nor UO_1799 (O_1799,N_29884,N_29945);
xor UO_1800 (O_1800,N_29849,N_29719);
nand UO_1801 (O_1801,N_29955,N_29630);
or UO_1802 (O_1802,N_29888,N_29538);
or UO_1803 (O_1803,N_29755,N_29734);
and UO_1804 (O_1804,N_29591,N_29879);
nor UO_1805 (O_1805,N_29621,N_29763);
nand UO_1806 (O_1806,N_29524,N_29646);
or UO_1807 (O_1807,N_29704,N_29922);
nand UO_1808 (O_1808,N_29857,N_29659);
and UO_1809 (O_1809,N_29839,N_29836);
nand UO_1810 (O_1810,N_29791,N_29503);
or UO_1811 (O_1811,N_29972,N_29608);
xor UO_1812 (O_1812,N_29709,N_29598);
nand UO_1813 (O_1813,N_29784,N_29547);
and UO_1814 (O_1814,N_29897,N_29639);
nor UO_1815 (O_1815,N_29963,N_29977);
nand UO_1816 (O_1816,N_29514,N_29714);
nand UO_1817 (O_1817,N_29597,N_29539);
nand UO_1818 (O_1818,N_29695,N_29998);
and UO_1819 (O_1819,N_29727,N_29916);
nor UO_1820 (O_1820,N_29780,N_29761);
and UO_1821 (O_1821,N_29513,N_29510);
or UO_1822 (O_1822,N_29821,N_29510);
or UO_1823 (O_1823,N_29902,N_29959);
and UO_1824 (O_1824,N_29799,N_29718);
nor UO_1825 (O_1825,N_29907,N_29519);
nor UO_1826 (O_1826,N_29580,N_29840);
nor UO_1827 (O_1827,N_29908,N_29603);
xnor UO_1828 (O_1828,N_29943,N_29683);
or UO_1829 (O_1829,N_29885,N_29874);
and UO_1830 (O_1830,N_29724,N_29848);
nor UO_1831 (O_1831,N_29895,N_29687);
nand UO_1832 (O_1832,N_29945,N_29541);
and UO_1833 (O_1833,N_29785,N_29839);
xnor UO_1834 (O_1834,N_29891,N_29582);
xnor UO_1835 (O_1835,N_29770,N_29725);
nand UO_1836 (O_1836,N_29568,N_29936);
xor UO_1837 (O_1837,N_29728,N_29642);
xor UO_1838 (O_1838,N_29681,N_29902);
nor UO_1839 (O_1839,N_29730,N_29582);
nor UO_1840 (O_1840,N_29867,N_29908);
or UO_1841 (O_1841,N_29772,N_29897);
and UO_1842 (O_1842,N_29844,N_29891);
and UO_1843 (O_1843,N_29988,N_29590);
or UO_1844 (O_1844,N_29885,N_29611);
nor UO_1845 (O_1845,N_29883,N_29780);
or UO_1846 (O_1846,N_29560,N_29773);
xor UO_1847 (O_1847,N_29649,N_29705);
nand UO_1848 (O_1848,N_29982,N_29942);
nand UO_1849 (O_1849,N_29893,N_29676);
or UO_1850 (O_1850,N_29842,N_29622);
xnor UO_1851 (O_1851,N_29790,N_29636);
xor UO_1852 (O_1852,N_29528,N_29569);
xnor UO_1853 (O_1853,N_29936,N_29543);
and UO_1854 (O_1854,N_29708,N_29852);
or UO_1855 (O_1855,N_29857,N_29841);
xnor UO_1856 (O_1856,N_29546,N_29972);
xnor UO_1857 (O_1857,N_29759,N_29752);
or UO_1858 (O_1858,N_29789,N_29864);
nand UO_1859 (O_1859,N_29709,N_29836);
xor UO_1860 (O_1860,N_29626,N_29799);
xor UO_1861 (O_1861,N_29934,N_29875);
or UO_1862 (O_1862,N_29585,N_29898);
nor UO_1863 (O_1863,N_29544,N_29643);
xor UO_1864 (O_1864,N_29961,N_29529);
xor UO_1865 (O_1865,N_29835,N_29543);
or UO_1866 (O_1866,N_29611,N_29659);
nor UO_1867 (O_1867,N_29564,N_29778);
xnor UO_1868 (O_1868,N_29987,N_29885);
nand UO_1869 (O_1869,N_29747,N_29653);
and UO_1870 (O_1870,N_29950,N_29577);
xor UO_1871 (O_1871,N_29923,N_29686);
and UO_1872 (O_1872,N_29632,N_29996);
nor UO_1873 (O_1873,N_29690,N_29936);
nor UO_1874 (O_1874,N_29816,N_29961);
nand UO_1875 (O_1875,N_29738,N_29736);
or UO_1876 (O_1876,N_29777,N_29722);
nand UO_1877 (O_1877,N_29743,N_29817);
nor UO_1878 (O_1878,N_29843,N_29940);
and UO_1879 (O_1879,N_29983,N_29688);
xnor UO_1880 (O_1880,N_29966,N_29978);
nor UO_1881 (O_1881,N_29816,N_29567);
nor UO_1882 (O_1882,N_29967,N_29942);
nor UO_1883 (O_1883,N_29760,N_29895);
or UO_1884 (O_1884,N_29615,N_29526);
nor UO_1885 (O_1885,N_29981,N_29631);
nor UO_1886 (O_1886,N_29699,N_29640);
nor UO_1887 (O_1887,N_29781,N_29739);
xnor UO_1888 (O_1888,N_29851,N_29957);
nor UO_1889 (O_1889,N_29932,N_29759);
and UO_1890 (O_1890,N_29745,N_29884);
nand UO_1891 (O_1891,N_29761,N_29806);
nor UO_1892 (O_1892,N_29784,N_29693);
xor UO_1893 (O_1893,N_29579,N_29689);
nand UO_1894 (O_1894,N_29750,N_29640);
xor UO_1895 (O_1895,N_29872,N_29927);
xnor UO_1896 (O_1896,N_29602,N_29688);
xnor UO_1897 (O_1897,N_29703,N_29623);
xnor UO_1898 (O_1898,N_29654,N_29735);
nor UO_1899 (O_1899,N_29578,N_29866);
nor UO_1900 (O_1900,N_29513,N_29653);
or UO_1901 (O_1901,N_29797,N_29576);
xor UO_1902 (O_1902,N_29639,N_29954);
and UO_1903 (O_1903,N_29844,N_29906);
or UO_1904 (O_1904,N_29672,N_29665);
nand UO_1905 (O_1905,N_29812,N_29792);
or UO_1906 (O_1906,N_29749,N_29582);
and UO_1907 (O_1907,N_29543,N_29996);
nor UO_1908 (O_1908,N_29752,N_29556);
nand UO_1909 (O_1909,N_29997,N_29920);
or UO_1910 (O_1910,N_29596,N_29945);
nand UO_1911 (O_1911,N_29854,N_29833);
xnor UO_1912 (O_1912,N_29631,N_29997);
xor UO_1913 (O_1913,N_29841,N_29617);
or UO_1914 (O_1914,N_29636,N_29537);
or UO_1915 (O_1915,N_29610,N_29614);
xnor UO_1916 (O_1916,N_29566,N_29658);
nor UO_1917 (O_1917,N_29862,N_29967);
nand UO_1918 (O_1918,N_29546,N_29813);
nand UO_1919 (O_1919,N_29975,N_29953);
or UO_1920 (O_1920,N_29505,N_29878);
nand UO_1921 (O_1921,N_29661,N_29573);
or UO_1922 (O_1922,N_29644,N_29904);
nor UO_1923 (O_1923,N_29674,N_29961);
xor UO_1924 (O_1924,N_29979,N_29740);
nand UO_1925 (O_1925,N_29831,N_29840);
or UO_1926 (O_1926,N_29837,N_29520);
nor UO_1927 (O_1927,N_29868,N_29708);
xnor UO_1928 (O_1928,N_29668,N_29759);
and UO_1929 (O_1929,N_29769,N_29826);
nand UO_1930 (O_1930,N_29587,N_29878);
xor UO_1931 (O_1931,N_29686,N_29860);
xor UO_1932 (O_1932,N_29922,N_29968);
nor UO_1933 (O_1933,N_29809,N_29598);
or UO_1934 (O_1934,N_29755,N_29723);
nand UO_1935 (O_1935,N_29538,N_29675);
nor UO_1936 (O_1936,N_29630,N_29853);
xor UO_1937 (O_1937,N_29709,N_29965);
xnor UO_1938 (O_1938,N_29983,N_29565);
nand UO_1939 (O_1939,N_29665,N_29972);
and UO_1940 (O_1940,N_29947,N_29987);
nor UO_1941 (O_1941,N_29604,N_29667);
or UO_1942 (O_1942,N_29688,N_29703);
nor UO_1943 (O_1943,N_29532,N_29769);
nor UO_1944 (O_1944,N_29727,N_29753);
and UO_1945 (O_1945,N_29963,N_29847);
xor UO_1946 (O_1946,N_29750,N_29837);
or UO_1947 (O_1947,N_29962,N_29683);
or UO_1948 (O_1948,N_29946,N_29819);
nor UO_1949 (O_1949,N_29841,N_29825);
or UO_1950 (O_1950,N_29896,N_29613);
nand UO_1951 (O_1951,N_29747,N_29540);
or UO_1952 (O_1952,N_29614,N_29750);
nand UO_1953 (O_1953,N_29927,N_29792);
nand UO_1954 (O_1954,N_29815,N_29681);
nand UO_1955 (O_1955,N_29782,N_29993);
and UO_1956 (O_1956,N_29882,N_29645);
nand UO_1957 (O_1957,N_29774,N_29972);
nand UO_1958 (O_1958,N_29951,N_29931);
xor UO_1959 (O_1959,N_29913,N_29794);
nor UO_1960 (O_1960,N_29617,N_29962);
and UO_1961 (O_1961,N_29565,N_29607);
nand UO_1962 (O_1962,N_29704,N_29823);
and UO_1963 (O_1963,N_29536,N_29720);
or UO_1964 (O_1964,N_29630,N_29755);
nor UO_1965 (O_1965,N_29996,N_29946);
and UO_1966 (O_1966,N_29628,N_29875);
nand UO_1967 (O_1967,N_29624,N_29775);
nand UO_1968 (O_1968,N_29545,N_29876);
nor UO_1969 (O_1969,N_29957,N_29874);
or UO_1970 (O_1970,N_29649,N_29598);
and UO_1971 (O_1971,N_29660,N_29917);
and UO_1972 (O_1972,N_29916,N_29918);
and UO_1973 (O_1973,N_29651,N_29974);
xor UO_1974 (O_1974,N_29849,N_29547);
or UO_1975 (O_1975,N_29813,N_29580);
and UO_1976 (O_1976,N_29688,N_29743);
xor UO_1977 (O_1977,N_29833,N_29837);
or UO_1978 (O_1978,N_29955,N_29510);
nor UO_1979 (O_1979,N_29536,N_29657);
and UO_1980 (O_1980,N_29879,N_29872);
nor UO_1981 (O_1981,N_29612,N_29883);
or UO_1982 (O_1982,N_29504,N_29950);
xnor UO_1983 (O_1983,N_29604,N_29852);
xor UO_1984 (O_1984,N_29782,N_29528);
xor UO_1985 (O_1985,N_29511,N_29502);
nor UO_1986 (O_1986,N_29504,N_29961);
nand UO_1987 (O_1987,N_29798,N_29668);
xor UO_1988 (O_1988,N_29881,N_29719);
nor UO_1989 (O_1989,N_29784,N_29773);
nor UO_1990 (O_1990,N_29932,N_29717);
nand UO_1991 (O_1991,N_29547,N_29633);
or UO_1992 (O_1992,N_29546,N_29708);
xor UO_1993 (O_1993,N_29730,N_29594);
nand UO_1994 (O_1994,N_29874,N_29593);
xor UO_1995 (O_1995,N_29613,N_29986);
or UO_1996 (O_1996,N_29900,N_29598);
or UO_1997 (O_1997,N_29656,N_29778);
xnor UO_1998 (O_1998,N_29957,N_29721);
or UO_1999 (O_1999,N_29913,N_29993);
nand UO_2000 (O_2000,N_29642,N_29830);
xnor UO_2001 (O_2001,N_29905,N_29799);
nor UO_2002 (O_2002,N_29646,N_29983);
nor UO_2003 (O_2003,N_29876,N_29874);
nand UO_2004 (O_2004,N_29713,N_29830);
nand UO_2005 (O_2005,N_29871,N_29960);
xnor UO_2006 (O_2006,N_29578,N_29550);
nand UO_2007 (O_2007,N_29682,N_29742);
xor UO_2008 (O_2008,N_29835,N_29895);
nor UO_2009 (O_2009,N_29868,N_29950);
nand UO_2010 (O_2010,N_29588,N_29987);
xor UO_2011 (O_2011,N_29833,N_29629);
nor UO_2012 (O_2012,N_29675,N_29635);
nand UO_2013 (O_2013,N_29911,N_29605);
nor UO_2014 (O_2014,N_29966,N_29909);
nor UO_2015 (O_2015,N_29537,N_29780);
xor UO_2016 (O_2016,N_29773,N_29650);
xor UO_2017 (O_2017,N_29640,N_29812);
nor UO_2018 (O_2018,N_29814,N_29520);
or UO_2019 (O_2019,N_29588,N_29566);
xnor UO_2020 (O_2020,N_29550,N_29735);
and UO_2021 (O_2021,N_29641,N_29915);
nor UO_2022 (O_2022,N_29769,N_29512);
or UO_2023 (O_2023,N_29721,N_29923);
xor UO_2024 (O_2024,N_29934,N_29815);
nor UO_2025 (O_2025,N_29735,N_29910);
nand UO_2026 (O_2026,N_29594,N_29609);
nand UO_2027 (O_2027,N_29636,N_29944);
nand UO_2028 (O_2028,N_29639,N_29857);
nand UO_2029 (O_2029,N_29910,N_29746);
and UO_2030 (O_2030,N_29692,N_29912);
nor UO_2031 (O_2031,N_29751,N_29599);
xnor UO_2032 (O_2032,N_29551,N_29512);
nand UO_2033 (O_2033,N_29691,N_29883);
nor UO_2034 (O_2034,N_29552,N_29970);
nand UO_2035 (O_2035,N_29595,N_29542);
nand UO_2036 (O_2036,N_29636,N_29729);
xnor UO_2037 (O_2037,N_29985,N_29798);
nor UO_2038 (O_2038,N_29647,N_29956);
nand UO_2039 (O_2039,N_29808,N_29709);
nor UO_2040 (O_2040,N_29643,N_29729);
or UO_2041 (O_2041,N_29857,N_29714);
or UO_2042 (O_2042,N_29536,N_29829);
nand UO_2043 (O_2043,N_29731,N_29895);
xor UO_2044 (O_2044,N_29746,N_29596);
nor UO_2045 (O_2045,N_29923,N_29517);
and UO_2046 (O_2046,N_29809,N_29581);
xnor UO_2047 (O_2047,N_29936,N_29962);
and UO_2048 (O_2048,N_29805,N_29846);
xor UO_2049 (O_2049,N_29645,N_29754);
and UO_2050 (O_2050,N_29536,N_29909);
xor UO_2051 (O_2051,N_29988,N_29999);
nand UO_2052 (O_2052,N_29866,N_29832);
xor UO_2053 (O_2053,N_29668,N_29591);
and UO_2054 (O_2054,N_29524,N_29605);
or UO_2055 (O_2055,N_29530,N_29907);
nor UO_2056 (O_2056,N_29940,N_29585);
xnor UO_2057 (O_2057,N_29559,N_29703);
xnor UO_2058 (O_2058,N_29581,N_29876);
and UO_2059 (O_2059,N_29778,N_29973);
or UO_2060 (O_2060,N_29633,N_29632);
nor UO_2061 (O_2061,N_29633,N_29726);
and UO_2062 (O_2062,N_29854,N_29874);
nand UO_2063 (O_2063,N_29793,N_29547);
nor UO_2064 (O_2064,N_29655,N_29992);
nand UO_2065 (O_2065,N_29820,N_29958);
and UO_2066 (O_2066,N_29843,N_29593);
nor UO_2067 (O_2067,N_29825,N_29568);
xnor UO_2068 (O_2068,N_29973,N_29585);
nor UO_2069 (O_2069,N_29958,N_29895);
nor UO_2070 (O_2070,N_29563,N_29515);
or UO_2071 (O_2071,N_29687,N_29719);
or UO_2072 (O_2072,N_29811,N_29852);
xor UO_2073 (O_2073,N_29669,N_29620);
or UO_2074 (O_2074,N_29728,N_29710);
xor UO_2075 (O_2075,N_29518,N_29888);
nand UO_2076 (O_2076,N_29871,N_29644);
or UO_2077 (O_2077,N_29520,N_29576);
and UO_2078 (O_2078,N_29969,N_29909);
nand UO_2079 (O_2079,N_29742,N_29658);
and UO_2080 (O_2080,N_29876,N_29628);
or UO_2081 (O_2081,N_29927,N_29776);
and UO_2082 (O_2082,N_29990,N_29555);
xor UO_2083 (O_2083,N_29580,N_29597);
nor UO_2084 (O_2084,N_29919,N_29658);
xnor UO_2085 (O_2085,N_29930,N_29571);
or UO_2086 (O_2086,N_29799,N_29981);
xor UO_2087 (O_2087,N_29677,N_29739);
nand UO_2088 (O_2088,N_29811,N_29862);
nor UO_2089 (O_2089,N_29652,N_29823);
nand UO_2090 (O_2090,N_29931,N_29983);
or UO_2091 (O_2091,N_29502,N_29535);
or UO_2092 (O_2092,N_29591,N_29913);
and UO_2093 (O_2093,N_29856,N_29844);
nor UO_2094 (O_2094,N_29921,N_29720);
xor UO_2095 (O_2095,N_29616,N_29875);
or UO_2096 (O_2096,N_29743,N_29608);
xnor UO_2097 (O_2097,N_29533,N_29779);
xnor UO_2098 (O_2098,N_29561,N_29591);
nor UO_2099 (O_2099,N_29583,N_29668);
nand UO_2100 (O_2100,N_29554,N_29536);
or UO_2101 (O_2101,N_29811,N_29694);
and UO_2102 (O_2102,N_29816,N_29578);
or UO_2103 (O_2103,N_29691,N_29674);
xnor UO_2104 (O_2104,N_29650,N_29501);
nand UO_2105 (O_2105,N_29652,N_29679);
nand UO_2106 (O_2106,N_29604,N_29547);
nand UO_2107 (O_2107,N_29651,N_29771);
nand UO_2108 (O_2108,N_29777,N_29951);
xor UO_2109 (O_2109,N_29824,N_29840);
xor UO_2110 (O_2110,N_29838,N_29752);
nor UO_2111 (O_2111,N_29907,N_29827);
nor UO_2112 (O_2112,N_29617,N_29796);
and UO_2113 (O_2113,N_29719,N_29636);
and UO_2114 (O_2114,N_29883,N_29841);
nor UO_2115 (O_2115,N_29590,N_29962);
nand UO_2116 (O_2116,N_29767,N_29509);
nand UO_2117 (O_2117,N_29947,N_29811);
xnor UO_2118 (O_2118,N_29988,N_29544);
nand UO_2119 (O_2119,N_29754,N_29786);
xnor UO_2120 (O_2120,N_29823,N_29760);
or UO_2121 (O_2121,N_29923,N_29546);
and UO_2122 (O_2122,N_29701,N_29545);
and UO_2123 (O_2123,N_29721,N_29699);
or UO_2124 (O_2124,N_29736,N_29575);
nand UO_2125 (O_2125,N_29745,N_29998);
nor UO_2126 (O_2126,N_29898,N_29568);
nand UO_2127 (O_2127,N_29538,N_29849);
and UO_2128 (O_2128,N_29958,N_29785);
nand UO_2129 (O_2129,N_29832,N_29682);
nand UO_2130 (O_2130,N_29951,N_29653);
xnor UO_2131 (O_2131,N_29706,N_29858);
xor UO_2132 (O_2132,N_29827,N_29704);
and UO_2133 (O_2133,N_29733,N_29905);
or UO_2134 (O_2134,N_29966,N_29726);
or UO_2135 (O_2135,N_29978,N_29986);
xor UO_2136 (O_2136,N_29751,N_29567);
and UO_2137 (O_2137,N_29881,N_29970);
and UO_2138 (O_2138,N_29790,N_29920);
xnor UO_2139 (O_2139,N_29606,N_29695);
or UO_2140 (O_2140,N_29927,N_29939);
or UO_2141 (O_2141,N_29512,N_29546);
or UO_2142 (O_2142,N_29741,N_29767);
and UO_2143 (O_2143,N_29985,N_29746);
nand UO_2144 (O_2144,N_29696,N_29693);
xnor UO_2145 (O_2145,N_29840,N_29588);
and UO_2146 (O_2146,N_29556,N_29797);
nor UO_2147 (O_2147,N_29899,N_29609);
nor UO_2148 (O_2148,N_29781,N_29683);
nor UO_2149 (O_2149,N_29595,N_29536);
and UO_2150 (O_2150,N_29909,N_29892);
or UO_2151 (O_2151,N_29544,N_29956);
nand UO_2152 (O_2152,N_29615,N_29547);
nand UO_2153 (O_2153,N_29508,N_29832);
nor UO_2154 (O_2154,N_29955,N_29803);
or UO_2155 (O_2155,N_29689,N_29934);
xor UO_2156 (O_2156,N_29836,N_29570);
nor UO_2157 (O_2157,N_29822,N_29910);
and UO_2158 (O_2158,N_29718,N_29724);
nor UO_2159 (O_2159,N_29792,N_29876);
nand UO_2160 (O_2160,N_29790,N_29558);
or UO_2161 (O_2161,N_29843,N_29690);
nor UO_2162 (O_2162,N_29521,N_29706);
and UO_2163 (O_2163,N_29739,N_29760);
nor UO_2164 (O_2164,N_29576,N_29825);
or UO_2165 (O_2165,N_29957,N_29609);
and UO_2166 (O_2166,N_29865,N_29753);
xor UO_2167 (O_2167,N_29620,N_29637);
and UO_2168 (O_2168,N_29504,N_29836);
xnor UO_2169 (O_2169,N_29859,N_29858);
xor UO_2170 (O_2170,N_29606,N_29642);
nand UO_2171 (O_2171,N_29705,N_29622);
nor UO_2172 (O_2172,N_29728,N_29840);
and UO_2173 (O_2173,N_29617,N_29891);
nand UO_2174 (O_2174,N_29724,N_29575);
and UO_2175 (O_2175,N_29625,N_29754);
nand UO_2176 (O_2176,N_29767,N_29657);
and UO_2177 (O_2177,N_29821,N_29859);
and UO_2178 (O_2178,N_29569,N_29505);
xnor UO_2179 (O_2179,N_29633,N_29906);
and UO_2180 (O_2180,N_29632,N_29621);
xor UO_2181 (O_2181,N_29787,N_29763);
or UO_2182 (O_2182,N_29983,N_29854);
nand UO_2183 (O_2183,N_29583,N_29545);
nand UO_2184 (O_2184,N_29588,N_29681);
nand UO_2185 (O_2185,N_29694,N_29940);
xor UO_2186 (O_2186,N_29734,N_29927);
xor UO_2187 (O_2187,N_29930,N_29681);
and UO_2188 (O_2188,N_29710,N_29592);
and UO_2189 (O_2189,N_29727,N_29553);
nand UO_2190 (O_2190,N_29865,N_29978);
nand UO_2191 (O_2191,N_29658,N_29511);
nor UO_2192 (O_2192,N_29749,N_29607);
or UO_2193 (O_2193,N_29722,N_29763);
or UO_2194 (O_2194,N_29959,N_29672);
or UO_2195 (O_2195,N_29657,N_29667);
xor UO_2196 (O_2196,N_29549,N_29633);
nand UO_2197 (O_2197,N_29888,N_29565);
nor UO_2198 (O_2198,N_29688,N_29647);
nor UO_2199 (O_2199,N_29976,N_29609);
nor UO_2200 (O_2200,N_29774,N_29997);
nor UO_2201 (O_2201,N_29737,N_29569);
xnor UO_2202 (O_2202,N_29704,N_29880);
nand UO_2203 (O_2203,N_29836,N_29546);
nor UO_2204 (O_2204,N_29595,N_29839);
and UO_2205 (O_2205,N_29727,N_29655);
nor UO_2206 (O_2206,N_29762,N_29786);
nand UO_2207 (O_2207,N_29963,N_29685);
nand UO_2208 (O_2208,N_29992,N_29575);
and UO_2209 (O_2209,N_29823,N_29693);
xor UO_2210 (O_2210,N_29886,N_29631);
nor UO_2211 (O_2211,N_29800,N_29759);
nand UO_2212 (O_2212,N_29503,N_29623);
nand UO_2213 (O_2213,N_29643,N_29652);
or UO_2214 (O_2214,N_29842,N_29850);
nor UO_2215 (O_2215,N_29732,N_29720);
xnor UO_2216 (O_2216,N_29660,N_29740);
nor UO_2217 (O_2217,N_29633,N_29566);
nor UO_2218 (O_2218,N_29831,N_29717);
xnor UO_2219 (O_2219,N_29828,N_29649);
nor UO_2220 (O_2220,N_29526,N_29540);
and UO_2221 (O_2221,N_29825,N_29865);
or UO_2222 (O_2222,N_29511,N_29628);
nand UO_2223 (O_2223,N_29522,N_29920);
and UO_2224 (O_2224,N_29824,N_29563);
xor UO_2225 (O_2225,N_29969,N_29973);
xnor UO_2226 (O_2226,N_29681,N_29743);
or UO_2227 (O_2227,N_29750,N_29656);
nor UO_2228 (O_2228,N_29969,N_29992);
nand UO_2229 (O_2229,N_29770,N_29955);
nand UO_2230 (O_2230,N_29823,N_29694);
nand UO_2231 (O_2231,N_29907,N_29696);
nand UO_2232 (O_2232,N_29603,N_29502);
or UO_2233 (O_2233,N_29743,N_29686);
nand UO_2234 (O_2234,N_29722,N_29918);
nand UO_2235 (O_2235,N_29756,N_29590);
or UO_2236 (O_2236,N_29792,N_29619);
nor UO_2237 (O_2237,N_29607,N_29906);
xnor UO_2238 (O_2238,N_29746,N_29628);
and UO_2239 (O_2239,N_29841,N_29683);
nor UO_2240 (O_2240,N_29633,N_29746);
and UO_2241 (O_2241,N_29822,N_29513);
xor UO_2242 (O_2242,N_29730,N_29812);
nor UO_2243 (O_2243,N_29519,N_29823);
or UO_2244 (O_2244,N_29968,N_29749);
nand UO_2245 (O_2245,N_29577,N_29580);
or UO_2246 (O_2246,N_29981,N_29585);
or UO_2247 (O_2247,N_29971,N_29967);
nor UO_2248 (O_2248,N_29990,N_29805);
nand UO_2249 (O_2249,N_29674,N_29631);
and UO_2250 (O_2250,N_29760,N_29916);
xor UO_2251 (O_2251,N_29695,N_29921);
nor UO_2252 (O_2252,N_29865,N_29603);
nor UO_2253 (O_2253,N_29652,N_29861);
nor UO_2254 (O_2254,N_29630,N_29726);
nor UO_2255 (O_2255,N_29989,N_29968);
nor UO_2256 (O_2256,N_29972,N_29904);
and UO_2257 (O_2257,N_29802,N_29943);
nand UO_2258 (O_2258,N_29995,N_29858);
nor UO_2259 (O_2259,N_29851,N_29840);
xor UO_2260 (O_2260,N_29845,N_29760);
xor UO_2261 (O_2261,N_29515,N_29938);
nor UO_2262 (O_2262,N_29822,N_29861);
and UO_2263 (O_2263,N_29979,N_29611);
xnor UO_2264 (O_2264,N_29528,N_29768);
and UO_2265 (O_2265,N_29906,N_29835);
xnor UO_2266 (O_2266,N_29990,N_29952);
or UO_2267 (O_2267,N_29916,N_29945);
and UO_2268 (O_2268,N_29697,N_29793);
nor UO_2269 (O_2269,N_29691,N_29636);
and UO_2270 (O_2270,N_29689,N_29762);
xor UO_2271 (O_2271,N_29638,N_29668);
or UO_2272 (O_2272,N_29546,N_29788);
nor UO_2273 (O_2273,N_29869,N_29928);
or UO_2274 (O_2274,N_29949,N_29577);
xnor UO_2275 (O_2275,N_29749,N_29657);
or UO_2276 (O_2276,N_29972,N_29718);
nand UO_2277 (O_2277,N_29991,N_29584);
and UO_2278 (O_2278,N_29749,N_29539);
xnor UO_2279 (O_2279,N_29658,N_29745);
and UO_2280 (O_2280,N_29835,N_29972);
nand UO_2281 (O_2281,N_29635,N_29669);
nor UO_2282 (O_2282,N_29840,N_29767);
nand UO_2283 (O_2283,N_29508,N_29933);
xor UO_2284 (O_2284,N_29596,N_29549);
xor UO_2285 (O_2285,N_29502,N_29620);
nor UO_2286 (O_2286,N_29592,N_29981);
xnor UO_2287 (O_2287,N_29544,N_29628);
or UO_2288 (O_2288,N_29843,N_29741);
nand UO_2289 (O_2289,N_29571,N_29598);
and UO_2290 (O_2290,N_29666,N_29509);
nand UO_2291 (O_2291,N_29504,N_29833);
and UO_2292 (O_2292,N_29980,N_29729);
nand UO_2293 (O_2293,N_29606,N_29812);
nand UO_2294 (O_2294,N_29963,N_29671);
or UO_2295 (O_2295,N_29732,N_29617);
nand UO_2296 (O_2296,N_29756,N_29865);
or UO_2297 (O_2297,N_29518,N_29990);
xor UO_2298 (O_2298,N_29712,N_29814);
or UO_2299 (O_2299,N_29698,N_29530);
xnor UO_2300 (O_2300,N_29881,N_29956);
nor UO_2301 (O_2301,N_29902,N_29853);
or UO_2302 (O_2302,N_29973,N_29847);
or UO_2303 (O_2303,N_29567,N_29559);
and UO_2304 (O_2304,N_29752,N_29950);
xor UO_2305 (O_2305,N_29506,N_29939);
nor UO_2306 (O_2306,N_29814,N_29553);
and UO_2307 (O_2307,N_29679,N_29829);
xnor UO_2308 (O_2308,N_29541,N_29663);
xnor UO_2309 (O_2309,N_29830,N_29529);
and UO_2310 (O_2310,N_29656,N_29751);
or UO_2311 (O_2311,N_29957,N_29617);
nor UO_2312 (O_2312,N_29650,N_29957);
nor UO_2313 (O_2313,N_29613,N_29752);
or UO_2314 (O_2314,N_29649,N_29721);
xor UO_2315 (O_2315,N_29657,N_29717);
xnor UO_2316 (O_2316,N_29759,N_29783);
and UO_2317 (O_2317,N_29783,N_29656);
and UO_2318 (O_2318,N_29671,N_29636);
xor UO_2319 (O_2319,N_29565,N_29764);
nor UO_2320 (O_2320,N_29796,N_29818);
nand UO_2321 (O_2321,N_29892,N_29778);
nor UO_2322 (O_2322,N_29905,N_29705);
or UO_2323 (O_2323,N_29647,N_29783);
or UO_2324 (O_2324,N_29663,N_29691);
nand UO_2325 (O_2325,N_29860,N_29629);
nor UO_2326 (O_2326,N_29821,N_29834);
nor UO_2327 (O_2327,N_29535,N_29842);
xor UO_2328 (O_2328,N_29977,N_29714);
and UO_2329 (O_2329,N_29811,N_29612);
nor UO_2330 (O_2330,N_29962,N_29619);
nand UO_2331 (O_2331,N_29623,N_29619);
nand UO_2332 (O_2332,N_29722,N_29594);
nor UO_2333 (O_2333,N_29784,N_29608);
xnor UO_2334 (O_2334,N_29976,N_29875);
and UO_2335 (O_2335,N_29995,N_29906);
or UO_2336 (O_2336,N_29976,N_29650);
nor UO_2337 (O_2337,N_29603,N_29946);
nand UO_2338 (O_2338,N_29849,N_29710);
nor UO_2339 (O_2339,N_29626,N_29629);
nor UO_2340 (O_2340,N_29777,N_29879);
or UO_2341 (O_2341,N_29804,N_29591);
nand UO_2342 (O_2342,N_29547,N_29679);
or UO_2343 (O_2343,N_29735,N_29761);
or UO_2344 (O_2344,N_29646,N_29557);
nand UO_2345 (O_2345,N_29667,N_29663);
or UO_2346 (O_2346,N_29525,N_29869);
and UO_2347 (O_2347,N_29619,N_29981);
nor UO_2348 (O_2348,N_29613,N_29981);
and UO_2349 (O_2349,N_29806,N_29745);
xor UO_2350 (O_2350,N_29625,N_29612);
xnor UO_2351 (O_2351,N_29969,N_29691);
xnor UO_2352 (O_2352,N_29981,N_29501);
nor UO_2353 (O_2353,N_29972,N_29919);
and UO_2354 (O_2354,N_29622,N_29514);
and UO_2355 (O_2355,N_29584,N_29823);
nand UO_2356 (O_2356,N_29632,N_29951);
and UO_2357 (O_2357,N_29912,N_29577);
xnor UO_2358 (O_2358,N_29759,N_29746);
nor UO_2359 (O_2359,N_29811,N_29800);
and UO_2360 (O_2360,N_29532,N_29531);
or UO_2361 (O_2361,N_29807,N_29946);
and UO_2362 (O_2362,N_29716,N_29818);
or UO_2363 (O_2363,N_29638,N_29819);
nor UO_2364 (O_2364,N_29664,N_29844);
nand UO_2365 (O_2365,N_29751,N_29564);
nor UO_2366 (O_2366,N_29797,N_29760);
nor UO_2367 (O_2367,N_29782,N_29913);
nor UO_2368 (O_2368,N_29773,N_29510);
and UO_2369 (O_2369,N_29903,N_29925);
or UO_2370 (O_2370,N_29933,N_29948);
xnor UO_2371 (O_2371,N_29563,N_29501);
nor UO_2372 (O_2372,N_29711,N_29862);
nor UO_2373 (O_2373,N_29882,N_29883);
and UO_2374 (O_2374,N_29843,N_29850);
and UO_2375 (O_2375,N_29508,N_29687);
xor UO_2376 (O_2376,N_29699,N_29548);
nor UO_2377 (O_2377,N_29781,N_29517);
nand UO_2378 (O_2378,N_29719,N_29958);
or UO_2379 (O_2379,N_29625,N_29637);
and UO_2380 (O_2380,N_29707,N_29564);
xnor UO_2381 (O_2381,N_29607,N_29660);
xnor UO_2382 (O_2382,N_29798,N_29960);
and UO_2383 (O_2383,N_29510,N_29634);
or UO_2384 (O_2384,N_29691,N_29503);
and UO_2385 (O_2385,N_29557,N_29869);
xor UO_2386 (O_2386,N_29584,N_29949);
or UO_2387 (O_2387,N_29616,N_29502);
nor UO_2388 (O_2388,N_29904,N_29910);
xor UO_2389 (O_2389,N_29561,N_29829);
and UO_2390 (O_2390,N_29826,N_29853);
or UO_2391 (O_2391,N_29764,N_29847);
nor UO_2392 (O_2392,N_29682,N_29715);
or UO_2393 (O_2393,N_29623,N_29708);
nor UO_2394 (O_2394,N_29881,N_29597);
nor UO_2395 (O_2395,N_29597,N_29708);
or UO_2396 (O_2396,N_29577,N_29772);
or UO_2397 (O_2397,N_29823,N_29610);
xor UO_2398 (O_2398,N_29929,N_29633);
nand UO_2399 (O_2399,N_29634,N_29939);
nand UO_2400 (O_2400,N_29620,N_29889);
xnor UO_2401 (O_2401,N_29636,N_29549);
xnor UO_2402 (O_2402,N_29975,N_29658);
or UO_2403 (O_2403,N_29580,N_29740);
or UO_2404 (O_2404,N_29857,N_29679);
nor UO_2405 (O_2405,N_29550,N_29796);
xnor UO_2406 (O_2406,N_29876,N_29700);
nand UO_2407 (O_2407,N_29884,N_29840);
xnor UO_2408 (O_2408,N_29605,N_29609);
nor UO_2409 (O_2409,N_29530,N_29886);
and UO_2410 (O_2410,N_29573,N_29886);
xor UO_2411 (O_2411,N_29631,N_29726);
nor UO_2412 (O_2412,N_29599,N_29768);
xor UO_2413 (O_2413,N_29960,N_29968);
or UO_2414 (O_2414,N_29721,N_29870);
and UO_2415 (O_2415,N_29991,N_29864);
xor UO_2416 (O_2416,N_29799,N_29909);
xnor UO_2417 (O_2417,N_29629,N_29843);
or UO_2418 (O_2418,N_29685,N_29944);
xor UO_2419 (O_2419,N_29616,N_29883);
xnor UO_2420 (O_2420,N_29657,N_29943);
nor UO_2421 (O_2421,N_29921,N_29769);
or UO_2422 (O_2422,N_29532,N_29833);
nor UO_2423 (O_2423,N_29614,N_29996);
nor UO_2424 (O_2424,N_29504,N_29612);
nor UO_2425 (O_2425,N_29511,N_29556);
and UO_2426 (O_2426,N_29595,N_29788);
and UO_2427 (O_2427,N_29584,N_29746);
xnor UO_2428 (O_2428,N_29702,N_29875);
nand UO_2429 (O_2429,N_29960,N_29928);
nor UO_2430 (O_2430,N_29593,N_29735);
nor UO_2431 (O_2431,N_29586,N_29511);
nand UO_2432 (O_2432,N_29726,N_29683);
or UO_2433 (O_2433,N_29519,N_29966);
nand UO_2434 (O_2434,N_29591,N_29924);
xnor UO_2435 (O_2435,N_29738,N_29785);
nor UO_2436 (O_2436,N_29847,N_29884);
nor UO_2437 (O_2437,N_29965,N_29792);
nor UO_2438 (O_2438,N_29916,N_29820);
nand UO_2439 (O_2439,N_29541,N_29695);
xor UO_2440 (O_2440,N_29970,N_29550);
nand UO_2441 (O_2441,N_29646,N_29899);
or UO_2442 (O_2442,N_29770,N_29951);
nor UO_2443 (O_2443,N_29672,N_29785);
or UO_2444 (O_2444,N_29986,N_29800);
and UO_2445 (O_2445,N_29867,N_29802);
or UO_2446 (O_2446,N_29956,N_29761);
or UO_2447 (O_2447,N_29743,N_29806);
xnor UO_2448 (O_2448,N_29524,N_29729);
and UO_2449 (O_2449,N_29805,N_29723);
nand UO_2450 (O_2450,N_29972,N_29710);
xor UO_2451 (O_2451,N_29582,N_29533);
or UO_2452 (O_2452,N_29959,N_29692);
nor UO_2453 (O_2453,N_29638,N_29782);
xor UO_2454 (O_2454,N_29825,N_29629);
or UO_2455 (O_2455,N_29598,N_29638);
nand UO_2456 (O_2456,N_29692,N_29678);
nand UO_2457 (O_2457,N_29756,N_29853);
or UO_2458 (O_2458,N_29583,N_29868);
or UO_2459 (O_2459,N_29937,N_29906);
xor UO_2460 (O_2460,N_29704,N_29792);
nor UO_2461 (O_2461,N_29641,N_29683);
nor UO_2462 (O_2462,N_29942,N_29936);
nand UO_2463 (O_2463,N_29516,N_29668);
xor UO_2464 (O_2464,N_29894,N_29915);
and UO_2465 (O_2465,N_29707,N_29508);
nor UO_2466 (O_2466,N_29941,N_29715);
nor UO_2467 (O_2467,N_29840,N_29848);
and UO_2468 (O_2468,N_29758,N_29745);
xor UO_2469 (O_2469,N_29722,N_29571);
nand UO_2470 (O_2470,N_29714,N_29896);
and UO_2471 (O_2471,N_29591,N_29893);
and UO_2472 (O_2472,N_29931,N_29879);
nand UO_2473 (O_2473,N_29809,N_29660);
or UO_2474 (O_2474,N_29657,N_29731);
and UO_2475 (O_2475,N_29734,N_29821);
nand UO_2476 (O_2476,N_29719,N_29655);
and UO_2477 (O_2477,N_29991,N_29842);
or UO_2478 (O_2478,N_29601,N_29777);
or UO_2479 (O_2479,N_29856,N_29789);
or UO_2480 (O_2480,N_29867,N_29845);
nand UO_2481 (O_2481,N_29578,N_29743);
or UO_2482 (O_2482,N_29918,N_29773);
xor UO_2483 (O_2483,N_29565,N_29550);
and UO_2484 (O_2484,N_29545,N_29881);
and UO_2485 (O_2485,N_29823,N_29701);
and UO_2486 (O_2486,N_29732,N_29643);
and UO_2487 (O_2487,N_29661,N_29526);
or UO_2488 (O_2488,N_29725,N_29881);
or UO_2489 (O_2489,N_29668,N_29684);
nand UO_2490 (O_2490,N_29577,N_29813);
nor UO_2491 (O_2491,N_29758,N_29709);
nand UO_2492 (O_2492,N_29542,N_29883);
nor UO_2493 (O_2493,N_29623,N_29525);
xnor UO_2494 (O_2494,N_29539,N_29954);
and UO_2495 (O_2495,N_29949,N_29687);
or UO_2496 (O_2496,N_29763,N_29532);
nand UO_2497 (O_2497,N_29530,N_29671);
or UO_2498 (O_2498,N_29715,N_29979);
nand UO_2499 (O_2499,N_29965,N_29779);
xor UO_2500 (O_2500,N_29611,N_29529);
xor UO_2501 (O_2501,N_29540,N_29649);
nand UO_2502 (O_2502,N_29960,N_29916);
xor UO_2503 (O_2503,N_29611,N_29522);
nand UO_2504 (O_2504,N_29668,N_29669);
and UO_2505 (O_2505,N_29893,N_29551);
xnor UO_2506 (O_2506,N_29531,N_29548);
nand UO_2507 (O_2507,N_29964,N_29545);
nor UO_2508 (O_2508,N_29980,N_29695);
xnor UO_2509 (O_2509,N_29770,N_29615);
xnor UO_2510 (O_2510,N_29695,N_29790);
nand UO_2511 (O_2511,N_29794,N_29977);
nor UO_2512 (O_2512,N_29867,N_29554);
and UO_2513 (O_2513,N_29784,N_29522);
nor UO_2514 (O_2514,N_29813,N_29635);
nand UO_2515 (O_2515,N_29883,N_29863);
nor UO_2516 (O_2516,N_29866,N_29764);
and UO_2517 (O_2517,N_29769,N_29578);
nand UO_2518 (O_2518,N_29919,N_29912);
xor UO_2519 (O_2519,N_29550,N_29760);
nand UO_2520 (O_2520,N_29931,N_29527);
nand UO_2521 (O_2521,N_29631,N_29823);
and UO_2522 (O_2522,N_29620,N_29934);
nand UO_2523 (O_2523,N_29817,N_29786);
xnor UO_2524 (O_2524,N_29833,N_29762);
nor UO_2525 (O_2525,N_29578,N_29883);
nor UO_2526 (O_2526,N_29853,N_29729);
nor UO_2527 (O_2527,N_29989,N_29509);
or UO_2528 (O_2528,N_29512,N_29741);
nor UO_2529 (O_2529,N_29700,N_29705);
and UO_2530 (O_2530,N_29913,N_29974);
and UO_2531 (O_2531,N_29884,N_29694);
nor UO_2532 (O_2532,N_29661,N_29628);
xnor UO_2533 (O_2533,N_29609,N_29630);
or UO_2534 (O_2534,N_29529,N_29923);
or UO_2535 (O_2535,N_29506,N_29863);
or UO_2536 (O_2536,N_29716,N_29764);
xnor UO_2537 (O_2537,N_29937,N_29568);
nand UO_2538 (O_2538,N_29577,N_29902);
or UO_2539 (O_2539,N_29577,N_29808);
nor UO_2540 (O_2540,N_29525,N_29867);
nor UO_2541 (O_2541,N_29854,N_29817);
xnor UO_2542 (O_2542,N_29798,N_29992);
nor UO_2543 (O_2543,N_29615,N_29879);
nor UO_2544 (O_2544,N_29859,N_29746);
nor UO_2545 (O_2545,N_29526,N_29603);
nor UO_2546 (O_2546,N_29810,N_29769);
or UO_2547 (O_2547,N_29853,N_29752);
xor UO_2548 (O_2548,N_29679,N_29735);
nor UO_2549 (O_2549,N_29570,N_29711);
nand UO_2550 (O_2550,N_29501,N_29917);
or UO_2551 (O_2551,N_29906,N_29917);
nor UO_2552 (O_2552,N_29678,N_29792);
nor UO_2553 (O_2553,N_29649,N_29833);
nand UO_2554 (O_2554,N_29960,N_29945);
xnor UO_2555 (O_2555,N_29504,N_29940);
nand UO_2556 (O_2556,N_29526,N_29776);
nand UO_2557 (O_2557,N_29865,N_29950);
xor UO_2558 (O_2558,N_29596,N_29814);
or UO_2559 (O_2559,N_29541,N_29605);
and UO_2560 (O_2560,N_29574,N_29531);
nor UO_2561 (O_2561,N_29989,N_29558);
or UO_2562 (O_2562,N_29523,N_29963);
and UO_2563 (O_2563,N_29907,N_29935);
xor UO_2564 (O_2564,N_29837,N_29836);
and UO_2565 (O_2565,N_29809,N_29758);
xor UO_2566 (O_2566,N_29840,N_29501);
or UO_2567 (O_2567,N_29990,N_29891);
nor UO_2568 (O_2568,N_29502,N_29583);
or UO_2569 (O_2569,N_29525,N_29912);
xnor UO_2570 (O_2570,N_29793,N_29980);
xor UO_2571 (O_2571,N_29725,N_29686);
and UO_2572 (O_2572,N_29742,N_29763);
nand UO_2573 (O_2573,N_29612,N_29896);
xnor UO_2574 (O_2574,N_29761,N_29535);
nand UO_2575 (O_2575,N_29854,N_29872);
and UO_2576 (O_2576,N_29974,N_29665);
nor UO_2577 (O_2577,N_29772,N_29556);
nand UO_2578 (O_2578,N_29531,N_29514);
xnor UO_2579 (O_2579,N_29913,N_29907);
or UO_2580 (O_2580,N_29792,N_29786);
xnor UO_2581 (O_2581,N_29835,N_29598);
or UO_2582 (O_2582,N_29930,N_29518);
or UO_2583 (O_2583,N_29620,N_29685);
xnor UO_2584 (O_2584,N_29645,N_29614);
and UO_2585 (O_2585,N_29988,N_29873);
xnor UO_2586 (O_2586,N_29876,N_29787);
nor UO_2587 (O_2587,N_29519,N_29940);
nor UO_2588 (O_2588,N_29684,N_29612);
nand UO_2589 (O_2589,N_29743,N_29828);
nand UO_2590 (O_2590,N_29613,N_29530);
nand UO_2591 (O_2591,N_29647,N_29579);
nand UO_2592 (O_2592,N_29573,N_29698);
nor UO_2593 (O_2593,N_29711,N_29500);
or UO_2594 (O_2594,N_29529,N_29594);
nor UO_2595 (O_2595,N_29951,N_29713);
nor UO_2596 (O_2596,N_29508,N_29617);
nand UO_2597 (O_2597,N_29883,N_29872);
nand UO_2598 (O_2598,N_29540,N_29851);
or UO_2599 (O_2599,N_29761,N_29616);
nor UO_2600 (O_2600,N_29672,N_29798);
xnor UO_2601 (O_2601,N_29707,N_29985);
xnor UO_2602 (O_2602,N_29801,N_29574);
and UO_2603 (O_2603,N_29849,N_29731);
nand UO_2604 (O_2604,N_29752,N_29662);
or UO_2605 (O_2605,N_29588,N_29809);
and UO_2606 (O_2606,N_29539,N_29559);
xor UO_2607 (O_2607,N_29761,N_29868);
nor UO_2608 (O_2608,N_29886,N_29838);
xor UO_2609 (O_2609,N_29978,N_29587);
xor UO_2610 (O_2610,N_29939,N_29732);
or UO_2611 (O_2611,N_29903,N_29652);
or UO_2612 (O_2612,N_29793,N_29524);
and UO_2613 (O_2613,N_29943,N_29826);
nand UO_2614 (O_2614,N_29870,N_29808);
nor UO_2615 (O_2615,N_29993,N_29523);
nor UO_2616 (O_2616,N_29785,N_29947);
xor UO_2617 (O_2617,N_29597,N_29868);
and UO_2618 (O_2618,N_29928,N_29796);
nand UO_2619 (O_2619,N_29802,N_29714);
nor UO_2620 (O_2620,N_29800,N_29863);
nand UO_2621 (O_2621,N_29789,N_29981);
nor UO_2622 (O_2622,N_29757,N_29500);
or UO_2623 (O_2623,N_29699,N_29562);
nor UO_2624 (O_2624,N_29619,N_29781);
nand UO_2625 (O_2625,N_29660,N_29588);
and UO_2626 (O_2626,N_29896,N_29584);
and UO_2627 (O_2627,N_29987,N_29761);
nor UO_2628 (O_2628,N_29572,N_29888);
or UO_2629 (O_2629,N_29677,N_29972);
or UO_2630 (O_2630,N_29632,N_29560);
nor UO_2631 (O_2631,N_29679,N_29902);
xnor UO_2632 (O_2632,N_29789,N_29674);
and UO_2633 (O_2633,N_29704,N_29860);
nand UO_2634 (O_2634,N_29918,N_29618);
xnor UO_2635 (O_2635,N_29829,N_29960);
xor UO_2636 (O_2636,N_29506,N_29588);
nand UO_2637 (O_2637,N_29738,N_29732);
and UO_2638 (O_2638,N_29787,N_29968);
nand UO_2639 (O_2639,N_29832,N_29896);
nand UO_2640 (O_2640,N_29861,N_29998);
nor UO_2641 (O_2641,N_29662,N_29798);
xor UO_2642 (O_2642,N_29538,N_29790);
nand UO_2643 (O_2643,N_29523,N_29930);
nand UO_2644 (O_2644,N_29573,N_29980);
or UO_2645 (O_2645,N_29665,N_29667);
xor UO_2646 (O_2646,N_29722,N_29627);
and UO_2647 (O_2647,N_29758,N_29666);
nor UO_2648 (O_2648,N_29917,N_29824);
nand UO_2649 (O_2649,N_29946,N_29613);
xnor UO_2650 (O_2650,N_29722,N_29878);
xnor UO_2651 (O_2651,N_29864,N_29878);
nand UO_2652 (O_2652,N_29865,N_29818);
or UO_2653 (O_2653,N_29750,N_29574);
and UO_2654 (O_2654,N_29841,N_29728);
nand UO_2655 (O_2655,N_29591,N_29679);
or UO_2656 (O_2656,N_29855,N_29556);
nand UO_2657 (O_2657,N_29619,N_29784);
and UO_2658 (O_2658,N_29814,N_29917);
xnor UO_2659 (O_2659,N_29775,N_29877);
and UO_2660 (O_2660,N_29652,N_29886);
xor UO_2661 (O_2661,N_29697,N_29820);
and UO_2662 (O_2662,N_29634,N_29521);
nand UO_2663 (O_2663,N_29928,N_29638);
or UO_2664 (O_2664,N_29849,N_29827);
nor UO_2665 (O_2665,N_29586,N_29925);
and UO_2666 (O_2666,N_29827,N_29664);
or UO_2667 (O_2667,N_29590,N_29700);
or UO_2668 (O_2668,N_29683,N_29800);
and UO_2669 (O_2669,N_29723,N_29536);
nand UO_2670 (O_2670,N_29977,N_29934);
and UO_2671 (O_2671,N_29680,N_29672);
nor UO_2672 (O_2672,N_29689,N_29967);
and UO_2673 (O_2673,N_29894,N_29889);
and UO_2674 (O_2674,N_29751,N_29589);
and UO_2675 (O_2675,N_29803,N_29546);
nand UO_2676 (O_2676,N_29896,N_29683);
nand UO_2677 (O_2677,N_29669,N_29991);
nand UO_2678 (O_2678,N_29785,N_29562);
nand UO_2679 (O_2679,N_29803,N_29964);
or UO_2680 (O_2680,N_29626,N_29952);
or UO_2681 (O_2681,N_29724,N_29767);
or UO_2682 (O_2682,N_29938,N_29878);
and UO_2683 (O_2683,N_29902,N_29869);
xor UO_2684 (O_2684,N_29861,N_29578);
nor UO_2685 (O_2685,N_29991,N_29971);
and UO_2686 (O_2686,N_29565,N_29698);
or UO_2687 (O_2687,N_29693,N_29842);
and UO_2688 (O_2688,N_29975,N_29885);
nor UO_2689 (O_2689,N_29923,N_29606);
xor UO_2690 (O_2690,N_29796,N_29540);
or UO_2691 (O_2691,N_29682,N_29642);
or UO_2692 (O_2692,N_29588,N_29616);
nand UO_2693 (O_2693,N_29966,N_29504);
nor UO_2694 (O_2694,N_29663,N_29811);
or UO_2695 (O_2695,N_29766,N_29692);
nand UO_2696 (O_2696,N_29926,N_29988);
nand UO_2697 (O_2697,N_29590,N_29874);
and UO_2698 (O_2698,N_29700,N_29568);
xnor UO_2699 (O_2699,N_29579,N_29767);
nor UO_2700 (O_2700,N_29743,N_29869);
and UO_2701 (O_2701,N_29521,N_29724);
or UO_2702 (O_2702,N_29792,N_29770);
nor UO_2703 (O_2703,N_29985,N_29816);
nor UO_2704 (O_2704,N_29679,N_29737);
nor UO_2705 (O_2705,N_29786,N_29708);
nand UO_2706 (O_2706,N_29761,N_29873);
nor UO_2707 (O_2707,N_29677,N_29572);
nor UO_2708 (O_2708,N_29741,N_29724);
and UO_2709 (O_2709,N_29911,N_29546);
or UO_2710 (O_2710,N_29659,N_29756);
xor UO_2711 (O_2711,N_29871,N_29806);
nand UO_2712 (O_2712,N_29711,N_29710);
and UO_2713 (O_2713,N_29697,N_29683);
or UO_2714 (O_2714,N_29624,N_29799);
nor UO_2715 (O_2715,N_29550,N_29554);
nor UO_2716 (O_2716,N_29922,N_29880);
xnor UO_2717 (O_2717,N_29704,N_29776);
or UO_2718 (O_2718,N_29943,N_29603);
xnor UO_2719 (O_2719,N_29544,N_29567);
and UO_2720 (O_2720,N_29583,N_29931);
nand UO_2721 (O_2721,N_29870,N_29851);
and UO_2722 (O_2722,N_29944,N_29666);
or UO_2723 (O_2723,N_29592,N_29529);
or UO_2724 (O_2724,N_29689,N_29544);
xnor UO_2725 (O_2725,N_29949,N_29677);
and UO_2726 (O_2726,N_29501,N_29809);
nand UO_2727 (O_2727,N_29805,N_29720);
and UO_2728 (O_2728,N_29874,N_29974);
and UO_2729 (O_2729,N_29735,N_29512);
or UO_2730 (O_2730,N_29666,N_29719);
xnor UO_2731 (O_2731,N_29630,N_29500);
nand UO_2732 (O_2732,N_29878,N_29793);
and UO_2733 (O_2733,N_29991,N_29809);
xor UO_2734 (O_2734,N_29889,N_29869);
nor UO_2735 (O_2735,N_29907,N_29992);
or UO_2736 (O_2736,N_29544,N_29909);
and UO_2737 (O_2737,N_29689,N_29589);
xnor UO_2738 (O_2738,N_29736,N_29683);
nor UO_2739 (O_2739,N_29862,N_29534);
and UO_2740 (O_2740,N_29826,N_29664);
xnor UO_2741 (O_2741,N_29993,N_29814);
and UO_2742 (O_2742,N_29797,N_29999);
or UO_2743 (O_2743,N_29515,N_29893);
nor UO_2744 (O_2744,N_29981,N_29717);
xnor UO_2745 (O_2745,N_29621,N_29753);
or UO_2746 (O_2746,N_29582,N_29971);
xor UO_2747 (O_2747,N_29810,N_29640);
nor UO_2748 (O_2748,N_29850,N_29515);
and UO_2749 (O_2749,N_29550,N_29653);
and UO_2750 (O_2750,N_29975,N_29700);
nor UO_2751 (O_2751,N_29838,N_29765);
or UO_2752 (O_2752,N_29936,N_29866);
nor UO_2753 (O_2753,N_29732,N_29681);
or UO_2754 (O_2754,N_29600,N_29750);
nand UO_2755 (O_2755,N_29860,N_29512);
nand UO_2756 (O_2756,N_29842,N_29879);
nand UO_2757 (O_2757,N_29767,N_29600);
xnor UO_2758 (O_2758,N_29612,N_29819);
nand UO_2759 (O_2759,N_29945,N_29568);
nand UO_2760 (O_2760,N_29819,N_29703);
nand UO_2761 (O_2761,N_29795,N_29653);
xor UO_2762 (O_2762,N_29624,N_29566);
or UO_2763 (O_2763,N_29918,N_29595);
or UO_2764 (O_2764,N_29817,N_29890);
nand UO_2765 (O_2765,N_29633,N_29802);
and UO_2766 (O_2766,N_29541,N_29866);
and UO_2767 (O_2767,N_29852,N_29897);
and UO_2768 (O_2768,N_29597,N_29689);
or UO_2769 (O_2769,N_29592,N_29827);
or UO_2770 (O_2770,N_29622,N_29922);
and UO_2771 (O_2771,N_29805,N_29552);
nor UO_2772 (O_2772,N_29795,N_29885);
xor UO_2773 (O_2773,N_29522,N_29994);
xor UO_2774 (O_2774,N_29887,N_29548);
nand UO_2775 (O_2775,N_29666,N_29578);
nor UO_2776 (O_2776,N_29712,N_29993);
nand UO_2777 (O_2777,N_29832,N_29537);
and UO_2778 (O_2778,N_29570,N_29509);
nand UO_2779 (O_2779,N_29971,N_29610);
nand UO_2780 (O_2780,N_29750,N_29586);
nand UO_2781 (O_2781,N_29884,N_29842);
xnor UO_2782 (O_2782,N_29638,N_29551);
nand UO_2783 (O_2783,N_29870,N_29702);
nor UO_2784 (O_2784,N_29841,N_29591);
nor UO_2785 (O_2785,N_29546,N_29952);
xor UO_2786 (O_2786,N_29664,N_29529);
nand UO_2787 (O_2787,N_29652,N_29781);
nor UO_2788 (O_2788,N_29740,N_29697);
and UO_2789 (O_2789,N_29868,N_29612);
nor UO_2790 (O_2790,N_29715,N_29974);
xor UO_2791 (O_2791,N_29591,N_29852);
and UO_2792 (O_2792,N_29859,N_29819);
xnor UO_2793 (O_2793,N_29725,N_29549);
nor UO_2794 (O_2794,N_29541,N_29750);
nand UO_2795 (O_2795,N_29848,N_29628);
xor UO_2796 (O_2796,N_29502,N_29585);
xnor UO_2797 (O_2797,N_29574,N_29984);
nor UO_2798 (O_2798,N_29704,N_29798);
and UO_2799 (O_2799,N_29670,N_29714);
xnor UO_2800 (O_2800,N_29511,N_29585);
or UO_2801 (O_2801,N_29914,N_29669);
nand UO_2802 (O_2802,N_29646,N_29593);
nand UO_2803 (O_2803,N_29679,N_29976);
xnor UO_2804 (O_2804,N_29532,N_29674);
or UO_2805 (O_2805,N_29978,N_29620);
nor UO_2806 (O_2806,N_29860,N_29998);
nand UO_2807 (O_2807,N_29882,N_29922);
nor UO_2808 (O_2808,N_29633,N_29501);
and UO_2809 (O_2809,N_29710,N_29921);
xnor UO_2810 (O_2810,N_29896,N_29707);
nand UO_2811 (O_2811,N_29739,N_29904);
and UO_2812 (O_2812,N_29540,N_29656);
nor UO_2813 (O_2813,N_29815,N_29835);
nor UO_2814 (O_2814,N_29809,N_29725);
nor UO_2815 (O_2815,N_29912,N_29994);
or UO_2816 (O_2816,N_29732,N_29985);
nor UO_2817 (O_2817,N_29917,N_29510);
nand UO_2818 (O_2818,N_29639,N_29606);
or UO_2819 (O_2819,N_29772,N_29989);
or UO_2820 (O_2820,N_29611,N_29706);
nand UO_2821 (O_2821,N_29843,N_29890);
nor UO_2822 (O_2822,N_29836,N_29770);
or UO_2823 (O_2823,N_29876,N_29747);
and UO_2824 (O_2824,N_29661,N_29675);
and UO_2825 (O_2825,N_29516,N_29903);
xnor UO_2826 (O_2826,N_29772,N_29838);
and UO_2827 (O_2827,N_29626,N_29787);
nand UO_2828 (O_2828,N_29656,N_29533);
nor UO_2829 (O_2829,N_29985,N_29742);
nand UO_2830 (O_2830,N_29533,N_29747);
or UO_2831 (O_2831,N_29800,N_29806);
nand UO_2832 (O_2832,N_29773,N_29606);
or UO_2833 (O_2833,N_29806,N_29972);
and UO_2834 (O_2834,N_29953,N_29978);
nor UO_2835 (O_2835,N_29993,N_29597);
nand UO_2836 (O_2836,N_29993,N_29770);
nand UO_2837 (O_2837,N_29538,N_29760);
nor UO_2838 (O_2838,N_29886,N_29671);
xor UO_2839 (O_2839,N_29737,N_29636);
or UO_2840 (O_2840,N_29676,N_29542);
nor UO_2841 (O_2841,N_29926,N_29776);
or UO_2842 (O_2842,N_29729,N_29962);
xnor UO_2843 (O_2843,N_29737,N_29710);
and UO_2844 (O_2844,N_29780,N_29625);
nand UO_2845 (O_2845,N_29920,N_29978);
or UO_2846 (O_2846,N_29578,N_29622);
or UO_2847 (O_2847,N_29650,N_29731);
xor UO_2848 (O_2848,N_29641,N_29866);
xnor UO_2849 (O_2849,N_29800,N_29626);
or UO_2850 (O_2850,N_29730,N_29656);
or UO_2851 (O_2851,N_29642,N_29836);
nand UO_2852 (O_2852,N_29928,N_29883);
xor UO_2853 (O_2853,N_29662,N_29594);
and UO_2854 (O_2854,N_29602,N_29790);
nand UO_2855 (O_2855,N_29697,N_29806);
or UO_2856 (O_2856,N_29956,N_29807);
xnor UO_2857 (O_2857,N_29740,N_29950);
and UO_2858 (O_2858,N_29598,N_29761);
or UO_2859 (O_2859,N_29562,N_29556);
nand UO_2860 (O_2860,N_29602,N_29828);
xnor UO_2861 (O_2861,N_29546,N_29897);
xor UO_2862 (O_2862,N_29853,N_29734);
nand UO_2863 (O_2863,N_29780,N_29712);
nand UO_2864 (O_2864,N_29911,N_29815);
nand UO_2865 (O_2865,N_29902,N_29586);
nand UO_2866 (O_2866,N_29829,N_29948);
xnor UO_2867 (O_2867,N_29715,N_29656);
nor UO_2868 (O_2868,N_29753,N_29751);
nor UO_2869 (O_2869,N_29754,N_29771);
xnor UO_2870 (O_2870,N_29667,N_29793);
xor UO_2871 (O_2871,N_29934,N_29502);
or UO_2872 (O_2872,N_29609,N_29606);
and UO_2873 (O_2873,N_29801,N_29734);
nor UO_2874 (O_2874,N_29538,N_29691);
or UO_2875 (O_2875,N_29880,N_29501);
and UO_2876 (O_2876,N_29640,N_29564);
or UO_2877 (O_2877,N_29982,N_29813);
nand UO_2878 (O_2878,N_29969,N_29590);
and UO_2879 (O_2879,N_29999,N_29831);
nand UO_2880 (O_2880,N_29900,N_29964);
and UO_2881 (O_2881,N_29974,N_29812);
or UO_2882 (O_2882,N_29887,N_29816);
nor UO_2883 (O_2883,N_29982,N_29909);
and UO_2884 (O_2884,N_29723,N_29695);
and UO_2885 (O_2885,N_29599,N_29869);
xor UO_2886 (O_2886,N_29774,N_29704);
nand UO_2887 (O_2887,N_29674,N_29764);
nand UO_2888 (O_2888,N_29843,N_29986);
and UO_2889 (O_2889,N_29673,N_29590);
nand UO_2890 (O_2890,N_29615,N_29631);
nor UO_2891 (O_2891,N_29949,N_29899);
nor UO_2892 (O_2892,N_29787,N_29691);
nand UO_2893 (O_2893,N_29675,N_29736);
nand UO_2894 (O_2894,N_29509,N_29969);
nor UO_2895 (O_2895,N_29601,N_29749);
nor UO_2896 (O_2896,N_29893,N_29901);
xor UO_2897 (O_2897,N_29542,N_29869);
nand UO_2898 (O_2898,N_29667,N_29756);
nor UO_2899 (O_2899,N_29924,N_29822);
or UO_2900 (O_2900,N_29571,N_29758);
nor UO_2901 (O_2901,N_29799,N_29873);
xor UO_2902 (O_2902,N_29999,N_29826);
nand UO_2903 (O_2903,N_29813,N_29778);
xor UO_2904 (O_2904,N_29566,N_29776);
and UO_2905 (O_2905,N_29743,N_29596);
or UO_2906 (O_2906,N_29835,N_29748);
xnor UO_2907 (O_2907,N_29860,N_29983);
and UO_2908 (O_2908,N_29875,N_29879);
or UO_2909 (O_2909,N_29954,N_29594);
and UO_2910 (O_2910,N_29515,N_29723);
nor UO_2911 (O_2911,N_29552,N_29933);
nand UO_2912 (O_2912,N_29701,N_29568);
nor UO_2913 (O_2913,N_29906,N_29776);
and UO_2914 (O_2914,N_29552,N_29611);
xor UO_2915 (O_2915,N_29912,N_29674);
nand UO_2916 (O_2916,N_29918,N_29555);
nand UO_2917 (O_2917,N_29770,N_29992);
nor UO_2918 (O_2918,N_29836,N_29524);
xor UO_2919 (O_2919,N_29843,N_29941);
xnor UO_2920 (O_2920,N_29953,N_29938);
nand UO_2921 (O_2921,N_29548,N_29811);
nor UO_2922 (O_2922,N_29926,N_29518);
nor UO_2923 (O_2923,N_29615,N_29818);
nor UO_2924 (O_2924,N_29963,N_29907);
nand UO_2925 (O_2925,N_29655,N_29652);
xor UO_2926 (O_2926,N_29898,N_29709);
xor UO_2927 (O_2927,N_29643,N_29594);
nand UO_2928 (O_2928,N_29991,N_29516);
and UO_2929 (O_2929,N_29584,N_29572);
xor UO_2930 (O_2930,N_29649,N_29514);
and UO_2931 (O_2931,N_29606,N_29900);
nor UO_2932 (O_2932,N_29889,N_29985);
nor UO_2933 (O_2933,N_29522,N_29837);
and UO_2934 (O_2934,N_29723,N_29954);
xor UO_2935 (O_2935,N_29846,N_29603);
or UO_2936 (O_2936,N_29794,N_29558);
or UO_2937 (O_2937,N_29507,N_29709);
xor UO_2938 (O_2938,N_29972,N_29701);
nand UO_2939 (O_2939,N_29948,N_29709);
nor UO_2940 (O_2940,N_29873,N_29651);
xor UO_2941 (O_2941,N_29505,N_29648);
or UO_2942 (O_2942,N_29627,N_29973);
nor UO_2943 (O_2943,N_29850,N_29753);
nand UO_2944 (O_2944,N_29857,N_29535);
and UO_2945 (O_2945,N_29960,N_29850);
and UO_2946 (O_2946,N_29605,N_29714);
or UO_2947 (O_2947,N_29522,N_29952);
and UO_2948 (O_2948,N_29953,N_29547);
nor UO_2949 (O_2949,N_29540,N_29912);
nor UO_2950 (O_2950,N_29794,N_29540);
xnor UO_2951 (O_2951,N_29933,N_29662);
nand UO_2952 (O_2952,N_29592,N_29857);
or UO_2953 (O_2953,N_29872,N_29542);
nand UO_2954 (O_2954,N_29764,N_29500);
nor UO_2955 (O_2955,N_29860,N_29973);
xor UO_2956 (O_2956,N_29719,N_29852);
nor UO_2957 (O_2957,N_29880,N_29720);
or UO_2958 (O_2958,N_29788,N_29772);
and UO_2959 (O_2959,N_29528,N_29533);
or UO_2960 (O_2960,N_29966,N_29948);
nor UO_2961 (O_2961,N_29682,N_29527);
nor UO_2962 (O_2962,N_29954,N_29934);
and UO_2963 (O_2963,N_29812,N_29633);
or UO_2964 (O_2964,N_29886,N_29617);
nor UO_2965 (O_2965,N_29731,N_29624);
and UO_2966 (O_2966,N_29670,N_29977);
nand UO_2967 (O_2967,N_29506,N_29790);
xnor UO_2968 (O_2968,N_29811,N_29913);
nand UO_2969 (O_2969,N_29806,N_29901);
and UO_2970 (O_2970,N_29665,N_29770);
or UO_2971 (O_2971,N_29688,N_29748);
and UO_2972 (O_2972,N_29644,N_29628);
and UO_2973 (O_2973,N_29913,N_29888);
nor UO_2974 (O_2974,N_29991,N_29868);
nand UO_2975 (O_2975,N_29723,N_29919);
or UO_2976 (O_2976,N_29553,N_29768);
xnor UO_2977 (O_2977,N_29756,N_29925);
xor UO_2978 (O_2978,N_29768,N_29959);
nand UO_2979 (O_2979,N_29545,N_29942);
or UO_2980 (O_2980,N_29554,N_29614);
or UO_2981 (O_2981,N_29605,N_29662);
nor UO_2982 (O_2982,N_29574,N_29714);
nand UO_2983 (O_2983,N_29976,N_29625);
xnor UO_2984 (O_2984,N_29731,N_29911);
xor UO_2985 (O_2985,N_29864,N_29736);
or UO_2986 (O_2986,N_29640,N_29874);
nor UO_2987 (O_2987,N_29790,N_29647);
nor UO_2988 (O_2988,N_29951,N_29624);
and UO_2989 (O_2989,N_29969,N_29688);
xor UO_2990 (O_2990,N_29930,N_29744);
and UO_2991 (O_2991,N_29750,N_29625);
nand UO_2992 (O_2992,N_29880,N_29636);
or UO_2993 (O_2993,N_29573,N_29849);
or UO_2994 (O_2994,N_29747,N_29788);
or UO_2995 (O_2995,N_29768,N_29852);
xor UO_2996 (O_2996,N_29820,N_29784);
nand UO_2997 (O_2997,N_29779,N_29825);
xor UO_2998 (O_2998,N_29832,N_29796);
and UO_2999 (O_2999,N_29743,N_29721);
or UO_3000 (O_3000,N_29671,N_29719);
and UO_3001 (O_3001,N_29952,N_29991);
nor UO_3002 (O_3002,N_29684,N_29831);
and UO_3003 (O_3003,N_29864,N_29868);
and UO_3004 (O_3004,N_29500,N_29717);
and UO_3005 (O_3005,N_29832,N_29620);
and UO_3006 (O_3006,N_29955,N_29506);
nor UO_3007 (O_3007,N_29861,N_29786);
nor UO_3008 (O_3008,N_29956,N_29694);
nor UO_3009 (O_3009,N_29790,N_29725);
xor UO_3010 (O_3010,N_29601,N_29785);
nor UO_3011 (O_3011,N_29688,N_29568);
and UO_3012 (O_3012,N_29983,N_29629);
or UO_3013 (O_3013,N_29871,N_29509);
nand UO_3014 (O_3014,N_29938,N_29552);
nand UO_3015 (O_3015,N_29758,N_29511);
xnor UO_3016 (O_3016,N_29614,N_29970);
xor UO_3017 (O_3017,N_29511,N_29612);
xor UO_3018 (O_3018,N_29751,N_29941);
or UO_3019 (O_3019,N_29568,N_29661);
and UO_3020 (O_3020,N_29988,N_29854);
xor UO_3021 (O_3021,N_29509,N_29855);
xnor UO_3022 (O_3022,N_29759,N_29778);
xnor UO_3023 (O_3023,N_29639,N_29514);
and UO_3024 (O_3024,N_29642,N_29514);
nor UO_3025 (O_3025,N_29604,N_29977);
or UO_3026 (O_3026,N_29763,N_29718);
xnor UO_3027 (O_3027,N_29545,N_29573);
xor UO_3028 (O_3028,N_29707,N_29804);
nand UO_3029 (O_3029,N_29964,N_29575);
nand UO_3030 (O_3030,N_29992,N_29536);
or UO_3031 (O_3031,N_29773,N_29529);
nand UO_3032 (O_3032,N_29679,N_29669);
and UO_3033 (O_3033,N_29714,N_29662);
or UO_3034 (O_3034,N_29914,N_29732);
or UO_3035 (O_3035,N_29858,N_29608);
nor UO_3036 (O_3036,N_29509,N_29765);
or UO_3037 (O_3037,N_29564,N_29654);
xor UO_3038 (O_3038,N_29838,N_29739);
and UO_3039 (O_3039,N_29865,N_29959);
nand UO_3040 (O_3040,N_29978,N_29816);
and UO_3041 (O_3041,N_29678,N_29534);
and UO_3042 (O_3042,N_29792,N_29532);
nand UO_3043 (O_3043,N_29880,N_29850);
nor UO_3044 (O_3044,N_29960,N_29799);
nand UO_3045 (O_3045,N_29846,N_29858);
and UO_3046 (O_3046,N_29645,N_29655);
xor UO_3047 (O_3047,N_29669,N_29525);
nor UO_3048 (O_3048,N_29917,N_29792);
nor UO_3049 (O_3049,N_29863,N_29788);
xnor UO_3050 (O_3050,N_29677,N_29655);
nor UO_3051 (O_3051,N_29558,N_29911);
and UO_3052 (O_3052,N_29546,N_29527);
nand UO_3053 (O_3053,N_29653,N_29655);
nand UO_3054 (O_3054,N_29800,N_29796);
nand UO_3055 (O_3055,N_29618,N_29789);
or UO_3056 (O_3056,N_29645,N_29806);
xor UO_3057 (O_3057,N_29802,N_29552);
nor UO_3058 (O_3058,N_29755,N_29641);
nand UO_3059 (O_3059,N_29906,N_29907);
nand UO_3060 (O_3060,N_29982,N_29949);
and UO_3061 (O_3061,N_29692,N_29873);
nor UO_3062 (O_3062,N_29696,N_29749);
and UO_3063 (O_3063,N_29587,N_29558);
nand UO_3064 (O_3064,N_29788,N_29633);
xor UO_3065 (O_3065,N_29711,N_29763);
nand UO_3066 (O_3066,N_29617,N_29986);
xnor UO_3067 (O_3067,N_29587,N_29538);
xnor UO_3068 (O_3068,N_29722,N_29805);
or UO_3069 (O_3069,N_29926,N_29996);
xnor UO_3070 (O_3070,N_29911,N_29985);
xor UO_3071 (O_3071,N_29937,N_29896);
xnor UO_3072 (O_3072,N_29549,N_29562);
nor UO_3073 (O_3073,N_29648,N_29789);
xor UO_3074 (O_3074,N_29721,N_29826);
or UO_3075 (O_3075,N_29728,N_29797);
xnor UO_3076 (O_3076,N_29787,N_29570);
nand UO_3077 (O_3077,N_29853,N_29929);
and UO_3078 (O_3078,N_29995,N_29754);
and UO_3079 (O_3079,N_29786,N_29721);
and UO_3080 (O_3080,N_29550,N_29651);
nor UO_3081 (O_3081,N_29513,N_29578);
nor UO_3082 (O_3082,N_29584,N_29652);
and UO_3083 (O_3083,N_29702,N_29877);
nand UO_3084 (O_3084,N_29697,N_29916);
and UO_3085 (O_3085,N_29547,N_29856);
or UO_3086 (O_3086,N_29751,N_29957);
xor UO_3087 (O_3087,N_29832,N_29831);
nand UO_3088 (O_3088,N_29793,N_29684);
nor UO_3089 (O_3089,N_29856,N_29575);
nor UO_3090 (O_3090,N_29698,N_29508);
or UO_3091 (O_3091,N_29743,N_29832);
nor UO_3092 (O_3092,N_29791,N_29890);
nor UO_3093 (O_3093,N_29643,N_29644);
or UO_3094 (O_3094,N_29897,N_29730);
nor UO_3095 (O_3095,N_29675,N_29916);
xor UO_3096 (O_3096,N_29570,N_29706);
and UO_3097 (O_3097,N_29538,N_29993);
nor UO_3098 (O_3098,N_29907,N_29945);
nor UO_3099 (O_3099,N_29996,N_29872);
nor UO_3100 (O_3100,N_29803,N_29548);
xnor UO_3101 (O_3101,N_29821,N_29732);
and UO_3102 (O_3102,N_29800,N_29656);
xnor UO_3103 (O_3103,N_29588,N_29947);
or UO_3104 (O_3104,N_29848,N_29608);
and UO_3105 (O_3105,N_29834,N_29890);
and UO_3106 (O_3106,N_29633,N_29949);
nand UO_3107 (O_3107,N_29971,N_29542);
nand UO_3108 (O_3108,N_29885,N_29617);
nand UO_3109 (O_3109,N_29896,N_29618);
xnor UO_3110 (O_3110,N_29824,N_29945);
nor UO_3111 (O_3111,N_29504,N_29795);
or UO_3112 (O_3112,N_29947,N_29646);
or UO_3113 (O_3113,N_29694,N_29958);
or UO_3114 (O_3114,N_29578,N_29791);
nand UO_3115 (O_3115,N_29640,N_29933);
nand UO_3116 (O_3116,N_29783,N_29762);
and UO_3117 (O_3117,N_29851,N_29507);
nor UO_3118 (O_3118,N_29667,N_29933);
and UO_3119 (O_3119,N_29632,N_29556);
xor UO_3120 (O_3120,N_29916,N_29650);
nand UO_3121 (O_3121,N_29829,N_29641);
and UO_3122 (O_3122,N_29936,N_29855);
xnor UO_3123 (O_3123,N_29791,N_29549);
xnor UO_3124 (O_3124,N_29808,N_29889);
nand UO_3125 (O_3125,N_29698,N_29585);
and UO_3126 (O_3126,N_29570,N_29960);
and UO_3127 (O_3127,N_29581,N_29751);
and UO_3128 (O_3128,N_29502,N_29655);
and UO_3129 (O_3129,N_29949,N_29806);
nor UO_3130 (O_3130,N_29679,N_29951);
xor UO_3131 (O_3131,N_29874,N_29939);
or UO_3132 (O_3132,N_29889,N_29659);
nand UO_3133 (O_3133,N_29894,N_29531);
xnor UO_3134 (O_3134,N_29639,N_29748);
xnor UO_3135 (O_3135,N_29711,N_29594);
xnor UO_3136 (O_3136,N_29979,N_29732);
or UO_3137 (O_3137,N_29908,N_29660);
or UO_3138 (O_3138,N_29579,N_29563);
xor UO_3139 (O_3139,N_29648,N_29835);
and UO_3140 (O_3140,N_29919,N_29921);
nand UO_3141 (O_3141,N_29976,N_29713);
or UO_3142 (O_3142,N_29663,N_29893);
or UO_3143 (O_3143,N_29646,N_29891);
xnor UO_3144 (O_3144,N_29637,N_29520);
or UO_3145 (O_3145,N_29829,N_29926);
xnor UO_3146 (O_3146,N_29907,N_29854);
xor UO_3147 (O_3147,N_29895,N_29634);
xnor UO_3148 (O_3148,N_29676,N_29839);
and UO_3149 (O_3149,N_29771,N_29643);
xnor UO_3150 (O_3150,N_29841,N_29714);
xor UO_3151 (O_3151,N_29950,N_29909);
nand UO_3152 (O_3152,N_29698,N_29982);
nor UO_3153 (O_3153,N_29979,N_29767);
and UO_3154 (O_3154,N_29833,N_29903);
and UO_3155 (O_3155,N_29576,N_29789);
or UO_3156 (O_3156,N_29915,N_29642);
nand UO_3157 (O_3157,N_29770,N_29685);
or UO_3158 (O_3158,N_29754,N_29775);
or UO_3159 (O_3159,N_29897,N_29535);
xor UO_3160 (O_3160,N_29591,N_29782);
nor UO_3161 (O_3161,N_29977,N_29661);
nand UO_3162 (O_3162,N_29625,N_29874);
nor UO_3163 (O_3163,N_29517,N_29675);
nand UO_3164 (O_3164,N_29553,N_29900);
xor UO_3165 (O_3165,N_29992,N_29773);
nand UO_3166 (O_3166,N_29861,N_29533);
nor UO_3167 (O_3167,N_29585,N_29777);
nand UO_3168 (O_3168,N_29842,N_29690);
and UO_3169 (O_3169,N_29796,N_29534);
nor UO_3170 (O_3170,N_29963,N_29660);
or UO_3171 (O_3171,N_29562,N_29703);
or UO_3172 (O_3172,N_29954,N_29899);
xor UO_3173 (O_3173,N_29823,N_29829);
or UO_3174 (O_3174,N_29648,N_29761);
or UO_3175 (O_3175,N_29518,N_29944);
or UO_3176 (O_3176,N_29801,N_29687);
nand UO_3177 (O_3177,N_29914,N_29573);
or UO_3178 (O_3178,N_29596,N_29564);
nor UO_3179 (O_3179,N_29871,N_29740);
xnor UO_3180 (O_3180,N_29648,N_29518);
nor UO_3181 (O_3181,N_29702,N_29996);
nor UO_3182 (O_3182,N_29570,N_29891);
and UO_3183 (O_3183,N_29608,N_29988);
nor UO_3184 (O_3184,N_29542,N_29755);
or UO_3185 (O_3185,N_29521,N_29892);
xor UO_3186 (O_3186,N_29529,N_29560);
xnor UO_3187 (O_3187,N_29645,N_29831);
and UO_3188 (O_3188,N_29838,N_29673);
nand UO_3189 (O_3189,N_29978,N_29681);
or UO_3190 (O_3190,N_29705,N_29540);
xnor UO_3191 (O_3191,N_29758,N_29573);
nand UO_3192 (O_3192,N_29980,N_29945);
or UO_3193 (O_3193,N_29510,N_29695);
nor UO_3194 (O_3194,N_29926,N_29675);
nand UO_3195 (O_3195,N_29760,N_29643);
xnor UO_3196 (O_3196,N_29931,N_29921);
xor UO_3197 (O_3197,N_29757,N_29895);
and UO_3198 (O_3198,N_29554,N_29611);
nand UO_3199 (O_3199,N_29752,N_29601);
xnor UO_3200 (O_3200,N_29877,N_29725);
and UO_3201 (O_3201,N_29742,N_29810);
nor UO_3202 (O_3202,N_29712,N_29510);
nor UO_3203 (O_3203,N_29561,N_29506);
nand UO_3204 (O_3204,N_29749,N_29920);
nor UO_3205 (O_3205,N_29806,N_29648);
or UO_3206 (O_3206,N_29915,N_29519);
and UO_3207 (O_3207,N_29694,N_29602);
nand UO_3208 (O_3208,N_29873,N_29547);
nor UO_3209 (O_3209,N_29656,N_29887);
nand UO_3210 (O_3210,N_29673,N_29878);
and UO_3211 (O_3211,N_29949,N_29683);
xnor UO_3212 (O_3212,N_29596,N_29851);
nand UO_3213 (O_3213,N_29521,N_29912);
nor UO_3214 (O_3214,N_29874,N_29777);
xor UO_3215 (O_3215,N_29643,N_29906);
nand UO_3216 (O_3216,N_29980,N_29999);
nor UO_3217 (O_3217,N_29796,N_29572);
xnor UO_3218 (O_3218,N_29548,N_29582);
and UO_3219 (O_3219,N_29915,N_29597);
and UO_3220 (O_3220,N_29724,N_29920);
and UO_3221 (O_3221,N_29601,N_29818);
and UO_3222 (O_3222,N_29768,N_29770);
or UO_3223 (O_3223,N_29525,N_29668);
nand UO_3224 (O_3224,N_29511,N_29549);
or UO_3225 (O_3225,N_29619,N_29769);
and UO_3226 (O_3226,N_29893,N_29615);
or UO_3227 (O_3227,N_29535,N_29714);
xor UO_3228 (O_3228,N_29648,N_29920);
or UO_3229 (O_3229,N_29841,N_29709);
or UO_3230 (O_3230,N_29971,N_29902);
nor UO_3231 (O_3231,N_29912,N_29833);
and UO_3232 (O_3232,N_29650,N_29897);
nor UO_3233 (O_3233,N_29634,N_29683);
xor UO_3234 (O_3234,N_29500,N_29804);
or UO_3235 (O_3235,N_29680,N_29738);
nor UO_3236 (O_3236,N_29858,N_29955);
nand UO_3237 (O_3237,N_29593,N_29939);
nor UO_3238 (O_3238,N_29827,N_29620);
or UO_3239 (O_3239,N_29900,N_29933);
nand UO_3240 (O_3240,N_29954,N_29880);
nand UO_3241 (O_3241,N_29589,N_29743);
or UO_3242 (O_3242,N_29675,N_29670);
and UO_3243 (O_3243,N_29868,N_29744);
xnor UO_3244 (O_3244,N_29998,N_29534);
nand UO_3245 (O_3245,N_29943,N_29997);
nor UO_3246 (O_3246,N_29808,N_29568);
nor UO_3247 (O_3247,N_29853,N_29981);
nand UO_3248 (O_3248,N_29519,N_29891);
and UO_3249 (O_3249,N_29600,N_29835);
xor UO_3250 (O_3250,N_29851,N_29681);
or UO_3251 (O_3251,N_29521,N_29734);
xor UO_3252 (O_3252,N_29707,N_29875);
xnor UO_3253 (O_3253,N_29876,N_29550);
and UO_3254 (O_3254,N_29832,N_29714);
nor UO_3255 (O_3255,N_29871,N_29938);
nand UO_3256 (O_3256,N_29555,N_29602);
and UO_3257 (O_3257,N_29842,N_29681);
or UO_3258 (O_3258,N_29613,N_29758);
and UO_3259 (O_3259,N_29671,N_29862);
and UO_3260 (O_3260,N_29606,N_29707);
nand UO_3261 (O_3261,N_29569,N_29759);
and UO_3262 (O_3262,N_29952,N_29731);
nor UO_3263 (O_3263,N_29919,N_29609);
nor UO_3264 (O_3264,N_29666,N_29925);
xnor UO_3265 (O_3265,N_29844,N_29953);
nor UO_3266 (O_3266,N_29774,N_29608);
or UO_3267 (O_3267,N_29897,N_29699);
xor UO_3268 (O_3268,N_29803,N_29520);
xnor UO_3269 (O_3269,N_29707,N_29834);
xnor UO_3270 (O_3270,N_29775,N_29752);
or UO_3271 (O_3271,N_29955,N_29866);
or UO_3272 (O_3272,N_29557,N_29673);
or UO_3273 (O_3273,N_29732,N_29688);
or UO_3274 (O_3274,N_29548,N_29869);
and UO_3275 (O_3275,N_29966,N_29566);
nand UO_3276 (O_3276,N_29850,N_29839);
xor UO_3277 (O_3277,N_29624,N_29800);
and UO_3278 (O_3278,N_29960,N_29543);
nand UO_3279 (O_3279,N_29562,N_29600);
nor UO_3280 (O_3280,N_29897,N_29759);
and UO_3281 (O_3281,N_29690,N_29990);
or UO_3282 (O_3282,N_29567,N_29611);
xor UO_3283 (O_3283,N_29875,N_29664);
nor UO_3284 (O_3284,N_29900,N_29672);
nor UO_3285 (O_3285,N_29618,N_29980);
xnor UO_3286 (O_3286,N_29817,N_29764);
xnor UO_3287 (O_3287,N_29989,N_29555);
or UO_3288 (O_3288,N_29620,N_29614);
nor UO_3289 (O_3289,N_29547,N_29833);
or UO_3290 (O_3290,N_29644,N_29562);
nor UO_3291 (O_3291,N_29714,N_29718);
or UO_3292 (O_3292,N_29916,N_29889);
nand UO_3293 (O_3293,N_29916,N_29819);
xor UO_3294 (O_3294,N_29872,N_29568);
or UO_3295 (O_3295,N_29948,N_29630);
xnor UO_3296 (O_3296,N_29570,N_29632);
or UO_3297 (O_3297,N_29802,N_29836);
and UO_3298 (O_3298,N_29687,N_29972);
or UO_3299 (O_3299,N_29634,N_29726);
nand UO_3300 (O_3300,N_29655,N_29586);
or UO_3301 (O_3301,N_29809,N_29937);
or UO_3302 (O_3302,N_29936,N_29814);
nand UO_3303 (O_3303,N_29820,N_29627);
and UO_3304 (O_3304,N_29877,N_29576);
nand UO_3305 (O_3305,N_29973,N_29877);
and UO_3306 (O_3306,N_29686,N_29639);
or UO_3307 (O_3307,N_29688,N_29510);
and UO_3308 (O_3308,N_29903,N_29565);
nor UO_3309 (O_3309,N_29807,N_29731);
nand UO_3310 (O_3310,N_29907,N_29923);
xor UO_3311 (O_3311,N_29631,N_29953);
nor UO_3312 (O_3312,N_29856,N_29670);
xor UO_3313 (O_3313,N_29758,N_29912);
xnor UO_3314 (O_3314,N_29873,N_29860);
nand UO_3315 (O_3315,N_29636,N_29510);
nor UO_3316 (O_3316,N_29509,N_29781);
and UO_3317 (O_3317,N_29861,N_29722);
or UO_3318 (O_3318,N_29881,N_29624);
xnor UO_3319 (O_3319,N_29850,N_29738);
and UO_3320 (O_3320,N_29816,N_29521);
nor UO_3321 (O_3321,N_29901,N_29685);
or UO_3322 (O_3322,N_29887,N_29657);
nand UO_3323 (O_3323,N_29740,N_29975);
nor UO_3324 (O_3324,N_29638,N_29697);
nand UO_3325 (O_3325,N_29618,N_29686);
xor UO_3326 (O_3326,N_29921,N_29865);
or UO_3327 (O_3327,N_29673,N_29640);
and UO_3328 (O_3328,N_29787,N_29776);
or UO_3329 (O_3329,N_29708,N_29917);
nand UO_3330 (O_3330,N_29573,N_29659);
or UO_3331 (O_3331,N_29643,N_29646);
nor UO_3332 (O_3332,N_29781,N_29557);
xnor UO_3333 (O_3333,N_29529,N_29615);
or UO_3334 (O_3334,N_29540,N_29678);
nand UO_3335 (O_3335,N_29626,N_29950);
or UO_3336 (O_3336,N_29611,N_29520);
nand UO_3337 (O_3337,N_29841,N_29748);
nand UO_3338 (O_3338,N_29919,N_29952);
xnor UO_3339 (O_3339,N_29736,N_29894);
xnor UO_3340 (O_3340,N_29674,N_29848);
or UO_3341 (O_3341,N_29532,N_29869);
nor UO_3342 (O_3342,N_29518,N_29625);
and UO_3343 (O_3343,N_29810,N_29634);
and UO_3344 (O_3344,N_29902,N_29650);
nor UO_3345 (O_3345,N_29518,N_29581);
xnor UO_3346 (O_3346,N_29537,N_29590);
and UO_3347 (O_3347,N_29532,N_29672);
nor UO_3348 (O_3348,N_29875,N_29674);
nor UO_3349 (O_3349,N_29977,N_29550);
nand UO_3350 (O_3350,N_29838,N_29865);
xnor UO_3351 (O_3351,N_29655,N_29567);
xnor UO_3352 (O_3352,N_29922,N_29508);
xor UO_3353 (O_3353,N_29962,N_29838);
xor UO_3354 (O_3354,N_29796,N_29575);
and UO_3355 (O_3355,N_29932,N_29780);
xnor UO_3356 (O_3356,N_29919,N_29780);
or UO_3357 (O_3357,N_29601,N_29784);
nor UO_3358 (O_3358,N_29595,N_29636);
or UO_3359 (O_3359,N_29830,N_29827);
and UO_3360 (O_3360,N_29881,N_29887);
or UO_3361 (O_3361,N_29532,N_29935);
nor UO_3362 (O_3362,N_29521,N_29990);
nor UO_3363 (O_3363,N_29594,N_29974);
or UO_3364 (O_3364,N_29678,N_29729);
nand UO_3365 (O_3365,N_29622,N_29946);
xor UO_3366 (O_3366,N_29502,N_29841);
nor UO_3367 (O_3367,N_29908,N_29923);
nor UO_3368 (O_3368,N_29845,N_29940);
nand UO_3369 (O_3369,N_29985,N_29876);
or UO_3370 (O_3370,N_29539,N_29826);
nand UO_3371 (O_3371,N_29780,N_29513);
and UO_3372 (O_3372,N_29910,N_29678);
or UO_3373 (O_3373,N_29844,N_29681);
and UO_3374 (O_3374,N_29882,N_29590);
xnor UO_3375 (O_3375,N_29551,N_29823);
nor UO_3376 (O_3376,N_29600,N_29525);
nor UO_3377 (O_3377,N_29524,N_29621);
nor UO_3378 (O_3378,N_29563,N_29525);
nor UO_3379 (O_3379,N_29698,N_29509);
nand UO_3380 (O_3380,N_29896,N_29634);
or UO_3381 (O_3381,N_29629,N_29813);
nor UO_3382 (O_3382,N_29683,N_29704);
nand UO_3383 (O_3383,N_29759,N_29619);
xor UO_3384 (O_3384,N_29942,N_29865);
nand UO_3385 (O_3385,N_29821,N_29832);
nand UO_3386 (O_3386,N_29969,N_29851);
xor UO_3387 (O_3387,N_29757,N_29820);
nor UO_3388 (O_3388,N_29660,N_29743);
or UO_3389 (O_3389,N_29917,N_29745);
or UO_3390 (O_3390,N_29579,N_29820);
or UO_3391 (O_3391,N_29527,N_29686);
xor UO_3392 (O_3392,N_29745,N_29895);
xnor UO_3393 (O_3393,N_29975,N_29908);
xor UO_3394 (O_3394,N_29510,N_29857);
nand UO_3395 (O_3395,N_29828,N_29502);
nand UO_3396 (O_3396,N_29506,N_29523);
and UO_3397 (O_3397,N_29987,N_29891);
or UO_3398 (O_3398,N_29949,N_29710);
xnor UO_3399 (O_3399,N_29659,N_29881);
and UO_3400 (O_3400,N_29886,N_29835);
nor UO_3401 (O_3401,N_29763,N_29746);
or UO_3402 (O_3402,N_29997,N_29676);
nor UO_3403 (O_3403,N_29990,N_29831);
and UO_3404 (O_3404,N_29732,N_29906);
and UO_3405 (O_3405,N_29864,N_29838);
nor UO_3406 (O_3406,N_29702,N_29685);
and UO_3407 (O_3407,N_29693,N_29550);
and UO_3408 (O_3408,N_29791,N_29556);
nor UO_3409 (O_3409,N_29791,N_29812);
xor UO_3410 (O_3410,N_29973,N_29524);
and UO_3411 (O_3411,N_29868,N_29644);
nor UO_3412 (O_3412,N_29916,N_29593);
and UO_3413 (O_3413,N_29679,N_29924);
nor UO_3414 (O_3414,N_29878,N_29781);
or UO_3415 (O_3415,N_29889,N_29813);
xor UO_3416 (O_3416,N_29783,N_29924);
xnor UO_3417 (O_3417,N_29848,N_29807);
xnor UO_3418 (O_3418,N_29649,N_29687);
nand UO_3419 (O_3419,N_29569,N_29656);
xor UO_3420 (O_3420,N_29980,N_29607);
nand UO_3421 (O_3421,N_29733,N_29846);
nor UO_3422 (O_3422,N_29818,N_29803);
or UO_3423 (O_3423,N_29542,N_29532);
or UO_3424 (O_3424,N_29632,N_29613);
nand UO_3425 (O_3425,N_29778,N_29547);
and UO_3426 (O_3426,N_29699,N_29572);
nor UO_3427 (O_3427,N_29993,N_29908);
xor UO_3428 (O_3428,N_29652,N_29509);
or UO_3429 (O_3429,N_29624,N_29903);
nor UO_3430 (O_3430,N_29863,N_29993);
nand UO_3431 (O_3431,N_29912,N_29810);
nor UO_3432 (O_3432,N_29915,N_29809);
nand UO_3433 (O_3433,N_29827,N_29507);
and UO_3434 (O_3434,N_29594,N_29587);
nand UO_3435 (O_3435,N_29539,N_29782);
and UO_3436 (O_3436,N_29999,N_29531);
and UO_3437 (O_3437,N_29921,N_29859);
xnor UO_3438 (O_3438,N_29522,N_29787);
nor UO_3439 (O_3439,N_29784,N_29722);
nor UO_3440 (O_3440,N_29855,N_29958);
and UO_3441 (O_3441,N_29520,N_29729);
nand UO_3442 (O_3442,N_29662,N_29676);
and UO_3443 (O_3443,N_29746,N_29897);
nand UO_3444 (O_3444,N_29537,N_29602);
or UO_3445 (O_3445,N_29919,N_29581);
nand UO_3446 (O_3446,N_29613,N_29667);
xnor UO_3447 (O_3447,N_29830,N_29572);
xor UO_3448 (O_3448,N_29924,N_29791);
and UO_3449 (O_3449,N_29991,N_29760);
nand UO_3450 (O_3450,N_29691,N_29659);
xnor UO_3451 (O_3451,N_29904,N_29915);
nand UO_3452 (O_3452,N_29640,N_29803);
nor UO_3453 (O_3453,N_29752,N_29799);
and UO_3454 (O_3454,N_29650,N_29935);
and UO_3455 (O_3455,N_29531,N_29620);
or UO_3456 (O_3456,N_29726,N_29713);
and UO_3457 (O_3457,N_29974,N_29704);
or UO_3458 (O_3458,N_29591,N_29646);
xor UO_3459 (O_3459,N_29811,N_29614);
or UO_3460 (O_3460,N_29790,N_29791);
nor UO_3461 (O_3461,N_29884,N_29856);
and UO_3462 (O_3462,N_29774,N_29830);
or UO_3463 (O_3463,N_29920,N_29636);
or UO_3464 (O_3464,N_29827,N_29938);
nor UO_3465 (O_3465,N_29793,N_29589);
nor UO_3466 (O_3466,N_29743,N_29768);
or UO_3467 (O_3467,N_29730,N_29844);
nand UO_3468 (O_3468,N_29983,N_29941);
nand UO_3469 (O_3469,N_29780,N_29903);
nand UO_3470 (O_3470,N_29967,N_29672);
xnor UO_3471 (O_3471,N_29833,N_29960);
nor UO_3472 (O_3472,N_29651,N_29601);
and UO_3473 (O_3473,N_29969,N_29984);
nor UO_3474 (O_3474,N_29599,N_29614);
and UO_3475 (O_3475,N_29959,N_29506);
nor UO_3476 (O_3476,N_29728,N_29508);
nor UO_3477 (O_3477,N_29558,N_29727);
or UO_3478 (O_3478,N_29990,N_29543);
and UO_3479 (O_3479,N_29831,N_29631);
xnor UO_3480 (O_3480,N_29648,N_29918);
nor UO_3481 (O_3481,N_29961,N_29701);
xnor UO_3482 (O_3482,N_29573,N_29687);
and UO_3483 (O_3483,N_29943,N_29999);
or UO_3484 (O_3484,N_29531,N_29768);
xor UO_3485 (O_3485,N_29962,N_29517);
nor UO_3486 (O_3486,N_29591,N_29579);
or UO_3487 (O_3487,N_29633,N_29560);
nor UO_3488 (O_3488,N_29799,N_29517);
xnor UO_3489 (O_3489,N_29930,N_29901);
xnor UO_3490 (O_3490,N_29651,N_29940);
xor UO_3491 (O_3491,N_29999,N_29845);
nor UO_3492 (O_3492,N_29693,N_29744);
xnor UO_3493 (O_3493,N_29612,N_29949);
nand UO_3494 (O_3494,N_29577,N_29855);
xor UO_3495 (O_3495,N_29862,N_29573);
xor UO_3496 (O_3496,N_29573,N_29929);
xnor UO_3497 (O_3497,N_29891,N_29777);
nor UO_3498 (O_3498,N_29975,N_29511);
nor UO_3499 (O_3499,N_29718,N_29826);
endmodule