module basic_500_3000_500_60_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_443,In_300);
or U1 (N_1,In_176,In_223);
nor U2 (N_2,In_413,In_315);
and U3 (N_3,In_138,In_425);
or U4 (N_4,In_8,In_310);
nor U5 (N_5,In_34,In_433);
nand U6 (N_6,In_452,In_25);
nand U7 (N_7,In_270,In_10);
xnor U8 (N_8,In_122,In_233);
nand U9 (N_9,In_330,In_370);
nor U10 (N_10,In_99,In_420);
or U11 (N_11,In_116,In_200);
xor U12 (N_12,In_202,In_195);
nand U13 (N_13,In_216,In_237);
and U14 (N_14,In_489,In_308);
and U15 (N_15,In_448,In_95);
and U16 (N_16,In_44,In_344);
or U17 (N_17,In_183,In_445);
and U18 (N_18,In_230,In_275);
or U19 (N_19,In_459,In_395);
nor U20 (N_20,In_153,In_212);
nor U21 (N_21,In_148,In_201);
and U22 (N_22,In_427,In_105);
nand U23 (N_23,In_389,In_328);
nor U24 (N_24,In_196,In_345);
or U25 (N_25,In_29,In_303);
nor U26 (N_26,In_426,In_170);
or U27 (N_27,In_188,In_410);
nand U28 (N_28,In_74,In_365);
xor U29 (N_29,In_393,In_273);
or U30 (N_30,In_262,In_278);
or U31 (N_31,In_15,In_467);
nor U32 (N_32,In_42,In_161);
and U33 (N_33,In_398,In_260);
nor U34 (N_34,In_31,In_451);
nor U35 (N_35,In_39,In_326);
or U36 (N_36,In_218,In_475);
and U37 (N_37,In_46,In_463);
or U38 (N_38,In_257,In_27);
and U39 (N_39,In_484,In_356);
xor U40 (N_40,In_63,In_460);
and U41 (N_41,In_65,In_479);
nand U42 (N_42,In_14,In_306);
nand U43 (N_43,In_43,In_2);
and U44 (N_44,In_305,In_182);
or U45 (N_45,In_431,In_444);
nand U46 (N_46,In_357,In_466);
and U47 (N_47,In_235,In_352);
and U48 (N_48,In_40,In_5);
or U49 (N_49,In_280,In_59);
nand U50 (N_50,In_491,In_107);
or U51 (N_51,In_418,In_386);
and U52 (N_52,In_104,In_387);
and U53 (N_53,In_89,In_341);
nand U54 (N_54,In_403,N_11);
nor U55 (N_55,In_258,In_261);
nor U56 (N_56,N_45,In_409);
nor U57 (N_57,In_368,In_132);
xnor U58 (N_58,In_391,In_343);
or U59 (N_59,In_19,In_347);
xnor U60 (N_60,In_55,In_332);
and U61 (N_61,In_259,In_400);
and U62 (N_62,In_423,N_24);
nor U63 (N_63,In_49,In_472);
nor U64 (N_64,In_4,N_44);
xor U65 (N_65,In_30,In_435);
and U66 (N_66,In_372,In_297);
nand U67 (N_67,In_399,In_139);
nand U68 (N_68,In_207,In_274);
nor U69 (N_69,In_458,In_87);
nor U70 (N_70,In_211,In_320);
and U71 (N_71,In_316,In_401);
nor U72 (N_72,N_32,In_497);
nand U73 (N_73,In_374,In_193);
nand U74 (N_74,In_494,In_162);
or U75 (N_75,In_119,In_487);
or U76 (N_76,In_392,In_1);
or U77 (N_77,In_437,In_100);
nor U78 (N_78,In_206,In_430);
or U79 (N_79,N_31,In_271);
or U80 (N_80,In_73,In_174);
and U81 (N_81,In_456,N_17);
nor U82 (N_82,In_252,In_247);
or U83 (N_83,In_84,In_377);
nand U84 (N_84,In_323,In_447);
nor U85 (N_85,N_43,In_92);
xnor U86 (N_86,In_208,In_441);
or U87 (N_87,In_376,In_428);
nor U88 (N_88,In_238,In_225);
nor U89 (N_89,In_419,In_301);
nor U90 (N_90,In_164,In_194);
nor U91 (N_91,In_322,In_239);
nor U92 (N_92,In_281,In_381);
xnor U93 (N_93,In_291,In_265);
nor U94 (N_94,In_470,In_351);
nor U95 (N_95,In_91,N_15);
nand U96 (N_96,In_429,In_312);
xnor U97 (N_97,In_33,In_492);
nand U98 (N_98,In_380,In_296);
nand U99 (N_99,In_408,In_78);
nand U100 (N_100,In_318,In_32);
or U101 (N_101,N_95,In_172);
or U102 (N_102,In_125,N_60);
nor U103 (N_103,In_465,In_244);
or U104 (N_104,N_79,In_112);
nand U105 (N_105,In_146,In_482);
or U106 (N_106,In_360,In_66);
nor U107 (N_107,In_254,In_402);
xnor U108 (N_108,In_163,N_23);
and U109 (N_109,In_75,In_128);
nor U110 (N_110,In_324,In_309);
and U111 (N_111,N_39,N_51);
nand U112 (N_112,In_284,In_52);
or U113 (N_113,N_49,N_68);
nand U114 (N_114,In_353,In_295);
xor U115 (N_115,In_285,N_42);
or U116 (N_116,In_106,In_342);
and U117 (N_117,In_455,In_269);
xnor U118 (N_118,N_3,In_179);
and U119 (N_119,In_129,N_99);
nor U120 (N_120,N_35,In_127);
or U121 (N_121,In_251,In_17);
or U122 (N_122,N_34,N_69);
nand U123 (N_123,In_362,In_80);
xor U124 (N_124,In_210,In_219);
or U125 (N_125,N_46,In_354);
nor U126 (N_126,N_9,In_255);
nor U127 (N_127,In_7,N_27);
and U128 (N_128,In_165,N_58);
and U129 (N_129,N_22,In_462);
and U130 (N_130,In_152,In_41);
and U131 (N_131,N_21,In_461);
xnor U132 (N_132,In_485,In_358);
or U133 (N_133,In_481,In_264);
or U134 (N_134,N_96,In_192);
xnor U135 (N_135,In_126,N_38);
and U136 (N_136,In_388,In_468);
and U137 (N_137,In_23,In_248);
and U138 (N_138,N_75,In_131);
and U139 (N_139,In_349,N_94);
nand U140 (N_140,In_147,In_187);
nand U141 (N_141,In_185,In_293);
and U142 (N_142,In_209,In_82);
nor U143 (N_143,In_217,In_151);
nor U144 (N_144,In_77,In_13);
nand U145 (N_145,In_22,N_90);
and U146 (N_146,In_286,In_0);
nor U147 (N_147,In_288,In_102);
or U148 (N_148,In_477,In_474);
nor U149 (N_149,In_340,In_53);
and U150 (N_150,In_68,In_317);
nor U151 (N_151,In_302,In_421);
xor U152 (N_152,In_12,In_375);
nor U153 (N_153,In_90,In_198);
or U154 (N_154,In_180,In_103);
and U155 (N_155,In_97,N_0);
xor U156 (N_156,In_72,In_457);
nand U157 (N_157,N_28,In_81);
xnor U158 (N_158,In_6,In_361);
or U159 (N_159,In_141,N_92);
nand U160 (N_160,In_11,In_268);
or U161 (N_161,In_416,In_136);
nor U162 (N_162,In_79,In_94);
and U163 (N_163,In_229,In_325);
nand U164 (N_164,In_486,In_442);
nor U165 (N_165,In_189,In_499);
nand U166 (N_166,In_167,In_50);
xor U167 (N_167,In_113,In_130);
and U168 (N_168,N_120,In_253);
or U169 (N_169,In_28,In_382);
nor U170 (N_170,N_73,In_114);
or U171 (N_171,N_66,N_82);
nor U172 (N_172,N_111,N_137);
and U173 (N_173,In_110,In_327);
nand U174 (N_174,In_204,In_294);
nand U175 (N_175,N_50,N_116);
and U176 (N_176,N_86,In_199);
or U177 (N_177,In_137,In_16);
or U178 (N_178,N_6,In_243);
nor U179 (N_179,In_57,N_105);
nor U180 (N_180,In_232,N_4);
nand U181 (N_181,In_490,In_85);
xnor U182 (N_182,N_89,In_405);
or U183 (N_183,In_236,In_51);
or U184 (N_184,In_234,In_145);
or U185 (N_185,In_115,In_21);
and U186 (N_186,N_140,In_173);
or U187 (N_187,In_394,In_96);
nor U188 (N_188,In_37,In_156);
or U189 (N_189,In_496,In_287);
or U190 (N_190,In_190,In_337);
or U191 (N_191,In_149,N_134);
or U192 (N_192,N_16,N_26);
and U193 (N_193,In_446,In_118);
or U194 (N_194,In_438,N_5);
and U195 (N_195,N_59,In_140);
xnor U196 (N_196,In_379,N_124);
nor U197 (N_197,In_93,N_104);
nand U198 (N_198,In_123,N_2);
and U199 (N_199,In_478,In_282);
and U200 (N_200,N_185,N_132);
and U201 (N_201,N_199,N_192);
and U202 (N_202,N_64,In_60);
xor U203 (N_203,N_67,In_142);
and U204 (N_204,In_277,In_440);
xor U205 (N_205,N_48,N_83);
and U206 (N_206,N_118,N_72);
and U207 (N_207,In_220,In_283);
and U208 (N_208,N_161,In_488);
xnor U209 (N_209,N_61,In_215);
and U210 (N_210,N_174,In_71);
or U211 (N_211,In_350,In_313);
and U212 (N_212,N_179,N_175);
and U213 (N_213,In_155,In_432);
or U214 (N_214,N_41,N_150);
nor U215 (N_215,In_249,N_53);
nand U216 (N_216,N_54,N_198);
and U217 (N_217,N_165,In_169);
nor U218 (N_218,In_469,In_133);
xor U219 (N_219,In_290,N_162);
nand U220 (N_220,N_20,N_80);
and U221 (N_221,N_178,In_267);
or U222 (N_222,In_120,In_334);
nor U223 (N_223,N_160,In_367);
nand U224 (N_224,N_98,In_240);
and U225 (N_225,N_87,N_109);
or U226 (N_226,N_189,N_148);
nand U227 (N_227,N_10,N_181);
or U228 (N_228,N_171,N_180);
nand U229 (N_229,In_54,N_8);
xor U230 (N_230,N_12,N_40);
or U231 (N_231,In_203,N_65);
and U232 (N_232,In_289,N_141);
and U233 (N_233,N_151,N_125);
nor U234 (N_234,N_85,N_146);
nor U235 (N_235,In_24,In_67);
nor U236 (N_236,N_25,In_221);
and U237 (N_237,In_333,In_58);
nor U238 (N_238,In_366,In_101);
and U239 (N_239,In_414,N_78);
or U240 (N_240,In_224,In_263);
and U241 (N_241,N_183,N_84);
or U242 (N_242,N_177,In_168);
nor U243 (N_243,N_88,In_35);
nand U244 (N_244,N_184,In_61);
or U245 (N_245,In_434,N_112);
and U246 (N_246,N_135,N_114);
xor U247 (N_247,N_47,N_97);
and U248 (N_248,N_106,In_64);
and U249 (N_249,N_7,N_138);
nor U250 (N_250,N_208,N_70);
nor U251 (N_251,In_348,In_157);
or U252 (N_252,In_396,N_164);
xnor U253 (N_253,N_220,N_123);
xnor U254 (N_254,In_412,In_417);
nand U255 (N_255,N_143,In_321);
nor U256 (N_256,N_103,In_48);
nor U257 (N_257,In_339,In_404);
and U258 (N_258,N_227,N_167);
or U259 (N_259,In_18,N_211);
or U260 (N_260,In_384,N_172);
or U261 (N_261,In_422,N_130);
and U262 (N_262,In_464,In_175);
xor U263 (N_263,In_373,N_19);
and U264 (N_264,In_205,In_159);
nand U265 (N_265,N_217,In_359);
and U266 (N_266,N_100,In_454);
nand U267 (N_267,In_378,In_498);
and U268 (N_268,N_93,In_36);
xnor U269 (N_269,In_62,N_126);
and U270 (N_270,In_449,N_243);
and U271 (N_271,N_195,In_453);
or U272 (N_272,In_355,N_62);
nand U273 (N_273,In_471,N_242);
or U274 (N_274,N_237,N_224);
and U275 (N_275,In_186,N_52);
nor U276 (N_276,In_397,N_245);
nand U277 (N_277,N_186,N_18);
or U278 (N_278,N_56,N_155);
nand U279 (N_279,N_115,N_210);
nor U280 (N_280,In_150,N_233);
and U281 (N_281,In_222,N_152);
nand U282 (N_282,N_240,In_184);
and U283 (N_283,In_276,N_156);
and U284 (N_284,N_57,In_228);
nand U285 (N_285,In_158,In_26);
or U286 (N_286,In_385,N_74);
nand U287 (N_287,In_439,N_81);
nand U288 (N_288,In_241,In_473);
nand U289 (N_289,N_158,In_266);
and U290 (N_290,N_207,In_407);
or U291 (N_291,N_222,In_166);
nor U292 (N_292,N_221,In_331);
nor U293 (N_293,N_215,In_88);
nand U294 (N_294,In_70,N_216);
or U295 (N_295,N_136,In_3);
xnor U296 (N_296,N_91,In_314);
and U297 (N_297,N_209,N_117);
and U298 (N_298,N_231,In_108);
nor U299 (N_299,In_480,N_37);
nor U300 (N_300,N_166,N_139);
nor U301 (N_301,N_246,N_280);
and U302 (N_302,N_203,In_178);
and U303 (N_303,N_133,N_241);
nand U304 (N_304,In_450,N_33);
and U305 (N_305,N_145,In_390);
nand U306 (N_306,N_236,In_86);
nand U307 (N_307,N_294,In_256);
and U308 (N_308,N_201,N_267);
nand U309 (N_309,N_204,N_29);
or U310 (N_310,N_234,N_170);
or U311 (N_311,In_299,N_107);
nand U312 (N_312,N_71,N_252);
nor U313 (N_313,N_249,N_144);
nand U314 (N_314,N_238,N_214);
and U315 (N_315,In_98,N_271);
nor U316 (N_316,In_231,N_127);
and U317 (N_317,In_83,N_258);
and U318 (N_318,N_30,N_1);
nor U319 (N_319,N_270,In_177);
xnor U320 (N_320,In_346,N_55);
nor U321 (N_321,N_176,N_278);
or U322 (N_322,In_242,In_436);
nor U323 (N_323,N_268,N_299);
nor U324 (N_324,N_292,N_229);
xor U325 (N_325,N_159,N_239);
xor U326 (N_326,N_259,N_122);
or U327 (N_327,N_119,N_190);
nand U328 (N_328,N_223,N_298);
nand U329 (N_329,In_143,In_20);
xor U330 (N_330,In_69,In_495);
or U331 (N_331,N_226,In_191);
and U332 (N_332,In_38,In_56);
nor U333 (N_333,N_36,In_213);
nor U334 (N_334,N_266,N_254);
and U335 (N_335,In_329,N_182);
or U336 (N_336,N_63,In_493);
and U337 (N_337,N_193,N_274);
or U338 (N_338,N_244,N_286);
and U339 (N_339,N_291,N_257);
or U340 (N_340,In_160,N_285);
nand U341 (N_341,In_304,N_197);
nand U342 (N_342,N_142,N_110);
nor U343 (N_343,In_144,N_250);
or U344 (N_344,In_319,In_47);
and U345 (N_345,In_411,N_213);
nor U346 (N_346,N_235,In_272);
nor U347 (N_347,N_14,In_154);
nor U348 (N_348,In_369,In_415);
nor U349 (N_349,N_297,In_371);
or U350 (N_350,N_349,N_279);
or U351 (N_351,N_272,N_188);
nand U352 (N_352,N_301,N_196);
nand U353 (N_353,N_101,In_197);
and U354 (N_354,N_191,N_338);
nand U355 (N_355,In_363,N_265);
xnor U356 (N_356,N_230,N_316);
or U357 (N_357,N_13,N_323);
and U358 (N_358,N_261,N_327);
and U359 (N_359,N_335,N_315);
nor U360 (N_360,N_228,In_135);
and U361 (N_361,In_9,N_77);
and U362 (N_362,N_232,In_245);
and U363 (N_363,N_248,N_283);
nor U364 (N_364,In_483,N_304);
nand U365 (N_365,In_111,N_318);
nor U366 (N_366,N_331,N_307);
nor U367 (N_367,In_424,N_308);
nor U368 (N_368,In_117,N_319);
xor U369 (N_369,N_269,N_342);
nor U370 (N_370,In_45,N_341);
nor U371 (N_371,In_383,N_153);
nor U372 (N_372,N_121,N_343);
or U373 (N_373,N_276,In_406);
and U374 (N_374,N_321,N_219);
nand U375 (N_375,N_287,N_346);
or U376 (N_376,N_154,N_337);
nor U377 (N_377,N_273,N_313);
or U378 (N_378,In_181,N_218);
xnor U379 (N_379,N_348,N_194);
nor U380 (N_380,In_335,N_317);
and U381 (N_381,N_324,In_246);
and U382 (N_382,N_168,N_340);
nand U383 (N_383,In_279,N_300);
xnor U384 (N_384,N_256,N_247);
and U385 (N_385,N_187,N_108);
and U386 (N_386,N_253,N_202);
nor U387 (N_387,In_338,N_333);
or U388 (N_388,In_336,N_289);
xor U389 (N_389,N_260,N_293);
nand U390 (N_390,In_171,In_307);
nand U391 (N_391,N_284,In_134);
nor U392 (N_392,N_147,N_131);
nand U393 (N_393,In_292,N_345);
and U394 (N_394,In_227,N_128);
nor U395 (N_395,N_329,N_336);
xnor U396 (N_396,In_476,N_263);
nor U397 (N_397,N_339,N_325);
xnor U398 (N_398,N_169,N_309);
or U399 (N_399,N_206,In_226);
or U400 (N_400,N_368,In_214);
and U401 (N_401,N_305,N_296);
nor U402 (N_402,N_360,N_384);
nand U403 (N_403,In_124,N_163);
and U404 (N_404,N_251,N_255);
nand U405 (N_405,N_330,N_389);
nand U406 (N_406,N_352,N_358);
xnor U407 (N_407,N_113,N_385);
and U408 (N_408,N_281,N_361);
and U409 (N_409,N_381,N_364);
nand U410 (N_410,N_295,N_372);
or U411 (N_411,N_351,N_356);
xnor U412 (N_412,N_225,In_250);
and U413 (N_413,N_379,N_303);
nor U414 (N_414,N_399,N_149);
or U415 (N_415,N_332,In_364);
and U416 (N_416,N_377,N_387);
nor U417 (N_417,N_350,N_392);
nor U418 (N_418,N_129,N_102);
and U419 (N_419,N_212,In_76);
or U420 (N_420,N_282,N_374);
nand U421 (N_421,N_376,N_383);
nor U422 (N_422,N_173,In_121);
and U423 (N_423,N_326,N_393);
or U424 (N_424,N_391,N_394);
nor U425 (N_425,N_395,N_200);
or U426 (N_426,N_322,N_320);
nor U427 (N_427,N_363,N_157);
and U428 (N_428,In_298,N_314);
and U429 (N_429,N_382,N_369);
or U430 (N_430,N_396,N_311);
and U431 (N_431,N_375,N_388);
or U432 (N_432,N_290,N_367);
and U433 (N_433,N_365,N_262);
nand U434 (N_434,N_362,N_355);
or U435 (N_435,N_366,N_353);
or U436 (N_436,N_310,N_354);
and U437 (N_437,N_264,N_378);
and U438 (N_438,N_277,N_357);
nor U439 (N_439,N_390,N_371);
nor U440 (N_440,N_288,N_380);
nor U441 (N_441,N_275,In_311);
and U442 (N_442,N_334,N_398);
nor U443 (N_443,N_373,N_302);
nand U444 (N_444,N_306,In_109);
nor U445 (N_445,N_397,N_344);
nand U446 (N_446,N_205,N_359);
or U447 (N_447,N_312,N_386);
and U448 (N_448,N_370,N_328);
nor U449 (N_449,N_76,N_347);
nor U450 (N_450,N_437,N_420);
or U451 (N_451,N_436,N_408);
or U452 (N_452,N_409,N_443);
nand U453 (N_453,N_444,N_400);
nor U454 (N_454,N_422,N_405);
and U455 (N_455,N_431,N_411);
or U456 (N_456,N_415,N_401);
nor U457 (N_457,N_403,N_435);
or U458 (N_458,N_414,N_438);
nand U459 (N_459,N_432,N_410);
nand U460 (N_460,N_434,N_419);
or U461 (N_461,N_428,N_426);
nor U462 (N_462,N_412,N_418);
nand U463 (N_463,N_442,N_448);
or U464 (N_464,N_446,N_407);
and U465 (N_465,N_402,N_430);
nor U466 (N_466,N_440,N_429);
and U467 (N_467,N_433,N_416);
nand U468 (N_468,N_417,N_439);
or U469 (N_469,N_424,N_449);
nor U470 (N_470,N_441,N_413);
and U471 (N_471,N_427,N_421);
nand U472 (N_472,N_404,N_445);
nor U473 (N_473,N_406,N_423);
and U474 (N_474,N_447,N_425);
and U475 (N_475,N_433,N_435);
nand U476 (N_476,N_422,N_417);
or U477 (N_477,N_421,N_435);
or U478 (N_478,N_423,N_433);
or U479 (N_479,N_433,N_430);
nor U480 (N_480,N_424,N_403);
nor U481 (N_481,N_434,N_436);
nand U482 (N_482,N_427,N_424);
nand U483 (N_483,N_416,N_445);
nor U484 (N_484,N_401,N_421);
nor U485 (N_485,N_403,N_433);
and U486 (N_486,N_419,N_427);
and U487 (N_487,N_430,N_432);
nand U488 (N_488,N_417,N_441);
xnor U489 (N_489,N_411,N_429);
or U490 (N_490,N_447,N_448);
xor U491 (N_491,N_441,N_447);
nand U492 (N_492,N_411,N_444);
or U493 (N_493,N_414,N_402);
nand U494 (N_494,N_441,N_402);
and U495 (N_495,N_427,N_442);
or U496 (N_496,N_431,N_439);
xor U497 (N_497,N_444,N_425);
or U498 (N_498,N_446,N_412);
or U499 (N_499,N_419,N_448);
xnor U500 (N_500,N_477,N_488);
nand U501 (N_501,N_476,N_453);
nor U502 (N_502,N_496,N_478);
nor U503 (N_503,N_469,N_460);
and U504 (N_504,N_455,N_481);
nand U505 (N_505,N_497,N_451);
nor U506 (N_506,N_468,N_466);
nand U507 (N_507,N_494,N_465);
and U508 (N_508,N_485,N_490);
or U509 (N_509,N_498,N_470);
nor U510 (N_510,N_487,N_499);
xor U511 (N_511,N_486,N_483);
and U512 (N_512,N_474,N_493);
or U513 (N_513,N_482,N_475);
or U514 (N_514,N_457,N_458);
nand U515 (N_515,N_492,N_464);
xnor U516 (N_516,N_484,N_489);
nand U517 (N_517,N_479,N_461);
or U518 (N_518,N_462,N_450);
or U519 (N_519,N_454,N_480);
nor U520 (N_520,N_471,N_456);
nand U521 (N_521,N_495,N_472);
and U522 (N_522,N_452,N_467);
and U523 (N_523,N_459,N_463);
nand U524 (N_524,N_473,N_491);
or U525 (N_525,N_453,N_470);
and U526 (N_526,N_486,N_454);
nor U527 (N_527,N_466,N_458);
and U528 (N_528,N_498,N_451);
nand U529 (N_529,N_494,N_452);
nor U530 (N_530,N_453,N_486);
or U531 (N_531,N_468,N_467);
nor U532 (N_532,N_474,N_476);
or U533 (N_533,N_499,N_497);
xnor U534 (N_534,N_458,N_489);
or U535 (N_535,N_489,N_486);
nand U536 (N_536,N_458,N_450);
nand U537 (N_537,N_480,N_450);
and U538 (N_538,N_461,N_480);
and U539 (N_539,N_484,N_494);
and U540 (N_540,N_471,N_463);
and U541 (N_541,N_478,N_484);
nor U542 (N_542,N_463,N_457);
or U543 (N_543,N_456,N_476);
nand U544 (N_544,N_458,N_478);
nor U545 (N_545,N_498,N_454);
and U546 (N_546,N_454,N_477);
nor U547 (N_547,N_470,N_477);
xor U548 (N_548,N_457,N_467);
nor U549 (N_549,N_490,N_457);
and U550 (N_550,N_503,N_545);
xor U551 (N_551,N_527,N_506);
or U552 (N_552,N_526,N_538);
nand U553 (N_553,N_543,N_510);
nand U554 (N_554,N_505,N_513);
or U555 (N_555,N_537,N_539);
nor U556 (N_556,N_523,N_528);
and U557 (N_557,N_547,N_500);
or U558 (N_558,N_520,N_546);
nand U559 (N_559,N_535,N_517);
or U560 (N_560,N_508,N_522);
xor U561 (N_561,N_533,N_544);
nor U562 (N_562,N_524,N_501);
or U563 (N_563,N_516,N_507);
and U564 (N_564,N_525,N_536);
or U565 (N_565,N_529,N_548);
or U566 (N_566,N_519,N_530);
and U567 (N_567,N_518,N_549);
nand U568 (N_568,N_502,N_531);
xor U569 (N_569,N_512,N_532);
nor U570 (N_570,N_504,N_534);
nand U571 (N_571,N_514,N_540);
nor U572 (N_572,N_515,N_542);
or U573 (N_573,N_521,N_509);
xnor U574 (N_574,N_511,N_541);
xor U575 (N_575,N_504,N_508);
nand U576 (N_576,N_531,N_510);
or U577 (N_577,N_507,N_544);
xnor U578 (N_578,N_511,N_545);
or U579 (N_579,N_526,N_530);
or U580 (N_580,N_527,N_534);
nor U581 (N_581,N_529,N_544);
or U582 (N_582,N_542,N_517);
or U583 (N_583,N_537,N_530);
nand U584 (N_584,N_520,N_511);
nor U585 (N_585,N_502,N_525);
or U586 (N_586,N_534,N_544);
nand U587 (N_587,N_506,N_518);
and U588 (N_588,N_538,N_511);
and U589 (N_589,N_540,N_517);
and U590 (N_590,N_543,N_539);
nor U591 (N_591,N_538,N_524);
nor U592 (N_592,N_539,N_541);
and U593 (N_593,N_533,N_527);
nand U594 (N_594,N_517,N_513);
nand U595 (N_595,N_508,N_501);
and U596 (N_596,N_500,N_545);
nand U597 (N_597,N_517,N_524);
and U598 (N_598,N_546,N_534);
nand U599 (N_599,N_508,N_513);
nand U600 (N_600,N_576,N_597);
nor U601 (N_601,N_590,N_566);
or U602 (N_602,N_575,N_587);
nor U603 (N_603,N_551,N_569);
nand U604 (N_604,N_561,N_558);
nor U605 (N_605,N_562,N_553);
or U606 (N_606,N_565,N_585);
xor U607 (N_607,N_552,N_598);
or U608 (N_608,N_579,N_555);
nand U609 (N_609,N_583,N_589);
and U610 (N_610,N_570,N_556);
and U611 (N_611,N_560,N_563);
nand U612 (N_612,N_564,N_584);
nand U613 (N_613,N_582,N_554);
and U614 (N_614,N_591,N_577);
and U615 (N_615,N_586,N_572);
nand U616 (N_616,N_595,N_592);
and U617 (N_617,N_588,N_574);
nor U618 (N_618,N_573,N_550);
and U619 (N_619,N_568,N_580);
nand U620 (N_620,N_594,N_593);
nand U621 (N_621,N_571,N_581);
or U622 (N_622,N_596,N_559);
and U623 (N_623,N_578,N_557);
or U624 (N_624,N_567,N_599);
nand U625 (N_625,N_588,N_597);
nor U626 (N_626,N_584,N_553);
or U627 (N_627,N_594,N_561);
nand U628 (N_628,N_584,N_555);
or U629 (N_629,N_552,N_586);
nand U630 (N_630,N_577,N_587);
or U631 (N_631,N_551,N_553);
and U632 (N_632,N_560,N_594);
and U633 (N_633,N_593,N_562);
nor U634 (N_634,N_597,N_550);
xnor U635 (N_635,N_585,N_586);
xor U636 (N_636,N_595,N_575);
nor U637 (N_637,N_593,N_577);
nand U638 (N_638,N_587,N_558);
nor U639 (N_639,N_577,N_589);
nand U640 (N_640,N_557,N_559);
or U641 (N_641,N_599,N_552);
xor U642 (N_642,N_563,N_577);
xnor U643 (N_643,N_565,N_577);
xnor U644 (N_644,N_559,N_582);
or U645 (N_645,N_588,N_583);
nor U646 (N_646,N_555,N_596);
or U647 (N_647,N_552,N_550);
nor U648 (N_648,N_555,N_595);
or U649 (N_649,N_595,N_593);
nor U650 (N_650,N_641,N_607);
or U651 (N_651,N_645,N_612);
xnor U652 (N_652,N_649,N_632);
and U653 (N_653,N_633,N_600);
nand U654 (N_654,N_631,N_614);
or U655 (N_655,N_606,N_642);
and U656 (N_656,N_628,N_638);
xnor U657 (N_657,N_613,N_644);
nand U658 (N_658,N_647,N_620);
xor U659 (N_659,N_601,N_626);
nand U660 (N_660,N_636,N_610);
or U661 (N_661,N_643,N_611);
and U662 (N_662,N_619,N_639);
or U663 (N_663,N_609,N_618);
or U664 (N_664,N_621,N_624);
nor U665 (N_665,N_608,N_646);
nor U666 (N_666,N_605,N_625);
xor U667 (N_667,N_629,N_635);
xnor U668 (N_668,N_640,N_630);
or U669 (N_669,N_615,N_637);
or U670 (N_670,N_616,N_623);
and U671 (N_671,N_603,N_627);
and U672 (N_672,N_617,N_604);
nor U673 (N_673,N_622,N_602);
or U674 (N_674,N_648,N_634);
and U675 (N_675,N_623,N_635);
or U676 (N_676,N_613,N_649);
and U677 (N_677,N_623,N_602);
nand U678 (N_678,N_604,N_608);
nor U679 (N_679,N_648,N_646);
or U680 (N_680,N_607,N_613);
nand U681 (N_681,N_642,N_641);
xnor U682 (N_682,N_636,N_619);
and U683 (N_683,N_640,N_617);
nand U684 (N_684,N_607,N_616);
or U685 (N_685,N_642,N_644);
nor U686 (N_686,N_640,N_627);
nor U687 (N_687,N_638,N_632);
and U688 (N_688,N_641,N_600);
and U689 (N_689,N_624,N_622);
and U690 (N_690,N_622,N_620);
nor U691 (N_691,N_638,N_649);
nand U692 (N_692,N_635,N_624);
and U693 (N_693,N_628,N_625);
nand U694 (N_694,N_602,N_604);
and U695 (N_695,N_623,N_604);
and U696 (N_696,N_634,N_649);
and U697 (N_697,N_626,N_648);
or U698 (N_698,N_641,N_608);
and U699 (N_699,N_614,N_641);
nand U700 (N_700,N_674,N_666);
and U701 (N_701,N_688,N_656);
or U702 (N_702,N_672,N_665);
nor U703 (N_703,N_686,N_676);
and U704 (N_704,N_694,N_658);
and U705 (N_705,N_664,N_690);
nor U706 (N_706,N_697,N_657);
and U707 (N_707,N_653,N_689);
nand U708 (N_708,N_685,N_696);
or U709 (N_709,N_673,N_682);
or U710 (N_710,N_663,N_680);
and U711 (N_711,N_692,N_678);
xnor U712 (N_712,N_651,N_668);
xnor U713 (N_713,N_660,N_655);
nand U714 (N_714,N_675,N_679);
nor U715 (N_715,N_652,N_695);
or U716 (N_716,N_677,N_691);
nor U717 (N_717,N_671,N_661);
and U718 (N_718,N_654,N_693);
nand U719 (N_719,N_687,N_698);
and U720 (N_720,N_669,N_681);
nor U721 (N_721,N_670,N_683);
and U722 (N_722,N_659,N_667);
and U723 (N_723,N_662,N_650);
xnor U724 (N_724,N_699,N_684);
nand U725 (N_725,N_673,N_689);
nor U726 (N_726,N_671,N_679);
xnor U727 (N_727,N_665,N_698);
nand U728 (N_728,N_672,N_658);
nand U729 (N_729,N_691,N_657);
nor U730 (N_730,N_696,N_660);
xnor U731 (N_731,N_655,N_673);
and U732 (N_732,N_667,N_684);
xnor U733 (N_733,N_687,N_681);
nor U734 (N_734,N_687,N_673);
and U735 (N_735,N_692,N_690);
or U736 (N_736,N_652,N_658);
or U737 (N_737,N_654,N_685);
xnor U738 (N_738,N_675,N_689);
and U739 (N_739,N_669,N_683);
or U740 (N_740,N_679,N_669);
and U741 (N_741,N_680,N_658);
nand U742 (N_742,N_662,N_680);
or U743 (N_743,N_689,N_691);
and U744 (N_744,N_653,N_677);
nand U745 (N_745,N_675,N_660);
and U746 (N_746,N_684,N_690);
nand U747 (N_747,N_686,N_692);
or U748 (N_748,N_657,N_661);
or U749 (N_749,N_688,N_687);
nor U750 (N_750,N_713,N_745);
xor U751 (N_751,N_710,N_744);
or U752 (N_752,N_706,N_715);
and U753 (N_753,N_711,N_735);
or U754 (N_754,N_732,N_727);
and U755 (N_755,N_733,N_712);
nand U756 (N_756,N_737,N_721);
or U757 (N_757,N_748,N_718);
or U758 (N_758,N_723,N_747);
xor U759 (N_759,N_728,N_742);
nor U760 (N_760,N_741,N_736);
or U761 (N_761,N_746,N_722);
and U762 (N_762,N_738,N_730);
nand U763 (N_763,N_717,N_716);
and U764 (N_764,N_704,N_725);
nor U765 (N_765,N_714,N_739);
or U766 (N_766,N_724,N_740);
nor U767 (N_767,N_708,N_702);
xnor U768 (N_768,N_749,N_729);
or U769 (N_769,N_726,N_700);
nor U770 (N_770,N_734,N_707);
nor U771 (N_771,N_703,N_709);
or U772 (N_772,N_701,N_720);
xor U773 (N_773,N_731,N_719);
nand U774 (N_774,N_705,N_743);
nand U775 (N_775,N_748,N_701);
nor U776 (N_776,N_712,N_707);
or U777 (N_777,N_747,N_738);
xnor U778 (N_778,N_744,N_748);
nor U779 (N_779,N_700,N_735);
nor U780 (N_780,N_743,N_732);
nand U781 (N_781,N_701,N_742);
and U782 (N_782,N_709,N_740);
xnor U783 (N_783,N_720,N_736);
or U784 (N_784,N_714,N_742);
nand U785 (N_785,N_706,N_720);
xnor U786 (N_786,N_739,N_709);
and U787 (N_787,N_706,N_728);
nand U788 (N_788,N_736,N_700);
and U789 (N_789,N_740,N_725);
or U790 (N_790,N_700,N_744);
and U791 (N_791,N_736,N_748);
or U792 (N_792,N_715,N_749);
nand U793 (N_793,N_729,N_708);
and U794 (N_794,N_743,N_704);
nor U795 (N_795,N_731,N_735);
nand U796 (N_796,N_747,N_734);
nor U797 (N_797,N_744,N_740);
and U798 (N_798,N_715,N_738);
nor U799 (N_799,N_715,N_724);
nand U800 (N_800,N_754,N_779);
and U801 (N_801,N_788,N_778);
nor U802 (N_802,N_758,N_798);
or U803 (N_803,N_785,N_792);
xnor U804 (N_804,N_761,N_768);
and U805 (N_805,N_751,N_781);
nand U806 (N_806,N_782,N_763);
or U807 (N_807,N_795,N_765);
or U808 (N_808,N_775,N_790);
or U809 (N_809,N_770,N_777);
and U810 (N_810,N_756,N_771);
or U811 (N_811,N_789,N_755);
and U812 (N_812,N_786,N_794);
nor U813 (N_813,N_772,N_762);
or U814 (N_814,N_773,N_774);
nand U815 (N_815,N_766,N_783);
nor U816 (N_816,N_753,N_780);
nand U817 (N_817,N_776,N_767);
xnor U818 (N_818,N_769,N_796);
xor U819 (N_819,N_760,N_750);
xnor U820 (N_820,N_793,N_797);
and U821 (N_821,N_787,N_791);
nor U822 (N_822,N_752,N_759);
nor U823 (N_823,N_784,N_799);
and U824 (N_824,N_757,N_764);
nand U825 (N_825,N_782,N_762);
and U826 (N_826,N_787,N_783);
nor U827 (N_827,N_763,N_757);
and U828 (N_828,N_770,N_795);
and U829 (N_829,N_753,N_785);
and U830 (N_830,N_781,N_778);
xnor U831 (N_831,N_793,N_764);
and U832 (N_832,N_780,N_793);
nor U833 (N_833,N_790,N_799);
xnor U834 (N_834,N_783,N_775);
or U835 (N_835,N_769,N_760);
and U836 (N_836,N_788,N_754);
and U837 (N_837,N_785,N_771);
or U838 (N_838,N_754,N_768);
or U839 (N_839,N_769,N_758);
nand U840 (N_840,N_773,N_768);
and U841 (N_841,N_787,N_798);
nor U842 (N_842,N_775,N_750);
nor U843 (N_843,N_765,N_775);
nor U844 (N_844,N_766,N_799);
or U845 (N_845,N_782,N_771);
xor U846 (N_846,N_766,N_797);
nand U847 (N_847,N_757,N_760);
and U848 (N_848,N_788,N_781);
or U849 (N_849,N_799,N_797);
or U850 (N_850,N_842,N_826);
and U851 (N_851,N_810,N_806);
nor U852 (N_852,N_813,N_833);
or U853 (N_853,N_824,N_821);
nand U854 (N_854,N_823,N_846);
and U855 (N_855,N_819,N_820);
and U856 (N_856,N_814,N_838);
nor U857 (N_857,N_836,N_828);
and U858 (N_858,N_849,N_804);
or U859 (N_859,N_840,N_839);
and U860 (N_860,N_811,N_802);
nor U861 (N_861,N_812,N_831);
nor U862 (N_862,N_808,N_817);
nand U863 (N_863,N_844,N_822);
or U864 (N_864,N_841,N_809);
and U865 (N_865,N_827,N_830);
nand U866 (N_866,N_847,N_834);
or U867 (N_867,N_835,N_829);
nand U868 (N_868,N_816,N_815);
nand U869 (N_869,N_848,N_843);
and U870 (N_870,N_832,N_800);
nand U871 (N_871,N_803,N_807);
and U872 (N_872,N_825,N_805);
xor U873 (N_873,N_845,N_837);
or U874 (N_874,N_818,N_801);
nand U875 (N_875,N_832,N_836);
nand U876 (N_876,N_845,N_824);
nor U877 (N_877,N_835,N_817);
or U878 (N_878,N_816,N_834);
and U879 (N_879,N_815,N_830);
xnor U880 (N_880,N_829,N_816);
or U881 (N_881,N_847,N_810);
and U882 (N_882,N_831,N_839);
nor U883 (N_883,N_841,N_808);
nand U884 (N_884,N_845,N_813);
xnor U885 (N_885,N_803,N_808);
and U886 (N_886,N_841,N_824);
and U887 (N_887,N_823,N_827);
and U888 (N_888,N_846,N_833);
nor U889 (N_889,N_800,N_804);
and U890 (N_890,N_829,N_837);
nand U891 (N_891,N_846,N_805);
or U892 (N_892,N_841,N_805);
xnor U893 (N_893,N_808,N_801);
or U894 (N_894,N_804,N_836);
nor U895 (N_895,N_808,N_843);
and U896 (N_896,N_815,N_819);
and U897 (N_897,N_813,N_817);
nor U898 (N_898,N_826,N_822);
nor U899 (N_899,N_818,N_843);
and U900 (N_900,N_899,N_880);
xnor U901 (N_901,N_864,N_866);
xnor U902 (N_902,N_873,N_856);
or U903 (N_903,N_883,N_869);
xnor U904 (N_904,N_885,N_875);
nand U905 (N_905,N_892,N_890);
xor U906 (N_906,N_886,N_888);
nand U907 (N_907,N_857,N_897);
and U908 (N_908,N_874,N_895);
xnor U909 (N_909,N_850,N_858);
or U910 (N_910,N_855,N_896);
and U911 (N_911,N_863,N_854);
nand U912 (N_912,N_878,N_865);
nand U913 (N_913,N_884,N_881);
nand U914 (N_914,N_887,N_876);
or U915 (N_915,N_853,N_859);
and U916 (N_916,N_877,N_872);
and U917 (N_917,N_889,N_894);
nor U918 (N_918,N_879,N_882);
xnor U919 (N_919,N_868,N_870);
and U920 (N_920,N_871,N_862);
and U921 (N_921,N_852,N_893);
nand U922 (N_922,N_860,N_851);
nand U923 (N_923,N_898,N_891);
and U924 (N_924,N_861,N_867);
and U925 (N_925,N_894,N_873);
or U926 (N_926,N_879,N_885);
and U927 (N_927,N_892,N_871);
and U928 (N_928,N_887,N_853);
and U929 (N_929,N_884,N_869);
nand U930 (N_930,N_886,N_859);
nand U931 (N_931,N_881,N_883);
or U932 (N_932,N_878,N_895);
and U933 (N_933,N_861,N_860);
and U934 (N_934,N_883,N_889);
and U935 (N_935,N_864,N_876);
or U936 (N_936,N_891,N_877);
xor U937 (N_937,N_870,N_873);
nand U938 (N_938,N_880,N_883);
or U939 (N_939,N_899,N_852);
nand U940 (N_940,N_886,N_892);
nor U941 (N_941,N_888,N_869);
nand U942 (N_942,N_875,N_894);
or U943 (N_943,N_850,N_865);
and U944 (N_944,N_877,N_865);
and U945 (N_945,N_873,N_872);
and U946 (N_946,N_879,N_886);
nor U947 (N_947,N_895,N_873);
or U948 (N_948,N_872,N_880);
xor U949 (N_949,N_887,N_863);
and U950 (N_950,N_917,N_921);
or U951 (N_951,N_909,N_903);
or U952 (N_952,N_919,N_918);
nand U953 (N_953,N_941,N_933);
or U954 (N_954,N_938,N_949);
nand U955 (N_955,N_911,N_915);
nand U956 (N_956,N_905,N_914);
or U957 (N_957,N_902,N_940);
and U958 (N_958,N_908,N_929);
nor U959 (N_959,N_936,N_939);
nor U960 (N_960,N_906,N_925);
nor U961 (N_961,N_920,N_943);
and U962 (N_962,N_907,N_934);
nor U963 (N_963,N_928,N_948);
nor U964 (N_964,N_924,N_901);
or U965 (N_965,N_932,N_904);
nand U966 (N_966,N_913,N_912);
nand U967 (N_967,N_916,N_944);
nand U968 (N_968,N_947,N_900);
nor U969 (N_969,N_930,N_931);
or U970 (N_970,N_946,N_922);
and U971 (N_971,N_945,N_927);
nand U972 (N_972,N_923,N_926);
xor U973 (N_973,N_937,N_942);
nand U974 (N_974,N_935,N_910);
nor U975 (N_975,N_933,N_925);
or U976 (N_976,N_901,N_903);
and U977 (N_977,N_912,N_930);
nor U978 (N_978,N_929,N_916);
and U979 (N_979,N_943,N_911);
or U980 (N_980,N_925,N_919);
nand U981 (N_981,N_918,N_930);
or U982 (N_982,N_931,N_905);
and U983 (N_983,N_936,N_927);
or U984 (N_984,N_902,N_933);
nand U985 (N_985,N_934,N_902);
nand U986 (N_986,N_908,N_935);
and U987 (N_987,N_919,N_930);
nand U988 (N_988,N_908,N_912);
or U989 (N_989,N_929,N_915);
nand U990 (N_990,N_948,N_916);
xnor U991 (N_991,N_949,N_936);
xnor U992 (N_992,N_928,N_902);
or U993 (N_993,N_935,N_939);
and U994 (N_994,N_900,N_907);
nor U995 (N_995,N_902,N_911);
nor U996 (N_996,N_929,N_937);
and U997 (N_997,N_905,N_927);
nor U998 (N_998,N_930,N_905);
nand U999 (N_999,N_943,N_916);
or U1000 (N_1000,N_998,N_995);
and U1001 (N_1001,N_983,N_973);
and U1002 (N_1002,N_980,N_962);
nor U1003 (N_1003,N_991,N_959);
and U1004 (N_1004,N_992,N_964);
nand U1005 (N_1005,N_982,N_999);
nor U1006 (N_1006,N_993,N_972);
and U1007 (N_1007,N_954,N_970);
and U1008 (N_1008,N_971,N_966);
or U1009 (N_1009,N_956,N_981);
nand U1010 (N_1010,N_987,N_965);
and U1011 (N_1011,N_952,N_996);
nor U1012 (N_1012,N_950,N_990);
xor U1013 (N_1013,N_994,N_997);
nor U1014 (N_1014,N_963,N_958);
and U1015 (N_1015,N_989,N_988);
nor U1016 (N_1016,N_967,N_978);
or U1017 (N_1017,N_979,N_961);
or U1018 (N_1018,N_975,N_955);
xnor U1019 (N_1019,N_984,N_953);
or U1020 (N_1020,N_969,N_985);
nor U1021 (N_1021,N_974,N_977);
nor U1022 (N_1022,N_976,N_968);
nor U1023 (N_1023,N_960,N_986);
xor U1024 (N_1024,N_957,N_951);
nand U1025 (N_1025,N_964,N_951);
nor U1026 (N_1026,N_954,N_979);
nand U1027 (N_1027,N_983,N_972);
nand U1028 (N_1028,N_997,N_962);
nand U1029 (N_1029,N_990,N_982);
nor U1030 (N_1030,N_966,N_990);
nand U1031 (N_1031,N_998,N_984);
xor U1032 (N_1032,N_957,N_992);
and U1033 (N_1033,N_985,N_982);
nor U1034 (N_1034,N_959,N_970);
nand U1035 (N_1035,N_968,N_958);
or U1036 (N_1036,N_964,N_972);
and U1037 (N_1037,N_990,N_972);
nand U1038 (N_1038,N_977,N_983);
nand U1039 (N_1039,N_950,N_962);
nand U1040 (N_1040,N_997,N_978);
or U1041 (N_1041,N_985,N_954);
and U1042 (N_1042,N_976,N_987);
and U1043 (N_1043,N_963,N_961);
xnor U1044 (N_1044,N_954,N_967);
or U1045 (N_1045,N_964,N_983);
xnor U1046 (N_1046,N_994,N_955);
nand U1047 (N_1047,N_999,N_976);
nor U1048 (N_1048,N_955,N_968);
and U1049 (N_1049,N_967,N_984);
xor U1050 (N_1050,N_1046,N_1008);
nand U1051 (N_1051,N_1035,N_1041);
or U1052 (N_1052,N_1039,N_1011);
or U1053 (N_1053,N_1036,N_1038);
nor U1054 (N_1054,N_1015,N_1049);
nor U1055 (N_1055,N_1048,N_1042);
or U1056 (N_1056,N_1045,N_1006);
and U1057 (N_1057,N_1021,N_1002);
nor U1058 (N_1058,N_1023,N_1017);
xor U1059 (N_1059,N_1016,N_1024);
and U1060 (N_1060,N_1040,N_1020);
and U1061 (N_1061,N_1029,N_1005);
or U1062 (N_1062,N_1009,N_1004);
nand U1063 (N_1063,N_1034,N_1018);
and U1064 (N_1064,N_1001,N_1030);
nand U1065 (N_1065,N_1047,N_1044);
xor U1066 (N_1066,N_1026,N_1019);
nor U1067 (N_1067,N_1028,N_1037);
or U1068 (N_1068,N_1022,N_1027);
or U1069 (N_1069,N_1013,N_1014);
xor U1070 (N_1070,N_1000,N_1032);
nor U1071 (N_1071,N_1031,N_1033);
nand U1072 (N_1072,N_1007,N_1043);
xor U1073 (N_1073,N_1025,N_1003);
nor U1074 (N_1074,N_1010,N_1012);
or U1075 (N_1075,N_1028,N_1036);
nand U1076 (N_1076,N_1000,N_1004);
nand U1077 (N_1077,N_1047,N_1028);
nand U1078 (N_1078,N_1021,N_1035);
and U1079 (N_1079,N_1046,N_1010);
nor U1080 (N_1080,N_1022,N_1008);
nand U1081 (N_1081,N_1006,N_1031);
nor U1082 (N_1082,N_1047,N_1041);
or U1083 (N_1083,N_1000,N_1011);
nor U1084 (N_1084,N_1003,N_1019);
or U1085 (N_1085,N_1043,N_1039);
or U1086 (N_1086,N_1003,N_1016);
xnor U1087 (N_1087,N_1045,N_1029);
xor U1088 (N_1088,N_1000,N_1006);
nand U1089 (N_1089,N_1047,N_1010);
and U1090 (N_1090,N_1044,N_1037);
nand U1091 (N_1091,N_1039,N_1048);
nor U1092 (N_1092,N_1025,N_1043);
xnor U1093 (N_1093,N_1033,N_1038);
nor U1094 (N_1094,N_1018,N_1016);
nand U1095 (N_1095,N_1001,N_1031);
nor U1096 (N_1096,N_1044,N_1031);
xnor U1097 (N_1097,N_1038,N_1022);
or U1098 (N_1098,N_1046,N_1038);
or U1099 (N_1099,N_1034,N_1011);
and U1100 (N_1100,N_1087,N_1083);
and U1101 (N_1101,N_1060,N_1056);
and U1102 (N_1102,N_1064,N_1081);
nor U1103 (N_1103,N_1057,N_1065);
xor U1104 (N_1104,N_1079,N_1093);
or U1105 (N_1105,N_1073,N_1097);
nor U1106 (N_1106,N_1091,N_1092);
nand U1107 (N_1107,N_1085,N_1052);
nand U1108 (N_1108,N_1053,N_1059);
nand U1109 (N_1109,N_1062,N_1090);
nor U1110 (N_1110,N_1088,N_1099);
nand U1111 (N_1111,N_1095,N_1072);
and U1112 (N_1112,N_1068,N_1075);
xnor U1113 (N_1113,N_1086,N_1070);
nand U1114 (N_1114,N_1063,N_1082);
nand U1115 (N_1115,N_1051,N_1084);
or U1116 (N_1116,N_1071,N_1098);
or U1117 (N_1117,N_1078,N_1058);
or U1118 (N_1118,N_1077,N_1080);
nand U1119 (N_1119,N_1074,N_1055);
and U1120 (N_1120,N_1076,N_1061);
nor U1121 (N_1121,N_1067,N_1089);
nand U1122 (N_1122,N_1094,N_1054);
or U1123 (N_1123,N_1050,N_1096);
or U1124 (N_1124,N_1069,N_1066);
nor U1125 (N_1125,N_1099,N_1058);
nand U1126 (N_1126,N_1081,N_1099);
or U1127 (N_1127,N_1089,N_1094);
nor U1128 (N_1128,N_1096,N_1099);
and U1129 (N_1129,N_1058,N_1053);
and U1130 (N_1130,N_1081,N_1097);
and U1131 (N_1131,N_1091,N_1052);
or U1132 (N_1132,N_1070,N_1097);
xnor U1133 (N_1133,N_1097,N_1079);
nand U1134 (N_1134,N_1091,N_1078);
and U1135 (N_1135,N_1091,N_1067);
nand U1136 (N_1136,N_1066,N_1074);
xnor U1137 (N_1137,N_1082,N_1094);
nand U1138 (N_1138,N_1053,N_1082);
nor U1139 (N_1139,N_1065,N_1066);
nand U1140 (N_1140,N_1050,N_1080);
and U1141 (N_1141,N_1069,N_1094);
nand U1142 (N_1142,N_1078,N_1086);
and U1143 (N_1143,N_1050,N_1065);
nand U1144 (N_1144,N_1098,N_1088);
nor U1145 (N_1145,N_1071,N_1061);
nor U1146 (N_1146,N_1089,N_1062);
nand U1147 (N_1147,N_1072,N_1061);
nor U1148 (N_1148,N_1071,N_1062);
and U1149 (N_1149,N_1064,N_1053);
or U1150 (N_1150,N_1137,N_1142);
or U1151 (N_1151,N_1131,N_1121);
and U1152 (N_1152,N_1107,N_1118);
nand U1153 (N_1153,N_1125,N_1119);
and U1154 (N_1154,N_1144,N_1130);
or U1155 (N_1155,N_1115,N_1146);
or U1156 (N_1156,N_1104,N_1128);
nand U1157 (N_1157,N_1106,N_1133);
nor U1158 (N_1158,N_1109,N_1143);
nand U1159 (N_1159,N_1135,N_1122);
nand U1160 (N_1160,N_1129,N_1145);
and U1161 (N_1161,N_1149,N_1127);
nor U1162 (N_1162,N_1140,N_1105);
or U1163 (N_1163,N_1116,N_1141);
nor U1164 (N_1164,N_1138,N_1117);
nor U1165 (N_1165,N_1103,N_1132);
xor U1166 (N_1166,N_1136,N_1113);
and U1167 (N_1167,N_1100,N_1102);
nand U1168 (N_1168,N_1120,N_1139);
and U1169 (N_1169,N_1111,N_1114);
and U1170 (N_1170,N_1101,N_1126);
nor U1171 (N_1171,N_1108,N_1134);
nand U1172 (N_1172,N_1124,N_1123);
nor U1173 (N_1173,N_1147,N_1110);
and U1174 (N_1174,N_1148,N_1112);
nand U1175 (N_1175,N_1122,N_1129);
xnor U1176 (N_1176,N_1107,N_1127);
nand U1177 (N_1177,N_1132,N_1123);
or U1178 (N_1178,N_1120,N_1138);
xor U1179 (N_1179,N_1146,N_1132);
nand U1180 (N_1180,N_1135,N_1104);
or U1181 (N_1181,N_1110,N_1140);
xnor U1182 (N_1182,N_1125,N_1116);
nor U1183 (N_1183,N_1131,N_1107);
nand U1184 (N_1184,N_1118,N_1145);
nor U1185 (N_1185,N_1132,N_1131);
and U1186 (N_1186,N_1106,N_1125);
and U1187 (N_1187,N_1104,N_1108);
nor U1188 (N_1188,N_1115,N_1121);
and U1189 (N_1189,N_1120,N_1143);
nand U1190 (N_1190,N_1124,N_1128);
and U1191 (N_1191,N_1118,N_1144);
nand U1192 (N_1192,N_1147,N_1108);
or U1193 (N_1193,N_1131,N_1106);
nand U1194 (N_1194,N_1123,N_1148);
nand U1195 (N_1195,N_1109,N_1103);
or U1196 (N_1196,N_1144,N_1149);
nand U1197 (N_1197,N_1146,N_1131);
nand U1198 (N_1198,N_1133,N_1126);
or U1199 (N_1199,N_1143,N_1145);
or U1200 (N_1200,N_1181,N_1169);
and U1201 (N_1201,N_1156,N_1185);
and U1202 (N_1202,N_1163,N_1170);
nand U1203 (N_1203,N_1153,N_1188);
or U1204 (N_1204,N_1162,N_1180);
nor U1205 (N_1205,N_1167,N_1178);
nand U1206 (N_1206,N_1189,N_1191);
and U1207 (N_1207,N_1174,N_1158);
or U1208 (N_1208,N_1194,N_1193);
and U1209 (N_1209,N_1197,N_1152);
and U1210 (N_1210,N_1184,N_1157);
and U1211 (N_1211,N_1175,N_1160);
or U1212 (N_1212,N_1192,N_1199);
nand U1213 (N_1213,N_1172,N_1182);
and U1214 (N_1214,N_1168,N_1198);
nor U1215 (N_1215,N_1161,N_1176);
and U1216 (N_1216,N_1155,N_1173);
nor U1217 (N_1217,N_1187,N_1159);
nand U1218 (N_1218,N_1179,N_1165);
nor U1219 (N_1219,N_1186,N_1151);
and U1220 (N_1220,N_1190,N_1195);
or U1221 (N_1221,N_1154,N_1171);
nor U1222 (N_1222,N_1166,N_1196);
and U1223 (N_1223,N_1183,N_1164);
and U1224 (N_1224,N_1150,N_1177);
and U1225 (N_1225,N_1164,N_1170);
nor U1226 (N_1226,N_1152,N_1199);
or U1227 (N_1227,N_1189,N_1165);
xnor U1228 (N_1228,N_1162,N_1184);
nor U1229 (N_1229,N_1157,N_1158);
and U1230 (N_1230,N_1152,N_1165);
nor U1231 (N_1231,N_1182,N_1195);
xor U1232 (N_1232,N_1179,N_1168);
xor U1233 (N_1233,N_1174,N_1172);
xnor U1234 (N_1234,N_1168,N_1150);
nand U1235 (N_1235,N_1167,N_1190);
or U1236 (N_1236,N_1162,N_1168);
and U1237 (N_1237,N_1160,N_1150);
nand U1238 (N_1238,N_1170,N_1182);
nand U1239 (N_1239,N_1161,N_1172);
or U1240 (N_1240,N_1173,N_1187);
xor U1241 (N_1241,N_1195,N_1162);
nor U1242 (N_1242,N_1159,N_1195);
nor U1243 (N_1243,N_1178,N_1182);
nand U1244 (N_1244,N_1192,N_1185);
nor U1245 (N_1245,N_1154,N_1164);
or U1246 (N_1246,N_1179,N_1167);
and U1247 (N_1247,N_1176,N_1188);
and U1248 (N_1248,N_1154,N_1186);
and U1249 (N_1249,N_1160,N_1156);
nor U1250 (N_1250,N_1224,N_1249);
and U1251 (N_1251,N_1245,N_1246);
and U1252 (N_1252,N_1226,N_1209);
nand U1253 (N_1253,N_1221,N_1239);
nand U1254 (N_1254,N_1206,N_1208);
or U1255 (N_1255,N_1232,N_1200);
nor U1256 (N_1256,N_1205,N_1238);
nor U1257 (N_1257,N_1233,N_1247);
nand U1258 (N_1258,N_1230,N_1236);
or U1259 (N_1259,N_1222,N_1248);
or U1260 (N_1260,N_1214,N_1210);
xor U1261 (N_1261,N_1225,N_1213);
nor U1262 (N_1262,N_1229,N_1201);
or U1263 (N_1263,N_1223,N_1212);
and U1264 (N_1264,N_1237,N_1244);
or U1265 (N_1265,N_1240,N_1241);
nand U1266 (N_1266,N_1234,N_1231);
and U1267 (N_1267,N_1203,N_1217);
or U1268 (N_1268,N_1204,N_1220);
nand U1269 (N_1269,N_1207,N_1219);
or U1270 (N_1270,N_1227,N_1216);
nand U1271 (N_1271,N_1215,N_1228);
or U1272 (N_1272,N_1235,N_1242);
nor U1273 (N_1273,N_1211,N_1218);
nor U1274 (N_1274,N_1202,N_1243);
nor U1275 (N_1275,N_1200,N_1241);
and U1276 (N_1276,N_1214,N_1247);
nand U1277 (N_1277,N_1229,N_1238);
nor U1278 (N_1278,N_1242,N_1237);
nand U1279 (N_1279,N_1210,N_1208);
and U1280 (N_1280,N_1214,N_1228);
nor U1281 (N_1281,N_1217,N_1226);
or U1282 (N_1282,N_1212,N_1234);
and U1283 (N_1283,N_1218,N_1230);
or U1284 (N_1284,N_1218,N_1216);
nand U1285 (N_1285,N_1210,N_1202);
and U1286 (N_1286,N_1240,N_1210);
or U1287 (N_1287,N_1239,N_1207);
nand U1288 (N_1288,N_1227,N_1239);
and U1289 (N_1289,N_1235,N_1226);
xnor U1290 (N_1290,N_1243,N_1237);
xor U1291 (N_1291,N_1222,N_1217);
and U1292 (N_1292,N_1245,N_1205);
or U1293 (N_1293,N_1215,N_1211);
nor U1294 (N_1294,N_1226,N_1238);
or U1295 (N_1295,N_1223,N_1206);
and U1296 (N_1296,N_1228,N_1234);
or U1297 (N_1297,N_1203,N_1249);
and U1298 (N_1298,N_1240,N_1219);
nor U1299 (N_1299,N_1231,N_1205);
xor U1300 (N_1300,N_1252,N_1297);
or U1301 (N_1301,N_1274,N_1291);
xnor U1302 (N_1302,N_1251,N_1276);
or U1303 (N_1303,N_1283,N_1292);
xor U1304 (N_1304,N_1270,N_1260);
or U1305 (N_1305,N_1294,N_1269);
nor U1306 (N_1306,N_1277,N_1271);
nand U1307 (N_1307,N_1280,N_1273);
nor U1308 (N_1308,N_1262,N_1256);
nor U1309 (N_1309,N_1289,N_1288);
nor U1310 (N_1310,N_1287,N_1266);
or U1311 (N_1311,N_1253,N_1275);
and U1312 (N_1312,N_1257,N_1255);
nor U1313 (N_1313,N_1281,N_1261);
nor U1314 (N_1314,N_1250,N_1263);
or U1315 (N_1315,N_1265,N_1267);
and U1316 (N_1316,N_1264,N_1282);
nor U1317 (N_1317,N_1299,N_1279);
nor U1318 (N_1318,N_1286,N_1295);
xor U1319 (N_1319,N_1258,N_1278);
nand U1320 (N_1320,N_1285,N_1254);
or U1321 (N_1321,N_1259,N_1268);
nor U1322 (N_1322,N_1293,N_1272);
and U1323 (N_1323,N_1284,N_1296);
or U1324 (N_1324,N_1290,N_1298);
nand U1325 (N_1325,N_1281,N_1253);
or U1326 (N_1326,N_1298,N_1281);
and U1327 (N_1327,N_1285,N_1265);
nor U1328 (N_1328,N_1265,N_1264);
and U1329 (N_1329,N_1266,N_1289);
or U1330 (N_1330,N_1271,N_1298);
nand U1331 (N_1331,N_1259,N_1273);
nor U1332 (N_1332,N_1261,N_1277);
nand U1333 (N_1333,N_1294,N_1268);
nor U1334 (N_1334,N_1277,N_1259);
nor U1335 (N_1335,N_1284,N_1297);
nand U1336 (N_1336,N_1294,N_1276);
and U1337 (N_1337,N_1259,N_1260);
xnor U1338 (N_1338,N_1262,N_1277);
nor U1339 (N_1339,N_1272,N_1253);
or U1340 (N_1340,N_1281,N_1287);
xor U1341 (N_1341,N_1285,N_1290);
nor U1342 (N_1342,N_1269,N_1296);
xnor U1343 (N_1343,N_1296,N_1259);
and U1344 (N_1344,N_1298,N_1280);
nand U1345 (N_1345,N_1277,N_1252);
nor U1346 (N_1346,N_1287,N_1252);
and U1347 (N_1347,N_1250,N_1293);
or U1348 (N_1348,N_1268,N_1284);
or U1349 (N_1349,N_1284,N_1267);
xnor U1350 (N_1350,N_1349,N_1340);
and U1351 (N_1351,N_1331,N_1304);
xor U1352 (N_1352,N_1306,N_1330);
nand U1353 (N_1353,N_1329,N_1346);
nand U1354 (N_1354,N_1300,N_1302);
nand U1355 (N_1355,N_1303,N_1301);
or U1356 (N_1356,N_1337,N_1320);
or U1357 (N_1357,N_1324,N_1343);
and U1358 (N_1358,N_1310,N_1338);
and U1359 (N_1359,N_1328,N_1347);
and U1360 (N_1360,N_1305,N_1344);
and U1361 (N_1361,N_1341,N_1307);
xor U1362 (N_1362,N_1313,N_1326);
or U1363 (N_1363,N_1339,N_1323);
nand U1364 (N_1364,N_1333,N_1312);
nand U1365 (N_1365,N_1332,N_1318);
nor U1366 (N_1366,N_1348,N_1316);
nand U1367 (N_1367,N_1322,N_1311);
nand U1368 (N_1368,N_1327,N_1342);
nor U1369 (N_1369,N_1308,N_1336);
and U1370 (N_1370,N_1325,N_1315);
nor U1371 (N_1371,N_1309,N_1317);
or U1372 (N_1372,N_1319,N_1345);
nand U1373 (N_1373,N_1334,N_1321);
xnor U1374 (N_1374,N_1335,N_1314);
xnor U1375 (N_1375,N_1332,N_1347);
or U1376 (N_1376,N_1342,N_1325);
or U1377 (N_1377,N_1323,N_1328);
or U1378 (N_1378,N_1324,N_1311);
nand U1379 (N_1379,N_1317,N_1323);
nand U1380 (N_1380,N_1323,N_1313);
nand U1381 (N_1381,N_1346,N_1321);
and U1382 (N_1382,N_1322,N_1347);
and U1383 (N_1383,N_1331,N_1338);
and U1384 (N_1384,N_1308,N_1335);
nand U1385 (N_1385,N_1300,N_1338);
nand U1386 (N_1386,N_1313,N_1317);
nor U1387 (N_1387,N_1335,N_1324);
nand U1388 (N_1388,N_1300,N_1315);
nor U1389 (N_1389,N_1302,N_1310);
nor U1390 (N_1390,N_1323,N_1318);
nand U1391 (N_1391,N_1346,N_1347);
nand U1392 (N_1392,N_1321,N_1343);
or U1393 (N_1393,N_1320,N_1310);
xnor U1394 (N_1394,N_1303,N_1321);
or U1395 (N_1395,N_1346,N_1304);
nand U1396 (N_1396,N_1321,N_1324);
and U1397 (N_1397,N_1326,N_1318);
and U1398 (N_1398,N_1322,N_1306);
nor U1399 (N_1399,N_1349,N_1310);
and U1400 (N_1400,N_1352,N_1354);
or U1401 (N_1401,N_1359,N_1377);
and U1402 (N_1402,N_1397,N_1388);
or U1403 (N_1403,N_1394,N_1382);
or U1404 (N_1404,N_1358,N_1392);
or U1405 (N_1405,N_1351,N_1389);
or U1406 (N_1406,N_1391,N_1380);
nor U1407 (N_1407,N_1375,N_1361);
or U1408 (N_1408,N_1378,N_1395);
nor U1409 (N_1409,N_1387,N_1365);
or U1410 (N_1410,N_1364,N_1393);
or U1411 (N_1411,N_1363,N_1369);
xor U1412 (N_1412,N_1353,N_1370);
or U1413 (N_1413,N_1350,N_1376);
and U1414 (N_1414,N_1367,N_1396);
nor U1415 (N_1415,N_1383,N_1373);
xor U1416 (N_1416,N_1385,N_1355);
and U1417 (N_1417,N_1374,N_1357);
nor U1418 (N_1418,N_1362,N_1371);
nor U1419 (N_1419,N_1360,N_1381);
nand U1420 (N_1420,N_1386,N_1368);
and U1421 (N_1421,N_1379,N_1390);
or U1422 (N_1422,N_1398,N_1356);
and U1423 (N_1423,N_1399,N_1366);
nand U1424 (N_1424,N_1372,N_1384);
nand U1425 (N_1425,N_1394,N_1351);
or U1426 (N_1426,N_1375,N_1350);
and U1427 (N_1427,N_1373,N_1350);
and U1428 (N_1428,N_1397,N_1363);
xnor U1429 (N_1429,N_1363,N_1378);
nor U1430 (N_1430,N_1395,N_1353);
nand U1431 (N_1431,N_1364,N_1362);
nor U1432 (N_1432,N_1383,N_1382);
nand U1433 (N_1433,N_1373,N_1396);
or U1434 (N_1434,N_1361,N_1350);
nand U1435 (N_1435,N_1362,N_1350);
or U1436 (N_1436,N_1394,N_1396);
or U1437 (N_1437,N_1386,N_1357);
or U1438 (N_1438,N_1365,N_1355);
and U1439 (N_1439,N_1360,N_1373);
or U1440 (N_1440,N_1358,N_1372);
nor U1441 (N_1441,N_1388,N_1396);
xor U1442 (N_1442,N_1358,N_1366);
nand U1443 (N_1443,N_1357,N_1353);
and U1444 (N_1444,N_1399,N_1387);
nand U1445 (N_1445,N_1397,N_1374);
nand U1446 (N_1446,N_1385,N_1366);
nand U1447 (N_1447,N_1391,N_1359);
and U1448 (N_1448,N_1355,N_1392);
nor U1449 (N_1449,N_1364,N_1390);
nand U1450 (N_1450,N_1411,N_1435);
nand U1451 (N_1451,N_1417,N_1414);
nor U1452 (N_1452,N_1401,N_1443);
nor U1453 (N_1453,N_1428,N_1405);
nand U1454 (N_1454,N_1409,N_1400);
nor U1455 (N_1455,N_1441,N_1430);
nor U1456 (N_1456,N_1406,N_1426);
nor U1457 (N_1457,N_1437,N_1404);
nand U1458 (N_1458,N_1449,N_1412);
and U1459 (N_1459,N_1416,N_1429);
nand U1460 (N_1460,N_1423,N_1440);
or U1461 (N_1461,N_1424,N_1420);
xnor U1462 (N_1462,N_1444,N_1407);
nand U1463 (N_1463,N_1445,N_1415);
xor U1464 (N_1464,N_1438,N_1447);
nand U1465 (N_1465,N_1403,N_1421);
or U1466 (N_1466,N_1446,N_1427);
and U1467 (N_1467,N_1434,N_1413);
xnor U1468 (N_1468,N_1408,N_1433);
or U1469 (N_1469,N_1439,N_1448);
or U1470 (N_1470,N_1422,N_1410);
nand U1471 (N_1471,N_1436,N_1431);
xor U1472 (N_1472,N_1442,N_1418);
and U1473 (N_1473,N_1432,N_1419);
nor U1474 (N_1474,N_1402,N_1425);
or U1475 (N_1475,N_1407,N_1419);
xnor U1476 (N_1476,N_1417,N_1419);
nor U1477 (N_1477,N_1434,N_1438);
or U1478 (N_1478,N_1441,N_1414);
or U1479 (N_1479,N_1414,N_1447);
and U1480 (N_1480,N_1429,N_1435);
nor U1481 (N_1481,N_1403,N_1411);
or U1482 (N_1482,N_1441,N_1410);
and U1483 (N_1483,N_1443,N_1439);
nor U1484 (N_1484,N_1426,N_1420);
xor U1485 (N_1485,N_1420,N_1410);
nand U1486 (N_1486,N_1404,N_1403);
or U1487 (N_1487,N_1426,N_1422);
or U1488 (N_1488,N_1416,N_1424);
nor U1489 (N_1489,N_1443,N_1414);
or U1490 (N_1490,N_1443,N_1404);
and U1491 (N_1491,N_1432,N_1448);
nor U1492 (N_1492,N_1424,N_1425);
and U1493 (N_1493,N_1403,N_1434);
nor U1494 (N_1494,N_1426,N_1438);
or U1495 (N_1495,N_1413,N_1446);
nor U1496 (N_1496,N_1432,N_1412);
nand U1497 (N_1497,N_1440,N_1421);
nor U1498 (N_1498,N_1445,N_1416);
nor U1499 (N_1499,N_1431,N_1401);
or U1500 (N_1500,N_1459,N_1462);
or U1501 (N_1501,N_1497,N_1457);
and U1502 (N_1502,N_1493,N_1486);
and U1503 (N_1503,N_1468,N_1481);
or U1504 (N_1504,N_1499,N_1464);
and U1505 (N_1505,N_1478,N_1488);
or U1506 (N_1506,N_1492,N_1466);
or U1507 (N_1507,N_1470,N_1463);
nor U1508 (N_1508,N_1451,N_1460);
or U1509 (N_1509,N_1474,N_1467);
nand U1510 (N_1510,N_1453,N_1482);
and U1511 (N_1511,N_1498,N_1469);
and U1512 (N_1512,N_1465,N_1484);
xnor U1513 (N_1513,N_1483,N_1458);
nand U1514 (N_1514,N_1495,N_1477);
xnor U1515 (N_1515,N_1485,N_1450);
or U1516 (N_1516,N_1455,N_1454);
or U1517 (N_1517,N_1479,N_1491);
nor U1518 (N_1518,N_1496,N_1490);
and U1519 (N_1519,N_1480,N_1473);
xor U1520 (N_1520,N_1487,N_1472);
or U1521 (N_1521,N_1494,N_1476);
xnor U1522 (N_1522,N_1456,N_1452);
nand U1523 (N_1523,N_1471,N_1475);
and U1524 (N_1524,N_1461,N_1489);
and U1525 (N_1525,N_1499,N_1476);
xnor U1526 (N_1526,N_1464,N_1472);
nor U1527 (N_1527,N_1497,N_1486);
and U1528 (N_1528,N_1482,N_1464);
nand U1529 (N_1529,N_1490,N_1482);
nor U1530 (N_1530,N_1495,N_1481);
nand U1531 (N_1531,N_1471,N_1458);
or U1532 (N_1532,N_1494,N_1484);
nor U1533 (N_1533,N_1492,N_1493);
and U1534 (N_1534,N_1454,N_1476);
and U1535 (N_1535,N_1491,N_1498);
or U1536 (N_1536,N_1492,N_1470);
or U1537 (N_1537,N_1460,N_1457);
and U1538 (N_1538,N_1494,N_1474);
xnor U1539 (N_1539,N_1475,N_1487);
nand U1540 (N_1540,N_1484,N_1460);
and U1541 (N_1541,N_1466,N_1459);
and U1542 (N_1542,N_1486,N_1480);
nand U1543 (N_1543,N_1451,N_1476);
or U1544 (N_1544,N_1496,N_1491);
nor U1545 (N_1545,N_1460,N_1489);
and U1546 (N_1546,N_1488,N_1490);
and U1547 (N_1547,N_1498,N_1489);
xnor U1548 (N_1548,N_1492,N_1471);
nor U1549 (N_1549,N_1492,N_1476);
and U1550 (N_1550,N_1533,N_1508);
nor U1551 (N_1551,N_1538,N_1536);
xnor U1552 (N_1552,N_1520,N_1545);
nand U1553 (N_1553,N_1544,N_1525);
or U1554 (N_1554,N_1511,N_1505);
nand U1555 (N_1555,N_1506,N_1528);
or U1556 (N_1556,N_1530,N_1543);
and U1557 (N_1557,N_1523,N_1503);
and U1558 (N_1558,N_1531,N_1534);
nand U1559 (N_1559,N_1542,N_1501);
xor U1560 (N_1560,N_1513,N_1541);
nand U1561 (N_1561,N_1507,N_1504);
and U1562 (N_1562,N_1539,N_1535);
nor U1563 (N_1563,N_1510,N_1502);
and U1564 (N_1564,N_1519,N_1516);
and U1565 (N_1565,N_1529,N_1524);
and U1566 (N_1566,N_1548,N_1526);
and U1567 (N_1567,N_1521,N_1500);
nand U1568 (N_1568,N_1512,N_1515);
nand U1569 (N_1569,N_1547,N_1514);
xnor U1570 (N_1570,N_1522,N_1527);
and U1571 (N_1571,N_1549,N_1532);
nand U1572 (N_1572,N_1537,N_1517);
nor U1573 (N_1573,N_1540,N_1546);
or U1574 (N_1574,N_1518,N_1509);
or U1575 (N_1575,N_1502,N_1543);
nor U1576 (N_1576,N_1506,N_1524);
or U1577 (N_1577,N_1513,N_1532);
nand U1578 (N_1578,N_1543,N_1547);
nor U1579 (N_1579,N_1546,N_1510);
xnor U1580 (N_1580,N_1542,N_1500);
xor U1581 (N_1581,N_1530,N_1520);
and U1582 (N_1582,N_1526,N_1521);
or U1583 (N_1583,N_1514,N_1528);
nor U1584 (N_1584,N_1534,N_1507);
xnor U1585 (N_1585,N_1523,N_1513);
and U1586 (N_1586,N_1520,N_1517);
or U1587 (N_1587,N_1540,N_1503);
xor U1588 (N_1588,N_1520,N_1549);
nand U1589 (N_1589,N_1511,N_1539);
nor U1590 (N_1590,N_1510,N_1500);
nand U1591 (N_1591,N_1514,N_1507);
and U1592 (N_1592,N_1502,N_1524);
and U1593 (N_1593,N_1530,N_1531);
xnor U1594 (N_1594,N_1531,N_1512);
or U1595 (N_1595,N_1537,N_1508);
nand U1596 (N_1596,N_1528,N_1535);
and U1597 (N_1597,N_1512,N_1504);
nor U1598 (N_1598,N_1547,N_1520);
or U1599 (N_1599,N_1518,N_1534);
or U1600 (N_1600,N_1583,N_1570);
nand U1601 (N_1601,N_1599,N_1594);
or U1602 (N_1602,N_1567,N_1559);
or U1603 (N_1603,N_1550,N_1565);
xor U1604 (N_1604,N_1577,N_1578);
nand U1605 (N_1605,N_1596,N_1584);
or U1606 (N_1606,N_1572,N_1566);
and U1607 (N_1607,N_1576,N_1580);
and U1608 (N_1608,N_1564,N_1569);
and U1609 (N_1609,N_1597,N_1553);
nor U1610 (N_1610,N_1561,N_1555);
and U1611 (N_1611,N_1551,N_1589);
or U1612 (N_1612,N_1593,N_1557);
and U1613 (N_1613,N_1563,N_1554);
nor U1614 (N_1614,N_1558,N_1574);
nor U1615 (N_1615,N_1575,N_1560);
nand U1616 (N_1616,N_1588,N_1591);
nor U1617 (N_1617,N_1582,N_1598);
and U1618 (N_1618,N_1552,N_1568);
nor U1619 (N_1619,N_1587,N_1579);
nor U1620 (N_1620,N_1595,N_1590);
nand U1621 (N_1621,N_1586,N_1581);
xnor U1622 (N_1622,N_1562,N_1573);
or U1623 (N_1623,N_1556,N_1571);
nor U1624 (N_1624,N_1585,N_1592);
or U1625 (N_1625,N_1584,N_1563);
or U1626 (N_1626,N_1584,N_1591);
or U1627 (N_1627,N_1598,N_1553);
nand U1628 (N_1628,N_1599,N_1557);
or U1629 (N_1629,N_1584,N_1574);
xnor U1630 (N_1630,N_1581,N_1599);
and U1631 (N_1631,N_1594,N_1577);
nor U1632 (N_1632,N_1555,N_1557);
and U1633 (N_1633,N_1578,N_1559);
and U1634 (N_1634,N_1579,N_1552);
nor U1635 (N_1635,N_1590,N_1574);
or U1636 (N_1636,N_1560,N_1576);
or U1637 (N_1637,N_1576,N_1574);
or U1638 (N_1638,N_1594,N_1579);
or U1639 (N_1639,N_1575,N_1586);
nor U1640 (N_1640,N_1577,N_1595);
and U1641 (N_1641,N_1588,N_1596);
nand U1642 (N_1642,N_1597,N_1589);
or U1643 (N_1643,N_1563,N_1558);
or U1644 (N_1644,N_1579,N_1592);
and U1645 (N_1645,N_1595,N_1589);
or U1646 (N_1646,N_1559,N_1585);
nor U1647 (N_1647,N_1570,N_1555);
nand U1648 (N_1648,N_1596,N_1572);
xnor U1649 (N_1649,N_1582,N_1591);
xnor U1650 (N_1650,N_1631,N_1621);
and U1651 (N_1651,N_1622,N_1613);
nor U1652 (N_1652,N_1610,N_1644);
nor U1653 (N_1653,N_1643,N_1627);
nand U1654 (N_1654,N_1602,N_1639);
or U1655 (N_1655,N_1600,N_1633);
nor U1656 (N_1656,N_1606,N_1635);
and U1657 (N_1657,N_1634,N_1620);
nor U1658 (N_1658,N_1628,N_1624);
xor U1659 (N_1659,N_1618,N_1632);
xor U1660 (N_1660,N_1607,N_1625);
xor U1661 (N_1661,N_1649,N_1647);
nor U1662 (N_1662,N_1638,N_1603);
and U1663 (N_1663,N_1616,N_1629);
nand U1664 (N_1664,N_1614,N_1605);
or U1665 (N_1665,N_1630,N_1642);
nor U1666 (N_1666,N_1636,N_1646);
nand U1667 (N_1667,N_1645,N_1619);
or U1668 (N_1668,N_1612,N_1641);
and U1669 (N_1669,N_1626,N_1617);
nor U1670 (N_1670,N_1611,N_1637);
nor U1671 (N_1671,N_1615,N_1640);
or U1672 (N_1672,N_1608,N_1609);
and U1673 (N_1673,N_1623,N_1604);
and U1674 (N_1674,N_1601,N_1648);
xor U1675 (N_1675,N_1635,N_1622);
and U1676 (N_1676,N_1612,N_1638);
nor U1677 (N_1677,N_1630,N_1629);
nand U1678 (N_1678,N_1604,N_1627);
xnor U1679 (N_1679,N_1606,N_1649);
nor U1680 (N_1680,N_1640,N_1621);
nand U1681 (N_1681,N_1639,N_1621);
and U1682 (N_1682,N_1611,N_1618);
or U1683 (N_1683,N_1645,N_1639);
or U1684 (N_1684,N_1604,N_1643);
xnor U1685 (N_1685,N_1649,N_1633);
or U1686 (N_1686,N_1629,N_1602);
nor U1687 (N_1687,N_1601,N_1610);
or U1688 (N_1688,N_1612,N_1632);
xnor U1689 (N_1689,N_1612,N_1643);
or U1690 (N_1690,N_1649,N_1641);
nor U1691 (N_1691,N_1615,N_1633);
nand U1692 (N_1692,N_1622,N_1632);
and U1693 (N_1693,N_1620,N_1629);
nand U1694 (N_1694,N_1617,N_1635);
nand U1695 (N_1695,N_1629,N_1623);
and U1696 (N_1696,N_1612,N_1600);
nor U1697 (N_1697,N_1605,N_1639);
and U1698 (N_1698,N_1614,N_1623);
and U1699 (N_1699,N_1605,N_1612);
nor U1700 (N_1700,N_1675,N_1650);
nand U1701 (N_1701,N_1687,N_1654);
nand U1702 (N_1702,N_1652,N_1676);
nor U1703 (N_1703,N_1699,N_1661);
nor U1704 (N_1704,N_1666,N_1653);
or U1705 (N_1705,N_1656,N_1669);
nand U1706 (N_1706,N_1668,N_1697);
nand U1707 (N_1707,N_1677,N_1664);
and U1708 (N_1708,N_1655,N_1671);
nand U1709 (N_1709,N_1688,N_1698);
nand U1710 (N_1710,N_1667,N_1663);
and U1711 (N_1711,N_1651,N_1696);
or U1712 (N_1712,N_1672,N_1673);
nand U1713 (N_1713,N_1691,N_1686);
or U1714 (N_1714,N_1693,N_1685);
or U1715 (N_1715,N_1659,N_1670);
xnor U1716 (N_1716,N_1689,N_1694);
xor U1717 (N_1717,N_1665,N_1692);
nor U1718 (N_1718,N_1684,N_1674);
or U1719 (N_1719,N_1680,N_1657);
or U1720 (N_1720,N_1678,N_1690);
nand U1721 (N_1721,N_1658,N_1683);
and U1722 (N_1722,N_1679,N_1682);
and U1723 (N_1723,N_1662,N_1695);
nand U1724 (N_1724,N_1660,N_1681);
nor U1725 (N_1725,N_1654,N_1657);
nor U1726 (N_1726,N_1691,N_1657);
nor U1727 (N_1727,N_1684,N_1679);
and U1728 (N_1728,N_1690,N_1697);
or U1729 (N_1729,N_1670,N_1672);
nand U1730 (N_1730,N_1661,N_1673);
nor U1731 (N_1731,N_1675,N_1688);
nand U1732 (N_1732,N_1657,N_1683);
and U1733 (N_1733,N_1697,N_1684);
or U1734 (N_1734,N_1657,N_1658);
nand U1735 (N_1735,N_1653,N_1651);
nor U1736 (N_1736,N_1653,N_1685);
nor U1737 (N_1737,N_1677,N_1650);
nand U1738 (N_1738,N_1667,N_1677);
nand U1739 (N_1739,N_1665,N_1688);
or U1740 (N_1740,N_1668,N_1695);
nand U1741 (N_1741,N_1695,N_1660);
or U1742 (N_1742,N_1662,N_1658);
nand U1743 (N_1743,N_1673,N_1658);
nand U1744 (N_1744,N_1659,N_1663);
xor U1745 (N_1745,N_1677,N_1698);
nor U1746 (N_1746,N_1660,N_1680);
or U1747 (N_1747,N_1677,N_1697);
and U1748 (N_1748,N_1684,N_1666);
nor U1749 (N_1749,N_1653,N_1663);
nor U1750 (N_1750,N_1746,N_1744);
or U1751 (N_1751,N_1707,N_1730);
nor U1752 (N_1752,N_1700,N_1733);
or U1753 (N_1753,N_1711,N_1710);
or U1754 (N_1754,N_1731,N_1708);
nand U1755 (N_1755,N_1738,N_1737);
nor U1756 (N_1756,N_1713,N_1705);
and U1757 (N_1757,N_1715,N_1709);
nand U1758 (N_1758,N_1743,N_1742);
nor U1759 (N_1759,N_1734,N_1712);
and U1760 (N_1760,N_1703,N_1741);
nor U1761 (N_1761,N_1719,N_1716);
nand U1762 (N_1762,N_1740,N_1736);
and U1763 (N_1763,N_1749,N_1728);
nor U1764 (N_1764,N_1717,N_1732);
or U1765 (N_1765,N_1701,N_1722);
nor U1766 (N_1766,N_1727,N_1745);
nor U1767 (N_1767,N_1739,N_1723);
nor U1768 (N_1768,N_1725,N_1748);
and U1769 (N_1769,N_1702,N_1735);
or U1770 (N_1770,N_1704,N_1729);
and U1771 (N_1771,N_1724,N_1718);
and U1772 (N_1772,N_1747,N_1706);
and U1773 (N_1773,N_1720,N_1726);
or U1774 (N_1774,N_1714,N_1721);
xor U1775 (N_1775,N_1708,N_1729);
or U1776 (N_1776,N_1743,N_1720);
or U1777 (N_1777,N_1731,N_1730);
nand U1778 (N_1778,N_1706,N_1705);
and U1779 (N_1779,N_1733,N_1748);
or U1780 (N_1780,N_1706,N_1717);
nor U1781 (N_1781,N_1732,N_1733);
and U1782 (N_1782,N_1719,N_1727);
and U1783 (N_1783,N_1733,N_1738);
nor U1784 (N_1784,N_1712,N_1702);
xnor U1785 (N_1785,N_1731,N_1733);
nand U1786 (N_1786,N_1720,N_1703);
or U1787 (N_1787,N_1728,N_1724);
or U1788 (N_1788,N_1731,N_1711);
nor U1789 (N_1789,N_1748,N_1714);
and U1790 (N_1790,N_1739,N_1702);
or U1791 (N_1791,N_1740,N_1749);
and U1792 (N_1792,N_1729,N_1734);
or U1793 (N_1793,N_1737,N_1731);
nor U1794 (N_1794,N_1723,N_1731);
or U1795 (N_1795,N_1724,N_1704);
nand U1796 (N_1796,N_1722,N_1702);
nor U1797 (N_1797,N_1716,N_1738);
and U1798 (N_1798,N_1722,N_1720);
nor U1799 (N_1799,N_1721,N_1700);
and U1800 (N_1800,N_1779,N_1784);
xnor U1801 (N_1801,N_1774,N_1771);
and U1802 (N_1802,N_1789,N_1782);
nand U1803 (N_1803,N_1787,N_1790);
nand U1804 (N_1804,N_1751,N_1770);
nand U1805 (N_1805,N_1781,N_1799);
nor U1806 (N_1806,N_1794,N_1793);
nor U1807 (N_1807,N_1785,N_1754);
nand U1808 (N_1808,N_1762,N_1768);
nor U1809 (N_1809,N_1760,N_1783);
nor U1810 (N_1810,N_1788,N_1776);
nor U1811 (N_1811,N_1758,N_1766);
and U1812 (N_1812,N_1753,N_1769);
nand U1813 (N_1813,N_1752,N_1764);
nand U1814 (N_1814,N_1798,N_1767);
nor U1815 (N_1815,N_1791,N_1755);
xor U1816 (N_1816,N_1763,N_1780);
nand U1817 (N_1817,N_1778,N_1792);
or U1818 (N_1818,N_1795,N_1761);
nor U1819 (N_1819,N_1765,N_1756);
nand U1820 (N_1820,N_1757,N_1773);
and U1821 (N_1821,N_1772,N_1796);
nand U1822 (N_1822,N_1786,N_1750);
or U1823 (N_1823,N_1759,N_1797);
nor U1824 (N_1824,N_1775,N_1777);
and U1825 (N_1825,N_1763,N_1760);
nand U1826 (N_1826,N_1781,N_1771);
xnor U1827 (N_1827,N_1763,N_1753);
or U1828 (N_1828,N_1755,N_1762);
xnor U1829 (N_1829,N_1754,N_1765);
nor U1830 (N_1830,N_1772,N_1786);
nand U1831 (N_1831,N_1759,N_1782);
nand U1832 (N_1832,N_1751,N_1790);
nand U1833 (N_1833,N_1773,N_1772);
nor U1834 (N_1834,N_1769,N_1789);
nand U1835 (N_1835,N_1772,N_1769);
xor U1836 (N_1836,N_1799,N_1784);
or U1837 (N_1837,N_1787,N_1776);
and U1838 (N_1838,N_1756,N_1784);
nand U1839 (N_1839,N_1761,N_1771);
or U1840 (N_1840,N_1777,N_1795);
or U1841 (N_1841,N_1760,N_1754);
nor U1842 (N_1842,N_1783,N_1750);
and U1843 (N_1843,N_1790,N_1762);
nor U1844 (N_1844,N_1767,N_1780);
or U1845 (N_1845,N_1760,N_1780);
nor U1846 (N_1846,N_1755,N_1785);
nor U1847 (N_1847,N_1757,N_1798);
and U1848 (N_1848,N_1788,N_1798);
or U1849 (N_1849,N_1795,N_1772);
nor U1850 (N_1850,N_1833,N_1809);
and U1851 (N_1851,N_1816,N_1840);
and U1852 (N_1852,N_1845,N_1813);
nand U1853 (N_1853,N_1801,N_1836);
and U1854 (N_1854,N_1846,N_1824);
nand U1855 (N_1855,N_1822,N_1832);
nor U1856 (N_1856,N_1821,N_1826);
or U1857 (N_1857,N_1819,N_1835);
and U1858 (N_1858,N_1815,N_1841);
nor U1859 (N_1859,N_1839,N_1827);
and U1860 (N_1860,N_1817,N_1802);
and U1861 (N_1861,N_1811,N_1834);
and U1862 (N_1862,N_1812,N_1847);
and U1863 (N_1863,N_1800,N_1825);
xor U1864 (N_1864,N_1803,N_1848);
nand U1865 (N_1865,N_1823,N_1829);
or U1866 (N_1866,N_1810,N_1820);
nand U1867 (N_1867,N_1818,N_1830);
or U1868 (N_1868,N_1805,N_1804);
or U1869 (N_1869,N_1843,N_1837);
and U1870 (N_1870,N_1838,N_1806);
nand U1871 (N_1871,N_1849,N_1814);
nand U1872 (N_1872,N_1808,N_1831);
nor U1873 (N_1873,N_1828,N_1842);
nor U1874 (N_1874,N_1807,N_1844);
and U1875 (N_1875,N_1827,N_1801);
and U1876 (N_1876,N_1803,N_1815);
nand U1877 (N_1877,N_1821,N_1835);
nor U1878 (N_1878,N_1803,N_1836);
nand U1879 (N_1879,N_1805,N_1842);
and U1880 (N_1880,N_1833,N_1834);
and U1881 (N_1881,N_1806,N_1849);
xnor U1882 (N_1882,N_1803,N_1800);
nand U1883 (N_1883,N_1802,N_1839);
nor U1884 (N_1884,N_1823,N_1846);
and U1885 (N_1885,N_1833,N_1846);
or U1886 (N_1886,N_1842,N_1848);
nand U1887 (N_1887,N_1812,N_1828);
xor U1888 (N_1888,N_1808,N_1811);
or U1889 (N_1889,N_1840,N_1849);
and U1890 (N_1890,N_1807,N_1808);
or U1891 (N_1891,N_1822,N_1844);
or U1892 (N_1892,N_1804,N_1835);
and U1893 (N_1893,N_1821,N_1804);
nand U1894 (N_1894,N_1835,N_1809);
and U1895 (N_1895,N_1803,N_1825);
and U1896 (N_1896,N_1801,N_1848);
nand U1897 (N_1897,N_1806,N_1825);
and U1898 (N_1898,N_1844,N_1821);
nor U1899 (N_1899,N_1803,N_1830);
and U1900 (N_1900,N_1861,N_1858);
or U1901 (N_1901,N_1876,N_1890);
and U1902 (N_1902,N_1898,N_1882);
nand U1903 (N_1903,N_1888,N_1862);
xnor U1904 (N_1904,N_1854,N_1850);
nand U1905 (N_1905,N_1892,N_1870);
or U1906 (N_1906,N_1885,N_1875);
or U1907 (N_1907,N_1879,N_1868);
or U1908 (N_1908,N_1897,N_1859);
and U1909 (N_1909,N_1884,N_1889);
or U1910 (N_1910,N_1872,N_1863);
and U1911 (N_1911,N_1865,N_1877);
and U1912 (N_1912,N_1873,N_1855);
and U1913 (N_1913,N_1893,N_1874);
or U1914 (N_1914,N_1851,N_1894);
or U1915 (N_1915,N_1871,N_1886);
or U1916 (N_1916,N_1896,N_1864);
and U1917 (N_1917,N_1883,N_1878);
or U1918 (N_1918,N_1891,N_1860);
nor U1919 (N_1919,N_1881,N_1866);
and U1920 (N_1920,N_1880,N_1857);
or U1921 (N_1921,N_1867,N_1852);
nor U1922 (N_1922,N_1856,N_1895);
nand U1923 (N_1923,N_1899,N_1869);
nand U1924 (N_1924,N_1887,N_1853);
or U1925 (N_1925,N_1861,N_1868);
xnor U1926 (N_1926,N_1864,N_1883);
nor U1927 (N_1927,N_1895,N_1884);
nor U1928 (N_1928,N_1890,N_1874);
or U1929 (N_1929,N_1867,N_1865);
or U1930 (N_1930,N_1858,N_1867);
and U1931 (N_1931,N_1877,N_1869);
and U1932 (N_1932,N_1890,N_1881);
nor U1933 (N_1933,N_1864,N_1878);
or U1934 (N_1934,N_1890,N_1889);
and U1935 (N_1935,N_1873,N_1883);
nor U1936 (N_1936,N_1894,N_1876);
nor U1937 (N_1937,N_1868,N_1886);
or U1938 (N_1938,N_1863,N_1860);
nor U1939 (N_1939,N_1898,N_1859);
or U1940 (N_1940,N_1854,N_1855);
and U1941 (N_1941,N_1854,N_1883);
and U1942 (N_1942,N_1890,N_1894);
or U1943 (N_1943,N_1858,N_1894);
xor U1944 (N_1944,N_1859,N_1886);
nor U1945 (N_1945,N_1859,N_1899);
nand U1946 (N_1946,N_1869,N_1865);
nand U1947 (N_1947,N_1891,N_1872);
nor U1948 (N_1948,N_1881,N_1879);
and U1949 (N_1949,N_1879,N_1899);
nand U1950 (N_1950,N_1905,N_1928);
nand U1951 (N_1951,N_1947,N_1931);
or U1952 (N_1952,N_1925,N_1915);
or U1953 (N_1953,N_1913,N_1901);
nand U1954 (N_1954,N_1924,N_1939);
or U1955 (N_1955,N_1923,N_1903);
xnor U1956 (N_1956,N_1910,N_1922);
and U1957 (N_1957,N_1934,N_1941);
or U1958 (N_1958,N_1926,N_1908);
or U1959 (N_1959,N_1937,N_1929);
or U1960 (N_1960,N_1919,N_1940);
xnor U1961 (N_1961,N_1932,N_1945);
nand U1962 (N_1962,N_1906,N_1911);
nand U1963 (N_1963,N_1943,N_1909);
nand U1964 (N_1964,N_1907,N_1918);
nor U1965 (N_1965,N_1935,N_1936);
or U1966 (N_1966,N_1946,N_1944);
and U1967 (N_1967,N_1914,N_1930);
or U1968 (N_1968,N_1948,N_1933);
nand U1969 (N_1969,N_1902,N_1927);
and U1970 (N_1970,N_1912,N_1904);
nor U1971 (N_1971,N_1938,N_1942);
nand U1972 (N_1972,N_1949,N_1917);
and U1973 (N_1973,N_1921,N_1920);
or U1974 (N_1974,N_1900,N_1916);
nand U1975 (N_1975,N_1939,N_1929);
or U1976 (N_1976,N_1932,N_1902);
and U1977 (N_1977,N_1905,N_1909);
or U1978 (N_1978,N_1907,N_1915);
nand U1979 (N_1979,N_1909,N_1917);
and U1980 (N_1980,N_1901,N_1909);
nor U1981 (N_1981,N_1910,N_1900);
or U1982 (N_1982,N_1943,N_1927);
nand U1983 (N_1983,N_1912,N_1930);
and U1984 (N_1984,N_1917,N_1938);
xnor U1985 (N_1985,N_1927,N_1923);
and U1986 (N_1986,N_1911,N_1919);
and U1987 (N_1987,N_1921,N_1922);
or U1988 (N_1988,N_1915,N_1944);
nor U1989 (N_1989,N_1902,N_1906);
and U1990 (N_1990,N_1925,N_1943);
and U1991 (N_1991,N_1947,N_1916);
or U1992 (N_1992,N_1942,N_1924);
nor U1993 (N_1993,N_1936,N_1902);
or U1994 (N_1994,N_1906,N_1931);
nand U1995 (N_1995,N_1901,N_1946);
nand U1996 (N_1996,N_1906,N_1913);
nor U1997 (N_1997,N_1923,N_1911);
xnor U1998 (N_1998,N_1944,N_1928);
nor U1999 (N_1999,N_1913,N_1910);
nor U2000 (N_2000,N_1988,N_1957);
nand U2001 (N_2001,N_1995,N_1951);
and U2002 (N_2002,N_1961,N_1982);
and U2003 (N_2003,N_1998,N_1977);
nor U2004 (N_2004,N_1990,N_1967);
or U2005 (N_2005,N_1978,N_1980);
or U2006 (N_2006,N_1973,N_1972);
and U2007 (N_2007,N_1976,N_1987);
or U2008 (N_2008,N_1962,N_1991);
xor U2009 (N_2009,N_1992,N_1999);
nand U2010 (N_2010,N_1952,N_1958);
or U2011 (N_2011,N_1983,N_1971);
or U2012 (N_2012,N_1989,N_1966);
or U2013 (N_2013,N_1963,N_1956);
or U2014 (N_2014,N_1959,N_1996);
nor U2015 (N_2015,N_1997,N_1974);
or U2016 (N_2016,N_1985,N_1984);
or U2017 (N_2017,N_1993,N_1981);
nor U2018 (N_2018,N_1994,N_1979);
nor U2019 (N_2019,N_1965,N_1953);
or U2020 (N_2020,N_1986,N_1964);
xor U2021 (N_2021,N_1954,N_1955);
or U2022 (N_2022,N_1968,N_1975);
nor U2023 (N_2023,N_1969,N_1950);
and U2024 (N_2024,N_1960,N_1970);
and U2025 (N_2025,N_1951,N_1953);
nor U2026 (N_2026,N_1980,N_1985);
and U2027 (N_2027,N_1997,N_1973);
nand U2028 (N_2028,N_1955,N_1961);
and U2029 (N_2029,N_1954,N_1998);
nand U2030 (N_2030,N_1998,N_1950);
or U2031 (N_2031,N_1987,N_1962);
nand U2032 (N_2032,N_1986,N_1969);
xnor U2033 (N_2033,N_1981,N_1986);
and U2034 (N_2034,N_1958,N_1977);
nor U2035 (N_2035,N_1983,N_1974);
xor U2036 (N_2036,N_1989,N_1976);
xnor U2037 (N_2037,N_1959,N_1994);
nand U2038 (N_2038,N_1998,N_1971);
nand U2039 (N_2039,N_1969,N_1993);
xor U2040 (N_2040,N_1955,N_1974);
or U2041 (N_2041,N_1981,N_1985);
or U2042 (N_2042,N_1997,N_1955);
nand U2043 (N_2043,N_1968,N_1988);
nor U2044 (N_2044,N_1976,N_1993);
nand U2045 (N_2045,N_1954,N_1966);
nand U2046 (N_2046,N_1964,N_1997);
nor U2047 (N_2047,N_1991,N_1958);
nor U2048 (N_2048,N_1962,N_1955);
nor U2049 (N_2049,N_1964,N_1966);
or U2050 (N_2050,N_2008,N_2036);
nand U2051 (N_2051,N_2045,N_2019);
xor U2052 (N_2052,N_2046,N_2012);
or U2053 (N_2053,N_2032,N_2021);
and U2054 (N_2054,N_2009,N_2033);
and U2055 (N_2055,N_2017,N_2040);
xor U2056 (N_2056,N_2001,N_2037);
and U2057 (N_2057,N_2005,N_2024);
nand U2058 (N_2058,N_2042,N_2010);
and U2059 (N_2059,N_2011,N_2006);
nor U2060 (N_2060,N_2003,N_2029);
or U2061 (N_2061,N_2025,N_2022);
and U2062 (N_2062,N_2002,N_2014);
nand U2063 (N_2063,N_2030,N_2035);
nand U2064 (N_2064,N_2041,N_2007);
nand U2065 (N_2065,N_2026,N_2020);
nand U2066 (N_2066,N_2018,N_2031);
nor U2067 (N_2067,N_2023,N_2049);
and U2068 (N_2068,N_2016,N_2004);
nor U2069 (N_2069,N_2048,N_2027);
nor U2070 (N_2070,N_2000,N_2034);
nand U2071 (N_2071,N_2044,N_2015);
or U2072 (N_2072,N_2039,N_2043);
xor U2073 (N_2073,N_2028,N_2038);
nor U2074 (N_2074,N_2047,N_2013);
nor U2075 (N_2075,N_2003,N_2018);
or U2076 (N_2076,N_2003,N_2021);
nor U2077 (N_2077,N_2029,N_2019);
nand U2078 (N_2078,N_2019,N_2011);
and U2079 (N_2079,N_2032,N_2039);
or U2080 (N_2080,N_2028,N_2030);
nor U2081 (N_2081,N_2021,N_2016);
nor U2082 (N_2082,N_2024,N_2023);
or U2083 (N_2083,N_2013,N_2044);
and U2084 (N_2084,N_2034,N_2042);
or U2085 (N_2085,N_2024,N_2038);
nor U2086 (N_2086,N_2004,N_2021);
nor U2087 (N_2087,N_2044,N_2008);
nor U2088 (N_2088,N_2047,N_2042);
nand U2089 (N_2089,N_2000,N_2007);
nor U2090 (N_2090,N_2014,N_2028);
and U2091 (N_2091,N_2012,N_2048);
and U2092 (N_2092,N_2012,N_2033);
and U2093 (N_2093,N_2010,N_2013);
nand U2094 (N_2094,N_2016,N_2008);
nand U2095 (N_2095,N_2021,N_2007);
xnor U2096 (N_2096,N_2025,N_2026);
nor U2097 (N_2097,N_2013,N_2049);
xor U2098 (N_2098,N_2010,N_2027);
or U2099 (N_2099,N_2006,N_2022);
and U2100 (N_2100,N_2064,N_2051);
nor U2101 (N_2101,N_2054,N_2060);
or U2102 (N_2102,N_2078,N_2062);
or U2103 (N_2103,N_2086,N_2091);
or U2104 (N_2104,N_2081,N_2073);
or U2105 (N_2105,N_2058,N_2092);
nand U2106 (N_2106,N_2050,N_2075);
xnor U2107 (N_2107,N_2067,N_2082);
or U2108 (N_2108,N_2098,N_2057);
nand U2109 (N_2109,N_2059,N_2071);
nor U2110 (N_2110,N_2095,N_2088);
nor U2111 (N_2111,N_2083,N_2063);
nand U2112 (N_2112,N_2085,N_2077);
or U2113 (N_2113,N_2089,N_2087);
nand U2114 (N_2114,N_2056,N_2093);
nand U2115 (N_2115,N_2099,N_2068);
nor U2116 (N_2116,N_2076,N_2079);
nor U2117 (N_2117,N_2061,N_2070);
and U2118 (N_2118,N_2066,N_2065);
or U2119 (N_2119,N_2072,N_2074);
nand U2120 (N_2120,N_2055,N_2052);
xor U2121 (N_2121,N_2094,N_2090);
xnor U2122 (N_2122,N_2080,N_2097);
or U2123 (N_2123,N_2053,N_2096);
nand U2124 (N_2124,N_2069,N_2084);
nor U2125 (N_2125,N_2098,N_2065);
nor U2126 (N_2126,N_2061,N_2068);
or U2127 (N_2127,N_2093,N_2086);
nand U2128 (N_2128,N_2082,N_2053);
or U2129 (N_2129,N_2071,N_2093);
and U2130 (N_2130,N_2086,N_2063);
or U2131 (N_2131,N_2086,N_2059);
and U2132 (N_2132,N_2061,N_2053);
nor U2133 (N_2133,N_2086,N_2075);
or U2134 (N_2134,N_2053,N_2060);
nand U2135 (N_2135,N_2052,N_2085);
nand U2136 (N_2136,N_2085,N_2057);
nor U2137 (N_2137,N_2068,N_2055);
nand U2138 (N_2138,N_2085,N_2068);
nand U2139 (N_2139,N_2064,N_2057);
xnor U2140 (N_2140,N_2077,N_2073);
and U2141 (N_2141,N_2082,N_2058);
nor U2142 (N_2142,N_2064,N_2075);
and U2143 (N_2143,N_2068,N_2095);
nand U2144 (N_2144,N_2053,N_2054);
nand U2145 (N_2145,N_2064,N_2071);
or U2146 (N_2146,N_2093,N_2070);
nand U2147 (N_2147,N_2089,N_2079);
and U2148 (N_2148,N_2072,N_2080);
nor U2149 (N_2149,N_2071,N_2095);
nand U2150 (N_2150,N_2146,N_2109);
nand U2151 (N_2151,N_2107,N_2121);
or U2152 (N_2152,N_2133,N_2112);
or U2153 (N_2153,N_2119,N_2130);
or U2154 (N_2154,N_2145,N_2116);
and U2155 (N_2155,N_2131,N_2101);
nor U2156 (N_2156,N_2128,N_2127);
nand U2157 (N_2157,N_2147,N_2126);
or U2158 (N_2158,N_2115,N_2134);
or U2159 (N_2159,N_2113,N_2102);
nor U2160 (N_2160,N_2143,N_2124);
nand U2161 (N_2161,N_2100,N_2118);
nand U2162 (N_2162,N_2136,N_2141);
and U2163 (N_2163,N_2142,N_2139);
nand U2164 (N_2164,N_2148,N_2123);
and U2165 (N_2165,N_2111,N_2103);
and U2166 (N_2166,N_2149,N_2138);
nor U2167 (N_2167,N_2106,N_2117);
and U2168 (N_2168,N_2135,N_2105);
or U2169 (N_2169,N_2104,N_2137);
xor U2170 (N_2170,N_2132,N_2129);
nand U2171 (N_2171,N_2110,N_2114);
nand U2172 (N_2172,N_2125,N_2140);
nor U2173 (N_2173,N_2144,N_2120);
nand U2174 (N_2174,N_2108,N_2122);
xor U2175 (N_2175,N_2117,N_2148);
and U2176 (N_2176,N_2133,N_2137);
and U2177 (N_2177,N_2148,N_2127);
xnor U2178 (N_2178,N_2117,N_2136);
xor U2179 (N_2179,N_2104,N_2136);
nand U2180 (N_2180,N_2101,N_2116);
or U2181 (N_2181,N_2119,N_2106);
nand U2182 (N_2182,N_2131,N_2129);
or U2183 (N_2183,N_2137,N_2127);
nor U2184 (N_2184,N_2120,N_2102);
and U2185 (N_2185,N_2133,N_2100);
nor U2186 (N_2186,N_2106,N_2142);
nor U2187 (N_2187,N_2142,N_2103);
nor U2188 (N_2188,N_2139,N_2126);
nand U2189 (N_2189,N_2138,N_2119);
nand U2190 (N_2190,N_2126,N_2119);
and U2191 (N_2191,N_2102,N_2139);
and U2192 (N_2192,N_2133,N_2127);
nor U2193 (N_2193,N_2148,N_2115);
nand U2194 (N_2194,N_2145,N_2123);
nand U2195 (N_2195,N_2136,N_2122);
nand U2196 (N_2196,N_2126,N_2145);
xnor U2197 (N_2197,N_2101,N_2144);
nand U2198 (N_2198,N_2144,N_2139);
nor U2199 (N_2199,N_2101,N_2124);
and U2200 (N_2200,N_2186,N_2166);
and U2201 (N_2201,N_2169,N_2163);
or U2202 (N_2202,N_2178,N_2150);
or U2203 (N_2203,N_2187,N_2160);
nor U2204 (N_2204,N_2165,N_2151);
xor U2205 (N_2205,N_2176,N_2198);
and U2206 (N_2206,N_2154,N_2177);
or U2207 (N_2207,N_2181,N_2173);
and U2208 (N_2208,N_2162,N_2194);
nand U2209 (N_2209,N_2184,N_2175);
nor U2210 (N_2210,N_2191,N_2199);
nor U2211 (N_2211,N_2189,N_2172);
and U2212 (N_2212,N_2159,N_2156);
and U2213 (N_2213,N_2168,N_2195);
or U2214 (N_2214,N_2185,N_2171);
or U2215 (N_2215,N_2170,N_2183);
or U2216 (N_2216,N_2196,N_2157);
or U2217 (N_2217,N_2192,N_2152);
nor U2218 (N_2218,N_2179,N_2174);
xnor U2219 (N_2219,N_2190,N_2167);
xnor U2220 (N_2220,N_2182,N_2197);
nand U2221 (N_2221,N_2153,N_2180);
nor U2222 (N_2222,N_2193,N_2155);
or U2223 (N_2223,N_2158,N_2188);
nor U2224 (N_2224,N_2164,N_2161);
or U2225 (N_2225,N_2178,N_2161);
nor U2226 (N_2226,N_2184,N_2150);
and U2227 (N_2227,N_2191,N_2172);
or U2228 (N_2228,N_2195,N_2193);
nand U2229 (N_2229,N_2191,N_2175);
and U2230 (N_2230,N_2196,N_2174);
and U2231 (N_2231,N_2191,N_2155);
and U2232 (N_2232,N_2155,N_2178);
nand U2233 (N_2233,N_2158,N_2174);
or U2234 (N_2234,N_2186,N_2199);
nor U2235 (N_2235,N_2161,N_2152);
or U2236 (N_2236,N_2189,N_2155);
nor U2237 (N_2237,N_2198,N_2170);
nor U2238 (N_2238,N_2170,N_2187);
or U2239 (N_2239,N_2167,N_2153);
nand U2240 (N_2240,N_2179,N_2150);
or U2241 (N_2241,N_2169,N_2179);
xnor U2242 (N_2242,N_2196,N_2193);
and U2243 (N_2243,N_2174,N_2177);
or U2244 (N_2244,N_2185,N_2155);
or U2245 (N_2245,N_2194,N_2180);
or U2246 (N_2246,N_2161,N_2160);
and U2247 (N_2247,N_2192,N_2165);
or U2248 (N_2248,N_2181,N_2160);
nor U2249 (N_2249,N_2176,N_2181);
and U2250 (N_2250,N_2242,N_2221);
and U2251 (N_2251,N_2224,N_2215);
nand U2252 (N_2252,N_2227,N_2213);
or U2253 (N_2253,N_2238,N_2214);
nand U2254 (N_2254,N_2204,N_2222);
nor U2255 (N_2255,N_2202,N_2231);
or U2256 (N_2256,N_2226,N_2237);
nor U2257 (N_2257,N_2235,N_2248);
nor U2258 (N_2258,N_2239,N_2206);
nand U2259 (N_2259,N_2244,N_2247);
or U2260 (N_2260,N_2245,N_2220);
xnor U2261 (N_2261,N_2216,N_2201);
and U2262 (N_2262,N_2208,N_2249);
nand U2263 (N_2263,N_2229,N_2236);
or U2264 (N_2264,N_2200,N_2225);
nor U2265 (N_2265,N_2219,N_2228);
nor U2266 (N_2266,N_2207,N_2218);
or U2267 (N_2267,N_2246,N_2211);
or U2268 (N_2268,N_2210,N_2203);
xnor U2269 (N_2269,N_2241,N_2217);
or U2270 (N_2270,N_2232,N_2240);
nor U2271 (N_2271,N_2209,N_2243);
and U2272 (N_2272,N_2212,N_2233);
nor U2273 (N_2273,N_2223,N_2234);
and U2274 (N_2274,N_2205,N_2230);
nand U2275 (N_2275,N_2220,N_2218);
and U2276 (N_2276,N_2218,N_2248);
and U2277 (N_2277,N_2237,N_2240);
xor U2278 (N_2278,N_2206,N_2217);
nor U2279 (N_2279,N_2227,N_2220);
nor U2280 (N_2280,N_2223,N_2214);
nor U2281 (N_2281,N_2240,N_2224);
or U2282 (N_2282,N_2213,N_2209);
nand U2283 (N_2283,N_2219,N_2203);
nor U2284 (N_2284,N_2206,N_2244);
and U2285 (N_2285,N_2235,N_2229);
nand U2286 (N_2286,N_2232,N_2214);
nand U2287 (N_2287,N_2213,N_2220);
nand U2288 (N_2288,N_2230,N_2228);
or U2289 (N_2289,N_2235,N_2222);
or U2290 (N_2290,N_2204,N_2214);
nor U2291 (N_2291,N_2230,N_2238);
and U2292 (N_2292,N_2206,N_2218);
or U2293 (N_2293,N_2224,N_2235);
xor U2294 (N_2294,N_2201,N_2242);
or U2295 (N_2295,N_2217,N_2233);
or U2296 (N_2296,N_2208,N_2229);
or U2297 (N_2297,N_2217,N_2249);
nor U2298 (N_2298,N_2204,N_2203);
nor U2299 (N_2299,N_2200,N_2208);
or U2300 (N_2300,N_2287,N_2273);
nand U2301 (N_2301,N_2299,N_2293);
or U2302 (N_2302,N_2252,N_2266);
nand U2303 (N_2303,N_2279,N_2278);
and U2304 (N_2304,N_2271,N_2270);
nor U2305 (N_2305,N_2280,N_2265);
or U2306 (N_2306,N_2263,N_2254);
xor U2307 (N_2307,N_2251,N_2275);
or U2308 (N_2308,N_2262,N_2264);
nand U2309 (N_2309,N_2259,N_2291);
nand U2310 (N_2310,N_2256,N_2282);
nand U2311 (N_2311,N_2288,N_2283);
xnor U2312 (N_2312,N_2289,N_2267);
nor U2313 (N_2313,N_2261,N_2295);
and U2314 (N_2314,N_2250,N_2296);
nand U2315 (N_2315,N_2255,N_2260);
nand U2316 (N_2316,N_2272,N_2269);
nor U2317 (N_2317,N_2284,N_2274);
nor U2318 (N_2318,N_2298,N_2281);
or U2319 (N_2319,N_2253,N_2276);
nand U2320 (N_2320,N_2258,N_2290);
and U2321 (N_2321,N_2292,N_2286);
or U2322 (N_2322,N_2297,N_2268);
and U2323 (N_2323,N_2294,N_2257);
nor U2324 (N_2324,N_2277,N_2285);
or U2325 (N_2325,N_2274,N_2283);
nor U2326 (N_2326,N_2266,N_2261);
and U2327 (N_2327,N_2291,N_2298);
nor U2328 (N_2328,N_2256,N_2294);
xor U2329 (N_2329,N_2289,N_2260);
xor U2330 (N_2330,N_2297,N_2286);
nor U2331 (N_2331,N_2278,N_2290);
nand U2332 (N_2332,N_2253,N_2268);
or U2333 (N_2333,N_2251,N_2263);
nand U2334 (N_2334,N_2283,N_2295);
or U2335 (N_2335,N_2286,N_2281);
and U2336 (N_2336,N_2265,N_2259);
and U2337 (N_2337,N_2298,N_2290);
or U2338 (N_2338,N_2263,N_2286);
nor U2339 (N_2339,N_2282,N_2290);
nor U2340 (N_2340,N_2263,N_2273);
and U2341 (N_2341,N_2287,N_2253);
and U2342 (N_2342,N_2288,N_2275);
nand U2343 (N_2343,N_2253,N_2271);
nor U2344 (N_2344,N_2289,N_2254);
nand U2345 (N_2345,N_2279,N_2274);
xnor U2346 (N_2346,N_2272,N_2275);
nand U2347 (N_2347,N_2272,N_2298);
and U2348 (N_2348,N_2285,N_2256);
xnor U2349 (N_2349,N_2268,N_2291);
nor U2350 (N_2350,N_2342,N_2319);
or U2351 (N_2351,N_2309,N_2316);
or U2352 (N_2352,N_2332,N_2328);
and U2353 (N_2353,N_2322,N_2315);
or U2354 (N_2354,N_2312,N_2317);
nor U2355 (N_2355,N_2302,N_2307);
xor U2356 (N_2356,N_2324,N_2327);
or U2357 (N_2357,N_2349,N_2318);
xor U2358 (N_2358,N_2321,N_2336);
nor U2359 (N_2359,N_2311,N_2310);
xor U2360 (N_2360,N_2340,N_2337);
and U2361 (N_2361,N_2335,N_2320);
nand U2362 (N_2362,N_2334,N_2339);
and U2363 (N_2363,N_2347,N_2314);
nor U2364 (N_2364,N_2300,N_2325);
and U2365 (N_2365,N_2338,N_2331);
nand U2366 (N_2366,N_2301,N_2305);
nor U2367 (N_2367,N_2348,N_2308);
and U2368 (N_2368,N_2313,N_2344);
nor U2369 (N_2369,N_2323,N_2306);
nor U2370 (N_2370,N_2341,N_2329);
nor U2371 (N_2371,N_2333,N_2303);
or U2372 (N_2372,N_2346,N_2326);
nor U2373 (N_2373,N_2304,N_2345);
and U2374 (N_2374,N_2343,N_2330);
nor U2375 (N_2375,N_2307,N_2309);
nand U2376 (N_2376,N_2321,N_2301);
nor U2377 (N_2377,N_2331,N_2307);
and U2378 (N_2378,N_2321,N_2345);
nor U2379 (N_2379,N_2323,N_2330);
nand U2380 (N_2380,N_2338,N_2323);
or U2381 (N_2381,N_2327,N_2319);
xor U2382 (N_2382,N_2344,N_2309);
nand U2383 (N_2383,N_2310,N_2349);
or U2384 (N_2384,N_2338,N_2310);
or U2385 (N_2385,N_2304,N_2305);
xnor U2386 (N_2386,N_2320,N_2332);
or U2387 (N_2387,N_2340,N_2318);
nor U2388 (N_2388,N_2317,N_2307);
or U2389 (N_2389,N_2339,N_2303);
nor U2390 (N_2390,N_2315,N_2328);
and U2391 (N_2391,N_2301,N_2315);
and U2392 (N_2392,N_2342,N_2331);
and U2393 (N_2393,N_2349,N_2331);
nor U2394 (N_2394,N_2336,N_2331);
nand U2395 (N_2395,N_2330,N_2303);
or U2396 (N_2396,N_2317,N_2316);
nor U2397 (N_2397,N_2314,N_2337);
xor U2398 (N_2398,N_2346,N_2340);
and U2399 (N_2399,N_2309,N_2308);
nand U2400 (N_2400,N_2391,N_2380);
and U2401 (N_2401,N_2394,N_2368);
nor U2402 (N_2402,N_2390,N_2386);
and U2403 (N_2403,N_2378,N_2372);
or U2404 (N_2404,N_2375,N_2392);
nand U2405 (N_2405,N_2358,N_2365);
or U2406 (N_2406,N_2393,N_2357);
nor U2407 (N_2407,N_2369,N_2356);
nand U2408 (N_2408,N_2355,N_2370);
and U2409 (N_2409,N_2371,N_2398);
or U2410 (N_2410,N_2383,N_2389);
and U2411 (N_2411,N_2387,N_2395);
nand U2412 (N_2412,N_2382,N_2363);
nor U2413 (N_2413,N_2350,N_2385);
nor U2414 (N_2414,N_2374,N_2352);
nand U2415 (N_2415,N_2366,N_2361);
nor U2416 (N_2416,N_2354,N_2396);
and U2417 (N_2417,N_2399,N_2379);
nand U2418 (N_2418,N_2367,N_2376);
nand U2419 (N_2419,N_2353,N_2377);
nor U2420 (N_2420,N_2364,N_2388);
and U2421 (N_2421,N_2397,N_2360);
and U2422 (N_2422,N_2351,N_2384);
nand U2423 (N_2423,N_2362,N_2359);
nand U2424 (N_2424,N_2381,N_2373);
nand U2425 (N_2425,N_2356,N_2378);
nand U2426 (N_2426,N_2380,N_2350);
xnor U2427 (N_2427,N_2353,N_2362);
xnor U2428 (N_2428,N_2350,N_2356);
or U2429 (N_2429,N_2389,N_2365);
nor U2430 (N_2430,N_2370,N_2350);
nor U2431 (N_2431,N_2395,N_2376);
nor U2432 (N_2432,N_2371,N_2394);
nand U2433 (N_2433,N_2356,N_2370);
nand U2434 (N_2434,N_2399,N_2352);
nand U2435 (N_2435,N_2370,N_2394);
and U2436 (N_2436,N_2353,N_2382);
or U2437 (N_2437,N_2386,N_2387);
nand U2438 (N_2438,N_2363,N_2365);
nor U2439 (N_2439,N_2354,N_2384);
nand U2440 (N_2440,N_2399,N_2383);
xnor U2441 (N_2441,N_2370,N_2357);
nor U2442 (N_2442,N_2358,N_2356);
nand U2443 (N_2443,N_2362,N_2373);
or U2444 (N_2444,N_2388,N_2383);
nor U2445 (N_2445,N_2378,N_2381);
and U2446 (N_2446,N_2367,N_2397);
nand U2447 (N_2447,N_2358,N_2357);
nand U2448 (N_2448,N_2367,N_2395);
xnor U2449 (N_2449,N_2380,N_2363);
or U2450 (N_2450,N_2412,N_2444);
nor U2451 (N_2451,N_2431,N_2421);
nand U2452 (N_2452,N_2428,N_2447);
or U2453 (N_2453,N_2402,N_2404);
nand U2454 (N_2454,N_2426,N_2449);
or U2455 (N_2455,N_2441,N_2434);
and U2456 (N_2456,N_2435,N_2429);
and U2457 (N_2457,N_2405,N_2445);
nand U2458 (N_2458,N_2420,N_2414);
xor U2459 (N_2459,N_2401,N_2439);
nor U2460 (N_2460,N_2427,N_2430);
nand U2461 (N_2461,N_2406,N_2413);
or U2462 (N_2462,N_2418,N_2443);
nand U2463 (N_2463,N_2411,N_2415);
nor U2464 (N_2464,N_2438,N_2417);
and U2465 (N_2465,N_2442,N_2433);
nand U2466 (N_2466,N_2448,N_2407);
nor U2467 (N_2467,N_2423,N_2409);
nor U2468 (N_2468,N_2410,N_2446);
and U2469 (N_2469,N_2408,N_2400);
or U2470 (N_2470,N_2422,N_2432);
or U2471 (N_2471,N_2436,N_2419);
or U2472 (N_2472,N_2424,N_2437);
nor U2473 (N_2473,N_2440,N_2425);
nand U2474 (N_2474,N_2416,N_2403);
xor U2475 (N_2475,N_2414,N_2416);
nand U2476 (N_2476,N_2424,N_2436);
or U2477 (N_2477,N_2442,N_2400);
nor U2478 (N_2478,N_2425,N_2419);
nor U2479 (N_2479,N_2432,N_2412);
nor U2480 (N_2480,N_2404,N_2400);
and U2481 (N_2481,N_2430,N_2419);
xnor U2482 (N_2482,N_2414,N_2430);
nand U2483 (N_2483,N_2441,N_2439);
and U2484 (N_2484,N_2438,N_2440);
nor U2485 (N_2485,N_2431,N_2445);
and U2486 (N_2486,N_2408,N_2426);
or U2487 (N_2487,N_2412,N_2422);
nor U2488 (N_2488,N_2410,N_2437);
and U2489 (N_2489,N_2447,N_2416);
or U2490 (N_2490,N_2404,N_2444);
and U2491 (N_2491,N_2404,N_2434);
nor U2492 (N_2492,N_2445,N_2408);
or U2493 (N_2493,N_2419,N_2443);
nor U2494 (N_2494,N_2414,N_2446);
nor U2495 (N_2495,N_2411,N_2402);
and U2496 (N_2496,N_2423,N_2427);
and U2497 (N_2497,N_2444,N_2426);
nor U2498 (N_2498,N_2445,N_2440);
or U2499 (N_2499,N_2446,N_2430);
and U2500 (N_2500,N_2496,N_2461);
or U2501 (N_2501,N_2464,N_2463);
or U2502 (N_2502,N_2488,N_2478);
nand U2503 (N_2503,N_2457,N_2460);
nor U2504 (N_2504,N_2471,N_2459);
or U2505 (N_2505,N_2450,N_2479);
and U2506 (N_2506,N_2476,N_2497);
and U2507 (N_2507,N_2495,N_2487);
nand U2508 (N_2508,N_2455,N_2482);
nor U2509 (N_2509,N_2489,N_2472);
nor U2510 (N_2510,N_2475,N_2486);
nor U2511 (N_2511,N_2481,N_2492);
or U2512 (N_2512,N_2473,N_2477);
or U2513 (N_2513,N_2494,N_2490);
or U2514 (N_2514,N_2468,N_2466);
nand U2515 (N_2515,N_2458,N_2453);
nand U2516 (N_2516,N_2470,N_2480);
and U2517 (N_2517,N_2469,N_2474);
or U2518 (N_2518,N_2452,N_2493);
nor U2519 (N_2519,N_2483,N_2454);
nand U2520 (N_2520,N_2462,N_2467);
nand U2521 (N_2521,N_2456,N_2451);
nor U2522 (N_2522,N_2491,N_2498);
or U2523 (N_2523,N_2484,N_2485);
or U2524 (N_2524,N_2465,N_2499);
nor U2525 (N_2525,N_2453,N_2476);
and U2526 (N_2526,N_2491,N_2475);
nand U2527 (N_2527,N_2462,N_2474);
or U2528 (N_2528,N_2471,N_2470);
xor U2529 (N_2529,N_2476,N_2487);
and U2530 (N_2530,N_2474,N_2484);
nor U2531 (N_2531,N_2491,N_2477);
or U2532 (N_2532,N_2495,N_2485);
nor U2533 (N_2533,N_2456,N_2482);
and U2534 (N_2534,N_2475,N_2476);
xor U2535 (N_2535,N_2460,N_2458);
or U2536 (N_2536,N_2484,N_2476);
and U2537 (N_2537,N_2490,N_2492);
xor U2538 (N_2538,N_2459,N_2491);
xnor U2539 (N_2539,N_2498,N_2454);
nor U2540 (N_2540,N_2480,N_2450);
and U2541 (N_2541,N_2461,N_2450);
or U2542 (N_2542,N_2494,N_2497);
nor U2543 (N_2543,N_2451,N_2480);
or U2544 (N_2544,N_2494,N_2477);
and U2545 (N_2545,N_2474,N_2468);
and U2546 (N_2546,N_2478,N_2498);
nand U2547 (N_2547,N_2485,N_2477);
nor U2548 (N_2548,N_2481,N_2452);
and U2549 (N_2549,N_2460,N_2450);
and U2550 (N_2550,N_2521,N_2540);
or U2551 (N_2551,N_2533,N_2505);
and U2552 (N_2552,N_2527,N_2542);
or U2553 (N_2553,N_2502,N_2548);
and U2554 (N_2554,N_2545,N_2526);
nand U2555 (N_2555,N_2538,N_2510);
nand U2556 (N_2556,N_2513,N_2537);
xnor U2557 (N_2557,N_2504,N_2508);
and U2558 (N_2558,N_2529,N_2523);
and U2559 (N_2559,N_2522,N_2547);
or U2560 (N_2560,N_2541,N_2532);
or U2561 (N_2561,N_2520,N_2539);
or U2562 (N_2562,N_2503,N_2519);
and U2563 (N_2563,N_2535,N_2530);
nor U2564 (N_2564,N_2525,N_2518);
nand U2565 (N_2565,N_2517,N_2534);
nor U2566 (N_2566,N_2528,N_2531);
nor U2567 (N_2567,N_2515,N_2536);
and U2568 (N_2568,N_2544,N_2516);
nor U2569 (N_2569,N_2507,N_2501);
or U2570 (N_2570,N_2543,N_2509);
or U2571 (N_2571,N_2512,N_2514);
nor U2572 (N_2572,N_2511,N_2549);
nor U2573 (N_2573,N_2546,N_2524);
nor U2574 (N_2574,N_2506,N_2500);
nand U2575 (N_2575,N_2531,N_2540);
xor U2576 (N_2576,N_2505,N_2545);
or U2577 (N_2577,N_2521,N_2509);
and U2578 (N_2578,N_2517,N_2548);
nand U2579 (N_2579,N_2526,N_2513);
nor U2580 (N_2580,N_2539,N_2529);
xnor U2581 (N_2581,N_2503,N_2547);
and U2582 (N_2582,N_2526,N_2501);
or U2583 (N_2583,N_2505,N_2531);
or U2584 (N_2584,N_2521,N_2507);
or U2585 (N_2585,N_2517,N_2540);
and U2586 (N_2586,N_2541,N_2539);
nand U2587 (N_2587,N_2504,N_2527);
or U2588 (N_2588,N_2507,N_2540);
xor U2589 (N_2589,N_2517,N_2539);
or U2590 (N_2590,N_2511,N_2533);
or U2591 (N_2591,N_2539,N_2514);
nand U2592 (N_2592,N_2517,N_2512);
nand U2593 (N_2593,N_2526,N_2522);
nand U2594 (N_2594,N_2517,N_2526);
nor U2595 (N_2595,N_2534,N_2532);
and U2596 (N_2596,N_2516,N_2545);
or U2597 (N_2597,N_2538,N_2504);
xnor U2598 (N_2598,N_2533,N_2507);
and U2599 (N_2599,N_2509,N_2516);
xor U2600 (N_2600,N_2564,N_2561);
nor U2601 (N_2601,N_2584,N_2594);
nor U2602 (N_2602,N_2558,N_2580);
nand U2603 (N_2603,N_2596,N_2572);
or U2604 (N_2604,N_2568,N_2595);
xor U2605 (N_2605,N_2554,N_2550);
nor U2606 (N_2606,N_2577,N_2555);
or U2607 (N_2607,N_2591,N_2581);
nand U2608 (N_2608,N_2579,N_2562);
nand U2609 (N_2609,N_2560,N_2556);
or U2610 (N_2610,N_2552,N_2557);
or U2611 (N_2611,N_2573,N_2588);
nand U2612 (N_2612,N_2574,N_2576);
or U2613 (N_2613,N_2583,N_2590);
and U2614 (N_2614,N_2593,N_2589);
and U2615 (N_2615,N_2565,N_2575);
nand U2616 (N_2616,N_2585,N_2570);
or U2617 (N_2617,N_2599,N_2559);
and U2618 (N_2618,N_2563,N_2578);
xnor U2619 (N_2619,N_2571,N_2592);
nor U2620 (N_2620,N_2586,N_2551);
or U2621 (N_2621,N_2582,N_2598);
nand U2622 (N_2622,N_2587,N_2567);
and U2623 (N_2623,N_2566,N_2569);
xor U2624 (N_2624,N_2597,N_2553);
nand U2625 (N_2625,N_2555,N_2568);
nor U2626 (N_2626,N_2565,N_2584);
or U2627 (N_2627,N_2594,N_2579);
nand U2628 (N_2628,N_2587,N_2576);
nand U2629 (N_2629,N_2597,N_2569);
nand U2630 (N_2630,N_2564,N_2550);
xnor U2631 (N_2631,N_2574,N_2596);
or U2632 (N_2632,N_2596,N_2552);
nor U2633 (N_2633,N_2565,N_2553);
nor U2634 (N_2634,N_2586,N_2570);
nor U2635 (N_2635,N_2594,N_2572);
or U2636 (N_2636,N_2557,N_2577);
xnor U2637 (N_2637,N_2566,N_2556);
nand U2638 (N_2638,N_2582,N_2556);
nor U2639 (N_2639,N_2561,N_2554);
nor U2640 (N_2640,N_2559,N_2554);
nor U2641 (N_2641,N_2591,N_2556);
and U2642 (N_2642,N_2557,N_2569);
xnor U2643 (N_2643,N_2574,N_2586);
and U2644 (N_2644,N_2571,N_2565);
nor U2645 (N_2645,N_2595,N_2596);
nor U2646 (N_2646,N_2566,N_2562);
nand U2647 (N_2647,N_2557,N_2586);
or U2648 (N_2648,N_2593,N_2558);
nand U2649 (N_2649,N_2577,N_2584);
nor U2650 (N_2650,N_2648,N_2642);
nor U2651 (N_2651,N_2604,N_2602);
nand U2652 (N_2652,N_2610,N_2632);
nand U2653 (N_2653,N_2607,N_2612);
and U2654 (N_2654,N_2621,N_2628);
or U2655 (N_2655,N_2609,N_2643);
nor U2656 (N_2656,N_2601,N_2629);
or U2657 (N_2657,N_2620,N_2647);
and U2658 (N_2658,N_2634,N_2616);
and U2659 (N_2659,N_2608,N_2613);
nor U2660 (N_2660,N_2624,N_2639);
and U2661 (N_2661,N_2619,N_2603);
or U2662 (N_2662,N_2649,N_2626);
nor U2663 (N_2663,N_2644,N_2611);
nand U2664 (N_2664,N_2618,N_2627);
nor U2665 (N_2665,N_2631,N_2623);
nand U2666 (N_2666,N_2638,N_2633);
or U2667 (N_2667,N_2600,N_2641);
nor U2668 (N_2668,N_2625,N_2640);
or U2669 (N_2669,N_2615,N_2646);
nand U2670 (N_2670,N_2614,N_2622);
and U2671 (N_2671,N_2617,N_2605);
nand U2672 (N_2672,N_2645,N_2606);
nor U2673 (N_2673,N_2630,N_2635);
or U2674 (N_2674,N_2637,N_2636);
nor U2675 (N_2675,N_2617,N_2625);
nor U2676 (N_2676,N_2628,N_2630);
nor U2677 (N_2677,N_2604,N_2639);
nand U2678 (N_2678,N_2648,N_2623);
or U2679 (N_2679,N_2644,N_2619);
and U2680 (N_2680,N_2624,N_2641);
nor U2681 (N_2681,N_2621,N_2616);
or U2682 (N_2682,N_2613,N_2617);
and U2683 (N_2683,N_2631,N_2649);
and U2684 (N_2684,N_2607,N_2634);
or U2685 (N_2685,N_2634,N_2638);
xor U2686 (N_2686,N_2621,N_2620);
nand U2687 (N_2687,N_2611,N_2632);
nor U2688 (N_2688,N_2629,N_2620);
nand U2689 (N_2689,N_2622,N_2625);
nand U2690 (N_2690,N_2624,N_2602);
or U2691 (N_2691,N_2621,N_2646);
or U2692 (N_2692,N_2618,N_2628);
nor U2693 (N_2693,N_2644,N_2618);
nor U2694 (N_2694,N_2620,N_2631);
and U2695 (N_2695,N_2639,N_2644);
or U2696 (N_2696,N_2619,N_2641);
or U2697 (N_2697,N_2600,N_2620);
nor U2698 (N_2698,N_2607,N_2635);
nor U2699 (N_2699,N_2616,N_2645);
nor U2700 (N_2700,N_2685,N_2667);
nand U2701 (N_2701,N_2675,N_2693);
or U2702 (N_2702,N_2686,N_2681);
xor U2703 (N_2703,N_2676,N_2687);
and U2704 (N_2704,N_2666,N_2697);
or U2705 (N_2705,N_2673,N_2694);
and U2706 (N_2706,N_2674,N_2658);
nand U2707 (N_2707,N_2662,N_2650);
and U2708 (N_2708,N_2664,N_2678);
nand U2709 (N_2709,N_2690,N_2689);
nor U2710 (N_2710,N_2669,N_2671);
nor U2711 (N_2711,N_2657,N_2659);
nand U2712 (N_2712,N_2699,N_2653);
nand U2713 (N_2713,N_2692,N_2696);
xor U2714 (N_2714,N_2698,N_2665);
and U2715 (N_2715,N_2651,N_2656);
and U2716 (N_2716,N_2677,N_2695);
or U2717 (N_2717,N_2680,N_2672);
or U2718 (N_2718,N_2663,N_2668);
nor U2719 (N_2719,N_2661,N_2679);
nor U2720 (N_2720,N_2684,N_2683);
nor U2721 (N_2721,N_2670,N_2691);
and U2722 (N_2722,N_2654,N_2652);
nand U2723 (N_2723,N_2682,N_2688);
nand U2724 (N_2724,N_2660,N_2655);
nand U2725 (N_2725,N_2694,N_2680);
nand U2726 (N_2726,N_2668,N_2677);
nor U2727 (N_2727,N_2659,N_2689);
and U2728 (N_2728,N_2665,N_2694);
xor U2729 (N_2729,N_2676,N_2657);
or U2730 (N_2730,N_2696,N_2687);
and U2731 (N_2731,N_2671,N_2664);
and U2732 (N_2732,N_2671,N_2655);
nand U2733 (N_2733,N_2659,N_2667);
xor U2734 (N_2734,N_2679,N_2669);
nand U2735 (N_2735,N_2669,N_2692);
or U2736 (N_2736,N_2650,N_2685);
nand U2737 (N_2737,N_2664,N_2691);
xnor U2738 (N_2738,N_2669,N_2688);
nor U2739 (N_2739,N_2683,N_2667);
nor U2740 (N_2740,N_2696,N_2680);
and U2741 (N_2741,N_2685,N_2655);
and U2742 (N_2742,N_2667,N_2675);
nand U2743 (N_2743,N_2698,N_2671);
and U2744 (N_2744,N_2679,N_2693);
nand U2745 (N_2745,N_2694,N_2668);
nor U2746 (N_2746,N_2685,N_2670);
or U2747 (N_2747,N_2677,N_2667);
nand U2748 (N_2748,N_2677,N_2683);
and U2749 (N_2749,N_2664,N_2657);
nand U2750 (N_2750,N_2734,N_2700);
and U2751 (N_2751,N_2709,N_2738);
or U2752 (N_2752,N_2741,N_2717);
nor U2753 (N_2753,N_2707,N_2711);
nand U2754 (N_2754,N_2739,N_2714);
or U2755 (N_2755,N_2731,N_2725);
or U2756 (N_2756,N_2730,N_2746);
or U2757 (N_2757,N_2735,N_2716);
nand U2758 (N_2758,N_2744,N_2710);
and U2759 (N_2759,N_2705,N_2732);
nand U2760 (N_2760,N_2726,N_2737);
nand U2761 (N_2761,N_2743,N_2701);
xor U2762 (N_2762,N_2702,N_2704);
nand U2763 (N_2763,N_2713,N_2736);
nor U2764 (N_2764,N_2749,N_2727);
nor U2765 (N_2765,N_2722,N_2728);
and U2766 (N_2766,N_2708,N_2729);
and U2767 (N_2767,N_2748,N_2723);
and U2768 (N_2768,N_2733,N_2719);
nand U2769 (N_2769,N_2720,N_2706);
xor U2770 (N_2770,N_2745,N_2724);
xor U2771 (N_2771,N_2715,N_2718);
and U2772 (N_2772,N_2712,N_2747);
or U2773 (N_2773,N_2703,N_2740);
nand U2774 (N_2774,N_2742,N_2721);
nand U2775 (N_2775,N_2717,N_2714);
or U2776 (N_2776,N_2725,N_2717);
nor U2777 (N_2777,N_2737,N_2728);
and U2778 (N_2778,N_2749,N_2744);
and U2779 (N_2779,N_2703,N_2739);
nor U2780 (N_2780,N_2744,N_2711);
xnor U2781 (N_2781,N_2747,N_2732);
or U2782 (N_2782,N_2734,N_2704);
nor U2783 (N_2783,N_2726,N_2708);
nor U2784 (N_2784,N_2734,N_2710);
or U2785 (N_2785,N_2729,N_2704);
nor U2786 (N_2786,N_2723,N_2731);
nand U2787 (N_2787,N_2723,N_2700);
nand U2788 (N_2788,N_2747,N_2703);
or U2789 (N_2789,N_2733,N_2707);
or U2790 (N_2790,N_2715,N_2714);
nor U2791 (N_2791,N_2716,N_2739);
nor U2792 (N_2792,N_2739,N_2735);
and U2793 (N_2793,N_2719,N_2722);
and U2794 (N_2794,N_2747,N_2735);
and U2795 (N_2795,N_2710,N_2735);
nand U2796 (N_2796,N_2714,N_2744);
and U2797 (N_2797,N_2727,N_2722);
nor U2798 (N_2798,N_2707,N_2732);
and U2799 (N_2799,N_2715,N_2729);
xnor U2800 (N_2800,N_2799,N_2755);
and U2801 (N_2801,N_2780,N_2775);
or U2802 (N_2802,N_2764,N_2784);
or U2803 (N_2803,N_2773,N_2751);
nand U2804 (N_2804,N_2792,N_2790);
nand U2805 (N_2805,N_2795,N_2797);
or U2806 (N_2806,N_2762,N_2789);
or U2807 (N_2807,N_2761,N_2791);
and U2808 (N_2808,N_2793,N_2788);
and U2809 (N_2809,N_2757,N_2772);
nor U2810 (N_2810,N_2754,N_2767);
or U2811 (N_2811,N_2796,N_2798);
xor U2812 (N_2812,N_2753,N_2760);
and U2813 (N_2813,N_2778,N_2768);
nand U2814 (N_2814,N_2781,N_2763);
or U2815 (N_2815,N_2765,N_2776);
nor U2816 (N_2816,N_2786,N_2787);
or U2817 (N_2817,N_2750,N_2794);
nor U2818 (N_2818,N_2777,N_2758);
nand U2819 (N_2819,N_2774,N_2785);
nor U2820 (N_2820,N_2770,N_2756);
and U2821 (N_2821,N_2782,N_2752);
nand U2822 (N_2822,N_2779,N_2766);
nand U2823 (N_2823,N_2769,N_2783);
xor U2824 (N_2824,N_2771,N_2759);
nor U2825 (N_2825,N_2772,N_2775);
nand U2826 (N_2826,N_2765,N_2760);
or U2827 (N_2827,N_2790,N_2795);
and U2828 (N_2828,N_2791,N_2778);
nor U2829 (N_2829,N_2793,N_2762);
nor U2830 (N_2830,N_2782,N_2770);
and U2831 (N_2831,N_2764,N_2757);
or U2832 (N_2832,N_2782,N_2789);
and U2833 (N_2833,N_2796,N_2772);
xor U2834 (N_2834,N_2758,N_2764);
nand U2835 (N_2835,N_2786,N_2770);
nor U2836 (N_2836,N_2757,N_2779);
and U2837 (N_2837,N_2799,N_2775);
or U2838 (N_2838,N_2797,N_2787);
nand U2839 (N_2839,N_2784,N_2778);
and U2840 (N_2840,N_2786,N_2751);
nor U2841 (N_2841,N_2791,N_2768);
nor U2842 (N_2842,N_2750,N_2788);
or U2843 (N_2843,N_2758,N_2780);
nand U2844 (N_2844,N_2796,N_2799);
and U2845 (N_2845,N_2753,N_2771);
nand U2846 (N_2846,N_2758,N_2789);
and U2847 (N_2847,N_2751,N_2775);
xor U2848 (N_2848,N_2765,N_2772);
nor U2849 (N_2849,N_2787,N_2792);
and U2850 (N_2850,N_2804,N_2823);
or U2851 (N_2851,N_2832,N_2835);
or U2852 (N_2852,N_2845,N_2830);
and U2853 (N_2853,N_2840,N_2822);
nor U2854 (N_2854,N_2816,N_2806);
nor U2855 (N_2855,N_2826,N_2838);
nand U2856 (N_2856,N_2817,N_2807);
nor U2857 (N_2857,N_2848,N_2836);
nand U2858 (N_2858,N_2801,N_2825);
and U2859 (N_2859,N_2833,N_2824);
and U2860 (N_2860,N_2828,N_2839);
and U2861 (N_2861,N_2829,N_2841);
nand U2862 (N_2862,N_2809,N_2831);
or U2863 (N_2863,N_2805,N_2849);
and U2864 (N_2864,N_2820,N_2837);
or U2865 (N_2865,N_2802,N_2847);
nor U2866 (N_2866,N_2810,N_2844);
xnor U2867 (N_2867,N_2818,N_2814);
nor U2868 (N_2868,N_2813,N_2843);
xnor U2869 (N_2869,N_2815,N_2834);
nor U2870 (N_2870,N_2811,N_2827);
xor U2871 (N_2871,N_2803,N_2819);
and U2872 (N_2872,N_2842,N_2846);
xor U2873 (N_2873,N_2800,N_2821);
nor U2874 (N_2874,N_2812,N_2808);
nand U2875 (N_2875,N_2837,N_2832);
xnor U2876 (N_2876,N_2817,N_2820);
or U2877 (N_2877,N_2847,N_2821);
nor U2878 (N_2878,N_2833,N_2840);
xor U2879 (N_2879,N_2840,N_2804);
nor U2880 (N_2880,N_2849,N_2801);
or U2881 (N_2881,N_2820,N_2809);
nor U2882 (N_2882,N_2823,N_2806);
nor U2883 (N_2883,N_2802,N_2817);
nand U2884 (N_2884,N_2808,N_2841);
nand U2885 (N_2885,N_2837,N_2836);
nor U2886 (N_2886,N_2844,N_2847);
and U2887 (N_2887,N_2834,N_2846);
or U2888 (N_2888,N_2823,N_2842);
nand U2889 (N_2889,N_2841,N_2844);
and U2890 (N_2890,N_2848,N_2820);
and U2891 (N_2891,N_2843,N_2811);
and U2892 (N_2892,N_2846,N_2800);
or U2893 (N_2893,N_2838,N_2821);
xor U2894 (N_2894,N_2840,N_2827);
nor U2895 (N_2895,N_2833,N_2848);
or U2896 (N_2896,N_2849,N_2812);
xor U2897 (N_2897,N_2832,N_2820);
nor U2898 (N_2898,N_2820,N_2807);
or U2899 (N_2899,N_2801,N_2808);
or U2900 (N_2900,N_2875,N_2898);
nand U2901 (N_2901,N_2881,N_2850);
nand U2902 (N_2902,N_2893,N_2890);
and U2903 (N_2903,N_2862,N_2892);
nor U2904 (N_2904,N_2894,N_2869);
nand U2905 (N_2905,N_2856,N_2899);
and U2906 (N_2906,N_2868,N_2879);
nand U2907 (N_2907,N_2863,N_2852);
or U2908 (N_2908,N_2865,N_2860);
nand U2909 (N_2909,N_2861,N_2870);
nand U2910 (N_2910,N_2853,N_2880);
and U2911 (N_2911,N_2872,N_2855);
nor U2912 (N_2912,N_2891,N_2882);
and U2913 (N_2913,N_2873,N_2897);
or U2914 (N_2914,N_2885,N_2888);
and U2915 (N_2915,N_2887,N_2877);
nor U2916 (N_2916,N_2866,N_2876);
xnor U2917 (N_2917,N_2886,N_2878);
nor U2918 (N_2918,N_2859,N_2884);
and U2919 (N_2919,N_2889,N_2864);
nor U2920 (N_2920,N_2874,N_2854);
nor U2921 (N_2921,N_2896,N_2858);
nor U2922 (N_2922,N_2895,N_2871);
and U2923 (N_2923,N_2857,N_2867);
and U2924 (N_2924,N_2883,N_2851);
and U2925 (N_2925,N_2860,N_2882);
nor U2926 (N_2926,N_2891,N_2853);
or U2927 (N_2927,N_2884,N_2892);
nor U2928 (N_2928,N_2864,N_2877);
xor U2929 (N_2929,N_2854,N_2886);
nor U2930 (N_2930,N_2877,N_2859);
and U2931 (N_2931,N_2856,N_2854);
nor U2932 (N_2932,N_2873,N_2890);
nand U2933 (N_2933,N_2865,N_2889);
nor U2934 (N_2934,N_2891,N_2856);
and U2935 (N_2935,N_2881,N_2890);
and U2936 (N_2936,N_2871,N_2857);
nand U2937 (N_2937,N_2881,N_2866);
xnor U2938 (N_2938,N_2871,N_2882);
and U2939 (N_2939,N_2861,N_2866);
nor U2940 (N_2940,N_2898,N_2855);
or U2941 (N_2941,N_2884,N_2878);
nand U2942 (N_2942,N_2859,N_2874);
and U2943 (N_2943,N_2891,N_2887);
nand U2944 (N_2944,N_2871,N_2875);
or U2945 (N_2945,N_2861,N_2853);
or U2946 (N_2946,N_2850,N_2875);
or U2947 (N_2947,N_2899,N_2898);
xnor U2948 (N_2948,N_2886,N_2865);
nor U2949 (N_2949,N_2893,N_2860);
or U2950 (N_2950,N_2946,N_2915);
nand U2951 (N_2951,N_2905,N_2908);
nand U2952 (N_2952,N_2940,N_2947);
nor U2953 (N_2953,N_2931,N_2937);
and U2954 (N_2954,N_2945,N_2930);
or U2955 (N_2955,N_2913,N_2929);
and U2956 (N_2956,N_2919,N_2906);
nor U2957 (N_2957,N_2901,N_2942);
xor U2958 (N_2958,N_2944,N_2927);
and U2959 (N_2959,N_2948,N_2911);
and U2960 (N_2960,N_2916,N_2939);
nand U2961 (N_2961,N_2918,N_2924);
and U2962 (N_2962,N_2907,N_2949);
nand U2963 (N_2963,N_2925,N_2936);
nand U2964 (N_2964,N_2933,N_2914);
and U2965 (N_2965,N_2935,N_2912);
nor U2966 (N_2966,N_2904,N_2910);
or U2967 (N_2967,N_2900,N_2902);
and U2968 (N_2968,N_2943,N_2928);
nor U2969 (N_2969,N_2903,N_2926);
or U2970 (N_2970,N_2934,N_2917);
nor U2971 (N_2971,N_2932,N_2922);
or U2972 (N_2972,N_2941,N_2938);
or U2973 (N_2973,N_2920,N_2921);
and U2974 (N_2974,N_2923,N_2909);
nand U2975 (N_2975,N_2949,N_2948);
and U2976 (N_2976,N_2932,N_2944);
nor U2977 (N_2977,N_2912,N_2904);
nand U2978 (N_2978,N_2924,N_2907);
or U2979 (N_2979,N_2906,N_2905);
and U2980 (N_2980,N_2925,N_2939);
nand U2981 (N_2981,N_2949,N_2928);
xor U2982 (N_2982,N_2909,N_2941);
and U2983 (N_2983,N_2929,N_2941);
or U2984 (N_2984,N_2901,N_2929);
or U2985 (N_2985,N_2935,N_2944);
nand U2986 (N_2986,N_2914,N_2917);
or U2987 (N_2987,N_2917,N_2918);
nand U2988 (N_2988,N_2924,N_2944);
or U2989 (N_2989,N_2949,N_2942);
or U2990 (N_2990,N_2947,N_2907);
xnor U2991 (N_2991,N_2907,N_2901);
nor U2992 (N_2992,N_2941,N_2926);
nand U2993 (N_2993,N_2931,N_2948);
nor U2994 (N_2994,N_2920,N_2931);
and U2995 (N_2995,N_2909,N_2907);
nand U2996 (N_2996,N_2939,N_2902);
and U2997 (N_2997,N_2901,N_2949);
and U2998 (N_2998,N_2913,N_2940);
or U2999 (N_2999,N_2929,N_2924);
or UO_0 (O_0,N_2992,N_2996);
nor UO_1 (O_1,N_2989,N_2963);
nor UO_2 (O_2,N_2973,N_2975);
or UO_3 (O_3,N_2953,N_2971);
or UO_4 (O_4,N_2954,N_2967);
and UO_5 (O_5,N_2986,N_2951);
or UO_6 (O_6,N_2974,N_2978);
nand UO_7 (O_7,N_2959,N_2970);
and UO_8 (O_8,N_2982,N_2950);
nand UO_9 (O_9,N_2956,N_2997);
nor UO_10 (O_10,N_2965,N_2972);
xnor UO_11 (O_11,N_2993,N_2961);
xnor UO_12 (O_12,N_2991,N_2969);
and UO_13 (O_13,N_2952,N_2955);
xnor UO_14 (O_14,N_2976,N_2962);
nor UO_15 (O_15,N_2968,N_2957);
and UO_16 (O_16,N_2990,N_2977);
nand UO_17 (O_17,N_2998,N_2985);
or UO_18 (O_18,N_2995,N_2979);
xnor UO_19 (O_19,N_2984,N_2980);
and UO_20 (O_20,N_2994,N_2988);
nand UO_21 (O_21,N_2983,N_2960);
or UO_22 (O_22,N_2958,N_2981);
nand UO_23 (O_23,N_2999,N_2966);
or UO_24 (O_24,N_2987,N_2964);
and UO_25 (O_25,N_2995,N_2967);
and UO_26 (O_26,N_2953,N_2964);
xor UO_27 (O_27,N_2983,N_2993);
xnor UO_28 (O_28,N_2989,N_2973);
xnor UO_29 (O_29,N_2954,N_2989);
xor UO_30 (O_30,N_2955,N_2954);
and UO_31 (O_31,N_2978,N_2972);
or UO_32 (O_32,N_2967,N_2976);
and UO_33 (O_33,N_2994,N_2958);
and UO_34 (O_34,N_2958,N_2950);
or UO_35 (O_35,N_2972,N_2988);
nor UO_36 (O_36,N_2980,N_2987);
nand UO_37 (O_37,N_2955,N_2994);
nor UO_38 (O_38,N_2958,N_2980);
and UO_39 (O_39,N_2973,N_2963);
or UO_40 (O_40,N_2951,N_2992);
nor UO_41 (O_41,N_2975,N_2987);
nand UO_42 (O_42,N_2997,N_2960);
nor UO_43 (O_43,N_2991,N_2982);
nand UO_44 (O_44,N_2958,N_2972);
and UO_45 (O_45,N_2970,N_2955);
nand UO_46 (O_46,N_2977,N_2992);
or UO_47 (O_47,N_2960,N_2954);
or UO_48 (O_48,N_2978,N_2997);
or UO_49 (O_49,N_2971,N_2962);
nand UO_50 (O_50,N_2986,N_2978);
nand UO_51 (O_51,N_2986,N_2962);
xor UO_52 (O_52,N_2975,N_2962);
and UO_53 (O_53,N_2995,N_2981);
nor UO_54 (O_54,N_2985,N_2983);
or UO_55 (O_55,N_2991,N_2967);
xnor UO_56 (O_56,N_2982,N_2953);
or UO_57 (O_57,N_2975,N_2950);
or UO_58 (O_58,N_2980,N_2985);
nor UO_59 (O_59,N_2971,N_2965);
nand UO_60 (O_60,N_2994,N_2976);
or UO_61 (O_61,N_2992,N_2993);
and UO_62 (O_62,N_2995,N_2969);
nor UO_63 (O_63,N_2950,N_2961);
and UO_64 (O_64,N_2981,N_2955);
or UO_65 (O_65,N_2970,N_2980);
or UO_66 (O_66,N_2969,N_2989);
and UO_67 (O_67,N_2987,N_2966);
nor UO_68 (O_68,N_2961,N_2984);
nand UO_69 (O_69,N_2987,N_2962);
nor UO_70 (O_70,N_2975,N_2963);
nand UO_71 (O_71,N_2959,N_2969);
and UO_72 (O_72,N_2985,N_2959);
nor UO_73 (O_73,N_2950,N_2987);
or UO_74 (O_74,N_2982,N_2956);
or UO_75 (O_75,N_2986,N_2953);
nand UO_76 (O_76,N_2984,N_2972);
and UO_77 (O_77,N_2954,N_2988);
or UO_78 (O_78,N_2968,N_2982);
nand UO_79 (O_79,N_2979,N_2971);
and UO_80 (O_80,N_2988,N_2965);
nor UO_81 (O_81,N_2957,N_2996);
nand UO_82 (O_82,N_2979,N_2981);
or UO_83 (O_83,N_2961,N_2960);
and UO_84 (O_84,N_2981,N_2997);
nor UO_85 (O_85,N_2959,N_2980);
nand UO_86 (O_86,N_2986,N_2959);
or UO_87 (O_87,N_2980,N_2994);
xor UO_88 (O_88,N_2969,N_2998);
xor UO_89 (O_89,N_2974,N_2999);
and UO_90 (O_90,N_2997,N_2985);
or UO_91 (O_91,N_2993,N_2965);
and UO_92 (O_92,N_2972,N_2987);
nand UO_93 (O_93,N_2973,N_2970);
and UO_94 (O_94,N_2967,N_2993);
nand UO_95 (O_95,N_2981,N_2994);
nor UO_96 (O_96,N_2972,N_2980);
xor UO_97 (O_97,N_2954,N_2971);
and UO_98 (O_98,N_2952,N_2981);
and UO_99 (O_99,N_2987,N_2968);
nor UO_100 (O_100,N_2994,N_2970);
nor UO_101 (O_101,N_2958,N_2969);
and UO_102 (O_102,N_2951,N_2999);
and UO_103 (O_103,N_2970,N_2992);
nor UO_104 (O_104,N_2953,N_2950);
nor UO_105 (O_105,N_2958,N_2952);
xor UO_106 (O_106,N_2964,N_2975);
nand UO_107 (O_107,N_2993,N_2998);
or UO_108 (O_108,N_2965,N_2991);
nand UO_109 (O_109,N_2990,N_2955);
nor UO_110 (O_110,N_2976,N_2989);
nor UO_111 (O_111,N_2971,N_2958);
nor UO_112 (O_112,N_2962,N_2973);
xnor UO_113 (O_113,N_2972,N_2981);
nand UO_114 (O_114,N_2984,N_2990);
nor UO_115 (O_115,N_2963,N_2966);
or UO_116 (O_116,N_2962,N_2972);
nand UO_117 (O_117,N_2955,N_2961);
and UO_118 (O_118,N_2963,N_2976);
or UO_119 (O_119,N_2952,N_2995);
xor UO_120 (O_120,N_2960,N_2967);
and UO_121 (O_121,N_2964,N_2965);
nand UO_122 (O_122,N_2977,N_2986);
nand UO_123 (O_123,N_2950,N_2992);
and UO_124 (O_124,N_2957,N_2964);
or UO_125 (O_125,N_2972,N_2960);
and UO_126 (O_126,N_2958,N_2990);
and UO_127 (O_127,N_2954,N_2965);
and UO_128 (O_128,N_2975,N_2953);
nand UO_129 (O_129,N_2958,N_2996);
and UO_130 (O_130,N_2984,N_2981);
nand UO_131 (O_131,N_2989,N_2979);
nand UO_132 (O_132,N_2951,N_2953);
xor UO_133 (O_133,N_2984,N_2966);
nand UO_134 (O_134,N_2997,N_2964);
nor UO_135 (O_135,N_2978,N_2950);
and UO_136 (O_136,N_2976,N_2977);
xor UO_137 (O_137,N_2985,N_2990);
or UO_138 (O_138,N_2981,N_2953);
or UO_139 (O_139,N_2990,N_2951);
or UO_140 (O_140,N_2994,N_2951);
nor UO_141 (O_141,N_2987,N_2984);
or UO_142 (O_142,N_2982,N_2964);
and UO_143 (O_143,N_2970,N_2953);
xnor UO_144 (O_144,N_2954,N_2958);
nand UO_145 (O_145,N_2976,N_2980);
nand UO_146 (O_146,N_2983,N_2962);
nand UO_147 (O_147,N_2996,N_2968);
or UO_148 (O_148,N_2966,N_2979);
and UO_149 (O_149,N_2968,N_2980);
and UO_150 (O_150,N_2997,N_2969);
nand UO_151 (O_151,N_2993,N_2973);
nor UO_152 (O_152,N_2968,N_2991);
xnor UO_153 (O_153,N_2981,N_2996);
and UO_154 (O_154,N_2958,N_2961);
or UO_155 (O_155,N_2984,N_2954);
or UO_156 (O_156,N_2971,N_2957);
nand UO_157 (O_157,N_2966,N_2982);
nor UO_158 (O_158,N_2959,N_2958);
or UO_159 (O_159,N_2952,N_2959);
nand UO_160 (O_160,N_2977,N_2952);
and UO_161 (O_161,N_2985,N_2984);
nor UO_162 (O_162,N_2972,N_2953);
and UO_163 (O_163,N_2989,N_2951);
nand UO_164 (O_164,N_2973,N_2988);
and UO_165 (O_165,N_2969,N_2954);
nor UO_166 (O_166,N_2988,N_2978);
nor UO_167 (O_167,N_2952,N_2969);
nand UO_168 (O_168,N_2960,N_2979);
or UO_169 (O_169,N_2961,N_2997);
nand UO_170 (O_170,N_2951,N_2970);
nor UO_171 (O_171,N_2950,N_2976);
nor UO_172 (O_172,N_2972,N_2983);
nor UO_173 (O_173,N_2967,N_2992);
nand UO_174 (O_174,N_2996,N_2960);
nand UO_175 (O_175,N_2971,N_2994);
or UO_176 (O_176,N_2986,N_2985);
nand UO_177 (O_177,N_2978,N_2987);
and UO_178 (O_178,N_2962,N_2964);
or UO_179 (O_179,N_2999,N_2972);
nand UO_180 (O_180,N_2969,N_2975);
xor UO_181 (O_181,N_2956,N_2981);
and UO_182 (O_182,N_2969,N_2996);
nor UO_183 (O_183,N_2985,N_2977);
or UO_184 (O_184,N_2982,N_2993);
xnor UO_185 (O_185,N_2969,N_2962);
and UO_186 (O_186,N_2963,N_2957);
or UO_187 (O_187,N_2967,N_2999);
or UO_188 (O_188,N_2956,N_2961);
or UO_189 (O_189,N_2967,N_2977);
xnor UO_190 (O_190,N_2998,N_2964);
nand UO_191 (O_191,N_2973,N_2976);
and UO_192 (O_192,N_2997,N_2996);
and UO_193 (O_193,N_2999,N_2996);
and UO_194 (O_194,N_2959,N_2954);
and UO_195 (O_195,N_2972,N_2982);
and UO_196 (O_196,N_2957,N_2983);
xnor UO_197 (O_197,N_2975,N_2977);
nor UO_198 (O_198,N_2963,N_2978);
xnor UO_199 (O_199,N_2992,N_2984);
and UO_200 (O_200,N_2975,N_2970);
and UO_201 (O_201,N_2970,N_2961);
nor UO_202 (O_202,N_2990,N_2966);
or UO_203 (O_203,N_2952,N_2973);
nand UO_204 (O_204,N_2954,N_2995);
nor UO_205 (O_205,N_2974,N_2967);
and UO_206 (O_206,N_2958,N_2983);
nand UO_207 (O_207,N_2994,N_2972);
nand UO_208 (O_208,N_2995,N_2985);
nor UO_209 (O_209,N_2999,N_2962);
xnor UO_210 (O_210,N_2997,N_2988);
and UO_211 (O_211,N_2950,N_2979);
or UO_212 (O_212,N_2974,N_2969);
or UO_213 (O_213,N_2987,N_2974);
nor UO_214 (O_214,N_2990,N_2973);
nor UO_215 (O_215,N_2961,N_2964);
nand UO_216 (O_216,N_2978,N_2976);
nand UO_217 (O_217,N_2998,N_2961);
or UO_218 (O_218,N_2953,N_2992);
and UO_219 (O_219,N_2974,N_2979);
nor UO_220 (O_220,N_2997,N_2983);
nand UO_221 (O_221,N_2992,N_2956);
and UO_222 (O_222,N_2988,N_2977);
nor UO_223 (O_223,N_2985,N_2989);
or UO_224 (O_224,N_2974,N_2989);
nor UO_225 (O_225,N_2991,N_2976);
nand UO_226 (O_226,N_2979,N_2964);
nand UO_227 (O_227,N_2991,N_2953);
nand UO_228 (O_228,N_2992,N_2980);
nand UO_229 (O_229,N_2996,N_2972);
and UO_230 (O_230,N_2955,N_2992);
nand UO_231 (O_231,N_2954,N_2972);
nor UO_232 (O_232,N_2954,N_2992);
nor UO_233 (O_233,N_2959,N_2973);
and UO_234 (O_234,N_2993,N_2981);
nor UO_235 (O_235,N_2969,N_2983);
nand UO_236 (O_236,N_2998,N_2971);
nand UO_237 (O_237,N_2967,N_2963);
or UO_238 (O_238,N_2998,N_2988);
and UO_239 (O_239,N_2970,N_2991);
or UO_240 (O_240,N_2962,N_2995);
and UO_241 (O_241,N_2951,N_2960);
and UO_242 (O_242,N_2992,N_2971);
nand UO_243 (O_243,N_2972,N_2979);
nand UO_244 (O_244,N_2995,N_2958);
nor UO_245 (O_245,N_2960,N_2999);
nand UO_246 (O_246,N_2995,N_2961);
nand UO_247 (O_247,N_2973,N_2968);
nor UO_248 (O_248,N_2995,N_2998);
or UO_249 (O_249,N_2979,N_2973);
nand UO_250 (O_250,N_2999,N_2970);
nor UO_251 (O_251,N_2969,N_2961);
nand UO_252 (O_252,N_2983,N_2967);
xnor UO_253 (O_253,N_2998,N_2965);
nand UO_254 (O_254,N_2958,N_2992);
nor UO_255 (O_255,N_2977,N_2973);
nor UO_256 (O_256,N_2999,N_2958);
or UO_257 (O_257,N_2985,N_2960);
nand UO_258 (O_258,N_2965,N_2997);
and UO_259 (O_259,N_2999,N_2995);
or UO_260 (O_260,N_2993,N_2963);
and UO_261 (O_261,N_2956,N_2955);
nand UO_262 (O_262,N_2991,N_2994);
or UO_263 (O_263,N_2955,N_2985);
or UO_264 (O_264,N_2990,N_2974);
or UO_265 (O_265,N_2995,N_2950);
nand UO_266 (O_266,N_2972,N_2952);
or UO_267 (O_267,N_2979,N_2953);
xnor UO_268 (O_268,N_2963,N_2987);
xor UO_269 (O_269,N_2966,N_2954);
and UO_270 (O_270,N_2965,N_2951);
nand UO_271 (O_271,N_2995,N_2991);
nand UO_272 (O_272,N_2986,N_2956);
or UO_273 (O_273,N_2984,N_2963);
or UO_274 (O_274,N_2982,N_2977);
nand UO_275 (O_275,N_2990,N_2986);
and UO_276 (O_276,N_2982,N_2961);
xnor UO_277 (O_277,N_2952,N_2991);
nand UO_278 (O_278,N_2986,N_2982);
nand UO_279 (O_279,N_2983,N_2996);
nand UO_280 (O_280,N_2961,N_2951);
nor UO_281 (O_281,N_2978,N_2965);
nand UO_282 (O_282,N_2981,N_2951);
nand UO_283 (O_283,N_2959,N_2955);
or UO_284 (O_284,N_2954,N_2961);
and UO_285 (O_285,N_2963,N_2959);
nand UO_286 (O_286,N_2973,N_2955);
nand UO_287 (O_287,N_2967,N_2966);
nand UO_288 (O_288,N_2987,N_2954);
or UO_289 (O_289,N_2961,N_2980);
and UO_290 (O_290,N_2959,N_2972);
and UO_291 (O_291,N_2956,N_2975);
nand UO_292 (O_292,N_2971,N_2966);
or UO_293 (O_293,N_2985,N_2963);
or UO_294 (O_294,N_2991,N_2951);
or UO_295 (O_295,N_2993,N_2955);
nor UO_296 (O_296,N_2998,N_2990);
nand UO_297 (O_297,N_2950,N_2971);
nand UO_298 (O_298,N_2982,N_2980);
or UO_299 (O_299,N_2980,N_2998);
or UO_300 (O_300,N_2969,N_2951);
nand UO_301 (O_301,N_2976,N_2968);
nand UO_302 (O_302,N_2957,N_2959);
nand UO_303 (O_303,N_2952,N_2988);
nand UO_304 (O_304,N_2962,N_2952);
nand UO_305 (O_305,N_2997,N_2989);
nor UO_306 (O_306,N_2991,N_2959);
and UO_307 (O_307,N_2973,N_2997);
nor UO_308 (O_308,N_2965,N_2957);
xor UO_309 (O_309,N_2995,N_2963);
or UO_310 (O_310,N_2960,N_2977);
or UO_311 (O_311,N_2996,N_2988);
nor UO_312 (O_312,N_2955,N_2982);
nand UO_313 (O_313,N_2964,N_2970);
and UO_314 (O_314,N_2962,N_2961);
xnor UO_315 (O_315,N_2954,N_2981);
nand UO_316 (O_316,N_2979,N_2956);
nor UO_317 (O_317,N_2964,N_2993);
nand UO_318 (O_318,N_2964,N_2963);
and UO_319 (O_319,N_2991,N_2999);
nor UO_320 (O_320,N_2950,N_2996);
xor UO_321 (O_321,N_2961,N_2952);
nand UO_322 (O_322,N_2995,N_2986);
nor UO_323 (O_323,N_2974,N_2993);
or UO_324 (O_324,N_2950,N_2969);
and UO_325 (O_325,N_2982,N_2974);
nor UO_326 (O_326,N_2957,N_2993);
nand UO_327 (O_327,N_2956,N_2974);
and UO_328 (O_328,N_2983,N_2971);
nor UO_329 (O_329,N_2998,N_2970);
nor UO_330 (O_330,N_2950,N_2951);
or UO_331 (O_331,N_2957,N_2974);
or UO_332 (O_332,N_2993,N_2954);
nand UO_333 (O_333,N_2963,N_2965);
or UO_334 (O_334,N_2973,N_2984);
and UO_335 (O_335,N_2996,N_2953);
nand UO_336 (O_336,N_2989,N_2971);
nand UO_337 (O_337,N_2983,N_2980);
nor UO_338 (O_338,N_2950,N_2964);
and UO_339 (O_339,N_2975,N_2957);
and UO_340 (O_340,N_2980,N_2952);
nand UO_341 (O_341,N_2963,N_2972);
or UO_342 (O_342,N_2986,N_2993);
and UO_343 (O_343,N_2963,N_2998);
and UO_344 (O_344,N_2998,N_2996);
nor UO_345 (O_345,N_2965,N_2986);
and UO_346 (O_346,N_2971,N_2961);
and UO_347 (O_347,N_2962,N_2990);
xnor UO_348 (O_348,N_2955,N_2971);
or UO_349 (O_349,N_2976,N_2992);
and UO_350 (O_350,N_2959,N_2982);
or UO_351 (O_351,N_2991,N_2990);
or UO_352 (O_352,N_2965,N_2994);
and UO_353 (O_353,N_2955,N_2999);
nor UO_354 (O_354,N_2986,N_2991);
nand UO_355 (O_355,N_2960,N_2982);
nand UO_356 (O_356,N_2975,N_2980);
nor UO_357 (O_357,N_2986,N_2998);
nor UO_358 (O_358,N_2988,N_2987);
or UO_359 (O_359,N_2956,N_2954);
nand UO_360 (O_360,N_2980,N_2988);
or UO_361 (O_361,N_2995,N_2971);
and UO_362 (O_362,N_2988,N_2969);
xnor UO_363 (O_363,N_2955,N_2997);
or UO_364 (O_364,N_2963,N_2951);
or UO_365 (O_365,N_2977,N_2953);
nor UO_366 (O_366,N_2992,N_2959);
xor UO_367 (O_367,N_2984,N_2976);
nand UO_368 (O_368,N_2954,N_2985);
and UO_369 (O_369,N_2987,N_2991);
and UO_370 (O_370,N_2987,N_2956);
or UO_371 (O_371,N_2976,N_2959);
nand UO_372 (O_372,N_2987,N_2996);
or UO_373 (O_373,N_2974,N_2977);
nand UO_374 (O_374,N_2974,N_2973);
nor UO_375 (O_375,N_2991,N_2966);
nor UO_376 (O_376,N_2968,N_2959);
xnor UO_377 (O_377,N_2990,N_2956);
xor UO_378 (O_378,N_2985,N_2996);
nor UO_379 (O_379,N_2961,N_2994);
or UO_380 (O_380,N_2975,N_2982);
or UO_381 (O_381,N_2988,N_2961);
nor UO_382 (O_382,N_2963,N_2992);
nand UO_383 (O_383,N_2990,N_2961);
nand UO_384 (O_384,N_2984,N_2959);
nand UO_385 (O_385,N_2968,N_2986);
nand UO_386 (O_386,N_2987,N_2970);
or UO_387 (O_387,N_2983,N_2976);
xor UO_388 (O_388,N_2951,N_2983);
and UO_389 (O_389,N_2978,N_2985);
and UO_390 (O_390,N_2952,N_2990);
or UO_391 (O_391,N_2998,N_2951);
nor UO_392 (O_392,N_2988,N_2950);
nand UO_393 (O_393,N_2997,N_2958);
xor UO_394 (O_394,N_2985,N_2962);
nor UO_395 (O_395,N_2952,N_2984);
nor UO_396 (O_396,N_2986,N_2961);
nor UO_397 (O_397,N_2976,N_2972);
nor UO_398 (O_398,N_2965,N_2961);
nor UO_399 (O_399,N_2957,N_2977);
nand UO_400 (O_400,N_2988,N_2971);
nand UO_401 (O_401,N_2955,N_2996);
and UO_402 (O_402,N_2960,N_2953);
nor UO_403 (O_403,N_2959,N_2995);
and UO_404 (O_404,N_2958,N_2989);
nor UO_405 (O_405,N_2985,N_2975);
xnor UO_406 (O_406,N_2950,N_2983);
xnor UO_407 (O_407,N_2999,N_2950);
or UO_408 (O_408,N_2991,N_2996);
xnor UO_409 (O_409,N_2978,N_2977);
nor UO_410 (O_410,N_2961,N_2976);
nor UO_411 (O_411,N_2969,N_2999);
nand UO_412 (O_412,N_2981,N_2988);
and UO_413 (O_413,N_2994,N_2987);
or UO_414 (O_414,N_2979,N_2969);
and UO_415 (O_415,N_2992,N_2979);
xnor UO_416 (O_416,N_2965,N_2983);
or UO_417 (O_417,N_2991,N_2989);
and UO_418 (O_418,N_2964,N_2958);
xor UO_419 (O_419,N_2990,N_2957);
or UO_420 (O_420,N_2968,N_2961);
and UO_421 (O_421,N_2962,N_2951);
nor UO_422 (O_422,N_2984,N_2998);
nor UO_423 (O_423,N_2989,N_2968);
xor UO_424 (O_424,N_2994,N_2986);
nand UO_425 (O_425,N_2970,N_2954);
nand UO_426 (O_426,N_2977,N_2966);
nor UO_427 (O_427,N_2998,N_2975);
nor UO_428 (O_428,N_2958,N_2988);
or UO_429 (O_429,N_2999,N_2979);
nand UO_430 (O_430,N_2955,N_2958);
nor UO_431 (O_431,N_2965,N_2979);
or UO_432 (O_432,N_2968,N_2997);
nor UO_433 (O_433,N_2999,N_2978);
and UO_434 (O_434,N_2995,N_2980);
or UO_435 (O_435,N_2970,N_2997);
nand UO_436 (O_436,N_2999,N_2953);
or UO_437 (O_437,N_2992,N_2983);
nand UO_438 (O_438,N_2980,N_2990);
nor UO_439 (O_439,N_2972,N_2964);
xor UO_440 (O_440,N_2970,N_2985);
nand UO_441 (O_441,N_2979,N_2998);
nor UO_442 (O_442,N_2964,N_2971);
or UO_443 (O_443,N_2961,N_2987);
or UO_444 (O_444,N_2972,N_2985);
and UO_445 (O_445,N_2995,N_2976);
nor UO_446 (O_446,N_2985,N_2952);
and UO_447 (O_447,N_2981,N_2982);
nor UO_448 (O_448,N_2957,N_2995);
and UO_449 (O_449,N_2961,N_2966);
and UO_450 (O_450,N_2978,N_2955);
xor UO_451 (O_451,N_2962,N_2974);
and UO_452 (O_452,N_2956,N_2959);
nor UO_453 (O_453,N_2958,N_2991);
xnor UO_454 (O_454,N_2993,N_2994);
nor UO_455 (O_455,N_2985,N_2971);
or UO_456 (O_456,N_2972,N_2993);
or UO_457 (O_457,N_2974,N_2952);
and UO_458 (O_458,N_2956,N_2971);
and UO_459 (O_459,N_2970,N_2984);
and UO_460 (O_460,N_2984,N_2962);
nand UO_461 (O_461,N_2964,N_2978);
and UO_462 (O_462,N_2954,N_2963);
and UO_463 (O_463,N_2975,N_2988);
or UO_464 (O_464,N_2950,N_2993);
and UO_465 (O_465,N_2975,N_2976);
nor UO_466 (O_466,N_2976,N_2955);
nand UO_467 (O_467,N_2984,N_2978);
nor UO_468 (O_468,N_2999,N_2975);
and UO_469 (O_469,N_2977,N_2950);
nor UO_470 (O_470,N_2974,N_2972);
nor UO_471 (O_471,N_2974,N_2971);
nor UO_472 (O_472,N_2961,N_2957);
and UO_473 (O_473,N_2952,N_2957);
and UO_474 (O_474,N_2961,N_2989);
and UO_475 (O_475,N_2975,N_2995);
nor UO_476 (O_476,N_2956,N_2962);
xnor UO_477 (O_477,N_2952,N_2978);
nor UO_478 (O_478,N_2993,N_2962);
nor UO_479 (O_479,N_2995,N_2993);
and UO_480 (O_480,N_2990,N_2963);
nor UO_481 (O_481,N_2986,N_2960);
nand UO_482 (O_482,N_2985,N_2950);
nor UO_483 (O_483,N_2993,N_2951);
or UO_484 (O_484,N_2961,N_2974);
and UO_485 (O_485,N_2966,N_2965);
xnor UO_486 (O_486,N_2975,N_2991);
nand UO_487 (O_487,N_2953,N_2952);
nand UO_488 (O_488,N_2952,N_2994);
xor UO_489 (O_489,N_2962,N_2980);
and UO_490 (O_490,N_2973,N_2966);
nor UO_491 (O_491,N_2988,N_2983);
or UO_492 (O_492,N_2960,N_2958);
and UO_493 (O_493,N_2968,N_2952);
and UO_494 (O_494,N_2968,N_2998);
and UO_495 (O_495,N_2991,N_2993);
nor UO_496 (O_496,N_2973,N_2992);
and UO_497 (O_497,N_2995,N_2955);
xor UO_498 (O_498,N_2957,N_2989);
or UO_499 (O_499,N_2950,N_2968);
endmodule