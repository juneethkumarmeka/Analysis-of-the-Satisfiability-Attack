module basic_500_3000_500_60_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_70,In_303);
and U1 (N_1,In_329,In_345);
or U2 (N_2,In_230,In_170);
or U3 (N_3,In_359,In_293);
nor U4 (N_4,In_256,In_200);
or U5 (N_5,In_182,In_415);
and U6 (N_6,In_444,In_31);
nor U7 (N_7,In_274,In_458);
and U8 (N_8,In_78,In_499);
nor U9 (N_9,In_349,In_355);
or U10 (N_10,In_314,In_111);
and U11 (N_11,In_337,In_72);
or U12 (N_12,In_203,In_442);
nand U13 (N_13,In_350,In_243);
or U14 (N_14,In_33,In_232);
nand U15 (N_15,In_65,In_172);
nand U16 (N_16,In_16,In_259);
nor U17 (N_17,In_432,In_177);
and U18 (N_18,In_436,In_235);
nor U19 (N_19,In_375,In_196);
or U20 (N_20,In_422,In_416);
or U21 (N_21,In_66,In_454);
nand U22 (N_22,In_231,In_245);
nand U23 (N_23,In_338,In_204);
nand U24 (N_24,In_282,In_437);
nor U25 (N_25,In_478,In_294);
nand U26 (N_26,In_205,In_276);
or U27 (N_27,In_175,In_41);
nand U28 (N_28,In_58,In_236);
or U29 (N_29,In_164,In_197);
or U30 (N_30,In_108,In_192);
nor U31 (N_31,In_138,In_174);
nand U32 (N_32,In_409,In_448);
and U33 (N_33,In_77,In_107);
and U34 (N_34,In_430,In_412);
nor U35 (N_35,In_456,In_250);
and U36 (N_36,In_191,In_494);
nand U37 (N_37,In_307,In_17);
or U38 (N_38,In_268,In_263);
nand U39 (N_39,In_424,In_308);
or U40 (N_40,In_91,In_376);
nand U41 (N_41,In_275,In_278);
nand U42 (N_42,In_149,In_301);
nand U43 (N_43,In_21,In_215);
nor U44 (N_44,In_207,In_106);
xnor U45 (N_45,In_486,In_98);
nand U46 (N_46,In_132,In_109);
or U47 (N_47,In_71,In_162);
nand U48 (N_48,In_300,In_488);
nor U49 (N_49,In_470,In_369);
nand U50 (N_50,In_96,In_285);
nand U51 (N_51,In_194,In_325);
and U52 (N_52,In_469,In_117);
nand U53 (N_53,In_403,In_311);
and U54 (N_54,In_479,In_52);
nor U55 (N_55,In_63,N_40);
or U56 (N_56,In_159,In_210);
and U57 (N_57,In_328,In_119);
or U58 (N_58,In_114,In_160);
and U59 (N_59,In_103,In_10);
or U60 (N_60,In_62,In_26);
or U61 (N_61,In_372,N_30);
or U62 (N_62,N_44,In_187);
nor U63 (N_63,In_11,In_9);
xnor U64 (N_64,In_429,In_116);
nor U65 (N_65,In_130,In_227);
nand U66 (N_66,In_397,In_356);
or U67 (N_67,N_41,In_330);
and U68 (N_68,In_90,In_425);
nand U69 (N_69,In_420,In_485);
and U70 (N_70,In_99,In_333);
or U71 (N_71,In_457,In_118);
nor U72 (N_72,In_441,In_241);
nand U73 (N_73,In_36,In_100);
or U74 (N_74,In_147,In_392);
nor U75 (N_75,In_321,N_38);
nand U76 (N_76,In_168,In_340);
nand U77 (N_77,In_343,In_380);
and U78 (N_78,In_451,In_377);
or U79 (N_79,In_497,In_83);
nor U80 (N_80,In_466,In_29);
nand U81 (N_81,In_51,In_59);
nand U82 (N_82,N_45,In_190);
nor U83 (N_83,N_19,In_292);
or U84 (N_84,In_492,In_133);
and U85 (N_85,In_223,In_153);
or U86 (N_86,In_411,In_89);
nor U87 (N_87,In_323,N_46);
nor U88 (N_88,In_439,In_453);
nand U89 (N_89,In_154,In_1);
and U90 (N_90,In_379,N_4);
nand U91 (N_91,In_296,In_125);
or U92 (N_92,In_348,In_25);
and U93 (N_93,In_87,In_84);
nand U94 (N_94,In_247,In_105);
nor U95 (N_95,In_265,In_421);
or U96 (N_96,In_319,In_487);
nor U97 (N_97,In_364,In_324);
nor U98 (N_98,In_94,In_352);
or U99 (N_99,N_3,In_463);
or U100 (N_100,In_68,In_0);
nor U101 (N_101,In_178,In_67);
nand U102 (N_102,In_316,In_326);
nor U103 (N_103,In_244,In_135);
nand U104 (N_104,In_13,In_373);
nand U105 (N_105,N_47,In_201);
and U106 (N_106,In_385,In_123);
and U107 (N_107,In_277,In_242);
or U108 (N_108,In_495,In_389);
nor U109 (N_109,N_2,In_490);
or U110 (N_110,N_98,In_279);
or U111 (N_111,In_28,In_185);
or U112 (N_112,In_295,N_60);
nor U113 (N_113,In_336,In_262);
nor U114 (N_114,In_370,In_95);
or U115 (N_115,In_386,In_347);
and U116 (N_116,In_237,N_62);
and U117 (N_117,In_433,N_7);
nor U118 (N_118,In_381,In_391);
or U119 (N_119,In_388,In_47);
nand U120 (N_120,N_27,N_31);
xor U121 (N_121,N_81,In_461);
nor U122 (N_122,N_33,In_408);
nor U123 (N_123,N_14,N_59);
nor U124 (N_124,In_428,In_334);
nand U125 (N_125,In_335,In_327);
nand U126 (N_126,In_60,N_8);
nand U127 (N_127,In_110,In_46);
and U128 (N_128,In_393,In_213);
nor U129 (N_129,In_53,In_155);
and U130 (N_130,N_28,In_362);
and U131 (N_131,In_418,N_56);
nand U132 (N_132,In_146,In_6);
nand U133 (N_133,In_360,In_30);
or U134 (N_134,In_248,In_88);
or U135 (N_135,N_93,In_158);
and U136 (N_136,N_99,N_69);
nand U137 (N_137,In_225,N_96);
nor U138 (N_138,In_413,In_73);
nand U139 (N_139,In_150,In_289);
and U140 (N_140,N_12,In_43);
and U141 (N_141,In_167,In_419);
nand U142 (N_142,In_198,In_3);
nor U143 (N_143,In_212,In_234);
nand U144 (N_144,In_404,In_214);
or U145 (N_145,In_179,In_183);
nor U146 (N_146,In_216,In_305);
nor U147 (N_147,N_76,In_86);
and U148 (N_148,In_208,In_222);
nor U149 (N_149,N_97,In_280);
nor U150 (N_150,In_417,In_4);
nand U151 (N_151,In_38,In_173);
nor U152 (N_152,In_383,In_131);
and U153 (N_153,N_89,N_29);
nor U154 (N_154,In_189,In_56);
nand U155 (N_155,In_465,In_396);
and U156 (N_156,In_140,N_71);
or U157 (N_157,In_332,N_13);
or U158 (N_158,In_122,N_142);
or U159 (N_159,In_440,In_163);
and U160 (N_160,In_474,In_137);
and U161 (N_161,In_165,In_407);
nor U162 (N_162,N_24,N_132);
nor U163 (N_163,N_91,In_134);
or U164 (N_164,N_139,In_42);
nor U165 (N_165,N_140,N_105);
nor U166 (N_166,N_135,In_384);
nand U167 (N_167,In_353,In_483);
and U168 (N_168,In_287,N_53);
or U169 (N_169,In_218,N_67);
or U170 (N_170,In_374,In_156);
and U171 (N_171,N_88,N_10);
nand U172 (N_172,In_450,In_171);
nor U173 (N_173,In_476,N_55);
nor U174 (N_174,In_166,N_123);
nand U175 (N_175,In_283,In_498);
nor U176 (N_176,In_2,In_446);
and U177 (N_177,In_272,In_310);
or U178 (N_178,N_74,In_306);
and U179 (N_179,In_5,In_447);
and U180 (N_180,In_127,N_43);
xnor U181 (N_181,N_79,In_239);
or U182 (N_182,In_129,In_217);
nor U183 (N_183,In_312,In_322);
or U184 (N_184,In_351,In_79);
nor U185 (N_185,In_142,In_493);
and U186 (N_186,In_102,N_136);
nor U187 (N_187,In_228,In_291);
and U188 (N_188,In_199,N_23);
and U189 (N_189,In_346,N_83);
or U190 (N_190,In_271,N_32);
nor U191 (N_191,In_115,N_108);
and U192 (N_192,In_368,In_249);
or U193 (N_193,In_423,N_149);
nand U194 (N_194,In_378,In_357);
nor U195 (N_195,N_94,In_240);
and U196 (N_196,N_6,In_206);
or U197 (N_197,In_258,In_452);
nor U198 (N_198,In_126,In_462);
nand U199 (N_199,In_286,In_169);
nor U200 (N_200,N_95,N_72);
and U201 (N_201,N_115,N_145);
and U202 (N_202,In_298,In_246);
nor U203 (N_203,In_69,In_35);
nand U204 (N_204,N_101,In_61);
and U205 (N_205,N_36,N_82);
or U206 (N_206,N_131,In_139);
nor U207 (N_207,N_18,In_220);
and U208 (N_208,In_226,N_78);
and U209 (N_209,In_398,In_431);
and U210 (N_210,In_434,In_24);
or U211 (N_211,In_64,In_7);
nand U212 (N_212,In_443,N_16);
nand U213 (N_213,In_57,In_75);
or U214 (N_214,In_85,N_117);
nor U215 (N_215,In_233,N_143);
or U216 (N_216,In_157,In_290);
nand U217 (N_217,In_427,N_63);
nand U218 (N_218,In_181,In_317);
and U219 (N_219,N_66,In_15);
and U220 (N_220,N_21,N_130);
or U221 (N_221,In_363,N_195);
or U222 (N_222,In_238,N_174);
and U223 (N_223,In_460,N_39);
nand U224 (N_224,In_395,N_154);
nor U225 (N_225,In_148,In_184);
nor U226 (N_226,In_54,In_401);
nor U227 (N_227,N_197,In_475);
xnor U228 (N_228,In_270,In_113);
and U229 (N_229,N_86,In_19);
and U230 (N_230,In_136,N_156);
nand U231 (N_231,N_17,N_118);
nand U232 (N_232,N_119,N_34);
or U233 (N_233,In_82,In_34);
nand U234 (N_234,N_150,In_315);
nor U235 (N_235,N_15,In_438);
nor U236 (N_236,N_172,In_406);
and U237 (N_237,In_44,In_101);
and U238 (N_238,In_331,In_55);
nor U239 (N_239,In_304,N_90);
nand U240 (N_240,In_18,N_58);
or U241 (N_241,N_198,N_193);
or U242 (N_242,N_80,In_354);
nand U243 (N_243,N_87,N_114);
nor U244 (N_244,In_124,N_102);
and U245 (N_245,In_161,In_382);
nor U246 (N_246,In_209,N_75);
and U247 (N_247,In_402,In_266);
nor U248 (N_248,In_477,N_129);
nand U249 (N_249,N_1,N_169);
nand U250 (N_250,N_122,N_121);
and U251 (N_251,In_313,In_358);
nor U252 (N_252,In_180,In_484);
and U253 (N_253,N_162,N_37);
and U254 (N_254,N_240,N_225);
and U255 (N_255,In_471,In_459);
or U256 (N_256,In_387,N_217);
or U257 (N_257,In_144,N_51);
nand U258 (N_258,N_220,N_109);
nor U259 (N_259,In_405,N_179);
nand U260 (N_260,N_168,N_227);
or U261 (N_261,N_104,In_297);
nand U262 (N_262,In_48,N_167);
or U263 (N_263,N_64,N_85);
nand U264 (N_264,N_20,N_232);
or U265 (N_265,N_222,N_247);
nand U266 (N_266,N_107,N_204);
nand U267 (N_267,In_202,N_180);
nand U268 (N_268,N_170,In_344);
and U269 (N_269,In_302,N_190);
or U270 (N_270,N_201,N_181);
or U271 (N_271,In_39,In_341);
nand U272 (N_272,N_185,In_467);
nand U273 (N_273,In_414,N_9);
nor U274 (N_274,N_157,In_219);
or U275 (N_275,N_236,N_235);
and U276 (N_276,In_50,N_160);
or U277 (N_277,In_472,In_253);
and U278 (N_278,In_40,In_361);
nor U279 (N_279,N_120,In_112);
nor U280 (N_280,In_27,In_320);
nand U281 (N_281,N_245,N_70);
or U282 (N_282,In_97,In_37);
and U283 (N_283,In_390,In_366);
or U284 (N_284,N_158,N_242);
nor U285 (N_285,In_81,N_147);
nand U286 (N_286,N_113,In_12);
and U287 (N_287,N_212,N_210);
nor U288 (N_288,N_183,N_228);
nand U289 (N_289,In_365,N_133);
and U290 (N_290,N_188,In_455);
nor U291 (N_291,N_249,In_141);
or U292 (N_292,N_22,In_257);
or U293 (N_293,N_112,In_254);
or U294 (N_294,In_435,N_239);
nand U295 (N_295,N_178,N_173);
or U296 (N_296,In_221,N_134);
nor U297 (N_297,In_152,N_126);
and U298 (N_298,N_208,N_244);
nor U299 (N_299,N_231,N_243);
xnor U300 (N_300,N_260,N_25);
or U301 (N_301,N_296,In_273);
nand U302 (N_302,In_464,In_318);
and U303 (N_303,In_473,N_148);
and U304 (N_304,N_233,N_237);
and U305 (N_305,N_229,N_138);
nor U306 (N_306,N_262,N_161);
or U307 (N_307,N_214,N_238);
nand U308 (N_308,In_128,N_137);
or U309 (N_309,N_146,N_152);
or U310 (N_310,In_20,N_230);
nor U311 (N_311,N_246,N_277);
or U312 (N_312,N_106,In_186);
nor U313 (N_313,N_209,N_290);
or U314 (N_314,N_186,N_287);
nor U315 (N_315,N_207,N_216);
and U316 (N_316,N_153,N_268);
and U317 (N_317,In_23,In_400);
nand U318 (N_318,N_298,N_92);
nor U319 (N_319,In_143,N_151);
nand U320 (N_320,In_145,N_276);
nand U321 (N_321,N_111,N_211);
nand U322 (N_322,In_426,N_289);
or U323 (N_323,N_282,N_255);
and U324 (N_324,In_399,N_166);
nand U325 (N_325,N_175,N_241);
nand U326 (N_326,In_22,N_159);
xnor U327 (N_327,N_73,N_253);
or U328 (N_328,In_371,In_480);
nor U329 (N_329,In_32,N_57);
nand U330 (N_330,N_199,In_489);
and U331 (N_331,In_482,N_219);
nor U332 (N_332,In_288,N_49);
nand U333 (N_333,N_294,N_125);
and U334 (N_334,N_250,In_491);
nand U335 (N_335,In_121,N_165);
and U336 (N_336,N_65,N_280);
nor U337 (N_337,N_61,N_110);
or U338 (N_338,N_256,N_77);
and U339 (N_339,N_295,N_144);
or U340 (N_340,N_297,In_260);
nor U341 (N_341,In_281,N_213);
nand U342 (N_342,N_215,In_188);
nor U343 (N_343,N_251,N_171);
nand U344 (N_344,N_35,N_155);
nor U345 (N_345,N_270,N_182);
and U346 (N_346,N_252,N_259);
and U347 (N_347,In_229,N_278);
or U348 (N_348,In_74,N_52);
and U349 (N_349,N_248,N_267);
and U350 (N_350,N_319,N_189);
and U351 (N_351,N_338,N_321);
or U352 (N_352,In_176,N_288);
nand U353 (N_353,N_336,In_151);
and U354 (N_354,N_283,N_347);
or U355 (N_355,N_272,In_195);
or U356 (N_356,N_324,In_468);
nor U357 (N_357,N_164,N_48);
and U358 (N_358,N_26,N_285);
or U359 (N_359,N_275,N_258);
nor U360 (N_360,N_325,N_0);
nor U361 (N_361,N_265,N_322);
or U362 (N_362,N_192,N_292);
nor U363 (N_363,N_42,N_263);
nand U364 (N_364,N_274,N_266);
nand U365 (N_365,N_330,In_76);
and U366 (N_366,In_267,In_299);
and U367 (N_367,N_320,In_252);
or U368 (N_368,N_346,N_286);
or U369 (N_369,In_445,In_93);
or U370 (N_370,N_218,N_5);
nor U371 (N_371,N_176,In_342);
or U372 (N_372,N_329,In_367);
and U373 (N_373,N_331,N_203);
or U374 (N_374,N_333,In_92);
and U375 (N_375,N_340,N_341);
nor U376 (N_376,N_317,N_221);
or U377 (N_377,N_206,N_348);
or U378 (N_378,N_163,N_54);
or U379 (N_379,N_327,In_120);
or U380 (N_380,N_307,N_226);
and U381 (N_381,N_128,N_343);
nor U382 (N_382,N_315,N_205);
or U383 (N_383,N_345,N_202);
nor U384 (N_384,N_187,N_284);
nor U385 (N_385,In_193,N_124);
nand U386 (N_386,N_300,In_104);
nand U387 (N_387,N_257,N_306);
nand U388 (N_388,N_339,N_271);
nand U389 (N_389,N_100,In_80);
and U390 (N_390,N_309,N_264);
and U391 (N_391,In_211,N_328);
nand U392 (N_392,In_410,N_184);
nand U393 (N_393,N_127,N_196);
nor U394 (N_394,In_264,N_141);
or U395 (N_395,N_299,N_68);
or U396 (N_396,N_84,N_191);
and U397 (N_397,N_308,In_309);
nor U398 (N_398,N_314,N_301);
and U399 (N_399,N_200,N_316);
and U400 (N_400,N_354,N_223);
and U401 (N_401,N_355,N_384);
and U402 (N_402,N_303,N_358);
nand U403 (N_403,N_360,N_305);
or U404 (N_404,In_481,N_273);
or U405 (N_405,N_385,N_312);
nand U406 (N_406,N_291,N_310);
and U407 (N_407,N_335,N_334);
or U408 (N_408,N_234,N_382);
or U409 (N_409,N_365,N_361);
nand U410 (N_410,N_372,In_49);
nor U411 (N_411,N_391,N_374);
nand U412 (N_412,In_269,N_387);
and U413 (N_413,N_376,N_375);
or U414 (N_414,N_381,N_386);
or U415 (N_415,N_395,In_284);
nand U416 (N_416,N_397,N_116);
or U417 (N_417,N_279,N_311);
or U418 (N_418,N_293,N_351);
nor U419 (N_419,N_370,N_367);
nand U420 (N_420,In_394,In_496);
nor U421 (N_421,In_261,In_251);
and U422 (N_422,N_302,N_326);
and U423 (N_423,N_396,N_362);
or U424 (N_424,N_254,N_379);
nand U425 (N_425,N_378,N_323);
or U426 (N_426,N_389,N_398);
nand U427 (N_427,N_224,N_380);
nor U428 (N_428,N_392,N_177);
nor U429 (N_429,N_342,N_364);
nor U430 (N_430,In_339,In_255);
or U431 (N_431,N_369,In_224);
or U432 (N_432,N_350,N_11);
or U433 (N_433,N_103,N_383);
nor U434 (N_434,N_332,N_353);
and U435 (N_435,N_269,N_352);
nor U436 (N_436,N_50,N_363);
nor U437 (N_437,In_14,N_281);
or U438 (N_438,N_388,N_394);
nor U439 (N_439,N_349,N_313);
nand U440 (N_440,N_368,N_390);
or U441 (N_441,N_359,N_304);
and U442 (N_442,N_377,N_366);
nand U443 (N_443,In_8,N_337);
or U444 (N_444,N_399,N_393);
nor U445 (N_445,In_45,N_318);
and U446 (N_446,N_357,N_371);
nand U447 (N_447,In_449,N_356);
or U448 (N_448,N_344,N_373);
nand U449 (N_449,N_194,N_261);
nand U450 (N_450,N_444,N_447);
nor U451 (N_451,N_434,N_436);
and U452 (N_452,N_449,N_407);
nor U453 (N_453,N_426,N_400);
nand U454 (N_454,N_440,N_419);
nor U455 (N_455,N_416,N_424);
nand U456 (N_456,N_420,N_405);
nand U457 (N_457,N_425,N_401);
and U458 (N_458,N_414,N_430);
nor U459 (N_459,N_442,N_415);
or U460 (N_460,N_417,N_432);
nor U461 (N_461,N_429,N_441);
or U462 (N_462,N_404,N_439);
nand U463 (N_463,N_410,N_437);
and U464 (N_464,N_408,N_445);
and U465 (N_465,N_431,N_448);
nand U466 (N_466,N_438,N_403);
and U467 (N_467,N_413,N_422);
nor U468 (N_468,N_443,N_418);
or U469 (N_469,N_446,N_402);
nand U470 (N_470,N_428,N_423);
nand U471 (N_471,N_435,N_433);
or U472 (N_472,N_409,N_406);
and U473 (N_473,N_412,N_411);
nor U474 (N_474,N_421,N_427);
and U475 (N_475,N_411,N_432);
nand U476 (N_476,N_429,N_414);
and U477 (N_477,N_446,N_433);
nor U478 (N_478,N_428,N_424);
nand U479 (N_479,N_402,N_440);
or U480 (N_480,N_407,N_421);
or U481 (N_481,N_432,N_425);
and U482 (N_482,N_445,N_427);
or U483 (N_483,N_404,N_402);
and U484 (N_484,N_413,N_438);
nand U485 (N_485,N_405,N_441);
and U486 (N_486,N_435,N_407);
nand U487 (N_487,N_414,N_410);
or U488 (N_488,N_434,N_407);
and U489 (N_489,N_419,N_437);
and U490 (N_490,N_417,N_408);
nand U491 (N_491,N_443,N_446);
nand U492 (N_492,N_444,N_446);
or U493 (N_493,N_428,N_448);
or U494 (N_494,N_428,N_427);
xor U495 (N_495,N_416,N_409);
or U496 (N_496,N_407,N_444);
and U497 (N_497,N_410,N_416);
xor U498 (N_498,N_417,N_434);
xor U499 (N_499,N_432,N_414);
or U500 (N_500,N_486,N_493);
nor U501 (N_501,N_482,N_459);
nor U502 (N_502,N_487,N_478);
and U503 (N_503,N_484,N_471);
nand U504 (N_504,N_480,N_460);
nor U505 (N_505,N_475,N_464);
or U506 (N_506,N_470,N_458);
nand U507 (N_507,N_455,N_463);
and U508 (N_508,N_479,N_473);
or U509 (N_509,N_497,N_495);
or U510 (N_510,N_476,N_467);
nor U511 (N_511,N_454,N_492);
nand U512 (N_512,N_466,N_468);
and U513 (N_513,N_477,N_450);
and U514 (N_514,N_474,N_491);
and U515 (N_515,N_481,N_457);
nand U516 (N_516,N_465,N_456);
xor U517 (N_517,N_498,N_485);
or U518 (N_518,N_488,N_499);
nand U519 (N_519,N_452,N_451);
nor U520 (N_520,N_496,N_472);
nand U521 (N_521,N_489,N_461);
nand U522 (N_522,N_462,N_469);
nor U523 (N_523,N_490,N_453);
nand U524 (N_524,N_483,N_494);
or U525 (N_525,N_454,N_499);
and U526 (N_526,N_466,N_493);
nor U527 (N_527,N_492,N_487);
or U528 (N_528,N_491,N_478);
or U529 (N_529,N_468,N_490);
or U530 (N_530,N_454,N_450);
and U531 (N_531,N_491,N_486);
or U532 (N_532,N_473,N_450);
nor U533 (N_533,N_494,N_491);
and U534 (N_534,N_483,N_469);
and U535 (N_535,N_493,N_463);
or U536 (N_536,N_475,N_499);
nand U537 (N_537,N_471,N_480);
and U538 (N_538,N_495,N_469);
and U539 (N_539,N_459,N_483);
or U540 (N_540,N_450,N_463);
or U541 (N_541,N_485,N_455);
and U542 (N_542,N_492,N_498);
and U543 (N_543,N_493,N_462);
nor U544 (N_544,N_489,N_496);
nand U545 (N_545,N_494,N_485);
nand U546 (N_546,N_469,N_484);
nor U547 (N_547,N_476,N_462);
nand U548 (N_548,N_479,N_483);
or U549 (N_549,N_494,N_484);
nand U550 (N_550,N_503,N_541);
or U551 (N_551,N_514,N_542);
nor U552 (N_552,N_529,N_540);
and U553 (N_553,N_546,N_531);
nor U554 (N_554,N_535,N_523);
nor U555 (N_555,N_534,N_533);
nor U556 (N_556,N_547,N_532);
nand U557 (N_557,N_513,N_522);
nor U558 (N_558,N_528,N_521);
or U559 (N_559,N_525,N_548);
xor U560 (N_560,N_519,N_527);
nor U561 (N_561,N_505,N_511);
nand U562 (N_562,N_549,N_536);
nor U563 (N_563,N_501,N_517);
or U564 (N_564,N_545,N_500);
nor U565 (N_565,N_543,N_516);
and U566 (N_566,N_539,N_504);
and U567 (N_567,N_538,N_537);
or U568 (N_568,N_508,N_526);
nor U569 (N_569,N_518,N_510);
nand U570 (N_570,N_515,N_512);
and U571 (N_571,N_506,N_524);
nand U572 (N_572,N_530,N_509);
or U573 (N_573,N_544,N_502);
nor U574 (N_574,N_520,N_507);
and U575 (N_575,N_515,N_535);
nor U576 (N_576,N_538,N_530);
or U577 (N_577,N_518,N_548);
and U578 (N_578,N_527,N_545);
and U579 (N_579,N_506,N_536);
and U580 (N_580,N_518,N_543);
or U581 (N_581,N_543,N_510);
nor U582 (N_582,N_517,N_523);
or U583 (N_583,N_529,N_521);
or U584 (N_584,N_545,N_516);
and U585 (N_585,N_544,N_510);
or U586 (N_586,N_527,N_539);
nand U587 (N_587,N_521,N_546);
and U588 (N_588,N_518,N_531);
nand U589 (N_589,N_520,N_527);
or U590 (N_590,N_503,N_500);
and U591 (N_591,N_526,N_533);
and U592 (N_592,N_543,N_500);
nand U593 (N_593,N_508,N_527);
and U594 (N_594,N_542,N_516);
nand U595 (N_595,N_539,N_511);
or U596 (N_596,N_542,N_549);
nand U597 (N_597,N_534,N_532);
and U598 (N_598,N_533,N_521);
nand U599 (N_599,N_545,N_530);
and U600 (N_600,N_551,N_589);
or U601 (N_601,N_590,N_550);
or U602 (N_602,N_594,N_593);
nor U603 (N_603,N_581,N_553);
or U604 (N_604,N_576,N_562);
nand U605 (N_605,N_554,N_586);
and U606 (N_606,N_575,N_570);
or U607 (N_607,N_556,N_573);
nor U608 (N_608,N_565,N_572);
nand U609 (N_609,N_574,N_587);
nand U610 (N_610,N_588,N_571);
and U611 (N_611,N_557,N_577);
nor U612 (N_612,N_569,N_591);
or U613 (N_613,N_596,N_592);
and U614 (N_614,N_583,N_558);
and U615 (N_615,N_598,N_579);
nand U616 (N_616,N_563,N_564);
nand U617 (N_617,N_566,N_552);
nor U618 (N_618,N_585,N_560);
nand U619 (N_619,N_568,N_555);
nor U620 (N_620,N_599,N_559);
nand U621 (N_621,N_561,N_595);
nor U622 (N_622,N_578,N_584);
nor U623 (N_623,N_580,N_597);
nor U624 (N_624,N_567,N_582);
or U625 (N_625,N_551,N_585);
nor U626 (N_626,N_553,N_579);
and U627 (N_627,N_587,N_572);
or U628 (N_628,N_575,N_563);
nand U629 (N_629,N_553,N_596);
nor U630 (N_630,N_562,N_561);
and U631 (N_631,N_592,N_594);
nand U632 (N_632,N_597,N_573);
nand U633 (N_633,N_553,N_582);
and U634 (N_634,N_591,N_588);
nor U635 (N_635,N_578,N_562);
or U636 (N_636,N_572,N_591);
nand U637 (N_637,N_591,N_555);
nor U638 (N_638,N_599,N_552);
nand U639 (N_639,N_561,N_559);
nor U640 (N_640,N_577,N_585);
or U641 (N_641,N_573,N_588);
nor U642 (N_642,N_596,N_586);
nor U643 (N_643,N_556,N_553);
nand U644 (N_644,N_577,N_574);
nor U645 (N_645,N_574,N_583);
nand U646 (N_646,N_595,N_569);
and U647 (N_647,N_590,N_568);
nand U648 (N_648,N_566,N_573);
or U649 (N_649,N_576,N_586);
nor U650 (N_650,N_643,N_613);
nand U651 (N_651,N_620,N_624);
or U652 (N_652,N_600,N_633);
or U653 (N_653,N_623,N_630);
nand U654 (N_654,N_635,N_646);
and U655 (N_655,N_638,N_602);
nand U656 (N_656,N_601,N_622);
and U657 (N_657,N_621,N_612);
nor U658 (N_658,N_618,N_609);
and U659 (N_659,N_617,N_627);
nand U660 (N_660,N_614,N_605);
nor U661 (N_661,N_644,N_639);
nor U662 (N_662,N_645,N_615);
or U663 (N_663,N_608,N_641);
nand U664 (N_664,N_642,N_603);
nand U665 (N_665,N_606,N_625);
and U666 (N_666,N_632,N_628);
nand U667 (N_667,N_634,N_648);
nand U668 (N_668,N_616,N_640);
or U669 (N_669,N_631,N_626);
nand U670 (N_670,N_647,N_637);
or U671 (N_671,N_636,N_611);
or U672 (N_672,N_619,N_604);
xnor U673 (N_673,N_629,N_649);
or U674 (N_674,N_610,N_607);
and U675 (N_675,N_619,N_643);
nand U676 (N_676,N_603,N_625);
or U677 (N_677,N_611,N_645);
or U678 (N_678,N_632,N_640);
and U679 (N_679,N_600,N_638);
nor U680 (N_680,N_633,N_611);
nor U681 (N_681,N_631,N_605);
or U682 (N_682,N_630,N_642);
and U683 (N_683,N_633,N_626);
nor U684 (N_684,N_607,N_620);
or U685 (N_685,N_642,N_643);
and U686 (N_686,N_646,N_612);
nand U687 (N_687,N_630,N_604);
nor U688 (N_688,N_607,N_633);
nand U689 (N_689,N_629,N_616);
nand U690 (N_690,N_636,N_642);
and U691 (N_691,N_649,N_626);
or U692 (N_692,N_601,N_640);
nand U693 (N_693,N_634,N_612);
and U694 (N_694,N_618,N_635);
or U695 (N_695,N_625,N_622);
and U696 (N_696,N_619,N_602);
and U697 (N_697,N_614,N_606);
or U698 (N_698,N_647,N_616);
nand U699 (N_699,N_639,N_645);
nor U700 (N_700,N_675,N_676);
and U701 (N_701,N_671,N_654);
and U702 (N_702,N_660,N_668);
or U703 (N_703,N_680,N_674);
or U704 (N_704,N_663,N_678);
and U705 (N_705,N_677,N_670);
or U706 (N_706,N_661,N_697);
nor U707 (N_707,N_653,N_679);
nand U708 (N_708,N_667,N_662);
and U709 (N_709,N_652,N_696);
or U710 (N_710,N_683,N_694);
and U711 (N_711,N_699,N_657);
nand U712 (N_712,N_655,N_673);
or U713 (N_713,N_682,N_651);
or U714 (N_714,N_664,N_698);
nor U715 (N_715,N_672,N_690);
and U716 (N_716,N_669,N_691);
or U717 (N_717,N_665,N_689);
or U718 (N_718,N_686,N_656);
or U719 (N_719,N_693,N_685);
nor U720 (N_720,N_650,N_684);
nor U721 (N_721,N_687,N_695);
nor U722 (N_722,N_666,N_681);
nand U723 (N_723,N_658,N_659);
and U724 (N_724,N_688,N_692);
nand U725 (N_725,N_688,N_667);
nand U726 (N_726,N_667,N_650);
and U727 (N_727,N_690,N_661);
nand U728 (N_728,N_686,N_678);
nor U729 (N_729,N_675,N_698);
and U730 (N_730,N_684,N_662);
and U731 (N_731,N_674,N_650);
or U732 (N_732,N_650,N_686);
nor U733 (N_733,N_696,N_662);
and U734 (N_734,N_698,N_693);
nand U735 (N_735,N_692,N_670);
or U736 (N_736,N_672,N_699);
and U737 (N_737,N_658,N_681);
nand U738 (N_738,N_666,N_698);
nand U739 (N_739,N_654,N_664);
nor U740 (N_740,N_670,N_655);
and U741 (N_741,N_655,N_681);
nand U742 (N_742,N_668,N_659);
nand U743 (N_743,N_662,N_654);
nor U744 (N_744,N_664,N_656);
nand U745 (N_745,N_690,N_675);
and U746 (N_746,N_677,N_686);
or U747 (N_747,N_696,N_675);
nor U748 (N_748,N_673,N_686);
nor U749 (N_749,N_678,N_666);
and U750 (N_750,N_728,N_746);
or U751 (N_751,N_726,N_715);
nand U752 (N_752,N_700,N_744);
or U753 (N_753,N_704,N_742);
and U754 (N_754,N_734,N_741);
or U755 (N_755,N_738,N_732);
nand U756 (N_756,N_703,N_747);
nor U757 (N_757,N_737,N_721);
nand U758 (N_758,N_727,N_709);
nor U759 (N_759,N_730,N_739);
and U760 (N_760,N_710,N_717);
nor U761 (N_761,N_712,N_722);
nor U762 (N_762,N_723,N_740);
nor U763 (N_763,N_705,N_713);
nand U764 (N_764,N_711,N_706);
nor U765 (N_765,N_731,N_720);
or U766 (N_766,N_724,N_749);
nand U767 (N_767,N_701,N_707);
and U768 (N_768,N_708,N_718);
nand U769 (N_769,N_733,N_736);
or U770 (N_770,N_714,N_716);
nand U771 (N_771,N_725,N_719);
nand U772 (N_772,N_748,N_735);
nand U773 (N_773,N_729,N_702);
xnor U774 (N_774,N_745,N_743);
or U775 (N_775,N_728,N_740);
or U776 (N_776,N_745,N_709);
and U777 (N_777,N_708,N_748);
nor U778 (N_778,N_721,N_734);
or U779 (N_779,N_740,N_730);
and U780 (N_780,N_716,N_703);
nand U781 (N_781,N_713,N_714);
nand U782 (N_782,N_709,N_735);
nand U783 (N_783,N_721,N_711);
nor U784 (N_784,N_742,N_726);
nor U785 (N_785,N_746,N_703);
or U786 (N_786,N_739,N_705);
and U787 (N_787,N_731,N_749);
or U788 (N_788,N_715,N_705);
nand U789 (N_789,N_710,N_716);
nor U790 (N_790,N_708,N_716);
nand U791 (N_791,N_725,N_730);
nor U792 (N_792,N_729,N_747);
nand U793 (N_793,N_732,N_727);
or U794 (N_794,N_745,N_713);
and U795 (N_795,N_747,N_709);
and U796 (N_796,N_745,N_719);
nor U797 (N_797,N_747,N_724);
and U798 (N_798,N_705,N_703);
or U799 (N_799,N_738,N_731);
nand U800 (N_800,N_799,N_788);
nand U801 (N_801,N_776,N_764);
nand U802 (N_802,N_786,N_771);
or U803 (N_803,N_793,N_781);
nand U804 (N_804,N_756,N_794);
nor U805 (N_805,N_765,N_782);
and U806 (N_806,N_766,N_790);
or U807 (N_807,N_780,N_785);
and U808 (N_808,N_783,N_774);
nor U809 (N_809,N_778,N_784);
or U810 (N_810,N_792,N_750);
nor U811 (N_811,N_761,N_757);
or U812 (N_812,N_796,N_791);
nand U813 (N_813,N_773,N_779);
nand U814 (N_814,N_753,N_775);
or U815 (N_815,N_798,N_760);
and U816 (N_816,N_795,N_752);
and U817 (N_817,N_755,N_762);
nand U818 (N_818,N_769,N_787);
nand U819 (N_819,N_751,N_759);
nand U820 (N_820,N_770,N_797);
or U821 (N_821,N_768,N_754);
or U822 (N_822,N_789,N_767);
and U823 (N_823,N_758,N_772);
or U824 (N_824,N_763,N_777);
or U825 (N_825,N_787,N_770);
nand U826 (N_826,N_779,N_759);
nand U827 (N_827,N_762,N_770);
nand U828 (N_828,N_764,N_781);
and U829 (N_829,N_761,N_783);
and U830 (N_830,N_787,N_764);
or U831 (N_831,N_763,N_779);
nor U832 (N_832,N_751,N_795);
or U833 (N_833,N_762,N_756);
and U834 (N_834,N_781,N_761);
nor U835 (N_835,N_775,N_755);
or U836 (N_836,N_787,N_782);
nand U837 (N_837,N_792,N_798);
or U838 (N_838,N_790,N_756);
nor U839 (N_839,N_777,N_752);
or U840 (N_840,N_778,N_777);
nor U841 (N_841,N_782,N_751);
nand U842 (N_842,N_764,N_763);
nand U843 (N_843,N_757,N_768);
nor U844 (N_844,N_767,N_775);
nand U845 (N_845,N_791,N_765);
or U846 (N_846,N_798,N_799);
nor U847 (N_847,N_755,N_779);
nand U848 (N_848,N_780,N_750);
or U849 (N_849,N_772,N_778);
nand U850 (N_850,N_803,N_843);
or U851 (N_851,N_849,N_816);
nand U852 (N_852,N_801,N_847);
or U853 (N_853,N_825,N_835);
and U854 (N_854,N_810,N_844);
nor U855 (N_855,N_808,N_815);
nand U856 (N_856,N_837,N_814);
nand U857 (N_857,N_845,N_846);
or U858 (N_858,N_820,N_827);
nor U859 (N_859,N_826,N_830);
or U860 (N_860,N_834,N_838);
nor U861 (N_861,N_817,N_805);
nand U862 (N_862,N_833,N_813);
nand U863 (N_863,N_823,N_839);
or U864 (N_864,N_831,N_821);
nand U865 (N_865,N_800,N_818);
nand U866 (N_866,N_822,N_804);
nand U867 (N_867,N_829,N_812);
xor U868 (N_868,N_811,N_807);
or U869 (N_869,N_806,N_841);
nor U870 (N_870,N_840,N_802);
or U871 (N_871,N_848,N_832);
nand U872 (N_872,N_842,N_836);
nand U873 (N_873,N_824,N_809);
or U874 (N_874,N_828,N_819);
and U875 (N_875,N_843,N_807);
nor U876 (N_876,N_801,N_813);
or U877 (N_877,N_842,N_823);
or U878 (N_878,N_810,N_827);
nand U879 (N_879,N_800,N_820);
or U880 (N_880,N_849,N_824);
nand U881 (N_881,N_826,N_816);
and U882 (N_882,N_805,N_803);
and U883 (N_883,N_813,N_808);
nand U884 (N_884,N_840,N_803);
nor U885 (N_885,N_821,N_822);
nand U886 (N_886,N_809,N_837);
and U887 (N_887,N_808,N_846);
nor U888 (N_888,N_818,N_808);
nor U889 (N_889,N_818,N_835);
nand U890 (N_890,N_810,N_816);
nand U891 (N_891,N_807,N_848);
or U892 (N_892,N_843,N_823);
or U893 (N_893,N_826,N_809);
or U894 (N_894,N_844,N_824);
and U895 (N_895,N_807,N_809);
and U896 (N_896,N_801,N_821);
nor U897 (N_897,N_805,N_845);
or U898 (N_898,N_839,N_804);
nor U899 (N_899,N_818,N_848);
and U900 (N_900,N_889,N_878);
and U901 (N_901,N_859,N_873);
and U902 (N_902,N_877,N_851);
nand U903 (N_903,N_881,N_895);
nor U904 (N_904,N_894,N_866);
or U905 (N_905,N_869,N_880);
or U906 (N_906,N_879,N_898);
and U907 (N_907,N_890,N_891);
and U908 (N_908,N_882,N_850);
and U909 (N_909,N_857,N_864);
nand U910 (N_910,N_855,N_896);
nand U911 (N_911,N_856,N_858);
nand U912 (N_912,N_892,N_875);
nand U913 (N_913,N_868,N_852);
nor U914 (N_914,N_853,N_865);
nor U915 (N_915,N_854,N_888);
and U916 (N_916,N_867,N_860);
xnor U917 (N_917,N_897,N_870);
and U918 (N_918,N_884,N_871);
nand U919 (N_919,N_862,N_861);
and U920 (N_920,N_885,N_876);
and U921 (N_921,N_893,N_887);
xor U922 (N_922,N_899,N_883);
nor U923 (N_923,N_872,N_874);
and U924 (N_924,N_886,N_863);
or U925 (N_925,N_869,N_855);
nand U926 (N_926,N_891,N_857);
nor U927 (N_927,N_893,N_891);
nor U928 (N_928,N_857,N_889);
nand U929 (N_929,N_879,N_856);
nor U930 (N_930,N_894,N_899);
or U931 (N_931,N_871,N_891);
and U932 (N_932,N_862,N_893);
nand U933 (N_933,N_881,N_890);
or U934 (N_934,N_884,N_895);
nor U935 (N_935,N_866,N_853);
nor U936 (N_936,N_876,N_867);
nand U937 (N_937,N_857,N_877);
and U938 (N_938,N_865,N_889);
nor U939 (N_939,N_873,N_852);
and U940 (N_940,N_883,N_882);
or U941 (N_941,N_893,N_858);
nor U942 (N_942,N_872,N_882);
or U943 (N_943,N_856,N_864);
nor U944 (N_944,N_894,N_887);
nand U945 (N_945,N_868,N_887);
nor U946 (N_946,N_869,N_887);
nor U947 (N_947,N_897,N_894);
nor U948 (N_948,N_873,N_892);
xnor U949 (N_949,N_864,N_882);
nor U950 (N_950,N_933,N_947);
nand U951 (N_951,N_944,N_915);
nand U952 (N_952,N_943,N_922);
nand U953 (N_953,N_917,N_936);
or U954 (N_954,N_905,N_910);
or U955 (N_955,N_901,N_945);
nor U956 (N_956,N_900,N_921);
and U957 (N_957,N_919,N_928);
and U958 (N_958,N_949,N_932);
nor U959 (N_959,N_912,N_906);
nand U960 (N_960,N_942,N_904);
nor U961 (N_961,N_924,N_940);
nand U962 (N_962,N_930,N_925);
nand U963 (N_963,N_941,N_926);
and U964 (N_964,N_931,N_914);
nand U965 (N_965,N_935,N_946);
and U966 (N_966,N_908,N_927);
nand U967 (N_967,N_937,N_918);
and U968 (N_968,N_929,N_920);
xor U969 (N_969,N_902,N_934);
nor U970 (N_970,N_911,N_907);
nor U971 (N_971,N_948,N_916);
nand U972 (N_972,N_938,N_923);
and U973 (N_973,N_939,N_903);
and U974 (N_974,N_909,N_913);
and U975 (N_975,N_924,N_922);
or U976 (N_976,N_907,N_930);
nor U977 (N_977,N_934,N_915);
nor U978 (N_978,N_925,N_905);
and U979 (N_979,N_926,N_909);
and U980 (N_980,N_917,N_915);
nor U981 (N_981,N_933,N_937);
or U982 (N_982,N_920,N_940);
and U983 (N_983,N_911,N_910);
or U984 (N_984,N_933,N_932);
and U985 (N_985,N_935,N_932);
and U986 (N_986,N_909,N_906);
or U987 (N_987,N_911,N_906);
and U988 (N_988,N_910,N_938);
nor U989 (N_989,N_930,N_949);
or U990 (N_990,N_934,N_941);
or U991 (N_991,N_942,N_920);
or U992 (N_992,N_909,N_940);
or U993 (N_993,N_911,N_908);
or U994 (N_994,N_901,N_908);
nor U995 (N_995,N_911,N_939);
nand U996 (N_996,N_936,N_941);
nand U997 (N_997,N_911,N_914);
or U998 (N_998,N_946,N_928);
or U999 (N_999,N_945,N_920);
and U1000 (N_1000,N_967,N_972);
nor U1001 (N_1001,N_973,N_960);
nand U1002 (N_1002,N_963,N_952);
or U1003 (N_1003,N_968,N_951);
nor U1004 (N_1004,N_987,N_990);
nor U1005 (N_1005,N_996,N_955);
and U1006 (N_1006,N_985,N_954);
nand U1007 (N_1007,N_964,N_991);
and U1008 (N_1008,N_988,N_957);
or U1009 (N_1009,N_998,N_980);
nor U1010 (N_1010,N_969,N_995);
nor U1011 (N_1011,N_974,N_999);
nand U1012 (N_1012,N_961,N_966);
nor U1013 (N_1013,N_994,N_981);
nor U1014 (N_1014,N_978,N_959);
nand U1015 (N_1015,N_984,N_989);
nor U1016 (N_1016,N_983,N_970);
nand U1017 (N_1017,N_962,N_977);
and U1018 (N_1018,N_971,N_997);
nor U1019 (N_1019,N_958,N_956);
nand U1020 (N_1020,N_982,N_953);
nor U1021 (N_1021,N_979,N_975);
and U1022 (N_1022,N_992,N_976);
or U1023 (N_1023,N_986,N_965);
nor U1024 (N_1024,N_993,N_950);
nand U1025 (N_1025,N_952,N_982);
and U1026 (N_1026,N_956,N_960);
or U1027 (N_1027,N_990,N_994);
or U1028 (N_1028,N_981,N_971);
xor U1029 (N_1029,N_983,N_995);
nor U1030 (N_1030,N_975,N_952);
nand U1031 (N_1031,N_987,N_978);
or U1032 (N_1032,N_958,N_989);
and U1033 (N_1033,N_999,N_992);
and U1034 (N_1034,N_976,N_984);
nor U1035 (N_1035,N_973,N_956);
nor U1036 (N_1036,N_959,N_990);
nand U1037 (N_1037,N_996,N_973);
nor U1038 (N_1038,N_979,N_960);
nand U1039 (N_1039,N_998,N_974);
and U1040 (N_1040,N_975,N_969);
or U1041 (N_1041,N_968,N_986);
and U1042 (N_1042,N_997,N_995);
nand U1043 (N_1043,N_970,N_964);
or U1044 (N_1044,N_974,N_970);
and U1045 (N_1045,N_987,N_995);
nor U1046 (N_1046,N_957,N_961);
and U1047 (N_1047,N_990,N_956);
nand U1048 (N_1048,N_993,N_982);
or U1049 (N_1049,N_988,N_966);
or U1050 (N_1050,N_1035,N_1016);
nand U1051 (N_1051,N_1030,N_1024);
nor U1052 (N_1052,N_1003,N_1040);
nand U1053 (N_1053,N_1048,N_1044);
nand U1054 (N_1054,N_1005,N_1017);
and U1055 (N_1055,N_1000,N_1036);
and U1056 (N_1056,N_1027,N_1034);
nor U1057 (N_1057,N_1032,N_1025);
nand U1058 (N_1058,N_1013,N_1014);
or U1059 (N_1059,N_1041,N_1037);
and U1060 (N_1060,N_1038,N_1043);
nand U1061 (N_1061,N_1011,N_1018);
and U1062 (N_1062,N_1020,N_1010);
and U1063 (N_1063,N_1033,N_1007);
nand U1064 (N_1064,N_1001,N_1012);
or U1065 (N_1065,N_1015,N_1049);
and U1066 (N_1066,N_1045,N_1006);
nand U1067 (N_1067,N_1029,N_1019);
nand U1068 (N_1068,N_1039,N_1031);
or U1069 (N_1069,N_1028,N_1023);
nand U1070 (N_1070,N_1047,N_1021);
and U1071 (N_1071,N_1022,N_1026);
nand U1072 (N_1072,N_1046,N_1008);
or U1073 (N_1073,N_1009,N_1004);
or U1074 (N_1074,N_1002,N_1042);
and U1075 (N_1075,N_1031,N_1038);
and U1076 (N_1076,N_1036,N_1023);
nand U1077 (N_1077,N_1037,N_1040);
and U1078 (N_1078,N_1041,N_1007);
and U1079 (N_1079,N_1003,N_1041);
and U1080 (N_1080,N_1026,N_1047);
nand U1081 (N_1081,N_1025,N_1046);
and U1082 (N_1082,N_1044,N_1027);
nor U1083 (N_1083,N_1004,N_1031);
or U1084 (N_1084,N_1045,N_1033);
nand U1085 (N_1085,N_1021,N_1048);
or U1086 (N_1086,N_1048,N_1020);
nand U1087 (N_1087,N_1006,N_1036);
nand U1088 (N_1088,N_1046,N_1017);
and U1089 (N_1089,N_1032,N_1036);
nand U1090 (N_1090,N_1031,N_1019);
or U1091 (N_1091,N_1025,N_1033);
nor U1092 (N_1092,N_1047,N_1028);
nand U1093 (N_1093,N_1001,N_1002);
or U1094 (N_1094,N_1031,N_1018);
and U1095 (N_1095,N_1029,N_1009);
and U1096 (N_1096,N_1005,N_1018);
and U1097 (N_1097,N_1048,N_1006);
and U1098 (N_1098,N_1043,N_1005);
nand U1099 (N_1099,N_1004,N_1013);
nor U1100 (N_1100,N_1067,N_1079);
or U1101 (N_1101,N_1053,N_1091);
nand U1102 (N_1102,N_1075,N_1087);
nand U1103 (N_1103,N_1098,N_1057);
nor U1104 (N_1104,N_1051,N_1059);
nor U1105 (N_1105,N_1061,N_1052);
and U1106 (N_1106,N_1095,N_1063);
nand U1107 (N_1107,N_1076,N_1097);
and U1108 (N_1108,N_1093,N_1078);
and U1109 (N_1109,N_1064,N_1086);
or U1110 (N_1110,N_1084,N_1055);
xnor U1111 (N_1111,N_1071,N_1070);
or U1112 (N_1112,N_1066,N_1099);
and U1113 (N_1113,N_1056,N_1062);
nor U1114 (N_1114,N_1082,N_1088);
and U1115 (N_1115,N_1054,N_1077);
nor U1116 (N_1116,N_1090,N_1050);
and U1117 (N_1117,N_1073,N_1085);
and U1118 (N_1118,N_1081,N_1068);
nor U1119 (N_1119,N_1069,N_1089);
nor U1120 (N_1120,N_1065,N_1094);
nand U1121 (N_1121,N_1058,N_1092);
or U1122 (N_1122,N_1060,N_1083);
nor U1123 (N_1123,N_1080,N_1074);
nand U1124 (N_1124,N_1096,N_1072);
or U1125 (N_1125,N_1060,N_1074);
nand U1126 (N_1126,N_1084,N_1080);
or U1127 (N_1127,N_1092,N_1070);
nor U1128 (N_1128,N_1063,N_1099);
nand U1129 (N_1129,N_1073,N_1062);
nand U1130 (N_1130,N_1065,N_1095);
and U1131 (N_1131,N_1073,N_1052);
nor U1132 (N_1132,N_1055,N_1058);
nand U1133 (N_1133,N_1052,N_1091);
nor U1134 (N_1134,N_1090,N_1092);
or U1135 (N_1135,N_1057,N_1066);
nor U1136 (N_1136,N_1083,N_1074);
and U1137 (N_1137,N_1089,N_1057);
and U1138 (N_1138,N_1058,N_1076);
nand U1139 (N_1139,N_1059,N_1064);
and U1140 (N_1140,N_1095,N_1050);
xnor U1141 (N_1141,N_1059,N_1076);
or U1142 (N_1142,N_1086,N_1052);
or U1143 (N_1143,N_1066,N_1095);
nand U1144 (N_1144,N_1073,N_1069);
or U1145 (N_1145,N_1086,N_1085);
nor U1146 (N_1146,N_1099,N_1072);
nand U1147 (N_1147,N_1053,N_1050);
or U1148 (N_1148,N_1056,N_1053);
nor U1149 (N_1149,N_1054,N_1078);
nand U1150 (N_1150,N_1100,N_1123);
or U1151 (N_1151,N_1101,N_1125);
nand U1152 (N_1152,N_1108,N_1106);
nor U1153 (N_1153,N_1140,N_1126);
nand U1154 (N_1154,N_1131,N_1127);
nor U1155 (N_1155,N_1109,N_1112);
or U1156 (N_1156,N_1111,N_1143);
or U1157 (N_1157,N_1144,N_1117);
and U1158 (N_1158,N_1118,N_1149);
or U1159 (N_1159,N_1138,N_1114);
and U1160 (N_1160,N_1119,N_1102);
nand U1161 (N_1161,N_1121,N_1103);
nand U1162 (N_1162,N_1122,N_1129);
and U1163 (N_1163,N_1104,N_1116);
or U1164 (N_1164,N_1142,N_1132);
nor U1165 (N_1165,N_1148,N_1128);
nor U1166 (N_1166,N_1141,N_1145);
nor U1167 (N_1167,N_1135,N_1113);
nand U1168 (N_1168,N_1137,N_1134);
nor U1169 (N_1169,N_1120,N_1146);
nand U1170 (N_1170,N_1147,N_1136);
nor U1171 (N_1171,N_1110,N_1105);
nand U1172 (N_1172,N_1133,N_1107);
nand U1173 (N_1173,N_1124,N_1130);
and U1174 (N_1174,N_1139,N_1115);
and U1175 (N_1175,N_1111,N_1118);
nand U1176 (N_1176,N_1100,N_1146);
nor U1177 (N_1177,N_1133,N_1141);
nand U1178 (N_1178,N_1118,N_1113);
or U1179 (N_1179,N_1101,N_1136);
and U1180 (N_1180,N_1147,N_1105);
and U1181 (N_1181,N_1144,N_1123);
and U1182 (N_1182,N_1134,N_1139);
and U1183 (N_1183,N_1116,N_1118);
xnor U1184 (N_1184,N_1135,N_1143);
nand U1185 (N_1185,N_1107,N_1124);
nand U1186 (N_1186,N_1108,N_1131);
nand U1187 (N_1187,N_1106,N_1122);
nor U1188 (N_1188,N_1117,N_1125);
or U1189 (N_1189,N_1110,N_1125);
or U1190 (N_1190,N_1104,N_1124);
nor U1191 (N_1191,N_1142,N_1111);
nor U1192 (N_1192,N_1130,N_1137);
or U1193 (N_1193,N_1145,N_1124);
or U1194 (N_1194,N_1142,N_1136);
nor U1195 (N_1195,N_1127,N_1138);
and U1196 (N_1196,N_1122,N_1139);
or U1197 (N_1197,N_1110,N_1109);
and U1198 (N_1198,N_1134,N_1111);
and U1199 (N_1199,N_1146,N_1101);
nand U1200 (N_1200,N_1165,N_1185);
nand U1201 (N_1201,N_1189,N_1163);
and U1202 (N_1202,N_1179,N_1190);
and U1203 (N_1203,N_1161,N_1157);
nand U1204 (N_1204,N_1177,N_1195);
and U1205 (N_1205,N_1150,N_1158);
nand U1206 (N_1206,N_1172,N_1175);
nand U1207 (N_1207,N_1151,N_1155);
xnor U1208 (N_1208,N_1162,N_1198);
nor U1209 (N_1209,N_1159,N_1170);
nor U1210 (N_1210,N_1178,N_1181);
nand U1211 (N_1211,N_1156,N_1180);
and U1212 (N_1212,N_1199,N_1168);
nor U1213 (N_1213,N_1191,N_1154);
or U1214 (N_1214,N_1152,N_1187);
nor U1215 (N_1215,N_1153,N_1164);
nand U1216 (N_1216,N_1188,N_1171);
and U1217 (N_1217,N_1173,N_1176);
nor U1218 (N_1218,N_1196,N_1194);
xnor U1219 (N_1219,N_1192,N_1169);
or U1220 (N_1220,N_1167,N_1197);
or U1221 (N_1221,N_1186,N_1183);
and U1222 (N_1222,N_1174,N_1184);
or U1223 (N_1223,N_1193,N_1160);
nor U1224 (N_1224,N_1182,N_1166);
or U1225 (N_1225,N_1163,N_1185);
nor U1226 (N_1226,N_1179,N_1183);
nor U1227 (N_1227,N_1156,N_1173);
nor U1228 (N_1228,N_1193,N_1168);
nor U1229 (N_1229,N_1184,N_1162);
or U1230 (N_1230,N_1198,N_1196);
nor U1231 (N_1231,N_1151,N_1193);
or U1232 (N_1232,N_1167,N_1159);
and U1233 (N_1233,N_1151,N_1189);
nand U1234 (N_1234,N_1198,N_1164);
and U1235 (N_1235,N_1167,N_1164);
and U1236 (N_1236,N_1171,N_1153);
nor U1237 (N_1237,N_1171,N_1154);
and U1238 (N_1238,N_1194,N_1195);
or U1239 (N_1239,N_1168,N_1173);
nand U1240 (N_1240,N_1189,N_1193);
or U1241 (N_1241,N_1151,N_1158);
or U1242 (N_1242,N_1189,N_1168);
or U1243 (N_1243,N_1180,N_1172);
nand U1244 (N_1244,N_1176,N_1160);
nand U1245 (N_1245,N_1154,N_1175);
nor U1246 (N_1246,N_1158,N_1178);
and U1247 (N_1247,N_1175,N_1177);
nor U1248 (N_1248,N_1165,N_1154);
nand U1249 (N_1249,N_1161,N_1192);
nor U1250 (N_1250,N_1242,N_1205);
or U1251 (N_1251,N_1220,N_1216);
or U1252 (N_1252,N_1206,N_1209);
nand U1253 (N_1253,N_1226,N_1204);
nand U1254 (N_1254,N_1230,N_1208);
nor U1255 (N_1255,N_1233,N_1238);
and U1256 (N_1256,N_1219,N_1234);
and U1257 (N_1257,N_1229,N_1218);
and U1258 (N_1258,N_1202,N_1246);
and U1259 (N_1259,N_1223,N_1240);
nand U1260 (N_1260,N_1222,N_1213);
and U1261 (N_1261,N_1210,N_1215);
nand U1262 (N_1262,N_1243,N_1247);
nand U1263 (N_1263,N_1224,N_1241);
nor U1264 (N_1264,N_1237,N_1201);
or U1265 (N_1265,N_1244,N_1235);
and U1266 (N_1266,N_1231,N_1232);
nand U1267 (N_1267,N_1212,N_1236);
or U1268 (N_1268,N_1221,N_1245);
and U1269 (N_1269,N_1239,N_1249);
or U1270 (N_1270,N_1207,N_1217);
and U1271 (N_1271,N_1248,N_1214);
and U1272 (N_1272,N_1227,N_1211);
nor U1273 (N_1273,N_1200,N_1225);
or U1274 (N_1274,N_1203,N_1228);
and U1275 (N_1275,N_1212,N_1201);
nor U1276 (N_1276,N_1231,N_1215);
and U1277 (N_1277,N_1213,N_1238);
nor U1278 (N_1278,N_1210,N_1221);
nand U1279 (N_1279,N_1232,N_1216);
nor U1280 (N_1280,N_1200,N_1223);
nand U1281 (N_1281,N_1229,N_1244);
and U1282 (N_1282,N_1232,N_1205);
or U1283 (N_1283,N_1219,N_1232);
and U1284 (N_1284,N_1241,N_1216);
and U1285 (N_1285,N_1201,N_1233);
and U1286 (N_1286,N_1206,N_1228);
nand U1287 (N_1287,N_1234,N_1217);
nor U1288 (N_1288,N_1245,N_1228);
nand U1289 (N_1289,N_1229,N_1208);
or U1290 (N_1290,N_1207,N_1213);
nand U1291 (N_1291,N_1214,N_1218);
nor U1292 (N_1292,N_1210,N_1249);
nor U1293 (N_1293,N_1215,N_1248);
and U1294 (N_1294,N_1201,N_1227);
or U1295 (N_1295,N_1239,N_1201);
nand U1296 (N_1296,N_1206,N_1203);
and U1297 (N_1297,N_1249,N_1235);
and U1298 (N_1298,N_1238,N_1231);
or U1299 (N_1299,N_1217,N_1221);
nor U1300 (N_1300,N_1288,N_1282);
or U1301 (N_1301,N_1258,N_1299);
nand U1302 (N_1302,N_1278,N_1251);
and U1303 (N_1303,N_1287,N_1262);
and U1304 (N_1304,N_1273,N_1265);
and U1305 (N_1305,N_1280,N_1298);
and U1306 (N_1306,N_1290,N_1269);
and U1307 (N_1307,N_1271,N_1296);
nor U1308 (N_1308,N_1266,N_1261);
and U1309 (N_1309,N_1270,N_1257);
or U1310 (N_1310,N_1294,N_1264);
nand U1311 (N_1311,N_1267,N_1250);
or U1312 (N_1312,N_1283,N_1286);
nor U1313 (N_1313,N_1253,N_1279);
xor U1314 (N_1314,N_1291,N_1255);
nand U1315 (N_1315,N_1277,N_1275);
nor U1316 (N_1316,N_1285,N_1252);
nand U1317 (N_1317,N_1289,N_1276);
xnor U1318 (N_1318,N_1274,N_1281);
nand U1319 (N_1319,N_1254,N_1295);
nand U1320 (N_1320,N_1297,N_1293);
nand U1321 (N_1321,N_1268,N_1256);
nor U1322 (N_1322,N_1284,N_1272);
nand U1323 (N_1323,N_1292,N_1260);
and U1324 (N_1324,N_1263,N_1259);
nor U1325 (N_1325,N_1277,N_1252);
nand U1326 (N_1326,N_1288,N_1276);
nand U1327 (N_1327,N_1289,N_1256);
or U1328 (N_1328,N_1277,N_1288);
nor U1329 (N_1329,N_1296,N_1268);
and U1330 (N_1330,N_1285,N_1269);
nor U1331 (N_1331,N_1269,N_1280);
and U1332 (N_1332,N_1251,N_1269);
nor U1333 (N_1333,N_1262,N_1289);
or U1334 (N_1334,N_1285,N_1254);
nand U1335 (N_1335,N_1284,N_1294);
nand U1336 (N_1336,N_1255,N_1271);
nand U1337 (N_1337,N_1280,N_1281);
or U1338 (N_1338,N_1265,N_1290);
or U1339 (N_1339,N_1280,N_1253);
nand U1340 (N_1340,N_1274,N_1288);
or U1341 (N_1341,N_1278,N_1264);
and U1342 (N_1342,N_1294,N_1250);
and U1343 (N_1343,N_1297,N_1288);
nor U1344 (N_1344,N_1256,N_1283);
nor U1345 (N_1345,N_1276,N_1268);
and U1346 (N_1346,N_1273,N_1299);
nor U1347 (N_1347,N_1266,N_1285);
and U1348 (N_1348,N_1281,N_1286);
nor U1349 (N_1349,N_1264,N_1255);
or U1350 (N_1350,N_1311,N_1316);
and U1351 (N_1351,N_1339,N_1313);
or U1352 (N_1352,N_1333,N_1325);
and U1353 (N_1353,N_1321,N_1305);
or U1354 (N_1354,N_1322,N_1349);
nand U1355 (N_1355,N_1301,N_1323);
nor U1356 (N_1356,N_1304,N_1310);
nand U1357 (N_1357,N_1335,N_1308);
or U1358 (N_1358,N_1327,N_1330);
nand U1359 (N_1359,N_1334,N_1328);
nor U1360 (N_1360,N_1338,N_1336);
or U1361 (N_1361,N_1317,N_1331);
or U1362 (N_1362,N_1329,N_1345);
and U1363 (N_1363,N_1318,N_1343);
nand U1364 (N_1364,N_1340,N_1306);
nand U1365 (N_1365,N_1344,N_1346);
or U1366 (N_1366,N_1337,N_1315);
and U1367 (N_1367,N_1309,N_1312);
nor U1368 (N_1368,N_1302,N_1348);
or U1369 (N_1369,N_1342,N_1326);
and U1370 (N_1370,N_1341,N_1300);
and U1371 (N_1371,N_1332,N_1320);
nor U1372 (N_1372,N_1314,N_1347);
nand U1373 (N_1373,N_1307,N_1319);
and U1374 (N_1374,N_1303,N_1324);
or U1375 (N_1375,N_1317,N_1322);
or U1376 (N_1376,N_1322,N_1345);
nand U1377 (N_1377,N_1349,N_1304);
nand U1378 (N_1378,N_1329,N_1338);
and U1379 (N_1379,N_1323,N_1334);
nand U1380 (N_1380,N_1345,N_1310);
nand U1381 (N_1381,N_1332,N_1330);
nand U1382 (N_1382,N_1335,N_1346);
and U1383 (N_1383,N_1323,N_1337);
or U1384 (N_1384,N_1340,N_1314);
and U1385 (N_1385,N_1318,N_1348);
and U1386 (N_1386,N_1323,N_1300);
nor U1387 (N_1387,N_1311,N_1307);
nor U1388 (N_1388,N_1323,N_1333);
or U1389 (N_1389,N_1309,N_1303);
and U1390 (N_1390,N_1332,N_1334);
and U1391 (N_1391,N_1306,N_1339);
and U1392 (N_1392,N_1314,N_1318);
nor U1393 (N_1393,N_1310,N_1320);
or U1394 (N_1394,N_1312,N_1301);
nand U1395 (N_1395,N_1318,N_1320);
or U1396 (N_1396,N_1313,N_1338);
or U1397 (N_1397,N_1339,N_1327);
nand U1398 (N_1398,N_1331,N_1319);
nor U1399 (N_1399,N_1318,N_1344);
nand U1400 (N_1400,N_1360,N_1362);
or U1401 (N_1401,N_1378,N_1361);
xor U1402 (N_1402,N_1376,N_1389);
nand U1403 (N_1403,N_1351,N_1352);
or U1404 (N_1404,N_1384,N_1398);
or U1405 (N_1405,N_1363,N_1366);
nor U1406 (N_1406,N_1355,N_1354);
or U1407 (N_1407,N_1381,N_1383);
or U1408 (N_1408,N_1373,N_1395);
nor U1409 (N_1409,N_1388,N_1394);
or U1410 (N_1410,N_1391,N_1399);
nand U1411 (N_1411,N_1365,N_1374);
and U1412 (N_1412,N_1369,N_1379);
or U1413 (N_1413,N_1359,N_1357);
or U1414 (N_1414,N_1386,N_1350);
nor U1415 (N_1415,N_1387,N_1371);
nor U1416 (N_1416,N_1353,N_1390);
and U1417 (N_1417,N_1358,N_1372);
nand U1418 (N_1418,N_1392,N_1368);
nor U1419 (N_1419,N_1396,N_1367);
or U1420 (N_1420,N_1370,N_1380);
and U1421 (N_1421,N_1364,N_1382);
nor U1422 (N_1422,N_1385,N_1393);
or U1423 (N_1423,N_1375,N_1397);
nor U1424 (N_1424,N_1356,N_1377);
nand U1425 (N_1425,N_1398,N_1366);
or U1426 (N_1426,N_1375,N_1353);
and U1427 (N_1427,N_1394,N_1371);
or U1428 (N_1428,N_1379,N_1399);
nor U1429 (N_1429,N_1390,N_1359);
nand U1430 (N_1430,N_1380,N_1376);
or U1431 (N_1431,N_1377,N_1362);
nand U1432 (N_1432,N_1379,N_1362);
nand U1433 (N_1433,N_1365,N_1353);
nand U1434 (N_1434,N_1358,N_1371);
and U1435 (N_1435,N_1358,N_1370);
nand U1436 (N_1436,N_1376,N_1370);
or U1437 (N_1437,N_1378,N_1367);
nand U1438 (N_1438,N_1373,N_1393);
or U1439 (N_1439,N_1373,N_1387);
nand U1440 (N_1440,N_1359,N_1386);
or U1441 (N_1441,N_1360,N_1369);
and U1442 (N_1442,N_1358,N_1378);
and U1443 (N_1443,N_1379,N_1377);
nor U1444 (N_1444,N_1386,N_1388);
or U1445 (N_1445,N_1365,N_1361);
and U1446 (N_1446,N_1395,N_1365);
nand U1447 (N_1447,N_1378,N_1387);
nand U1448 (N_1448,N_1371,N_1365);
nor U1449 (N_1449,N_1357,N_1398);
or U1450 (N_1450,N_1427,N_1437);
nor U1451 (N_1451,N_1439,N_1402);
or U1452 (N_1452,N_1407,N_1413);
or U1453 (N_1453,N_1418,N_1425);
and U1454 (N_1454,N_1412,N_1438);
nand U1455 (N_1455,N_1429,N_1431);
or U1456 (N_1456,N_1449,N_1415);
nor U1457 (N_1457,N_1433,N_1432);
nand U1458 (N_1458,N_1442,N_1419);
nand U1459 (N_1459,N_1408,N_1424);
and U1460 (N_1460,N_1445,N_1406);
nor U1461 (N_1461,N_1446,N_1400);
and U1462 (N_1462,N_1414,N_1436);
nand U1463 (N_1463,N_1401,N_1420);
and U1464 (N_1464,N_1434,N_1403);
nor U1465 (N_1465,N_1416,N_1443);
nand U1466 (N_1466,N_1409,N_1423);
and U1467 (N_1467,N_1422,N_1440);
nor U1468 (N_1468,N_1405,N_1430);
or U1469 (N_1469,N_1441,N_1404);
or U1470 (N_1470,N_1428,N_1411);
nor U1471 (N_1471,N_1421,N_1417);
or U1472 (N_1472,N_1447,N_1426);
nand U1473 (N_1473,N_1444,N_1435);
or U1474 (N_1474,N_1448,N_1410);
nand U1475 (N_1475,N_1443,N_1401);
nor U1476 (N_1476,N_1407,N_1444);
or U1477 (N_1477,N_1447,N_1430);
nand U1478 (N_1478,N_1412,N_1427);
and U1479 (N_1479,N_1445,N_1436);
nor U1480 (N_1480,N_1431,N_1435);
nand U1481 (N_1481,N_1437,N_1429);
nor U1482 (N_1482,N_1425,N_1400);
nand U1483 (N_1483,N_1403,N_1438);
and U1484 (N_1484,N_1423,N_1445);
or U1485 (N_1485,N_1408,N_1420);
nand U1486 (N_1486,N_1441,N_1448);
or U1487 (N_1487,N_1433,N_1429);
or U1488 (N_1488,N_1435,N_1432);
xor U1489 (N_1489,N_1413,N_1447);
nor U1490 (N_1490,N_1436,N_1428);
or U1491 (N_1491,N_1433,N_1439);
and U1492 (N_1492,N_1413,N_1419);
or U1493 (N_1493,N_1436,N_1409);
or U1494 (N_1494,N_1403,N_1404);
nand U1495 (N_1495,N_1423,N_1403);
nand U1496 (N_1496,N_1443,N_1446);
and U1497 (N_1497,N_1421,N_1445);
nand U1498 (N_1498,N_1407,N_1426);
or U1499 (N_1499,N_1437,N_1449);
nand U1500 (N_1500,N_1484,N_1476);
nor U1501 (N_1501,N_1462,N_1471);
nand U1502 (N_1502,N_1452,N_1490);
and U1503 (N_1503,N_1498,N_1486);
or U1504 (N_1504,N_1497,N_1463);
nor U1505 (N_1505,N_1453,N_1485);
nor U1506 (N_1506,N_1475,N_1460);
or U1507 (N_1507,N_1492,N_1451);
and U1508 (N_1508,N_1470,N_1466);
nand U1509 (N_1509,N_1450,N_1482);
nor U1510 (N_1510,N_1491,N_1456);
nor U1511 (N_1511,N_1457,N_1469);
nand U1512 (N_1512,N_1495,N_1468);
or U1513 (N_1513,N_1483,N_1472);
nand U1514 (N_1514,N_1479,N_1493);
xor U1515 (N_1515,N_1461,N_1494);
nor U1516 (N_1516,N_1478,N_1464);
and U1517 (N_1517,N_1477,N_1474);
nand U1518 (N_1518,N_1458,N_1467);
and U1519 (N_1519,N_1499,N_1496);
nand U1520 (N_1520,N_1459,N_1481);
nand U1521 (N_1521,N_1487,N_1473);
and U1522 (N_1522,N_1480,N_1454);
nor U1523 (N_1523,N_1465,N_1455);
nor U1524 (N_1524,N_1488,N_1489);
and U1525 (N_1525,N_1470,N_1478);
nand U1526 (N_1526,N_1478,N_1469);
or U1527 (N_1527,N_1458,N_1466);
nor U1528 (N_1528,N_1455,N_1495);
nand U1529 (N_1529,N_1452,N_1458);
or U1530 (N_1530,N_1490,N_1451);
nor U1531 (N_1531,N_1478,N_1460);
and U1532 (N_1532,N_1486,N_1464);
nand U1533 (N_1533,N_1470,N_1469);
nand U1534 (N_1534,N_1489,N_1487);
or U1535 (N_1535,N_1453,N_1454);
nor U1536 (N_1536,N_1481,N_1484);
and U1537 (N_1537,N_1452,N_1475);
or U1538 (N_1538,N_1450,N_1498);
and U1539 (N_1539,N_1488,N_1485);
or U1540 (N_1540,N_1473,N_1497);
or U1541 (N_1541,N_1456,N_1455);
nor U1542 (N_1542,N_1457,N_1484);
nor U1543 (N_1543,N_1483,N_1468);
nand U1544 (N_1544,N_1489,N_1478);
and U1545 (N_1545,N_1469,N_1477);
and U1546 (N_1546,N_1473,N_1452);
nand U1547 (N_1547,N_1488,N_1498);
or U1548 (N_1548,N_1486,N_1490);
and U1549 (N_1549,N_1494,N_1475);
nand U1550 (N_1550,N_1546,N_1509);
and U1551 (N_1551,N_1531,N_1525);
nand U1552 (N_1552,N_1512,N_1542);
xor U1553 (N_1553,N_1528,N_1515);
or U1554 (N_1554,N_1527,N_1500);
or U1555 (N_1555,N_1533,N_1510);
nor U1556 (N_1556,N_1540,N_1514);
nor U1557 (N_1557,N_1536,N_1504);
or U1558 (N_1558,N_1549,N_1539);
nand U1559 (N_1559,N_1511,N_1535);
nor U1560 (N_1560,N_1519,N_1543);
nor U1561 (N_1561,N_1530,N_1545);
nor U1562 (N_1562,N_1541,N_1501);
and U1563 (N_1563,N_1505,N_1547);
or U1564 (N_1564,N_1516,N_1517);
nor U1565 (N_1565,N_1534,N_1523);
or U1566 (N_1566,N_1506,N_1513);
nor U1567 (N_1567,N_1529,N_1518);
or U1568 (N_1568,N_1532,N_1507);
nand U1569 (N_1569,N_1537,N_1508);
nor U1570 (N_1570,N_1520,N_1548);
nand U1571 (N_1571,N_1538,N_1502);
or U1572 (N_1572,N_1544,N_1522);
nand U1573 (N_1573,N_1503,N_1524);
nor U1574 (N_1574,N_1521,N_1526);
or U1575 (N_1575,N_1508,N_1529);
nor U1576 (N_1576,N_1519,N_1537);
or U1577 (N_1577,N_1521,N_1549);
and U1578 (N_1578,N_1540,N_1544);
or U1579 (N_1579,N_1505,N_1513);
nand U1580 (N_1580,N_1529,N_1505);
nor U1581 (N_1581,N_1530,N_1540);
nand U1582 (N_1582,N_1501,N_1519);
or U1583 (N_1583,N_1502,N_1517);
or U1584 (N_1584,N_1536,N_1524);
nand U1585 (N_1585,N_1507,N_1533);
nand U1586 (N_1586,N_1511,N_1527);
nor U1587 (N_1587,N_1548,N_1500);
nand U1588 (N_1588,N_1517,N_1533);
or U1589 (N_1589,N_1542,N_1532);
and U1590 (N_1590,N_1522,N_1510);
nand U1591 (N_1591,N_1525,N_1538);
nand U1592 (N_1592,N_1547,N_1549);
and U1593 (N_1593,N_1525,N_1515);
nand U1594 (N_1594,N_1522,N_1507);
and U1595 (N_1595,N_1530,N_1502);
nor U1596 (N_1596,N_1548,N_1541);
nand U1597 (N_1597,N_1500,N_1549);
nand U1598 (N_1598,N_1549,N_1538);
nor U1599 (N_1599,N_1526,N_1533);
nand U1600 (N_1600,N_1581,N_1572);
or U1601 (N_1601,N_1562,N_1568);
and U1602 (N_1602,N_1573,N_1576);
nand U1603 (N_1603,N_1586,N_1585);
nand U1604 (N_1604,N_1558,N_1593);
nor U1605 (N_1605,N_1587,N_1599);
nand U1606 (N_1606,N_1574,N_1580);
or U1607 (N_1607,N_1566,N_1596);
nand U1608 (N_1608,N_1592,N_1570);
nand U1609 (N_1609,N_1567,N_1565);
nand U1610 (N_1610,N_1561,N_1550);
or U1611 (N_1611,N_1591,N_1582);
nand U1612 (N_1612,N_1575,N_1589);
nand U1613 (N_1613,N_1554,N_1557);
or U1614 (N_1614,N_1598,N_1569);
nand U1615 (N_1615,N_1577,N_1579);
nand U1616 (N_1616,N_1551,N_1556);
nor U1617 (N_1617,N_1559,N_1563);
and U1618 (N_1618,N_1584,N_1552);
or U1619 (N_1619,N_1555,N_1564);
or U1620 (N_1620,N_1597,N_1553);
or U1621 (N_1621,N_1595,N_1571);
nor U1622 (N_1622,N_1578,N_1588);
and U1623 (N_1623,N_1594,N_1560);
or U1624 (N_1624,N_1590,N_1583);
or U1625 (N_1625,N_1564,N_1582);
or U1626 (N_1626,N_1556,N_1596);
or U1627 (N_1627,N_1588,N_1556);
or U1628 (N_1628,N_1566,N_1568);
and U1629 (N_1629,N_1567,N_1559);
or U1630 (N_1630,N_1550,N_1583);
or U1631 (N_1631,N_1552,N_1575);
nand U1632 (N_1632,N_1591,N_1574);
nand U1633 (N_1633,N_1581,N_1592);
and U1634 (N_1634,N_1567,N_1556);
nor U1635 (N_1635,N_1583,N_1598);
and U1636 (N_1636,N_1597,N_1556);
nand U1637 (N_1637,N_1552,N_1586);
or U1638 (N_1638,N_1590,N_1552);
or U1639 (N_1639,N_1555,N_1578);
nor U1640 (N_1640,N_1570,N_1583);
nor U1641 (N_1641,N_1564,N_1571);
or U1642 (N_1642,N_1589,N_1591);
or U1643 (N_1643,N_1560,N_1590);
and U1644 (N_1644,N_1574,N_1592);
nand U1645 (N_1645,N_1570,N_1559);
nor U1646 (N_1646,N_1568,N_1575);
or U1647 (N_1647,N_1585,N_1572);
or U1648 (N_1648,N_1557,N_1562);
or U1649 (N_1649,N_1597,N_1562);
and U1650 (N_1650,N_1639,N_1630);
nor U1651 (N_1651,N_1644,N_1608);
nand U1652 (N_1652,N_1610,N_1648);
or U1653 (N_1653,N_1634,N_1619);
nand U1654 (N_1654,N_1628,N_1645);
nor U1655 (N_1655,N_1600,N_1614);
and U1656 (N_1656,N_1641,N_1635);
and U1657 (N_1657,N_1642,N_1637);
nor U1658 (N_1658,N_1612,N_1621);
nand U1659 (N_1659,N_1631,N_1616);
or U1660 (N_1660,N_1605,N_1606);
nor U1661 (N_1661,N_1649,N_1601);
and U1662 (N_1662,N_1627,N_1646);
or U1663 (N_1663,N_1633,N_1611);
or U1664 (N_1664,N_1602,N_1622);
and U1665 (N_1665,N_1624,N_1638);
nor U1666 (N_1666,N_1603,N_1618);
nand U1667 (N_1667,N_1623,N_1615);
and U1668 (N_1668,N_1607,N_1643);
or U1669 (N_1669,N_1629,N_1640);
nor U1670 (N_1670,N_1609,N_1636);
or U1671 (N_1671,N_1613,N_1626);
or U1672 (N_1672,N_1632,N_1625);
and U1673 (N_1673,N_1647,N_1617);
or U1674 (N_1674,N_1620,N_1604);
nor U1675 (N_1675,N_1616,N_1645);
nand U1676 (N_1676,N_1600,N_1613);
and U1677 (N_1677,N_1619,N_1616);
and U1678 (N_1678,N_1627,N_1622);
or U1679 (N_1679,N_1631,N_1637);
nand U1680 (N_1680,N_1614,N_1639);
or U1681 (N_1681,N_1609,N_1604);
nor U1682 (N_1682,N_1619,N_1641);
and U1683 (N_1683,N_1631,N_1630);
nor U1684 (N_1684,N_1640,N_1646);
and U1685 (N_1685,N_1608,N_1607);
nand U1686 (N_1686,N_1635,N_1609);
nand U1687 (N_1687,N_1616,N_1643);
nand U1688 (N_1688,N_1610,N_1632);
or U1689 (N_1689,N_1637,N_1633);
and U1690 (N_1690,N_1616,N_1640);
and U1691 (N_1691,N_1630,N_1637);
or U1692 (N_1692,N_1603,N_1601);
and U1693 (N_1693,N_1649,N_1644);
and U1694 (N_1694,N_1601,N_1647);
nand U1695 (N_1695,N_1648,N_1613);
nand U1696 (N_1696,N_1625,N_1601);
and U1697 (N_1697,N_1639,N_1610);
or U1698 (N_1698,N_1606,N_1615);
nand U1699 (N_1699,N_1621,N_1616);
nor U1700 (N_1700,N_1675,N_1652);
or U1701 (N_1701,N_1683,N_1684);
or U1702 (N_1702,N_1687,N_1662);
nor U1703 (N_1703,N_1661,N_1678);
and U1704 (N_1704,N_1668,N_1672);
and U1705 (N_1705,N_1688,N_1660);
nor U1706 (N_1706,N_1663,N_1671);
nor U1707 (N_1707,N_1682,N_1673);
nor U1708 (N_1708,N_1679,N_1653);
nor U1709 (N_1709,N_1697,N_1681);
or U1710 (N_1710,N_1696,N_1693);
nor U1711 (N_1711,N_1674,N_1689);
and U1712 (N_1712,N_1664,N_1698);
or U1713 (N_1713,N_1695,N_1670);
and U1714 (N_1714,N_1665,N_1676);
nor U1715 (N_1715,N_1667,N_1659);
nor U1716 (N_1716,N_1654,N_1690);
or U1717 (N_1717,N_1699,N_1657);
or U1718 (N_1718,N_1651,N_1658);
or U1719 (N_1719,N_1650,N_1692);
and U1720 (N_1720,N_1656,N_1666);
nand U1721 (N_1721,N_1685,N_1686);
and U1722 (N_1722,N_1669,N_1680);
nand U1723 (N_1723,N_1691,N_1694);
nand U1724 (N_1724,N_1677,N_1655);
nor U1725 (N_1725,N_1661,N_1686);
xor U1726 (N_1726,N_1660,N_1659);
nand U1727 (N_1727,N_1664,N_1691);
nor U1728 (N_1728,N_1673,N_1694);
and U1729 (N_1729,N_1665,N_1658);
or U1730 (N_1730,N_1652,N_1673);
nor U1731 (N_1731,N_1659,N_1668);
nor U1732 (N_1732,N_1699,N_1661);
and U1733 (N_1733,N_1663,N_1674);
and U1734 (N_1734,N_1657,N_1659);
nand U1735 (N_1735,N_1663,N_1669);
and U1736 (N_1736,N_1659,N_1671);
or U1737 (N_1737,N_1683,N_1657);
or U1738 (N_1738,N_1698,N_1675);
and U1739 (N_1739,N_1695,N_1697);
nand U1740 (N_1740,N_1656,N_1680);
or U1741 (N_1741,N_1684,N_1659);
and U1742 (N_1742,N_1656,N_1689);
and U1743 (N_1743,N_1668,N_1690);
and U1744 (N_1744,N_1673,N_1693);
or U1745 (N_1745,N_1674,N_1650);
nand U1746 (N_1746,N_1679,N_1664);
nand U1747 (N_1747,N_1672,N_1676);
or U1748 (N_1748,N_1689,N_1680);
and U1749 (N_1749,N_1660,N_1662);
or U1750 (N_1750,N_1731,N_1718);
nand U1751 (N_1751,N_1706,N_1700);
nor U1752 (N_1752,N_1743,N_1704);
nor U1753 (N_1753,N_1702,N_1709);
and U1754 (N_1754,N_1708,N_1723);
nand U1755 (N_1755,N_1736,N_1712);
and U1756 (N_1756,N_1714,N_1710);
and U1757 (N_1757,N_1746,N_1705);
nand U1758 (N_1758,N_1703,N_1720);
or U1759 (N_1759,N_1707,N_1716);
nor U1760 (N_1760,N_1726,N_1739);
nand U1761 (N_1761,N_1715,N_1722);
nor U1762 (N_1762,N_1744,N_1734);
nand U1763 (N_1763,N_1711,N_1738);
nor U1764 (N_1764,N_1724,N_1737);
and U1765 (N_1765,N_1729,N_1728);
and U1766 (N_1766,N_1733,N_1725);
or U1767 (N_1767,N_1717,N_1727);
and U1768 (N_1768,N_1741,N_1732);
or U1769 (N_1769,N_1747,N_1701);
nor U1770 (N_1770,N_1735,N_1740);
nor U1771 (N_1771,N_1719,N_1748);
and U1772 (N_1772,N_1730,N_1749);
nor U1773 (N_1773,N_1745,N_1742);
nor U1774 (N_1774,N_1713,N_1721);
nand U1775 (N_1775,N_1747,N_1704);
nand U1776 (N_1776,N_1701,N_1705);
or U1777 (N_1777,N_1715,N_1704);
nor U1778 (N_1778,N_1704,N_1731);
nand U1779 (N_1779,N_1717,N_1749);
and U1780 (N_1780,N_1738,N_1712);
or U1781 (N_1781,N_1726,N_1723);
nor U1782 (N_1782,N_1747,N_1727);
xor U1783 (N_1783,N_1702,N_1714);
and U1784 (N_1784,N_1705,N_1713);
and U1785 (N_1785,N_1745,N_1707);
and U1786 (N_1786,N_1728,N_1702);
or U1787 (N_1787,N_1727,N_1719);
or U1788 (N_1788,N_1711,N_1736);
nor U1789 (N_1789,N_1702,N_1721);
or U1790 (N_1790,N_1739,N_1704);
or U1791 (N_1791,N_1733,N_1740);
and U1792 (N_1792,N_1745,N_1709);
and U1793 (N_1793,N_1748,N_1725);
nand U1794 (N_1794,N_1725,N_1742);
nor U1795 (N_1795,N_1711,N_1709);
nand U1796 (N_1796,N_1730,N_1741);
and U1797 (N_1797,N_1715,N_1733);
nand U1798 (N_1798,N_1746,N_1704);
nor U1799 (N_1799,N_1732,N_1734);
nor U1800 (N_1800,N_1781,N_1766);
or U1801 (N_1801,N_1793,N_1784);
and U1802 (N_1802,N_1767,N_1770);
and U1803 (N_1803,N_1768,N_1794);
nand U1804 (N_1804,N_1755,N_1772);
nand U1805 (N_1805,N_1752,N_1762);
nand U1806 (N_1806,N_1751,N_1789);
nor U1807 (N_1807,N_1795,N_1750);
or U1808 (N_1808,N_1760,N_1754);
nor U1809 (N_1809,N_1765,N_1771);
nand U1810 (N_1810,N_1796,N_1764);
nand U1811 (N_1811,N_1792,N_1758);
nor U1812 (N_1812,N_1763,N_1790);
and U1813 (N_1813,N_1782,N_1774);
nand U1814 (N_1814,N_1775,N_1753);
or U1815 (N_1815,N_1778,N_1779);
and U1816 (N_1816,N_1785,N_1786);
nand U1817 (N_1817,N_1761,N_1799);
and U1818 (N_1818,N_1756,N_1798);
or U1819 (N_1819,N_1769,N_1776);
nand U1820 (N_1820,N_1791,N_1788);
or U1821 (N_1821,N_1787,N_1773);
and U1822 (N_1822,N_1780,N_1783);
and U1823 (N_1823,N_1797,N_1777);
or U1824 (N_1824,N_1757,N_1759);
or U1825 (N_1825,N_1753,N_1787);
or U1826 (N_1826,N_1776,N_1792);
nor U1827 (N_1827,N_1784,N_1799);
and U1828 (N_1828,N_1753,N_1772);
and U1829 (N_1829,N_1781,N_1786);
or U1830 (N_1830,N_1753,N_1762);
or U1831 (N_1831,N_1776,N_1777);
nor U1832 (N_1832,N_1767,N_1774);
nor U1833 (N_1833,N_1791,N_1779);
and U1834 (N_1834,N_1769,N_1786);
and U1835 (N_1835,N_1756,N_1759);
and U1836 (N_1836,N_1789,N_1756);
and U1837 (N_1837,N_1772,N_1756);
nor U1838 (N_1838,N_1791,N_1777);
and U1839 (N_1839,N_1792,N_1779);
nand U1840 (N_1840,N_1778,N_1774);
nand U1841 (N_1841,N_1796,N_1756);
and U1842 (N_1842,N_1751,N_1757);
nor U1843 (N_1843,N_1790,N_1775);
nor U1844 (N_1844,N_1767,N_1772);
nor U1845 (N_1845,N_1775,N_1791);
nor U1846 (N_1846,N_1788,N_1798);
nand U1847 (N_1847,N_1769,N_1795);
nand U1848 (N_1848,N_1795,N_1781);
and U1849 (N_1849,N_1780,N_1759);
nand U1850 (N_1850,N_1839,N_1847);
nor U1851 (N_1851,N_1841,N_1833);
and U1852 (N_1852,N_1810,N_1820);
nor U1853 (N_1853,N_1819,N_1835);
nor U1854 (N_1854,N_1823,N_1843);
or U1855 (N_1855,N_1824,N_1836);
or U1856 (N_1856,N_1821,N_1844);
nand U1857 (N_1857,N_1825,N_1804);
nand U1858 (N_1858,N_1818,N_1827);
nor U1859 (N_1859,N_1826,N_1848);
or U1860 (N_1860,N_1815,N_1840);
nor U1861 (N_1861,N_1802,N_1800);
nand U1862 (N_1862,N_1814,N_1816);
nand U1863 (N_1863,N_1849,N_1830);
and U1864 (N_1864,N_1811,N_1837);
nand U1865 (N_1865,N_1801,N_1813);
nand U1866 (N_1866,N_1838,N_1807);
and U1867 (N_1867,N_1845,N_1806);
and U1868 (N_1868,N_1809,N_1846);
and U1869 (N_1869,N_1822,N_1812);
and U1870 (N_1870,N_1834,N_1831);
nand U1871 (N_1871,N_1803,N_1805);
and U1872 (N_1872,N_1832,N_1829);
or U1873 (N_1873,N_1817,N_1808);
nor U1874 (N_1874,N_1842,N_1828);
or U1875 (N_1875,N_1828,N_1824);
nand U1876 (N_1876,N_1845,N_1819);
nor U1877 (N_1877,N_1800,N_1839);
nor U1878 (N_1878,N_1839,N_1803);
nand U1879 (N_1879,N_1803,N_1828);
and U1880 (N_1880,N_1844,N_1818);
nand U1881 (N_1881,N_1805,N_1813);
and U1882 (N_1882,N_1811,N_1843);
nand U1883 (N_1883,N_1826,N_1822);
and U1884 (N_1884,N_1805,N_1807);
or U1885 (N_1885,N_1839,N_1808);
nor U1886 (N_1886,N_1829,N_1809);
nor U1887 (N_1887,N_1828,N_1825);
and U1888 (N_1888,N_1819,N_1836);
and U1889 (N_1889,N_1803,N_1810);
nor U1890 (N_1890,N_1828,N_1806);
or U1891 (N_1891,N_1818,N_1835);
nor U1892 (N_1892,N_1844,N_1825);
or U1893 (N_1893,N_1800,N_1822);
or U1894 (N_1894,N_1808,N_1830);
nand U1895 (N_1895,N_1812,N_1826);
and U1896 (N_1896,N_1819,N_1815);
and U1897 (N_1897,N_1842,N_1821);
or U1898 (N_1898,N_1835,N_1846);
or U1899 (N_1899,N_1814,N_1846);
nand U1900 (N_1900,N_1852,N_1854);
nand U1901 (N_1901,N_1896,N_1882);
or U1902 (N_1902,N_1862,N_1880);
and U1903 (N_1903,N_1895,N_1897);
or U1904 (N_1904,N_1879,N_1868);
and U1905 (N_1905,N_1884,N_1885);
nand U1906 (N_1906,N_1876,N_1898);
nor U1907 (N_1907,N_1891,N_1865);
or U1908 (N_1908,N_1887,N_1893);
nor U1909 (N_1909,N_1875,N_1871);
and U1910 (N_1910,N_1873,N_1899);
or U1911 (N_1911,N_1851,N_1853);
and U1912 (N_1912,N_1881,N_1883);
nand U1913 (N_1913,N_1861,N_1850);
nand U1914 (N_1914,N_1860,N_1892);
and U1915 (N_1915,N_1872,N_1855);
or U1916 (N_1916,N_1874,N_1878);
nor U1917 (N_1917,N_1857,N_1889);
nor U1918 (N_1918,N_1863,N_1894);
nand U1919 (N_1919,N_1866,N_1859);
or U1920 (N_1920,N_1890,N_1886);
and U1921 (N_1921,N_1877,N_1856);
or U1922 (N_1922,N_1888,N_1858);
nor U1923 (N_1923,N_1864,N_1869);
or U1924 (N_1924,N_1867,N_1870);
nor U1925 (N_1925,N_1868,N_1891);
nor U1926 (N_1926,N_1876,N_1851);
nor U1927 (N_1927,N_1850,N_1858);
nor U1928 (N_1928,N_1870,N_1871);
nand U1929 (N_1929,N_1885,N_1867);
nor U1930 (N_1930,N_1877,N_1875);
nand U1931 (N_1931,N_1870,N_1878);
nor U1932 (N_1932,N_1861,N_1897);
and U1933 (N_1933,N_1877,N_1854);
nor U1934 (N_1934,N_1873,N_1876);
and U1935 (N_1935,N_1893,N_1889);
nand U1936 (N_1936,N_1872,N_1868);
nor U1937 (N_1937,N_1878,N_1850);
or U1938 (N_1938,N_1870,N_1898);
nor U1939 (N_1939,N_1883,N_1859);
xnor U1940 (N_1940,N_1871,N_1886);
nor U1941 (N_1941,N_1861,N_1894);
and U1942 (N_1942,N_1878,N_1851);
or U1943 (N_1943,N_1858,N_1853);
nand U1944 (N_1944,N_1891,N_1874);
nand U1945 (N_1945,N_1870,N_1862);
or U1946 (N_1946,N_1881,N_1850);
and U1947 (N_1947,N_1870,N_1874);
nor U1948 (N_1948,N_1888,N_1885);
nand U1949 (N_1949,N_1876,N_1857);
nand U1950 (N_1950,N_1921,N_1902);
or U1951 (N_1951,N_1926,N_1903);
nand U1952 (N_1952,N_1909,N_1949);
or U1953 (N_1953,N_1927,N_1932);
nand U1954 (N_1954,N_1904,N_1924);
or U1955 (N_1955,N_1944,N_1910);
nand U1956 (N_1956,N_1933,N_1907);
or U1957 (N_1957,N_1919,N_1928);
nand U1958 (N_1958,N_1915,N_1935);
nor U1959 (N_1959,N_1941,N_1934);
nand U1960 (N_1960,N_1943,N_1937);
nor U1961 (N_1961,N_1947,N_1930);
nand U1962 (N_1962,N_1905,N_1906);
or U1963 (N_1963,N_1946,N_1918);
or U1964 (N_1964,N_1916,N_1939);
nand U1965 (N_1965,N_1908,N_1917);
or U1966 (N_1966,N_1911,N_1900);
nor U1967 (N_1967,N_1936,N_1901);
nand U1968 (N_1968,N_1925,N_1923);
or U1969 (N_1969,N_1938,N_1922);
and U1970 (N_1970,N_1912,N_1945);
nand U1971 (N_1971,N_1940,N_1929);
and U1972 (N_1972,N_1914,N_1948);
nand U1973 (N_1973,N_1931,N_1942);
nor U1974 (N_1974,N_1920,N_1913);
and U1975 (N_1975,N_1941,N_1920);
nor U1976 (N_1976,N_1913,N_1935);
and U1977 (N_1977,N_1928,N_1929);
nand U1978 (N_1978,N_1925,N_1930);
and U1979 (N_1979,N_1948,N_1906);
nor U1980 (N_1980,N_1905,N_1926);
or U1981 (N_1981,N_1946,N_1940);
or U1982 (N_1982,N_1910,N_1938);
nand U1983 (N_1983,N_1943,N_1907);
or U1984 (N_1984,N_1944,N_1931);
or U1985 (N_1985,N_1905,N_1901);
nand U1986 (N_1986,N_1905,N_1945);
nor U1987 (N_1987,N_1901,N_1919);
or U1988 (N_1988,N_1901,N_1930);
nand U1989 (N_1989,N_1901,N_1926);
nand U1990 (N_1990,N_1901,N_1920);
or U1991 (N_1991,N_1942,N_1933);
and U1992 (N_1992,N_1935,N_1941);
and U1993 (N_1993,N_1944,N_1948);
nand U1994 (N_1994,N_1931,N_1940);
or U1995 (N_1995,N_1922,N_1919);
nand U1996 (N_1996,N_1919,N_1904);
nor U1997 (N_1997,N_1928,N_1945);
nand U1998 (N_1998,N_1934,N_1940);
and U1999 (N_1999,N_1937,N_1944);
nor U2000 (N_2000,N_1953,N_1998);
and U2001 (N_2001,N_1962,N_1972);
or U2002 (N_2002,N_1952,N_1993);
nor U2003 (N_2003,N_1987,N_1967);
and U2004 (N_2004,N_1985,N_1988);
and U2005 (N_2005,N_1996,N_1963);
and U2006 (N_2006,N_1980,N_1991);
and U2007 (N_2007,N_1951,N_1982);
nand U2008 (N_2008,N_1956,N_1955);
nand U2009 (N_2009,N_1957,N_1970);
or U2010 (N_2010,N_1994,N_1999);
or U2011 (N_2011,N_1986,N_1997);
and U2012 (N_2012,N_1974,N_1969);
nor U2013 (N_2013,N_1954,N_1965);
nand U2014 (N_2014,N_1971,N_1976);
or U2015 (N_2015,N_1990,N_1978);
nor U2016 (N_2016,N_1966,N_1959);
or U2017 (N_2017,N_1964,N_1975);
nor U2018 (N_2018,N_1950,N_1960);
or U2019 (N_2019,N_1958,N_1981);
nor U2020 (N_2020,N_1992,N_1961);
nand U2021 (N_2021,N_1995,N_1977);
and U2022 (N_2022,N_1968,N_1984);
nand U2023 (N_2023,N_1973,N_1989);
and U2024 (N_2024,N_1979,N_1983);
nor U2025 (N_2025,N_1971,N_1972);
nand U2026 (N_2026,N_1976,N_1982);
and U2027 (N_2027,N_1963,N_1998);
and U2028 (N_2028,N_1993,N_1960);
nand U2029 (N_2029,N_1981,N_1966);
and U2030 (N_2030,N_1991,N_1984);
and U2031 (N_2031,N_1995,N_1980);
or U2032 (N_2032,N_1951,N_1972);
nand U2033 (N_2033,N_1976,N_1994);
nor U2034 (N_2034,N_1954,N_1990);
or U2035 (N_2035,N_1994,N_1967);
or U2036 (N_2036,N_1954,N_1963);
nor U2037 (N_2037,N_1962,N_1986);
and U2038 (N_2038,N_1951,N_1955);
nor U2039 (N_2039,N_1952,N_1998);
or U2040 (N_2040,N_1993,N_1969);
nor U2041 (N_2041,N_1969,N_1962);
and U2042 (N_2042,N_1986,N_1958);
and U2043 (N_2043,N_1989,N_1999);
and U2044 (N_2044,N_1959,N_1960);
and U2045 (N_2045,N_1969,N_1990);
or U2046 (N_2046,N_1958,N_1972);
and U2047 (N_2047,N_1975,N_1997);
nor U2048 (N_2048,N_1983,N_1997);
nor U2049 (N_2049,N_1958,N_1989);
nand U2050 (N_2050,N_2009,N_2036);
nand U2051 (N_2051,N_2010,N_2006);
and U2052 (N_2052,N_2021,N_2028);
nand U2053 (N_2053,N_2044,N_2038);
and U2054 (N_2054,N_2004,N_2035);
or U2055 (N_2055,N_2029,N_2048);
nor U2056 (N_2056,N_2005,N_2003);
or U2057 (N_2057,N_2008,N_2014);
and U2058 (N_2058,N_2027,N_2011);
and U2059 (N_2059,N_2030,N_2034);
and U2060 (N_2060,N_2041,N_2017);
nand U2061 (N_2061,N_2007,N_2001);
nor U2062 (N_2062,N_2023,N_2016);
or U2063 (N_2063,N_2026,N_2049);
nand U2064 (N_2064,N_2046,N_2033);
or U2065 (N_2065,N_2039,N_2045);
nand U2066 (N_2066,N_2018,N_2000);
and U2067 (N_2067,N_2032,N_2002);
and U2068 (N_2068,N_2047,N_2043);
nor U2069 (N_2069,N_2019,N_2015);
or U2070 (N_2070,N_2040,N_2025);
and U2071 (N_2071,N_2020,N_2042);
and U2072 (N_2072,N_2022,N_2037);
nor U2073 (N_2073,N_2012,N_2013);
nand U2074 (N_2074,N_2031,N_2024);
nor U2075 (N_2075,N_2041,N_2046);
or U2076 (N_2076,N_2008,N_2021);
and U2077 (N_2077,N_2039,N_2032);
nand U2078 (N_2078,N_2019,N_2036);
nor U2079 (N_2079,N_2044,N_2036);
or U2080 (N_2080,N_2016,N_2036);
nor U2081 (N_2081,N_2027,N_2029);
or U2082 (N_2082,N_2028,N_2033);
or U2083 (N_2083,N_2025,N_2007);
nor U2084 (N_2084,N_2038,N_2010);
nor U2085 (N_2085,N_2002,N_2008);
nand U2086 (N_2086,N_2041,N_2039);
or U2087 (N_2087,N_2017,N_2039);
nand U2088 (N_2088,N_2039,N_2026);
nor U2089 (N_2089,N_2011,N_2013);
nand U2090 (N_2090,N_2008,N_2022);
or U2091 (N_2091,N_2024,N_2044);
and U2092 (N_2092,N_2001,N_2048);
or U2093 (N_2093,N_2015,N_2039);
nor U2094 (N_2094,N_2042,N_2002);
nor U2095 (N_2095,N_2003,N_2016);
nand U2096 (N_2096,N_2038,N_2013);
nor U2097 (N_2097,N_2009,N_2021);
and U2098 (N_2098,N_2048,N_2008);
or U2099 (N_2099,N_2001,N_2035);
nor U2100 (N_2100,N_2073,N_2052);
and U2101 (N_2101,N_2096,N_2054);
nor U2102 (N_2102,N_2084,N_2056);
and U2103 (N_2103,N_2093,N_2079);
nand U2104 (N_2104,N_2088,N_2072);
nor U2105 (N_2105,N_2083,N_2095);
or U2106 (N_2106,N_2076,N_2075);
and U2107 (N_2107,N_2092,N_2067);
xnor U2108 (N_2108,N_2078,N_2094);
or U2109 (N_2109,N_2050,N_2066);
and U2110 (N_2110,N_2065,N_2081);
nor U2111 (N_2111,N_2085,N_2090);
and U2112 (N_2112,N_2069,N_2068);
and U2113 (N_2113,N_2098,N_2059);
and U2114 (N_2114,N_2070,N_2086);
and U2115 (N_2115,N_2080,N_2053);
or U2116 (N_2116,N_2057,N_2060);
or U2117 (N_2117,N_2082,N_2071);
and U2118 (N_2118,N_2089,N_2087);
nor U2119 (N_2119,N_2097,N_2099);
and U2120 (N_2120,N_2077,N_2062);
and U2121 (N_2121,N_2091,N_2074);
or U2122 (N_2122,N_2061,N_2051);
or U2123 (N_2123,N_2063,N_2058);
or U2124 (N_2124,N_2064,N_2055);
and U2125 (N_2125,N_2066,N_2077);
nand U2126 (N_2126,N_2065,N_2058);
nor U2127 (N_2127,N_2082,N_2079);
or U2128 (N_2128,N_2060,N_2098);
nor U2129 (N_2129,N_2059,N_2052);
or U2130 (N_2130,N_2090,N_2094);
or U2131 (N_2131,N_2060,N_2076);
and U2132 (N_2132,N_2089,N_2084);
nor U2133 (N_2133,N_2051,N_2093);
and U2134 (N_2134,N_2078,N_2067);
or U2135 (N_2135,N_2077,N_2065);
nor U2136 (N_2136,N_2089,N_2076);
and U2137 (N_2137,N_2056,N_2077);
nand U2138 (N_2138,N_2083,N_2068);
nand U2139 (N_2139,N_2052,N_2089);
and U2140 (N_2140,N_2083,N_2050);
and U2141 (N_2141,N_2075,N_2083);
nor U2142 (N_2142,N_2089,N_2099);
nor U2143 (N_2143,N_2086,N_2075);
nand U2144 (N_2144,N_2062,N_2088);
nand U2145 (N_2145,N_2084,N_2082);
and U2146 (N_2146,N_2072,N_2056);
and U2147 (N_2147,N_2060,N_2052);
nor U2148 (N_2148,N_2099,N_2096);
and U2149 (N_2149,N_2064,N_2074);
or U2150 (N_2150,N_2116,N_2105);
or U2151 (N_2151,N_2128,N_2149);
nand U2152 (N_2152,N_2125,N_2123);
nor U2153 (N_2153,N_2118,N_2108);
or U2154 (N_2154,N_2111,N_2135);
nor U2155 (N_2155,N_2109,N_2112);
or U2156 (N_2156,N_2148,N_2138);
nor U2157 (N_2157,N_2121,N_2106);
nand U2158 (N_2158,N_2114,N_2131);
or U2159 (N_2159,N_2113,N_2142);
and U2160 (N_2160,N_2101,N_2102);
nand U2161 (N_2161,N_2139,N_2129);
nand U2162 (N_2162,N_2133,N_2134);
xor U2163 (N_2163,N_2126,N_2127);
xor U2164 (N_2164,N_2145,N_2140);
or U2165 (N_2165,N_2146,N_2104);
or U2166 (N_2166,N_2119,N_2130);
and U2167 (N_2167,N_2132,N_2143);
nor U2168 (N_2168,N_2136,N_2117);
or U2169 (N_2169,N_2100,N_2107);
and U2170 (N_2170,N_2147,N_2122);
or U2171 (N_2171,N_2120,N_2144);
and U2172 (N_2172,N_2141,N_2110);
and U2173 (N_2173,N_2124,N_2115);
and U2174 (N_2174,N_2103,N_2137);
nand U2175 (N_2175,N_2111,N_2138);
nor U2176 (N_2176,N_2135,N_2118);
or U2177 (N_2177,N_2120,N_2147);
and U2178 (N_2178,N_2133,N_2132);
and U2179 (N_2179,N_2105,N_2114);
nor U2180 (N_2180,N_2108,N_2111);
nand U2181 (N_2181,N_2109,N_2148);
nor U2182 (N_2182,N_2111,N_2140);
nand U2183 (N_2183,N_2102,N_2136);
nand U2184 (N_2184,N_2131,N_2121);
nor U2185 (N_2185,N_2135,N_2143);
nand U2186 (N_2186,N_2130,N_2123);
nor U2187 (N_2187,N_2143,N_2141);
nand U2188 (N_2188,N_2144,N_2115);
nor U2189 (N_2189,N_2104,N_2130);
or U2190 (N_2190,N_2109,N_2137);
or U2191 (N_2191,N_2127,N_2144);
nand U2192 (N_2192,N_2113,N_2143);
or U2193 (N_2193,N_2122,N_2144);
nand U2194 (N_2194,N_2112,N_2146);
and U2195 (N_2195,N_2116,N_2125);
nor U2196 (N_2196,N_2110,N_2111);
nor U2197 (N_2197,N_2142,N_2137);
nor U2198 (N_2198,N_2102,N_2119);
and U2199 (N_2199,N_2119,N_2120);
or U2200 (N_2200,N_2198,N_2167);
nor U2201 (N_2201,N_2197,N_2175);
or U2202 (N_2202,N_2199,N_2181);
nor U2203 (N_2203,N_2150,N_2183);
nor U2204 (N_2204,N_2180,N_2170);
nor U2205 (N_2205,N_2195,N_2156);
or U2206 (N_2206,N_2162,N_2164);
nand U2207 (N_2207,N_2159,N_2182);
or U2208 (N_2208,N_2165,N_2186);
nor U2209 (N_2209,N_2155,N_2174);
or U2210 (N_2210,N_2158,N_2187);
and U2211 (N_2211,N_2185,N_2191);
nand U2212 (N_2212,N_2184,N_2193);
and U2213 (N_2213,N_2196,N_2153);
and U2214 (N_2214,N_2179,N_2177);
or U2215 (N_2215,N_2189,N_2192);
or U2216 (N_2216,N_2188,N_2173);
nand U2217 (N_2217,N_2151,N_2157);
and U2218 (N_2218,N_2178,N_2171);
nor U2219 (N_2219,N_2168,N_2169);
and U2220 (N_2220,N_2194,N_2152);
nor U2221 (N_2221,N_2190,N_2176);
xnor U2222 (N_2222,N_2161,N_2172);
or U2223 (N_2223,N_2163,N_2154);
nand U2224 (N_2224,N_2166,N_2160);
nor U2225 (N_2225,N_2177,N_2181);
or U2226 (N_2226,N_2193,N_2180);
nand U2227 (N_2227,N_2178,N_2162);
or U2228 (N_2228,N_2190,N_2158);
and U2229 (N_2229,N_2195,N_2162);
nand U2230 (N_2230,N_2174,N_2156);
or U2231 (N_2231,N_2164,N_2199);
and U2232 (N_2232,N_2179,N_2185);
nor U2233 (N_2233,N_2167,N_2183);
nand U2234 (N_2234,N_2154,N_2150);
and U2235 (N_2235,N_2175,N_2161);
nand U2236 (N_2236,N_2196,N_2157);
nand U2237 (N_2237,N_2188,N_2197);
or U2238 (N_2238,N_2158,N_2162);
nor U2239 (N_2239,N_2170,N_2175);
nand U2240 (N_2240,N_2183,N_2161);
and U2241 (N_2241,N_2183,N_2199);
or U2242 (N_2242,N_2175,N_2182);
nor U2243 (N_2243,N_2189,N_2174);
and U2244 (N_2244,N_2170,N_2167);
nand U2245 (N_2245,N_2185,N_2156);
and U2246 (N_2246,N_2164,N_2194);
or U2247 (N_2247,N_2183,N_2158);
and U2248 (N_2248,N_2150,N_2192);
nand U2249 (N_2249,N_2169,N_2181);
nor U2250 (N_2250,N_2211,N_2245);
nor U2251 (N_2251,N_2229,N_2203);
nand U2252 (N_2252,N_2212,N_2226);
and U2253 (N_2253,N_2215,N_2243);
nand U2254 (N_2254,N_2224,N_2221);
or U2255 (N_2255,N_2209,N_2202);
or U2256 (N_2256,N_2210,N_2208);
nand U2257 (N_2257,N_2241,N_2220);
nand U2258 (N_2258,N_2238,N_2235);
nor U2259 (N_2259,N_2223,N_2232);
or U2260 (N_2260,N_2244,N_2225);
or U2261 (N_2261,N_2204,N_2200);
nor U2262 (N_2262,N_2214,N_2218);
nand U2263 (N_2263,N_2216,N_2239);
nor U2264 (N_2264,N_2233,N_2213);
nor U2265 (N_2265,N_2228,N_2217);
and U2266 (N_2266,N_2201,N_2237);
nor U2267 (N_2267,N_2246,N_2234);
nand U2268 (N_2268,N_2236,N_2230);
and U2269 (N_2269,N_2219,N_2205);
nand U2270 (N_2270,N_2222,N_2242);
nand U2271 (N_2271,N_2248,N_2207);
nor U2272 (N_2272,N_2206,N_2249);
or U2273 (N_2273,N_2231,N_2227);
nand U2274 (N_2274,N_2247,N_2240);
and U2275 (N_2275,N_2220,N_2219);
or U2276 (N_2276,N_2247,N_2238);
nor U2277 (N_2277,N_2209,N_2214);
nor U2278 (N_2278,N_2236,N_2202);
nand U2279 (N_2279,N_2245,N_2207);
nor U2280 (N_2280,N_2217,N_2245);
and U2281 (N_2281,N_2201,N_2206);
nand U2282 (N_2282,N_2204,N_2217);
nand U2283 (N_2283,N_2227,N_2235);
or U2284 (N_2284,N_2209,N_2213);
nand U2285 (N_2285,N_2245,N_2202);
and U2286 (N_2286,N_2232,N_2200);
or U2287 (N_2287,N_2243,N_2209);
and U2288 (N_2288,N_2204,N_2212);
or U2289 (N_2289,N_2221,N_2248);
nand U2290 (N_2290,N_2235,N_2220);
nor U2291 (N_2291,N_2221,N_2229);
nand U2292 (N_2292,N_2235,N_2202);
nor U2293 (N_2293,N_2220,N_2215);
and U2294 (N_2294,N_2217,N_2244);
nor U2295 (N_2295,N_2233,N_2205);
or U2296 (N_2296,N_2235,N_2223);
nor U2297 (N_2297,N_2235,N_2225);
and U2298 (N_2298,N_2212,N_2210);
and U2299 (N_2299,N_2242,N_2201);
and U2300 (N_2300,N_2279,N_2256);
nor U2301 (N_2301,N_2297,N_2275);
nand U2302 (N_2302,N_2261,N_2262);
or U2303 (N_2303,N_2265,N_2295);
nor U2304 (N_2304,N_2250,N_2287);
and U2305 (N_2305,N_2264,N_2253);
or U2306 (N_2306,N_2291,N_2282);
or U2307 (N_2307,N_2259,N_2252);
or U2308 (N_2308,N_2271,N_2251);
nor U2309 (N_2309,N_2272,N_2292);
and U2310 (N_2310,N_2273,N_2270);
nor U2311 (N_2311,N_2257,N_2268);
nand U2312 (N_2312,N_2278,N_2276);
nor U2313 (N_2313,N_2280,N_2296);
or U2314 (N_2314,N_2263,N_2298);
nand U2315 (N_2315,N_2290,N_2255);
nand U2316 (N_2316,N_2285,N_2269);
or U2317 (N_2317,N_2293,N_2260);
nor U2318 (N_2318,N_2274,N_2289);
and U2319 (N_2319,N_2294,N_2283);
and U2320 (N_2320,N_2299,N_2267);
nor U2321 (N_2321,N_2258,N_2266);
or U2322 (N_2322,N_2281,N_2284);
nor U2323 (N_2323,N_2254,N_2288);
or U2324 (N_2324,N_2277,N_2286);
and U2325 (N_2325,N_2267,N_2260);
nand U2326 (N_2326,N_2273,N_2289);
nand U2327 (N_2327,N_2277,N_2267);
and U2328 (N_2328,N_2258,N_2256);
nor U2329 (N_2329,N_2299,N_2271);
nand U2330 (N_2330,N_2255,N_2275);
or U2331 (N_2331,N_2292,N_2299);
or U2332 (N_2332,N_2268,N_2283);
or U2333 (N_2333,N_2263,N_2258);
nand U2334 (N_2334,N_2255,N_2282);
or U2335 (N_2335,N_2272,N_2288);
nand U2336 (N_2336,N_2251,N_2262);
nand U2337 (N_2337,N_2281,N_2276);
and U2338 (N_2338,N_2298,N_2281);
nand U2339 (N_2339,N_2253,N_2274);
and U2340 (N_2340,N_2282,N_2280);
or U2341 (N_2341,N_2274,N_2254);
and U2342 (N_2342,N_2292,N_2254);
and U2343 (N_2343,N_2297,N_2271);
nand U2344 (N_2344,N_2294,N_2275);
nor U2345 (N_2345,N_2266,N_2280);
nand U2346 (N_2346,N_2268,N_2281);
or U2347 (N_2347,N_2267,N_2263);
and U2348 (N_2348,N_2286,N_2269);
nor U2349 (N_2349,N_2298,N_2260);
or U2350 (N_2350,N_2325,N_2345);
nand U2351 (N_2351,N_2346,N_2330);
or U2352 (N_2352,N_2342,N_2349);
and U2353 (N_2353,N_2316,N_2323);
or U2354 (N_2354,N_2320,N_2313);
and U2355 (N_2355,N_2339,N_2329);
or U2356 (N_2356,N_2309,N_2331);
nand U2357 (N_2357,N_2311,N_2315);
nor U2358 (N_2358,N_2333,N_2338);
nand U2359 (N_2359,N_2317,N_2306);
nand U2360 (N_2360,N_2305,N_2301);
nand U2361 (N_2361,N_2347,N_2310);
or U2362 (N_2362,N_2328,N_2344);
or U2363 (N_2363,N_2318,N_2341);
nand U2364 (N_2364,N_2302,N_2337);
and U2365 (N_2365,N_2343,N_2322);
and U2366 (N_2366,N_2307,N_2326);
and U2367 (N_2367,N_2304,N_2334);
and U2368 (N_2368,N_2321,N_2332);
nor U2369 (N_2369,N_2312,N_2335);
and U2370 (N_2370,N_2319,N_2300);
and U2371 (N_2371,N_2324,N_2348);
nand U2372 (N_2372,N_2303,N_2336);
xor U2373 (N_2373,N_2327,N_2308);
nand U2374 (N_2374,N_2340,N_2314);
or U2375 (N_2375,N_2341,N_2324);
and U2376 (N_2376,N_2333,N_2348);
or U2377 (N_2377,N_2310,N_2321);
and U2378 (N_2378,N_2345,N_2323);
and U2379 (N_2379,N_2303,N_2328);
and U2380 (N_2380,N_2346,N_2337);
and U2381 (N_2381,N_2313,N_2321);
or U2382 (N_2382,N_2305,N_2315);
nand U2383 (N_2383,N_2327,N_2317);
and U2384 (N_2384,N_2336,N_2324);
nand U2385 (N_2385,N_2338,N_2335);
or U2386 (N_2386,N_2313,N_2342);
nand U2387 (N_2387,N_2304,N_2310);
nor U2388 (N_2388,N_2338,N_2304);
and U2389 (N_2389,N_2320,N_2335);
or U2390 (N_2390,N_2340,N_2315);
or U2391 (N_2391,N_2342,N_2337);
nand U2392 (N_2392,N_2301,N_2329);
or U2393 (N_2393,N_2333,N_2331);
nor U2394 (N_2394,N_2301,N_2328);
nand U2395 (N_2395,N_2326,N_2308);
nand U2396 (N_2396,N_2339,N_2334);
nor U2397 (N_2397,N_2312,N_2324);
nor U2398 (N_2398,N_2340,N_2344);
nor U2399 (N_2399,N_2336,N_2307);
xor U2400 (N_2400,N_2393,N_2351);
or U2401 (N_2401,N_2373,N_2381);
and U2402 (N_2402,N_2360,N_2353);
nand U2403 (N_2403,N_2366,N_2371);
or U2404 (N_2404,N_2380,N_2398);
or U2405 (N_2405,N_2355,N_2364);
or U2406 (N_2406,N_2375,N_2391);
nor U2407 (N_2407,N_2363,N_2396);
and U2408 (N_2408,N_2357,N_2394);
nand U2409 (N_2409,N_2372,N_2395);
nand U2410 (N_2410,N_2387,N_2379);
nor U2411 (N_2411,N_2397,N_2359);
or U2412 (N_2412,N_2352,N_2368);
or U2413 (N_2413,N_2385,N_2369);
nor U2414 (N_2414,N_2376,N_2378);
and U2415 (N_2415,N_2370,N_2358);
and U2416 (N_2416,N_2384,N_2361);
or U2417 (N_2417,N_2390,N_2386);
nor U2418 (N_2418,N_2354,N_2382);
or U2419 (N_2419,N_2350,N_2389);
nand U2420 (N_2420,N_2362,N_2377);
nand U2421 (N_2421,N_2356,N_2399);
nor U2422 (N_2422,N_2388,N_2365);
nand U2423 (N_2423,N_2383,N_2367);
nor U2424 (N_2424,N_2374,N_2392);
and U2425 (N_2425,N_2363,N_2385);
nor U2426 (N_2426,N_2367,N_2350);
nor U2427 (N_2427,N_2372,N_2377);
nand U2428 (N_2428,N_2352,N_2379);
or U2429 (N_2429,N_2354,N_2387);
nor U2430 (N_2430,N_2391,N_2393);
and U2431 (N_2431,N_2389,N_2374);
nand U2432 (N_2432,N_2379,N_2380);
nand U2433 (N_2433,N_2352,N_2365);
or U2434 (N_2434,N_2359,N_2388);
and U2435 (N_2435,N_2398,N_2362);
nor U2436 (N_2436,N_2398,N_2396);
or U2437 (N_2437,N_2380,N_2355);
and U2438 (N_2438,N_2391,N_2395);
and U2439 (N_2439,N_2350,N_2395);
and U2440 (N_2440,N_2397,N_2375);
and U2441 (N_2441,N_2388,N_2383);
nor U2442 (N_2442,N_2350,N_2364);
nand U2443 (N_2443,N_2384,N_2396);
or U2444 (N_2444,N_2363,N_2394);
or U2445 (N_2445,N_2394,N_2393);
nor U2446 (N_2446,N_2390,N_2379);
xor U2447 (N_2447,N_2370,N_2355);
nor U2448 (N_2448,N_2387,N_2368);
or U2449 (N_2449,N_2363,N_2360);
and U2450 (N_2450,N_2449,N_2435);
xor U2451 (N_2451,N_2420,N_2416);
nor U2452 (N_2452,N_2423,N_2424);
nor U2453 (N_2453,N_2402,N_2414);
and U2454 (N_2454,N_2413,N_2443);
or U2455 (N_2455,N_2410,N_2418);
or U2456 (N_2456,N_2401,N_2427);
nor U2457 (N_2457,N_2429,N_2422);
nand U2458 (N_2458,N_2448,N_2415);
nor U2459 (N_2459,N_2400,N_2408);
or U2460 (N_2460,N_2428,N_2445);
and U2461 (N_2461,N_2430,N_2431);
nor U2462 (N_2462,N_2409,N_2438);
or U2463 (N_2463,N_2447,N_2437);
nor U2464 (N_2464,N_2406,N_2405);
nand U2465 (N_2465,N_2425,N_2417);
and U2466 (N_2466,N_2439,N_2434);
nor U2467 (N_2467,N_2446,N_2432);
nor U2468 (N_2468,N_2412,N_2421);
nor U2469 (N_2469,N_2411,N_2433);
and U2470 (N_2470,N_2440,N_2426);
nor U2471 (N_2471,N_2403,N_2404);
or U2472 (N_2472,N_2441,N_2436);
and U2473 (N_2473,N_2442,N_2419);
or U2474 (N_2474,N_2407,N_2444);
or U2475 (N_2475,N_2439,N_2402);
or U2476 (N_2476,N_2449,N_2431);
and U2477 (N_2477,N_2407,N_2428);
nand U2478 (N_2478,N_2427,N_2416);
nor U2479 (N_2479,N_2403,N_2406);
nor U2480 (N_2480,N_2428,N_2413);
and U2481 (N_2481,N_2427,N_2409);
nand U2482 (N_2482,N_2406,N_2422);
nor U2483 (N_2483,N_2448,N_2425);
nor U2484 (N_2484,N_2446,N_2404);
nand U2485 (N_2485,N_2440,N_2423);
or U2486 (N_2486,N_2401,N_2422);
or U2487 (N_2487,N_2410,N_2441);
nor U2488 (N_2488,N_2418,N_2430);
nand U2489 (N_2489,N_2420,N_2407);
nor U2490 (N_2490,N_2415,N_2405);
nand U2491 (N_2491,N_2436,N_2434);
or U2492 (N_2492,N_2421,N_2424);
and U2493 (N_2493,N_2411,N_2435);
nand U2494 (N_2494,N_2436,N_2411);
and U2495 (N_2495,N_2411,N_2437);
nand U2496 (N_2496,N_2401,N_2407);
and U2497 (N_2497,N_2409,N_2439);
or U2498 (N_2498,N_2447,N_2405);
nor U2499 (N_2499,N_2411,N_2409);
and U2500 (N_2500,N_2465,N_2458);
or U2501 (N_2501,N_2490,N_2464);
nor U2502 (N_2502,N_2478,N_2472);
nor U2503 (N_2503,N_2494,N_2496);
and U2504 (N_2504,N_2477,N_2469);
nor U2505 (N_2505,N_2452,N_2468);
and U2506 (N_2506,N_2454,N_2484);
or U2507 (N_2507,N_2479,N_2488);
and U2508 (N_2508,N_2491,N_2470);
and U2509 (N_2509,N_2483,N_2451);
and U2510 (N_2510,N_2460,N_2467);
and U2511 (N_2511,N_2497,N_2492);
nand U2512 (N_2512,N_2485,N_2473);
or U2513 (N_2513,N_2493,N_2471);
or U2514 (N_2514,N_2450,N_2475);
nor U2515 (N_2515,N_2474,N_2462);
or U2516 (N_2516,N_2456,N_2495);
and U2517 (N_2517,N_2476,N_2481);
nand U2518 (N_2518,N_2489,N_2457);
and U2519 (N_2519,N_2463,N_2499);
nor U2520 (N_2520,N_2453,N_2498);
or U2521 (N_2521,N_2480,N_2455);
nor U2522 (N_2522,N_2466,N_2459);
or U2523 (N_2523,N_2482,N_2487);
and U2524 (N_2524,N_2461,N_2486);
or U2525 (N_2525,N_2462,N_2475);
nand U2526 (N_2526,N_2482,N_2456);
and U2527 (N_2527,N_2496,N_2486);
nor U2528 (N_2528,N_2490,N_2458);
nor U2529 (N_2529,N_2493,N_2487);
nand U2530 (N_2530,N_2484,N_2479);
nand U2531 (N_2531,N_2477,N_2454);
nand U2532 (N_2532,N_2467,N_2451);
or U2533 (N_2533,N_2460,N_2478);
or U2534 (N_2534,N_2492,N_2457);
and U2535 (N_2535,N_2475,N_2473);
nor U2536 (N_2536,N_2496,N_2459);
or U2537 (N_2537,N_2472,N_2471);
or U2538 (N_2538,N_2478,N_2494);
and U2539 (N_2539,N_2459,N_2454);
and U2540 (N_2540,N_2484,N_2475);
nand U2541 (N_2541,N_2465,N_2496);
nor U2542 (N_2542,N_2480,N_2488);
nand U2543 (N_2543,N_2478,N_2473);
and U2544 (N_2544,N_2463,N_2477);
nand U2545 (N_2545,N_2488,N_2451);
or U2546 (N_2546,N_2468,N_2487);
nand U2547 (N_2547,N_2474,N_2481);
nor U2548 (N_2548,N_2450,N_2489);
nor U2549 (N_2549,N_2456,N_2484);
or U2550 (N_2550,N_2525,N_2537);
nor U2551 (N_2551,N_2517,N_2514);
or U2552 (N_2552,N_2541,N_2504);
and U2553 (N_2553,N_2500,N_2538);
and U2554 (N_2554,N_2507,N_2531);
and U2555 (N_2555,N_2547,N_2535);
nand U2556 (N_2556,N_2509,N_2527);
and U2557 (N_2557,N_2521,N_2530);
and U2558 (N_2558,N_2518,N_2524);
or U2559 (N_2559,N_2512,N_2528);
nor U2560 (N_2560,N_2522,N_2545);
nand U2561 (N_2561,N_2532,N_2536);
nand U2562 (N_2562,N_2506,N_2542);
nand U2563 (N_2563,N_2533,N_2529);
nand U2564 (N_2564,N_2502,N_2503);
or U2565 (N_2565,N_2544,N_2516);
and U2566 (N_2566,N_2539,N_2513);
nand U2567 (N_2567,N_2510,N_2508);
and U2568 (N_2568,N_2511,N_2515);
nand U2569 (N_2569,N_2526,N_2523);
nor U2570 (N_2570,N_2534,N_2543);
nand U2571 (N_2571,N_2520,N_2519);
or U2572 (N_2572,N_2540,N_2546);
or U2573 (N_2573,N_2501,N_2549);
and U2574 (N_2574,N_2548,N_2505);
nand U2575 (N_2575,N_2516,N_2549);
nor U2576 (N_2576,N_2520,N_2544);
nand U2577 (N_2577,N_2537,N_2540);
or U2578 (N_2578,N_2543,N_2504);
and U2579 (N_2579,N_2501,N_2512);
and U2580 (N_2580,N_2509,N_2514);
nor U2581 (N_2581,N_2519,N_2501);
nor U2582 (N_2582,N_2531,N_2512);
nor U2583 (N_2583,N_2514,N_2519);
nand U2584 (N_2584,N_2526,N_2500);
nor U2585 (N_2585,N_2535,N_2508);
nand U2586 (N_2586,N_2514,N_2546);
nor U2587 (N_2587,N_2531,N_2539);
or U2588 (N_2588,N_2524,N_2519);
nand U2589 (N_2589,N_2532,N_2537);
nand U2590 (N_2590,N_2503,N_2519);
and U2591 (N_2591,N_2534,N_2544);
or U2592 (N_2592,N_2533,N_2510);
nand U2593 (N_2593,N_2530,N_2522);
or U2594 (N_2594,N_2538,N_2522);
nand U2595 (N_2595,N_2526,N_2528);
xor U2596 (N_2596,N_2541,N_2536);
and U2597 (N_2597,N_2534,N_2518);
or U2598 (N_2598,N_2548,N_2515);
or U2599 (N_2599,N_2525,N_2515);
nand U2600 (N_2600,N_2581,N_2567);
nand U2601 (N_2601,N_2588,N_2552);
and U2602 (N_2602,N_2561,N_2577);
or U2603 (N_2603,N_2571,N_2592);
nor U2604 (N_2604,N_2560,N_2597);
nand U2605 (N_2605,N_2591,N_2565);
nand U2606 (N_2606,N_2579,N_2587);
nand U2607 (N_2607,N_2582,N_2596);
or U2608 (N_2608,N_2550,N_2583);
nor U2609 (N_2609,N_2558,N_2557);
nand U2610 (N_2610,N_2568,N_2573);
nand U2611 (N_2611,N_2563,N_2559);
or U2612 (N_2612,N_2595,N_2555);
nand U2613 (N_2613,N_2556,N_2585);
nand U2614 (N_2614,N_2578,N_2594);
and U2615 (N_2615,N_2598,N_2569);
nand U2616 (N_2616,N_2554,N_2551);
or U2617 (N_2617,N_2590,N_2566);
or U2618 (N_2618,N_2584,N_2593);
and U2619 (N_2619,N_2589,N_2564);
or U2620 (N_2620,N_2553,N_2570);
nor U2621 (N_2621,N_2562,N_2575);
and U2622 (N_2622,N_2572,N_2580);
or U2623 (N_2623,N_2599,N_2586);
nand U2624 (N_2624,N_2574,N_2576);
nand U2625 (N_2625,N_2560,N_2553);
nor U2626 (N_2626,N_2585,N_2560);
nand U2627 (N_2627,N_2571,N_2599);
or U2628 (N_2628,N_2582,N_2567);
nor U2629 (N_2629,N_2560,N_2578);
nand U2630 (N_2630,N_2552,N_2554);
nor U2631 (N_2631,N_2574,N_2577);
nor U2632 (N_2632,N_2583,N_2597);
nand U2633 (N_2633,N_2583,N_2566);
nor U2634 (N_2634,N_2565,N_2575);
and U2635 (N_2635,N_2552,N_2587);
nand U2636 (N_2636,N_2555,N_2569);
and U2637 (N_2637,N_2550,N_2573);
and U2638 (N_2638,N_2582,N_2578);
nand U2639 (N_2639,N_2573,N_2593);
or U2640 (N_2640,N_2550,N_2585);
and U2641 (N_2641,N_2567,N_2569);
nand U2642 (N_2642,N_2559,N_2550);
or U2643 (N_2643,N_2558,N_2552);
and U2644 (N_2644,N_2580,N_2588);
nand U2645 (N_2645,N_2594,N_2562);
and U2646 (N_2646,N_2562,N_2581);
and U2647 (N_2647,N_2596,N_2561);
nand U2648 (N_2648,N_2581,N_2554);
nor U2649 (N_2649,N_2586,N_2567);
xnor U2650 (N_2650,N_2629,N_2603);
nor U2651 (N_2651,N_2649,N_2611);
and U2652 (N_2652,N_2616,N_2642);
nand U2653 (N_2653,N_2627,N_2631);
nor U2654 (N_2654,N_2610,N_2632);
nand U2655 (N_2655,N_2620,N_2615);
nor U2656 (N_2656,N_2606,N_2612);
and U2657 (N_2657,N_2628,N_2645);
or U2658 (N_2658,N_2604,N_2617);
and U2659 (N_2659,N_2647,N_2637);
nor U2660 (N_2660,N_2636,N_2613);
or U2661 (N_2661,N_2635,N_2634);
nor U2662 (N_2662,N_2605,N_2646);
or U2663 (N_2663,N_2633,N_2601);
and U2664 (N_2664,N_2641,N_2623);
nand U2665 (N_2665,N_2643,N_2622);
nor U2666 (N_2666,N_2640,N_2624);
and U2667 (N_2667,N_2619,N_2626);
or U2668 (N_2668,N_2621,N_2609);
nand U2669 (N_2669,N_2608,N_2607);
and U2670 (N_2670,N_2630,N_2648);
nand U2671 (N_2671,N_2614,N_2600);
or U2672 (N_2672,N_2644,N_2618);
and U2673 (N_2673,N_2638,N_2639);
or U2674 (N_2674,N_2602,N_2625);
or U2675 (N_2675,N_2615,N_2638);
nand U2676 (N_2676,N_2620,N_2640);
or U2677 (N_2677,N_2612,N_2636);
or U2678 (N_2678,N_2630,N_2634);
nand U2679 (N_2679,N_2616,N_2604);
xnor U2680 (N_2680,N_2648,N_2647);
nand U2681 (N_2681,N_2625,N_2647);
and U2682 (N_2682,N_2631,N_2638);
nand U2683 (N_2683,N_2637,N_2646);
and U2684 (N_2684,N_2620,N_2633);
nand U2685 (N_2685,N_2642,N_2644);
nand U2686 (N_2686,N_2608,N_2638);
or U2687 (N_2687,N_2623,N_2626);
or U2688 (N_2688,N_2649,N_2647);
and U2689 (N_2689,N_2606,N_2642);
nor U2690 (N_2690,N_2621,N_2633);
or U2691 (N_2691,N_2600,N_2646);
and U2692 (N_2692,N_2631,N_2605);
nand U2693 (N_2693,N_2608,N_2625);
or U2694 (N_2694,N_2649,N_2638);
and U2695 (N_2695,N_2615,N_2607);
nand U2696 (N_2696,N_2622,N_2628);
and U2697 (N_2697,N_2647,N_2608);
nor U2698 (N_2698,N_2600,N_2641);
nand U2699 (N_2699,N_2630,N_2621);
or U2700 (N_2700,N_2674,N_2650);
and U2701 (N_2701,N_2662,N_2665);
nand U2702 (N_2702,N_2688,N_2660);
nor U2703 (N_2703,N_2655,N_2664);
or U2704 (N_2704,N_2669,N_2651);
or U2705 (N_2705,N_2698,N_2656);
nor U2706 (N_2706,N_2676,N_2696);
and U2707 (N_2707,N_2654,N_2687);
or U2708 (N_2708,N_2658,N_2683);
or U2709 (N_2709,N_2661,N_2670);
or U2710 (N_2710,N_2668,N_2657);
nand U2711 (N_2711,N_2666,N_2671);
nand U2712 (N_2712,N_2695,N_2692);
or U2713 (N_2713,N_2685,N_2697);
nand U2714 (N_2714,N_2653,N_2684);
and U2715 (N_2715,N_2673,N_2678);
or U2716 (N_2716,N_2652,N_2691);
nand U2717 (N_2717,N_2667,N_2675);
nor U2718 (N_2718,N_2679,N_2663);
and U2719 (N_2719,N_2659,N_2699);
or U2720 (N_2720,N_2680,N_2672);
nor U2721 (N_2721,N_2690,N_2682);
nand U2722 (N_2722,N_2686,N_2694);
nor U2723 (N_2723,N_2677,N_2693);
and U2724 (N_2724,N_2681,N_2689);
or U2725 (N_2725,N_2680,N_2659);
nor U2726 (N_2726,N_2654,N_2671);
nor U2727 (N_2727,N_2654,N_2679);
nand U2728 (N_2728,N_2655,N_2671);
and U2729 (N_2729,N_2661,N_2672);
and U2730 (N_2730,N_2668,N_2692);
and U2731 (N_2731,N_2688,N_2677);
or U2732 (N_2732,N_2662,N_2684);
nand U2733 (N_2733,N_2650,N_2665);
nor U2734 (N_2734,N_2689,N_2694);
and U2735 (N_2735,N_2660,N_2694);
or U2736 (N_2736,N_2675,N_2659);
nand U2737 (N_2737,N_2678,N_2698);
nand U2738 (N_2738,N_2665,N_2676);
nand U2739 (N_2739,N_2688,N_2681);
nor U2740 (N_2740,N_2696,N_2678);
nor U2741 (N_2741,N_2659,N_2658);
nand U2742 (N_2742,N_2662,N_2658);
or U2743 (N_2743,N_2678,N_2669);
and U2744 (N_2744,N_2693,N_2662);
and U2745 (N_2745,N_2680,N_2654);
nand U2746 (N_2746,N_2678,N_2670);
or U2747 (N_2747,N_2683,N_2688);
or U2748 (N_2748,N_2677,N_2672);
and U2749 (N_2749,N_2682,N_2668);
or U2750 (N_2750,N_2704,N_2706);
or U2751 (N_2751,N_2712,N_2734);
and U2752 (N_2752,N_2740,N_2709);
and U2753 (N_2753,N_2726,N_2747);
nor U2754 (N_2754,N_2718,N_2703);
or U2755 (N_2755,N_2736,N_2707);
nand U2756 (N_2756,N_2732,N_2719);
nand U2757 (N_2757,N_2721,N_2743);
nor U2758 (N_2758,N_2723,N_2737);
or U2759 (N_2759,N_2730,N_2700);
nor U2760 (N_2760,N_2715,N_2711);
and U2761 (N_2761,N_2705,N_2716);
nor U2762 (N_2762,N_2741,N_2701);
nor U2763 (N_2763,N_2745,N_2713);
and U2764 (N_2764,N_2727,N_2733);
nand U2765 (N_2765,N_2748,N_2739);
or U2766 (N_2766,N_2714,N_2722);
or U2767 (N_2767,N_2731,N_2717);
or U2768 (N_2768,N_2702,N_2708);
nor U2769 (N_2769,N_2746,N_2749);
or U2770 (N_2770,N_2724,N_2742);
nand U2771 (N_2771,N_2729,N_2744);
and U2772 (N_2772,N_2738,N_2710);
nor U2773 (N_2773,N_2720,N_2728);
nor U2774 (N_2774,N_2725,N_2735);
or U2775 (N_2775,N_2712,N_2746);
nor U2776 (N_2776,N_2718,N_2716);
nand U2777 (N_2777,N_2726,N_2748);
and U2778 (N_2778,N_2732,N_2711);
nor U2779 (N_2779,N_2724,N_2709);
nand U2780 (N_2780,N_2729,N_2740);
and U2781 (N_2781,N_2720,N_2744);
nand U2782 (N_2782,N_2711,N_2729);
and U2783 (N_2783,N_2705,N_2717);
nor U2784 (N_2784,N_2713,N_2704);
nor U2785 (N_2785,N_2730,N_2719);
nand U2786 (N_2786,N_2723,N_2704);
or U2787 (N_2787,N_2723,N_2713);
or U2788 (N_2788,N_2726,N_2742);
and U2789 (N_2789,N_2748,N_2707);
and U2790 (N_2790,N_2708,N_2707);
or U2791 (N_2791,N_2739,N_2732);
or U2792 (N_2792,N_2722,N_2723);
or U2793 (N_2793,N_2727,N_2718);
nor U2794 (N_2794,N_2710,N_2745);
or U2795 (N_2795,N_2721,N_2706);
nor U2796 (N_2796,N_2729,N_2727);
nor U2797 (N_2797,N_2740,N_2746);
nand U2798 (N_2798,N_2736,N_2727);
nor U2799 (N_2799,N_2704,N_2745);
nand U2800 (N_2800,N_2791,N_2767);
nor U2801 (N_2801,N_2755,N_2789);
nor U2802 (N_2802,N_2783,N_2772);
nand U2803 (N_2803,N_2761,N_2781);
and U2804 (N_2804,N_2790,N_2794);
nand U2805 (N_2805,N_2753,N_2759);
nand U2806 (N_2806,N_2752,N_2793);
nand U2807 (N_2807,N_2758,N_2774);
nand U2808 (N_2808,N_2750,N_2769);
or U2809 (N_2809,N_2766,N_2751);
nor U2810 (N_2810,N_2787,N_2785);
and U2811 (N_2811,N_2760,N_2780);
or U2812 (N_2812,N_2778,N_2797);
and U2813 (N_2813,N_2754,N_2796);
nor U2814 (N_2814,N_2756,N_2792);
nor U2815 (N_2815,N_2779,N_2773);
and U2816 (N_2816,N_2784,N_2762);
nor U2817 (N_2817,N_2799,N_2777);
and U2818 (N_2818,N_2770,N_2771);
or U2819 (N_2819,N_2798,N_2765);
and U2820 (N_2820,N_2763,N_2775);
nor U2821 (N_2821,N_2788,N_2757);
and U2822 (N_2822,N_2786,N_2768);
nor U2823 (N_2823,N_2782,N_2764);
nand U2824 (N_2824,N_2776,N_2795);
nor U2825 (N_2825,N_2785,N_2798);
and U2826 (N_2826,N_2789,N_2762);
nand U2827 (N_2827,N_2786,N_2774);
nand U2828 (N_2828,N_2759,N_2774);
and U2829 (N_2829,N_2793,N_2792);
nor U2830 (N_2830,N_2766,N_2784);
or U2831 (N_2831,N_2780,N_2770);
nor U2832 (N_2832,N_2775,N_2752);
and U2833 (N_2833,N_2785,N_2791);
or U2834 (N_2834,N_2787,N_2794);
or U2835 (N_2835,N_2786,N_2762);
or U2836 (N_2836,N_2768,N_2781);
or U2837 (N_2837,N_2781,N_2790);
nor U2838 (N_2838,N_2779,N_2778);
nand U2839 (N_2839,N_2766,N_2758);
or U2840 (N_2840,N_2787,N_2772);
nor U2841 (N_2841,N_2772,N_2752);
nor U2842 (N_2842,N_2783,N_2794);
or U2843 (N_2843,N_2783,N_2760);
nor U2844 (N_2844,N_2773,N_2795);
and U2845 (N_2845,N_2776,N_2793);
or U2846 (N_2846,N_2771,N_2787);
and U2847 (N_2847,N_2791,N_2774);
and U2848 (N_2848,N_2796,N_2791);
and U2849 (N_2849,N_2772,N_2764);
or U2850 (N_2850,N_2803,N_2843);
nor U2851 (N_2851,N_2831,N_2835);
and U2852 (N_2852,N_2813,N_2829);
and U2853 (N_2853,N_2810,N_2818);
nand U2854 (N_2854,N_2809,N_2802);
or U2855 (N_2855,N_2837,N_2820);
or U2856 (N_2856,N_2825,N_2833);
nand U2857 (N_2857,N_2847,N_2840);
nor U2858 (N_2858,N_2814,N_2832);
nand U2859 (N_2859,N_2822,N_2821);
and U2860 (N_2860,N_2806,N_2836);
or U2861 (N_2861,N_2808,N_2804);
and U2862 (N_2862,N_2848,N_2817);
or U2863 (N_2863,N_2801,N_2841);
nand U2864 (N_2864,N_2828,N_2842);
or U2865 (N_2865,N_2819,N_2834);
nand U2866 (N_2866,N_2826,N_2845);
or U2867 (N_2867,N_2839,N_2805);
nor U2868 (N_2868,N_2812,N_2800);
nor U2869 (N_2869,N_2838,N_2823);
nor U2870 (N_2870,N_2815,N_2811);
nand U2871 (N_2871,N_2849,N_2816);
or U2872 (N_2872,N_2807,N_2844);
nor U2873 (N_2873,N_2846,N_2827);
and U2874 (N_2874,N_2830,N_2824);
or U2875 (N_2875,N_2814,N_2823);
nor U2876 (N_2876,N_2832,N_2819);
nand U2877 (N_2877,N_2815,N_2814);
nor U2878 (N_2878,N_2811,N_2819);
nor U2879 (N_2879,N_2807,N_2835);
nor U2880 (N_2880,N_2819,N_2842);
nand U2881 (N_2881,N_2844,N_2804);
nand U2882 (N_2882,N_2806,N_2801);
and U2883 (N_2883,N_2847,N_2849);
nor U2884 (N_2884,N_2808,N_2810);
and U2885 (N_2885,N_2802,N_2815);
or U2886 (N_2886,N_2801,N_2831);
nor U2887 (N_2887,N_2823,N_2804);
nor U2888 (N_2888,N_2809,N_2801);
nor U2889 (N_2889,N_2804,N_2819);
nor U2890 (N_2890,N_2848,N_2834);
and U2891 (N_2891,N_2803,N_2801);
and U2892 (N_2892,N_2806,N_2813);
nand U2893 (N_2893,N_2837,N_2845);
nor U2894 (N_2894,N_2834,N_2839);
and U2895 (N_2895,N_2834,N_2824);
or U2896 (N_2896,N_2816,N_2845);
nand U2897 (N_2897,N_2842,N_2812);
nor U2898 (N_2898,N_2805,N_2842);
xnor U2899 (N_2899,N_2824,N_2841);
nor U2900 (N_2900,N_2879,N_2893);
nor U2901 (N_2901,N_2890,N_2870);
nor U2902 (N_2902,N_2882,N_2884);
and U2903 (N_2903,N_2871,N_2850);
xnor U2904 (N_2904,N_2873,N_2862);
nand U2905 (N_2905,N_2876,N_2854);
nor U2906 (N_2906,N_2898,N_2894);
or U2907 (N_2907,N_2851,N_2863);
and U2908 (N_2908,N_2888,N_2864);
nor U2909 (N_2909,N_2869,N_2896);
nand U2910 (N_2910,N_2860,N_2880);
or U2911 (N_2911,N_2866,N_2856);
nor U2912 (N_2912,N_2899,N_2881);
or U2913 (N_2913,N_2878,N_2886);
or U2914 (N_2914,N_2877,N_2858);
nand U2915 (N_2915,N_2855,N_2865);
and U2916 (N_2916,N_2895,N_2892);
and U2917 (N_2917,N_2891,N_2897);
or U2918 (N_2918,N_2857,N_2874);
and U2919 (N_2919,N_2889,N_2852);
nand U2920 (N_2920,N_2867,N_2861);
and U2921 (N_2921,N_2859,N_2883);
nor U2922 (N_2922,N_2887,N_2868);
and U2923 (N_2923,N_2853,N_2885);
or U2924 (N_2924,N_2875,N_2872);
nand U2925 (N_2925,N_2890,N_2884);
nand U2926 (N_2926,N_2890,N_2871);
nor U2927 (N_2927,N_2884,N_2879);
and U2928 (N_2928,N_2898,N_2861);
and U2929 (N_2929,N_2889,N_2871);
or U2930 (N_2930,N_2869,N_2857);
nand U2931 (N_2931,N_2876,N_2890);
nor U2932 (N_2932,N_2868,N_2896);
and U2933 (N_2933,N_2864,N_2884);
or U2934 (N_2934,N_2888,N_2890);
nor U2935 (N_2935,N_2873,N_2889);
nand U2936 (N_2936,N_2895,N_2853);
nor U2937 (N_2937,N_2873,N_2899);
or U2938 (N_2938,N_2878,N_2864);
nor U2939 (N_2939,N_2888,N_2857);
nand U2940 (N_2940,N_2888,N_2852);
nor U2941 (N_2941,N_2862,N_2872);
nor U2942 (N_2942,N_2874,N_2863);
and U2943 (N_2943,N_2869,N_2893);
and U2944 (N_2944,N_2856,N_2895);
nand U2945 (N_2945,N_2871,N_2875);
and U2946 (N_2946,N_2896,N_2872);
and U2947 (N_2947,N_2895,N_2878);
or U2948 (N_2948,N_2895,N_2896);
or U2949 (N_2949,N_2878,N_2877);
nor U2950 (N_2950,N_2912,N_2909);
nand U2951 (N_2951,N_2928,N_2920);
or U2952 (N_2952,N_2914,N_2936);
or U2953 (N_2953,N_2934,N_2902);
or U2954 (N_2954,N_2903,N_2905);
or U2955 (N_2955,N_2901,N_2938);
nor U2956 (N_2956,N_2910,N_2923);
and U2957 (N_2957,N_2916,N_2939);
nand U2958 (N_2958,N_2940,N_2933);
or U2959 (N_2959,N_2935,N_2949);
nand U2960 (N_2960,N_2917,N_2913);
and U2961 (N_2961,N_2915,N_2926);
nand U2962 (N_2962,N_2932,N_2948);
and U2963 (N_2963,N_2921,N_2919);
or U2964 (N_2964,N_2929,N_2942);
or U2965 (N_2965,N_2922,N_2918);
nand U2966 (N_2966,N_2945,N_2911);
nand U2967 (N_2967,N_2931,N_2943);
nand U2968 (N_2968,N_2946,N_2907);
or U2969 (N_2969,N_2924,N_2941);
nor U2970 (N_2970,N_2925,N_2904);
nand U2971 (N_2971,N_2944,N_2908);
or U2972 (N_2972,N_2937,N_2927);
or U2973 (N_2973,N_2906,N_2930);
nor U2974 (N_2974,N_2947,N_2900);
or U2975 (N_2975,N_2919,N_2901);
or U2976 (N_2976,N_2938,N_2936);
or U2977 (N_2977,N_2901,N_2915);
nand U2978 (N_2978,N_2948,N_2919);
and U2979 (N_2979,N_2902,N_2907);
or U2980 (N_2980,N_2909,N_2948);
and U2981 (N_2981,N_2914,N_2949);
and U2982 (N_2982,N_2914,N_2910);
nand U2983 (N_2983,N_2911,N_2905);
and U2984 (N_2984,N_2912,N_2949);
and U2985 (N_2985,N_2920,N_2947);
and U2986 (N_2986,N_2913,N_2911);
and U2987 (N_2987,N_2930,N_2936);
or U2988 (N_2988,N_2924,N_2901);
and U2989 (N_2989,N_2914,N_2931);
nor U2990 (N_2990,N_2921,N_2935);
and U2991 (N_2991,N_2943,N_2926);
or U2992 (N_2992,N_2932,N_2910);
nor U2993 (N_2993,N_2910,N_2919);
nand U2994 (N_2994,N_2926,N_2913);
nor U2995 (N_2995,N_2948,N_2949);
nand U2996 (N_2996,N_2948,N_2904);
or U2997 (N_2997,N_2941,N_2917);
nand U2998 (N_2998,N_2925,N_2912);
nand U2999 (N_2999,N_2901,N_2943);
nor UO_0 (O_0,N_2997,N_2980);
and UO_1 (O_1,N_2968,N_2956);
nor UO_2 (O_2,N_2961,N_2972);
and UO_3 (O_3,N_2969,N_2979);
or UO_4 (O_4,N_2976,N_2996);
or UO_5 (O_5,N_2966,N_2965);
and UO_6 (O_6,N_2984,N_2987);
nor UO_7 (O_7,N_2981,N_2994);
nor UO_8 (O_8,N_2974,N_2975);
nor UO_9 (O_9,N_2953,N_2998);
nor UO_10 (O_10,N_2995,N_2977);
and UO_11 (O_11,N_2999,N_2991);
nor UO_12 (O_12,N_2954,N_2967);
and UO_13 (O_13,N_2951,N_2959);
nor UO_14 (O_14,N_2964,N_2960);
nor UO_15 (O_15,N_2992,N_2978);
nand UO_16 (O_16,N_2973,N_2990);
nor UO_17 (O_17,N_2950,N_2957);
nand UO_18 (O_18,N_2983,N_2989);
nand UO_19 (O_19,N_2955,N_2988);
and UO_20 (O_20,N_2971,N_2986);
nand UO_21 (O_21,N_2952,N_2985);
and UO_22 (O_22,N_2982,N_2962);
or UO_23 (O_23,N_2970,N_2963);
nor UO_24 (O_24,N_2993,N_2958);
nand UO_25 (O_25,N_2974,N_2953);
and UO_26 (O_26,N_2992,N_2979);
or UO_27 (O_27,N_2987,N_2962);
and UO_28 (O_28,N_2959,N_2968);
nor UO_29 (O_29,N_2969,N_2951);
and UO_30 (O_30,N_2994,N_2976);
and UO_31 (O_31,N_2995,N_2999);
nor UO_32 (O_32,N_2979,N_2955);
nand UO_33 (O_33,N_2950,N_2969);
or UO_34 (O_34,N_2997,N_2989);
and UO_35 (O_35,N_2994,N_2968);
nor UO_36 (O_36,N_2982,N_2990);
nand UO_37 (O_37,N_2976,N_2964);
nand UO_38 (O_38,N_2991,N_2975);
and UO_39 (O_39,N_2979,N_2953);
nand UO_40 (O_40,N_2983,N_2999);
nand UO_41 (O_41,N_2984,N_2960);
and UO_42 (O_42,N_2962,N_2979);
nand UO_43 (O_43,N_2990,N_2958);
nor UO_44 (O_44,N_2996,N_2966);
and UO_45 (O_45,N_2984,N_2994);
or UO_46 (O_46,N_2980,N_2999);
nand UO_47 (O_47,N_2965,N_2984);
or UO_48 (O_48,N_2992,N_2963);
or UO_49 (O_49,N_2978,N_2981);
nor UO_50 (O_50,N_2953,N_2981);
or UO_51 (O_51,N_2985,N_2982);
nor UO_52 (O_52,N_2993,N_2976);
nor UO_53 (O_53,N_2981,N_2998);
and UO_54 (O_54,N_2996,N_2990);
or UO_55 (O_55,N_2959,N_2953);
nor UO_56 (O_56,N_2979,N_2960);
and UO_57 (O_57,N_2999,N_2977);
and UO_58 (O_58,N_2963,N_2967);
nand UO_59 (O_59,N_2998,N_2962);
nand UO_60 (O_60,N_2978,N_2967);
nand UO_61 (O_61,N_2966,N_2957);
nand UO_62 (O_62,N_2950,N_2952);
nand UO_63 (O_63,N_2969,N_2973);
nand UO_64 (O_64,N_2993,N_2966);
and UO_65 (O_65,N_2968,N_2985);
nand UO_66 (O_66,N_2961,N_2995);
or UO_67 (O_67,N_2978,N_2953);
nor UO_68 (O_68,N_2988,N_2974);
and UO_69 (O_69,N_2977,N_2979);
nand UO_70 (O_70,N_2970,N_2998);
nor UO_71 (O_71,N_2959,N_2981);
or UO_72 (O_72,N_2953,N_2992);
or UO_73 (O_73,N_2979,N_2980);
or UO_74 (O_74,N_2956,N_2994);
or UO_75 (O_75,N_2964,N_2961);
or UO_76 (O_76,N_2959,N_2958);
nor UO_77 (O_77,N_2974,N_2996);
and UO_78 (O_78,N_2987,N_2998);
nor UO_79 (O_79,N_2986,N_2973);
nand UO_80 (O_80,N_2973,N_2956);
nor UO_81 (O_81,N_2998,N_2971);
or UO_82 (O_82,N_2992,N_2973);
nor UO_83 (O_83,N_2950,N_2953);
or UO_84 (O_84,N_2968,N_2987);
or UO_85 (O_85,N_2977,N_2953);
nor UO_86 (O_86,N_2979,N_2990);
or UO_87 (O_87,N_2954,N_2990);
or UO_88 (O_88,N_2960,N_2968);
nand UO_89 (O_89,N_2967,N_2990);
nor UO_90 (O_90,N_2997,N_2964);
and UO_91 (O_91,N_2955,N_2996);
nand UO_92 (O_92,N_2962,N_2983);
nand UO_93 (O_93,N_2951,N_2950);
nand UO_94 (O_94,N_2997,N_2951);
nor UO_95 (O_95,N_2987,N_2972);
and UO_96 (O_96,N_2999,N_2982);
nand UO_97 (O_97,N_2986,N_2998);
nand UO_98 (O_98,N_2978,N_2997);
nor UO_99 (O_99,N_2992,N_2988);
nand UO_100 (O_100,N_2962,N_2951);
and UO_101 (O_101,N_2976,N_2967);
or UO_102 (O_102,N_2978,N_2971);
nor UO_103 (O_103,N_2979,N_2981);
nor UO_104 (O_104,N_2957,N_2956);
nor UO_105 (O_105,N_2957,N_2976);
nor UO_106 (O_106,N_2957,N_2993);
nand UO_107 (O_107,N_2997,N_2995);
nor UO_108 (O_108,N_2980,N_2984);
and UO_109 (O_109,N_2963,N_2991);
nand UO_110 (O_110,N_2971,N_2989);
and UO_111 (O_111,N_2955,N_2987);
or UO_112 (O_112,N_2952,N_2983);
or UO_113 (O_113,N_2980,N_2983);
or UO_114 (O_114,N_2997,N_2987);
and UO_115 (O_115,N_2967,N_2953);
or UO_116 (O_116,N_2970,N_2969);
or UO_117 (O_117,N_2964,N_2991);
nand UO_118 (O_118,N_2974,N_2994);
nand UO_119 (O_119,N_2980,N_2976);
or UO_120 (O_120,N_2989,N_2990);
nand UO_121 (O_121,N_2992,N_2998);
nand UO_122 (O_122,N_2971,N_2987);
nor UO_123 (O_123,N_2963,N_2952);
nor UO_124 (O_124,N_2986,N_2985);
nor UO_125 (O_125,N_2998,N_2955);
nor UO_126 (O_126,N_2980,N_2982);
nor UO_127 (O_127,N_2999,N_2986);
xor UO_128 (O_128,N_2961,N_2965);
nand UO_129 (O_129,N_2959,N_2986);
nor UO_130 (O_130,N_2994,N_2961);
and UO_131 (O_131,N_2975,N_2996);
and UO_132 (O_132,N_2995,N_2950);
or UO_133 (O_133,N_2951,N_2973);
nor UO_134 (O_134,N_2950,N_2982);
or UO_135 (O_135,N_2994,N_2972);
nand UO_136 (O_136,N_2993,N_2977);
nand UO_137 (O_137,N_2969,N_2980);
or UO_138 (O_138,N_2976,N_2968);
nand UO_139 (O_139,N_2956,N_2971);
nand UO_140 (O_140,N_2997,N_2988);
or UO_141 (O_141,N_2951,N_2980);
or UO_142 (O_142,N_2982,N_2974);
or UO_143 (O_143,N_2984,N_2950);
or UO_144 (O_144,N_2985,N_2962);
nor UO_145 (O_145,N_2958,N_2965);
nor UO_146 (O_146,N_2964,N_2968);
nor UO_147 (O_147,N_2952,N_2975);
nor UO_148 (O_148,N_2952,N_2964);
and UO_149 (O_149,N_2993,N_2961);
or UO_150 (O_150,N_2985,N_2988);
nor UO_151 (O_151,N_2964,N_2978);
nor UO_152 (O_152,N_2999,N_2974);
nor UO_153 (O_153,N_2985,N_2996);
nor UO_154 (O_154,N_2999,N_2955);
nor UO_155 (O_155,N_2968,N_2999);
and UO_156 (O_156,N_2967,N_2985);
nand UO_157 (O_157,N_2978,N_2952);
or UO_158 (O_158,N_2957,N_2973);
nand UO_159 (O_159,N_2997,N_2952);
and UO_160 (O_160,N_2983,N_2993);
nor UO_161 (O_161,N_2976,N_2954);
or UO_162 (O_162,N_2974,N_2952);
nand UO_163 (O_163,N_2984,N_2973);
nor UO_164 (O_164,N_2964,N_2992);
and UO_165 (O_165,N_2999,N_2954);
or UO_166 (O_166,N_2951,N_2995);
nand UO_167 (O_167,N_2963,N_2956);
nand UO_168 (O_168,N_2958,N_2968);
nand UO_169 (O_169,N_2952,N_2973);
and UO_170 (O_170,N_2960,N_2985);
or UO_171 (O_171,N_2956,N_2988);
or UO_172 (O_172,N_2954,N_2958);
nand UO_173 (O_173,N_2968,N_2970);
or UO_174 (O_174,N_2990,N_2976);
and UO_175 (O_175,N_2986,N_2956);
nand UO_176 (O_176,N_2951,N_2970);
nand UO_177 (O_177,N_2979,N_2967);
nor UO_178 (O_178,N_2964,N_2975);
nor UO_179 (O_179,N_2954,N_2964);
or UO_180 (O_180,N_2968,N_2997);
or UO_181 (O_181,N_2984,N_2996);
or UO_182 (O_182,N_2982,N_2988);
nor UO_183 (O_183,N_2981,N_2991);
nor UO_184 (O_184,N_2997,N_2984);
nor UO_185 (O_185,N_2950,N_2971);
and UO_186 (O_186,N_2959,N_2995);
nand UO_187 (O_187,N_2992,N_2969);
nor UO_188 (O_188,N_2999,N_2963);
or UO_189 (O_189,N_2966,N_2977);
or UO_190 (O_190,N_2960,N_2967);
nand UO_191 (O_191,N_2981,N_2988);
and UO_192 (O_192,N_2962,N_2986);
nand UO_193 (O_193,N_2999,N_2981);
nand UO_194 (O_194,N_2976,N_2952);
or UO_195 (O_195,N_2994,N_2975);
and UO_196 (O_196,N_2960,N_2976);
and UO_197 (O_197,N_2986,N_2961);
nor UO_198 (O_198,N_2955,N_2968);
or UO_199 (O_199,N_2997,N_2983);
and UO_200 (O_200,N_2975,N_2995);
nand UO_201 (O_201,N_2967,N_2984);
or UO_202 (O_202,N_2998,N_2980);
or UO_203 (O_203,N_2994,N_2983);
and UO_204 (O_204,N_2969,N_2974);
and UO_205 (O_205,N_2988,N_2990);
nand UO_206 (O_206,N_2998,N_2959);
nor UO_207 (O_207,N_2997,N_2990);
nor UO_208 (O_208,N_2976,N_2972);
and UO_209 (O_209,N_2980,N_2996);
nor UO_210 (O_210,N_2990,N_2962);
or UO_211 (O_211,N_2976,N_2989);
nor UO_212 (O_212,N_2979,N_2954);
nor UO_213 (O_213,N_2988,N_2970);
or UO_214 (O_214,N_2960,N_2998);
nand UO_215 (O_215,N_2996,N_2999);
or UO_216 (O_216,N_2950,N_2974);
nor UO_217 (O_217,N_2984,N_2952);
and UO_218 (O_218,N_2982,N_2964);
nor UO_219 (O_219,N_2970,N_2958);
nor UO_220 (O_220,N_2979,N_2986);
nor UO_221 (O_221,N_2951,N_2981);
nand UO_222 (O_222,N_2986,N_2958);
nor UO_223 (O_223,N_2966,N_2971);
nand UO_224 (O_224,N_2992,N_2950);
nand UO_225 (O_225,N_2957,N_2959);
and UO_226 (O_226,N_2960,N_2993);
or UO_227 (O_227,N_2977,N_2967);
nand UO_228 (O_228,N_2991,N_2973);
or UO_229 (O_229,N_2961,N_2958);
or UO_230 (O_230,N_2992,N_2999);
nand UO_231 (O_231,N_2971,N_2985);
and UO_232 (O_232,N_2965,N_2974);
nor UO_233 (O_233,N_2996,N_2967);
or UO_234 (O_234,N_2962,N_2994);
or UO_235 (O_235,N_2963,N_2976);
nor UO_236 (O_236,N_2977,N_2975);
and UO_237 (O_237,N_2956,N_2950);
nand UO_238 (O_238,N_2984,N_2968);
or UO_239 (O_239,N_2973,N_2963);
or UO_240 (O_240,N_2981,N_2950);
nand UO_241 (O_241,N_2984,N_2951);
or UO_242 (O_242,N_2958,N_2950);
and UO_243 (O_243,N_2988,N_2963);
and UO_244 (O_244,N_2989,N_2981);
nor UO_245 (O_245,N_2981,N_2971);
nand UO_246 (O_246,N_2992,N_2993);
nand UO_247 (O_247,N_2998,N_2982);
nor UO_248 (O_248,N_2976,N_2995);
and UO_249 (O_249,N_2980,N_2990);
or UO_250 (O_250,N_2955,N_2980);
xor UO_251 (O_251,N_2970,N_2993);
nor UO_252 (O_252,N_2968,N_2986);
nand UO_253 (O_253,N_2989,N_2955);
nor UO_254 (O_254,N_2961,N_2968);
nand UO_255 (O_255,N_2983,N_2986);
nand UO_256 (O_256,N_2973,N_2979);
nand UO_257 (O_257,N_2994,N_2963);
and UO_258 (O_258,N_2963,N_2950);
nor UO_259 (O_259,N_2970,N_2982);
and UO_260 (O_260,N_2950,N_2975);
nand UO_261 (O_261,N_2973,N_2999);
nand UO_262 (O_262,N_2983,N_2996);
xor UO_263 (O_263,N_2967,N_2956);
nor UO_264 (O_264,N_2971,N_2995);
nand UO_265 (O_265,N_2974,N_2992);
nor UO_266 (O_266,N_2980,N_2964);
or UO_267 (O_267,N_2981,N_2993);
nand UO_268 (O_268,N_2999,N_2989);
nor UO_269 (O_269,N_2989,N_2965);
or UO_270 (O_270,N_2986,N_2963);
nand UO_271 (O_271,N_2997,N_2985);
and UO_272 (O_272,N_2974,N_2958);
or UO_273 (O_273,N_2971,N_2965);
or UO_274 (O_274,N_2970,N_2985);
nand UO_275 (O_275,N_2969,N_2967);
or UO_276 (O_276,N_2991,N_2993);
and UO_277 (O_277,N_2978,N_2966);
or UO_278 (O_278,N_2981,N_2984);
and UO_279 (O_279,N_2974,N_2990);
and UO_280 (O_280,N_2957,N_2981);
nor UO_281 (O_281,N_2973,N_2987);
or UO_282 (O_282,N_2972,N_2995);
nor UO_283 (O_283,N_2972,N_2954);
nor UO_284 (O_284,N_2996,N_2978);
and UO_285 (O_285,N_2962,N_2960);
nand UO_286 (O_286,N_2991,N_2984);
and UO_287 (O_287,N_2983,N_2990);
and UO_288 (O_288,N_2979,N_2998);
and UO_289 (O_289,N_2960,N_2978);
or UO_290 (O_290,N_2996,N_2988);
nor UO_291 (O_291,N_2953,N_2984);
xnor UO_292 (O_292,N_2998,N_2954);
and UO_293 (O_293,N_2973,N_2964);
nor UO_294 (O_294,N_2981,N_2969);
and UO_295 (O_295,N_2955,N_2953);
nor UO_296 (O_296,N_2986,N_2978);
nand UO_297 (O_297,N_2992,N_2995);
nand UO_298 (O_298,N_2997,N_2970);
nand UO_299 (O_299,N_2966,N_2953);
nand UO_300 (O_300,N_2951,N_2975);
nand UO_301 (O_301,N_2969,N_2997);
nand UO_302 (O_302,N_2953,N_2952);
and UO_303 (O_303,N_2986,N_2960);
nand UO_304 (O_304,N_2994,N_2960);
nand UO_305 (O_305,N_2995,N_2979);
nor UO_306 (O_306,N_2972,N_2983);
or UO_307 (O_307,N_2984,N_2954);
xor UO_308 (O_308,N_2995,N_2987);
or UO_309 (O_309,N_2970,N_2960);
nor UO_310 (O_310,N_2971,N_2999);
nor UO_311 (O_311,N_2956,N_2987);
and UO_312 (O_312,N_2991,N_2997);
nand UO_313 (O_313,N_2964,N_2985);
nand UO_314 (O_314,N_2953,N_2987);
and UO_315 (O_315,N_2962,N_2966);
and UO_316 (O_316,N_2991,N_2956);
nor UO_317 (O_317,N_2987,N_2963);
and UO_318 (O_318,N_2958,N_2967);
and UO_319 (O_319,N_2956,N_2959);
and UO_320 (O_320,N_2953,N_2999);
nor UO_321 (O_321,N_2990,N_2951);
or UO_322 (O_322,N_2971,N_2955);
nor UO_323 (O_323,N_2994,N_2998);
nand UO_324 (O_324,N_2983,N_2954);
or UO_325 (O_325,N_2994,N_2990);
nor UO_326 (O_326,N_2993,N_2955);
nor UO_327 (O_327,N_2977,N_2997);
nand UO_328 (O_328,N_2979,N_2970);
or UO_329 (O_329,N_2986,N_2955);
nand UO_330 (O_330,N_2998,N_2961);
xnor UO_331 (O_331,N_2975,N_2985);
nand UO_332 (O_332,N_2952,N_2967);
xnor UO_333 (O_333,N_2973,N_2971);
and UO_334 (O_334,N_2972,N_2978);
and UO_335 (O_335,N_2962,N_2981);
or UO_336 (O_336,N_2971,N_2979);
nor UO_337 (O_337,N_2982,N_2969);
nor UO_338 (O_338,N_2964,N_2986);
nand UO_339 (O_339,N_2977,N_2976);
and UO_340 (O_340,N_2984,N_2969);
nand UO_341 (O_341,N_2956,N_2989);
nor UO_342 (O_342,N_2957,N_2985);
nor UO_343 (O_343,N_2954,N_2953);
and UO_344 (O_344,N_2989,N_2961);
nor UO_345 (O_345,N_2992,N_2952);
nor UO_346 (O_346,N_2959,N_2961);
nor UO_347 (O_347,N_2987,N_2982);
and UO_348 (O_348,N_2963,N_2981);
or UO_349 (O_349,N_2989,N_2962);
or UO_350 (O_350,N_2963,N_2996);
and UO_351 (O_351,N_2953,N_2986);
nor UO_352 (O_352,N_2998,N_2968);
nor UO_353 (O_353,N_2990,N_2964);
nand UO_354 (O_354,N_2988,N_2951);
nand UO_355 (O_355,N_2952,N_2960);
and UO_356 (O_356,N_2976,N_2961);
and UO_357 (O_357,N_2974,N_2987);
or UO_358 (O_358,N_2968,N_2969);
or UO_359 (O_359,N_2997,N_2965);
nand UO_360 (O_360,N_2971,N_2961);
xnor UO_361 (O_361,N_2981,N_2987);
nor UO_362 (O_362,N_2977,N_2984);
nand UO_363 (O_363,N_2954,N_2950);
or UO_364 (O_364,N_2978,N_2973);
and UO_365 (O_365,N_2999,N_2966);
and UO_366 (O_366,N_2967,N_2964);
or UO_367 (O_367,N_2956,N_2976);
and UO_368 (O_368,N_2974,N_2968);
nand UO_369 (O_369,N_2956,N_2965);
nand UO_370 (O_370,N_2996,N_2961);
nor UO_371 (O_371,N_2952,N_2999);
and UO_372 (O_372,N_2959,N_2994);
or UO_373 (O_373,N_2996,N_2995);
nor UO_374 (O_374,N_2954,N_2989);
nor UO_375 (O_375,N_2990,N_2966);
or UO_376 (O_376,N_2989,N_2988);
nand UO_377 (O_377,N_2995,N_2990);
nand UO_378 (O_378,N_2974,N_2955);
nand UO_379 (O_379,N_2965,N_2967);
nand UO_380 (O_380,N_2971,N_2984);
or UO_381 (O_381,N_2998,N_2964);
nand UO_382 (O_382,N_2954,N_2987);
or UO_383 (O_383,N_2988,N_2984);
or UO_384 (O_384,N_2961,N_2957);
nor UO_385 (O_385,N_2952,N_2982);
nand UO_386 (O_386,N_2959,N_2963);
nand UO_387 (O_387,N_2984,N_2978);
nor UO_388 (O_388,N_2963,N_2961);
nand UO_389 (O_389,N_2959,N_2983);
nor UO_390 (O_390,N_2997,N_2956);
nor UO_391 (O_391,N_2953,N_2989);
or UO_392 (O_392,N_2976,N_2991);
nor UO_393 (O_393,N_2983,N_2978);
nor UO_394 (O_394,N_2952,N_2961);
nand UO_395 (O_395,N_2952,N_2970);
and UO_396 (O_396,N_2980,N_2986);
and UO_397 (O_397,N_2993,N_2968);
nand UO_398 (O_398,N_2991,N_2962);
nand UO_399 (O_399,N_2974,N_2972);
nand UO_400 (O_400,N_2961,N_2982);
nor UO_401 (O_401,N_2997,N_2961);
nand UO_402 (O_402,N_2987,N_2977);
nand UO_403 (O_403,N_2964,N_2950);
nand UO_404 (O_404,N_2977,N_2958);
nor UO_405 (O_405,N_2999,N_2975);
nor UO_406 (O_406,N_2960,N_2980);
and UO_407 (O_407,N_2985,N_2961);
or UO_408 (O_408,N_2986,N_2992);
nor UO_409 (O_409,N_2952,N_2969);
nand UO_410 (O_410,N_2997,N_2999);
or UO_411 (O_411,N_2968,N_2966);
nor UO_412 (O_412,N_2994,N_2964);
nand UO_413 (O_413,N_2977,N_2955);
and UO_414 (O_414,N_2974,N_2966);
and UO_415 (O_415,N_2980,N_2995);
and UO_416 (O_416,N_2967,N_2966);
or UO_417 (O_417,N_2957,N_2971);
and UO_418 (O_418,N_2990,N_2998);
nand UO_419 (O_419,N_2994,N_2988);
nor UO_420 (O_420,N_2987,N_2967);
nor UO_421 (O_421,N_2990,N_2977);
xor UO_422 (O_422,N_2971,N_2954);
nand UO_423 (O_423,N_2984,N_2957);
nand UO_424 (O_424,N_2995,N_2978);
nand UO_425 (O_425,N_2988,N_2993);
nor UO_426 (O_426,N_2974,N_2962);
nand UO_427 (O_427,N_2970,N_2978);
or UO_428 (O_428,N_2957,N_2952);
nor UO_429 (O_429,N_2968,N_2983);
and UO_430 (O_430,N_2975,N_2973);
nand UO_431 (O_431,N_2978,N_2998);
nand UO_432 (O_432,N_2950,N_2955);
nand UO_433 (O_433,N_2956,N_2984);
or UO_434 (O_434,N_2973,N_2965);
or UO_435 (O_435,N_2975,N_2966);
or UO_436 (O_436,N_2956,N_2964);
nand UO_437 (O_437,N_2967,N_2983);
and UO_438 (O_438,N_2956,N_2996);
and UO_439 (O_439,N_2966,N_2969);
nand UO_440 (O_440,N_2979,N_2957);
or UO_441 (O_441,N_2977,N_2962);
and UO_442 (O_442,N_2990,N_2981);
or UO_443 (O_443,N_2992,N_2972);
and UO_444 (O_444,N_2966,N_2954);
nor UO_445 (O_445,N_2991,N_2983);
nand UO_446 (O_446,N_2956,N_2953);
nand UO_447 (O_447,N_2986,N_2965);
nor UO_448 (O_448,N_2969,N_2986);
and UO_449 (O_449,N_2993,N_2975);
or UO_450 (O_450,N_2973,N_2983);
nor UO_451 (O_451,N_2969,N_2965);
and UO_452 (O_452,N_2977,N_2974);
or UO_453 (O_453,N_2961,N_2969);
and UO_454 (O_454,N_2985,N_2966);
and UO_455 (O_455,N_2984,N_2970);
or UO_456 (O_456,N_2987,N_2990);
and UO_457 (O_457,N_2973,N_2988);
xor UO_458 (O_458,N_2989,N_2974);
nand UO_459 (O_459,N_2965,N_2955);
and UO_460 (O_460,N_2984,N_2963);
nand UO_461 (O_461,N_2959,N_2992);
nand UO_462 (O_462,N_2997,N_2986);
and UO_463 (O_463,N_2952,N_2959);
nand UO_464 (O_464,N_2970,N_2974);
xor UO_465 (O_465,N_2983,N_2979);
and UO_466 (O_466,N_2970,N_2986);
or UO_467 (O_467,N_2979,N_2952);
or UO_468 (O_468,N_2952,N_2986);
and UO_469 (O_469,N_2951,N_2963);
and UO_470 (O_470,N_2985,N_2959);
or UO_471 (O_471,N_2995,N_2973);
or UO_472 (O_472,N_2998,N_2985);
or UO_473 (O_473,N_2984,N_2961);
nand UO_474 (O_474,N_2979,N_2985);
or UO_475 (O_475,N_2982,N_2983);
nand UO_476 (O_476,N_2987,N_2951);
nand UO_477 (O_477,N_2985,N_2973);
nor UO_478 (O_478,N_2956,N_2978);
or UO_479 (O_479,N_2968,N_2957);
nand UO_480 (O_480,N_2995,N_2983);
or UO_481 (O_481,N_2960,N_2977);
and UO_482 (O_482,N_2955,N_2969);
nor UO_483 (O_483,N_2957,N_2975);
or UO_484 (O_484,N_2988,N_2979);
or UO_485 (O_485,N_2999,N_2985);
or UO_486 (O_486,N_2967,N_2968);
nor UO_487 (O_487,N_2985,N_2974);
and UO_488 (O_488,N_2957,N_2955);
nand UO_489 (O_489,N_2952,N_2994);
or UO_490 (O_490,N_2986,N_2977);
nor UO_491 (O_491,N_2974,N_2954);
and UO_492 (O_492,N_2988,N_2977);
and UO_493 (O_493,N_2976,N_2998);
and UO_494 (O_494,N_2978,N_2962);
nor UO_495 (O_495,N_2955,N_2984);
nor UO_496 (O_496,N_2978,N_2991);
xor UO_497 (O_497,N_2962,N_2984);
and UO_498 (O_498,N_2954,N_2970);
nand UO_499 (O_499,N_2965,N_2985);
endmodule