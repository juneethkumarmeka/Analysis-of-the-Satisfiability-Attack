module basic_500_3000_500_5_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_109,In_208);
nor U1 (N_1,In_418,In_363);
and U2 (N_2,In_341,In_125);
nor U3 (N_3,In_280,In_374);
and U4 (N_4,In_93,In_173);
nor U5 (N_5,In_314,In_259);
nor U6 (N_6,In_372,In_117);
xnor U7 (N_7,In_453,In_420);
nand U8 (N_8,In_142,In_178);
nand U9 (N_9,In_346,In_450);
nand U10 (N_10,In_229,In_486);
xnor U11 (N_11,In_238,In_277);
and U12 (N_12,In_114,In_237);
or U13 (N_13,In_215,In_218);
nand U14 (N_14,In_38,In_2);
nand U15 (N_15,In_386,In_56);
nor U16 (N_16,In_6,In_22);
xnor U17 (N_17,In_451,In_454);
or U18 (N_18,In_42,In_433);
xnor U19 (N_19,In_477,In_26);
nand U20 (N_20,In_211,In_65);
or U21 (N_21,In_74,In_312);
nor U22 (N_22,In_171,In_269);
and U23 (N_23,In_449,In_70);
and U24 (N_24,In_1,In_424);
nand U25 (N_25,In_223,In_20);
nor U26 (N_26,In_416,In_319);
nand U27 (N_27,In_204,In_321);
nand U28 (N_28,In_214,In_139);
or U29 (N_29,In_465,In_7);
and U30 (N_30,In_325,In_92);
or U31 (N_31,In_138,In_481);
nand U32 (N_32,In_193,In_87);
nor U33 (N_33,In_73,In_91);
and U34 (N_34,In_345,In_355);
xnor U35 (N_35,In_428,In_216);
nor U36 (N_36,In_60,In_313);
nor U37 (N_37,In_198,In_226);
and U38 (N_38,In_133,In_236);
and U39 (N_39,In_83,In_69);
or U40 (N_40,In_279,In_360);
nand U41 (N_41,In_164,In_52);
and U42 (N_42,In_232,In_63);
or U43 (N_43,In_28,In_258);
nand U44 (N_44,In_48,In_320);
xor U45 (N_45,In_268,In_482);
or U46 (N_46,In_468,In_409);
and U47 (N_47,In_108,In_163);
nand U48 (N_48,In_336,In_426);
nor U49 (N_49,In_86,In_414);
nand U50 (N_50,In_412,In_287);
nor U51 (N_51,In_227,In_396);
or U52 (N_52,In_288,In_122);
nor U53 (N_53,In_478,In_471);
or U54 (N_54,In_407,In_489);
and U55 (N_55,In_398,In_121);
and U56 (N_56,In_435,In_202);
nand U57 (N_57,In_473,In_191);
nand U58 (N_58,In_281,In_487);
nand U59 (N_59,In_493,In_188);
and U60 (N_60,In_431,In_421);
nor U61 (N_61,In_290,In_298);
nor U62 (N_62,In_67,In_434);
nor U63 (N_63,In_102,In_131);
nor U64 (N_64,In_350,In_79);
nor U65 (N_65,In_463,In_490);
nor U66 (N_66,In_152,In_101);
or U67 (N_67,In_370,In_353);
nand U68 (N_68,In_221,In_359);
and U69 (N_69,In_495,In_395);
and U70 (N_70,In_408,In_172);
nor U71 (N_71,In_301,In_305);
or U72 (N_72,In_252,In_273);
nor U73 (N_73,In_385,In_242);
nand U74 (N_74,In_240,In_246);
and U75 (N_75,In_187,In_456);
or U76 (N_76,In_75,In_103);
or U77 (N_77,In_306,In_464);
nand U78 (N_78,In_417,In_41);
nor U79 (N_79,In_224,In_383);
nand U80 (N_80,In_123,In_285);
nor U81 (N_81,In_339,In_207);
nor U82 (N_82,In_179,In_194);
nand U83 (N_83,In_496,In_272);
nand U84 (N_84,In_439,In_254);
xnor U85 (N_85,In_12,In_82);
nand U86 (N_86,In_352,In_241);
and U87 (N_87,In_452,In_61);
nand U88 (N_88,In_327,In_384);
nand U89 (N_89,In_64,In_243);
nand U90 (N_90,In_497,In_154);
and U91 (N_91,In_53,In_54);
or U92 (N_92,In_366,In_239);
or U93 (N_93,In_380,In_120);
nand U94 (N_94,In_334,In_399);
nand U95 (N_95,In_441,In_488);
nand U96 (N_96,In_335,In_257);
xnor U97 (N_97,In_78,In_310);
and U98 (N_98,In_50,In_161);
or U99 (N_99,In_442,In_222);
or U100 (N_100,In_181,In_177);
or U101 (N_101,In_40,In_157);
nor U102 (N_102,In_403,In_84);
and U103 (N_103,In_467,In_205);
or U104 (N_104,In_19,In_419);
nor U105 (N_105,In_112,In_14);
and U106 (N_106,In_24,In_391);
nor U107 (N_107,In_499,In_309);
nor U108 (N_108,In_302,In_381);
nor U109 (N_109,In_199,In_357);
nand U110 (N_110,In_382,In_213);
nor U111 (N_111,In_183,In_485);
and U112 (N_112,In_343,In_361);
and U113 (N_113,In_21,In_104);
nand U114 (N_114,In_462,In_30);
and U115 (N_115,In_167,In_155);
or U116 (N_116,In_429,In_225);
nor U117 (N_117,In_349,In_255);
and U118 (N_118,In_127,In_480);
or U119 (N_119,In_51,In_295);
nor U120 (N_120,In_494,In_37);
nor U121 (N_121,In_264,In_168);
or U122 (N_122,In_315,In_176);
nand U123 (N_123,In_146,In_333);
nor U124 (N_124,In_230,In_362);
and U125 (N_125,In_351,In_15);
and U126 (N_126,In_27,In_220);
and U127 (N_127,In_106,In_99);
nand U128 (N_128,In_95,In_201);
nand U129 (N_129,In_265,In_143);
or U130 (N_130,In_76,In_77);
or U131 (N_131,In_356,In_165);
or U132 (N_132,In_260,In_251);
and U133 (N_133,In_136,In_389);
or U134 (N_134,In_44,In_141);
or U135 (N_135,In_270,In_43);
nand U136 (N_136,In_25,In_369);
nor U137 (N_137,In_10,In_189);
or U138 (N_138,In_250,In_184);
nor U139 (N_139,In_34,In_46);
nor U140 (N_140,In_322,In_85);
nand U141 (N_141,In_145,In_342);
or U142 (N_142,In_447,In_192);
and U143 (N_143,In_348,In_401);
or U144 (N_144,In_248,In_275);
nor U145 (N_145,In_308,In_159);
nand U146 (N_146,In_459,In_368);
and U147 (N_147,In_185,In_115);
and U148 (N_148,In_466,In_455);
xnor U149 (N_149,In_197,In_413);
nor U150 (N_150,In_387,In_16);
and U151 (N_151,In_234,In_11);
nand U152 (N_152,In_49,In_457);
or U153 (N_153,In_397,In_150);
or U154 (N_154,In_423,In_90);
nand U155 (N_155,In_303,In_347);
nor U156 (N_156,In_58,In_261);
nor U157 (N_157,In_94,In_461);
nor U158 (N_158,In_17,In_323);
nand U159 (N_159,In_492,In_406);
and U160 (N_160,In_97,In_375);
and U161 (N_161,In_262,In_330);
nor U162 (N_162,In_276,In_151);
nand U163 (N_163,In_256,In_3);
and U164 (N_164,In_200,In_317);
nor U165 (N_165,In_166,In_98);
and U166 (N_166,In_328,In_444);
nor U167 (N_167,In_411,In_116);
nand U168 (N_168,In_289,In_235);
and U169 (N_169,In_284,In_118);
nand U170 (N_170,In_68,In_231);
or U171 (N_171,In_160,In_66);
or U172 (N_172,In_458,In_460);
nand U173 (N_173,In_175,In_286);
nand U174 (N_174,In_324,In_124);
and U175 (N_175,In_81,In_5);
nor U176 (N_176,In_344,In_0);
or U177 (N_177,In_100,In_358);
and U178 (N_178,In_402,In_267);
or U179 (N_179,In_140,In_186);
nor U180 (N_180,In_249,In_217);
nand U181 (N_181,In_195,In_296);
or U182 (N_182,In_32,In_326);
or U183 (N_183,In_437,In_89);
nand U184 (N_184,In_329,In_293);
nand U185 (N_185,In_206,In_47);
nor U186 (N_186,In_432,In_233);
nor U187 (N_187,In_110,In_427);
and U188 (N_188,In_271,In_316);
and U189 (N_189,In_491,In_162);
nand U190 (N_190,In_113,In_170);
nand U191 (N_191,In_470,In_144);
or U192 (N_192,In_445,In_88);
nand U193 (N_193,In_158,In_156);
nand U194 (N_194,In_394,In_469);
nand U195 (N_195,In_404,In_210);
and U196 (N_196,In_476,In_291);
xnor U197 (N_197,In_62,In_283);
or U198 (N_198,In_196,In_57);
or U199 (N_199,In_134,In_180);
and U200 (N_200,In_130,In_245);
and U201 (N_201,In_297,In_148);
nand U202 (N_202,In_436,In_484);
or U203 (N_203,In_174,In_483);
and U204 (N_204,In_209,In_149);
and U205 (N_205,In_55,In_263);
or U206 (N_206,In_96,In_425);
nand U207 (N_207,In_137,In_266);
or U208 (N_208,In_311,In_9);
or U209 (N_209,In_182,In_247);
nor U210 (N_210,In_80,In_244);
nand U211 (N_211,In_365,In_318);
nor U212 (N_212,In_274,In_364);
nor U213 (N_213,In_107,In_390);
and U214 (N_214,In_111,In_190);
or U215 (N_215,In_18,In_400);
or U216 (N_216,In_39,In_446);
nand U217 (N_217,In_371,In_338);
nor U218 (N_218,In_367,In_438);
nor U219 (N_219,In_72,In_23);
or U220 (N_220,In_373,In_128);
nand U221 (N_221,In_392,In_299);
nand U222 (N_222,In_29,In_212);
nand U223 (N_223,In_36,In_35);
or U224 (N_224,In_475,In_410);
nor U225 (N_225,In_282,In_498);
and U226 (N_226,In_332,In_4);
nand U227 (N_227,In_31,In_203);
xor U228 (N_228,In_430,In_119);
or U229 (N_229,In_129,In_169);
nand U230 (N_230,In_304,In_479);
and U231 (N_231,In_405,In_422);
xnor U232 (N_232,In_219,In_378);
nor U233 (N_233,In_415,In_105);
nor U234 (N_234,In_448,In_8);
nand U235 (N_235,In_376,In_379);
nor U236 (N_236,In_294,In_71);
nor U237 (N_237,In_135,In_153);
nand U238 (N_238,In_126,In_354);
or U239 (N_239,In_59,In_393);
xnor U240 (N_240,In_278,In_331);
or U241 (N_241,In_132,In_45);
nor U242 (N_242,In_340,In_253);
or U243 (N_243,In_474,In_472);
nor U244 (N_244,In_443,In_33);
or U245 (N_245,In_337,In_388);
or U246 (N_246,In_377,In_228);
nor U247 (N_247,In_13,In_147);
nand U248 (N_248,In_300,In_292);
nand U249 (N_249,In_307,In_440);
and U250 (N_250,In_398,In_381);
nor U251 (N_251,In_383,In_381);
nand U252 (N_252,In_301,In_151);
nand U253 (N_253,In_148,In_48);
and U254 (N_254,In_279,In_438);
nand U255 (N_255,In_313,In_471);
nor U256 (N_256,In_77,In_118);
nor U257 (N_257,In_255,In_82);
or U258 (N_258,In_377,In_472);
nand U259 (N_259,In_331,In_342);
and U260 (N_260,In_28,In_330);
and U261 (N_261,In_112,In_5);
or U262 (N_262,In_440,In_161);
nor U263 (N_263,In_337,In_492);
nor U264 (N_264,In_97,In_493);
nor U265 (N_265,In_473,In_303);
or U266 (N_266,In_173,In_349);
xnor U267 (N_267,In_320,In_309);
nor U268 (N_268,In_391,In_85);
nor U269 (N_269,In_407,In_145);
nand U270 (N_270,In_371,In_204);
or U271 (N_271,In_320,In_399);
and U272 (N_272,In_420,In_296);
nand U273 (N_273,In_66,In_346);
nor U274 (N_274,In_288,In_192);
nor U275 (N_275,In_94,In_90);
nor U276 (N_276,In_140,In_478);
nand U277 (N_277,In_131,In_120);
nand U278 (N_278,In_472,In_365);
nor U279 (N_279,In_456,In_458);
nor U280 (N_280,In_375,In_244);
or U281 (N_281,In_399,In_341);
nor U282 (N_282,In_483,In_93);
and U283 (N_283,In_108,In_6);
and U284 (N_284,In_27,In_364);
xnor U285 (N_285,In_84,In_250);
nand U286 (N_286,In_194,In_36);
nor U287 (N_287,In_46,In_388);
nor U288 (N_288,In_432,In_197);
or U289 (N_289,In_313,In_437);
or U290 (N_290,In_137,In_8);
and U291 (N_291,In_420,In_150);
and U292 (N_292,In_216,In_320);
and U293 (N_293,In_162,In_476);
and U294 (N_294,In_156,In_237);
nand U295 (N_295,In_498,In_93);
or U296 (N_296,In_101,In_283);
nor U297 (N_297,In_286,In_7);
nand U298 (N_298,In_462,In_116);
nand U299 (N_299,In_229,In_116);
and U300 (N_300,In_389,In_400);
or U301 (N_301,In_340,In_329);
nor U302 (N_302,In_28,In_103);
nand U303 (N_303,In_93,In_228);
nand U304 (N_304,In_375,In_29);
nand U305 (N_305,In_138,In_296);
and U306 (N_306,In_299,In_24);
and U307 (N_307,In_312,In_157);
and U308 (N_308,In_151,In_220);
nand U309 (N_309,In_438,In_90);
and U310 (N_310,In_162,In_168);
and U311 (N_311,In_383,In_432);
nand U312 (N_312,In_100,In_259);
and U313 (N_313,In_8,In_174);
and U314 (N_314,In_39,In_407);
or U315 (N_315,In_152,In_413);
nand U316 (N_316,In_6,In_261);
and U317 (N_317,In_371,In_220);
nor U318 (N_318,In_225,In_425);
and U319 (N_319,In_28,In_192);
xor U320 (N_320,In_213,In_494);
nand U321 (N_321,In_198,In_330);
or U322 (N_322,In_354,In_414);
nand U323 (N_323,In_454,In_461);
nand U324 (N_324,In_108,In_294);
and U325 (N_325,In_358,In_118);
or U326 (N_326,In_330,In_123);
nor U327 (N_327,In_155,In_356);
nor U328 (N_328,In_493,In_233);
nand U329 (N_329,In_361,In_395);
nor U330 (N_330,In_50,In_181);
nand U331 (N_331,In_256,In_398);
nor U332 (N_332,In_258,In_15);
nand U333 (N_333,In_493,In_313);
and U334 (N_334,In_145,In_174);
and U335 (N_335,In_398,In_353);
and U336 (N_336,In_126,In_362);
or U337 (N_337,In_427,In_216);
and U338 (N_338,In_158,In_390);
nor U339 (N_339,In_425,In_367);
and U340 (N_340,In_16,In_250);
and U341 (N_341,In_334,In_172);
or U342 (N_342,In_168,In_87);
and U343 (N_343,In_83,In_385);
nor U344 (N_344,In_194,In_267);
and U345 (N_345,In_460,In_130);
and U346 (N_346,In_367,In_423);
or U347 (N_347,In_493,In_24);
or U348 (N_348,In_88,In_387);
xnor U349 (N_349,In_428,In_340);
or U350 (N_350,In_327,In_400);
nand U351 (N_351,In_337,In_392);
or U352 (N_352,In_68,In_113);
or U353 (N_353,In_406,In_204);
and U354 (N_354,In_70,In_415);
nor U355 (N_355,In_126,In_10);
and U356 (N_356,In_157,In_418);
and U357 (N_357,In_188,In_319);
xnor U358 (N_358,In_483,In_38);
and U359 (N_359,In_159,In_494);
nor U360 (N_360,In_310,In_0);
nand U361 (N_361,In_34,In_274);
or U362 (N_362,In_268,In_13);
and U363 (N_363,In_92,In_423);
nor U364 (N_364,In_21,In_150);
or U365 (N_365,In_133,In_245);
and U366 (N_366,In_277,In_78);
nand U367 (N_367,In_318,In_266);
nand U368 (N_368,In_275,In_117);
nand U369 (N_369,In_178,In_459);
nor U370 (N_370,In_369,In_200);
or U371 (N_371,In_113,In_356);
nand U372 (N_372,In_233,In_389);
nor U373 (N_373,In_483,In_338);
nor U374 (N_374,In_89,In_301);
and U375 (N_375,In_91,In_100);
and U376 (N_376,In_120,In_270);
and U377 (N_377,In_130,In_468);
nor U378 (N_378,In_13,In_207);
and U379 (N_379,In_315,In_244);
nand U380 (N_380,In_295,In_468);
and U381 (N_381,In_333,In_457);
nor U382 (N_382,In_154,In_190);
nand U383 (N_383,In_180,In_57);
or U384 (N_384,In_25,In_172);
or U385 (N_385,In_441,In_282);
and U386 (N_386,In_164,In_27);
nand U387 (N_387,In_311,In_297);
and U388 (N_388,In_29,In_273);
nor U389 (N_389,In_346,In_446);
or U390 (N_390,In_135,In_186);
or U391 (N_391,In_342,In_52);
nor U392 (N_392,In_246,In_374);
nor U393 (N_393,In_213,In_61);
and U394 (N_394,In_1,In_73);
nor U395 (N_395,In_226,In_376);
and U396 (N_396,In_289,In_198);
or U397 (N_397,In_454,In_208);
nor U398 (N_398,In_155,In_203);
nor U399 (N_399,In_211,In_130);
or U400 (N_400,In_286,In_14);
nand U401 (N_401,In_370,In_364);
and U402 (N_402,In_88,In_81);
and U403 (N_403,In_360,In_337);
nor U404 (N_404,In_445,In_219);
and U405 (N_405,In_152,In_203);
nor U406 (N_406,In_25,In_118);
and U407 (N_407,In_412,In_145);
nor U408 (N_408,In_67,In_379);
and U409 (N_409,In_35,In_257);
or U410 (N_410,In_361,In_30);
nand U411 (N_411,In_226,In_359);
or U412 (N_412,In_463,In_478);
or U413 (N_413,In_136,In_43);
nand U414 (N_414,In_345,In_378);
or U415 (N_415,In_480,In_400);
and U416 (N_416,In_30,In_144);
or U417 (N_417,In_216,In_389);
nor U418 (N_418,In_30,In_229);
nand U419 (N_419,In_108,In_461);
or U420 (N_420,In_234,In_17);
nor U421 (N_421,In_218,In_312);
and U422 (N_422,In_12,In_21);
xor U423 (N_423,In_170,In_144);
or U424 (N_424,In_198,In_458);
nand U425 (N_425,In_456,In_38);
nand U426 (N_426,In_265,In_297);
nand U427 (N_427,In_283,In_272);
nand U428 (N_428,In_492,In_316);
nor U429 (N_429,In_104,In_310);
or U430 (N_430,In_27,In_352);
nor U431 (N_431,In_293,In_235);
nand U432 (N_432,In_333,In_45);
and U433 (N_433,In_400,In_267);
and U434 (N_434,In_243,In_188);
nor U435 (N_435,In_136,In_332);
or U436 (N_436,In_160,In_76);
nand U437 (N_437,In_79,In_439);
nand U438 (N_438,In_287,In_233);
nor U439 (N_439,In_286,In_454);
nor U440 (N_440,In_338,In_181);
and U441 (N_441,In_141,In_232);
and U442 (N_442,In_344,In_245);
or U443 (N_443,In_484,In_399);
nand U444 (N_444,In_422,In_342);
and U445 (N_445,In_85,In_46);
or U446 (N_446,In_247,In_361);
or U447 (N_447,In_247,In_457);
nor U448 (N_448,In_436,In_487);
and U449 (N_449,In_469,In_325);
or U450 (N_450,In_397,In_100);
nor U451 (N_451,In_350,In_97);
nand U452 (N_452,In_136,In_393);
nor U453 (N_453,In_485,In_1);
or U454 (N_454,In_474,In_453);
nand U455 (N_455,In_338,In_159);
nor U456 (N_456,In_413,In_83);
nand U457 (N_457,In_185,In_81);
nand U458 (N_458,In_152,In_19);
and U459 (N_459,In_290,In_173);
and U460 (N_460,In_428,In_227);
nand U461 (N_461,In_230,In_62);
nand U462 (N_462,In_401,In_23);
nor U463 (N_463,In_92,In_6);
nand U464 (N_464,In_227,In_363);
and U465 (N_465,In_82,In_5);
and U466 (N_466,In_332,In_264);
nand U467 (N_467,In_440,In_408);
or U468 (N_468,In_398,In_102);
xnor U469 (N_469,In_203,In_313);
nor U470 (N_470,In_321,In_486);
or U471 (N_471,In_212,In_407);
nor U472 (N_472,In_172,In_267);
xor U473 (N_473,In_102,In_347);
nand U474 (N_474,In_266,In_264);
or U475 (N_475,In_344,In_55);
and U476 (N_476,In_473,In_171);
nor U477 (N_477,In_33,In_146);
nand U478 (N_478,In_25,In_348);
or U479 (N_479,In_248,In_257);
and U480 (N_480,In_275,In_41);
xor U481 (N_481,In_428,In_465);
nand U482 (N_482,In_437,In_343);
and U483 (N_483,In_313,In_490);
and U484 (N_484,In_430,In_448);
or U485 (N_485,In_149,In_263);
and U486 (N_486,In_296,In_95);
nand U487 (N_487,In_184,In_199);
or U488 (N_488,In_309,In_489);
or U489 (N_489,In_127,In_347);
or U490 (N_490,In_109,In_227);
nor U491 (N_491,In_356,In_439);
nor U492 (N_492,In_23,In_213);
xnor U493 (N_493,In_33,In_332);
nor U494 (N_494,In_48,In_497);
xor U495 (N_495,In_0,In_476);
nand U496 (N_496,In_469,In_267);
nor U497 (N_497,In_396,In_416);
xnor U498 (N_498,In_432,In_484);
or U499 (N_499,In_33,In_204);
nor U500 (N_500,In_430,In_471);
and U501 (N_501,In_338,In_319);
nand U502 (N_502,In_411,In_199);
or U503 (N_503,In_466,In_82);
nor U504 (N_504,In_302,In_109);
nand U505 (N_505,In_118,In_326);
or U506 (N_506,In_120,In_253);
and U507 (N_507,In_60,In_273);
nor U508 (N_508,In_292,In_351);
and U509 (N_509,In_166,In_24);
or U510 (N_510,In_436,In_267);
nand U511 (N_511,In_321,In_23);
nand U512 (N_512,In_69,In_95);
and U513 (N_513,In_259,In_481);
and U514 (N_514,In_187,In_11);
nor U515 (N_515,In_285,In_280);
nand U516 (N_516,In_219,In_279);
nor U517 (N_517,In_70,In_6);
and U518 (N_518,In_97,In_28);
nand U519 (N_519,In_478,In_28);
and U520 (N_520,In_386,In_282);
and U521 (N_521,In_94,In_11);
and U522 (N_522,In_17,In_254);
nor U523 (N_523,In_258,In_493);
nor U524 (N_524,In_367,In_427);
or U525 (N_525,In_156,In_42);
nor U526 (N_526,In_114,In_251);
or U527 (N_527,In_328,In_235);
and U528 (N_528,In_145,In_14);
or U529 (N_529,In_382,In_284);
or U530 (N_530,In_148,In_432);
or U531 (N_531,In_14,In_380);
or U532 (N_532,In_52,In_475);
nor U533 (N_533,In_416,In_385);
and U534 (N_534,In_474,In_19);
nand U535 (N_535,In_286,In_292);
or U536 (N_536,In_189,In_365);
nor U537 (N_537,In_66,In_310);
or U538 (N_538,In_442,In_301);
or U539 (N_539,In_77,In_452);
nor U540 (N_540,In_469,In_387);
and U541 (N_541,In_17,In_21);
nor U542 (N_542,In_102,In_133);
nor U543 (N_543,In_44,In_226);
nand U544 (N_544,In_492,In_475);
and U545 (N_545,In_172,In_412);
or U546 (N_546,In_77,In_63);
xor U547 (N_547,In_161,In_369);
or U548 (N_548,In_295,In_88);
or U549 (N_549,In_67,In_391);
nand U550 (N_550,In_198,In_294);
nor U551 (N_551,In_451,In_221);
nor U552 (N_552,In_307,In_387);
or U553 (N_553,In_315,In_338);
or U554 (N_554,In_346,In_200);
nand U555 (N_555,In_269,In_311);
nand U556 (N_556,In_388,In_36);
and U557 (N_557,In_444,In_268);
or U558 (N_558,In_239,In_393);
nand U559 (N_559,In_109,In_198);
nor U560 (N_560,In_444,In_352);
nand U561 (N_561,In_441,In_2);
nor U562 (N_562,In_28,In_353);
and U563 (N_563,In_213,In_100);
and U564 (N_564,In_358,In_281);
or U565 (N_565,In_381,In_438);
or U566 (N_566,In_234,In_358);
and U567 (N_567,In_187,In_215);
and U568 (N_568,In_194,In_23);
and U569 (N_569,In_359,In_461);
and U570 (N_570,In_480,In_499);
or U571 (N_571,In_80,In_412);
and U572 (N_572,In_410,In_22);
nor U573 (N_573,In_77,In_257);
nand U574 (N_574,In_86,In_244);
nand U575 (N_575,In_185,In_447);
or U576 (N_576,In_265,In_122);
or U577 (N_577,In_198,In_422);
and U578 (N_578,In_284,In_398);
nand U579 (N_579,In_96,In_108);
nor U580 (N_580,In_64,In_429);
and U581 (N_581,In_28,In_177);
and U582 (N_582,In_108,In_368);
and U583 (N_583,In_249,In_273);
nand U584 (N_584,In_52,In_467);
nand U585 (N_585,In_3,In_386);
nor U586 (N_586,In_144,In_296);
and U587 (N_587,In_285,In_377);
or U588 (N_588,In_489,In_244);
or U589 (N_589,In_473,In_401);
and U590 (N_590,In_434,In_347);
or U591 (N_591,In_283,In_54);
nor U592 (N_592,In_291,In_364);
nor U593 (N_593,In_406,In_111);
nand U594 (N_594,In_344,In_200);
and U595 (N_595,In_172,In_164);
and U596 (N_596,In_199,In_455);
and U597 (N_597,In_239,In_378);
nand U598 (N_598,In_350,In_284);
or U599 (N_599,In_284,In_157);
or U600 (N_600,N_124,N_442);
and U601 (N_601,N_317,N_375);
xor U602 (N_602,N_7,N_172);
or U603 (N_603,N_544,N_198);
or U604 (N_604,N_483,N_186);
or U605 (N_605,N_68,N_246);
or U606 (N_606,N_484,N_521);
nor U607 (N_607,N_540,N_518);
or U608 (N_608,N_423,N_162);
and U609 (N_609,N_86,N_188);
nand U610 (N_610,N_24,N_335);
nand U611 (N_611,N_531,N_383);
nor U612 (N_612,N_201,N_574);
and U613 (N_613,N_178,N_507);
nor U614 (N_614,N_353,N_42);
or U615 (N_615,N_242,N_181);
and U616 (N_616,N_366,N_318);
nand U617 (N_617,N_435,N_545);
nand U618 (N_618,N_1,N_476);
and U619 (N_619,N_529,N_412);
and U620 (N_620,N_490,N_347);
nor U621 (N_621,N_241,N_16);
nor U622 (N_622,N_33,N_527);
or U623 (N_623,N_314,N_326);
nor U624 (N_624,N_421,N_216);
nand U625 (N_625,N_313,N_520);
nor U626 (N_626,N_228,N_420);
and U627 (N_627,N_297,N_323);
or U628 (N_628,N_495,N_104);
or U629 (N_629,N_582,N_332);
and U630 (N_630,N_4,N_372);
or U631 (N_631,N_103,N_199);
nor U632 (N_632,N_105,N_530);
and U633 (N_633,N_194,N_338);
nor U634 (N_634,N_248,N_143);
and U635 (N_635,N_398,N_340);
or U636 (N_636,N_163,N_380);
nand U637 (N_637,N_66,N_191);
nand U638 (N_638,N_404,N_283);
nand U639 (N_639,N_496,N_35);
or U640 (N_640,N_559,N_110);
nor U641 (N_641,N_570,N_126);
nor U642 (N_642,N_477,N_171);
or U643 (N_643,N_277,N_400);
or U644 (N_644,N_355,N_387);
nand U645 (N_645,N_217,N_377);
or U646 (N_646,N_38,N_526);
nor U647 (N_647,N_367,N_593);
nor U648 (N_648,N_436,N_14);
or U649 (N_649,N_364,N_352);
nor U650 (N_650,N_385,N_28);
nor U651 (N_651,N_243,N_362);
nor U652 (N_652,N_500,N_413);
nor U653 (N_653,N_206,N_63);
nand U654 (N_654,N_179,N_461);
nand U655 (N_655,N_99,N_374);
and U656 (N_656,N_272,N_575);
nand U657 (N_657,N_341,N_46);
nor U658 (N_658,N_184,N_113);
nor U659 (N_659,N_269,N_43);
or U660 (N_660,N_11,N_254);
or U661 (N_661,N_2,N_312);
nor U662 (N_662,N_503,N_293);
and U663 (N_663,N_137,N_93);
or U664 (N_664,N_357,N_263);
or U665 (N_665,N_433,N_8);
or U666 (N_666,N_96,N_345);
nand U667 (N_667,N_21,N_169);
nand U668 (N_668,N_252,N_295);
nor U669 (N_669,N_480,N_514);
and U670 (N_670,N_118,N_462);
nor U671 (N_671,N_108,N_552);
or U672 (N_672,N_543,N_549);
nor U673 (N_673,N_557,N_90);
or U674 (N_674,N_239,N_139);
and U675 (N_675,N_13,N_394);
nand U676 (N_676,N_273,N_571);
nand U677 (N_677,N_210,N_251);
nor U678 (N_678,N_53,N_233);
nor U679 (N_679,N_390,N_524);
and U680 (N_680,N_258,N_359);
or U681 (N_681,N_382,N_379);
nor U682 (N_682,N_300,N_418);
and U683 (N_683,N_197,N_454);
and U684 (N_684,N_510,N_158);
nand U685 (N_685,N_261,N_114);
or U686 (N_686,N_222,N_81);
or U687 (N_687,N_26,N_146);
nor U688 (N_688,N_384,N_342);
xnor U689 (N_689,N_350,N_465);
and U690 (N_690,N_505,N_72);
or U691 (N_691,N_112,N_185);
or U692 (N_692,N_537,N_441);
xor U693 (N_693,N_55,N_349);
xnor U694 (N_694,N_591,N_472);
nor U695 (N_695,N_174,N_266);
or U696 (N_696,N_419,N_513);
or U697 (N_697,N_170,N_502);
nand U698 (N_698,N_31,N_9);
or U699 (N_699,N_488,N_506);
or U700 (N_700,N_159,N_393);
and U701 (N_701,N_523,N_459);
and U702 (N_702,N_265,N_29);
and U703 (N_703,N_406,N_361);
and U704 (N_704,N_528,N_561);
nor U705 (N_705,N_234,N_44);
nor U706 (N_706,N_147,N_79);
nor U707 (N_707,N_17,N_123);
or U708 (N_708,N_539,N_597);
or U709 (N_709,N_111,N_84);
nor U710 (N_710,N_65,N_449);
and U711 (N_711,N_89,N_152);
and U712 (N_712,N_80,N_471);
and U713 (N_713,N_280,N_94);
xor U714 (N_714,N_386,N_583);
nand U715 (N_715,N_535,N_221);
and U716 (N_716,N_565,N_27);
or U717 (N_717,N_148,N_240);
or U718 (N_718,N_532,N_52);
or U719 (N_719,N_308,N_450);
nor U720 (N_720,N_223,N_20);
nand U721 (N_721,N_285,N_207);
nand U722 (N_722,N_426,N_294);
or U723 (N_723,N_492,N_373);
or U724 (N_724,N_316,N_401);
and U725 (N_725,N_284,N_101);
nor U726 (N_726,N_3,N_85);
nand U727 (N_727,N_566,N_204);
and U728 (N_728,N_303,N_125);
nor U729 (N_729,N_439,N_363);
xor U730 (N_730,N_381,N_235);
and U731 (N_731,N_516,N_10);
and U732 (N_732,N_253,N_180);
nor U733 (N_733,N_209,N_551);
or U734 (N_734,N_424,N_276);
or U735 (N_735,N_573,N_219);
nor U736 (N_736,N_224,N_167);
nor U737 (N_737,N_213,N_60);
nand U738 (N_738,N_238,N_329);
or U739 (N_739,N_183,N_227);
and U740 (N_740,N_208,N_30);
and U741 (N_741,N_346,N_37);
nand U742 (N_742,N_493,N_331);
or U743 (N_743,N_376,N_156);
and U744 (N_744,N_304,N_91);
and U745 (N_745,N_494,N_431);
nor U746 (N_746,N_195,N_555);
xnor U747 (N_747,N_250,N_414);
and U748 (N_748,N_149,N_212);
nand U749 (N_749,N_173,N_120);
and U750 (N_750,N_556,N_411);
nand U751 (N_751,N_75,N_460);
or U752 (N_752,N_330,N_554);
nand U753 (N_753,N_517,N_368);
and U754 (N_754,N_469,N_452);
nor U755 (N_755,N_370,N_260);
and U756 (N_756,N_579,N_324);
or U757 (N_757,N_515,N_572);
nand U758 (N_758,N_508,N_344);
nor U759 (N_759,N_562,N_278);
and U760 (N_760,N_290,N_215);
nor U761 (N_761,N_56,N_161);
nand U762 (N_762,N_481,N_533);
nor U763 (N_763,N_407,N_425);
and U764 (N_764,N_391,N_0);
nor U765 (N_765,N_339,N_422);
nand U766 (N_766,N_82,N_164);
nand U767 (N_767,N_291,N_47);
or U768 (N_768,N_232,N_356);
or U769 (N_769,N_15,N_457);
nor U770 (N_770,N_512,N_130);
or U771 (N_771,N_98,N_226);
nor U772 (N_772,N_117,N_131);
or U773 (N_773,N_74,N_32);
and U774 (N_774,N_542,N_586);
xor U775 (N_775,N_354,N_585);
nor U776 (N_776,N_129,N_497);
nand U777 (N_777,N_546,N_41);
nand U778 (N_778,N_87,N_595);
nor U779 (N_779,N_189,N_203);
nand U780 (N_780,N_102,N_133);
nand U781 (N_781,N_548,N_564);
nand U782 (N_782,N_190,N_321);
and U783 (N_783,N_154,N_54);
nand U784 (N_784,N_62,N_358);
and U785 (N_785,N_473,N_150);
and U786 (N_786,N_444,N_417);
xnor U787 (N_787,N_220,N_351);
nor U788 (N_788,N_64,N_145);
nand U789 (N_789,N_218,N_447);
nand U790 (N_790,N_311,N_519);
nand U791 (N_791,N_175,N_140);
or U792 (N_792,N_399,N_187);
and U793 (N_793,N_51,N_282);
and U794 (N_794,N_588,N_470);
nand U795 (N_795,N_270,N_109);
nor U796 (N_796,N_408,N_153);
nand U797 (N_797,N_580,N_305);
nand U798 (N_798,N_67,N_231);
nor U799 (N_799,N_100,N_416);
nor U800 (N_800,N_36,N_327);
nand U801 (N_801,N_596,N_88);
or U802 (N_802,N_491,N_205);
and U803 (N_803,N_19,N_486);
and U804 (N_804,N_39,N_77);
nor U805 (N_805,N_309,N_225);
or U806 (N_806,N_107,N_166);
nor U807 (N_807,N_409,N_236);
nand U808 (N_808,N_434,N_577);
nand U809 (N_809,N_534,N_71);
or U810 (N_810,N_334,N_360);
or U811 (N_811,N_83,N_443);
nand U812 (N_812,N_455,N_92);
nor U813 (N_813,N_440,N_45);
or U814 (N_814,N_135,N_287);
or U815 (N_815,N_589,N_501);
or U816 (N_816,N_581,N_498);
xnor U817 (N_817,N_511,N_116);
or U818 (N_818,N_333,N_49);
nand U819 (N_819,N_453,N_522);
or U820 (N_820,N_410,N_299);
xnor U821 (N_821,N_478,N_292);
or U822 (N_822,N_138,N_275);
and U823 (N_823,N_568,N_550);
and U824 (N_824,N_302,N_474);
nand U825 (N_825,N_467,N_428);
nor U826 (N_826,N_245,N_429);
and U827 (N_827,N_165,N_415);
and U828 (N_828,N_567,N_132);
or U829 (N_829,N_468,N_177);
nor U830 (N_830,N_525,N_151);
nor U831 (N_831,N_590,N_448);
nor U832 (N_832,N_463,N_6);
or U833 (N_833,N_237,N_563);
and U834 (N_834,N_247,N_430);
and U835 (N_835,N_259,N_97);
and U836 (N_836,N_504,N_487);
nor U837 (N_837,N_121,N_427);
nand U838 (N_838,N_50,N_115);
nand U839 (N_839,N_288,N_397);
or U840 (N_840,N_456,N_48);
xnor U841 (N_841,N_378,N_192);
nor U842 (N_842,N_509,N_451);
or U843 (N_843,N_59,N_279);
and U844 (N_844,N_298,N_594);
or U845 (N_845,N_211,N_395);
nand U846 (N_846,N_445,N_365);
nor U847 (N_847,N_319,N_23);
nand U848 (N_848,N_134,N_271);
nor U849 (N_849,N_182,N_466);
or U850 (N_850,N_122,N_446);
and U851 (N_851,N_144,N_403);
and U852 (N_852,N_22,N_482);
nand U853 (N_853,N_320,N_541);
nand U854 (N_854,N_34,N_155);
and U855 (N_855,N_599,N_229);
nor U856 (N_856,N_547,N_343);
nor U857 (N_857,N_202,N_587);
nand U858 (N_858,N_274,N_25);
and U859 (N_859,N_40,N_322);
nand U860 (N_860,N_286,N_244);
nor U861 (N_861,N_598,N_142);
nor U862 (N_862,N_200,N_306);
nand U863 (N_863,N_264,N_73);
and U864 (N_864,N_69,N_578);
nand U865 (N_865,N_475,N_12);
or U866 (N_866,N_262,N_257);
nand U867 (N_867,N_76,N_325);
nor U868 (N_868,N_5,N_119);
nand U869 (N_869,N_336,N_584);
nand U870 (N_870,N_405,N_18);
nand U871 (N_871,N_396,N_281);
nand U872 (N_872,N_538,N_157);
or U873 (N_873,N_289,N_348);
nor U874 (N_874,N_214,N_437);
nor U875 (N_875,N_307,N_489);
xnor U876 (N_876,N_301,N_310);
and U877 (N_877,N_536,N_553);
nor U878 (N_878,N_136,N_141);
nand U879 (N_879,N_371,N_255);
and U880 (N_880,N_558,N_256);
nor U881 (N_881,N_57,N_328);
or U882 (N_882,N_249,N_268);
nor U883 (N_883,N_369,N_176);
xor U884 (N_884,N_388,N_458);
nand U885 (N_885,N_78,N_230);
or U886 (N_886,N_432,N_389);
nor U887 (N_887,N_499,N_392);
nor U888 (N_888,N_127,N_479);
nand U889 (N_889,N_485,N_438);
nor U890 (N_890,N_296,N_592);
nor U891 (N_891,N_402,N_464);
nor U892 (N_892,N_196,N_576);
or U893 (N_893,N_193,N_106);
and U894 (N_894,N_95,N_569);
nand U895 (N_895,N_315,N_560);
nand U896 (N_896,N_128,N_61);
nor U897 (N_897,N_168,N_70);
and U898 (N_898,N_267,N_337);
nand U899 (N_899,N_58,N_160);
nand U900 (N_900,N_585,N_321);
and U901 (N_901,N_375,N_414);
and U902 (N_902,N_173,N_169);
nand U903 (N_903,N_126,N_121);
nor U904 (N_904,N_464,N_159);
or U905 (N_905,N_274,N_13);
and U906 (N_906,N_479,N_356);
and U907 (N_907,N_432,N_274);
or U908 (N_908,N_362,N_160);
nand U909 (N_909,N_549,N_207);
and U910 (N_910,N_528,N_136);
nand U911 (N_911,N_18,N_142);
nor U912 (N_912,N_208,N_16);
and U913 (N_913,N_68,N_595);
nand U914 (N_914,N_138,N_479);
nor U915 (N_915,N_183,N_95);
or U916 (N_916,N_510,N_587);
or U917 (N_917,N_68,N_96);
or U918 (N_918,N_337,N_77);
or U919 (N_919,N_337,N_27);
nor U920 (N_920,N_549,N_472);
nor U921 (N_921,N_197,N_344);
and U922 (N_922,N_70,N_5);
nor U923 (N_923,N_107,N_211);
nand U924 (N_924,N_233,N_459);
nor U925 (N_925,N_469,N_141);
xnor U926 (N_926,N_199,N_189);
or U927 (N_927,N_591,N_418);
or U928 (N_928,N_37,N_167);
or U929 (N_929,N_219,N_38);
nand U930 (N_930,N_252,N_376);
and U931 (N_931,N_92,N_355);
and U932 (N_932,N_195,N_6);
and U933 (N_933,N_378,N_371);
nand U934 (N_934,N_391,N_168);
nor U935 (N_935,N_216,N_486);
or U936 (N_936,N_351,N_411);
and U937 (N_937,N_523,N_157);
and U938 (N_938,N_479,N_36);
nand U939 (N_939,N_503,N_26);
nand U940 (N_940,N_316,N_37);
nand U941 (N_941,N_83,N_597);
or U942 (N_942,N_587,N_271);
nor U943 (N_943,N_289,N_440);
nor U944 (N_944,N_370,N_174);
nand U945 (N_945,N_598,N_322);
or U946 (N_946,N_10,N_177);
or U947 (N_947,N_29,N_371);
or U948 (N_948,N_307,N_370);
or U949 (N_949,N_258,N_364);
xnor U950 (N_950,N_56,N_174);
nor U951 (N_951,N_358,N_513);
and U952 (N_952,N_100,N_581);
nor U953 (N_953,N_254,N_192);
or U954 (N_954,N_45,N_39);
xor U955 (N_955,N_497,N_5);
nor U956 (N_956,N_289,N_568);
nor U957 (N_957,N_219,N_495);
and U958 (N_958,N_378,N_2);
nand U959 (N_959,N_269,N_387);
or U960 (N_960,N_536,N_568);
nor U961 (N_961,N_510,N_115);
or U962 (N_962,N_458,N_301);
or U963 (N_963,N_586,N_203);
nand U964 (N_964,N_215,N_55);
nand U965 (N_965,N_216,N_249);
or U966 (N_966,N_29,N_574);
nor U967 (N_967,N_384,N_505);
or U968 (N_968,N_470,N_18);
nor U969 (N_969,N_406,N_466);
or U970 (N_970,N_77,N_462);
nand U971 (N_971,N_215,N_552);
nor U972 (N_972,N_51,N_165);
nand U973 (N_973,N_69,N_214);
or U974 (N_974,N_336,N_408);
nand U975 (N_975,N_444,N_132);
nor U976 (N_976,N_87,N_356);
xnor U977 (N_977,N_245,N_390);
and U978 (N_978,N_248,N_519);
or U979 (N_979,N_231,N_236);
nor U980 (N_980,N_94,N_445);
nand U981 (N_981,N_509,N_7);
nand U982 (N_982,N_461,N_8);
or U983 (N_983,N_552,N_299);
and U984 (N_984,N_263,N_140);
nor U985 (N_985,N_454,N_40);
or U986 (N_986,N_88,N_265);
nand U987 (N_987,N_82,N_193);
or U988 (N_988,N_528,N_458);
and U989 (N_989,N_39,N_472);
nor U990 (N_990,N_106,N_382);
nor U991 (N_991,N_390,N_225);
nor U992 (N_992,N_528,N_396);
nor U993 (N_993,N_477,N_445);
nand U994 (N_994,N_522,N_66);
and U995 (N_995,N_580,N_283);
or U996 (N_996,N_554,N_528);
nor U997 (N_997,N_341,N_160);
or U998 (N_998,N_413,N_156);
or U999 (N_999,N_104,N_469);
nor U1000 (N_1000,N_282,N_52);
or U1001 (N_1001,N_101,N_405);
nand U1002 (N_1002,N_293,N_585);
nor U1003 (N_1003,N_320,N_123);
or U1004 (N_1004,N_66,N_89);
nand U1005 (N_1005,N_270,N_429);
nand U1006 (N_1006,N_340,N_293);
nand U1007 (N_1007,N_383,N_190);
nand U1008 (N_1008,N_98,N_221);
or U1009 (N_1009,N_133,N_515);
nor U1010 (N_1010,N_70,N_233);
or U1011 (N_1011,N_520,N_482);
nand U1012 (N_1012,N_244,N_201);
and U1013 (N_1013,N_452,N_269);
xnor U1014 (N_1014,N_254,N_370);
nor U1015 (N_1015,N_589,N_107);
nand U1016 (N_1016,N_409,N_557);
or U1017 (N_1017,N_464,N_104);
nor U1018 (N_1018,N_489,N_510);
and U1019 (N_1019,N_249,N_195);
nand U1020 (N_1020,N_190,N_275);
or U1021 (N_1021,N_239,N_198);
nand U1022 (N_1022,N_110,N_596);
nor U1023 (N_1023,N_476,N_291);
nor U1024 (N_1024,N_334,N_216);
nor U1025 (N_1025,N_225,N_211);
and U1026 (N_1026,N_57,N_198);
and U1027 (N_1027,N_267,N_190);
nand U1028 (N_1028,N_151,N_241);
or U1029 (N_1029,N_173,N_453);
nor U1030 (N_1030,N_394,N_225);
or U1031 (N_1031,N_69,N_428);
nor U1032 (N_1032,N_499,N_183);
and U1033 (N_1033,N_407,N_489);
nand U1034 (N_1034,N_325,N_537);
and U1035 (N_1035,N_257,N_151);
or U1036 (N_1036,N_410,N_405);
nor U1037 (N_1037,N_27,N_110);
or U1038 (N_1038,N_263,N_455);
and U1039 (N_1039,N_343,N_373);
nor U1040 (N_1040,N_574,N_193);
or U1041 (N_1041,N_320,N_212);
nor U1042 (N_1042,N_5,N_386);
nand U1043 (N_1043,N_433,N_256);
or U1044 (N_1044,N_227,N_409);
and U1045 (N_1045,N_410,N_94);
and U1046 (N_1046,N_264,N_410);
or U1047 (N_1047,N_544,N_545);
nor U1048 (N_1048,N_361,N_402);
and U1049 (N_1049,N_433,N_407);
nand U1050 (N_1050,N_271,N_411);
nor U1051 (N_1051,N_325,N_477);
or U1052 (N_1052,N_270,N_214);
nand U1053 (N_1053,N_131,N_520);
nand U1054 (N_1054,N_2,N_161);
nor U1055 (N_1055,N_597,N_428);
or U1056 (N_1056,N_481,N_595);
or U1057 (N_1057,N_90,N_381);
or U1058 (N_1058,N_387,N_491);
and U1059 (N_1059,N_438,N_395);
or U1060 (N_1060,N_286,N_195);
nand U1061 (N_1061,N_350,N_42);
or U1062 (N_1062,N_569,N_44);
nor U1063 (N_1063,N_70,N_258);
nand U1064 (N_1064,N_468,N_259);
or U1065 (N_1065,N_372,N_86);
or U1066 (N_1066,N_355,N_34);
nor U1067 (N_1067,N_477,N_237);
or U1068 (N_1068,N_345,N_559);
and U1069 (N_1069,N_221,N_475);
nand U1070 (N_1070,N_119,N_175);
nand U1071 (N_1071,N_480,N_497);
and U1072 (N_1072,N_513,N_141);
nand U1073 (N_1073,N_114,N_227);
nand U1074 (N_1074,N_387,N_542);
or U1075 (N_1075,N_427,N_76);
nand U1076 (N_1076,N_356,N_27);
and U1077 (N_1077,N_487,N_503);
nor U1078 (N_1078,N_562,N_57);
nand U1079 (N_1079,N_68,N_92);
nand U1080 (N_1080,N_425,N_157);
nor U1081 (N_1081,N_517,N_217);
nor U1082 (N_1082,N_181,N_313);
nor U1083 (N_1083,N_459,N_228);
nand U1084 (N_1084,N_576,N_308);
and U1085 (N_1085,N_222,N_414);
nand U1086 (N_1086,N_529,N_294);
or U1087 (N_1087,N_336,N_384);
nand U1088 (N_1088,N_382,N_401);
or U1089 (N_1089,N_175,N_438);
nor U1090 (N_1090,N_508,N_88);
and U1091 (N_1091,N_94,N_516);
nand U1092 (N_1092,N_218,N_339);
or U1093 (N_1093,N_545,N_90);
and U1094 (N_1094,N_598,N_468);
nor U1095 (N_1095,N_365,N_337);
nand U1096 (N_1096,N_146,N_51);
or U1097 (N_1097,N_498,N_37);
or U1098 (N_1098,N_138,N_317);
or U1099 (N_1099,N_394,N_194);
or U1100 (N_1100,N_271,N_261);
or U1101 (N_1101,N_314,N_527);
nor U1102 (N_1102,N_30,N_353);
or U1103 (N_1103,N_250,N_137);
nor U1104 (N_1104,N_98,N_26);
or U1105 (N_1105,N_183,N_164);
and U1106 (N_1106,N_539,N_373);
or U1107 (N_1107,N_258,N_230);
or U1108 (N_1108,N_369,N_44);
xor U1109 (N_1109,N_20,N_513);
nor U1110 (N_1110,N_429,N_431);
and U1111 (N_1111,N_153,N_196);
or U1112 (N_1112,N_131,N_4);
or U1113 (N_1113,N_366,N_589);
nor U1114 (N_1114,N_553,N_394);
or U1115 (N_1115,N_82,N_261);
and U1116 (N_1116,N_217,N_266);
nor U1117 (N_1117,N_265,N_507);
nor U1118 (N_1118,N_581,N_576);
and U1119 (N_1119,N_284,N_152);
or U1120 (N_1120,N_33,N_235);
or U1121 (N_1121,N_376,N_24);
and U1122 (N_1122,N_527,N_108);
nor U1123 (N_1123,N_587,N_481);
and U1124 (N_1124,N_127,N_487);
and U1125 (N_1125,N_207,N_580);
and U1126 (N_1126,N_18,N_53);
nand U1127 (N_1127,N_234,N_452);
nand U1128 (N_1128,N_1,N_583);
and U1129 (N_1129,N_193,N_241);
or U1130 (N_1130,N_471,N_571);
nand U1131 (N_1131,N_3,N_227);
nand U1132 (N_1132,N_199,N_396);
nor U1133 (N_1133,N_94,N_79);
nor U1134 (N_1134,N_312,N_519);
and U1135 (N_1135,N_166,N_73);
or U1136 (N_1136,N_427,N_372);
nor U1137 (N_1137,N_309,N_110);
nand U1138 (N_1138,N_302,N_424);
and U1139 (N_1139,N_83,N_503);
nor U1140 (N_1140,N_452,N_282);
and U1141 (N_1141,N_450,N_319);
nor U1142 (N_1142,N_47,N_219);
and U1143 (N_1143,N_597,N_167);
nand U1144 (N_1144,N_387,N_486);
nand U1145 (N_1145,N_565,N_253);
or U1146 (N_1146,N_102,N_66);
and U1147 (N_1147,N_496,N_426);
nand U1148 (N_1148,N_87,N_208);
nor U1149 (N_1149,N_518,N_224);
or U1150 (N_1150,N_482,N_35);
and U1151 (N_1151,N_38,N_0);
nand U1152 (N_1152,N_531,N_510);
or U1153 (N_1153,N_589,N_202);
and U1154 (N_1154,N_194,N_172);
and U1155 (N_1155,N_284,N_588);
and U1156 (N_1156,N_599,N_101);
xor U1157 (N_1157,N_401,N_91);
nor U1158 (N_1158,N_9,N_401);
and U1159 (N_1159,N_250,N_597);
or U1160 (N_1160,N_69,N_110);
nor U1161 (N_1161,N_582,N_462);
nor U1162 (N_1162,N_436,N_85);
nand U1163 (N_1163,N_204,N_187);
nor U1164 (N_1164,N_301,N_281);
and U1165 (N_1165,N_555,N_431);
or U1166 (N_1166,N_566,N_125);
or U1167 (N_1167,N_340,N_436);
or U1168 (N_1168,N_172,N_227);
nand U1169 (N_1169,N_507,N_529);
or U1170 (N_1170,N_405,N_21);
or U1171 (N_1171,N_109,N_572);
nor U1172 (N_1172,N_12,N_590);
or U1173 (N_1173,N_464,N_282);
nand U1174 (N_1174,N_290,N_441);
and U1175 (N_1175,N_435,N_36);
nand U1176 (N_1176,N_55,N_343);
nand U1177 (N_1177,N_202,N_368);
or U1178 (N_1178,N_571,N_44);
nand U1179 (N_1179,N_387,N_534);
nand U1180 (N_1180,N_84,N_349);
and U1181 (N_1181,N_521,N_103);
or U1182 (N_1182,N_145,N_47);
nor U1183 (N_1183,N_465,N_93);
and U1184 (N_1184,N_224,N_318);
or U1185 (N_1185,N_127,N_432);
or U1186 (N_1186,N_530,N_177);
and U1187 (N_1187,N_546,N_142);
or U1188 (N_1188,N_59,N_27);
and U1189 (N_1189,N_26,N_576);
nand U1190 (N_1190,N_524,N_426);
nand U1191 (N_1191,N_15,N_58);
or U1192 (N_1192,N_328,N_23);
nor U1193 (N_1193,N_372,N_449);
xnor U1194 (N_1194,N_4,N_293);
or U1195 (N_1195,N_238,N_163);
or U1196 (N_1196,N_6,N_237);
nand U1197 (N_1197,N_110,N_286);
nor U1198 (N_1198,N_75,N_264);
nor U1199 (N_1199,N_260,N_216);
and U1200 (N_1200,N_891,N_993);
and U1201 (N_1201,N_1000,N_652);
nand U1202 (N_1202,N_1179,N_991);
nor U1203 (N_1203,N_1114,N_853);
xor U1204 (N_1204,N_1007,N_833);
xnor U1205 (N_1205,N_619,N_631);
or U1206 (N_1206,N_675,N_1149);
nand U1207 (N_1207,N_963,N_986);
nand U1208 (N_1208,N_695,N_712);
or U1209 (N_1209,N_831,N_682);
nand U1210 (N_1210,N_733,N_813);
nor U1211 (N_1211,N_753,N_697);
nand U1212 (N_1212,N_1145,N_776);
and U1213 (N_1213,N_601,N_1096);
and U1214 (N_1214,N_981,N_724);
or U1215 (N_1215,N_613,N_1083);
nand U1216 (N_1216,N_1090,N_961);
nor U1217 (N_1217,N_1069,N_901);
nand U1218 (N_1218,N_691,N_1188);
nor U1219 (N_1219,N_795,N_842);
nand U1220 (N_1220,N_706,N_932);
nor U1221 (N_1221,N_827,N_1061);
or U1222 (N_1222,N_714,N_1056);
nor U1223 (N_1223,N_726,N_1146);
and U1224 (N_1224,N_1139,N_1196);
xor U1225 (N_1225,N_994,N_838);
or U1226 (N_1226,N_990,N_1162);
and U1227 (N_1227,N_1059,N_738);
and U1228 (N_1228,N_851,N_1161);
nor U1229 (N_1229,N_925,N_1077);
and U1230 (N_1230,N_1022,N_1187);
nand U1231 (N_1231,N_600,N_686);
nand U1232 (N_1232,N_717,N_1137);
nand U1233 (N_1233,N_974,N_629);
nor U1234 (N_1234,N_657,N_1078);
nand U1235 (N_1235,N_926,N_905);
or U1236 (N_1236,N_782,N_1042);
nand U1237 (N_1237,N_823,N_1154);
nor U1238 (N_1238,N_1140,N_1191);
or U1239 (N_1239,N_933,N_903);
and U1240 (N_1240,N_760,N_667);
or U1241 (N_1241,N_972,N_1067);
or U1242 (N_1242,N_1173,N_856);
nor U1243 (N_1243,N_1117,N_650);
nor U1244 (N_1244,N_1144,N_989);
nor U1245 (N_1245,N_1047,N_958);
or U1246 (N_1246,N_966,N_704);
nand U1247 (N_1247,N_1171,N_718);
and U1248 (N_1248,N_895,N_1138);
nor U1249 (N_1249,N_1102,N_946);
nor U1250 (N_1250,N_1091,N_832);
nand U1251 (N_1251,N_900,N_1118);
nand U1252 (N_1252,N_790,N_984);
nand U1253 (N_1253,N_1031,N_936);
nor U1254 (N_1254,N_1073,N_744);
nand U1255 (N_1255,N_767,N_956);
and U1256 (N_1256,N_638,N_954);
nor U1257 (N_1257,N_747,N_935);
or U1258 (N_1258,N_672,N_834);
or U1259 (N_1259,N_1155,N_939);
and U1260 (N_1260,N_996,N_1160);
nand U1261 (N_1261,N_916,N_1098);
nand U1262 (N_1262,N_1040,N_713);
nor U1263 (N_1263,N_668,N_907);
nand U1264 (N_1264,N_1027,N_847);
or U1265 (N_1265,N_983,N_766);
nand U1266 (N_1266,N_729,N_752);
nor U1267 (N_1267,N_978,N_693);
or U1268 (N_1268,N_878,N_858);
or U1269 (N_1269,N_772,N_844);
nand U1270 (N_1270,N_977,N_950);
or U1271 (N_1271,N_1029,N_841);
nor U1272 (N_1272,N_642,N_985);
or U1273 (N_1273,N_1026,N_666);
nand U1274 (N_1274,N_783,N_1051);
nand U1275 (N_1275,N_787,N_734);
nand U1276 (N_1276,N_799,N_1112);
and U1277 (N_1277,N_988,N_623);
or U1278 (N_1278,N_618,N_867);
and U1279 (N_1279,N_775,N_997);
and U1280 (N_1280,N_865,N_982);
nand U1281 (N_1281,N_725,N_1108);
nand U1282 (N_1282,N_1038,N_641);
or U1283 (N_1283,N_645,N_1133);
nor U1284 (N_1284,N_845,N_883);
nand U1285 (N_1285,N_625,N_882);
and U1286 (N_1286,N_944,N_816);
nand U1287 (N_1287,N_801,N_611);
xnor U1288 (N_1288,N_980,N_1192);
and U1289 (N_1289,N_646,N_622);
or U1290 (N_1290,N_605,N_931);
and U1291 (N_1291,N_1184,N_949);
xnor U1292 (N_1292,N_890,N_880);
or U1293 (N_1293,N_665,N_1158);
xnor U1294 (N_1294,N_751,N_971);
and U1295 (N_1295,N_929,N_952);
nor U1296 (N_1296,N_1055,N_617);
or U1297 (N_1297,N_1064,N_948);
and U1298 (N_1298,N_736,N_1034);
nand U1299 (N_1299,N_941,N_648);
or U1300 (N_1300,N_943,N_1082);
and U1301 (N_1301,N_877,N_1036);
nor U1302 (N_1302,N_679,N_959);
nor U1303 (N_1303,N_1121,N_764);
nor U1304 (N_1304,N_1057,N_788);
nand U1305 (N_1305,N_859,N_663);
or U1306 (N_1306,N_830,N_1185);
nor U1307 (N_1307,N_659,N_1186);
nor U1308 (N_1308,N_633,N_615);
nand U1309 (N_1309,N_771,N_1001);
and U1310 (N_1310,N_1014,N_694);
nand U1311 (N_1311,N_967,N_1157);
nor U1312 (N_1312,N_715,N_762);
or U1313 (N_1313,N_1103,N_635);
nand U1314 (N_1314,N_904,N_849);
or U1315 (N_1315,N_873,N_870);
or U1316 (N_1316,N_720,N_683);
or U1317 (N_1317,N_909,N_1089);
and U1318 (N_1318,N_1039,N_848);
nand U1319 (N_1319,N_1127,N_604);
and U1320 (N_1320,N_864,N_1141);
nand U1321 (N_1321,N_857,N_892);
and U1322 (N_1322,N_721,N_1130);
nand U1323 (N_1323,N_784,N_746);
or U1324 (N_1324,N_808,N_1018);
nand U1325 (N_1325,N_837,N_653);
nor U1326 (N_1326,N_1088,N_1166);
nor U1327 (N_1327,N_1104,N_866);
nand U1328 (N_1328,N_1156,N_962);
and U1329 (N_1329,N_850,N_1052);
and U1330 (N_1330,N_1068,N_1150);
or U1331 (N_1331,N_1107,N_942);
nand U1332 (N_1332,N_698,N_1165);
and U1333 (N_1333,N_610,N_687);
or U1334 (N_1334,N_681,N_658);
nor U1335 (N_1335,N_781,N_976);
and U1336 (N_1336,N_1004,N_1116);
nor U1337 (N_1337,N_1147,N_822);
nand U1338 (N_1338,N_701,N_937);
or U1339 (N_1339,N_1198,N_1050);
and U1340 (N_1340,N_829,N_1076);
nand U1341 (N_1341,N_602,N_624);
and U1342 (N_1342,N_777,N_758);
or U1343 (N_1343,N_1013,N_1005);
and U1344 (N_1344,N_1066,N_894);
or U1345 (N_1345,N_1016,N_908);
and U1346 (N_1346,N_906,N_616);
nand U1347 (N_1347,N_1062,N_1123);
nand U1348 (N_1348,N_1169,N_1093);
nor U1349 (N_1349,N_912,N_999);
nand U1350 (N_1350,N_780,N_940);
or U1351 (N_1351,N_709,N_1106);
or U1352 (N_1352,N_1135,N_1010);
nor U1353 (N_1353,N_921,N_674);
or U1354 (N_1354,N_1177,N_632);
nor U1355 (N_1355,N_1105,N_710);
nor U1356 (N_1356,N_1041,N_647);
nor U1357 (N_1357,N_608,N_1087);
nor U1358 (N_1358,N_868,N_913);
or U1359 (N_1359,N_1129,N_627);
or U1360 (N_1360,N_732,N_910);
and U1361 (N_1361,N_819,N_885);
nand U1362 (N_1362,N_798,N_620);
or U1363 (N_1363,N_1136,N_696);
nand U1364 (N_1364,N_1178,N_1113);
and U1365 (N_1365,N_1125,N_778);
nor U1366 (N_1366,N_745,N_951);
nor U1367 (N_1367,N_1019,N_1190);
and U1368 (N_1368,N_804,N_998);
and U1369 (N_1369,N_1080,N_930);
and U1370 (N_1370,N_728,N_1070);
nand U1371 (N_1371,N_793,N_785);
nand U1372 (N_1372,N_970,N_992);
and U1373 (N_1373,N_684,N_651);
and U1374 (N_1374,N_1170,N_1058);
or U1375 (N_1375,N_923,N_810);
nor U1376 (N_1376,N_1115,N_1167);
nand U1377 (N_1377,N_737,N_1028);
or U1378 (N_1378,N_973,N_1189);
nor U1379 (N_1379,N_680,N_1100);
nand U1380 (N_1380,N_609,N_671);
or U1381 (N_1381,N_769,N_914);
nand U1382 (N_1382,N_664,N_741);
nand U1383 (N_1383,N_626,N_1037);
and U1384 (N_1384,N_750,N_630);
or U1385 (N_1385,N_662,N_1194);
nand U1386 (N_1386,N_874,N_723);
or U1387 (N_1387,N_655,N_792);
or U1388 (N_1388,N_805,N_628);
nor U1389 (N_1389,N_1152,N_1111);
nor U1390 (N_1390,N_1151,N_881);
and U1391 (N_1391,N_828,N_897);
or U1392 (N_1392,N_794,N_1148);
and U1393 (N_1393,N_779,N_1181);
nand U1394 (N_1394,N_1099,N_898);
and U1395 (N_1395,N_1126,N_1163);
xnor U1396 (N_1396,N_824,N_614);
and U1397 (N_1397,N_634,N_700);
nor U1398 (N_1398,N_708,N_995);
nand U1399 (N_1399,N_654,N_739);
nand U1400 (N_1400,N_786,N_1164);
nor U1401 (N_1401,N_884,N_705);
and U1402 (N_1402,N_1048,N_748);
or U1403 (N_1403,N_927,N_869);
and U1404 (N_1404,N_922,N_742);
nor U1405 (N_1405,N_643,N_670);
nand U1406 (N_1406,N_644,N_975);
nand U1407 (N_1407,N_768,N_1006);
and U1408 (N_1408,N_773,N_1095);
nand U1409 (N_1409,N_863,N_789);
or U1410 (N_1410,N_1176,N_1053);
nor U1411 (N_1411,N_1109,N_1197);
nor U1412 (N_1412,N_1046,N_835);
nand U1413 (N_1413,N_1092,N_1024);
nor U1414 (N_1414,N_1044,N_957);
and U1415 (N_1415,N_920,N_756);
nand U1416 (N_1416,N_919,N_802);
or U1417 (N_1417,N_1097,N_1025);
or U1418 (N_1418,N_678,N_757);
or U1419 (N_1419,N_699,N_1049);
nor U1420 (N_1420,N_1180,N_814);
nand U1421 (N_1421,N_839,N_1182);
nor U1422 (N_1422,N_915,N_702);
or U1423 (N_1423,N_888,N_676);
or U1424 (N_1424,N_1065,N_812);
and U1425 (N_1425,N_1045,N_1128);
nand U1426 (N_1426,N_797,N_918);
or U1427 (N_1427,N_862,N_1183);
xnor U1428 (N_1428,N_1075,N_924);
nor U1429 (N_1429,N_1074,N_1168);
nor U1430 (N_1430,N_1009,N_1193);
xnor U1431 (N_1431,N_879,N_917);
and U1432 (N_1432,N_843,N_807);
and U1433 (N_1433,N_1085,N_1119);
nor U1434 (N_1434,N_763,N_612);
nor U1435 (N_1435,N_1017,N_1079);
or U1436 (N_1436,N_637,N_938);
nor U1437 (N_1437,N_1134,N_673);
nor U1438 (N_1438,N_755,N_1120);
nor U1439 (N_1439,N_953,N_1143);
nand U1440 (N_1440,N_1008,N_1003);
and U1441 (N_1441,N_1033,N_719);
xor U1442 (N_1442,N_886,N_902);
or U1443 (N_1443,N_735,N_722);
nor U1444 (N_1444,N_1174,N_1035);
nand U1445 (N_1445,N_660,N_1086);
nand U1446 (N_1446,N_796,N_846);
or U1447 (N_1447,N_821,N_911);
and U1448 (N_1448,N_1175,N_955);
nor U1449 (N_1449,N_690,N_759);
and U1450 (N_1450,N_945,N_607);
nor U1451 (N_1451,N_934,N_854);
nand U1452 (N_1452,N_876,N_688);
and U1453 (N_1453,N_852,N_899);
nor U1454 (N_1454,N_711,N_603);
and U1455 (N_1455,N_1084,N_656);
and U1456 (N_1456,N_1021,N_1159);
nor U1457 (N_1457,N_871,N_964);
nor U1458 (N_1458,N_749,N_639);
or U1459 (N_1459,N_987,N_893);
or U1460 (N_1460,N_928,N_730);
nor U1461 (N_1461,N_969,N_818);
nand U1462 (N_1462,N_685,N_1132);
nand U1463 (N_1463,N_743,N_806);
nor U1464 (N_1464,N_1142,N_1094);
and U1465 (N_1465,N_765,N_836);
nand U1466 (N_1466,N_661,N_731);
nand U1467 (N_1467,N_1015,N_1060);
xor U1468 (N_1468,N_875,N_826);
nand U1469 (N_1469,N_968,N_1054);
xor U1470 (N_1470,N_803,N_855);
or U1471 (N_1471,N_1030,N_809);
or U1472 (N_1472,N_1110,N_640);
nor U1473 (N_1473,N_1081,N_861);
and U1474 (N_1474,N_1002,N_1131);
or U1475 (N_1475,N_1020,N_825);
nand U1476 (N_1476,N_1195,N_947);
or U1477 (N_1477,N_811,N_815);
or U1478 (N_1478,N_979,N_1063);
and U1479 (N_1479,N_791,N_860);
nor U1480 (N_1480,N_716,N_1124);
and U1481 (N_1481,N_840,N_761);
nand U1482 (N_1482,N_800,N_896);
nand U1483 (N_1483,N_1071,N_960);
nand U1484 (N_1484,N_677,N_606);
or U1485 (N_1485,N_727,N_889);
nand U1486 (N_1486,N_965,N_669);
xnor U1487 (N_1487,N_1101,N_1032);
nand U1488 (N_1488,N_621,N_754);
nand U1489 (N_1489,N_817,N_707);
xor U1490 (N_1490,N_689,N_692);
or U1491 (N_1491,N_740,N_1153);
or U1492 (N_1492,N_872,N_774);
nand U1493 (N_1493,N_1072,N_1023);
nor U1494 (N_1494,N_820,N_1199);
nand U1495 (N_1495,N_1012,N_770);
or U1496 (N_1496,N_649,N_1011);
or U1497 (N_1497,N_1122,N_887);
or U1498 (N_1498,N_1172,N_1043);
xor U1499 (N_1499,N_636,N_703);
or U1500 (N_1500,N_965,N_934);
and U1501 (N_1501,N_1160,N_1185);
and U1502 (N_1502,N_728,N_842);
nand U1503 (N_1503,N_1031,N_901);
nand U1504 (N_1504,N_613,N_929);
nor U1505 (N_1505,N_948,N_873);
nand U1506 (N_1506,N_928,N_1070);
nand U1507 (N_1507,N_864,N_731);
nand U1508 (N_1508,N_681,N_1171);
nor U1509 (N_1509,N_619,N_801);
or U1510 (N_1510,N_879,N_834);
or U1511 (N_1511,N_955,N_1166);
nor U1512 (N_1512,N_744,N_697);
nand U1513 (N_1513,N_1091,N_1050);
nand U1514 (N_1514,N_652,N_662);
nor U1515 (N_1515,N_925,N_930);
or U1516 (N_1516,N_1100,N_1003);
or U1517 (N_1517,N_1134,N_1010);
nand U1518 (N_1518,N_680,N_872);
nor U1519 (N_1519,N_619,N_660);
or U1520 (N_1520,N_1064,N_1006);
nand U1521 (N_1521,N_681,N_1005);
or U1522 (N_1522,N_788,N_730);
nor U1523 (N_1523,N_1168,N_1008);
or U1524 (N_1524,N_912,N_674);
xor U1525 (N_1525,N_1067,N_1148);
xor U1526 (N_1526,N_817,N_1016);
xnor U1527 (N_1527,N_1106,N_982);
nor U1528 (N_1528,N_1050,N_1058);
and U1529 (N_1529,N_652,N_954);
and U1530 (N_1530,N_1176,N_944);
nand U1531 (N_1531,N_899,N_901);
nand U1532 (N_1532,N_623,N_1126);
nor U1533 (N_1533,N_800,N_769);
nor U1534 (N_1534,N_1043,N_1133);
and U1535 (N_1535,N_1104,N_953);
nand U1536 (N_1536,N_1183,N_846);
and U1537 (N_1537,N_1115,N_1102);
nand U1538 (N_1538,N_954,N_739);
nor U1539 (N_1539,N_971,N_659);
nor U1540 (N_1540,N_859,N_645);
or U1541 (N_1541,N_1118,N_623);
or U1542 (N_1542,N_974,N_862);
nor U1543 (N_1543,N_685,N_756);
nand U1544 (N_1544,N_725,N_732);
and U1545 (N_1545,N_1053,N_808);
nand U1546 (N_1546,N_847,N_795);
nand U1547 (N_1547,N_977,N_737);
nor U1548 (N_1548,N_852,N_989);
nor U1549 (N_1549,N_1092,N_662);
nand U1550 (N_1550,N_1168,N_839);
and U1551 (N_1551,N_1094,N_629);
and U1552 (N_1552,N_953,N_755);
or U1553 (N_1553,N_976,N_1033);
nor U1554 (N_1554,N_1184,N_765);
nand U1555 (N_1555,N_1046,N_1075);
nand U1556 (N_1556,N_885,N_1028);
and U1557 (N_1557,N_1083,N_684);
and U1558 (N_1558,N_646,N_744);
and U1559 (N_1559,N_1022,N_1146);
nor U1560 (N_1560,N_613,N_1148);
nor U1561 (N_1561,N_836,N_1060);
nor U1562 (N_1562,N_1148,N_737);
nand U1563 (N_1563,N_672,N_765);
nand U1564 (N_1564,N_1067,N_950);
nor U1565 (N_1565,N_1169,N_715);
nand U1566 (N_1566,N_753,N_724);
nor U1567 (N_1567,N_708,N_971);
and U1568 (N_1568,N_926,N_603);
nand U1569 (N_1569,N_1060,N_926);
nor U1570 (N_1570,N_943,N_793);
nand U1571 (N_1571,N_886,N_1089);
and U1572 (N_1572,N_1170,N_841);
nor U1573 (N_1573,N_736,N_617);
xor U1574 (N_1574,N_1048,N_910);
or U1575 (N_1575,N_647,N_1115);
nand U1576 (N_1576,N_606,N_868);
and U1577 (N_1577,N_1027,N_791);
and U1578 (N_1578,N_615,N_1159);
or U1579 (N_1579,N_781,N_1139);
nor U1580 (N_1580,N_1118,N_1106);
or U1581 (N_1581,N_1150,N_845);
nand U1582 (N_1582,N_1183,N_1187);
and U1583 (N_1583,N_1111,N_842);
nor U1584 (N_1584,N_816,N_621);
and U1585 (N_1585,N_1038,N_1004);
nand U1586 (N_1586,N_820,N_1083);
nor U1587 (N_1587,N_834,N_646);
and U1588 (N_1588,N_1119,N_1075);
or U1589 (N_1589,N_786,N_1191);
and U1590 (N_1590,N_763,N_843);
nor U1591 (N_1591,N_1018,N_1001);
and U1592 (N_1592,N_749,N_744);
nand U1593 (N_1593,N_646,N_685);
and U1594 (N_1594,N_915,N_709);
or U1595 (N_1595,N_808,N_1042);
and U1596 (N_1596,N_802,N_668);
nor U1597 (N_1597,N_873,N_885);
or U1598 (N_1598,N_835,N_1041);
or U1599 (N_1599,N_791,N_1117);
nor U1600 (N_1600,N_1140,N_1182);
and U1601 (N_1601,N_917,N_853);
or U1602 (N_1602,N_1147,N_912);
nand U1603 (N_1603,N_753,N_814);
nor U1604 (N_1604,N_860,N_970);
nand U1605 (N_1605,N_1061,N_736);
and U1606 (N_1606,N_1056,N_743);
and U1607 (N_1607,N_847,N_934);
and U1608 (N_1608,N_675,N_870);
or U1609 (N_1609,N_1103,N_629);
nand U1610 (N_1610,N_1070,N_1032);
xnor U1611 (N_1611,N_1017,N_772);
and U1612 (N_1612,N_1187,N_624);
or U1613 (N_1613,N_1067,N_709);
nor U1614 (N_1614,N_604,N_755);
and U1615 (N_1615,N_1156,N_721);
or U1616 (N_1616,N_754,N_897);
and U1617 (N_1617,N_1006,N_1162);
and U1618 (N_1618,N_661,N_936);
nor U1619 (N_1619,N_763,N_1030);
or U1620 (N_1620,N_1160,N_821);
nor U1621 (N_1621,N_627,N_1080);
nor U1622 (N_1622,N_1103,N_1061);
or U1623 (N_1623,N_956,N_684);
nand U1624 (N_1624,N_617,N_1081);
or U1625 (N_1625,N_862,N_1148);
nand U1626 (N_1626,N_722,N_1102);
nand U1627 (N_1627,N_616,N_996);
or U1628 (N_1628,N_785,N_827);
nor U1629 (N_1629,N_1007,N_791);
nor U1630 (N_1630,N_958,N_908);
nor U1631 (N_1631,N_653,N_838);
nand U1632 (N_1632,N_816,N_918);
or U1633 (N_1633,N_982,N_827);
and U1634 (N_1634,N_1092,N_940);
nand U1635 (N_1635,N_702,N_1188);
and U1636 (N_1636,N_706,N_1016);
or U1637 (N_1637,N_1150,N_763);
xnor U1638 (N_1638,N_813,N_808);
or U1639 (N_1639,N_837,N_1138);
or U1640 (N_1640,N_612,N_1194);
nand U1641 (N_1641,N_738,N_1028);
xor U1642 (N_1642,N_1033,N_843);
or U1643 (N_1643,N_1189,N_970);
xnor U1644 (N_1644,N_765,N_1054);
and U1645 (N_1645,N_1146,N_623);
nor U1646 (N_1646,N_857,N_669);
nand U1647 (N_1647,N_1122,N_866);
nand U1648 (N_1648,N_682,N_1149);
and U1649 (N_1649,N_1096,N_1024);
nor U1650 (N_1650,N_616,N_1123);
and U1651 (N_1651,N_688,N_828);
nor U1652 (N_1652,N_1124,N_1080);
and U1653 (N_1653,N_859,N_1164);
nand U1654 (N_1654,N_1141,N_1074);
xnor U1655 (N_1655,N_1083,N_765);
nor U1656 (N_1656,N_620,N_684);
nand U1657 (N_1657,N_653,N_778);
or U1658 (N_1658,N_963,N_747);
nor U1659 (N_1659,N_1160,N_709);
nor U1660 (N_1660,N_710,N_1100);
nor U1661 (N_1661,N_720,N_772);
nor U1662 (N_1662,N_1100,N_718);
xor U1663 (N_1663,N_785,N_662);
nor U1664 (N_1664,N_1141,N_771);
nor U1665 (N_1665,N_961,N_819);
and U1666 (N_1666,N_1032,N_656);
nor U1667 (N_1667,N_1152,N_1159);
nor U1668 (N_1668,N_658,N_1171);
or U1669 (N_1669,N_989,N_821);
nor U1670 (N_1670,N_720,N_827);
or U1671 (N_1671,N_730,N_1059);
nand U1672 (N_1672,N_934,N_1065);
nand U1673 (N_1673,N_902,N_601);
or U1674 (N_1674,N_1134,N_1052);
nand U1675 (N_1675,N_1096,N_851);
or U1676 (N_1676,N_1139,N_1021);
and U1677 (N_1677,N_718,N_729);
nand U1678 (N_1678,N_1063,N_615);
nor U1679 (N_1679,N_1053,N_623);
nor U1680 (N_1680,N_1100,N_698);
and U1681 (N_1681,N_738,N_1036);
nand U1682 (N_1682,N_1097,N_1193);
nand U1683 (N_1683,N_1084,N_601);
and U1684 (N_1684,N_982,N_932);
nor U1685 (N_1685,N_854,N_935);
nand U1686 (N_1686,N_820,N_950);
nor U1687 (N_1687,N_661,N_877);
and U1688 (N_1688,N_977,N_894);
or U1689 (N_1689,N_1196,N_1174);
nand U1690 (N_1690,N_770,N_862);
or U1691 (N_1691,N_958,N_1000);
or U1692 (N_1692,N_1199,N_773);
or U1693 (N_1693,N_968,N_1129);
and U1694 (N_1694,N_800,N_858);
and U1695 (N_1695,N_918,N_837);
nand U1696 (N_1696,N_1183,N_1182);
and U1697 (N_1697,N_929,N_1163);
nand U1698 (N_1698,N_1168,N_1157);
nand U1699 (N_1699,N_714,N_900);
or U1700 (N_1700,N_1168,N_790);
nand U1701 (N_1701,N_824,N_1138);
and U1702 (N_1702,N_838,N_620);
nand U1703 (N_1703,N_906,N_1141);
nand U1704 (N_1704,N_742,N_946);
nand U1705 (N_1705,N_734,N_1172);
nor U1706 (N_1706,N_986,N_664);
nor U1707 (N_1707,N_854,N_644);
or U1708 (N_1708,N_948,N_1011);
nand U1709 (N_1709,N_1016,N_616);
nand U1710 (N_1710,N_1145,N_961);
or U1711 (N_1711,N_743,N_809);
or U1712 (N_1712,N_1179,N_1149);
or U1713 (N_1713,N_1088,N_739);
or U1714 (N_1714,N_1000,N_711);
or U1715 (N_1715,N_621,N_710);
nand U1716 (N_1716,N_843,N_647);
nand U1717 (N_1717,N_996,N_700);
or U1718 (N_1718,N_1158,N_663);
nand U1719 (N_1719,N_897,N_805);
nor U1720 (N_1720,N_1175,N_1197);
nor U1721 (N_1721,N_1014,N_793);
nand U1722 (N_1722,N_660,N_919);
and U1723 (N_1723,N_925,N_828);
or U1724 (N_1724,N_1073,N_1092);
nand U1725 (N_1725,N_886,N_1078);
and U1726 (N_1726,N_659,N_777);
nand U1727 (N_1727,N_1022,N_650);
nor U1728 (N_1728,N_606,N_729);
and U1729 (N_1729,N_691,N_1112);
nand U1730 (N_1730,N_1132,N_892);
nor U1731 (N_1731,N_1131,N_867);
or U1732 (N_1732,N_862,N_887);
nand U1733 (N_1733,N_1165,N_1133);
nor U1734 (N_1734,N_1089,N_1010);
or U1735 (N_1735,N_1194,N_759);
or U1736 (N_1736,N_979,N_995);
or U1737 (N_1737,N_1131,N_893);
or U1738 (N_1738,N_865,N_1156);
and U1739 (N_1739,N_621,N_699);
nand U1740 (N_1740,N_1098,N_929);
and U1741 (N_1741,N_882,N_1020);
nand U1742 (N_1742,N_790,N_775);
nor U1743 (N_1743,N_880,N_1091);
nand U1744 (N_1744,N_611,N_1109);
and U1745 (N_1745,N_615,N_842);
nor U1746 (N_1746,N_628,N_1067);
nand U1747 (N_1747,N_678,N_635);
or U1748 (N_1748,N_773,N_863);
or U1749 (N_1749,N_1176,N_975);
or U1750 (N_1750,N_738,N_1149);
and U1751 (N_1751,N_1033,N_868);
nor U1752 (N_1752,N_962,N_899);
and U1753 (N_1753,N_702,N_1108);
and U1754 (N_1754,N_1075,N_891);
and U1755 (N_1755,N_623,N_870);
and U1756 (N_1756,N_1087,N_1055);
nand U1757 (N_1757,N_1047,N_927);
nor U1758 (N_1758,N_785,N_1054);
nor U1759 (N_1759,N_981,N_955);
and U1760 (N_1760,N_1193,N_641);
nand U1761 (N_1761,N_896,N_724);
and U1762 (N_1762,N_1036,N_610);
or U1763 (N_1763,N_1136,N_736);
or U1764 (N_1764,N_1158,N_960);
nor U1765 (N_1765,N_1188,N_878);
nor U1766 (N_1766,N_1157,N_1185);
and U1767 (N_1767,N_658,N_1139);
xnor U1768 (N_1768,N_967,N_800);
nor U1769 (N_1769,N_627,N_978);
or U1770 (N_1770,N_933,N_1180);
nor U1771 (N_1771,N_941,N_705);
nor U1772 (N_1772,N_843,N_677);
xnor U1773 (N_1773,N_1040,N_673);
nand U1774 (N_1774,N_1066,N_863);
xnor U1775 (N_1775,N_712,N_745);
or U1776 (N_1776,N_971,N_944);
or U1777 (N_1777,N_815,N_645);
and U1778 (N_1778,N_1097,N_677);
nand U1779 (N_1779,N_749,N_703);
nand U1780 (N_1780,N_952,N_752);
nand U1781 (N_1781,N_631,N_739);
and U1782 (N_1782,N_635,N_992);
nor U1783 (N_1783,N_898,N_1113);
or U1784 (N_1784,N_836,N_828);
nand U1785 (N_1785,N_1087,N_663);
or U1786 (N_1786,N_607,N_1001);
or U1787 (N_1787,N_893,N_1171);
nand U1788 (N_1788,N_991,N_601);
nand U1789 (N_1789,N_1001,N_972);
or U1790 (N_1790,N_1172,N_920);
and U1791 (N_1791,N_778,N_907);
or U1792 (N_1792,N_1122,N_888);
nand U1793 (N_1793,N_781,N_801);
nand U1794 (N_1794,N_653,N_1109);
nor U1795 (N_1795,N_1164,N_911);
nand U1796 (N_1796,N_1190,N_935);
xor U1797 (N_1797,N_1185,N_987);
nor U1798 (N_1798,N_1149,N_1035);
nand U1799 (N_1799,N_967,N_864);
and U1800 (N_1800,N_1697,N_1515);
nand U1801 (N_1801,N_1357,N_1304);
nor U1802 (N_1802,N_1762,N_1696);
nor U1803 (N_1803,N_1590,N_1373);
nor U1804 (N_1804,N_1300,N_1636);
nor U1805 (N_1805,N_1754,N_1608);
nand U1806 (N_1806,N_1435,N_1535);
or U1807 (N_1807,N_1688,N_1501);
nor U1808 (N_1808,N_1690,N_1629);
nor U1809 (N_1809,N_1581,N_1283);
nand U1810 (N_1810,N_1242,N_1232);
and U1811 (N_1811,N_1675,N_1423);
nor U1812 (N_1812,N_1322,N_1459);
and U1813 (N_1813,N_1781,N_1390);
or U1814 (N_1814,N_1551,N_1292);
or U1815 (N_1815,N_1352,N_1479);
nand U1816 (N_1816,N_1389,N_1396);
and U1817 (N_1817,N_1585,N_1750);
and U1818 (N_1818,N_1529,N_1611);
and U1819 (N_1819,N_1673,N_1603);
nand U1820 (N_1820,N_1470,N_1455);
and U1821 (N_1821,N_1260,N_1271);
and U1822 (N_1822,N_1453,N_1214);
or U1823 (N_1823,N_1244,N_1667);
and U1824 (N_1824,N_1538,N_1202);
and U1825 (N_1825,N_1285,N_1741);
or U1826 (N_1826,N_1561,N_1384);
and U1827 (N_1827,N_1262,N_1496);
or U1828 (N_1828,N_1481,N_1719);
and U1829 (N_1829,N_1513,N_1734);
and U1830 (N_1830,N_1647,N_1744);
nand U1831 (N_1831,N_1256,N_1446);
or U1832 (N_1832,N_1722,N_1520);
nor U1833 (N_1833,N_1691,N_1649);
nor U1834 (N_1834,N_1725,N_1707);
and U1835 (N_1835,N_1245,N_1503);
and U1836 (N_1836,N_1703,N_1718);
and U1837 (N_1837,N_1411,N_1648);
nor U1838 (N_1838,N_1668,N_1205);
and U1839 (N_1839,N_1249,N_1445);
or U1840 (N_1840,N_1223,N_1494);
nand U1841 (N_1841,N_1358,N_1272);
and U1842 (N_1842,N_1536,N_1444);
and U1843 (N_1843,N_1758,N_1577);
and U1844 (N_1844,N_1493,N_1278);
and U1845 (N_1845,N_1416,N_1462);
nand U1846 (N_1846,N_1364,N_1442);
or U1847 (N_1847,N_1452,N_1236);
or U1848 (N_1848,N_1213,N_1710);
nand U1849 (N_1849,N_1631,N_1708);
nor U1850 (N_1850,N_1557,N_1552);
nor U1851 (N_1851,N_1316,N_1227);
or U1852 (N_1852,N_1517,N_1568);
or U1853 (N_1853,N_1425,N_1458);
and U1854 (N_1854,N_1429,N_1628);
nand U1855 (N_1855,N_1349,N_1763);
and U1856 (N_1856,N_1752,N_1778);
or U1857 (N_1857,N_1676,N_1642);
nor U1858 (N_1858,N_1487,N_1461);
nand U1859 (N_1859,N_1367,N_1267);
nand U1860 (N_1860,N_1702,N_1477);
nor U1861 (N_1861,N_1619,N_1408);
or U1862 (N_1862,N_1525,N_1790);
nand U1863 (N_1863,N_1595,N_1254);
and U1864 (N_1864,N_1243,N_1397);
nand U1865 (N_1865,N_1341,N_1250);
nand U1866 (N_1866,N_1468,N_1201);
nand U1867 (N_1867,N_1726,N_1749);
or U1868 (N_1868,N_1692,N_1622);
and U1869 (N_1869,N_1712,N_1465);
nor U1870 (N_1870,N_1727,N_1414);
or U1871 (N_1871,N_1216,N_1701);
and U1872 (N_1872,N_1606,N_1544);
and U1873 (N_1873,N_1645,N_1366);
nand U1874 (N_1874,N_1514,N_1545);
or U1875 (N_1875,N_1251,N_1559);
nand U1876 (N_1876,N_1303,N_1774);
nand U1877 (N_1877,N_1344,N_1296);
nand U1878 (N_1878,N_1746,N_1208);
nand U1879 (N_1879,N_1368,N_1728);
nand U1880 (N_1880,N_1795,N_1263);
and U1881 (N_1881,N_1714,N_1456);
and U1882 (N_1882,N_1314,N_1681);
and U1883 (N_1883,N_1342,N_1761);
and U1884 (N_1884,N_1679,N_1571);
or U1885 (N_1885,N_1365,N_1313);
nand U1886 (N_1886,N_1660,N_1326);
nor U1887 (N_1887,N_1471,N_1247);
or U1888 (N_1888,N_1755,N_1788);
nand U1889 (N_1889,N_1388,N_1226);
or U1890 (N_1890,N_1351,N_1683);
or U1891 (N_1891,N_1584,N_1343);
or U1892 (N_1892,N_1320,N_1640);
nand U1893 (N_1893,N_1522,N_1632);
nor U1894 (N_1894,N_1293,N_1532);
nor U1895 (N_1895,N_1682,N_1400);
nor U1896 (N_1896,N_1666,N_1233);
nand U1897 (N_1897,N_1528,N_1252);
and U1898 (N_1898,N_1488,N_1518);
nand U1899 (N_1899,N_1580,N_1328);
nand U1900 (N_1900,N_1258,N_1424);
or U1901 (N_1901,N_1508,N_1653);
and U1902 (N_1902,N_1530,N_1792);
and U1903 (N_1903,N_1554,N_1705);
nand U1904 (N_1904,N_1420,N_1486);
nand U1905 (N_1905,N_1583,N_1588);
nand U1906 (N_1906,N_1777,N_1434);
nor U1907 (N_1907,N_1637,N_1253);
and U1908 (N_1908,N_1573,N_1484);
and U1909 (N_1909,N_1467,N_1402);
and U1910 (N_1910,N_1599,N_1586);
nand U1911 (N_1911,N_1268,N_1562);
and U1912 (N_1912,N_1711,N_1549);
or U1913 (N_1913,N_1224,N_1785);
nor U1914 (N_1914,N_1298,N_1410);
or U1915 (N_1915,N_1371,N_1312);
nand U1916 (N_1916,N_1264,N_1541);
nor U1917 (N_1917,N_1421,N_1597);
xor U1918 (N_1918,N_1569,N_1798);
and U1919 (N_1919,N_1533,N_1780);
nand U1920 (N_1920,N_1413,N_1685);
nor U1921 (N_1921,N_1346,N_1572);
nand U1922 (N_1922,N_1306,N_1759);
nor U1923 (N_1923,N_1394,N_1497);
and U1924 (N_1924,N_1500,N_1209);
nand U1925 (N_1925,N_1732,N_1553);
nand U1926 (N_1926,N_1560,N_1650);
or U1927 (N_1927,N_1512,N_1450);
or U1928 (N_1928,N_1436,N_1729);
nor U1929 (N_1929,N_1475,N_1651);
nor U1930 (N_1930,N_1449,N_1624);
nand U1931 (N_1931,N_1724,N_1335);
and U1932 (N_1932,N_1381,N_1439);
nand U1933 (N_1933,N_1219,N_1318);
or U1934 (N_1934,N_1787,N_1451);
nand U1935 (N_1935,N_1638,N_1221);
nand U1936 (N_1936,N_1279,N_1354);
nand U1937 (N_1937,N_1212,N_1524);
nand U1938 (N_1938,N_1684,N_1600);
nand U1939 (N_1939,N_1401,N_1526);
or U1940 (N_1940,N_1796,N_1495);
nand U1941 (N_1941,N_1626,N_1558);
and U1942 (N_1942,N_1231,N_1229);
or U1943 (N_1943,N_1793,N_1745);
nand U1944 (N_1944,N_1203,N_1234);
and U1945 (N_1945,N_1259,N_1672);
nor U1946 (N_1946,N_1376,N_1677);
and U1947 (N_1947,N_1621,N_1776);
nand U1948 (N_1948,N_1771,N_1215);
or U1949 (N_1949,N_1634,N_1548);
nor U1950 (N_1950,N_1789,N_1274);
or U1951 (N_1951,N_1395,N_1472);
nand U1952 (N_1952,N_1598,N_1720);
and U1953 (N_1953,N_1294,N_1321);
nand U1954 (N_1954,N_1620,N_1578);
nand U1955 (N_1955,N_1307,N_1625);
and U1956 (N_1956,N_1669,N_1363);
nor U1957 (N_1957,N_1204,N_1345);
and U1958 (N_1958,N_1257,N_1301);
nor U1959 (N_1959,N_1616,N_1731);
nor U1960 (N_1960,N_1299,N_1540);
and U1961 (N_1961,N_1399,N_1733);
nand U1962 (N_1962,N_1700,N_1612);
or U1963 (N_1963,N_1469,N_1506);
and U1964 (N_1964,N_1398,N_1330);
nor U1965 (N_1965,N_1613,N_1695);
or U1966 (N_1966,N_1654,N_1288);
or U1967 (N_1967,N_1255,N_1239);
nor U1968 (N_1968,N_1510,N_1412);
or U1969 (N_1969,N_1238,N_1735);
and U1970 (N_1970,N_1543,N_1768);
or U1971 (N_1971,N_1633,N_1430);
or U1972 (N_1972,N_1483,N_1379);
and U1973 (N_1973,N_1601,N_1406);
nor U1974 (N_1974,N_1658,N_1457);
and U1975 (N_1975,N_1609,N_1337);
and U1976 (N_1976,N_1786,N_1375);
nand U1977 (N_1977,N_1441,N_1309);
nand U1978 (N_1978,N_1225,N_1721);
nand U1979 (N_1979,N_1448,N_1564);
or U1980 (N_1980,N_1280,N_1478);
nand U1981 (N_1981,N_1615,N_1407);
or U1982 (N_1982,N_1419,N_1607);
and U1983 (N_1983,N_1767,N_1217);
nand U1984 (N_1984,N_1431,N_1531);
nor U1985 (N_1985,N_1547,N_1218);
and U1986 (N_1986,N_1499,N_1686);
and U1987 (N_1987,N_1207,N_1291);
nor U1988 (N_1988,N_1383,N_1360);
nor U1989 (N_1989,N_1630,N_1485);
nor U1990 (N_1990,N_1556,N_1523);
nor U1991 (N_1991,N_1534,N_1610);
and U1992 (N_1992,N_1505,N_1327);
and U1993 (N_1993,N_1290,N_1386);
and U1994 (N_1994,N_1438,N_1593);
and U1995 (N_1995,N_1220,N_1378);
or U1996 (N_1996,N_1519,N_1241);
or U1997 (N_1997,N_1338,N_1374);
and U1998 (N_1998,N_1334,N_1305);
and U1999 (N_1999,N_1511,N_1287);
and U2000 (N_2000,N_1286,N_1656);
or U2001 (N_2001,N_1646,N_1466);
or U2002 (N_2002,N_1706,N_1332);
nand U2003 (N_2003,N_1694,N_1775);
and U2004 (N_2004,N_1211,N_1655);
nand U2005 (N_2005,N_1716,N_1644);
or U2006 (N_2006,N_1769,N_1605);
nor U2007 (N_2007,N_1403,N_1282);
nor U2008 (N_2008,N_1325,N_1333);
and U2009 (N_2009,N_1704,N_1773);
and U2010 (N_2010,N_1361,N_1340);
or U2011 (N_2011,N_1235,N_1579);
and U2012 (N_2012,N_1269,N_1418);
or U2013 (N_2013,N_1489,N_1210);
nor U2014 (N_2014,N_1427,N_1276);
nand U2015 (N_2015,N_1794,N_1743);
or U2016 (N_2016,N_1261,N_1504);
nand U2017 (N_2017,N_1392,N_1550);
nor U2018 (N_2018,N_1555,N_1738);
nand U2019 (N_2019,N_1369,N_1492);
or U2020 (N_2020,N_1302,N_1507);
nor U2021 (N_2021,N_1372,N_1473);
and U2022 (N_2022,N_1240,N_1490);
or U2023 (N_2023,N_1228,N_1324);
or U2024 (N_2024,N_1678,N_1385);
nand U2025 (N_2025,N_1464,N_1362);
and U2026 (N_2026,N_1281,N_1652);
nor U2027 (N_2027,N_1440,N_1230);
nand U2028 (N_2028,N_1737,N_1766);
and U2029 (N_2029,N_1336,N_1589);
or U2030 (N_2030,N_1270,N_1689);
or U2031 (N_2031,N_1592,N_1756);
xor U2032 (N_2032,N_1663,N_1331);
and U2033 (N_2033,N_1200,N_1657);
or U2034 (N_2034,N_1665,N_1757);
and U2035 (N_2035,N_1447,N_1317);
nor U2036 (N_2036,N_1742,N_1591);
nand U2037 (N_2037,N_1509,N_1680);
and U2038 (N_2038,N_1248,N_1614);
nand U2039 (N_2039,N_1779,N_1339);
nand U2040 (N_2040,N_1635,N_1347);
nand U2041 (N_2041,N_1687,N_1753);
nor U2042 (N_2042,N_1308,N_1246);
or U2043 (N_2043,N_1311,N_1723);
or U2044 (N_2044,N_1370,N_1623);
and U2045 (N_2045,N_1480,N_1206);
and U2046 (N_2046,N_1350,N_1432);
and U2047 (N_2047,N_1319,N_1491);
xor U2048 (N_2048,N_1641,N_1409);
or U2049 (N_2049,N_1782,N_1391);
or U2050 (N_2050,N_1751,N_1784);
and U2051 (N_2051,N_1516,N_1415);
or U2052 (N_2052,N_1387,N_1382);
or U2053 (N_2053,N_1618,N_1566);
nand U2054 (N_2054,N_1604,N_1498);
nor U2055 (N_2055,N_1627,N_1348);
or U2056 (N_2056,N_1428,N_1546);
or U2057 (N_2057,N_1422,N_1265);
nand U2058 (N_2058,N_1359,N_1799);
and U2059 (N_2059,N_1730,N_1567);
or U2060 (N_2060,N_1323,N_1765);
or U2061 (N_2061,N_1740,N_1393);
nand U2062 (N_2062,N_1222,N_1315);
or U2063 (N_2063,N_1404,N_1502);
nor U2064 (N_2064,N_1289,N_1594);
nor U2065 (N_2065,N_1310,N_1463);
and U2066 (N_2066,N_1443,N_1437);
nor U2067 (N_2067,N_1709,N_1377);
or U2068 (N_2068,N_1791,N_1674);
or U2069 (N_2069,N_1783,N_1659);
and U2070 (N_2070,N_1574,N_1275);
or U2071 (N_2071,N_1563,N_1454);
nand U2072 (N_2072,N_1575,N_1699);
and U2073 (N_2073,N_1474,N_1715);
or U2074 (N_2074,N_1670,N_1380);
or U2075 (N_2075,N_1295,N_1664);
and U2076 (N_2076,N_1539,N_1639);
nor U2077 (N_2077,N_1713,N_1356);
nor U2078 (N_2078,N_1671,N_1662);
nand U2079 (N_2079,N_1460,N_1570);
and U2080 (N_2080,N_1329,N_1277);
and U2081 (N_2081,N_1770,N_1426);
nor U2082 (N_2082,N_1596,N_1297);
nand U2083 (N_2083,N_1760,N_1772);
or U2084 (N_2084,N_1284,N_1693);
nor U2085 (N_2085,N_1748,N_1521);
nor U2086 (N_2086,N_1527,N_1617);
nor U2087 (N_2087,N_1273,N_1739);
or U2088 (N_2088,N_1565,N_1405);
nand U2089 (N_2089,N_1717,N_1537);
nor U2090 (N_2090,N_1747,N_1602);
or U2091 (N_2091,N_1353,N_1587);
nor U2092 (N_2092,N_1576,N_1736);
or U2093 (N_2093,N_1643,N_1266);
nand U2094 (N_2094,N_1417,N_1764);
nor U2095 (N_2095,N_1355,N_1797);
and U2096 (N_2096,N_1433,N_1582);
nand U2097 (N_2097,N_1698,N_1476);
nor U2098 (N_2098,N_1542,N_1237);
nor U2099 (N_2099,N_1661,N_1482);
nand U2100 (N_2100,N_1464,N_1314);
nand U2101 (N_2101,N_1453,N_1337);
nor U2102 (N_2102,N_1415,N_1778);
and U2103 (N_2103,N_1585,N_1434);
nand U2104 (N_2104,N_1578,N_1505);
nor U2105 (N_2105,N_1775,N_1731);
or U2106 (N_2106,N_1592,N_1740);
nand U2107 (N_2107,N_1383,N_1551);
nor U2108 (N_2108,N_1722,N_1471);
or U2109 (N_2109,N_1261,N_1431);
nand U2110 (N_2110,N_1642,N_1719);
nor U2111 (N_2111,N_1542,N_1207);
nor U2112 (N_2112,N_1359,N_1711);
nand U2113 (N_2113,N_1359,N_1216);
nand U2114 (N_2114,N_1744,N_1610);
or U2115 (N_2115,N_1695,N_1407);
and U2116 (N_2116,N_1360,N_1395);
or U2117 (N_2117,N_1799,N_1301);
and U2118 (N_2118,N_1456,N_1410);
nand U2119 (N_2119,N_1239,N_1287);
and U2120 (N_2120,N_1232,N_1471);
and U2121 (N_2121,N_1562,N_1791);
nor U2122 (N_2122,N_1411,N_1512);
nor U2123 (N_2123,N_1238,N_1604);
nor U2124 (N_2124,N_1700,N_1248);
or U2125 (N_2125,N_1681,N_1345);
nor U2126 (N_2126,N_1689,N_1571);
or U2127 (N_2127,N_1319,N_1664);
nor U2128 (N_2128,N_1487,N_1608);
nand U2129 (N_2129,N_1612,N_1567);
nor U2130 (N_2130,N_1225,N_1358);
or U2131 (N_2131,N_1669,N_1704);
nand U2132 (N_2132,N_1636,N_1495);
or U2133 (N_2133,N_1202,N_1722);
and U2134 (N_2134,N_1526,N_1249);
nor U2135 (N_2135,N_1607,N_1363);
and U2136 (N_2136,N_1352,N_1509);
xor U2137 (N_2137,N_1466,N_1465);
nand U2138 (N_2138,N_1724,N_1246);
nand U2139 (N_2139,N_1542,N_1611);
nor U2140 (N_2140,N_1537,N_1342);
and U2141 (N_2141,N_1739,N_1393);
or U2142 (N_2142,N_1295,N_1490);
nor U2143 (N_2143,N_1693,N_1219);
or U2144 (N_2144,N_1792,N_1436);
and U2145 (N_2145,N_1553,N_1258);
nand U2146 (N_2146,N_1520,N_1521);
nor U2147 (N_2147,N_1298,N_1732);
nor U2148 (N_2148,N_1695,N_1522);
nand U2149 (N_2149,N_1736,N_1748);
nand U2150 (N_2150,N_1690,N_1550);
or U2151 (N_2151,N_1653,N_1324);
or U2152 (N_2152,N_1286,N_1642);
nor U2153 (N_2153,N_1348,N_1397);
nor U2154 (N_2154,N_1591,N_1796);
nand U2155 (N_2155,N_1649,N_1456);
nor U2156 (N_2156,N_1547,N_1351);
nand U2157 (N_2157,N_1451,N_1366);
or U2158 (N_2158,N_1699,N_1751);
nand U2159 (N_2159,N_1721,N_1765);
or U2160 (N_2160,N_1642,N_1200);
or U2161 (N_2161,N_1236,N_1717);
or U2162 (N_2162,N_1246,N_1309);
and U2163 (N_2163,N_1434,N_1346);
or U2164 (N_2164,N_1756,N_1739);
or U2165 (N_2165,N_1304,N_1527);
nor U2166 (N_2166,N_1378,N_1579);
xor U2167 (N_2167,N_1656,N_1227);
and U2168 (N_2168,N_1485,N_1472);
or U2169 (N_2169,N_1715,N_1329);
nand U2170 (N_2170,N_1205,N_1506);
or U2171 (N_2171,N_1231,N_1292);
nand U2172 (N_2172,N_1500,N_1770);
and U2173 (N_2173,N_1279,N_1709);
or U2174 (N_2174,N_1769,N_1422);
and U2175 (N_2175,N_1209,N_1270);
nor U2176 (N_2176,N_1743,N_1426);
nor U2177 (N_2177,N_1363,N_1207);
and U2178 (N_2178,N_1617,N_1771);
and U2179 (N_2179,N_1410,N_1427);
and U2180 (N_2180,N_1224,N_1711);
or U2181 (N_2181,N_1309,N_1232);
or U2182 (N_2182,N_1594,N_1480);
nand U2183 (N_2183,N_1690,N_1509);
or U2184 (N_2184,N_1465,N_1456);
nor U2185 (N_2185,N_1644,N_1329);
xor U2186 (N_2186,N_1604,N_1686);
and U2187 (N_2187,N_1556,N_1290);
or U2188 (N_2188,N_1408,N_1751);
and U2189 (N_2189,N_1203,N_1591);
nand U2190 (N_2190,N_1747,N_1790);
nand U2191 (N_2191,N_1583,N_1523);
nand U2192 (N_2192,N_1462,N_1518);
and U2193 (N_2193,N_1309,N_1429);
and U2194 (N_2194,N_1535,N_1455);
and U2195 (N_2195,N_1662,N_1395);
or U2196 (N_2196,N_1512,N_1588);
nand U2197 (N_2197,N_1330,N_1565);
nor U2198 (N_2198,N_1494,N_1290);
nor U2199 (N_2199,N_1406,N_1242);
or U2200 (N_2200,N_1405,N_1762);
or U2201 (N_2201,N_1446,N_1362);
nor U2202 (N_2202,N_1528,N_1772);
nand U2203 (N_2203,N_1451,N_1326);
or U2204 (N_2204,N_1444,N_1378);
nand U2205 (N_2205,N_1307,N_1679);
or U2206 (N_2206,N_1668,N_1214);
nor U2207 (N_2207,N_1317,N_1690);
or U2208 (N_2208,N_1575,N_1636);
or U2209 (N_2209,N_1622,N_1205);
and U2210 (N_2210,N_1405,N_1444);
nor U2211 (N_2211,N_1721,N_1774);
nor U2212 (N_2212,N_1558,N_1773);
nor U2213 (N_2213,N_1620,N_1417);
nand U2214 (N_2214,N_1760,N_1399);
nor U2215 (N_2215,N_1368,N_1544);
nor U2216 (N_2216,N_1793,N_1657);
nand U2217 (N_2217,N_1445,N_1300);
and U2218 (N_2218,N_1300,N_1465);
nor U2219 (N_2219,N_1588,N_1732);
nand U2220 (N_2220,N_1392,N_1228);
or U2221 (N_2221,N_1482,N_1629);
and U2222 (N_2222,N_1690,N_1481);
nor U2223 (N_2223,N_1745,N_1578);
and U2224 (N_2224,N_1530,N_1583);
and U2225 (N_2225,N_1389,N_1645);
and U2226 (N_2226,N_1775,N_1457);
nand U2227 (N_2227,N_1304,N_1742);
nand U2228 (N_2228,N_1455,N_1515);
and U2229 (N_2229,N_1627,N_1503);
nand U2230 (N_2230,N_1399,N_1221);
xor U2231 (N_2231,N_1411,N_1456);
and U2232 (N_2232,N_1684,N_1751);
and U2233 (N_2233,N_1638,N_1205);
nand U2234 (N_2234,N_1372,N_1716);
nand U2235 (N_2235,N_1407,N_1576);
nor U2236 (N_2236,N_1606,N_1470);
or U2237 (N_2237,N_1473,N_1338);
or U2238 (N_2238,N_1232,N_1731);
or U2239 (N_2239,N_1776,N_1779);
nand U2240 (N_2240,N_1567,N_1649);
and U2241 (N_2241,N_1623,N_1241);
nand U2242 (N_2242,N_1716,N_1444);
nand U2243 (N_2243,N_1776,N_1313);
nor U2244 (N_2244,N_1489,N_1714);
or U2245 (N_2245,N_1712,N_1452);
xor U2246 (N_2246,N_1640,N_1517);
and U2247 (N_2247,N_1403,N_1749);
and U2248 (N_2248,N_1374,N_1520);
nor U2249 (N_2249,N_1456,N_1308);
and U2250 (N_2250,N_1505,N_1537);
nor U2251 (N_2251,N_1609,N_1288);
and U2252 (N_2252,N_1426,N_1535);
nand U2253 (N_2253,N_1381,N_1491);
and U2254 (N_2254,N_1708,N_1538);
nor U2255 (N_2255,N_1403,N_1717);
nor U2256 (N_2256,N_1430,N_1628);
and U2257 (N_2257,N_1324,N_1322);
and U2258 (N_2258,N_1489,N_1773);
or U2259 (N_2259,N_1699,N_1345);
and U2260 (N_2260,N_1598,N_1333);
or U2261 (N_2261,N_1370,N_1301);
and U2262 (N_2262,N_1444,N_1671);
nand U2263 (N_2263,N_1710,N_1695);
and U2264 (N_2264,N_1358,N_1450);
nand U2265 (N_2265,N_1467,N_1376);
xnor U2266 (N_2266,N_1225,N_1690);
and U2267 (N_2267,N_1235,N_1301);
nand U2268 (N_2268,N_1332,N_1567);
nand U2269 (N_2269,N_1775,N_1759);
or U2270 (N_2270,N_1696,N_1570);
nor U2271 (N_2271,N_1709,N_1481);
nor U2272 (N_2272,N_1383,N_1540);
nor U2273 (N_2273,N_1611,N_1754);
nor U2274 (N_2274,N_1700,N_1470);
nand U2275 (N_2275,N_1692,N_1736);
and U2276 (N_2276,N_1569,N_1577);
or U2277 (N_2277,N_1414,N_1784);
nand U2278 (N_2278,N_1238,N_1372);
nand U2279 (N_2279,N_1271,N_1525);
and U2280 (N_2280,N_1613,N_1202);
and U2281 (N_2281,N_1207,N_1429);
nand U2282 (N_2282,N_1665,N_1491);
and U2283 (N_2283,N_1724,N_1382);
and U2284 (N_2284,N_1545,N_1329);
and U2285 (N_2285,N_1786,N_1517);
or U2286 (N_2286,N_1422,N_1632);
nor U2287 (N_2287,N_1737,N_1640);
or U2288 (N_2288,N_1436,N_1747);
nand U2289 (N_2289,N_1397,N_1792);
nand U2290 (N_2290,N_1705,N_1623);
nand U2291 (N_2291,N_1642,N_1472);
nand U2292 (N_2292,N_1240,N_1339);
and U2293 (N_2293,N_1559,N_1535);
or U2294 (N_2294,N_1650,N_1483);
or U2295 (N_2295,N_1450,N_1793);
nor U2296 (N_2296,N_1692,N_1446);
nor U2297 (N_2297,N_1272,N_1252);
nand U2298 (N_2298,N_1499,N_1645);
nand U2299 (N_2299,N_1317,N_1693);
and U2300 (N_2300,N_1551,N_1508);
and U2301 (N_2301,N_1518,N_1396);
and U2302 (N_2302,N_1432,N_1561);
or U2303 (N_2303,N_1342,N_1523);
and U2304 (N_2304,N_1654,N_1658);
nand U2305 (N_2305,N_1410,N_1217);
or U2306 (N_2306,N_1648,N_1282);
or U2307 (N_2307,N_1384,N_1574);
nor U2308 (N_2308,N_1218,N_1594);
and U2309 (N_2309,N_1388,N_1228);
nor U2310 (N_2310,N_1594,N_1572);
or U2311 (N_2311,N_1344,N_1306);
xor U2312 (N_2312,N_1720,N_1650);
or U2313 (N_2313,N_1787,N_1400);
or U2314 (N_2314,N_1645,N_1644);
or U2315 (N_2315,N_1599,N_1393);
and U2316 (N_2316,N_1364,N_1546);
or U2317 (N_2317,N_1410,N_1250);
or U2318 (N_2318,N_1791,N_1510);
or U2319 (N_2319,N_1377,N_1355);
nor U2320 (N_2320,N_1437,N_1560);
nand U2321 (N_2321,N_1346,N_1695);
nand U2322 (N_2322,N_1639,N_1426);
or U2323 (N_2323,N_1450,N_1544);
nand U2324 (N_2324,N_1234,N_1585);
nand U2325 (N_2325,N_1658,N_1661);
nand U2326 (N_2326,N_1656,N_1255);
nand U2327 (N_2327,N_1592,N_1791);
and U2328 (N_2328,N_1423,N_1334);
and U2329 (N_2329,N_1266,N_1616);
and U2330 (N_2330,N_1722,N_1210);
nor U2331 (N_2331,N_1789,N_1747);
and U2332 (N_2332,N_1245,N_1648);
nand U2333 (N_2333,N_1468,N_1435);
nor U2334 (N_2334,N_1479,N_1400);
nor U2335 (N_2335,N_1759,N_1799);
and U2336 (N_2336,N_1786,N_1667);
nand U2337 (N_2337,N_1765,N_1399);
or U2338 (N_2338,N_1600,N_1276);
or U2339 (N_2339,N_1533,N_1569);
and U2340 (N_2340,N_1668,N_1256);
or U2341 (N_2341,N_1501,N_1300);
nand U2342 (N_2342,N_1595,N_1421);
nor U2343 (N_2343,N_1609,N_1593);
nor U2344 (N_2344,N_1447,N_1621);
and U2345 (N_2345,N_1353,N_1432);
or U2346 (N_2346,N_1637,N_1787);
and U2347 (N_2347,N_1427,N_1446);
nand U2348 (N_2348,N_1608,N_1581);
nand U2349 (N_2349,N_1429,N_1593);
nor U2350 (N_2350,N_1733,N_1405);
and U2351 (N_2351,N_1217,N_1720);
xnor U2352 (N_2352,N_1638,N_1639);
nor U2353 (N_2353,N_1738,N_1565);
or U2354 (N_2354,N_1410,N_1404);
or U2355 (N_2355,N_1622,N_1392);
and U2356 (N_2356,N_1666,N_1303);
and U2357 (N_2357,N_1301,N_1237);
or U2358 (N_2358,N_1583,N_1533);
nand U2359 (N_2359,N_1450,N_1751);
nand U2360 (N_2360,N_1748,N_1229);
or U2361 (N_2361,N_1631,N_1286);
xnor U2362 (N_2362,N_1737,N_1730);
nor U2363 (N_2363,N_1442,N_1236);
nand U2364 (N_2364,N_1457,N_1614);
or U2365 (N_2365,N_1444,N_1735);
nand U2366 (N_2366,N_1738,N_1755);
or U2367 (N_2367,N_1756,N_1390);
nand U2368 (N_2368,N_1345,N_1410);
and U2369 (N_2369,N_1243,N_1713);
nand U2370 (N_2370,N_1423,N_1275);
and U2371 (N_2371,N_1658,N_1413);
and U2372 (N_2372,N_1451,N_1334);
xor U2373 (N_2373,N_1619,N_1516);
and U2374 (N_2374,N_1553,N_1686);
or U2375 (N_2375,N_1311,N_1271);
or U2376 (N_2376,N_1355,N_1606);
nor U2377 (N_2377,N_1573,N_1499);
or U2378 (N_2378,N_1415,N_1222);
nor U2379 (N_2379,N_1628,N_1761);
or U2380 (N_2380,N_1325,N_1295);
nor U2381 (N_2381,N_1281,N_1220);
nand U2382 (N_2382,N_1766,N_1400);
or U2383 (N_2383,N_1658,N_1499);
and U2384 (N_2384,N_1315,N_1332);
nor U2385 (N_2385,N_1427,N_1675);
or U2386 (N_2386,N_1391,N_1749);
or U2387 (N_2387,N_1427,N_1496);
nand U2388 (N_2388,N_1362,N_1705);
or U2389 (N_2389,N_1612,N_1348);
nand U2390 (N_2390,N_1582,N_1469);
or U2391 (N_2391,N_1366,N_1226);
or U2392 (N_2392,N_1748,N_1581);
nor U2393 (N_2393,N_1632,N_1445);
or U2394 (N_2394,N_1461,N_1789);
nor U2395 (N_2395,N_1793,N_1492);
nand U2396 (N_2396,N_1216,N_1639);
and U2397 (N_2397,N_1298,N_1260);
xor U2398 (N_2398,N_1443,N_1271);
and U2399 (N_2399,N_1580,N_1406);
nand U2400 (N_2400,N_2023,N_2302);
and U2401 (N_2401,N_2055,N_2300);
and U2402 (N_2402,N_2316,N_1918);
nor U2403 (N_2403,N_1899,N_1934);
nor U2404 (N_2404,N_2178,N_1915);
or U2405 (N_2405,N_1879,N_2298);
or U2406 (N_2406,N_2326,N_2174);
or U2407 (N_2407,N_2371,N_1809);
and U2408 (N_2408,N_1895,N_2160);
or U2409 (N_2409,N_2012,N_2346);
or U2410 (N_2410,N_1960,N_1803);
nand U2411 (N_2411,N_2170,N_2111);
nand U2412 (N_2412,N_2365,N_1961);
nand U2413 (N_2413,N_2325,N_2275);
nor U2414 (N_2414,N_2211,N_1976);
nor U2415 (N_2415,N_1945,N_2212);
and U2416 (N_2416,N_2051,N_1812);
and U2417 (N_2417,N_2224,N_2279);
or U2418 (N_2418,N_2022,N_1862);
nor U2419 (N_2419,N_1957,N_1848);
nand U2420 (N_2420,N_2353,N_1914);
nor U2421 (N_2421,N_1996,N_2159);
nor U2422 (N_2422,N_2031,N_2216);
or U2423 (N_2423,N_2167,N_2054);
and U2424 (N_2424,N_1906,N_2362);
or U2425 (N_2425,N_1837,N_1897);
nor U2426 (N_2426,N_2359,N_1890);
nor U2427 (N_2427,N_2336,N_2273);
and U2428 (N_2428,N_1911,N_2120);
or U2429 (N_2429,N_1875,N_2377);
nor U2430 (N_2430,N_2204,N_2315);
and U2431 (N_2431,N_1968,N_2002);
nand U2432 (N_2432,N_2364,N_2009);
nand U2433 (N_2433,N_2322,N_2102);
or U2434 (N_2434,N_2208,N_2263);
and U2435 (N_2435,N_2114,N_1905);
nand U2436 (N_2436,N_2147,N_1807);
nor U2437 (N_2437,N_1988,N_2317);
and U2438 (N_2438,N_1815,N_2179);
and U2439 (N_2439,N_2343,N_2255);
or U2440 (N_2440,N_2324,N_1943);
nor U2441 (N_2441,N_2063,N_2245);
nand U2442 (N_2442,N_2184,N_2376);
or U2443 (N_2443,N_2235,N_2254);
or U2444 (N_2444,N_2121,N_1922);
nor U2445 (N_2445,N_2073,N_2360);
nor U2446 (N_2446,N_1978,N_1883);
nand U2447 (N_2447,N_2194,N_2161);
xnor U2448 (N_2448,N_2189,N_2248);
and U2449 (N_2449,N_2110,N_2366);
nor U2450 (N_2450,N_2112,N_2361);
nand U2451 (N_2451,N_2039,N_1871);
and U2452 (N_2452,N_1937,N_2020);
or U2453 (N_2453,N_2086,N_2210);
or U2454 (N_2454,N_1884,N_2152);
or U2455 (N_2455,N_2081,N_1924);
or U2456 (N_2456,N_2129,N_1855);
or U2457 (N_2457,N_2043,N_2265);
nand U2458 (N_2458,N_1912,N_1870);
and U2459 (N_2459,N_1965,N_2187);
nand U2460 (N_2460,N_2010,N_1808);
nor U2461 (N_2461,N_2383,N_2100);
or U2462 (N_2462,N_2358,N_2215);
nand U2463 (N_2463,N_2146,N_2270);
nand U2464 (N_2464,N_2319,N_2027);
or U2465 (N_2465,N_2108,N_2278);
and U2466 (N_2466,N_1834,N_2250);
nand U2467 (N_2467,N_2351,N_1856);
nand U2468 (N_2468,N_2028,N_1810);
or U2469 (N_2469,N_1923,N_1865);
nor U2470 (N_2470,N_2374,N_2091);
nand U2471 (N_2471,N_1970,N_2140);
xor U2472 (N_2472,N_2075,N_1824);
and U2473 (N_2473,N_2378,N_1946);
and U2474 (N_2474,N_2149,N_1839);
nand U2475 (N_2475,N_2329,N_2069);
or U2476 (N_2476,N_2045,N_1830);
nor U2477 (N_2477,N_2372,N_1832);
nor U2478 (N_2478,N_2044,N_1847);
nor U2479 (N_2479,N_2084,N_2180);
or U2480 (N_2480,N_2172,N_2328);
or U2481 (N_2481,N_2087,N_2192);
and U2482 (N_2482,N_2274,N_2037);
or U2483 (N_2483,N_1902,N_1880);
nand U2484 (N_2484,N_2201,N_1829);
nand U2485 (N_2485,N_2320,N_2017);
nand U2486 (N_2486,N_1938,N_2284);
or U2487 (N_2487,N_2134,N_2330);
or U2488 (N_2488,N_1842,N_2218);
nor U2489 (N_2489,N_2107,N_1941);
nor U2490 (N_2490,N_1853,N_2082);
or U2491 (N_2491,N_2321,N_1985);
nor U2492 (N_2492,N_2047,N_2025);
and U2493 (N_2493,N_2234,N_2391);
nand U2494 (N_2494,N_2034,N_2005);
nand U2495 (N_2495,N_1944,N_2079);
nand U2496 (N_2496,N_2150,N_1995);
or U2497 (N_2497,N_1889,N_1826);
nor U2498 (N_2498,N_1953,N_2006);
nor U2499 (N_2499,N_2390,N_2141);
or U2500 (N_2500,N_1981,N_1999);
nor U2501 (N_2501,N_2199,N_2165);
nor U2502 (N_2502,N_1949,N_1958);
nor U2503 (N_2503,N_2223,N_2264);
nand U2504 (N_2504,N_1989,N_2356);
nor U2505 (N_2505,N_1869,N_2342);
nor U2506 (N_2506,N_2058,N_1909);
nand U2507 (N_2507,N_2029,N_1992);
or U2508 (N_2508,N_2318,N_2038);
or U2509 (N_2509,N_2389,N_2333);
and U2510 (N_2510,N_1823,N_2231);
nand U2511 (N_2511,N_2209,N_1919);
or U2512 (N_2512,N_2222,N_1936);
and U2513 (N_2513,N_2276,N_2345);
nor U2514 (N_2514,N_2296,N_2239);
nand U2515 (N_2515,N_1952,N_2357);
nand U2516 (N_2516,N_2185,N_2243);
and U2517 (N_2517,N_2143,N_2387);
or U2518 (N_2518,N_2236,N_2132);
nor U2519 (N_2519,N_2203,N_2094);
or U2520 (N_2520,N_1888,N_2097);
and U2521 (N_2521,N_2313,N_2188);
or U2522 (N_2522,N_2101,N_2042);
nand U2523 (N_2523,N_2238,N_2018);
nor U2524 (N_2524,N_2092,N_2327);
and U2525 (N_2525,N_2397,N_2013);
nand U2526 (N_2526,N_2065,N_2220);
and U2527 (N_2527,N_1857,N_1959);
or U2528 (N_2528,N_1866,N_2256);
nor U2529 (N_2529,N_2303,N_2059);
and U2530 (N_2530,N_2154,N_1802);
nor U2531 (N_2531,N_2335,N_1963);
or U2532 (N_2532,N_1872,N_1806);
nand U2533 (N_2533,N_1966,N_2289);
nor U2534 (N_2534,N_2261,N_2145);
and U2535 (N_2535,N_2014,N_2016);
nand U2536 (N_2536,N_2190,N_2214);
nand U2537 (N_2537,N_2287,N_2370);
and U2538 (N_2538,N_1825,N_2341);
nor U2539 (N_2539,N_2367,N_1930);
or U2540 (N_2540,N_2118,N_2206);
and U2541 (N_2541,N_1878,N_2375);
nand U2542 (N_2542,N_2021,N_2309);
or U2543 (N_2543,N_2237,N_2127);
nand U2544 (N_2544,N_1813,N_2380);
nand U2545 (N_2545,N_2306,N_2153);
or U2546 (N_2546,N_1898,N_1851);
or U2547 (N_2547,N_2252,N_1972);
xnor U2548 (N_2548,N_1986,N_2177);
nand U2549 (N_2549,N_2057,N_2019);
or U2550 (N_2550,N_1836,N_2080);
xor U2551 (N_2551,N_1892,N_2048);
nand U2552 (N_2552,N_1877,N_1843);
and U2553 (N_2553,N_2314,N_2007);
and U2554 (N_2554,N_1935,N_1971);
nor U2555 (N_2555,N_1967,N_2137);
and U2556 (N_2556,N_2297,N_2003);
nand U2557 (N_2557,N_2219,N_1840);
and U2558 (N_2558,N_1983,N_2310);
nand U2559 (N_2559,N_2136,N_1821);
nor U2560 (N_2560,N_2379,N_1954);
or U2561 (N_2561,N_2156,N_2354);
nor U2562 (N_2562,N_1801,N_2240);
nor U2563 (N_2563,N_2163,N_2304);
and U2564 (N_2564,N_2227,N_2171);
and U2565 (N_2565,N_1916,N_1849);
nor U2566 (N_2566,N_1881,N_1841);
nand U2567 (N_2567,N_1833,N_2392);
xnor U2568 (N_2568,N_2259,N_2077);
and U2569 (N_2569,N_2035,N_1827);
nor U2570 (N_2570,N_2186,N_2133);
xnor U2571 (N_2571,N_2125,N_1928);
and U2572 (N_2572,N_2232,N_2226);
nand U2573 (N_2573,N_1800,N_1858);
nand U2574 (N_2574,N_2001,N_2126);
and U2575 (N_2575,N_2229,N_2083);
or U2576 (N_2576,N_2205,N_2332);
and U2577 (N_2577,N_1868,N_1926);
or U2578 (N_2578,N_2244,N_2228);
nor U2579 (N_2579,N_1993,N_2338);
nand U2580 (N_2580,N_1901,N_2288);
nand U2581 (N_2581,N_2225,N_2036);
or U2582 (N_2582,N_2266,N_1850);
and U2583 (N_2583,N_1876,N_2040);
nor U2584 (N_2584,N_1974,N_2130);
and U2585 (N_2585,N_1817,N_1900);
nor U2586 (N_2586,N_1859,N_2337);
xor U2587 (N_2587,N_1882,N_1844);
nor U2588 (N_2588,N_1863,N_2307);
and U2589 (N_2589,N_1907,N_1997);
and U2590 (N_2590,N_1927,N_1894);
nand U2591 (N_2591,N_2271,N_1933);
or U2592 (N_2592,N_1964,N_1908);
or U2593 (N_2593,N_2061,N_2066);
or U2594 (N_2594,N_2071,N_2363);
nand U2595 (N_2595,N_2116,N_2246);
or U2596 (N_2596,N_2060,N_1893);
and U2597 (N_2597,N_2122,N_2000);
nand U2598 (N_2598,N_1835,N_2340);
and U2599 (N_2599,N_2308,N_2384);
nor U2600 (N_2600,N_2202,N_2024);
nor U2601 (N_2601,N_2368,N_2272);
or U2602 (N_2602,N_2088,N_1860);
nor U2603 (N_2603,N_2323,N_2249);
nand U2604 (N_2604,N_2182,N_2056);
and U2605 (N_2605,N_2128,N_2176);
and U2606 (N_2606,N_2350,N_2173);
nor U2607 (N_2607,N_1925,N_2241);
nor U2608 (N_2608,N_2193,N_2280);
or U2609 (N_2609,N_1805,N_1948);
nand U2610 (N_2610,N_1984,N_1987);
or U2611 (N_2611,N_2242,N_1921);
nor U2612 (N_2612,N_2181,N_2217);
nand U2613 (N_2613,N_2334,N_2033);
nand U2614 (N_2614,N_2262,N_1816);
nor U2615 (N_2615,N_2292,N_1913);
and U2616 (N_2616,N_1982,N_1940);
and U2617 (N_2617,N_2183,N_2131);
nand U2618 (N_2618,N_2089,N_2169);
and U2619 (N_2619,N_2098,N_2074);
nand U2620 (N_2620,N_2339,N_2299);
or U2621 (N_2621,N_2195,N_1956);
nand U2622 (N_2622,N_2026,N_2049);
nor U2623 (N_2623,N_1929,N_2119);
nand U2624 (N_2624,N_1979,N_1854);
nand U2625 (N_2625,N_2115,N_2197);
or U2626 (N_2626,N_1874,N_2164);
or U2627 (N_2627,N_2344,N_2162);
and U2628 (N_2628,N_1962,N_2157);
and U2629 (N_2629,N_2293,N_2200);
nand U2630 (N_2630,N_2070,N_2064);
nor U2631 (N_2631,N_2175,N_2247);
nor U2632 (N_2632,N_2004,N_2155);
nand U2633 (N_2633,N_1820,N_2233);
and U2634 (N_2634,N_2294,N_1819);
nor U2635 (N_2635,N_1811,N_1885);
xor U2636 (N_2636,N_2076,N_2139);
and U2637 (N_2637,N_2369,N_2277);
and U2638 (N_2638,N_2103,N_1994);
nor U2639 (N_2639,N_2085,N_2046);
or U2640 (N_2640,N_2381,N_2396);
nor U2641 (N_2641,N_1977,N_1822);
nor U2642 (N_2642,N_1951,N_2373);
and U2643 (N_2643,N_1861,N_2386);
and U2644 (N_2644,N_2078,N_2251);
or U2645 (N_2645,N_2305,N_1939);
nand U2646 (N_2646,N_1991,N_2267);
nor U2647 (N_2647,N_1804,N_1998);
or U2648 (N_2648,N_2258,N_1814);
or U2649 (N_2649,N_2388,N_2311);
and U2650 (N_2650,N_2269,N_2158);
nor U2651 (N_2651,N_1980,N_2191);
nor U2652 (N_2652,N_1932,N_1886);
nand U2653 (N_2653,N_2090,N_2260);
or U2654 (N_2654,N_2253,N_2124);
nand U2655 (N_2655,N_2072,N_2291);
nand U2656 (N_2656,N_1867,N_1990);
nand U2657 (N_2657,N_2382,N_1864);
and U2658 (N_2658,N_1903,N_2398);
and U2659 (N_2659,N_2331,N_2295);
or U2660 (N_2660,N_1942,N_2301);
or U2661 (N_2661,N_1845,N_2104);
and U2662 (N_2662,N_2062,N_2352);
or U2663 (N_2663,N_2347,N_2008);
nor U2664 (N_2664,N_1910,N_2283);
nor U2665 (N_2665,N_2168,N_2067);
or U2666 (N_2666,N_2394,N_2138);
and U2667 (N_2667,N_2011,N_1887);
xor U2668 (N_2668,N_2151,N_2105);
and U2669 (N_2669,N_2095,N_1896);
nand U2670 (N_2670,N_2096,N_1920);
nand U2671 (N_2671,N_2257,N_2015);
or U2672 (N_2672,N_2312,N_2053);
or U2673 (N_2673,N_2221,N_2385);
and U2674 (N_2674,N_2068,N_2030);
nand U2675 (N_2675,N_2281,N_1975);
nand U2676 (N_2676,N_2268,N_2399);
and U2677 (N_2677,N_1828,N_2213);
or U2678 (N_2678,N_2050,N_1950);
xnor U2679 (N_2679,N_1846,N_2106);
or U2680 (N_2680,N_2282,N_1947);
or U2681 (N_2681,N_2395,N_2198);
nand U2682 (N_2682,N_2286,N_2393);
nand U2683 (N_2683,N_2113,N_1838);
nand U2684 (N_2684,N_1904,N_1955);
nor U2685 (N_2685,N_2207,N_2142);
or U2686 (N_2686,N_2285,N_2117);
xnor U2687 (N_2687,N_2148,N_1973);
nand U2688 (N_2688,N_2052,N_2109);
nand U2689 (N_2689,N_2123,N_2348);
and U2690 (N_2690,N_1852,N_2032);
nor U2691 (N_2691,N_1818,N_2355);
or U2692 (N_2692,N_1969,N_1891);
nor U2693 (N_2693,N_2349,N_1931);
nand U2694 (N_2694,N_1873,N_2196);
nor U2695 (N_2695,N_2041,N_2099);
nor U2696 (N_2696,N_2093,N_2135);
or U2697 (N_2697,N_2166,N_2144);
and U2698 (N_2698,N_1917,N_1831);
nor U2699 (N_2699,N_2290,N_2230);
nand U2700 (N_2700,N_1943,N_2073);
or U2701 (N_2701,N_2316,N_1879);
or U2702 (N_2702,N_1937,N_2307);
and U2703 (N_2703,N_2161,N_1943);
or U2704 (N_2704,N_1891,N_1956);
and U2705 (N_2705,N_1900,N_1939);
nor U2706 (N_2706,N_2249,N_2111);
nand U2707 (N_2707,N_1916,N_1833);
and U2708 (N_2708,N_1931,N_1961);
nand U2709 (N_2709,N_2264,N_2049);
or U2710 (N_2710,N_2090,N_1885);
nand U2711 (N_2711,N_1886,N_1910);
and U2712 (N_2712,N_2225,N_2372);
nor U2713 (N_2713,N_1846,N_2060);
nor U2714 (N_2714,N_2394,N_2271);
and U2715 (N_2715,N_1950,N_2231);
nand U2716 (N_2716,N_2143,N_2295);
and U2717 (N_2717,N_2193,N_2005);
or U2718 (N_2718,N_1958,N_1889);
xor U2719 (N_2719,N_1807,N_1870);
nand U2720 (N_2720,N_2210,N_2155);
nor U2721 (N_2721,N_2119,N_2319);
nand U2722 (N_2722,N_1817,N_2013);
nor U2723 (N_2723,N_2060,N_1875);
nor U2724 (N_2724,N_1811,N_1958);
or U2725 (N_2725,N_1894,N_1851);
and U2726 (N_2726,N_2131,N_2208);
nand U2727 (N_2727,N_2081,N_2379);
nor U2728 (N_2728,N_2023,N_1862);
or U2729 (N_2729,N_2096,N_2097);
xnor U2730 (N_2730,N_1921,N_2392);
nand U2731 (N_2731,N_2014,N_1883);
nor U2732 (N_2732,N_1870,N_2012);
and U2733 (N_2733,N_2081,N_1995);
nor U2734 (N_2734,N_2121,N_2186);
nand U2735 (N_2735,N_1962,N_2253);
or U2736 (N_2736,N_2128,N_2056);
nand U2737 (N_2737,N_1865,N_2297);
and U2738 (N_2738,N_2121,N_2003);
nand U2739 (N_2739,N_1986,N_2011);
and U2740 (N_2740,N_2289,N_2139);
nor U2741 (N_2741,N_1903,N_2335);
and U2742 (N_2742,N_2317,N_2305);
nor U2743 (N_2743,N_2051,N_2103);
nor U2744 (N_2744,N_2379,N_1879);
and U2745 (N_2745,N_2009,N_1945);
and U2746 (N_2746,N_2377,N_2203);
and U2747 (N_2747,N_1938,N_1835);
and U2748 (N_2748,N_2287,N_1872);
and U2749 (N_2749,N_1956,N_2118);
and U2750 (N_2750,N_2255,N_2176);
nand U2751 (N_2751,N_2282,N_2129);
and U2752 (N_2752,N_2097,N_1893);
and U2753 (N_2753,N_2044,N_2314);
nand U2754 (N_2754,N_1982,N_2001);
or U2755 (N_2755,N_2263,N_1884);
and U2756 (N_2756,N_1918,N_2307);
and U2757 (N_2757,N_2134,N_1857);
and U2758 (N_2758,N_2194,N_2293);
or U2759 (N_2759,N_2190,N_2238);
nor U2760 (N_2760,N_2121,N_2154);
xnor U2761 (N_2761,N_2351,N_2347);
or U2762 (N_2762,N_2302,N_2149);
and U2763 (N_2763,N_2304,N_2003);
and U2764 (N_2764,N_2294,N_2365);
nand U2765 (N_2765,N_2163,N_1851);
nand U2766 (N_2766,N_2028,N_2277);
or U2767 (N_2767,N_2020,N_1800);
nor U2768 (N_2768,N_1960,N_2050);
nor U2769 (N_2769,N_2387,N_2091);
and U2770 (N_2770,N_2324,N_2070);
nand U2771 (N_2771,N_1845,N_1904);
and U2772 (N_2772,N_1953,N_2227);
or U2773 (N_2773,N_2380,N_1806);
or U2774 (N_2774,N_2180,N_2354);
nand U2775 (N_2775,N_2388,N_1816);
or U2776 (N_2776,N_2374,N_2193);
nor U2777 (N_2777,N_2000,N_1919);
or U2778 (N_2778,N_2228,N_2366);
nand U2779 (N_2779,N_2256,N_1953);
nor U2780 (N_2780,N_2256,N_1957);
nand U2781 (N_2781,N_2178,N_2395);
nand U2782 (N_2782,N_2344,N_2345);
and U2783 (N_2783,N_2245,N_1815);
and U2784 (N_2784,N_2118,N_2023);
nor U2785 (N_2785,N_2252,N_2263);
nor U2786 (N_2786,N_2329,N_2269);
or U2787 (N_2787,N_2133,N_2180);
nor U2788 (N_2788,N_2127,N_2057);
and U2789 (N_2789,N_1853,N_2358);
or U2790 (N_2790,N_2314,N_2295);
nand U2791 (N_2791,N_2375,N_1933);
and U2792 (N_2792,N_2253,N_1801);
nor U2793 (N_2793,N_2311,N_1946);
nor U2794 (N_2794,N_1969,N_2183);
or U2795 (N_2795,N_2333,N_2275);
nor U2796 (N_2796,N_2298,N_2094);
and U2797 (N_2797,N_2166,N_2013);
nand U2798 (N_2798,N_2333,N_2353);
and U2799 (N_2799,N_2245,N_2184);
and U2800 (N_2800,N_2396,N_1912);
nor U2801 (N_2801,N_2309,N_2025);
nand U2802 (N_2802,N_1900,N_1933);
nor U2803 (N_2803,N_2369,N_2093);
or U2804 (N_2804,N_1962,N_2130);
nor U2805 (N_2805,N_1953,N_2269);
and U2806 (N_2806,N_2381,N_2183);
nand U2807 (N_2807,N_2104,N_1973);
or U2808 (N_2808,N_2059,N_2148);
nand U2809 (N_2809,N_2282,N_1871);
nor U2810 (N_2810,N_2138,N_2099);
nand U2811 (N_2811,N_1867,N_2302);
and U2812 (N_2812,N_1982,N_2090);
or U2813 (N_2813,N_1925,N_2373);
nand U2814 (N_2814,N_2306,N_2108);
nand U2815 (N_2815,N_2211,N_1921);
or U2816 (N_2816,N_2163,N_2204);
or U2817 (N_2817,N_1812,N_1860);
or U2818 (N_2818,N_2365,N_1832);
nor U2819 (N_2819,N_1895,N_2385);
and U2820 (N_2820,N_1850,N_2330);
nor U2821 (N_2821,N_2246,N_2085);
and U2822 (N_2822,N_1818,N_2134);
nor U2823 (N_2823,N_2285,N_2288);
nand U2824 (N_2824,N_2034,N_2370);
or U2825 (N_2825,N_1969,N_2115);
nand U2826 (N_2826,N_1812,N_1909);
nor U2827 (N_2827,N_1993,N_1922);
or U2828 (N_2828,N_1809,N_1864);
and U2829 (N_2829,N_2340,N_2158);
or U2830 (N_2830,N_2334,N_2288);
nor U2831 (N_2831,N_2110,N_1998);
nand U2832 (N_2832,N_1830,N_1836);
or U2833 (N_2833,N_1981,N_2261);
nor U2834 (N_2834,N_2142,N_2070);
or U2835 (N_2835,N_2317,N_2241);
nand U2836 (N_2836,N_2255,N_1908);
nor U2837 (N_2837,N_2056,N_2127);
and U2838 (N_2838,N_2363,N_2313);
and U2839 (N_2839,N_2287,N_1901);
nor U2840 (N_2840,N_2157,N_2283);
xor U2841 (N_2841,N_1831,N_1955);
nor U2842 (N_2842,N_2249,N_2338);
nor U2843 (N_2843,N_1867,N_2193);
nor U2844 (N_2844,N_1823,N_1956);
and U2845 (N_2845,N_1837,N_2160);
nand U2846 (N_2846,N_2115,N_2232);
or U2847 (N_2847,N_2156,N_2161);
nor U2848 (N_2848,N_2219,N_2314);
nand U2849 (N_2849,N_2079,N_1809);
or U2850 (N_2850,N_2067,N_2286);
and U2851 (N_2851,N_2149,N_2345);
and U2852 (N_2852,N_1853,N_2220);
nand U2853 (N_2853,N_1977,N_1931);
nor U2854 (N_2854,N_2239,N_2254);
or U2855 (N_2855,N_2349,N_2174);
and U2856 (N_2856,N_2345,N_2220);
or U2857 (N_2857,N_2024,N_1898);
or U2858 (N_2858,N_2272,N_1817);
nor U2859 (N_2859,N_2189,N_1943);
or U2860 (N_2860,N_2151,N_2037);
or U2861 (N_2861,N_1876,N_2303);
nand U2862 (N_2862,N_2074,N_1997);
nand U2863 (N_2863,N_2204,N_2245);
or U2864 (N_2864,N_2374,N_1877);
or U2865 (N_2865,N_2283,N_2063);
or U2866 (N_2866,N_2160,N_2047);
nand U2867 (N_2867,N_2337,N_2193);
or U2868 (N_2868,N_2364,N_1987);
nor U2869 (N_2869,N_2125,N_2051);
or U2870 (N_2870,N_2192,N_2371);
nor U2871 (N_2871,N_2340,N_2206);
or U2872 (N_2872,N_2309,N_2033);
nand U2873 (N_2873,N_1820,N_2330);
or U2874 (N_2874,N_2281,N_2106);
or U2875 (N_2875,N_2320,N_2329);
nand U2876 (N_2876,N_1972,N_2107);
or U2877 (N_2877,N_2076,N_2314);
and U2878 (N_2878,N_1978,N_1841);
and U2879 (N_2879,N_1971,N_1812);
or U2880 (N_2880,N_1802,N_2277);
nand U2881 (N_2881,N_2327,N_1810);
nand U2882 (N_2882,N_1856,N_1926);
nand U2883 (N_2883,N_2030,N_2201);
or U2884 (N_2884,N_2230,N_2112);
and U2885 (N_2885,N_2042,N_2125);
or U2886 (N_2886,N_2262,N_2070);
or U2887 (N_2887,N_2011,N_2320);
or U2888 (N_2888,N_1888,N_2283);
nand U2889 (N_2889,N_2365,N_1887);
nand U2890 (N_2890,N_1991,N_1918);
and U2891 (N_2891,N_2098,N_2360);
and U2892 (N_2892,N_1883,N_2196);
xnor U2893 (N_2893,N_2268,N_2296);
or U2894 (N_2894,N_2233,N_2174);
and U2895 (N_2895,N_1820,N_1844);
nor U2896 (N_2896,N_1804,N_2122);
nor U2897 (N_2897,N_2039,N_2048);
or U2898 (N_2898,N_1819,N_2127);
nand U2899 (N_2899,N_2183,N_1841);
or U2900 (N_2900,N_2393,N_2297);
nor U2901 (N_2901,N_1842,N_1937);
nand U2902 (N_2902,N_2234,N_1906);
nand U2903 (N_2903,N_2027,N_2174);
nor U2904 (N_2904,N_2047,N_1821);
nand U2905 (N_2905,N_2144,N_2108);
nand U2906 (N_2906,N_2266,N_2306);
and U2907 (N_2907,N_2120,N_1825);
nor U2908 (N_2908,N_2201,N_2262);
nor U2909 (N_2909,N_2033,N_1869);
nand U2910 (N_2910,N_1834,N_2317);
or U2911 (N_2911,N_1942,N_1833);
and U2912 (N_2912,N_2008,N_2250);
nor U2913 (N_2913,N_2047,N_2004);
and U2914 (N_2914,N_2271,N_2154);
and U2915 (N_2915,N_2399,N_1943);
and U2916 (N_2916,N_1967,N_2173);
nor U2917 (N_2917,N_1803,N_1908);
or U2918 (N_2918,N_1815,N_2320);
and U2919 (N_2919,N_2271,N_2372);
nor U2920 (N_2920,N_2243,N_1840);
and U2921 (N_2921,N_1868,N_1985);
nor U2922 (N_2922,N_2301,N_2331);
and U2923 (N_2923,N_2141,N_2041);
nor U2924 (N_2924,N_1850,N_1802);
nor U2925 (N_2925,N_2151,N_2009);
and U2926 (N_2926,N_2117,N_2303);
nor U2927 (N_2927,N_2354,N_2084);
xnor U2928 (N_2928,N_1967,N_1884);
and U2929 (N_2929,N_2316,N_2086);
nand U2930 (N_2930,N_1934,N_1884);
and U2931 (N_2931,N_1900,N_1929);
nand U2932 (N_2932,N_2152,N_2161);
and U2933 (N_2933,N_2352,N_2369);
xnor U2934 (N_2934,N_1861,N_2003);
xor U2935 (N_2935,N_1999,N_2199);
or U2936 (N_2936,N_2191,N_1968);
nand U2937 (N_2937,N_2160,N_2166);
nor U2938 (N_2938,N_2023,N_1881);
or U2939 (N_2939,N_2159,N_2316);
or U2940 (N_2940,N_1883,N_2074);
and U2941 (N_2941,N_1836,N_2215);
nor U2942 (N_2942,N_1939,N_2031);
nand U2943 (N_2943,N_1809,N_1960);
or U2944 (N_2944,N_2166,N_2168);
and U2945 (N_2945,N_2353,N_1988);
and U2946 (N_2946,N_2202,N_2261);
nand U2947 (N_2947,N_2176,N_2118);
and U2948 (N_2948,N_1872,N_2222);
or U2949 (N_2949,N_1877,N_2187);
nor U2950 (N_2950,N_2050,N_1871);
and U2951 (N_2951,N_2122,N_2344);
nand U2952 (N_2952,N_2087,N_2165);
or U2953 (N_2953,N_2001,N_2176);
xor U2954 (N_2954,N_2213,N_1858);
or U2955 (N_2955,N_1946,N_2362);
nor U2956 (N_2956,N_1934,N_2171);
and U2957 (N_2957,N_2088,N_2272);
or U2958 (N_2958,N_2368,N_2354);
and U2959 (N_2959,N_1980,N_2324);
nand U2960 (N_2960,N_2375,N_2295);
and U2961 (N_2961,N_2239,N_1850);
nand U2962 (N_2962,N_1969,N_2292);
and U2963 (N_2963,N_1994,N_2044);
or U2964 (N_2964,N_1931,N_2279);
nand U2965 (N_2965,N_2079,N_2338);
nand U2966 (N_2966,N_2375,N_2096);
and U2967 (N_2967,N_1908,N_2092);
and U2968 (N_2968,N_2222,N_2054);
and U2969 (N_2969,N_1822,N_2238);
nor U2970 (N_2970,N_2284,N_2392);
and U2971 (N_2971,N_1860,N_2321);
nor U2972 (N_2972,N_2207,N_2069);
or U2973 (N_2973,N_2023,N_1858);
nand U2974 (N_2974,N_2202,N_2219);
nor U2975 (N_2975,N_2118,N_2295);
nand U2976 (N_2976,N_2075,N_1809);
nor U2977 (N_2977,N_2100,N_2065);
nor U2978 (N_2978,N_2329,N_2145);
and U2979 (N_2979,N_2217,N_2085);
or U2980 (N_2980,N_2049,N_2268);
nor U2981 (N_2981,N_2114,N_2272);
or U2982 (N_2982,N_2149,N_1961);
nand U2983 (N_2983,N_2385,N_1884);
and U2984 (N_2984,N_2171,N_2243);
and U2985 (N_2985,N_1918,N_2265);
nand U2986 (N_2986,N_2134,N_2308);
nand U2987 (N_2987,N_1986,N_2152);
nor U2988 (N_2988,N_2361,N_1856);
and U2989 (N_2989,N_2191,N_2131);
nor U2990 (N_2990,N_2286,N_2371);
or U2991 (N_2991,N_2204,N_2213);
or U2992 (N_2992,N_2101,N_1925);
nand U2993 (N_2993,N_2248,N_2266);
nand U2994 (N_2994,N_1809,N_1973);
xnor U2995 (N_2995,N_2149,N_2215);
and U2996 (N_2996,N_1800,N_1977);
nand U2997 (N_2997,N_1923,N_2306);
nand U2998 (N_2998,N_2044,N_2204);
nand U2999 (N_2999,N_1975,N_1890);
and UO_0 (O_0,N_2456,N_2427);
xor UO_1 (O_1,N_2947,N_2508);
and UO_2 (O_2,N_2678,N_2664);
nor UO_3 (O_3,N_2729,N_2716);
nand UO_4 (O_4,N_2577,N_2615);
xnor UO_5 (O_5,N_2590,N_2932);
xor UO_6 (O_6,N_2765,N_2707);
or UO_7 (O_7,N_2694,N_2758);
or UO_8 (O_8,N_2500,N_2683);
xnor UO_9 (O_9,N_2816,N_2492);
or UO_10 (O_10,N_2679,N_2677);
or UO_11 (O_11,N_2647,N_2708);
nand UO_12 (O_12,N_2988,N_2878);
nand UO_13 (O_13,N_2790,N_2803);
and UO_14 (O_14,N_2489,N_2857);
and UO_15 (O_15,N_2888,N_2520);
nand UO_16 (O_16,N_2948,N_2566);
nor UO_17 (O_17,N_2778,N_2941);
nand UO_18 (O_18,N_2451,N_2616);
nor UO_19 (O_19,N_2513,N_2808);
nand UO_20 (O_20,N_2749,N_2518);
and UO_21 (O_21,N_2580,N_2735);
nor UO_22 (O_22,N_2632,N_2562);
or UO_23 (O_23,N_2732,N_2811);
or UO_24 (O_24,N_2424,N_2917);
xor UO_25 (O_25,N_2431,N_2969);
nand UO_26 (O_26,N_2416,N_2884);
or UO_27 (O_27,N_2859,N_2675);
nand UO_28 (O_28,N_2776,N_2463);
nor UO_29 (O_29,N_2497,N_2618);
nand UO_30 (O_30,N_2833,N_2641);
nor UO_31 (O_31,N_2505,N_2871);
and UO_32 (O_32,N_2959,N_2845);
xor UO_33 (O_33,N_2662,N_2648);
and UO_34 (O_34,N_2660,N_2759);
and UO_35 (O_35,N_2853,N_2982);
nand UO_36 (O_36,N_2402,N_2799);
nor UO_37 (O_37,N_2997,N_2980);
or UO_38 (O_38,N_2691,N_2401);
nor UO_39 (O_39,N_2529,N_2928);
nor UO_40 (O_40,N_2481,N_2898);
nor UO_41 (O_41,N_2530,N_2668);
nor UO_42 (O_42,N_2583,N_2432);
and UO_43 (O_43,N_2455,N_2835);
and UO_44 (O_44,N_2998,N_2830);
nor UO_45 (O_45,N_2957,N_2579);
nand UO_46 (O_46,N_2843,N_2686);
or UO_47 (O_47,N_2558,N_2512);
or UO_48 (O_48,N_2547,N_2659);
and UO_49 (O_49,N_2715,N_2796);
or UO_50 (O_50,N_2999,N_2777);
nor UO_51 (O_51,N_2847,N_2739);
xnor UO_52 (O_52,N_2990,N_2746);
or UO_53 (O_53,N_2541,N_2439);
or UO_54 (O_54,N_2960,N_2839);
nand UO_55 (O_55,N_2991,N_2755);
or UO_56 (O_56,N_2696,N_2996);
and UO_57 (O_57,N_2470,N_2719);
or UO_58 (O_58,N_2511,N_2464);
or UO_59 (O_59,N_2491,N_2544);
nor UO_60 (O_60,N_2929,N_2894);
and UO_61 (O_61,N_2435,N_2597);
nor UO_62 (O_62,N_2922,N_2901);
nor UO_63 (O_63,N_2724,N_2798);
nor UO_64 (O_64,N_2935,N_2426);
nor UO_65 (O_65,N_2567,N_2551);
and UO_66 (O_66,N_2542,N_2412);
or UO_67 (O_67,N_2961,N_2634);
nand UO_68 (O_68,N_2437,N_2587);
or UO_69 (O_69,N_2493,N_2419);
or UO_70 (O_70,N_2653,N_2625);
nor UO_71 (O_71,N_2697,N_2892);
and UO_72 (O_72,N_2975,N_2534);
and UO_73 (O_73,N_2767,N_2726);
nand UO_74 (O_74,N_2410,N_2594);
xor UO_75 (O_75,N_2779,N_2537);
nand UO_76 (O_76,N_2766,N_2768);
nand UO_77 (O_77,N_2971,N_2831);
nand UO_78 (O_78,N_2868,N_2501);
or UO_79 (O_79,N_2723,N_2797);
nand UO_80 (O_80,N_2494,N_2775);
nand UO_81 (O_81,N_2771,N_2792);
nand UO_82 (O_82,N_2731,N_2883);
or UO_83 (O_83,N_2822,N_2661);
nand UO_84 (O_84,N_2554,N_2930);
nand UO_85 (O_85,N_2946,N_2821);
or UO_86 (O_86,N_2612,N_2546);
nor UO_87 (O_87,N_2478,N_2667);
and UO_88 (O_88,N_2820,N_2896);
nand UO_89 (O_89,N_2860,N_2549);
or UO_90 (O_90,N_2890,N_2876);
nor UO_91 (O_91,N_2657,N_2858);
and UO_92 (O_92,N_2899,N_2571);
nand UO_93 (O_93,N_2656,N_2442);
or UO_94 (O_94,N_2962,N_2965);
nand UO_95 (O_95,N_2613,N_2469);
nor UO_96 (O_96,N_2944,N_2786);
and UO_97 (O_97,N_2411,N_2690);
or UO_98 (O_98,N_2815,N_2670);
nand UO_99 (O_99,N_2733,N_2563);
or UO_100 (O_100,N_2879,N_2606);
nand UO_101 (O_101,N_2842,N_2519);
and UO_102 (O_102,N_2800,N_2882);
nand UO_103 (O_103,N_2674,N_2573);
nor UO_104 (O_104,N_2744,N_2526);
nand UO_105 (O_105,N_2406,N_2807);
nor UO_106 (O_106,N_2806,N_2630);
nor UO_107 (O_107,N_2623,N_2599);
nand UO_108 (O_108,N_2963,N_2784);
and UO_109 (O_109,N_2742,N_2728);
nand UO_110 (O_110,N_2440,N_2722);
or UO_111 (O_111,N_2914,N_2408);
and UO_112 (O_112,N_2994,N_2730);
nor UO_113 (O_113,N_2918,N_2977);
and UO_114 (O_114,N_2757,N_2791);
and UO_115 (O_115,N_2923,N_2595);
nand UO_116 (O_116,N_2752,N_2569);
or UO_117 (O_117,N_2617,N_2507);
or UO_118 (O_118,N_2403,N_2450);
and UO_119 (O_119,N_2514,N_2480);
nor UO_120 (O_120,N_2976,N_2773);
nor UO_121 (O_121,N_2881,N_2684);
nor UO_122 (O_122,N_2651,N_2874);
nor UO_123 (O_123,N_2737,N_2958);
nor UO_124 (O_124,N_2655,N_2973);
or UO_125 (O_125,N_2702,N_2638);
nand UO_126 (O_126,N_2665,N_2885);
or UO_127 (O_127,N_2851,N_2578);
nor UO_128 (O_128,N_2772,N_2504);
nor UO_129 (O_129,N_2717,N_2433);
nand UO_130 (O_130,N_2666,N_2781);
nand UO_131 (O_131,N_2814,N_2747);
nand UO_132 (O_132,N_2785,N_2938);
and UO_133 (O_133,N_2591,N_2531);
or UO_134 (O_134,N_2624,N_2787);
or UO_135 (O_135,N_2693,N_2564);
nor UO_136 (O_136,N_2495,N_2951);
or UO_137 (O_137,N_2561,N_2966);
and UO_138 (O_138,N_2762,N_2704);
nor UO_139 (O_139,N_2940,N_2605);
and UO_140 (O_140,N_2793,N_2510);
and UO_141 (O_141,N_2636,N_2818);
and UO_142 (O_142,N_2650,N_2908);
or UO_143 (O_143,N_2925,N_2688);
nand UO_144 (O_144,N_2499,N_2872);
nand UO_145 (O_145,N_2837,N_2949);
or UO_146 (O_146,N_2956,N_2770);
or UO_147 (O_147,N_2886,N_2865);
and UO_148 (O_148,N_2409,N_2745);
xnor UO_149 (O_149,N_2600,N_2974);
nand UO_150 (O_150,N_2644,N_2407);
and UO_151 (O_151,N_2447,N_2490);
and UO_152 (O_152,N_2629,N_2671);
or UO_153 (O_153,N_2588,N_2673);
nand UO_154 (O_154,N_2453,N_2711);
nand UO_155 (O_155,N_2524,N_2698);
and UO_156 (O_156,N_2756,N_2841);
nor UO_157 (O_157,N_2610,N_2780);
nor UO_158 (O_158,N_2523,N_2596);
nand UO_159 (O_159,N_2483,N_2631);
and UO_160 (O_160,N_2795,N_2627);
and UO_161 (O_161,N_2642,N_2931);
nand UO_162 (O_162,N_2992,N_2515);
or UO_163 (O_163,N_2443,N_2718);
and UO_164 (O_164,N_2919,N_2856);
nor UO_165 (O_165,N_2895,N_2517);
or UO_166 (O_166,N_2414,N_2754);
or UO_167 (O_167,N_2829,N_2826);
nand UO_168 (O_168,N_2415,N_2875);
nand UO_169 (O_169,N_2533,N_2472);
and UO_170 (O_170,N_2989,N_2813);
nand UO_171 (O_171,N_2584,N_2911);
nand UO_172 (O_172,N_2474,N_2819);
nor UO_173 (O_173,N_2404,N_2788);
nor UO_174 (O_174,N_2713,N_2701);
and UO_175 (O_175,N_2903,N_2855);
nor UO_176 (O_176,N_2649,N_2984);
nand UO_177 (O_177,N_2710,N_2750);
nand UO_178 (O_178,N_2817,N_2676);
nand UO_179 (O_179,N_2769,N_2485);
or UO_180 (O_180,N_2457,N_2985);
nand UO_181 (O_181,N_2852,N_2942);
and UO_182 (O_182,N_2761,N_2425);
nand UO_183 (O_183,N_2748,N_2628);
nand UO_184 (O_184,N_2934,N_2905);
nor UO_185 (O_185,N_2699,N_2645);
and UO_186 (O_186,N_2421,N_2955);
and UO_187 (O_187,N_2565,N_2672);
or UO_188 (O_188,N_2794,N_2654);
and UO_189 (O_189,N_2446,N_2608);
or UO_190 (O_190,N_2950,N_2640);
nand UO_191 (O_191,N_2598,N_2838);
or UO_192 (O_192,N_2601,N_2979);
or UO_193 (O_193,N_2986,N_2589);
nand UO_194 (O_194,N_2943,N_2516);
or UO_195 (O_195,N_2405,N_2525);
nand UO_196 (O_196,N_2482,N_2834);
nand UO_197 (O_197,N_2604,N_2459);
xor UO_198 (O_198,N_2873,N_2789);
and UO_199 (O_199,N_2552,N_2585);
nand UO_200 (O_200,N_2945,N_2926);
nor UO_201 (O_201,N_2467,N_2486);
nor UO_202 (O_202,N_2909,N_2652);
nor UO_203 (O_203,N_2418,N_2477);
nand UO_204 (O_204,N_2887,N_2607);
nand UO_205 (O_205,N_2462,N_2417);
nand UO_206 (O_206,N_2720,N_2827);
and UO_207 (O_207,N_2967,N_2559);
nor UO_208 (O_208,N_2706,N_2428);
or UO_209 (O_209,N_2915,N_2832);
and UO_210 (O_210,N_2709,N_2863);
or UO_211 (O_211,N_2441,N_2849);
and UO_212 (O_212,N_2738,N_2970);
nand UO_213 (O_213,N_2669,N_2968);
or UO_214 (O_214,N_2452,N_2538);
nor UO_215 (O_215,N_2471,N_2614);
nor UO_216 (O_216,N_2540,N_2586);
nor UO_217 (O_217,N_2692,N_2658);
nand UO_218 (O_218,N_2560,N_2920);
and UO_219 (O_219,N_2689,N_2438);
or UO_220 (O_220,N_2476,N_2736);
nor UO_221 (O_221,N_2705,N_2413);
nand UO_222 (O_222,N_2740,N_2861);
and UO_223 (O_223,N_2528,N_2498);
nand UO_224 (O_224,N_2712,N_2854);
xor UO_225 (O_225,N_2557,N_2473);
or UO_226 (O_226,N_2420,N_2550);
and UO_227 (O_227,N_2581,N_2445);
or UO_228 (O_228,N_2870,N_2488);
nor UO_229 (O_229,N_2907,N_2866);
nand UO_230 (O_230,N_2805,N_2620);
and UO_231 (O_231,N_2621,N_2809);
nand UO_232 (O_232,N_2864,N_2576);
nor UO_233 (O_233,N_2436,N_2633);
nor UO_234 (O_234,N_2700,N_2913);
or UO_235 (O_235,N_2869,N_2422);
or UO_236 (O_236,N_2850,N_2619);
or UO_237 (O_237,N_2727,N_2602);
nor UO_238 (O_238,N_2695,N_2897);
nor UO_239 (O_239,N_2527,N_2637);
and UO_240 (O_240,N_2466,N_2430);
xnor UO_241 (O_241,N_2993,N_2609);
nand UO_242 (O_242,N_2714,N_2880);
or UO_243 (O_243,N_2681,N_2902);
nor UO_244 (O_244,N_2862,N_2622);
and UO_245 (O_245,N_2454,N_2953);
xor UO_246 (O_246,N_2900,N_2475);
and UO_247 (O_247,N_2812,N_2891);
and UO_248 (O_248,N_2939,N_2836);
and UO_249 (O_249,N_2646,N_2964);
nor UO_250 (O_250,N_2912,N_2825);
or UO_251 (O_251,N_2906,N_2444);
nor UO_252 (O_252,N_2522,N_2555);
and UO_253 (O_253,N_2924,N_2933);
nand UO_254 (O_254,N_2954,N_2801);
nand UO_255 (O_255,N_2506,N_2536);
nor UO_256 (O_256,N_2643,N_2844);
nand UO_257 (O_257,N_2487,N_2810);
and UO_258 (O_258,N_2782,N_2592);
nand UO_259 (O_259,N_2978,N_2867);
nand UO_260 (O_260,N_2828,N_2572);
nand UO_261 (O_261,N_2936,N_2448);
nand UO_262 (O_262,N_2937,N_2543);
nor UO_263 (O_263,N_2458,N_2823);
and UO_264 (O_264,N_2995,N_2981);
nor UO_265 (O_265,N_2582,N_2535);
nor UO_266 (O_266,N_2804,N_2764);
nor UO_267 (O_267,N_2916,N_2741);
or UO_268 (O_268,N_2889,N_2568);
nand UO_269 (O_269,N_2753,N_2783);
or UO_270 (O_270,N_2556,N_2983);
and UO_271 (O_271,N_2952,N_2496);
nand UO_272 (O_272,N_2703,N_2509);
nor UO_273 (O_273,N_2460,N_2721);
xnor UO_274 (O_274,N_2910,N_2877);
or UO_275 (O_275,N_2893,N_2521);
and UO_276 (O_276,N_2611,N_2921);
nor UO_277 (O_277,N_2434,N_2680);
and UO_278 (O_278,N_2479,N_2532);
nor UO_279 (O_279,N_2423,N_2848);
xor UO_280 (O_280,N_2626,N_2639);
or UO_281 (O_281,N_2429,N_2751);
and UO_282 (O_282,N_2539,N_2734);
nand UO_283 (O_283,N_2840,N_2987);
nor UO_284 (O_284,N_2575,N_2972);
nor UO_285 (O_285,N_2846,N_2548);
and UO_286 (O_286,N_2682,N_2468);
nor UO_287 (O_287,N_2663,N_2545);
nand UO_288 (O_288,N_2760,N_2593);
nor UO_289 (O_289,N_2743,N_2802);
nor UO_290 (O_290,N_2687,N_2484);
and UO_291 (O_291,N_2685,N_2502);
and UO_292 (O_292,N_2927,N_2570);
and UO_293 (O_293,N_2635,N_2503);
nand UO_294 (O_294,N_2400,N_2449);
xor UO_295 (O_295,N_2465,N_2904);
or UO_296 (O_296,N_2824,N_2574);
nor UO_297 (O_297,N_2774,N_2603);
nor UO_298 (O_298,N_2461,N_2763);
nand UO_299 (O_299,N_2725,N_2553);
nand UO_300 (O_300,N_2576,N_2936);
nor UO_301 (O_301,N_2870,N_2774);
or UO_302 (O_302,N_2880,N_2628);
and UO_303 (O_303,N_2528,N_2938);
nor UO_304 (O_304,N_2929,N_2566);
nor UO_305 (O_305,N_2857,N_2677);
nor UO_306 (O_306,N_2612,N_2594);
nand UO_307 (O_307,N_2634,N_2574);
nand UO_308 (O_308,N_2513,N_2696);
nand UO_309 (O_309,N_2552,N_2859);
and UO_310 (O_310,N_2930,N_2932);
nand UO_311 (O_311,N_2861,N_2400);
or UO_312 (O_312,N_2999,N_2960);
nor UO_313 (O_313,N_2801,N_2447);
nor UO_314 (O_314,N_2488,N_2577);
or UO_315 (O_315,N_2736,N_2945);
or UO_316 (O_316,N_2666,N_2648);
or UO_317 (O_317,N_2587,N_2549);
nand UO_318 (O_318,N_2854,N_2801);
nand UO_319 (O_319,N_2536,N_2419);
nand UO_320 (O_320,N_2842,N_2880);
and UO_321 (O_321,N_2919,N_2758);
xor UO_322 (O_322,N_2408,N_2463);
xnor UO_323 (O_323,N_2812,N_2844);
nor UO_324 (O_324,N_2746,N_2663);
or UO_325 (O_325,N_2465,N_2444);
nor UO_326 (O_326,N_2925,N_2943);
xnor UO_327 (O_327,N_2614,N_2730);
or UO_328 (O_328,N_2628,N_2947);
and UO_329 (O_329,N_2454,N_2586);
nand UO_330 (O_330,N_2503,N_2445);
xor UO_331 (O_331,N_2863,N_2557);
or UO_332 (O_332,N_2891,N_2568);
nand UO_333 (O_333,N_2615,N_2654);
and UO_334 (O_334,N_2594,N_2944);
nor UO_335 (O_335,N_2896,N_2893);
nand UO_336 (O_336,N_2557,N_2717);
nand UO_337 (O_337,N_2945,N_2413);
nor UO_338 (O_338,N_2555,N_2607);
nor UO_339 (O_339,N_2810,N_2499);
and UO_340 (O_340,N_2457,N_2641);
and UO_341 (O_341,N_2580,N_2495);
nand UO_342 (O_342,N_2495,N_2633);
nor UO_343 (O_343,N_2993,N_2815);
or UO_344 (O_344,N_2458,N_2501);
nand UO_345 (O_345,N_2899,N_2601);
or UO_346 (O_346,N_2756,N_2958);
nand UO_347 (O_347,N_2445,N_2401);
nor UO_348 (O_348,N_2419,N_2547);
and UO_349 (O_349,N_2862,N_2845);
or UO_350 (O_350,N_2906,N_2748);
or UO_351 (O_351,N_2492,N_2567);
and UO_352 (O_352,N_2400,N_2917);
nand UO_353 (O_353,N_2973,N_2906);
and UO_354 (O_354,N_2425,N_2685);
and UO_355 (O_355,N_2483,N_2689);
nor UO_356 (O_356,N_2964,N_2781);
nor UO_357 (O_357,N_2795,N_2712);
nand UO_358 (O_358,N_2761,N_2753);
or UO_359 (O_359,N_2588,N_2890);
xor UO_360 (O_360,N_2834,N_2672);
or UO_361 (O_361,N_2444,N_2466);
nand UO_362 (O_362,N_2524,N_2714);
or UO_363 (O_363,N_2648,N_2471);
nand UO_364 (O_364,N_2905,N_2983);
or UO_365 (O_365,N_2475,N_2516);
and UO_366 (O_366,N_2561,N_2746);
or UO_367 (O_367,N_2514,N_2881);
or UO_368 (O_368,N_2832,N_2890);
and UO_369 (O_369,N_2523,N_2480);
nor UO_370 (O_370,N_2644,N_2847);
or UO_371 (O_371,N_2791,N_2467);
nand UO_372 (O_372,N_2969,N_2421);
nand UO_373 (O_373,N_2430,N_2661);
and UO_374 (O_374,N_2429,N_2589);
nor UO_375 (O_375,N_2883,N_2766);
and UO_376 (O_376,N_2785,N_2403);
or UO_377 (O_377,N_2846,N_2989);
and UO_378 (O_378,N_2830,N_2806);
nor UO_379 (O_379,N_2556,N_2428);
xor UO_380 (O_380,N_2673,N_2573);
or UO_381 (O_381,N_2672,N_2547);
and UO_382 (O_382,N_2999,N_2919);
and UO_383 (O_383,N_2716,N_2633);
or UO_384 (O_384,N_2790,N_2768);
nand UO_385 (O_385,N_2557,N_2961);
nand UO_386 (O_386,N_2469,N_2466);
nand UO_387 (O_387,N_2761,N_2903);
nand UO_388 (O_388,N_2972,N_2557);
nor UO_389 (O_389,N_2858,N_2867);
or UO_390 (O_390,N_2979,N_2437);
or UO_391 (O_391,N_2755,N_2915);
nand UO_392 (O_392,N_2525,N_2816);
or UO_393 (O_393,N_2918,N_2489);
nand UO_394 (O_394,N_2731,N_2859);
or UO_395 (O_395,N_2469,N_2873);
nand UO_396 (O_396,N_2735,N_2839);
or UO_397 (O_397,N_2843,N_2453);
nor UO_398 (O_398,N_2734,N_2753);
nand UO_399 (O_399,N_2931,N_2621);
or UO_400 (O_400,N_2779,N_2709);
nand UO_401 (O_401,N_2487,N_2712);
and UO_402 (O_402,N_2572,N_2655);
and UO_403 (O_403,N_2439,N_2566);
nor UO_404 (O_404,N_2668,N_2624);
and UO_405 (O_405,N_2714,N_2571);
and UO_406 (O_406,N_2804,N_2808);
or UO_407 (O_407,N_2474,N_2492);
nand UO_408 (O_408,N_2804,N_2542);
nor UO_409 (O_409,N_2516,N_2886);
and UO_410 (O_410,N_2564,N_2946);
nand UO_411 (O_411,N_2704,N_2456);
nor UO_412 (O_412,N_2676,N_2928);
nor UO_413 (O_413,N_2747,N_2648);
nor UO_414 (O_414,N_2471,N_2792);
or UO_415 (O_415,N_2960,N_2571);
nand UO_416 (O_416,N_2543,N_2961);
or UO_417 (O_417,N_2602,N_2718);
nor UO_418 (O_418,N_2421,N_2846);
and UO_419 (O_419,N_2968,N_2915);
and UO_420 (O_420,N_2510,N_2987);
or UO_421 (O_421,N_2700,N_2706);
nand UO_422 (O_422,N_2527,N_2677);
or UO_423 (O_423,N_2744,N_2987);
and UO_424 (O_424,N_2721,N_2735);
or UO_425 (O_425,N_2750,N_2813);
nand UO_426 (O_426,N_2630,N_2696);
nand UO_427 (O_427,N_2506,N_2780);
and UO_428 (O_428,N_2888,N_2961);
or UO_429 (O_429,N_2773,N_2701);
or UO_430 (O_430,N_2519,N_2928);
or UO_431 (O_431,N_2412,N_2906);
or UO_432 (O_432,N_2623,N_2558);
nor UO_433 (O_433,N_2927,N_2558);
nor UO_434 (O_434,N_2498,N_2974);
and UO_435 (O_435,N_2912,N_2700);
and UO_436 (O_436,N_2933,N_2869);
nand UO_437 (O_437,N_2470,N_2816);
nand UO_438 (O_438,N_2765,N_2831);
or UO_439 (O_439,N_2651,N_2663);
or UO_440 (O_440,N_2472,N_2679);
or UO_441 (O_441,N_2754,N_2962);
nand UO_442 (O_442,N_2708,N_2826);
and UO_443 (O_443,N_2626,N_2545);
nor UO_444 (O_444,N_2445,N_2676);
nand UO_445 (O_445,N_2840,N_2950);
or UO_446 (O_446,N_2730,N_2533);
nor UO_447 (O_447,N_2857,N_2554);
nor UO_448 (O_448,N_2536,N_2963);
and UO_449 (O_449,N_2486,N_2427);
and UO_450 (O_450,N_2803,N_2730);
and UO_451 (O_451,N_2597,N_2546);
nor UO_452 (O_452,N_2551,N_2455);
nand UO_453 (O_453,N_2780,N_2421);
and UO_454 (O_454,N_2686,N_2497);
or UO_455 (O_455,N_2506,N_2503);
nand UO_456 (O_456,N_2841,N_2902);
or UO_457 (O_457,N_2715,N_2603);
or UO_458 (O_458,N_2924,N_2995);
nor UO_459 (O_459,N_2787,N_2461);
or UO_460 (O_460,N_2517,N_2644);
and UO_461 (O_461,N_2507,N_2762);
or UO_462 (O_462,N_2689,N_2448);
nand UO_463 (O_463,N_2427,N_2584);
nor UO_464 (O_464,N_2525,N_2615);
or UO_465 (O_465,N_2920,N_2772);
nand UO_466 (O_466,N_2733,N_2869);
and UO_467 (O_467,N_2920,N_2479);
and UO_468 (O_468,N_2792,N_2447);
and UO_469 (O_469,N_2598,N_2652);
and UO_470 (O_470,N_2917,N_2742);
and UO_471 (O_471,N_2923,N_2673);
xnor UO_472 (O_472,N_2541,N_2940);
nand UO_473 (O_473,N_2453,N_2448);
nor UO_474 (O_474,N_2987,N_2732);
xor UO_475 (O_475,N_2584,N_2732);
nand UO_476 (O_476,N_2783,N_2645);
and UO_477 (O_477,N_2699,N_2688);
or UO_478 (O_478,N_2446,N_2510);
nor UO_479 (O_479,N_2441,N_2819);
and UO_480 (O_480,N_2800,N_2420);
nand UO_481 (O_481,N_2655,N_2718);
and UO_482 (O_482,N_2470,N_2879);
nand UO_483 (O_483,N_2768,N_2749);
nand UO_484 (O_484,N_2406,N_2737);
or UO_485 (O_485,N_2893,N_2795);
or UO_486 (O_486,N_2904,N_2725);
nor UO_487 (O_487,N_2863,N_2414);
or UO_488 (O_488,N_2415,N_2713);
nor UO_489 (O_489,N_2491,N_2677);
or UO_490 (O_490,N_2748,N_2792);
nand UO_491 (O_491,N_2724,N_2615);
or UO_492 (O_492,N_2571,N_2580);
and UO_493 (O_493,N_2675,N_2913);
nand UO_494 (O_494,N_2401,N_2663);
and UO_495 (O_495,N_2867,N_2643);
and UO_496 (O_496,N_2560,N_2582);
nand UO_497 (O_497,N_2924,N_2940);
nand UO_498 (O_498,N_2570,N_2689);
and UO_499 (O_499,N_2997,N_2516);
endmodule