module basic_500_3000_500_60_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_66,In_205);
and U1 (N_1,In_375,In_429);
and U2 (N_2,In_399,In_37);
and U3 (N_3,In_463,In_123);
nor U4 (N_4,In_306,In_42);
or U5 (N_5,In_326,In_422);
xor U6 (N_6,In_359,In_269);
nand U7 (N_7,In_0,In_394);
or U8 (N_8,In_459,In_278);
or U9 (N_9,In_391,In_264);
or U10 (N_10,In_469,In_353);
or U11 (N_11,In_413,In_136);
and U12 (N_12,In_168,In_193);
nand U13 (N_13,In_18,In_20);
and U14 (N_14,In_164,In_292);
and U15 (N_15,In_54,In_84);
nor U16 (N_16,In_285,In_144);
nor U17 (N_17,In_129,In_266);
nor U18 (N_18,In_94,In_36);
and U19 (N_19,In_287,In_320);
or U20 (N_20,In_448,In_156);
or U21 (N_21,In_6,In_308);
nor U22 (N_22,In_152,In_442);
or U23 (N_23,In_171,In_361);
nor U24 (N_24,In_108,In_402);
nand U25 (N_25,In_208,In_484);
nor U26 (N_26,In_11,In_176);
and U27 (N_27,In_215,In_455);
nand U28 (N_28,In_179,In_410);
nor U29 (N_29,In_95,In_293);
and U30 (N_30,In_403,In_387);
xor U31 (N_31,In_104,In_126);
nand U32 (N_32,In_134,In_440);
nand U33 (N_33,In_240,In_158);
nand U34 (N_34,In_295,In_177);
or U35 (N_35,In_302,In_336);
and U36 (N_36,In_113,In_196);
nor U37 (N_37,In_55,In_393);
nand U38 (N_38,In_321,In_43);
xor U39 (N_39,In_253,In_451);
nor U40 (N_40,In_453,In_119);
and U41 (N_41,In_339,In_38);
xor U42 (N_42,In_207,In_351);
or U43 (N_43,In_76,In_186);
and U44 (N_44,In_227,In_187);
nor U45 (N_45,In_250,In_405);
nand U46 (N_46,In_314,In_226);
nand U47 (N_47,In_230,In_338);
nor U48 (N_48,In_460,In_198);
nor U49 (N_49,In_334,In_323);
or U50 (N_50,In_157,In_335);
nor U51 (N_51,In_404,In_221);
nor U52 (N_52,In_499,In_344);
nor U53 (N_53,In_409,In_172);
nor U54 (N_54,In_19,In_213);
and U55 (N_55,In_98,In_46);
nand U56 (N_56,In_89,In_224);
nand U57 (N_57,In_23,In_56);
nor U58 (N_58,In_189,In_452);
nand U59 (N_59,N_5,In_97);
or U60 (N_60,In_496,In_232);
and U61 (N_61,In_420,In_112);
nor U62 (N_62,In_234,In_162);
nand U63 (N_63,In_255,N_33);
nand U64 (N_64,In_72,In_426);
nand U65 (N_65,In_472,In_457);
xor U66 (N_66,In_454,In_125);
or U67 (N_67,In_280,In_461);
nor U68 (N_68,In_7,In_376);
or U69 (N_69,In_277,In_163);
and U70 (N_70,In_450,In_333);
and U71 (N_71,In_282,N_28);
and U72 (N_72,In_78,In_90);
or U73 (N_73,In_325,In_70);
and U74 (N_74,In_245,In_309);
nand U75 (N_75,In_236,In_33);
or U76 (N_76,In_329,In_83);
nand U77 (N_77,In_366,In_211);
and U78 (N_78,N_31,N_42);
nor U79 (N_79,In_133,In_290);
nor U80 (N_80,In_50,In_27);
nand U81 (N_81,In_148,In_32);
nand U82 (N_82,In_279,In_401);
nor U83 (N_83,In_485,In_217);
nand U84 (N_84,In_74,In_256);
xor U85 (N_85,In_433,In_203);
and U86 (N_86,In_53,In_464);
and U87 (N_87,In_99,In_223);
and U88 (N_88,N_17,In_380);
nand U89 (N_89,N_19,In_478);
and U90 (N_90,N_11,In_270);
xor U91 (N_91,In_300,In_117);
or U92 (N_92,In_182,In_267);
xor U93 (N_93,N_44,In_350);
and U94 (N_94,In_180,In_102);
nor U95 (N_95,In_465,In_346);
nor U96 (N_96,In_13,In_142);
or U97 (N_97,In_437,N_13);
and U98 (N_98,In_170,In_101);
or U99 (N_99,In_151,In_28);
nand U100 (N_100,In_297,In_384);
nor U101 (N_101,N_57,In_58);
nor U102 (N_102,In_327,In_424);
nand U103 (N_103,In_204,In_341);
or U104 (N_104,In_438,In_31);
or U105 (N_105,N_79,N_29);
or U106 (N_106,In_17,In_291);
nor U107 (N_107,In_425,In_35);
or U108 (N_108,In_367,In_114);
and U109 (N_109,In_388,In_109);
nor U110 (N_110,In_87,In_468);
nand U111 (N_111,In_75,In_483);
nand U112 (N_112,In_286,In_299);
xor U113 (N_113,In_482,N_75);
nand U114 (N_114,In_120,In_283);
nor U115 (N_115,In_276,In_337);
or U116 (N_116,In_247,In_145);
nand U117 (N_117,N_30,In_386);
nor U118 (N_118,In_110,In_486);
nor U119 (N_119,N_51,N_89);
nand U120 (N_120,In_385,In_408);
and U121 (N_121,In_428,In_246);
and U122 (N_122,In_155,In_103);
and U123 (N_123,In_490,In_79);
or U124 (N_124,In_59,In_441);
xor U125 (N_125,N_98,In_195);
or U126 (N_126,In_439,In_233);
xor U127 (N_127,N_7,In_175);
and U128 (N_128,In_248,In_435);
nor U129 (N_129,In_199,In_322);
nand U130 (N_130,In_141,In_495);
xnor U131 (N_131,In_197,In_487);
or U132 (N_132,In_492,In_273);
nand U133 (N_133,In_184,In_192);
nor U134 (N_134,In_105,In_34);
xnor U135 (N_135,N_53,In_445);
nor U136 (N_136,N_78,In_372);
or U137 (N_137,In_16,In_150);
or U138 (N_138,In_392,In_173);
or U139 (N_139,In_470,N_10);
xor U140 (N_140,N_69,In_190);
or U141 (N_141,In_271,N_91);
xor U142 (N_142,In_48,N_23);
and U143 (N_143,In_49,In_167);
and U144 (N_144,In_2,In_249);
and U145 (N_145,N_43,In_443);
nor U146 (N_146,In_132,N_52);
nor U147 (N_147,In_15,N_87);
nor U148 (N_148,In_310,In_191);
or U149 (N_149,In_476,In_462);
or U150 (N_150,In_206,N_131);
or U151 (N_151,In_364,In_477);
or U152 (N_152,N_50,N_58);
nor U153 (N_153,In_319,In_382);
nor U154 (N_154,In_317,N_38);
or U155 (N_155,N_70,In_434);
xnor U156 (N_156,N_1,In_218);
and U157 (N_157,In_288,In_122);
nand U158 (N_158,N_110,In_378);
nor U159 (N_159,In_82,N_101);
nand U160 (N_160,In_243,In_118);
nand U161 (N_161,In_354,N_72);
nor U162 (N_162,In_357,In_96);
xnor U163 (N_163,N_96,In_412);
nor U164 (N_164,N_104,In_165);
or U165 (N_165,In_258,N_60);
and U166 (N_166,In_12,In_106);
and U167 (N_167,N_105,N_26);
and U168 (N_168,In_396,In_491);
nor U169 (N_169,N_56,In_489);
and U170 (N_170,N_100,In_307);
xor U171 (N_171,In_449,In_235);
xnor U172 (N_172,In_369,N_88);
and U173 (N_173,In_398,N_68);
nand U174 (N_174,In_91,N_24);
or U175 (N_175,In_92,N_147);
nand U176 (N_176,N_4,N_71);
nor U177 (N_177,In_222,N_49);
and U178 (N_178,In_260,In_362);
or U179 (N_179,In_471,In_368);
nand U180 (N_180,In_415,N_3);
nand U181 (N_181,In_365,In_124);
nand U182 (N_182,N_63,In_254);
and U183 (N_183,In_360,In_411);
nor U184 (N_184,In_436,In_458);
xnor U185 (N_185,In_474,In_183);
and U186 (N_186,In_284,In_446);
nor U187 (N_187,In_14,N_118);
or U188 (N_188,N_21,In_47);
and U189 (N_189,N_113,In_261);
nand U190 (N_190,In_416,In_40);
nor U191 (N_191,In_301,N_35);
nand U192 (N_192,N_59,In_395);
nand U193 (N_193,N_106,In_24);
and U194 (N_194,N_102,In_447);
nor U195 (N_195,N_92,In_242);
nand U196 (N_196,In_257,In_44);
nand U197 (N_197,N_114,N_129);
xnor U198 (N_198,In_348,In_330);
nor U199 (N_199,In_111,N_64);
nor U200 (N_200,N_195,In_116);
nor U201 (N_201,In_340,In_418);
or U202 (N_202,In_377,N_36);
and U203 (N_203,In_275,N_194);
xor U204 (N_204,N_192,N_128);
nor U205 (N_205,In_373,In_400);
or U206 (N_206,N_45,N_90);
or U207 (N_207,N_95,N_139);
nor U208 (N_208,In_494,In_169);
and U209 (N_209,In_188,In_274);
nand U210 (N_210,In_417,N_148);
xor U211 (N_211,N_144,In_289);
xor U212 (N_212,N_116,N_73);
or U213 (N_213,N_61,N_46);
nand U214 (N_214,In_239,In_430);
nor U215 (N_215,N_8,In_374);
or U216 (N_216,N_186,N_12);
or U217 (N_217,N_163,N_166);
nor U218 (N_218,In_128,N_182);
xor U219 (N_219,N_165,In_332);
and U220 (N_220,In_147,N_161);
or U221 (N_221,N_108,In_8);
or U222 (N_222,In_154,N_193);
nor U223 (N_223,In_363,In_209);
or U224 (N_224,N_146,In_212);
xor U225 (N_225,In_1,N_76);
nor U226 (N_226,In_131,N_55);
xor U227 (N_227,In_480,N_112);
and U228 (N_228,N_14,N_85);
or U229 (N_229,N_18,N_48);
nor U230 (N_230,N_184,N_160);
and U231 (N_231,N_169,N_180);
nand U232 (N_232,In_30,N_149);
or U233 (N_233,In_29,In_39);
and U234 (N_234,In_107,N_142);
or U235 (N_235,N_74,In_80);
nor U236 (N_236,In_479,N_117);
xor U237 (N_237,N_156,In_159);
nor U238 (N_238,N_170,N_39);
or U239 (N_239,N_188,In_21);
and U240 (N_240,In_259,N_162);
nor U241 (N_241,N_121,In_347);
nand U242 (N_242,N_168,N_155);
xnor U243 (N_243,In_251,N_20);
nor U244 (N_244,In_139,In_160);
nand U245 (N_245,In_22,In_5);
or U246 (N_246,In_370,In_143);
nand U247 (N_247,N_93,N_62);
and U248 (N_248,In_26,In_265);
xnor U249 (N_249,N_120,In_130);
or U250 (N_250,N_213,N_22);
and U251 (N_251,N_15,N_223);
nor U252 (N_252,N_119,N_111);
nor U253 (N_253,In_3,N_54);
and U254 (N_254,N_80,In_65);
nor U255 (N_255,N_240,N_99);
nor U256 (N_256,N_199,In_303);
and U257 (N_257,In_315,N_154);
or U258 (N_258,N_222,N_229);
nand U259 (N_259,N_83,In_238);
and U260 (N_260,N_175,In_296);
or U261 (N_261,In_481,N_143);
or U262 (N_262,N_231,In_488);
nand U263 (N_263,N_221,In_140);
and U264 (N_264,In_414,N_32);
nor U265 (N_265,N_94,In_45);
nor U266 (N_266,In_345,N_137);
nor U267 (N_267,In_153,In_178);
nand U268 (N_268,N_205,N_174);
and U269 (N_269,In_444,In_64);
and U270 (N_270,In_383,N_77);
or U271 (N_271,In_61,In_200);
xnor U272 (N_272,N_236,In_355);
and U273 (N_273,In_466,N_132);
nand U274 (N_274,In_81,In_57);
nand U275 (N_275,In_63,In_298);
nor U276 (N_276,In_268,In_210);
and U277 (N_277,In_77,N_16);
xnor U278 (N_278,N_201,In_328);
nor U279 (N_279,In_214,N_216);
and U280 (N_280,In_10,N_217);
and U281 (N_281,In_294,In_86);
and U282 (N_282,N_173,N_41);
and U283 (N_283,In_252,In_51);
nor U284 (N_284,In_231,N_40);
nor U285 (N_285,N_189,N_239);
and U286 (N_286,In_166,In_318);
and U287 (N_287,In_311,N_67);
xnor U288 (N_288,N_158,In_407);
and U289 (N_289,N_133,In_85);
and U290 (N_290,N_210,N_81);
xnor U291 (N_291,N_181,In_194);
and U292 (N_292,In_9,In_381);
nor U293 (N_293,N_176,In_121);
xnor U294 (N_294,N_25,N_66);
or U295 (N_295,In_237,In_304);
or U296 (N_296,In_352,In_202);
nand U297 (N_297,N_97,N_204);
or U298 (N_298,N_157,In_493);
and U299 (N_299,N_230,N_238);
xor U300 (N_300,N_268,N_286);
or U301 (N_301,In_149,N_187);
and U302 (N_302,In_312,N_297);
nand U303 (N_303,N_256,N_284);
or U304 (N_304,N_296,N_244);
nor U305 (N_305,In_263,In_219);
nor U306 (N_306,N_277,In_356);
and U307 (N_307,N_84,In_421);
nand U308 (N_308,In_73,N_37);
or U309 (N_309,N_215,In_137);
nand U310 (N_310,In_220,N_135);
or U311 (N_311,N_293,In_93);
xnor U312 (N_312,N_269,N_126);
xnor U313 (N_313,N_218,N_233);
xnor U314 (N_314,N_212,In_427);
nand U315 (N_315,N_265,N_249);
and U316 (N_316,N_260,N_276);
nand U317 (N_317,In_431,N_130);
nand U318 (N_318,N_242,N_292);
nor U319 (N_319,In_379,In_371);
nand U320 (N_320,In_342,N_295);
and U321 (N_321,N_0,N_262);
and U322 (N_322,N_235,N_257);
nor U323 (N_323,In_397,N_275);
xnor U324 (N_324,N_298,N_299);
and U325 (N_325,N_124,In_467);
or U326 (N_326,N_232,N_272);
or U327 (N_327,N_266,In_241);
xnor U328 (N_328,N_123,N_274);
nor U329 (N_329,N_152,N_289);
or U330 (N_330,N_228,In_358);
nor U331 (N_331,N_243,N_6);
nor U332 (N_332,N_115,In_324);
nor U333 (N_333,N_171,In_88);
xor U334 (N_334,In_497,In_225);
and U335 (N_335,In_138,N_219);
nor U336 (N_336,N_47,N_267);
or U337 (N_337,N_291,In_343);
and U338 (N_338,N_185,In_406);
xnor U339 (N_339,In_181,N_177);
and U340 (N_340,N_34,N_141);
or U341 (N_341,N_248,In_69);
nand U342 (N_342,In_4,N_224);
and U343 (N_343,N_246,N_255);
xnor U344 (N_344,N_159,In_174);
nand U345 (N_345,N_178,In_389);
or U346 (N_346,In_229,N_27);
and U347 (N_347,In_115,N_264);
or U348 (N_348,N_2,N_287);
and U349 (N_349,In_216,In_68);
nor U350 (N_350,N_247,N_107);
nand U351 (N_351,In_62,N_337);
or U352 (N_352,N_339,N_172);
and U353 (N_353,N_340,In_331);
or U354 (N_354,N_167,N_317);
or U355 (N_355,N_203,In_432);
nand U356 (N_356,N_282,N_197);
nand U357 (N_357,In_305,N_103);
and U358 (N_358,In_244,N_211);
nor U359 (N_359,N_288,N_273);
nor U360 (N_360,N_323,N_328);
and U361 (N_361,In_185,In_272);
nand U362 (N_362,In_262,N_145);
nor U363 (N_363,N_302,In_475);
and U364 (N_364,N_138,N_279);
nand U365 (N_365,N_254,N_209);
xnor U366 (N_366,N_310,N_342);
nand U367 (N_367,N_311,N_136);
nand U368 (N_368,N_301,N_322);
nand U369 (N_369,N_306,N_191);
or U370 (N_370,In_201,N_324);
nand U371 (N_371,N_225,N_261);
nor U372 (N_372,N_253,N_140);
nand U373 (N_373,N_252,N_227);
and U374 (N_374,N_283,N_250);
or U375 (N_375,N_259,N_300);
nor U376 (N_376,N_305,N_206);
xor U377 (N_377,N_285,N_303);
nor U378 (N_378,In_456,N_346);
or U379 (N_379,In_419,In_423);
nor U380 (N_380,N_332,In_60);
and U381 (N_381,N_220,N_330);
nor U382 (N_382,N_341,N_226);
nor U383 (N_383,N_320,N_82);
and U384 (N_384,In_498,N_179);
nand U385 (N_385,In_161,N_200);
nand U386 (N_386,N_208,In_228);
and U387 (N_387,N_65,N_349);
nand U388 (N_388,N_307,N_316);
or U389 (N_389,N_334,N_151);
or U390 (N_390,N_348,N_214);
nor U391 (N_391,In_67,In_52);
nor U392 (N_392,N_321,N_280);
or U393 (N_393,N_294,N_331);
or U394 (N_394,N_318,N_304);
nand U395 (N_395,N_333,In_71);
xnor U396 (N_396,In_313,N_315);
and U397 (N_397,N_245,N_258);
nand U398 (N_398,N_314,N_325);
or U399 (N_399,N_345,N_134);
or U400 (N_400,N_384,N_198);
and U401 (N_401,N_313,In_146);
nor U402 (N_402,N_202,N_368);
nand U403 (N_403,N_364,N_355);
nand U404 (N_404,N_9,N_373);
or U405 (N_405,N_396,N_326);
and U406 (N_406,N_354,N_391);
nand U407 (N_407,N_122,N_366);
or U408 (N_408,N_164,N_390);
and U409 (N_409,N_352,N_329);
and U410 (N_410,N_371,N_234);
and U411 (N_411,N_369,N_290);
xnor U412 (N_412,N_393,N_361);
nand U413 (N_413,In_100,N_263);
and U414 (N_414,N_399,N_312);
and U415 (N_415,N_356,N_270);
nand U416 (N_416,N_353,In_25);
nor U417 (N_417,N_359,N_382);
or U418 (N_418,In_349,N_377);
nand U419 (N_419,In_127,N_336);
and U420 (N_420,N_380,N_381);
and U421 (N_421,In_473,N_357);
and U422 (N_422,N_308,N_347);
xnor U423 (N_423,N_362,N_338);
and U424 (N_424,N_370,N_372);
and U425 (N_425,N_153,N_365);
nor U426 (N_426,N_358,N_150);
nand U427 (N_427,N_351,N_395);
and U428 (N_428,N_196,N_374);
nand U429 (N_429,N_190,In_281);
or U430 (N_430,N_127,N_309);
nor U431 (N_431,N_344,N_271);
nor U432 (N_432,N_360,N_335);
nand U433 (N_433,N_367,In_316);
or U434 (N_434,N_376,In_390);
nand U435 (N_435,In_41,N_375);
nand U436 (N_436,N_241,N_379);
nand U437 (N_437,N_251,N_392);
or U438 (N_438,N_383,N_378);
or U439 (N_439,N_386,N_387);
nand U440 (N_440,N_86,N_350);
nand U441 (N_441,N_385,N_109);
nor U442 (N_442,N_237,N_278);
and U443 (N_443,N_207,N_343);
and U444 (N_444,N_327,N_183);
or U445 (N_445,N_281,N_388);
nor U446 (N_446,N_389,N_363);
or U447 (N_447,N_394,N_398);
nand U448 (N_448,N_319,N_397);
and U449 (N_449,In_135,N_125);
nor U450 (N_450,N_428,N_420);
and U451 (N_451,N_415,N_422);
nor U452 (N_452,N_409,N_430);
nand U453 (N_453,N_410,N_431);
or U454 (N_454,N_421,N_401);
and U455 (N_455,N_411,N_424);
nand U456 (N_456,N_447,N_402);
nor U457 (N_457,N_436,N_429);
nand U458 (N_458,N_407,N_433);
or U459 (N_459,N_416,N_426);
xnor U460 (N_460,N_423,N_425);
nand U461 (N_461,N_406,N_440);
nand U462 (N_462,N_443,N_417);
and U463 (N_463,N_439,N_446);
nor U464 (N_464,N_441,N_405);
nor U465 (N_465,N_413,N_419);
nor U466 (N_466,N_404,N_449);
or U467 (N_467,N_408,N_403);
and U468 (N_468,N_442,N_437);
or U469 (N_469,N_414,N_448);
nor U470 (N_470,N_432,N_427);
nand U471 (N_471,N_435,N_418);
or U472 (N_472,N_434,N_412);
nand U473 (N_473,N_445,N_400);
nand U474 (N_474,N_438,N_444);
and U475 (N_475,N_434,N_436);
nand U476 (N_476,N_445,N_401);
nor U477 (N_477,N_428,N_441);
nand U478 (N_478,N_412,N_413);
nand U479 (N_479,N_427,N_400);
nand U480 (N_480,N_405,N_436);
or U481 (N_481,N_441,N_446);
nand U482 (N_482,N_447,N_429);
nand U483 (N_483,N_418,N_407);
and U484 (N_484,N_431,N_432);
or U485 (N_485,N_421,N_400);
and U486 (N_486,N_426,N_408);
and U487 (N_487,N_411,N_408);
or U488 (N_488,N_415,N_437);
nor U489 (N_489,N_419,N_429);
nand U490 (N_490,N_430,N_424);
xor U491 (N_491,N_429,N_403);
nor U492 (N_492,N_408,N_414);
nand U493 (N_493,N_404,N_435);
nand U494 (N_494,N_433,N_427);
and U495 (N_495,N_441,N_421);
and U496 (N_496,N_445,N_405);
and U497 (N_497,N_444,N_431);
and U498 (N_498,N_436,N_426);
and U499 (N_499,N_424,N_443);
or U500 (N_500,N_490,N_498);
nor U501 (N_501,N_451,N_491);
or U502 (N_502,N_467,N_474);
and U503 (N_503,N_473,N_497);
or U504 (N_504,N_478,N_450);
or U505 (N_505,N_492,N_476);
or U506 (N_506,N_459,N_454);
nand U507 (N_507,N_460,N_494);
nand U508 (N_508,N_487,N_493);
nor U509 (N_509,N_489,N_499);
nor U510 (N_510,N_479,N_470);
nor U511 (N_511,N_486,N_466);
nand U512 (N_512,N_455,N_465);
and U513 (N_513,N_477,N_452);
or U514 (N_514,N_469,N_472);
or U515 (N_515,N_480,N_463);
nor U516 (N_516,N_485,N_462);
or U517 (N_517,N_496,N_495);
xor U518 (N_518,N_464,N_488);
or U519 (N_519,N_483,N_484);
nand U520 (N_520,N_468,N_475);
and U521 (N_521,N_461,N_471);
nor U522 (N_522,N_457,N_482);
or U523 (N_523,N_481,N_456);
and U524 (N_524,N_458,N_453);
nand U525 (N_525,N_480,N_484);
and U526 (N_526,N_450,N_477);
or U527 (N_527,N_455,N_484);
nand U528 (N_528,N_472,N_497);
nand U529 (N_529,N_464,N_456);
nand U530 (N_530,N_464,N_495);
nor U531 (N_531,N_485,N_488);
or U532 (N_532,N_489,N_481);
nand U533 (N_533,N_476,N_483);
and U534 (N_534,N_462,N_453);
nand U535 (N_535,N_468,N_451);
nand U536 (N_536,N_450,N_490);
or U537 (N_537,N_458,N_484);
nand U538 (N_538,N_464,N_498);
nor U539 (N_539,N_486,N_465);
xnor U540 (N_540,N_460,N_458);
nor U541 (N_541,N_478,N_452);
nor U542 (N_542,N_460,N_497);
and U543 (N_543,N_450,N_489);
or U544 (N_544,N_486,N_474);
nand U545 (N_545,N_482,N_460);
and U546 (N_546,N_474,N_471);
nand U547 (N_547,N_484,N_466);
nor U548 (N_548,N_487,N_465);
or U549 (N_549,N_473,N_465);
and U550 (N_550,N_520,N_503);
nand U551 (N_551,N_527,N_524);
or U552 (N_552,N_517,N_508);
nor U553 (N_553,N_521,N_548);
and U554 (N_554,N_515,N_540);
nand U555 (N_555,N_537,N_505);
nand U556 (N_556,N_528,N_516);
nand U557 (N_557,N_549,N_538);
nor U558 (N_558,N_543,N_512);
nand U559 (N_559,N_501,N_547);
nor U560 (N_560,N_518,N_514);
and U561 (N_561,N_541,N_506);
or U562 (N_562,N_534,N_523);
nor U563 (N_563,N_504,N_510);
or U564 (N_564,N_511,N_513);
or U565 (N_565,N_530,N_525);
and U566 (N_566,N_526,N_509);
and U567 (N_567,N_507,N_539);
and U568 (N_568,N_532,N_533);
or U569 (N_569,N_519,N_529);
or U570 (N_570,N_502,N_545);
xnor U571 (N_571,N_536,N_500);
and U572 (N_572,N_544,N_522);
and U573 (N_573,N_542,N_531);
xor U574 (N_574,N_535,N_546);
nor U575 (N_575,N_525,N_529);
and U576 (N_576,N_510,N_515);
nand U577 (N_577,N_533,N_510);
nand U578 (N_578,N_542,N_504);
or U579 (N_579,N_516,N_522);
or U580 (N_580,N_530,N_506);
and U581 (N_581,N_528,N_529);
nand U582 (N_582,N_547,N_503);
or U583 (N_583,N_526,N_525);
or U584 (N_584,N_511,N_523);
nor U585 (N_585,N_532,N_544);
and U586 (N_586,N_531,N_516);
nand U587 (N_587,N_538,N_537);
xor U588 (N_588,N_513,N_503);
nor U589 (N_589,N_512,N_514);
nor U590 (N_590,N_526,N_501);
nor U591 (N_591,N_500,N_541);
or U592 (N_592,N_510,N_532);
xor U593 (N_593,N_543,N_508);
and U594 (N_594,N_516,N_512);
and U595 (N_595,N_546,N_539);
xnor U596 (N_596,N_542,N_526);
nand U597 (N_597,N_532,N_514);
xor U598 (N_598,N_501,N_511);
and U599 (N_599,N_540,N_521);
and U600 (N_600,N_592,N_586);
nand U601 (N_601,N_594,N_588);
nor U602 (N_602,N_591,N_578);
and U603 (N_603,N_573,N_576);
nand U604 (N_604,N_585,N_562);
nor U605 (N_605,N_550,N_560);
nor U606 (N_606,N_564,N_561);
nand U607 (N_607,N_599,N_587);
and U608 (N_608,N_566,N_574);
nand U609 (N_609,N_577,N_552);
or U610 (N_610,N_595,N_571);
xor U611 (N_611,N_554,N_581);
xor U612 (N_612,N_569,N_579);
nor U613 (N_613,N_575,N_583);
xnor U614 (N_614,N_559,N_568);
and U615 (N_615,N_598,N_582);
or U616 (N_616,N_589,N_551);
or U617 (N_617,N_565,N_597);
nor U618 (N_618,N_584,N_590);
nand U619 (N_619,N_553,N_563);
nor U620 (N_620,N_556,N_593);
nand U621 (N_621,N_580,N_567);
nand U622 (N_622,N_557,N_558);
nor U623 (N_623,N_555,N_596);
nor U624 (N_624,N_570,N_572);
nor U625 (N_625,N_596,N_552);
nand U626 (N_626,N_567,N_577);
nor U627 (N_627,N_553,N_565);
nor U628 (N_628,N_576,N_557);
nor U629 (N_629,N_568,N_591);
or U630 (N_630,N_565,N_557);
and U631 (N_631,N_593,N_594);
nand U632 (N_632,N_599,N_597);
nor U633 (N_633,N_551,N_587);
nand U634 (N_634,N_564,N_579);
nor U635 (N_635,N_595,N_577);
xor U636 (N_636,N_596,N_581);
nand U637 (N_637,N_562,N_567);
nand U638 (N_638,N_597,N_556);
and U639 (N_639,N_581,N_563);
nor U640 (N_640,N_559,N_583);
nand U641 (N_641,N_591,N_562);
nor U642 (N_642,N_589,N_565);
nor U643 (N_643,N_586,N_553);
nor U644 (N_644,N_579,N_580);
nand U645 (N_645,N_584,N_580);
nor U646 (N_646,N_557,N_562);
nand U647 (N_647,N_550,N_573);
and U648 (N_648,N_590,N_553);
nor U649 (N_649,N_597,N_569);
nand U650 (N_650,N_607,N_624);
nor U651 (N_651,N_615,N_619);
nor U652 (N_652,N_642,N_649);
nand U653 (N_653,N_614,N_626);
nand U654 (N_654,N_617,N_613);
and U655 (N_655,N_629,N_608);
and U656 (N_656,N_644,N_621);
nand U657 (N_657,N_605,N_637);
and U658 (N_658,N_609,N_640);
and U659 (N_659,N_632,N_628);
xor U660 (N_660,N_643,N_645);
nand U661 (N_661,N_603,N_639);
and U662 (N_662,N_646,N_631);
and U663 (N_663,N_630,N_604);
nand U664 (N_664,N_610,N_622);
and U665 (N_665,N_612,N_623);
and U666 (N_666,N_611,N_616);
nand U667 (N_667,N_601,N_633);
nand U668 (N_668,N_636,N_627);
or U669 (N_669,N_625,N_647);
and U670 (N_670,N_648,N_620);
nor U671 (N_671,N_638,N_618);
nor U672 (N_672,N_600,N_602);
nand U673 (N_673,N_641,N_635);
nand U674 (N_674,N_634,N_606);
or U675 (N_675,N_644,N_615);
xor U676 (N_676,N_631,N_633);
or U677 (N_677,N_611,N_636);
and U678 (N_678,N_633,N_639);
xor U679 (N_679,N_646,N_636);
nor U680 (N_680,N_618,N_604);
or U681 (N_681,N_601,N_605);
nor U682 (N_682,N_623,N_610);
xnor U683 (N_683,N_649,N_614);
xor U684 (N_684,N_639,N_605);
nand U685 (N_685,N_611,N_631);
nor U686 (N_686,N_628,N_601);
and U687 (N_687,N_602,N_633);
nor U688 (N_688,N_636,N_600);
nor U689 (N_689,N_634,N_642);
nand U690 (N_690,N_623,N_622);
nand U691 (N_691,N_607,N_612);
and U692 (N_692,N_645,N_642);
nand U693 (N_693,N_617,N_640);
xor U694 (N_694,N_637,N_638);
xor U695 (N_695,N_648,N_636);
nand U696 (N_696,N_615,N_635);
and U697 (N_697,N_640,N_607);
or U698 (N_698,N_603,N_631);
nand U699 (N_699,N_636,N_623);
xnor U700 (N_700,N_663,N_692);
nor U701 (N_701,N_676,N_695);
and U702 (N_702,N_654,N_688);
xnor U703 (N_703,N_694,N_671);
nand U704 (N_704,N_689,N_667);
nand U705 (N_705,N_666,N_650);
xor U706 (N_706,N_673,N_655);
nand U707 (N_707,N_686,N_658);
nand U708 (N_708,N_698,N_685);
and U709 (N_709,N_664,N_669);
nand U710 (N_710,N_677,N_687);
and U711 (N_711,N_660,N_681);
nand U712 (N_712,N_670,N_651);
nand U713 (N_713,N_674,N_690);
nor U714 (N_714,N_668,N_656);
and U715 (N_715,N_672,N_679);
or U716 (N_716,N_696,N_653);
and U717 (N_717,N_678,N_680);
nor U718 (N_718,N_699,N_684);
nor U719 (N_719,N_682,N_675);
and U720 (N_720,N_661,N_691);
and U721 (N_721,N_657,N_665);
nand U722 (N_722,N_697,N_652);
and U723 (N_723,N_659,N_683);
and U724 (N_724,N_693,N_662);
nor U725 (N_725,N_689,N_696);
nand U726 (N_726,N_673,N_653);
nand U727 (N_727,N_684,N_688);
xor U728 (N_728,N_653,N_670);
and U729 (N_729,N_677,N_668);
nor U730 (N_730,N_655,N_685);
nor U731 (N_731,N_662,N_687);
or U732 (N_732,N_673,N_683);
or U733 (N_733,N_699,N_673);
or U734 (N_734,N_689,N_684);
nand U735 (N_735,N_650,N_694);
nand U736 (N_736,N_666,N_679);
nor U737 (N_737,N_655,N_690);
or U738 (N_738,N_651,N_675);
nand U739 (N_739,N_681,N_668);
nor U740 (N_740,N_650,N_670);
or U741 (N_741,N_673,N_688);
or U742 (N_742,N_680,N_689);
or U743 (N_743,N_689,N_686);
nor U744 (N_744,N_655,N_693);
nand U745 (N_745,N_654,N_660);
or U746 (N_746,N_688,N_655);
nand U747 (N_747,N_656,N_681);
or U748 (N_748,N_674,N_672);
and U749 (N_749,N_650,N_699);
and U750 (N_750,N_706,N_705);
nand U751 (N_751,N_737,N_728);
nand U752 (N_752,N_741,N_723);
and U753 (N_753,N_715,N_712);
and U754 (N_754,N_725,N_707);
xor U755 (N_755,N_721,N_745);
nor U756 (N_756,N_719,N_704);
xor U757 (N_757,N_731,N_717);
nor U758 (N_758,N_746,N_714);
nor U759 (N_759,N_711,N_722);
and U760 (N_760,N_739,N_749);
and U761 (N_761,N_702,N_727);
nand U762 (N_762,N_732,N_740);
or U763 (N_763,N_733,N_735);
nand U764 (N_764,N_724,N_744);
or U765 (N_765,N_718,N_716);
or U766 (N_766,N_700,N_720);
and U767 (N_767,N_736,N_703);
nor U768 (N_768,N_710,N_730);
xnor U769 (N_769,N_709,N_743);
nor U770 (N_770,N_713,N_748);
or U771 (N_771,N_729,N_742);
nor U772 (N_772,N_708,N_734);
xnor U773 (N_773,N_738,N_726);
xor U774 (N_774,N_747,N_701);
xnor U775 (N_775,N_705,N_708);
or U776 (N_776,N_708,N_700);
nor U777 (N_777,N_716,N_733);
xor U778 (N_778,N_739,N_717);
and U779 (N_779,N_721,N_746);
and U780 (N_780,N_709,N_704);
nand U781 (N_781,N_704,N_707);
nand U782 (N_782,N_717,N_706);
nor U783 (N_783,N_725,N_727);
nand U784 (N_784,N_731,N_712);
nor U785 (N_785,N_724,N_712);
xnor U786 (N_786,N_733,N_747);
and U787 (N_787,N_727,N_749);
nand U788 (N_788,N_734,N_726);
and U789 (N_789,N_723,N_734);
nor U790 (N_790,N_723,N_737);
or U791 (N_791,N_743,N_700);
nand U792 (N_792,N_735,N_726);
xor U793 (N_793,N_730,N_701);
and U794 (N_794,N_719,N_744);
or U795 (N_795,N_743,N_730);
and U796 (N_796,N_735,N_721);
nand U797 (N_797,N_709,N_713);
xnor U798 (N_798,N_731,N_744);
or U799 (N_799,N_703,N_731);
and U800 (N_800,N_777,N_767);
nand U801 (N_801,N_794,N_757);
xor U802 (N_802,N_766,N_774);
and U803 (N_803,N_750,N_763);
xnor U804 (N_804,N_770,N_792);
or U805 (N_805,N_754,N_759);
and U806 (N_806,N_797,N_799);
nor U807 (N_807,N_793,N_764);
nand U808 (N_808,N_756,N_758);
and U809 (N_809,N_755,N_761);
nor U810 (N_810,N_778,N_785);
nor U811 (N_811,N_786,N_791);
nand U812 (N_812,N_772,N_788);
and U813 (N_813,N_779,N_765);
nor U814 (N_814,N_783,N_768);
nor U815 (N_815,N_760,N_780);
or U816 (N_816,N_795,N_769);
nor U817 (N_817,N_781,N_782);
nand U818 (N_818,N_784,N_787);
or U819 (N_819,N_762,N_775);
nand U820 (N_820,N_751,N_776);
or U821 (N_821,N_752,N_753);
or U822 (N_822,N_798,N_789);
nand U823 (N_823,N_796,N_771);
nor U824 (N_824,N_773,N_790);
or U825 (N_825,N_754,N_776);
nand U826 (N_826,N_791,N_768);
xnor U827 (N_827,N_795,N_762);
and U828 (N_828,N_758,N_773);
and U829 (N_829,N_754,N_792);
and U830 (N_830,N_787,N_766);
and U831 (N_831,N_773,N_754);
nor U832 (N_832,N_794,N_777);
nand U833 (N_833,N_799,N_796);
or U834 (N_834,N_789,N_776);
nand U835 (N_835,N_784,N_765);
xor U836 (N_836,N_766,N_789);
or U837 (N_837,N_775,N_756);
nor U838 (N_838,N_760,N_789);
or U839 (N_839,N_778,N_780);
nand U840 (N_840,N_778,N_767);
nor U841 (N_841,N_795,N_753);
and U842 (N_842,N_789,N_777);
or U843 (N_843,N_776,N_791);
nand U844 (N_844,N_796,N_761);
or U845 (N_845,N_794,N_755);
nand U846 (N_846,N_794,N_789);
xnor U847 (N_847,N_757,N_751);
and U848 (N_848,N_762,N_793);
xor U849 (N_849,N_788,N_754);
nor U850 (N_850,N_848,N_806);
or U851 (N_851,N_805,N_821);
nand U852 (N_852,N_849,N_816);
and U853 (N_853,N_809,N_801);
nor U854 (N_854,N_813,N_815);
or U855 (N_855,N_826,N_825);
or U856 (N_856,N_807,N_808);
nor U857 (N_857,N_804,N_847);
or U858 (N_858,N_828,N_800);
nand U859 (N_859,N_811,N_842);
nor U860 (N_860,N_840,N_833);
nor U861 (N_861,N_803,N_817);
and U862 (N_862,N_838,N_812);
nand U863 (N_863,N_814,N_823);
nor U864 (N_864,N_818,N_829);
nand U865 (N_865,N_834,N_827);
nor U866 (N_866,N_832,N_810);
nor U867 (N_867,N_835,N_836);
xor U868 (N_868,N_830,N_839);
or U869 (N_869,N_819,N_844);
nor U870 (N_870,N_822,N_846);
and U871 (N_871,N_837,N_802);
or U872 (N_872,N_824,N_845);
nand U873 (N_873,N_820,N_843);
and U874 (N_874,N_831,N_841);
or U875 (N_875,N_843,N_846);
nor U876 (N_876,N_819,N_825);
or U877 (N_877,N_807,N_800);
xor U878 (N_878,N_809,N_802);
nor U879 (N_879,N_825,N_832);
nor U880 (N_880,N_838,N_806);
xor U881 (N_881,N_809,N_818);
or U882 (N_882,N_814,N_849);
and U883 (N_883,N_834,N_820);
nor U884 (N_884,N_823,N_839);
or U885 (N_885,N_812,N_828);
or U886 (N_886,N_809,N_830);
nand U887 (N_887,N_841,N_810);
and U888 (N_888,N_840,N_821);
or U889 (N_889,N_832,N_838);
or U890 (N_890,N_849,N_811);
nor U891 (N_891,N_808,N_834);
nor U892 (N_892,N_829,N_806);
and U893 (N_893,N_820,N_805);
or U894 (N_894,N_800,N_848);
or U895 (N_895,N_819,N_812);
or U896 (N_896,N_834,N_846);
nand U897 (N_897,N_847,N_809);
nor U898 (N_898,N_840,N_828);
nand U899 (N_899,N_826,N_819);
and U900 (N_900,N_867,N_897);
or U901 (N_901,N_862,N_859);
nor U902 (N_902,N_880,N_852);
nor U903 (N_903,N_873,N_875);
nand U904 (N_904,N_855,N_883);
and U905 (N_905,N_868,N_896);
nand U906 (N_906,N_885,N_853);
or U907 (N_907,N_895,N_856);
and U908 (N_908,N_886,N_863);
or U909 (N_909,N_891,N_884);
nor U910 (N_910,N_864,N_858);
or U911 (N_911,N_877,N_851);
or U912 (N_912,N_865,N_866);
and U913 (N_913,N_894,N_861);
and U914 (N_914,N_892,N_898);
nor U915 (N_915,N_893,N_899);
and U916 (N_916,N_879,N_860);
and U917 (N_917,N_874,N_882);
nor U918 (N_918,N_889,N_871);
nand U919 (N_919,N_872,N_857);
nor U920 (N_920,N_878,N_881);
and U921 (N_921,N_870,N_854);
nand U922 (N_922,N_876,N_869);
or U923 (N_923,N_888,N_890);
nand U924 (N_924,N_850,N_887);
and U925 (N_925,N_877,N_882);
and U926 (N_926,N_898,N_853);
nor U927 (N_927,N_896,N_875);
or U928 (N_928,N_883,N_893);
nor U929 (N_929,N_870,N_859);
and U930 (N_930,N_882,N_872);
or U931 (N_931,N_896,N_895);
nor U932 (N_932,N_884,N_887);
and U933 (N_933,N_884,N_867);
nor U934 (N_934,N_850,N_867);
or U935 (N_935,N_875,N_871);
or U936 (N_936,N_855,N_880);
and U937 (N_937,N_858,N_868);
xor U938 (N_938,N_898,N_854);
nor U939 (N_939,N_855,N_876);
nor U940 (N_940,N_868,N_899);
and U941 (N_941,N_861,N_895);
or U942 (N_942,N_872,N_866);
nor U943 (N_943,N_889,N_865);
nor U944 (N_944,N_864,N_888);
or U945 (N_945,N_851,N_880);
or U946 (N_946,N_880,N_872);
nor U947 (N_947,N_869,N_858);
nand U948 (N_948,N_861,N_859);
and U949 (N_949,N_895,N_869);
nor U950 (N_950,N_937,N_914);
or U951 (N_951,N_925,N_934);
or U952 (N_952,N_921,N_930);
nand U953 (N_953,N_944,N_917);
or U954 (N_954,N_948,N_920);
nor U955 (N_955,N_928,N_904);
nor U956 (N_956,N_940,N_946);
or U957 (N_957,N_902,N_912);
nor U958 (N_958,N_933,N_939);
or U959 (N_959,N_935,N_922);
xnor U960 (N_960,N_938,N_910);
xor U961 (N_961,N_941,N_909);
and U962 (N_962,N_936,N_932);
nor U963 (N_963,N_919,N_916);
nor U964 (N_964,N_949,N_913);
nor U965 (N_965,N_911,N_947);
and U966 (N_966,N_943,N_915);
nor U967 (N_967,N_907,N_926);
and U968 (N_968,N_901,N_931);
nand U969 (N_969,N_900,N_927);
and U970 (N_970,N_905,N_923);
or U971 (N_971,N_924,N_942);
and U972 (N_972,N_906,N_908);
xor U973 (N_973,N_903,N_918);
and U974 (N_974,N_929,N_945);
or U975 (N_975,N_907,N_947);
and U976 (N_976,N_948,N_918);
nand U977 (N_977,N_942,N_927);
nor U978 (N_978,N_901,N_904);
nor U979 (N_979,N_929,N_948);
nor U980 (N_980,N_922,N_908);
xnor U981 (N_981,N_908,N_944);
and U982 (N_982,N_938,N_906);
nand U983 (N_983,N_937,N_923);
xnor U984 (N_984,N_937,N_944);
nand U985 (N_985,N_929,N_923);
nor U986 (N_986,N_930,N_922);
or U987 (N_987,N_921,N_946);
nand U988 (N_988,N_920,N_942);
or U989 (N_989,N_907,N_906);
nand U990 (N_990,N_911,N_945);
nor U991 (N_991,N_902,N_905);
or U992 (N_992,N_913,N_900);
xnor U993 (N_993,N_943,N_924);
nand U994 (N_994,N_912,N_922);
nand U995 (N_995,N_948,N_904);
xor U996 (N_996,N_908,N_948);
nor U997 (N_997,N_940,N_912);
or U998 (N_998,N_936,N_916);
or U999 (N_999,N_909,N_932);
and U1000 (N_1000,N_971,N_970);
or U1001 (N_1001,N_962,N_976);
nor U1002 (N_1002,N_969,N_993);
and U1003 (N_1003,N_963,N_958);
nor U1004 (N_1004,N_974,N_973);
nand U1005 (N_1005,N_966,N_984);
nor U1006 (N_1006,N_982,N_953);
nor U1007 (N_1007,N_952,N_990);
xnor U1008 (N_1008,N_989,N_988);
xor U1009 (N_1009,N_998,N_995);
nor U1010 (N_1010,N_950,N_959);
nor U1011 (N_1011,N_961,N_972);
xor U1012 (N_1012,N_999,N_978);
nand U1013 (N_1013,N_975,N_956);
and U1014 (N_1014,N_980,N_965);
nor U1015 (N_1015,N_985,N_957);
and U1016 (N_1016,N_977,N_994);
and U1017 (N_1017,N_992,N_964);
nor U1018 (N_1018,N_951,N_987);
nand U1019 (N_1019,N_997,N_979);
nand U1020 (N_1020,N_986,N_983);
xor U1021 (N_1021,N_954,N_991);
or U1022 (N_1022,N_981,N_968);
nand U1023 (N_1023,N_960,N_996);
and U1024 (N_1024,N_955,N_967);
nor U1025 (N_1025,N_999,N_975);
nor U1026 (N_1026,N_988,N_992);
or U1027 (N_1027,N_952,N_998);
nand U1028 (N_1028,N_999,N_991);
nand U1029 (N_1029,N_950,N_979);
nor U1030 (N_1030,N_989,N_976);
nand U1031 (N_1031,N_966,N_990);
and U1032 (N_1032,N_958,N_971);
or U1033 (N_1033,N_986,N_966);
or U1034 (N_1034,N_976,N_997);
or U1035 (N_1035,N_975,N_955);
nand U1036 (N_1036,N_989,N_957);
nand U1037 (N_1037,N_964,N_976);
or U1038 (N_1038,N_986,N_954);
nand U1039 (N_1039,N_978,N_979);
and U1040 (N_1040,N_992,N_977);
and U1041 (N_1041,N_984,N_986);
nor U1042 (N_1042,N_989,N_998);
and U1043 (N_1043,N_998,N_993);
or U1044 (N_1044,N_970,N_976);
and U1045 (N_1045,N_988,N_974);
and U1046 (N_1046,N_962,N_995);
nand U1047 (N_1047,N_954,N_995);
nand U1048 (N_1048,N_965,N_979);
nand U1049 (N_1049,N_973,N_976);
nor U1050 (N_1050,N_1004,N_1040);
xor U1051 (N_1051,N_1045,N_1003);
nand U1052 (N_1052,N_1032,N_1024);
nand U1053 (N_1053,N_1039,N_1001);
nand U1054 (N_1054,N_1027,N_1006);
or U1055 (N_1055,N_1025,N_1046);
nor U1056 (N_1056,N_1012,N_1020);
xnor U1057 (N_1057,N_1037,N_1023);
nand U1058 (N_1058,N_1034,N_1047);
nor U1059 (N_1059,N_1017,N_1030);
nor U1060 (N_1060,N_1033,N_1013);
or U1061 (N_1061,N_1038,N_1019);
nand U1062 (N_1062,N_1011,N_1041);
nor U1063 (N_1063,N_1009,N_1021);
or U1064 (N_1064,N_1016,N_1028);
and U1065 (N_1065,N_1007,N_1022);
and U1066 (N_1066,N_1049,N_1014);
nand U1067 (N_1067,N_1029,N_1031);
nand U1068 (N_1068,N_1008,N_1035);
nand U1069 (N_1069,N_1018,N_1010);
nor U1070 (N_1070,N_1043,N_1044);
and U1071 (N_1071,N_1015,N_1000);
nand U1072 (N_1072,N_1005,N_1002);
and U1073 (N_1073,N_1048,N_1036);
nand U1074 (N_1074,N_1042,N_1026);
nor U1075 (N_1075,N_1035,N_1010);
and U1076 (N_1076,N_1038,N_1045);
nand U1077 (N_1077,N_1028,N_1000);
nor U1078 (N_1078,N_1030,N_1001);
or U1079 (N_1079,N_1013,N_1049);
nand U1080 (N_1080,N_1008,N_1027);
nand U1081 (N_1081,N_1024,N_1025);
or U1082 (N_1082,N_1015,N_1012);
or U1083 (N_1083,N_1010,N_1031);
and U1084 (N_1084,N_1011,N_1046);
and U1085 (N_1085,N_1047,N_1030);
nand U1086 (N_1086,N_1047,N_1009);
nor U1087 (N_1087,N_1027,N_1034);
xnor U1088 (N_1088,N_1003,N_1034);
or U1089 (N_1089,N_1018,N_1049);
nand U1090 (N_1090,N_1043,N_1021);
nand U1091 (N_1091,N_1035,N_1045);
nor U1092 (N_1092,N_1014,N_1038);
or U1093 (N_1093,N_1045,N_1008);
nor U1094 (N_1094,N_1005,N_1007);
xnor U1095 (N_1095,N_1048,N_1035);
or U1096 (N_1096,N_1017,N_1022);
or U1097 (N_1097,N_1023,N_1028);
xor U1098 (N_1098,N_1010,N_1041);
xor U1099 (N_1099,N_1018,N_1006);
nor U1100 (N_1100,N_1079,N_1070);
xnor U1101 (N_1101,N_1089,N_1094);
or U1102 (N_1102,N_1097,N_1087);
and U1103 (N_1103,N_1091,N_1095);
and U1104 (N_1104,N_1061,N_1057);
and U1105 (N_1105,N_1053,N_1072);
nand U1106 (N_1106,N_1075,N_1096);
xor U1107 (N_1107,N_1051,N_1063);
or U1108 (N_1108,N_1050,N_1078);
and U1109 (N_1109,N_1082,N_1066);
nand U1110 (N_1110,N_1058,N_1062);
and U1111 (N_1111,N_1081,N_1088);
nand U1112 (N_1112,N_1060,N_1067);
nor U1113 (N_1113,N_1052,N_1085);
nor U1114 (N_1114,N_1077,N_1090);
and U1115 (N_1115,N_1098,N_1065);
nor U1116 (N_1116,N_1099,N_1055);
nor U1117 (N_1117,N_1092,N_1093);
nor U1118 (N_1118,N_1076,N_1073);
and U1119 (N_1119,N_1068,N_1056);
nor U1120 (N_1120,N_1064,N_1086);
or U1121 (N_1121,N_1071,N_1084);
nor U1122 (N_1122,N_1054,N_1083);
and U1123 (N_1123,N_1059,N_1080);
or U1124 (N_1124,N_1074,N_1069);
and U1125 (N_1125,N_1093,N_1069);
or U1126 (N_1126,N_1052,N_1092);
and U1127 (N_1127,N_1052,N_1089);
nor U1128 (N_1128,N_1080,N_1090);
nor U1129 (N_1129,N_1094,N_1097);
or U1130 (N_1130,N_1068,N_1083);
nor U1131 (N_1131,N_1080,N_1063);
xor U1132 (N_1132,N_1093,N_1073);
and U1133 (N_1133,N_1062,N_1092);
and U1134 (N_1134,N_1073,N_1077);
or U1135 (N_1135,N_1079,N_1098);
and U1136 (N_1136,N_1076,N_1063);
nor U1137 (N_1137,N_1080,N_1058);
nand U1138 (N_1138,N_1051,N_1054);
or U1139 (N_1139,N_1050,N_1099);
or U1140 (N_1140,N_1062,N_1059);
and U1141 (N_1141,N_1061,N_1085);
and U1142 (N_1142,N_1078,N_1093);
and U1143 (N_1143,N_1086,N_1085);
nand U1144 (N_1144,N_1074,N_1071);
xnor U1145 (N_1145,N_1086,N_1066);
or U1146 (N_1146,N_1082,N_1088);
nor U1147 (N_1147,N_1089,N_1096);
nor U1148 (N_1148,N_1091,N_1081);
or U1149 (N_1149,N_1074,N_1084);
nor U1150 (N_1150,N_1124,N_1141);
and U1151 (N_1151,N_1111,N_1103);
and U1152 (N_1152,N_1112,N_1121);
nor U1153 (N_1153,N_1122,N_1127);
and U1154 (N_1154,N_1139,N_1123);
or U1155 (N_1155,N_1108,N_1142);
xor U1156 (N_1156,N_1101,N_1106);
nand U1157 (N_1157,N_1119,N_1125);
nor U1158 (N_1158,N_1131,N_1128);
or U1159 (N_1159,N_1104,N_1115);
or U1160 (N_1160,N_1135,N_1120);
and U1161 (N_1161,N_1130,N_1118);
or U1162 (N_1162,N_1117,N_1100);
and U1163 (N_1163,N_1140,N_1116);
nand U1164 (N_1164,N_1143,N_1129);
and U1165 (N_1165,N_1147,N_1145);
nor U1166 (N_1166,N_1107,N_1126);
or U1167 (N_1167,N_1110,N_1109);
or U1168 (N_1168,N_1146,N_1148);
xnor U1169 (N_1169,N_1149,N_1102);
xnor U1170 (N_1170,N_1144,N_1132);
nand U1171 (N_1171,N_1114,N_1136);
or U1172 (N_1172,N_1137,N_1138);
or U1173 (N_1173,N_1134,N_1105);
nand U1174 (N_1174,N_1133,N_1113);
and U1175 (N_1175,N_1144,N_1122);
or U1176 (N_1176,N_1133,N_1119);
or U1177 (N_1177,N_1132,N_1112);
nand U1178 (N_1178,N_1140,N_1129);
or U1179 (N_1179,N_1105,N_1114);
and U1180 (N_1180,N_1141,N_1142);
or U1181 (N_1181,N_1143,N_1100);
and U1182 (N_1182,N_1138,N_1142);
and U1183 (N_1183,N_1139,N_1102);
nor U1184 (N_1184,N_1124,N_1145);
nand U1185 (N_1185,N_1133,N_1118);
and U1186 (N_1186,N_1131,N_1100);
or U1187 (N_1187,N_1128,N_1126);
nor U1188 (N_1188,N_1138,N_1112);
or U1189 (N_1189,N_1138,N_1145);
nand U1190 (N_1190,N_1114,N_1121);
or U1191 (N_1191,N_1123,N_1104);
nor U1192 (N_1192,N_1103,N_1105);
xnor U1193 (N_1193,N_1116,N_1130);
and U1194 (N_1194,N_1115,N_1111);
nor U1195 (N_1195,N_1103,N_1110);
and U1196 (N_1196,N_1138,N_1116);
or U1197 (N_1197,N_1121,N_1145);
nor U1198 (N_1198,N_1117,N_1113);
or U1199 (N_1199,N_1146,N_1112);
nand U1200 (N_1200,N_1169,N_1181);
nor U1201 (N_1201,N_1161,N_1185);
and U1202 (N_1202,N_1150,N_1157);
nand U1203 (N_1203,N_1166,N_1198);
nor U1204 (N_1204,N_1183,N_1177);
xnor U1205 (N_1205,N_1182,N_1197);
xor U1206 (N_1206,N_1179,N_1175);
nand U1207 (N_1207,N_1187,N_1195);
xor U1208 (N_1208,N_1190,N_1156);
nor U1209 (N_1209,N_1151,N_1180);
xor U1210 (N_1210,N_1170,N_1154);
and U1211 (N_1211,N_1152,N_1159);
nand U1212 (N_1212,N_1165,N_1171);
xnor U1213 (N_1213,N_1192,N_1193);
xnor U1214 (N_1214,N_1194,N_1167);
and U1215 (N_1215,N_1155,N_1158);
and U1216 (N_1216,N_1172,N_1164);
xor U1217 (N_1217,N_1196,N_1160);
nand U1218 (N_1218,N_1188,N_1199);
nand U1219 (N_1219,N_1184,N_1176);
nand U1220 (N_1220,N_1186,N_1173);
nand U1221 (N_1221,N_1168,N_1174);
and U1222 (N_1222,N_1189,N_1162);
or U1223 (N_1223,N_1178,N_1163);
and U1224 (N_1224,N_1191,N_1153);
and U1225 (N_1225,N_1183,N_1188);
nor U1226 (N_1226,N_1180,N_1186);
or U1227 (N_1227,N_1193,N_1155);
nand U1228 (N_1228,N_1198,N_1199);
and U1229 (N_1229,N_1191,N_1192);
nor U1230 (N_1230,N_1166,N_1150);
or U1231 (N_1231,N_1175,N_1167);
or U1232 (N_1232,N_1185,N_1164);
nor U1233 (N_1233,N_1170,N_1160);
nand U1234 (N_1234,N_1194,N_1197);
and U1235 (N_1235,N_1163,N_1164);
or U1236 (N_1236,N_1172,N_1178);
nand U1237 (N_1237,N_1165,N_1192);
nor U1238 (N_1238,N_1151,N_1158);
and U1239 (N_1239,N_1183,N_1167);
nand U1240 (N_1240,N_1184,N_1174);
nor U1241 (N_1241,N_1180,N_1183);
or U1242 (N_1242,N_1170,N_1158);
nand U1243 (N_1243,N_1189,N_1185);
xnor U1244 (N_1244,N_1184,N_1158);
or U1245 (N_1245,N_1190,N_1185);
nand U1246 (N_1246,N_1152,N_1190);
or U1247 (N_1247,N_1152,N_1169);
and U1248 (N_1248,N_1163,N_1188);
or U1249 (N_1249,N_1159,N_1155);
and U1250 (N_1250,N_1210,N_1217);
and U1251 (N_1251,N_1226,N_1225);
and U1252 (N_1252,N_1227,N_1215);
or U1253 (N_1253,N_1239,N_1220);
or U1254 (N_1254,N_1230,N_1248);
or U1255 (N_1255,N_1203,N_1204);
nor U1256 (N_1256,N_1221,N_1249);
nand U1257 (N_1257,N_1208,N_1201);
nand U1258 (N_1258,N_1232,N_1216);
nand U1259 (N_1259,N_1241,N_1209);
and U1260 (N_1260,N_1231,N_1237);
nand U1261 (N_1261,N_1234,N_1211);
or U1262 (N_1262,N_1223,N_1205);
or U1263 (N_1263,N_1212,N_1246);
or U1264 (N_1264,N_1244,N_1218);
nand U1265 (N_1265,N_1213,N_1247);
nor U1266 (N_1266,N_1228,N_1243);
and U1267 (N_1267,N_1222,N_1238);
nand U1268 (N_1268,N_1206,N_1242);
or U1269 (N_1269,N_1219,N_1245);
and U1270 (N_1270,N_1240,N_1214);
or U1271 (N_1271,N_1200,N_1229);
nor U1272 (N_1272,N_1202,N_1236);
nor U1273 (N_1273,N_1233,N_1224);
xnor U1274 (N_1274,N_1235,N_1207);
and U1275 (N_1275,N_1206,N_1236);
nand U1276 (N_1276,N_1215,N_1208);
nor U1277 (N_1277,N_1243,N_1211);
or U1278 (N_1278,N_1213,N_1234);
nor U1279 (N_1279,N_1234,N_1223);
and U1280 (N_1280,N_1208,N_1218);
and U1281 (N_1281,N_1217,N_1228);
xnor U1282 (N_1282,N_1243,N_1205);
nand U1283 (N_1283,N_1247,N_1214);
nand U1284 (N_1284,N_1204,N_1222);
xor U1285 (N_1285,N_1207,N_1205);
and U1286 (N_1286,N_1211,N_1203);
and U1287 (N_1287,N_1231,N_1215);
nor U1288 (N_1288,N_1249,N_1205);
or U1289 (N_1289,N_1204,N_1210);
xor U1290 (N_1290,N_1232,N_1234);
nor U1291 (N_1291,N_1207,N_1200);
and U1292 (N_1292,N_1209,N_1206);
xnor U1293 (N_1293,N_1225,N_1223);
and U1294 (N_1294,N_1248,N_1222);
nor U1295 (N_1295,N_1237,N_1224);
nor U1296 (N_1296,N_1213,N_1243);
or U1297 (N_1297,N_1240,N_1202);
nor U1298 (N_1298,N_1214,N_1246);
or U1299 (N_1299,N_1218,N_1229);
or U1300 (N_1300,N_1288,N_1289);
xor U1301 (N_1301,N_1277,N_1281);
or U1302 (N_1302,N_1270,N_1258);
nor U1303 (N_1303,N_1296,N_1265);
nor U1304 (N_1304,N_1278,N_1268);
nand U1305 (N_1305,N_1276,N_1294);
or U1306 (N_1306,N_1252,N_1263);
and U1307 (N_1307,N_1297,N_1272);
and U1308 (N_1308,N_1266,N_1250);
nand U1309 (N_1309,N_1280,N_1271);
and U1310 (N_1310,N_1275,N_1257);
or U1311 (N_1311,N_1290,N_1256);
and U1312 (N_1312,N_1253,N_1273);
or U1313 (N_1313,N_1283,N_1262);
or U1314 (N_1314,N_1254,N_1285);
nor U1315 (N_1315,N_1282,N_1255);
nor U1316 (N_1316,N_1292,N_1293);
nand U1317 (N_1317,N_1295,N_1269);
or U1318 (N_1318,N_1284,N_1287);
nor U1319 (N_1319,N_1261,N_1259);
or U1320 (N_1320,N_1299,N_1260);
nor U1321 (N_1321,N_1274,N_1279);
xnor U1322 (N_1322,N_1267,N_1264);
nor U1323 (N_1323,N_1286,N_1291);
nand U1324 (N_1324,N_1251,N_1298);
xor U1325 (N_1325,N_1297,N_1251);
and U1326 (N_1326,N_1291,N_1252);
or U1327 (N_1327,N_1264,N_1284);
xnor U1328 (N_1328,N_1277,N_1252);
nand U1329 (N_1329,N_1289,N_1279);
or U1330 (N_1330,N_1272,N_1289);
or U1331 (N_1331,N_1281,N_1250);
nor U1332 (N_1332,N_1256,N_1265);
or U1333 (N_1333,N_1281,N_1287);
nor U1334 (N_1334,N_1266,N_1284);
nor U1335 (N_1335,N_1276,N_1280);
and U1336 (N_1336,N_1261,N_1264);
nor U1337 (N_1337,N_1290,N_1273);
or U1338 (N_1338,N_1274,N_1291);
and U1339 (N_1339,N_1278,N_1295);
nor U1340 (N_1340,N_1288,N_1252);
and U1341 (N_1341,N_1273,N_1299);
nand U1342 (N_1342,N_1265,N_1262);
nand U1343 (N_1343,N_1299,N_1288);
and U1344 (N_1344,N_1282,N_1279);
or U1345 (N_1345,N_1272,N_1284);
nand U1346 (N_1346,N_1294,N_1252);
nor U1347 (N_1347,N_1290,N_1250);
nand U1348 (N_1348,N_1273,N_1277);
xor U1349 (N_1349,N_1277,N_1264);
nor U1350 (N_1350,N_1338,N_1313);
and U1351 (N_1351,N_1342,N_1346);
nand U1352 (N_1352,N_1305,N_1323);
or U1353 (N_1353,N_1320,N_1303);
or U1354 (N_1354,N_1332,N_1324);
nor U1355 (N_1355,N_1339,N_1343);
or U1356 (N_1356,N_1306,N_1318);
nor U1357 (N_1357,N_1341,N_1344);
nor U1358 (N_1358,N_1331,N_1326);
and U1359 (N_1359,N_1314,N_1304);
or U1360 (N_1360,N_1302,N_1307);
or U1361 (N_1361,N_1300,N_1321);
nor U1362 (N_1362,N_1322,N_1301);
xor U1363 (N_1363,N_1311,N_1348);
nand U1364 (N_1364,N_1315,N_1309);
xnor U1365 (N_1365,N_1319,N_1310);
and U1366 (N_1366,N_1336,N_1308);
and U1367 (N_1367,N_1334,N_1312);
nand U1368 (N_1368,N_1317,N_1330);
or U1369 (N_1369,N_1337,N_1328);
nand U1370 (N_1370,N_1349,N_1347);
nor U1371 (N_1371,N_1335,N_1316);
nor U1372 (N_1372,N_1325,N_1345);
or U1373 (N_1373,N_1329,N_1333);
or U1374 (N_1374,N_1327,N_1340);
xnor U1375 (N_1375,N_1309,N_1338);
nand U1376 (N_1376,N_1327,N_1324);
or U1377 (N_1377,N_1345,N_1330);
and U1378 (N_1378,N_1323,N_1302);
nor U1379 (N_1379,N_1328,N_1308);
nand U1380 (N_1380,N_1348,N_1326);
or U1381 (N_1381,N_1346,N_1344);
nand U1382 (N_1382,N_1313,N_1330);
nor U1383 (N_1383,N_1318,N_1327);
nor U1384 (N_1384,N_1330,N_1319);
nor U1385 (N_1385,N_1337,N_1309);
or U1386 (N_1386,N_1334,N_1310);
xnor U1387 (N_1387,N_1322,N_1349);
and U1388 (N_1388,N_1312,N_1339);
and U1389 (N_1389,N_1312,N_1310);
nor U1390 (N_1390,N_1312,N_1321);
nand U1391 (N_1391,N_1339,N_1303);
and U1392 (N_1392,N_1333,N_1330);
nand U1393 (N_1393,N_1344,N_1339);
and U1394 (N_1394,N_1315,N_1323);
or U1395 (N_1395,N_1339,N_1346);
nand U1396 (N_1396,N_1338,N_1308);
nand U1397 (N_1397,N_1325,N_1319);
and U1398 (N_1398,N_1345,N_1347);
or U1399 (N_1399,N_1306,N_1328);
and U1400 (N_1400,N_1397,N_1356);
and U1401 (N_1401,N_1371,N_1350);
and U1402 (N_1402,N_1399,N_1389);
and U1403 (N_1403,N_1380,N_1384);
nand U1404 (N_1404,N_1374,N_1396);
nor U1405 (N_1405,N_1369,N_1357);
nand U1406 (N_1406,N_1362,N_1372);
nand U1407 (N_1407,N_1375,N_1354);
or U1408 (N_1408,N_1391,N_1378);
nor U1409 (N_1409,N_1383,N_1353);
and U1410 (N_1410,N_1367,N_1359);
xor U1411 (N_1411,N_1382,N_1394);
or U1412 (N_1412,N_1386,N_1388);
and U1413 (N_1413,N_1398,N_1392);
or U1414 (N_1414,N_1363,N_1377);
and U1415 (N_1415,N_1376,N_1379);
and U1416 (N_1416,N_1352,N_1390);
or U1417 (N_1417,N_1361,N_1395);
or U1418 (N_1418,N_1366,N_1364);
or U1419 (N_1419,N_1360,N_1373);
nand U1420 (N_1420,N_1368,N_1393);
and U1421 (N_1421,N_1385,N_1358);
nand U1422 (N_1422,N_1355,N_1381);
nor U1423 (N_1423,N_1387,N_1351);
nand U1424 (N_1424,N_1365,N_1370);
nor U1425 (N_1425,N_1394,N_1393);
nand U1426 (N_1426,N_1386,N_1393);
or U1427 (N_1427,N_1353,N_1369);
nor U1428 (N_1428,N_1378,N_1389);
and U1429 (N_1429,N_1399,N_1367);
nor U1430 (N_1430,N_1368,N_1371);
and U1431 (N_1431,N_1373,N_1361);
or U1432 (N_1432,N_1370,N_1389);
nand U1433 (N_1433,N_1391,N_1394);
nand U1434 (N_1434,N_1375,N_1394);
nand U1435 (N_1435,N_1381,N_1391);
xor U1436 (N_1436,N_1382,N_1352);
xor U1437 (N_1437,N_1373,N_1358);
and U1438 (N_1438,N_1375,N_1360);
or U1439 (N_1439,N_1387,N_1390);
xnor U1440 (N_1440,N_1371,N_1367);
and U1441 (N_1441,N_1392,N_1386);
nand U1442 (N_1442,N_1384,N_1378);
xnor U1443 (N_1443,N_1390,N_1355);
nor U1444 (N_1444,N_1383,N_1350);
nand U1445 (N_1445,N_1361,N_1362);
or U1446 (N_1446,N_1368,N_1373);
or U1447 (N_1447,N_1355,N_1378);
and U1448 (N_1448,N_1360,N_1387);
nor U1449 (N_1449,N_1372,N_1381);
xor U1450 (N_1450,N_1440,N_1433);
nor U1451 (N_1451,N_1429,N_1422);
and U1452 (N_1452,N_1442,N_1435);
or U1453 (N_1453,N_1445,N_1401);
nor U1454 (N_1454,N_1409,N_1404);
nand U1455 (N_1455,N_1431,N_1411);
or U1456 (N_1456,N_1423,N_1439);
nor U1457 (N_1457,N_1418,N_1412);
nor U1458 (N_1458,N_1419,N_1416);
or U1459 (N_1459,N_1446,N_1408);
or U1460 (N_1460,N_1405,N_1448);
nor U1461 (N_1461,N_1427,N_1434);
xnor U1462 (N_1462,N_1402,N_1430);
xnor U1463 (N_1463,N_1403,N_1428);
and U1464 (N_1464,N_1413,N_1424);
nor U1465 (N_1465,N_1406,N_1449);
nor U1466 (N_1466,N_1400,N_1407);
nand U1467 (N_1467,N_1414,N_1415);
and U1468 (N_1468,N_1438,N_1443);
and U1469 (N_1469,N_1437,N_1432);
or U1470 (N_1470,N_1417,N_1447);
or U1471 (N_1471,N_1410,N_1436);
nand U1472 (N_1472,N_1441,N_1420);
nand U1473 (N_1473,N_1444,N_1421);
or U1474 (N_1474,N_1425,N_1426);
and U1475 (N_1475,N_1407,N_1446);
and U1476 (N_1476,N_1447,N_1414);
nor U1477 (N_1477,N_1401,N_1425);
nand U1478 (N_1478,N_1405,N_1442);
or U1479 (N_1479,N_1426,N_1408);
nand U1480 (N_1480,N_1429,N_1440);
or U1481 (N_1481,N_1422,N_1425);
nor U1482 (N_1482,N_1402,N_1431);
or U1483 (N_1483,N_1423,N_1426);
and U1484 (N_1484,N_1418,N_1415);
nor U1485 (N_1485,N_1412,N_1400);
and U1486 (N_1486,N_1438,N_1408);
xnor U1487 (N_1487,N_1409,N_1407);
nor U1488 (N_1488,N_1438,N_1406);
and U1489 (N_1489,N_1443,N_1445);
xnor U1490 (N_1490,N_1401,N_1411);
and U1491 (N_1491,N_1415,N_1428);
nand U1492 (N_1492,N_1440,N_1438);
nand U1493 (N_1493,N_1435,N_1440);
xor U1494 (N_1494,N_1412,N_1407);
and U1495 (N_1495,N_1440,N_1447);
or U1496 (N_1496,N_1407,N_1425);
or U1497 (N_1497,N_1437,N_1422);
nor U1498 (N_1498,N_1414,N_1421);
nor U1499 (N_1499,N_1412,N_1437);
or U1500 (N_1500,N_1455,N_1470);
nand U1501 (N_1501,N_1467,N_1471);
nor U1502 (N_1502,N_1474,N_1459);
xnor U1503 (N_1503,N_1468,N_1458);
or U1504 (N_1504,N_1484,N_1464);
nor U1505 (N_1505,N_1476,N_1486);
and U1506 (N_1506,N_1485,N_1489);
nand U1507 (N_1507,N_1450,N_1483);
or U1508 (N_1508,N_1498,N_1496);
nor U1509 (N_1509,N_1457,N_1481);
and U1510 (N_1510,N_1475,N_1478);
nor U1511 (N_1511,N_1488,N_1466);
and U1512 (N_1512,N_1454,N_1463);
and U1513 (N_1513,N_1461,N_1465);
xor U1514 (N_1514,N_1456,N_1472);
and U1515 (N_1515,N_1473,N_1492);
or U1516 (N_1516,N_1479,N_1451);
or U1517 (N_1517,N_1495,N_1487);
and U1518 (N_1518,N_1482,N_1469);
or U1519 (N_1519,N_1497,N_1494);
or U1520 (N_1520,N_1480,N_1477);
nor U1521 (N_1521,N_1460,N_1490);
nor U1522 (N_1522,N_1462,N_1493);
xor U1523 (N_1523,N_1491,N_1453);
nor U1524 (N_1524,N_1499,N_1452);
or U1525 (N_1525,N_1489,N_1473);
xnor U1526 (N_1526,N_1468,N_1482);
nand U1527 (N_1527,N_1452,N_1462);
and U1528 (N_1528,N_1458,N_1453);
and U1529 (N_1529,N_1460,N_1484);
and U1530 (N_1530,N_1485,N_1498);
or U1531 (N_1531,N_1495,N_1484);
or U1532 (N_1532,N_1469,N_1477);
or U1533 (N_1533,N_1475,N_1485);
xor U1534 (N_1534,N_1497,N_1464);
nand U1535 (N_1535,N_1470,N_1468);
or U1536 (N_1536,N_1485,N_1496);
nand U1537 (N_1537,N_1499,N_1483);
and U1538 (N_1538,N_1460,N_1470);
and U1539 (N_1539,N_1472,N_1487);
and U1540 (N_1540,N_1454,N_1460);
nor U1541 (N_1541,N_1491,N_1462);
or U1542 (N_1542,N_1499,N_1466);
nor U1543 (N_1543,N_1476,N_1461);
nor U1544 (N_1544,N_1497,N_1466);
nor U1545 (N_1545,N_1456,N_1467);
nand U1546 (N_1546,N_1486,N_1487);
and U1547 (N_1547,N_1470,N_1497);
nand U1548 (N_1548,N_1467,N_1452);
and U1549 (N_1549,N_1473,N_1454);
or U1550 (N_1550,N_1517,N_1527);
or U1551 (N_1551,N_1530,N_1531);
and U1552 (N_1552,N_1523,N_1504);
nand U1553 (N_1553,N_1532,N_1500);
xor U1554 (N_1554,N_1542,N_1501);
nand U1555 (N_1555,N_1529,N_1522);
or U1556 (N_1556,N_1545,N_1503);
or U1557 (N_1557,N_1538,N_1524);
nand U1558 (N_1558,N_1510,N_1508);
or U1559 (N_1559,N_1546,N_1549);
nand U1560 (N_1560,N_1543,N_1533);
or U1561 (N_1561,N_1536,N_1547);
or U1562 (N_1562,N_1514,N_1502);
or U1563 (N_1563,N_1539,N_1534);
nor U1564 (N_1564,N_1540,N_1528);
nand U1565 (N_1565,N_1505,N_1548);
or U1566 (N_1566,N_1509,N_1535);
nand U1567 (N_1567,N_1511,N_1526);
or U1568 (N_1568,N_1521,N_1525);
nor U1569 (N_1569,N_1518,N_1541);
or U1570 (N_1570,N_1515,N_1520);
nand U1571 (N_1571,N_1506,N_1507);
nand U1572 (N_1572,N_1513,N_1519);
or U1573 (N_1573,N_1512,N_1544);
nor U1574 (N_1574,N_1516,N_1537);
nand U1575 (N_1575,N_1537,N_1501);
xor U1576 (N_1576,N_1537,N_1504);
nand U1577 (N_1577,N_1546,N_1507);
and U1578 (N_1578,N_1544,N_1547);
nor U1579 (N_1579,N_1537,N_1523);
and U1580 (N_1580,N_1519,N_1508);
or U1581 (N_1581,N_1507,N_1517);
nand U1582 (N_1582,N_1509,N_1522);
nand U1583 (N_1583,N_1544,N_1522);
xnor U1584 (N_1584,N_1503,N_1531);
and U1585 (N_1585,N_1537,N_1538);
and U1586 (N_1586,N_1507,N_1509);
nor U1587 (N_1587,N_1512,N_1533);
nand U1588 (N_1588,N_1533,N_1516);
or U1589 (N_1589,N_1501,N_1524);
and U1590 (N_1590,N_1530,N_1540);
and U1591 (N_1591,N_1508,N_1534);
or U1592 (N_1592,N_1512,N_1507);
or U1593 (N_1593,N_1521,N_1503);
and U1594 (N_1594,N_1519,N_1535);
nor U1595 (N_1595,N_1500,N_1529);
and U1596 (N_1596,N_1532,N_1517);
and U1597 (N_1597,N_1520,N_1506);
nor U1598 (N_1598,N_1502,N_1546);
or U1599 (N_1599,N_1516,N_1502);
and U1600 (N_1600,N_1588,N_1581);
and U1601 (N_1601,N_1576,N_1567);
and U1602 (N_1602,N_1598,N_1555);
nand U1603 (N_1603,N_1582,N_1557);
and U1604 (N_1604,N_1589,N_1596);
xnor U1605 (N_1605,N_1561,N_1595);
or U1606 (N_1606,N_1571,N_1554);
nand U1607 (N_1607,N_1550,N_1594);
nand U1608 (N_1608,N_1578,N_1579);
or U1609 (N_1609,N_1570,N_1558);
and U1610 (N_1610,N_1593,N_1569);
nor U1611 (N_1611,N_1551,N_1586);
nand U1612 (N_1612,N_1559,N_1575);
nand U1613 (N_1613,N_1580,N_1584);
and U1614 (N_1614,N_1572,N_1583);
nor U1615 (N_1615,N_1574,N_1560);
and U1616 (N_1616,N_1556,N_1597);
nor U1617 (N_1617,N_1587,N_1599);
nand U1618 (N_1618,N_1585,N_1552);
xor U1619 (N_1619,N_1577,N_1568);
or U1620 (N_1620,N_1553,N_1590);
xor U1621 (N_1621,N_1566,N_1562);
and U1622 (N_1622,N_1564,N_1592);
xnor U1623 (N_1623,N_1563,N_1591);
and U1624 (N_1624,N_1573,N_1565);
or U1625 (N_1625,N_1554,N_1552);
nand U1626 (N_1626,N_1565,N_1592);
nor U1627 (N_1627,N_1578,N_1582);
and U1628 (N_1628,N_1593,N_1582);
nor U1629 (N_1629,N_1565,N_1560);
and U1630 (N_1630,N_1575,N_1597);
nor U1631 (N_1631,N_1586,N_1595);
nor U1632 (N_1632,N_1586,N_1589);
xor U1633 (N_1633,N_1593,N_1599);
and U1634 (N_1634,N_1579,N_1593);
or U1635 (N_1635,N_1571,N_1565);
and U1636 (N_1636,N_1581,N_1557);
or U1637 (N_1637,N_1598,N_1560);
or U1638 (N_1638,N_1570,N_1577);
or U1639 (N_1639,N_1564,N_1581);
and U1640 (N_1640,N_1569,N_1597);
nand U1641 (N_1641,N_1557,N_1598);
and U1642 (N_1642,N_1579,N_1573);
or U1643 (N_1643,N_1560,N_1597);
nand U1644 (N_1644,N_1596,N_1556);
and U1645 (N_1645,N_1555,N_1596);
xnor U1646 (N_1646,N_1564,N_1561);
xnor U1647 (N_1647,N_1598,N_1593);
nor U1648 (N_1648,N_1572,N_1587);
and U1649 (N_1649,N_1595,N_1566);
xor U1650 (N_1650,N_1601,N_1607);
or U1651 (N_1651,N_1623,N_1612);
and U1652 (N_1652,N_1631,N_1622);
or U1653 (N_1653,N_1625,N_1621);
and U1654 (N_1654,N_1602,N_1608);
nand U1655 (N_1655,N_1635,N_1628);
or U1656 (N_1656,N_1637,N_1606);
and U1657 (N_1657,N_1649,N_1603);
nor U1658 (N_1658,N_1604,N_1624);
nand U1659 (N_1659,N_1615,N_1626);
or U1660 (N_1660,N_1647,N_1643);
and U1661 (N_1661,N_1613,N_1632);
nor U1662 (N_1662,N_1609,N_1648);
and U1663 (N_1663,N_1640,N_1630);
nor U1664 (N_1664,N_1645,N_1634);
and U1665 (N_1665,N_1618,N_1641);
nand U1666 (N_1666,N_1605,N_1614);
xnor U1667 (N_1667,N_1610,N_1642);
nor U1668 (N_1668,N_1636,N_1617);
and U1669 (N_1669,N_1619,N_1638);
and U1670 (N_1670,N_1639,N_1611);
nor U1671 (N_1671,N_1620,N_1627);
and U1672 (N_1672,N_1629,N_1646);
nor U1673 (N_1673,N_1633,N_1616);
or U1674 (N_1674,N_1600,N_1644);
nand U1675 (N_1675,N_1634,N_1614);
or U1676 (N_1676,N_1621,N_1627);
nand U1677 (N_1677,N_1644,N_1646);
nand U1678 (N_1678,N_1641,N_1607);
nand U1679 (N_1679,N_1601,N_1616);
and U1680 (N_1680,N_1630,N_1618);
nand U1681 (N_1681,N_1600,N_1643);
or U1682 (N_1682,N_1619,N_1620);
nand U1683 (N_1683,N_1644,N_1632);
and U1684 (N_1684,N_1648,N_1627);
and U1685 (N_1685,N_1625,N_1617);
nor U1686 (N_1686,N_1615,N_1631);
or U1687 (N_1687,N_1612,N_1601);
or U1688 (N_1688,N_1620,N_1640);
nor U1689 (N_1689,N_1635,N_1648);
nand U1690 (N_1690,N_1649,N_1637);
nand U1691 (N_1691,N_1601,N_1610);
nor U1692 (N_1692,N_1640,N_1616);
nor U1693 (N_1693,N_1612,N_1647);
and U1694 (N_1694,N_1611,N_1602);
nand U1695 (N_1695,N_1643,N_1615);
nand U1696 (N_1696,N_1649,N_1607);
xor U1697 (N_1697,N_1614,N_1638);
and U1698 (N_1698,N_1634,N_1630);
or U1699 (N_1699,N_1612,N_1604);
or U1700 (N_1700,N_1671,N_1688);
or U1701 (N_1701,N_1653,N_1669);
nand U1702 (N_1702,N_1683,N_1663);
and U1703 (N_1703,N_1696,N_1691);
nor U1704 (N_1704,N_1687,N_1660);
xnor U1705 (N_1705,N_1667,N_1686);
nor U1706 (N_1706,N_1665,N_1697);
or U1707 (N_1707,N_1680,N_1659);
and U1708 (N_1708,N_1664,N_1666);
nand U1709 (N_1709,N_1679,N_1672);
nor U1710 (N_1710,N_1651,N_1658);
nand U1711 (N_1711,N_1661,N_1650);
xnor U1712 (N_1712,N_1673,N_1690);
or U1713 (N_1713,N_1674,N_1675);
nor U1714 (N_1714,N_1662,N_1677);
nor U1715 (N_1715,N_1698,N_1681);
and U1716 (N_1716,N_1655,N_1693);
nand U1717 (N_1717,N_1676,N_1695);
and U1718 (N_1718,N_1656,N_1699);
or U1719 (N_1719,N_1689,N_1668);
or U1720 (N_1720,N_1692,N_1685);
and U1721 (N_1721,N_1694,N_1682);
nand U1722 (N_1722,N_1652,N_1670);
nor U1723 (N_1723,N_1684,N_1678);
nor U1724 (N_1724,N_1654,N_1657);
or U1725 (N_1725,N_1661,N_1683);
nand U1726 (N_1726,N_1667,N_1657);
nor U1727 (N_1727,N_1699,N_1665);
xor U1728 (N_1728,N_1677,N_1652);
nor U1729 (N_1729,N_1655,N_1658);
nor U1730 (N_1730,N_1681,N_1663);
and U1731 (N_1731,N_1680,N_1672);
nand U1732 (N_1732,N_1682,N_1687);
xnor U1733 (N_1733,N_1675,N_1661);
and U1734 (N_1734,N_1666,N_1677);
nor U1735 (N_1735,N_1653,N_1676);
nand U1736 (N_1736,N_1678,N_1669);
nor U1737 (N_1737,N_1671,N_1655);
nand U1738 (N_1738,N_1684,N_1652);
or U1739 (N_1739,N_1680,N_1653);
nor U1740 (N_1740,N_1682,N_1662);
or U1741 (N_1741,N_1673,N_1683);
xor U1742 (N_1742,N_1669,N_1664);
and U1743 (N_1743,N_1689,N_1657);
and U1744 (N_1744,N_1666,N_1654);
xnor U1745 (N_1745,N_1652,N_1674);
nand U1746 (N_1746,N_1664,N_1685);
nor U1747 (N_1747,N_1672,N_1697);
and U1748 (N_1748,N_1681,N_1664);
and U1749 (N_1749,N_1667,N_1665);
or U1750 (N_1750,N_1749,N_1722);
xnor U1751 (N_1751,N_1725,N_1709);
nor U1752 (N_1752,N_1726,N_1728);
or U1753 (N_1753,N_1731,N_1704);
or U1754 (N_1754,N_1707,N_1740);
or U1755 (N_1755,N_1714,N_1713);
or U1756 (N_1756,N_1717,N_1746);
and U1757 (N_1757,N_1734,N_1724);
and U1758 (N_1758,N_1738,N_1711);
nand U1759 (N_1759,N_1729,N_1737);
nor U1760 (N_1760,N_1742,N_1747);
nor U1761 (N_1761,N_1702,N_1708);
nand U1762 (N_1762,N_1712,N_1735);
or U1763 (N_1763,N_1745,N_1716);
or U1764 (N_1764,N_1727,N_1733);
and U1765 (N_1765,N_1723,N_1718);
nor U1766 (N_1766,N_1744,N_1706);
nand U1767 (N_1767,N_1705,N_1721);
or U1768 (N_1768,N_1703,N_1701);
or U1769 (N_1769,N_1736,N_1743);
nor U1770 (N_1770,N_1710,N_1730);
nor U1771 (N_1771,N_1748,N_1720);
or U1772 (N_1772,N_1715,N_1700);
and U1773 (N_1773,N_1741,N_1732);
and U1774 (N_1774,N_1739,N_1719);
and U1775 (N_1775,N_1716,N_1705);
nor U1776 (N_1776,N_1734,N_1720);
nand U1777 (N_1777,N_1700,N_1748);
nand U1778 (N_1778,N_1729,N_1701);
or U1779 (N_1779,N_1733,N_1734);
nor U1780 (N_1780,N_1701,N_1747);
nor U1781 (N_1781,N_1744,N_1740);
nand U1782 (N_1782,N_1726,N_1702);
nand U1783 (N_1783,N_1749,N_1700);
and U1784 (N_1784,N_1700,N_1727);
and U1785 (N_1785,N_1721,N_1733);
and U1786 (N_1786,N_1742,N_1706);
or U1787 (N_1787,N_1729,N_1735);
nand U1788 (N_1788,N_1703,N_1725);
or U1789 (N_1789,N_1722,N_1729);
nor U1790 (N_1790,N_1703,N_1710);
xnor U1791 (N_1791,N_1721,N_1724);
and U1792 (N_1792,N_1734,N_1700);
or U1793 (N_1793,N_1734,N_1747);
nand U1794 (N_1794,N_1715,N_1712);
nor U1795 (N_1795,N_1711,N_1707);
and U1796 (N_1796,N_1717,N_1719);
nand U1797 (N_1797,N_1700,N_1709);
nor U1798 (N_1798,N_1707,N_1721);
nor U1799 (N_1799,N_1723,N_1743);
or U1800 (N_1800,N_1758,N_1766);
and U1801 (N_1801,N_1781,N_1757);
nand U1802 (N_1802,N_1754,N_1761);
nor U1803 (N_1803,N_1774,N_1768);
and U1804 (N_1804,N_1777,N_1750);
xnor U1805 (N_1805,N_1798,N_1759);
nor U1806 (N_1806,N_1775,N_1788);
nand U1807 (N_1807,N_1796,N_1787);
or U1808 (N_1808,N_1791,N_1793);
and U1809 (N_1809,N_1785,N_1795);
nor U1810 (N_1810,N_1760,N_1769);
and U1811 (N_1811,N_1756,N_1779);
nor U1812 (N_1812,N_1794,N_1772);
nand U1813 (N_1813,N_1780,N_1762);
nand U1814 (N_1814,N_1776,N_1790);
or U1815 (N_1815,N_1752,N_1784);
nand U1816 (N_1816,N_1799,N_1765);
nor U1817 (N_1817,N_1773,N_1770);
and U1818 (N_1818,N_1792,N_1751);
nand U1819 (N_1819,N_1786,N_1767);
nor U1820 (N_1820,N_1771,N_1782);
xor U1821 (N_1821,N_1753,N_1764);
nand U1822 (N_1822,N_1797,N_1783);
or U1823 (N_1823,N_1789,N_1778);
or U1824 (N_1824,N_1763,N_1755);
nand U1825 (N_1825,N_1798,N_1752);
and U1826 (N_1826,N_1753,N_1773);
or U1827 (N_1827,N_1797,N_1758);
and U1828 (N_1828,N_1772,N_1775);
or U1829 (N_1829,N_1799,N_1766);
nand U1830 (N_1830,N_1792,N_1782);
nand U1831 (N_1831,N_1755,N_1785);
or U1832 (N_1832,N_1780,N_1760);
and U1833 (N_1833,N_1763,N_1759);
nor U1834 (N_1834,N_1766,N_1790);
nand U1835 (N_1835,N_1756,N_1761);
xnor U1836 (N_1836,N_1757,N_1769);
nand U1837 (N_1837,N_1787,N_1767);
nand U1838 (N_1838,N_1779,N_1769);
or U1839 (N_1839,N_1750,N_1755);
and U1840 (N_1840,N_1764,N_1765);
xnor U1841 (N_1841,N_1796,N_1789);
and U1842 (N_1842,N_1755,N_1769);
xor U1843 (N_1843,N_1770,N_1798);
and U1844 (N_1844,N_1775,N_1778);
and U1845 (N_1845,N_1778,N_1781);
nor U1846 (N_1846,N_1789,N_1794);
nand U1847 (N_1847,N_1762,N_1761);
nand U1848 (N_1848,N_1766,N_1777);
or U1849 (N_1849,N_1789,N_1772);
and U1850 (N_1850,N_1839,N_1801);
and U1851 (N_1851,N_1805,N_1842);
and U1852 (N_1852,N_1831,N_1809);
nand U1853 (N_1853,N_1823,N_1816);
or U1854 (N_1854,N_1811,N_1848);
or U1855 (N_1855,N_1837,N_1840);
nor U1856 (N_1856,N_1836,N_1829);
nand U1857 (N_1857,N_1802,N_1846);
xnor U1858 (N_1858,N_1844,N_1813);
and U1859 (N_1859,N_1822,N_1834);
nand U1860 (N_1860,N_1818,N_1845);
nor U1861 (N_1861,N_1827,N_1843);
nor U1862 (N_1862,N_1804,N_1815);
nor U1863 (N_1863,N_1819,N_1814);
nor U1864 (N_1864,N_1800,N_1833);
and U1865 (N_1865,N_1812,N_1832);
and U1866 (N_1866,N_1825,N_1830);
or U1867 (N_1867,N_1807,N_1803);
nand U1868 (N_1868,N_1841,N_1821);
nor U1869 (N_1869,N_1806,N_1820);
or U1870 (N_1870,N_1808,N_1810);
xnor U1871 (N_1871,N_1838,N_1817);
and U1872 (N_1872,N_1835,N_1847);
and U1873 (N_1873,N_1826,N_1824);
nor U1874 (N_1874,N_1828,N_1849);
nor U1875 (N_1875,N_1822,N_1821);
nor U1876 (N_1876,N_1839,N_1817);
nor U1877 (N_1877,N_1826,N_1812);
nand U1878 (N_1878,N_1809,N_1814);
nor U1879 (N_1879,N_1805,N_1840);
nor U1880 (N_1880,N_1821,N_1825);
xor U1881 (N_1881,N_1830,N_1817);
nor U1882 (N_1882,N_1846,N_1832);
nand U1883 (N_1883,N_1830,N_1848);
or U1884 (N_1884,N_1805,N_1801);
and U1885 (N_1885,N_1843,N_1801);
xor U1886 (N_1886,N_1803,N_1812);
and U1887 (N_1887,N_1819,N_1810);
xor U1888 (N_1888,N_1824,N_1828);
nand U1889 (N_1889,N_1803,N_1817);
nor U1890 (N_1890,N_1806,N_1812);
nor U1891 (N_1891,N_1837,N_1828);
xnor U1892 (N_1892,N_1819,N_1846);
nand U1893 (N_1893,N_1807,N_1818);
nand U1894 (N_1894,N_1813,N_1814);
and U1895 (N_1895,N_1815,N_1833);
nor U1896 (N_1896,N_1825,N_1800);
or U1897 (N_1897,N_1845,N_1827);
nor U1898 (N_1898,N_1806,N_1828);
nand U1899 (N_1899,N_1848,N_1821);
xor U1900 (N_1900,N_1883,N_1862);
and U1901 (N_1901,N_1889,N_1866);
nor U1902 (N_1902,N_1893,N_1877);
nor U1903 (N_1903,N_1867,N_1852);
xor U1904 (N_1904,N_1888,N_1887);
and U1905 (N_1905,N_1881,N_1864);
or U1906 (N_1906,N_1882,N_1884);
nand U1907 (N_1907,N_1873,N_1899);
and U1908 (N_1908,N_1851,N_1880);
or U1909 (N_1909,N_1850,N_1886);
xnor U1910 (N_1910,N_1885,N_1863);
and U1911 (N_1911,N_1856,N_1898);
and U1912 (N_1912,N_1857,N_1860);
nand U1913 (N_1913,N_1894,N_1854);
or U1914 (N_1914,N_1869,N_1891);
or U1915 (N_1915,N_1858,N_1874);
nand U1916 (N_1916,N_1897,N_1890);
and U1917 (N_1917,N_1879,N_1861);
xnor U1918 (N_1918,N_1855,N_1875);
nand U1919 (N_1919,N_1878,N_1876);
or U1920 (N_1920,N_1868,N_1871);
nor U1921 (N_1921,N_1896,N_1853);
nor U1922 (N_1922,N_1892,N_1859);
nor U1923 (N_1923,N_1895,N_1865);
nor U1924 (N_1924,N_1872,N_1870);
or U1925 (N_1925,N_1851,N_1883);
or U1926 (N_1926,N_1871,N_1878);
or U1927 (N_1927,N_1860,N_1889);
nor U1928 (N_1928,N_1869,N_1872);
or U1929 (N_1929,N_1868,N_1898);
or U1930 (N_1930,N_1874,N_1851);
and U1931 (N_1931,N_1860,N_1898);
and U1932 (N_1932,N_1888,N_1873);
nor U1933 (N_1933,N_1894,N_1890);
and U1934 (N_1934,N_1857,N_1876);
nor U1935 (N_1935,N_1864,N_1897);
nor U1936 (N_1936,N_1892,N_1878);
or U1937 (N_1937,N_1855,N_1899);
nor U1938 (N_1938,N_1868,N_1860);
and U1939 (N_1939,N_1859,N_1866);
nand U1940 (N_1940,N_1876,N_1883);
and U1941 (N_1941,N_1862,N_1865);
or U1942 (N_1942,N_1865,N_1882);
nand U1943 (N_1943,N_1854,N_1870);
xnor U1944 (N_1944,N_1870,N_1865);
or U1945 (N_1945,N_1859,N_1885);
or U1946 (N_1946,N_1853,N_1871);
or U1947 (N_1947,N_1879,N_1883);
nand U1948 (N_1948,N_1872,N_1888);
or U1949 (N_1949,N_1874,N_1888);
nand U1950 (N_1950,N_1945,N_1905);
and U1951 (N_1951,N_1913,N_1923);
nand U1952 (N_1952,N_1948,N_1947);
or U1953 (N_1953,N_1944,N_1933);
nor U1954 (N_1954,N_1937,N_1911);
nand U1955 (N_1955,N_1918,N_1949);
or U1956 (N_1956,N_1921,N_1939);
or U1957 (N_1957,N_1930,N_1926);
nand U1958 (N_1958,N_1919,N_1925);
xor U1959 (N_1959,N_1936,N_1932);
nor U1960 (N_1960,N_1941,N_1927);
nand U1961 (N_1961,N_1931,N_1914);
and U1962 (N_1962,N_1942,N_1912);
and U1963 (N_1963,N_1929,N_1917);
or U1964 (N_1964,N_1935,N_1910);
xnor U1965 (N_1965,N_1909,N_1916);
nor U1966 (N_1966,N_1946,N_1902);
nand U1967 (N_1967,N_1922,N_1924);
xor U1968 (N_1968,N_1906,N_1904);
nor U1969 (N_1969,N_1903,N_1915);
or U1970 (N_1970,N_1900,N_1938);
and U1971 (N_1971,N_1920,N_1908);
nand U1972 (N_1972,N_1928,N_1907);
or U1973 (N_1973,N_1940,N_1901);
and U1974 (N_1974,N_1934,N_1943);
nor U1975 (N_1975,N_1909,N_1931);
and U1976 (N_1976,N_1923,N_1919);
nand U1977 (N_1977,N_1901,N_1937);
and U1978 (N_1978,N_1939,N_1922);
or U1979 (N_1979,N_1945,N_1932);
or U1980 (N_1980,N_1935,N_1928);
or U1981 (N_1981,N_1912,N_1925);
nand U1982 (N_1982,N_1942,N_1947);
or U1983 (N_1983,N_1905,N_1929);
and U1984 (N_1984,N_1925,N_1939);
and U1985 (N_1985,N_1930,N_1949);
nand U1986 (N_1986,N_1928,N_1936);
nor U1987 (N_1987,N_1941,N_1938);
nor U1988 (N_1988,N_1903,N_1927);
or U1989 (N_1989,N_1934,N_1922);
and U1990 (N_1990,N_1946,N_1932);
nor U1991 (N_1991,N_1918,N_1920);
or U1992 (N_1992,N_1910,N_1917);
nor U1993 (N_1993,N_1902,N_1932);
and U1994 (N_1994,N_1909,N_1925);
and U1995 (N_1995,N_1918,N_1924);
and U1996 (N_1996,N_1937,N_1938);
or U1997 (N_1997,N_1907,N_1918);
and U1998 (N_1998,N_1940,N_1930);
nand U1999 (N_1999,N_1919,N_1926);
nand U2000 (N_2000,N_1997,N_1992);
nor U2001 (N_2001,N_1991,N_1973);
nand U2002 (N_2002,N_1983,N_1967);
and U2003 (N_2003,N_1995,N_1987);
or U2004 (N_2004,N_1954,N_1958);
nor U2005 (N_2005,N_1981,N_1968);
nor U2006 (N_2006,N_1955,N_1972);
nor U2007 (N_2007,N_1979,N_1977);
nor U2008 (N_2008,N_1980,N_1963);
and U2009 (N_2009,N_1952,N_1998);
or U2010 (N_2010,N_1984,N_1985);
nand U2011 (N_2011,N_1976,N_1990);
or U2012 (N_2012,N_1960,N_1971);
and U2013 (N_2013,N_1982,N_1950);
and U2014 (N_2014,N_1962,N_1989);
nor U2015 (N_2015,N_1988,N_1957);
nand U2016 (N_2016,N_1994,N_1996);
nand U2017 (N_2017,N_1953,N_1993);
nor U2018 (N_2018,N_1969,N_1974);
nand U2019 (N_2019,N_1965,N_1964);
and U2020 (N_2020,N_1961,N_1978);
nor U2021 (N_2021,N_1999,N_1951);
or U2022 (N_2022,N_1975,N_1956);
or U2023 (N_2023,N_1970,N_1959);
xor U2024 (N_2024,N_1966,N_1986);
xnor U2025 (N_2025,N_1991,N_1986);
nor U2026 (N_2026,N_1958,N_1957);
and U2027 (N_2027,N_1991,N_1989);
and U2028 (N_2028,N_1958,N_1986);
xor U2029 (N_2029,N_1975,N_1993);
nor U2030 (N_2030,N_1979,N_1972);
nand U2031 (N_2031,N_1991,N_1985);
nand U2032 (N_2032,N_1979,N_1964);
xor U2033 (N_2033,N_1951,N_1968);
nand U2034 (N_2034,N_1980,N_1979);
or U2035 (N_2035,N_1983,N_1969);
nand U2036 (N_2036,N_1997,N_1958);
xnor U2037 (N_2037,N_1982,N_1951);
nor U2038 (N_2038,N_1975,N_1994);
and U2039 (N_2039,N_1963,N_1972);
nor U2040 (N_2040,N_1974,N_1950);
nand U2041 (N_2041,N_1992,N_1950);
xor U2042 (N_2042,N_1975,N_1967);
and U2043 (N_2043,N_1980,N_1971);
nand U2044 (N_2044,N_1962,N_1975);
nand U2045 (N_2045,N_1962,N_1990);
nor U2046 (N_2046,N_1967,N_1951);
or U2047 (N_2047,N_1974,N_1965);
nand U2048 (N_2048,N_1983,N_1975);
and U2049 (N_2049,N_1991,N_1988);
nor U2050 (N_2050,N_2012,N_2031);
nand U2051 (N_2051,N_2029,N_2020);
nand U2052 (N_2052,N_2003,N_2024);
nand U2053 (N_2053,N_2042,N_2019);
or U2054 (N_2054,N_2001,N_2023);
nor U2055 (N_2055,N_2009,N_2045);
nand U2056 (N_2056,N_2010,N_2005);
nand U2057 (N_2057,N_2048,N_2040);
or U2058 (N_2058,N_2006,N_2034);
nor U2059 (N_2059,N_2037,N_2028);
nand U2060 (N_2060,N_2033,N_2002);
nor U2061 (N_2061,N_2014,N_2018);
nand U2062 (N_2062,N_2022,N_2008);
or U2063 (N_2063,N_2021,N_2004);
xnor U2064 (N_2064,N_2030,N_2011);
nand U2065 (N_2065,N_2046,N_2041);
nor U2066 (N_2066,N_2044,N_2049);
or U2067 (N_2067,N_2016,N_2000);
nor U2068 (N_2068,N_2035,N_2039);
nor U2069 (N_2069,N_2036,N_2017);
nand U2070 (N_2070,N_2043,N_2047);
or U2071 (N_2071,N_2027,N_2038);
or U2072 (N_2072,N_2026,N_2025);
nand U2073 (N_2073,N_2032,N_2015);
or U2074 (N_2074,N_2013,N_2007);
or U2075 (N_2075,N_2046,N_2011);
nand U2076 (N_2076,N_2029,N_2031);
and U2077 (N_2077,N_2007,N_2039);
nor U2078 (N_2078,N_2049,N_2029);
nand U2079 (N_2079,N_2028,N_2035);
nor U2080 (N_2080,N_2013,N_2039);
nor U2081 (N_2081,N_2020,N_2044);
nor U2082 (N_2082,N_2010,N_2014);
and U2083 (N_2083,N_2020,N_2046);
nand U2084 (N_2084,N_2036,N_2008);
nand U2085 (N_2085,N_2041,N_2007);
and U2086 (N_2086,N_2042,N_2003);
nand U2087 (N_2087,N_2027,N_2044);
and U2088 (N_2088,N_2003,N_2006);
nor U2089 (N_2089,N_2033,N_2001);
or U2090 (N_2090,N_2027,N_2002);
nand U2091 (N_2091,N_2040,N_2037);
nor U2092 (N_2092,N_2013,N_2019);
xor U2093 (N_2093,N_2017,N_2022);
and U2094 (N_2094,N_2035,N_2019);
or U2095 (N_2095,N_2027,N_2001);
xor U2096 (N_2096,N_2038,N_2005);
or U2097 (N_2097,N_2033,N_2026);
and U2098 (N_2098,N_2019,N_2020);
nor U2099 (N_2099,N_2000,N_2027);
and U2100 (N_2100,N_2063,N_2060);
and U2101 (N_2101,N_2054,N_2077);
and U2102 (N_2102,N_2058,N_2050);
nor U2103 (N_2103,N_2092,N_2078);
or U2104 (N_2104,N_2080,N_2086);
nor U2105 (N_2105,N_2074,N_2084);
nand U2106 (N_2106,N_2091,N_2089);
or U2107 (N_2107,N_2061,N_2066);
or U2108 (N_2108,N_2098,N_2087);
and U2109 (N_2109,N_2070,N_2072);
xnor U2110 (N_2110,N_2099,N_2055);
nand U2111 (N_2111,N_2095,N_2088);
and U2112 (N_2112,N_2085,N_2056);
nand U2113 (N_2113,N_2071,N_2079);
xnor U2114 (N_2114,N_2068,N_2051);
nor U2115 (N_2115,N_2067,N_2062);
or U2116 (N_2116,N_2082,N_2065);
nor U2117 (N_2117,N_2097,N_2075);
nand U2118 (N_2118,N_2094,N_2090);
and U2119 (N_2119,N_2057,N_2081);
nor U2120 (N_2120,N_2064,N_2059);
or U2121 (N_2121,N_2052,N_2076);
or U2122 (N_2122,N_2073,N_2069);
or U2123 (N_2123,N_2083,N_2096);
xor U2124 (N_2124,N_2093,N_2053);
xnor U2125 (N_2125,N_2081,N_2061);
nand U2126 (N_2126,N_2095,N_2070);
nor U2127 (N_2127,N_2070,N_2097);
and U2128 (N_2128,N_2058,N_2070);
nor U2129 (N_2129,N_2081,N_2070);
nand U2130 (N_2130,N_2098,N_2064);
nand U2131 (N_2131,N_2068,N_2069);
and U2132 (N_2132,N_2055,N_2066);
and U2133 (N_2133,N_2080,N_2064);
nor U2134 (N_2134,N_2071,N_2086);
and U2135 (N_2135,N_2091,N_2083);
xor U2136 (N_2136,N_2071,N_2058);
nor U2137 (N_2137,N_2076,N_2054);
nand U2138 (N_2138,N_2086,N_2062);
nand U2139 (N_2139,N_2092,N_2095);
or U2140 (N_2140,N_2055,N_2051);
nor U2141 (N_2141,N_2058,N_2082);
and U2142 (N_2142,N_2067,N_2072);
and U2143 (N_2143,N_2076,N_2074);
nor U2144 (N_2144,N_2080,N_2054);
nor U2145 (N_2145,N_2075,N_2086);
or U2146 (N_2146,N_2056,N_2062);
xnor U2147 (N_2147,N_2061,N_2094);
or U2148 (N_2148,N_2084,N_2091);
nor U2149 (N_2149,N_2076,N_2079);
or U2150 (N_2150,N_2145,N_2126);
nor U2151 (N_2151,N_2143,N_2106);
and U2152 (N_2152,N_2133,N_2112);
nand U2153 (N_2153,N_2134,N_2104);
nand U2154 (N_2154,N_2119,N_2125);
xor U2155 (N_2155,N_2120,N_2123);
or U2156 (N_2156,N_2130,N_2121);
or U2157 (N_2157,N_2131,N_2144);
nand U2158 (N_2158,N_2117,N_2103);
nor U2159 (N_2159,N_2128,N_2108);
or U2160 (N_2160,N_2102,N_2146);
and U2161 (N_2161,N_2109,N_2141);
and U2162 (N_2162,N_2118,N_2111);
or U2163 (N_2163,N_2113,N_2139);
or U2164 (N_2164,N_2149,N_2127);
nor U2165 (N_2165,N_2124,N_2115);
or U2166 (N_2166,N_2116,N_2110);
or U2167 (N_2167,N_2137,N_2101);
and U2168 (N_2168,N_2132,N_2122);
or U2169 (N_2169,N_2105,N_2129);
nand U2170 (N_2170,N_2138,N_2147);
and U2171 (N_2171,N_2114,N_2107);
nand U2172 (N_2172,N_2135,N_2136);
nand U2173 (N_2173,N_2100,N_2142);
and U2174 (N_2174,N_2148,N_2140);
and U2175 (N_2175,N_2104,N_2123);
nand U2176 (N_2176,N_2120,N_2113);
and U2177 (N_2177,N_2133,N_2131);
or U2178 (N_2178,N_2149,N_2131);
and U2179 (N_2179,N_2104,N_2147);
and U2180 (N_2180,N_2148,N_2104);
or U2181 (N_2181,N_2130,N_2107);
nand U2182 (N_2182,N_2129,N_2119);
nor U2183 (N_2183,N_2127,N_2126);
and U2184 (N_2184,N_2138,N_2140);
nand U2185 (N_2185,N_2136,N_2113);
nand U2186 (N_2186,N_2101,N_2132);
and U2187 (N_2187,N_2140,N_2126);
or U2188 (N_2188,N_2132,N_2130);
or U2189 (N_2189,N_2100,N_2104);
nor U2190 (N_2190,N_2148,N_2109);
nand U2191 (N_2191,N_2143,N_2138);
or U2192 (N_2192,N_2122,N_2102);
nand U2193 (N_2193,N_2128,N_2141);
or U2194 (N_2194,N_2139,N_2125);
or U2195 (N_2195,N_2126,N_2115);
xnor U2196 (N_2196,N_2123,N_2132);
or U2197 (N_2197,N_2135,N_2124);
or U2198 (N_2198,N_2135,N_2104);
or U2199 (N_2199,N_2143,N_2119);
or U2200 (N_2200,N_2173,N_2161);
nand U2201 (N_2201,N_2189,N_2177);
or U2202 (N_2202,N_2155,N_2166);
and U2203 (N_2203,N_2170,N_2164);
nor U2204 (N_2204,N_2190,N_2152);
nor U2205 (N_2205,N_2192,N_2181);
and U2206 (N_2206,N_2187,N_2154);
and U2207 (N_2207,N_2162,N_2188);
or U2208 (N_2208,N_2172,N_2197);
nand U2209 (N_2209,N_2186,N_2178);
or U2210 (N_2210,N_2163,N_2176);
or U2211 (N_2211,N_2158,N_2182);
nor U2212 (N_2212,N_2175,N_2198);
nor U2213 (N_2213,N_2199,N_2179);
or U2214 (N_2214,N_2157,N_2156);
or U2215 (N_2215,N_2196,N_2167);
nand U2216 (N_2216,N_2153,N_2183);
nor U2217 (N_2217,N_2193,N_2165);
nand U2218 (N_2218,N_2194,N_2150);
xnor U2219 (N_2219,N_2168,N_2185);
or U2220 (N_2220,N_2174,N_2169);
xnor U2221 (N_2221,N_2160,N_2184);
and U2222 (N_2222,N_2191,N_2180);
xnor U2223 (N_2223,N_2151,N_2171);
nand U2224 (N_2224,N_2159,N_2195);
and U2225 (N_2225,N_2153,N_2195);
or U2226 (N_2226,N_2199,N_2189);
nor U2227 (N_2227,N_2172,N_2160);
nor U2228 (N_2228,N_2153,N_2185);
nor U2229 (N_2229,N_2198,N_2171);
and U2230 (N_2230,N_2150,N_2171);
or U2231 (N_2231,N_2190,N_2191);
and U2232 (N_2232,N_2193,N_2182);
or U2233 (N_2233,N_2158,N_2163);
and U2234 (N_2234,N_2191,N_2183);
or U2235 (N_2235,N_2162,N_2185);
or U2236 (N_2236,N_2174,N_2157);
and U2237 (N_2237,N_2176,N_2161);
and U2238 (N_2238,N_2177,N_2173);
nor U2239 (N_2239,N_2197,N_2181);
or U2240 (N_2240,N_2194,N_2160);
nor U2241 (N_2241,N_2184,N_2185);
nor U2242 (N_2242,N_2176,N_2199);
and U2243 (N_2243,N_2176,N_2174);
nand U2244 (N_2244,N_2152,N_2199);
and U2245 (N_2245,N_2197,N_2183);
or U2246 (N_2246,N_2170,N_2173);
xor U2247 (N_2247,N_2158,N_2188);
nor U2248 (N_2248,N_2179,N_2183);
nand U2249 (N_2249,N_2159,N_2193);
nand U2250 (N_2250,N_2209,N_2232);
and U2251 (N_2251,N_2216,N_2218);
or U2252 (N_2252,N_2238,N_2231);
nand U2253 (N_2253,N_2215,N_2230);
nand U2254 (N_2254,N_2233,N_2223);
nand U2255 (N_2255,N_2239,N_2249);
or U2256 (N_2256,N_2212,N_2242);
nand U2257 (N_2257,N_2246,N_2247);
nand U2258 (N_2258,N_2205,N_2227);
and U2259 (N_2259,N_2213,N_2225);
nor U2260 (N_2260,N_2222,N_2217);
or U2261 (N_2261,N_2203,N_2210);
nand U2262 (N_2262,N_2200,N_2206);
nand U2263 (N_2263,N_2229,N_2245);
nand U2264 (N_2264,N_2243,N_2214);
nand U2265 (N_2265,N_2234,N_2237);
or U2266 (N_2266,N_2202,N_2236);
or U2267 (N_2267,N_2208,N_2201);
xnor U2268 (N_2268,N_2241,N_2235);
and U2269 (N_2269,N_2240,N_2220);
nand U2270 (N_2270,N_2248,N_2204);
nand U2271 (N_2271,N_2221,N_2224);
nor U2272 (N_2272,N_2226,N_2211);
nor U2273 (N_2273,N_2219,N_2244);
nor U2274 (N_2274,N_2207,N_2228);
and U2275 (N_2275,N_2217,N_2211);
or U2276 (N_2276,N_2232,N_2223);
nand U2277 (N_2277,N_2217,N_2210);
nand U2278 (N_2278,N_2212,N_2240);
nor U2279 (N_2279,N_2246,N_2208);
or U2280 (N_2280,N_2244,N_2200);
nand U2281 (N_2281,N_2230,N_2218);
and U2282 (N_2282,N_2208,N_2228);
or U2283 (N_2283,N_2221,N_2243);
nor U2284 (N_2284,N_2224,N_2230);
or U2285 (N_2285,N_2229,N_2233);
nor U2286 (N_2286,N_2206,N_2218);
and U2287 (N_2287,N_2217,N_2219);
or U2288 (N_2288,N_2207,N_2238);
and U2289 (N_2289,N_2238,N_2201);
or U2290 (N_2290,N_2205,N_2232);
and U2291 (N_2291,N_2209,N_2233);
and U2292 (N_2292,N_2209,N_2247);
and U2293 (N_2293,N_2211,N_2214);
and U2294 (N_2294,N_2247,N_2201);
nor U2295 (N_2295,N_2205,N_2228);
nor U2296 (N_2296,N_2202,N_2215);
xnor U2297 (N_2297,N_2221,N_2244);
or U2298 (N_2298,N_2207,N_2245);
nand U2299 (N_2299,N_2200,N_2208);
nor U2300 (N_2300,N_2254,N_2272);
and U2301 (N_2301,N_2286,N_2285);
xor U2302 (N_2302,N_2298,N_2260);
nand U2303 (N_2303,N_2282,N_2275);
and U2304 (N_2304,N_2288,N_2263);
and U2305 (N_2305,N_2261,N_2297);
and U2306 (N_2306,N_2293,N_2280);
and U2307 (N_2307,N_2281,N_2256);
nor U2308 (N_2308,N_2252,N_2292);
or U2309 (N_2309,N_2267,N_2287);
nor U2310 (N_2310,N_2294,N_2290);
and U2311 (N_2311,N_2250,N_2259);
nor U2312 (N_2312,N_2266,N_2295);
nor U2313 (N_2313,N_2283,N_2278);
nor U2314 (N_2314,N_2257,N_2264);
nor U2315 (N_2315,N_2251,N_2270);
or U2316 (N_2316,N_2276,N_2289);
xor U2317 (N_2317,N_2273,N_2277);
nand U2318 (N_2318,N_2279,N_2258);
or U2319 (N_2319,N_2253,N_2271);
nand U2320 (N_2320,N_2274,N_2268);
nor U2321 (N_2321,N_2269,N_2299);
or U2322 (N_2322,N_2284,N_2265);
nor U2323 (N_2323,N_2255,N_2291);
and U2324 (N_2324,N_2262,N_2296);
nand U2325 (N_2325,N_2269,N_2250);
or U2326 (N_2326,N_2262,N_2277);
and U2327 (N_2327,N_2274,N_2262);
or U2328 (N_2328,N_2296,N_2290);
and U2329 (N_2329,N_2255,N_2267);
or U2330 (N_2330,N_2290,N_2252);
xor U2331 (N_2331,N_2270,N_2292);
nand U2332 (N_2332,N_2286,N_2250);
or U2333 (N_2333,N_2253,N_2282);
and U2334 (N_2334,N_2274,N_2284);
or U2335 (N_2335,N_2278,N_2251);
nand U2336 (N_2336,N_2270,N_2285);
or U2337 (N_2337,N_2291,N_2295);
nor U2338 (N_2338,N_2282,N_2297);
nand U2339 (N_2339,N_2258,N_2292);
xnor U2340 (N_2340,N_2252,N_2257);
or U2341 (N_2341,N_2282,N_2254);
xor U2342 (N_2342,N_2263,N_2290);
nand U2343 (N_2343,N_2261,N_2258);
nor U2344 (N_2344,N_2252,N_2278);
and U2345 (N_2345,N_2273,N_2252);
and U2346 (N_2346,N_2284,N_2264);
and U2347 (N_2347,N_2280,N_2289);
and U2348 (N_2348,N_2254,N_2283);
nor U2349 (N_2349,N_2294,N_2269);
nor U2350 (N_2350,N_2314,N_2330);
and U2351 (N_2351,N_2307,N_2349);
and U2352 (N_2352,N_2305,N_2343);
and U2353 (N_2353,N_2332,N_2312);
and U2354 (N_2354,N_2334,N_2338);
and U2355 (N_2355,N_2313,N_2316);
and U2356 (N_2356,N_2309,N_2348);
nand U2357 (N_2357,N_2331,N_2323);
or U2358 (N_2358,N_2319,N_2344);
nand U2359 (N_2359,N_2327,N_2341);
xnor U2360 (N_2360,N_2339,N_2337);
xor U2361 (N_2361,N_2318,N_2345);
xnor U2362 (N_2362,N_2310,N_2321);
or U2363 (N_2363,N_2317,N_2328);
or U2364 (N_2364,N_2306,N_2335);
xnor U2365 (N_2365,N_2308,N_2336);
and U2366 (N_2366,N_2303,N_2342);
nand U2367 (N_2367,N_2325,N_2311);
nor U2368 (N_2368,N_2322,N_2347);
or U2369 (N_2369,N_2329,N_2301);
nor U2370 (N_2370,N_2333,N_2346);
xnor U2371 (N_2371,N_2340,N_2326);
nand U2372 (N_2372,N_2324,N_2320);
or U2373 (N_2373,N_2300,N_2315);
nor U2374 (N_2374,N_2302,N_2304);
nand U2375 (N_2375,N_2342,N_2332);
or U2376 (N_2376,N_2331,N_2339);
xor U2377 (N_2377,N_2327,N_2309);
or U2378 (N_2378,N_2310,N_2324);
and U2379 (N_2379,N_2347,N_2319);
and U2380 (N_2380,N_2316,N_2333);
or U2381 (N_2381,N_2301,N_2311);
nor U2382 (N_2382,N_2321,N_2307);
nor U2383 (N_2383,N_2314,N_2302);
nand U2384 (N_2384,N_2308,N_2305);
and U2385 (N_2385,N_2322,N_2339);
nor U2386 (N_2386,N_2349,N_2339);
nor U2387 (N_2387,N_2326,N_2344);
or U2388 (N_2388,N_2303,N_2318);
nand U2389 (N_2389,N_2304,N_2335);
nor U2390 (N_2390,N_2345,N_2317);
nand U2391 (N_2391,N_2347,N_2333);
nor U2392 (N_2392,N_2309,N_2315);
and U2393 (N_2393,N_2346,N_2319);
nor U2394 (N_2394,N_2315,N_2327);
and U2395 (N_2395,N_2325,N_2304);
or U2396 (N_2396,N_2312,N_2333);
and U2397 (N_2397,N_2307,N_2331);
or U2398 (N_2398,N_2328,N_2348);
nor U2399 (N_2399,N_2315,N_2337);
or U2400 (N_2400,N_2386,N_2387);
and U2401 (N_2401,N_2359,N_2395);
nor U2402 (N_2402,N_2376,N_2374);
nand U2403 (N_2403,N_2379,N_2383);
nand U2404 (N_2404,N_2396,N_2369);
nand U2405 (N_2405,N_2390,N_2394);
or U2406 (N_2406,N_2375,N_2377);
nor U2407 (N_2407,N_2372,N_2361);
nor U2408 (N_2408,N_2365,N_2371);
or U2409 (N_2409,N_2367,N_2360);
nor U2410 (N_2410,N_2356,N_2385);
nand U2411 (N_2411,N_2357,N_2373);
nor U2412 (N_2412,N_2363,N_2354);
xnor U2413 (N_2413,N_2382,N_2368);
nand U2414 (N_2414,N_2384,N_2391);
nor U2415 (N_2415,N_2397,N_2358);
nand U2416 (N_2416,N_2355,N_2378);
nor U2417 (N_2417,N_2389,N_2380);
and U2418 (N_2418,N_2351,N_2353);
nor U2419 (N_2419,N_2366,N_2350);
nor U2420 (N_2420,N_2352,N_2364);
xnor U2421 (N_2421,N_2370,N_2362);
nand U2422 (N_2422,N_2392,N_2388);
and U2423 (N_2423,N_2399,N_2393);
nand U2424 (N_2424,N_2381,N_2398);
and U2425 (N_2425,N_2365,N_2372);
nand U2426 (N_2426,N_2372,N_2378);
xor U2427 (N_2427,N_2390,N_2393);
and U2428 (N_2428,N_2365,N_2399);
and U2429 (N_2429,N_2381,N_2365);
nand U2430 (N_2430,N_2368,N_2383);
or U2431 (N_2431,N_2367,N_2353);
or U2432 (N_2432,N_2386,N_2366);
nor U2433 (N_2433,N_2353,N_2364);
or U2434 (N_2434,N_2358,N_2362);
nand U2435 (N_2435,N_2386,N_2399);
and U2436 (N_2436,N_2392,N_2369);
nand U2437 (N_2437,N_2388,N_2360);
and U2438 (N_2438,N_2385,N_2367);
or U2439 (N_2439,N_2375,N_2368);
and U2440 (N_2440,N_2353,N_2386);
xnor U2441 (N_2441,N_2368,N_2385);
or U2442 (N_2442,N_2390,N_2381);
xnor U2443 (N_2443,N_2371,N_2356);
nand U2444 (N_2444,N_2361,N_2363);
or U2445 (N_2445,N_2373,N_2375);
or U2446 (N_2446,N_2369,N_2361);
nor U2447 (N_2447,N_2354,N_2352);
and U2448 (N_2448,N_2350,N_2388);
xor U2449 (N_2449,N_2366,N_2384);
xor U2450 (N_2450,N_2416,N_2417);
nor U2451 (N_2451,N_2422,N_2434);
or U2452 (N_2452,N_2425,N_2447);
and U2453 (N_2453,N_2446,N_2409);
nor U2454 (N_2454,N_2420,N_2405);
nor U2455 (N_2455,N_2440,N_2407);
and U2456 (N_2456,N_2431,N_2439);
and U2457 (N_2457,N_2402,N_2412);
nand U2458 (N_2458,N_2408,N_2438);
and U2459 (N_2459,N_2411,N_2444);
and U2460 (N_2460,N_2421,N_2404);
or U2461 (N_2461,N_2449,N_2403);
and U2462 (N_2462,N_2448,N_2445);
nor U2463 (N_2463,N_2424,N_2415);
and U2464 (N_2464,N_2435,N_2428);
nand U2465 (N_2465,N_2419,N_2430);
or U2466 (N_2466,N_2441,N_2414);
nand U2467 (N_2467,N_2400,N_2401);
nand U2468 (N_2468,N_2426,N_2436);
or U2469 (N_2469,N_2442,N_2413);
and U2470 (N_2470,N_2429,N_2433);
nand U2471 (N_2471,N_2427,N_2443);
or U2472 (N_2472,N_2432,N_2418);
and U2473 (N_2473,N_2437,N_2410);
or U2474 (N_2474,N_2406,N_2423);
or U2475 (N_2475,N_2428,N_2410);
nor U2476 (N_2476,N_2423,N_2414);
or U2477 (N_2477,N_2426,N_2441);
or U2478 (N_2478,N_2428,N_2430);
xor U2479 (N_2479,N_2437,N_2430);
and U2480 (N_2480,N_2407,N_2444);
nand U2481 (N_2481,N_2437,N_2434);
nand U2482 (N_2482,N_2402,N_2407);
nor U2483 (N_2483,N_2402,N_2436);
nand U2484 (N_2484,N_2442,N_2421);
nand U2485 (N_2485,N_2426,N_2432);
and U2486 (N_2486,N_2431,N_2448);
and U2487 (N_2487,N_2406,N_2407);
or U2488 (N_2488,N_2437,N_2408);
nand U2489 (N_2489,N_2417,N_2418);
nor U2490 (N_2490,N_2408,N_2401);
nand U2491 (N_2491,N_2405,N_2417);
and U2492 (N_2492,N_2447,N_2418);
and U2493 (N_2493,N_2448,N_2442);
and U2494 (N_2494,N_2402,N_2415);
nand U2495 (N_2495,N_2424,N_2443);
or U2496 (N_2496,N_2444,N_2442);
nor U2497 (N_2497,N_2403,N_2441);
or U2498 (N_2498,N_2422,N_2412);
and U2499 (N_2499,N_2414,N_2419);
nor U2500 (N_2500,N_2453,N_2461);
or U2501 (N_2501,N_2480,N_2495);
or U2502 (N_2502,N_2488,N_2491);
nor U2503 (N_2503,N_2494,N_2459);
nand U2504 (N_2504,N_2477,N_2458);
or U2505 (N_2505,N_2470,N_2463);
nor U2506 (N_2506,N_2473,N_2469);
nor U2507 (N_2507,N_2468,N_2479);
or U2508 (N_2508,N_2451,N_2478);
nand U2509 (N_2509,N_2452,N_2466);
nand U2510 (N_2510,N_2457,N_2496);
or U2511 (N_2511,N_2456,N_2493);
or U2512 (N_2512,N_2465,N_2462);
and U2513 (N_2513,N_2497,N_2455);
nor U2514 (N_2514,N_2490,N_2471);
nor U2515 (N_2515,N_2485,N_2450);
xnor U2516 (N_2516,N_2481,N_2467);
and U2517 (N_2517,N_2492,N_2464);
and U2518 (N_2518,N_2487,N_2484);
xor U2519 (N_2519,N_2472,N_2489);
or U2520 (N_2520,N_2474,N_2460);
nor U2521 (N_2521,N_2475,N_2454);
or U2522 (N_2522,N_2482,N_2486);
nand U2523 (N_2523,N_2476,N_2499);
and U2524 (N_2524,N_2483,N_2498);
nor U2525 (N_2525,N_2483,N_2462);
or U2526 (N_2526,N_2466,N_2455);
nand U2527 (N_2527,N_2462,N_2452);
nand U2528 (N_2528,N_2474,N_2464);
nand U2529 (N_2529,N_2454,N_2455);
nor U2530 (N_2530,N_2490,N_2474);
and U2531 (N_2531,N_2461,N_2473);
nor U2532 (N_2532,N_2457,N_2498);
nor U2533 (N_2533,N_2481,N_2492);
xnor U2534 (N_2534,N_2494,N_2484);
or U2535 (N_2535,N_2480,N_2455);
and U2536 (N_2536,N_2493,N_2484);
xnor U2537 (N_2537,N_2453,N_2466);
and U2538 (N_2538,N_2479,N_2494);
nor U2539 (N_2539,N_2473,N_2480);
and U2540 (N_2540,N_2497,N_2461);
or U2541 (N_2541,N_2459,N_2485);
or U2542 (N_2542,N_2494,N_2488);
and U2543 (N_2543,N_2461,N_2464);
nor U2544 (N_2544,N_2455,N_2478);
nor U2545 (N_2545,N_2462,N_2475);
nor U2546 (N_2546,N_2486,N_2487);
and U2547 (N_2547,N_2490,N_2460);
nand U2548 (N_2548,N_2480,N_2486);
nor U2549 (N_2549,N_2464,N_2456);
nor U2550 (N_2550,N_2548,N_2543);
nand U2551 (N_2551,N_2541,N_2542);
xor U2552 (N_2552,N_2512,N_2518);
nor U2553 (N_2553,N_2519,N_2501);
nand U2554 (N_2554,N_2546,N_2523);
xnor U2555 (N_2555,N_2530,N_2517);
nor U2556 (N_2556,N_2503,N_2540);
or U2557 (N_2557,N_2527,N_2524);
or U2558 (N_2558,N_2505,N_2545);
xor U2559 (N_2559,N_2521,N_2538);
and U2560 (N_2560,N_2502,N_2513);
nor U2561 (N_2561,N_2511,N_2507);
or U2562 (N_2562,N_2510,N_2544);
nand U2563 (N_2563,N_2514,N_2547);
nor U2564 (N_2564,N_2522,N_2534);
nand U2565 (N_2565,N_2539,N_2525);
nand U2566 (N_2566,N_2549,N_2531);
or U2567 (N_2567,N_2515,N_2526);
nor U2568 (N_2568,N_2506,N_2532);
and U2569 (N_2569,N_2508,N_2504);
or U2570 (N_2570,N_2500,N_2535);
nor U2571 (N_2571,N_2533,N_2509);
nor U2572 (N_2572,N_2516,N_2528);
or U2573 (N_2573,N_2520,N_2536);
and U2574 (N_2574,N_2537,N_2529);
xnor U2575 (N_2575,N_2534,N_2533);
and U2576 (N_2576,N_2530,N_2532);
xor U2577 (N_2577,N_2502,N_2530);
nand U2578 (N_2578,N_2511,N_2503);
nor U2579 (N_2579,N_2525,N_2534);
nor U2580 (N_2580,N_2528,N_2524);
xnor U2581 (N_2581,N_2534,N_2531);
nand U2582 (N_2582,N_2528,N_2548);
nand U2583 (N_2583,N_2521,N_2536);
nand U2584 (N_2584,N_2523,N_2511);
nand U2585 (N_2585,N_2541,N_2544);
nor U2586 (N_2586,N_2537,N_2508);
nor U2587 (N_2587,N_2538,N_2503);
nand U2588 (N_2588,N_2502,N_2537);
nand U2589 (N_2589,N_2510,N_2543);
or U2590 (N_2590,N_2504,N_2513);
nand U2591 (N_2591,N_2547,N_2515);
xnor U2592 (N_2592,N_2507,N_2513);
and U2593 (N_2593,N_2515,N_2502);
nand U2594 (N_2594,N_2526,N_2506);
and U2595 (N_2595,N_2538,N_2513);
nand U2596 (N_2596,N_2512,N_2506);
or U2597 (N_2597,N_2516,N_2529);
or U2598 (N_2598,N_2507,N_2521);
nor U2599 (N_2599,N_2543,N_2545);
or U2600 (N_2600,N_2580,N_2566);
nor U2601 (N_2601,N_2598,N_2599);
and U2602 (N_2602,N_2565,N_2584);
nand U2603 (N_2603,N_2556,N_2555);
or U2604 (N_2604,N_2559,N_2593);
and U2605 (N_2605,N_2581,N_2564);
and U2606 (N_2606,N_2554,N_2563);
nand U2607 (N_2607,N_2560,N_2577);
nor U2608 (N_2608,N_2586,N_2569);
and U2609 (N_2609,N_2590,N_2585);
nor U2610 (N_2610,N_2592,N_2595);
or U2611 (N_2611,N_2596,N_2550);
nand U2612 (N_2612,N_2588,N_2572);
nand U2613 (N_2613,N_2576,N_2573);
or U2614 (N_2614,N_2591,N_2552);
and U2615 (N_2615,N_2567,N_2582);
or U2616 (N_2616,N_2551,N_2575);
nand U2617 (N_2617,N_2597,N_2571);
nand U2618 (N_2618,N_2558,N_2562);
nor U2619 (N_2619,N_2561,N_2574);
nor U2620 (N_2620,N_2568,N_2579);
and U2621 (N_2621,N_2557,N_2570);
and U2622 (N_2622,N_2594,N_2578);
and U2623 (N_2623,N_2589,N_2583);
nor U2624 (N_2624,N_2587,N_2553);
xnor U2625 (N_2625,N_2590,N_2594);
and U2626 (N_2626,N_2577,N_2578);
nor U2627 (N_2627,N_2590,N_2564);
nand U2628 (N_2628,N_2566,N_2592);
and U2629 (N_2629,N_2593,N_2583);
and U2630 (N_2630,N_2587,N_2583);
xor U2631 (N_2631,N_2591,N_2573);
nor U2632 (N_2632,N_2550,N_2599);
or U2633 (N_2633,N_2571,N_2593);
nor U2634 (N_2634,N_2588,N_2574);
nor U2635 (N_2635,N_2563,N_2581);
nor U2636 (N_2636,N_2558,N_2596);
and U2637 (N_2637,N_2571,N_2555);
or U2638 (N_2638,N_2587,N_2595);
or U2639 (N_2639,N_2551,N_2562);
nand U2640 (N_2640,N_2591,N_2582);
and U2641 (N_2641,N_2563,N_2550);
xor U2642 (N_2642,N_2569,N_2568);
xnor U2643 (N_2643,N_2583,N_2553);
nor U2644 (N_2644,N_2597,N_2577);
xor U2645 (N_2645,N_2557,N_2553);
nand U2646 (N_2646,N_2558,N_2582);
or U2647 (N_2647,N_2566,N_2567);
nor U2648 (N_2648,N_2583,N_2576);
nand U2649 (N_2649,N_2569,N_2577);
and U2650 (N_2650,N_2643,N_2638);
or U2651 (N_2651,N_2607,N_2640);
or U2652 (N_2652,N_2644,N_2633);
nand U2653 (N_2653,N_2642,N_2616);
nor U2654 (N_2654,N_2641,N_2617);
or U2655 (N_2655,N_2632,N_2615);
nand U2656 (N_2656,N_2623,N_2624);
nand U2657 (N_2657,N_2602,N_2637);
or U2658 (N_2658,N_2627,N_2619);
nand U2659 (N_2659,N_2649,N_2625);
nand U2660 (N_2660,N_2647,N_2612);
or U2661 (N_2661,N_2608,N_2622);
nand U2662 (N_2662,N_2645,N_2628);
or U2663 (N_2663,N_2603,N_2606);
and U2664 (N_2664,N_2600,N_2630);
or U2665 (N_2665,N_2639,N_2636);
nand U2666 (N_2666,N_2618,N_2631);
xor U2667 (N_2667,N_2621,N_2610);
nor U2668 (N_2668,N_2634,N_2635);
nand U2669 (N_2669,N_2629,N_2611);
nand U2670 (N_2670,N_2626,N_2614);
nand U2671 (N_2671,N_2604,N_2613);
nor U2672 (N_2672,N_2605,N_2620);
nand U2673 (N_2673,N_2648,N_2609);
or U2674 (N_2674,N_2601,N_2646);
and U2675 (N_2675,N_2614,N_2616);
and U2676 (N_2676,N_2606,N_2639);
or U2677 (N_2677,N_2610,N_2640);
and U2678 (N_2678,N_2646,N_2625);
xor U2679 (N_2679,N_2608,N_2647);
or U2680 (N_2680,N_2602,N_2648);
xnor U2681 (N_2681,N_2611,N_2614);
nand U2682 (N_2682,N_2610,N_2603);
or U2683 (N_2683,N_2626,N_2605);
and U2684 (N_2684,N_2648,N_2616);
and U2685 (N_2685,N_2606,N_2628);
or U2686 (N_2686,N_2619,N_2628);
nor U2687 (N_2687,N_2602,N_2631);
nand U2688 (N_2688,N_2630,N_2627);
nor U2689 (N_2689,N_2627,N_2607);
xor U2690 (N_2690,N_2617,N_2628);
or U2691 (N_2691,N_2613,N_2627);
nand U2692 (N_2692,N_2608,N_2636);
nor U2693 (N_2693,N_2628,N_2621);
nor U2694 (N_2694,N_2646,N_2649);
and U2695 (N_2695,N_2630,N_2602);
nand U2696 (N_2696,N_2640,N_2611);
and U2697 (N_2697,N_2642,N_2607);
and U2698 (N_2698,N_2637,N_2617);
nand U2699 (N_2699,N_2606,N_2636);
nor U2700 (N_2700,N_2664,N_2699);
and U2701 (N_2701,N_2665,N_2674);
nand U2702 (N_2702,N_2690,N_2669);
nor U2703 (N_2703,N_2650,N_2670);
nor U2704 (N_2704,N_2675,N_2676);
nor U2705 (N_2705,N_2677,N_2684);
and U2706 (N_2706,N_2652,N_2658);
nand U2707 (N_2707,N_2698,N_2679);
or U2708 (N_2708,N_2667,N_2693);
and U2709 (N_2709,N_2668,N_2678);
xor U2710 (N_2710,N_2687,N_2657);
xnor U2711 (N_2711,N_2660,N_2681);
or U2712 (N_2712,N_2683,N_2691);
nor U2713 (N_2713,N_2672,N_2685);
nand U2714 (N_2714,N_2651,N_2662);
xnor U2715 (N_2715,N_2682,N_2659);
nand U2716 (N_2716,N_2695,N_2686);
and U2717 (N_2717,N_2688,N_2697);
or U2718 (N_2718,N_2671,N_2656);
and U2719 (N_2719,N_2689,N_2654);
nor U2720 (N_2720,N_2673,N_2696);
xor U2721 (N_2721,N_2653,N_2661);
nand U2722 (N_2722,N_2692,N_2680);
nand U2723 (N_2723,N_2663,N_2655);
nand U2724 (N_2724,N_2666,N_2694);
or U2725 (N_2725,N_2674,N_2650);
nor U2726 (N_2726,N_2685,N_2683);
or U2727 (N_2727,N_2686,N_2674);
and U2728 (N_2728,N_2680,N_2677);
xnor U2729 (N_2729,N_2682,N_2691);
nand U2730 (N_2730,N_2652,N_2671);
nand U2731 (N_2731,N_2680,N_2655);
or U2732 (N_2732,N_2666,N_2682);
nand U2733 (N_2733,N_2658,N_2667);
and U2734 (N_2734,N_2691,N_2678);
or U2735 (N_2735,N_2654,N_2683);
or U2736 (N_2736,N_2653,N_2694);
or U2737 (N_2737,N_2655,N_2682);
nand U2738 (N_2738,N_2659,N_2657);
nand U2739 (N_2739,N_2691,N_2654);
xor U2740 (N_2740,N_2663,N_2661);
or U2741 (N_2741,N_2671,N_2683);
or U2742 (N_2742,N_2678,N_2685);
nor U2743 (N_2743,N_2651,N_2650);
xor U2744 (N_2744,N_2698,N_2665);
or U2745 (N_2745,N_2684,N_2693);
xnor U2746 (N_2746,N_2686,N_2676);
or U2747 (N_2747,N_2698,N_2696);
and U2748 (N_2748,N_2686,N_2681);
and U2749 (N_2749,N_2653,N_2683);
and U2750 (N_2750,N_2740,N_2731);
nand U2751 (N_2751,N_2747,N_2713);
and U2752 (N_2752,N_2708,N_2706);
and U2753 (N_2753,N_2729,N_2725);
and U2754 (N_2754,N_2738,N_2724);
xnor U2755 (N_2755,N_2728,N_2744);
and U2756 (N_2756,N_2727,N_2720);
xor U2757 (N_2757,N_2736,N_2704);
or U2758 (N_2758,N_2748,N_2719);
and U2759 (N_2759,N_2735,N_2703);
nand U2760 (N_2760,N_2712,N_2739);
and U2761 (N_2761,N_2723,N_2726);
or U2762 (N_2762,N_2710,N_2717);
xor U2763 (N_2763,N_2714,N_2742);
nor U2764 (N_2764,N_2746,N_2741);
or U2765 (N_2765,N_2711,N_2749);
nand U2766 (N_2766,N_2730,N_2722);
or U2767 (N_2767,N_2732,N_2734);
and U2768 (N_2768,N_2721,N_2705);
nor U2769 (N_2769,N_2737,N_2718);
xnor U2770 (N_2770,N_2745,N_2701);
and U2771 (N_2771,N_2733,N_2709);
xnor U2772 (N_2772,N_2700,N_2743);
or U2773 (N_2773,N_2707,N_2715);
nor U2774 (N_2774,N_2716,N_2702);
or U2775 (N_2775,N_2708,N_2712);
nor U2776 (N_2776,N_2701,N_2715);
nor U2777 (N_2777,N_2712,N_2722);
xor U2778 (N_2778,N_2729,N_2722);
xnor U2779 (N_2779,N_2742,N_2728);
nor U2780 (N_2780,N_2715,N_2726);
xnor U2781 (N_2781,N_2704,N_2707);
xor U2782 (N_2782,N_2716,N_2709);
or U2783 (N_2783,N_2708,N_2711);
nand U2784 (N_2784,N_2712,N_2726);
or U2785 (N_2785,N_2714,N_2725);
nand U2786 (N_2786,N_2729,N_2700);
nor U2787 (N_2787,N_2715,N_2735);
nor U2788 (N_2788,N_2741,N_2723);
or U2789 (N_2789,N_2710,N_2740);
nand U2790 (N_2790,N_2708,N_2718);
and U2791 (N_2791,N_2707,N_2744);
nor U2792 (N_2792,N_2748,N_2726);
and U2793 (N_2793,N_2739,N_2743);
and U2794 (N_2794,N_2732,N_2748);
and U2795 (N_2795,N_2739,N_2748);
and U2796 (N_2796,N_2703,N_2724);
xor U2797 (N_2797,N_2717,N_2703);
or U2798 (N_2798,N_2726,N_2730);
and U2799 (N_2799,N_2705,N_2719);
or U2800 (N_2800,N_2784,N_2780);
and U2801 (N_2801,N_2765,N_2753);
nand U2802 (N_2802,N_2792,N_2754);
or U2803 (N_2803,N_2761,N_2799);
nand U2804 (N_2804,N_2797,N_2786);
nor U2805 (N_2805,N_2785,N_2766);
nor U2806 (N_2806,N_2758,N_2751);
nand U2807 (N_2807,N_2788,N_2782);
or U2808 (N_2808,N_2759,N_2762);
xor U2809 (N_2809,N_2770,N_2763);
nand U2810 (N_2810,N_2794,N_2772);
and U2811 (N_2811,N_2771,N_2756);
or U2812 (N_2812,N_2760,N_2790);
or U2813 (N_2813,N_2779,N_2798);
nand U2814 (N_2814,N_2781,N_2776);
and U2815 (N_2815,N_2752,N_2783);
or U2816 (N_2816,N_2778,N_2769);
nand U2817 (N_2817,N_2757,N_2791);
nor U2818 (N_2818,N_2767,N_2787);
and U2819 (N_2819,N_2768,N_2773);
nor U2820 (N_2820,N_2796,N_2777);
nor U2821 (N_2821,N_2775,N_2793);
nand U2822 (N_2822,N_2755,N_2795);
or U2823 (N_2823,N_2750,N_2764);
nor U2824 (N_2824,N_2774,N_2789);
or U2825 (N_2825,N_2761,N_2773);
and U2826 (N_2826,N_2766,N_2787);
nor U2827 (N_2827,N_2792,N_2767);
xnor U2828 (N_2828,N_2794,N_2758);
or U2829 (N_2829,N_2775,N_2766);
nand U2830 (N_2830,N_2779,N_2751);
nor U2831 (N_2831,N_2798,N_2781);
or U2832 (N_2832,N_2785,N_2768);
and U2833 (N_2833,N_2764,N_2780);
xnor U2834 (N_2834,N_2782,N_2799);
or U2835 (N_2835,N_2795,N_2757);
nand U2836 (N_2836,N_2755,N_2789);
and U2837 (N_2837,N_2789,N_2752);
and U2838 (N_2838,N_2758,N_2783);
or U2839 (N_2839,N_2785,N_2792);
nand U2840 (N_2840,N_2792,N_2797);
nand U2841 (N_2841,N_2765,N_2764);
nor U2842 (N_2842,N_2768,N_2775);
nor U2843 (N_2843,N_2795,N_2780);
nor U2844 (N_2844,N_2756,N_2778);
and U2845 (N_2845,N_2751,N_2754);
or U2846 (N_2846,N_2775,N_2781);
and U2847 (N_2847,N_2765,N_2792);
or U2848 (N_2848,N_2798,N_2750);
xnor U2849 (N_2849,N_2776,N_2769);
xnor U2850 (N_2850,N_2831,N_2809);
nand U2851 (N_2851,N_2846,N_2844);
nor U2852 (N_2852,N_2818,N_2800);
or U2853 (N_2853,N_2842,N_2807);
or U2854 (N_2854,N_2813,N_2811);
and U2855 (N_2855,N_2812,N_2821);
nand U2856 (N_2856,N_2833,N_2822);
nor U2857 (N_2857,N_2802,N_2806);
xor U2858 (N_2858,N_2835,N_2803);
and U2859 (N_2859,N_2836,N_2823);
nand U2860 (N_2860,N_2843,N_2815);
or U2861 (N_2861,N_2847,N_2801);
and U2862 (N_2862,N_2808,N_2841);
and U2863 (N_2863,N_2814,N_2832);
or U2864 (N_2864,N_2838,N_2819);
nand U2865 (N_2865,N_2827,N_2834);
and U2866 (N_2866,N_2826,N_2805);
and U2867 (N_2867,N_2830,N_2837);
nor U2868 (N_2868,N_2828,N_2804);
nand U2869 (N_2869,N_2848,N_2840);
or U2870 (N_2870,N_2820,N_2839);
nand U2871 (N_2871,N_2810,N_2845);
nand U2872 (N_2872,N_2829,N_2824);
nand U2873 (N_2873,N_2825,N_2817);
nand U2874 (N_2874,N_2849,N_2816);
nor U2875 (N_2875,N_2845,N_2816);
and U2876 (N_2876,N_2829,N_2839);
or U2877 (N_2877,N_2806,N_2834);
or U2878 (N_2878,N_2842,N_2839);
and U2879 (N_2879,N_2808,N_2829);
xnor U2880 (N_2880,N_2803,N_2833);
and U2881 (N_2881,N_2837,N_2812);
nand U2882 (N_2882,N_2815,N_2813);
nand U2883 (N_2883,N_2828,N_2831);
nand U2884 (N_2884,N_2805,N_2848);
nand U2885 (N_2885,N_2848,N_2837);
nand U2886 (N_2886,N_2823,N_2818);
nor U2887 (N_2887,N_2804,N_2849);
xor U2888 (N_2888,N_2846,N_2845);
nor U2889 (N_2889,N_2836,N_2804);
nor U2890 (N_2890,N_2839,N_2806);
nand U2891 (N_2891,N_2809,N_2806);
nor U2892 (N_2892,N_2827,N_2814);
nand U2893 (N_2893,N_2814,N_2818);
xnor U2894 (N_2894,N_2827,N_2803);
nand U2895 (N_2895,N_2832,N_2845);
nor U2896 (N_2896,N_2825,N_2810);
nand U2897 (N_2897,N_2812,N_2801);
nor U2898 (N_2898,N_2844,N_2810);
nor U2899 (N_2899,N_2814,N_2804);
nor U2900 (N_2900,N_2880,N_2892);
and U2901 (N_2901,N_2866,N_2851);
or U2902 (N_2902,N_2858,N_2864);
or U2903 (N_2903,N_2897,N_2859);
or U2904 (N_2904,N_2889,N_2890);
xor U2905 (N_2905,N_2876,N_2856);
and U2906 (N_2906,N_2853,N_2857);
or U2907 (N_2907,N_2881,N_2863);
nand U2908 (N_2908,N_2868,N_2875);
nand U2909 (N_2909,N_2852,N_2877);
xnor U2910 (N_2910,N_2898,N_2861);
and U2911 (N_2911,N_2893,N_2899);
nor U2912 (N_2912,N_2882,N_2867);
nand U2913 (N_2913,N_2872,N_2888);
nor U2914 (N_2914,N_2879,N_2887);
and U2915 (N_2915,N_2865,N_2870);
or U2916 (N_2916,N_2891,N_2855);
and U2917 (N_2917,N_2854,N_2894);
or U2918 (N_2918,N_2873,N_2878);
and U2919 (N_2919,N_2895,N_2871);
nand U2920 (N_2920,N_2896,N_2883);
nor U2921 (N_2921,N_2874,N_2886);
and U2922 (N_2922,N_2850,N_2885);
nand U2923 (N_2923,N_2862,N_2884);
and U2924 (N_2924,N_2869,N_2860);
or U2925 (N_2925,N_2889,N_2857);
or U2926 (N_2926,N_2867,N_2876);
nor U2927 (N_2927,N_2894,N_2852);
and U2928 (N_2928,N_2868,N_2850);
xnor U2929 (N_2929,N_2858,N_2852);
or U2930 (N_2930,N_2854,N_2879);
nor U2931 (N_2931,N_2884,N_2865);
and U2932 (N_2932,N_2853,N_2888);
nand U2933 (N_2933,N_2860,N_2884);
nand U2934 (N_2934,N_2886,N_2854);
xor U2935 (N_2935,N_2863,N_2871);
and U2936 (N_2936,N_2868,N_2897);
or U2937 (N_2937,N_2890,N_2858);
nand U2938 (N_2938,N_2850,N_2893);
and U2939 (N_2939,N_2860,N_2883);
nor U2940 (N_2940,N_2859,N_2871);
nand U2941 (N_2941,N_2867,N_2862);
and U2942 (N_2942,N_2856,N_2883);
nor U2943 (N_2943,N_2854,N_2887);
xor U2944 (N_2944,N_2862,N_2852);
nand U2945 (N_2945,N_2887,N_2890);
nand U2946 (N_2946,N_2864,N_2869);
and U2947 (N_2947,N_2882,N_2861);
nand U2948 (N_2948,N_2862,N_2854);
nor U2949 (N_2949,N_2888,N_2884);
and U2950 (N_2950,N_2908,N_2936);
nand U2951 (N_2951,N_2907,N_2929);
and U2952 (N_2952,N_2928,N_2935);
or U2953 (N_2953,N_2941,N_2911);
or U2954 (N_2954,N_2934,N_2932);
and U2955 (N_2955,N_2901,N_2900);
nor U2956 (N_2956,N_2942,N_2910);
and U2957 (N_2957,N_2903,N_2919);
or U2958 (N_2958,N_2902,N_2922);
or U2959 (N_2959,N_2906,N_2905);
or U2960 (N_2960,N_2915,N_2913);
nor U2961 (N_2961,N_2943,N_2930);
or U2962 (N_2962,N_2904,N_2916);
nand U2963 (N_2963,N_2945,N_2927);
nor U2964 (N_2964,N_2946,N_2920);
or U2965 (N_2965,N_2909,N_2925);
nor U2966 (N_2966,N_2938,N_2924);
nand U2967 (N_2967,N_2914,N_2937);
or U2968 (N_2968,N_2921,N_2940);
nor U2969 (N_2969,N_2917,N_2933);
nand U2970 (N_2970,N_2944,N_2931);
nand U2971 (N_2971,N_2923,N_2926);
nand U2972 (N_2972,N_2918,N_2947);
and U2973 (N_2973,N_2948,N_2939);
and U2974 (N_2974,N_2912,N_2949);
and U2975 (N_2975,N_2913,N_2918);
nor U2976 (N_2976,N_2943,N_2908);
and U2977 (N_2977,N_2925,N_2901);
nor U2978 (N_2978,N_2921,N_2919);
nand U2979 (N_2979,N_2914,N_2902);
xor U2980 (N_2980,N_2915,N_2921);
xnor U2981 (N_2981,N_2927,N_2910);
and U2982 (N_2982,N_2929,N_2927);
nand U2983 (N_2983,N_2918,N_2927);
nand U2984 (N_2984,N_2942,N_2933);
nor U2985 (N_2985,N_2938,N_2915);
and U2986 (N_2986,N_2908,N_2922);
nand U2987 (N_2987,N_2945,N_2924);
or U2988 (N_2988,N_2926,N_2920);
nand U2989 (N_2989,N_2939,N_2907);
xnor U2990 (N_2990,N_2902,N_2948);
nand U2991 (N_2991,N_2945,N_2933);
nand U2992 (N_2992,N_2911,N_2940);
or U2993 (N_2993,N_2941,N_2923);
nand U2994 (N_2994,N_2920,N_2925);
and U2995 (N_2995,N_2900,N_2922);
nand U2996 (N_2996,N_2940,N_2900);
and U2997 (N_2997,N_2947,N_2926);
and U2998 (N_2998,N_2938,N_2919);
nor U2999 (N_2999,N_2946,N_2942);
and UO_0 (O_0,N_2971,N_2978);
nor UO_1 (O_1,N_2973,N_2981);
nand UO_2 (O_2,N_2965,N_2985);
nand UO_3 (O_3,N_2970,N_2984);
xnor UO_4 (O_4,N_2986,N_2991);
nor UO_5 (O_5,N_2962,N_2963);
and UO_6 (O_6,N_2972,N_2976);
or UO_7 (O_7,N_2952,N_2992);
nand UO_8 (O_8,N_2964,N_2989);
nand UO_9 (O_9,N_2960,N_2956);
nand UO_10 (O_10,N_2994,N_2951);
xor UO_11 (O_11,N_2959,N_2950);
and UO_12 (O_12,N_2974,N_2997);
nor UO_13 (O_13,N_2993,N_2977);
nor UO_14 (O_14,N_2987,N_2957);
nand UO_15 (O_15,N_2969,N_2996);
nand UO_16 (O_16,N_2955,N_2966);
or UO_17 (O_17,N_2954,N_2953);
nor UO_18 (O_18,N_2988,N_2990);
xnor UO_19 (O_19,N_2980,N_2975);
nor UO_20 (O_20,N_2983,N_2958);
or UO_21 (O_21,N_2998,N_2968);
and UO_22 (O_22,N_2999,N_2967);
or UO_23 (O_23,N_2995,N_2982);
nand UO_24 (O_24,N_2979,N_2961);
nand UO_25 (O_25,N_2997,N_2971);
and UO_26 (O_26,N_2950,N_2974);
nand UO_27 (O_27,N_2960,N_2953);
nand UO_28 (O_28,N_2970,N_2981);
nand UO_29 (O_29,N_2981,N_2956);
and UO_30 (O_30,N_2984,N_2989);
and UO_31 (O_31,N_2983,N_2981);
or UO_32 (O_32,N_2989,N_2956);
or UO_33 (O_33,N_2951,N_2991);
xnor UO_34 (O_34,N_2982,N_2986);
or UO_35 (O_35,N_2965,N_2974);
or UO_36 (O_36,N_2973,N_2974);
xor UO_37 (O_37,N_2984,N_2977);
nor UO_38 (O_38,N_2997,N_2985);
nor UO_39 (O_39,N_2990,N_2959);
nor UO_40 (O_40,N_2969,N_2959);
nor UO_41 (O_41,N_2967,N_2982);
and UO_42 (O_42,N_2979,N_2973);
and UO_43 (O_43,N_2984,N_2991);
nor UO_44 (O_44,N_2997,N_2989);
nand UO_45 (O_45,N_2979,N_2994);
and UO_46 (O_46,N_2975,N_2956);
or UO_47 (O_47,N_2971,N_2963);
nand UO_48 (O_48,N_2987,N_2982);
and UO_49 (O_49,N_2953,N_2992);
nand UO_50 (O_50,N_2978,N_2988);
xor UO_51 (O_51,N_2963,N_2983);
and UO_52 (O_52,N_2967,N_2969);
or UO_53 (O_53,N_2957,N_2996);
and UO_54 (O_54,N_2958,N_2967);
xnor UO_55 (O_55,N_2965,N_2989);
nor UO_56 (O_56,N_2982,N_2961);
nor UO_57 (O_57,N_2991,N_2955);
or UO_58 (O_58,N_2961,N_2966);
and UO_59 (O_59,N_2981,N_2991);
xnor UO_60 (O_60,N_2999,N_2995);
or UO_61 (O_61,N_2965,N_2992);
nand UO_62 (O_62,N_2976,N_2955);
and UO_63 (O_63,N_2954,N_2989);
nand UO_64 (O_64,N_2986,N_2958);
nand UO_65 (O_65,N_2968,N_2993);
xor UO_66 (O_66,N_2985,N_2996);
and UO_67 (O_67,N_2983,N_2961);
xor UO_68 (O_68,N_2986,N_2992);
and UO_69 (O_69,N_2992,N_2972);
and UO_70 (O_70,N_2979,N_2964);
nor UO_71 (O_71,N_2951,N_2984);
nand UO_72 (O_72,N_2967,N_2979);
nor UO_73 (O_73,N_2996,N_2975);
and UO_74 (O_74,N_2975,N_2955);
or UO_75 (O_75,N_2979,N_2960);
and UO_76 (O_76,N_2971,N_2973);
and UO_77 (O_77,N_2987,N_2964);
or UO_78 (O_78,N_2957,N_2965);
nand UO_79 (O_79,N_2987,N_2990);
nand UO_80 (O_80,N_2996,N_2987);
and UO_81 (O_81,N_2967,N_2960);
nand UO_82 (O_82,N_2980,N_2955);
and UO_83 (O_83,N_2979,N_2968);
or UO_84 (O_84,N_2950,N_2989);
nor UO_85 (O_85,N_2970,N_2977);
xnor UO_86 (O_86,N_2957,N_2974);
and UO_87 (O_87,N_2952,N_2999);
xnor UO_88 (O_88,N_2956,N_2994);
nor UO_89 (O_89,N_2976,N_2966);
nor UO_90 (O_90,N_2990,N_2992);
nor UO_91 (O_91,N_2994,N_2974);
nor UO_92 (O_92,N_2987,N_2983);
nor UO_93 (O_93,N_2961,N_2992);
xor UO_94 (O_94,N_2956,N_2970);
or UO_95 (O_95,N_2950,N_2994);
nand UO_96 (O_96,N_2986,N_2988);
or UO_97 (O_97,N_2987,N_2963);
or UO_98 (O_98,N_2956,N_2991);
and UO_99 (O_99,N_2977,N_2959);
or UO_100 (O_100,N_2955,N_2974);
nand UO_101 (O_101,N_2964,N_2994);
nor UO_102 (O_102,N_2955,N_2954);
nor UO_103 (O_103,N_2965,N_2980);
nor UO_104 (O_104,N_2990,N_2964);
nor UO_105 (O_105,N_2982,N_2983);
and UO_106 (O_106,N_2978,N_2975);
nand UO_107 (O_107,N_2950,N_2951);
xnor UO_108 (O_108,N_2992,N_2950);
xnor UO_109 (O_109,N_2975,N_2986);
and UO_110 (O_110,N_2974,N_2979);
or UO_111 (O_111,N_2950,N_2985);
xnor UO_112 (O_112,N_2961,N_2998);
or UO_113 (O_113,N_2971,N_2962);
nor UO_114 (O_114,N_2968,N_2955);
and UO_115 (O_115,N_2956,N_2963);
or UO_116 (O_116,N_2973,N_2950);
nand UO_117 (O_117,N_2979,N_2996);
nor UO_118 (O_118,N_2988,N_2981);
nand UO_119 (O_119,N_2992,N_2966);
nor UO_120 (O_120,N_2983,N_2976);
or UO_121 (O_121,N_2966,N_2993);
xor UO_122 (O_122,N_2966,N_2999);
xor UO_123 (O_123,N_2963,N_2992);
and UO_124 (O_124,N_2976,N_2963);
nand UO_125 (O_125,N_2953,N_2983);
and UO_126 (O_126,N_2994,N_2980);
xor UO_127 (O_127,N_2956,N_2964);
xnor UO_128 (O_128,N_2986,N_2970);
nor UO_129 (O_129,N_2950,N_2991);
or UO_130 (O_130,N_2953,N_2973);
nor UO_131 (O_131,N_2981,N_2990);
and UO_132 (O_132,N_2957,N_2954);
xor UO_133 (O_133,N_2982,N_2985);
or UO_134 (O_134,N_2996,N_2991);
nor UO_135 (O_135,N_2979,N_2998);
and UO_136 (O_136,N_2999,N_2996);
and UO_137 (O_137,N_2995,N_2997);
or UO_138 (O_138,N_2983,N_2997);
nand UO_139 (O_139,N_2998,N_2985);
nand UO_140 (O_140,N_2958,N_2973);
nor UO_141 (O_141,N_2956,N_2995);
or UO_142 (O_142,N_2993,N_2954);
nand UO_143 (O_143,N_2968,N_2958);
nand UO_144 (O_144,N_2959,N_2974);
or UO_145 (O_145,N_2986,N_2967);
and UO_146 (O_146,N_2973,N_2964);
or UO_147 (O_147,N_2952,N_2961);
nand UO_148 (O_148,N_2981,N_2977);
nand UO_149 (O_149,N_2953,N_2955);
and UO_150 (O_150,N_2985,N_2971);
nand UO_151 (O_151,N_2962,N_2985);
xnor UO_152 (O_152,N_2974,N_2956);
or UO_153 (O_153,N_2955,N_2973);
or UO_154 (O_154,N_2957,N_2971);
or UO_155 (O_155,N_2996,N_2997);
nor UO_156 (O_156,N_2959,N_2963);
nand UO_157 (O_157,N_2964,N_2961);
and UO_158 (O_158,N_2968,N_2974);
and UO_159 (O_159,N_2996,N_2950);
or UO_160 (O_160,N_2959,N_2965);
xnor UO_161 (O_161,N_2962,N_2967);
and UO_162 (O_162,N_2982,N_2955);
or UO_163 (O_163,N_2958,N_2953);
nor UO_164 (O_164,N_2973,N_2993);
nor UO_165 (O_165,N_2961,N_2969);
and UO_166 (O_166,N_2967,N_2970);
and UO_167 (O_167,N_2966,N_2951);
nand UO_168 (O_168,N_2988,N_2992);
xor UO_169 (O_169,N_2950,N_2966);
or UO_170 (O_170,N_2997,N_2967);
nor UO_171 (O_171,N_2985,N_2979);
and UO_172 (O_172,N_2950,N_2995);
or UO_173 (O_173,N_2952,N_2970);
nand UO_174 (O_174,N_2958,N_2981);
xor UO_175 (O_175,N_2993,N_2970);
and UO_176 (O_176,N_2970,N_2966);
and UO_177 (O_177,N_2965,N_2986);
and UO_178 (O_178,N_2987,N_2993);
or UO_179 (O_179,N_2998,N_2969);
nand UO_180 (O_180,N_2983,N_2965);
nor UO_181 (O_181,N_2979,N_2981);
nor UO_182 (O_182,N_2983,N_2975);
and UO_183 (O_183,N_2999,N_2975);
nand UO_184 (O_184,N_2991,N_2982);
and UO_185 (O_185,N_2967,N_2952);
nand UO_186 (O_186,N_2960,N_2993);
nor UO_187 (O_187,N_2988,N_2979);
nor UO_188 (O_188,N_2958,N_2997);
xnor UO_189 (O_189,N_2954,N_2972);
and UO_190 (O_190,N_2992,N_2977);
nor UO_191 (O_191,N_2967,N_2973);
nor UO_192 (O_192,N_2994,N_2999);
nand UO_193 (O_193,N_2986,N_2997);
xnor UO_194 (O_194,N_2972,N_2981);
nand UO_195 (O_195,N_2972,N_2973);
nor UO_196 (O_196,N_2996,N_2968);
and UO_197 (O_197,N_2980,N_2990);
nand UO_198 (O_198,N_2961,N_2958);
and UO_199 (O_199,N_2997,N_2959);
nor UO_200 (O_200,N_2966,N_2978);
and UO_201 (O_201,N_2987,N_2968);
xor UO_202 (O_202,N_2959,N_2973);
and UO_203 (O_203,N_2987,N_2978);
nor UO_204 (O_204,N_2953,N_2961);
or UO_205 (O_205,N_2953,N_2957);
and UO_206 (O_206,N_2984,N_2997);
or UO_207 (O_207,N_2964,N_2968);
nand UO_208 (O_208,N_2990,N_2952);
or UO_209 (O_209,N_2961,N_2993);
or UO_210 (O_210,N_2984,N_2952);
and UO_211 (O_211,N_2966,N_2994);
nand UO_212 (O_212,N_2951,N_2996);
and UO_213 (O_213,N_2956,N_2997);
nand UO_214 (O_214,N_2969,N_2963);
nand UO_215 (O_215,N_2957,N_2966);
or UO_216 (O_216,N_2958,N_2978);
and UO_217 (O_217,N_2979,N_2952);
nand UO_218 (O_218,N_2988,N_2957);
or UO_219 (O_219,N_2965,N_2982);
nand UO_220 (O_220,N_2957,N_2983);
nand UO_221 (O_221,N_2986,N_2974);
nand UO_222 (O_222,N_2969,N_2964);
or UO_223 (O_223,N_2972,N_2971);
nand UO_224 (O_224,N_2966,N_2988);
and UO_225 (O_225,N_2971,N_2952);
xnor UO_226 (O_226,N_2951,N_2999);
nor UO_227 (O_227,N_2983,N_2955);
nor UO_228 (O_228,N_2995,N_2970);
or UO_229 (O_229,N_2965,N_2958);
or UO_230 (O_230,N_2978,N_2973);
or UO_231 (O_231,N_2951,N_2963);
nor UO_232 (O_232,N_2969,N_2989);
xnor UO_233 (O_233,N_2976,N_2960);
or UO_234 (O_234,N_2969,N_2952);
nor UO_235 (O_235,N_2962,N_2953);
nand UO_236 (O_236,N_2990,N_2951);
nand UO_237 (O_237,N_2972,N_2959);
nand UO_238 (O_238,N_2965,N_2998);
nor UO_239 (O_239,N_2963,N_2972);
and UO_240 (O_240,N_2967,N_2966);
nor UO_241 (O_241,N_2960,N_2969);
and UO_242 (O_242,N_2990,N_2955);
xor UO_243 (O_243,N_2951,N_2978);
or UO_244 (O_244,N_2953,N_2978);
and UO_245 (O_245,N_2990,N_2984);
and UO_246 (O_246,N_2994,N_2960);
or UO_247 (O_247,N_2954,N_2971);
nor UO_248 (O_248,N_2971,N_2991);
and UO_249 (O_249,N_2973,N_2984);
nor UO_250 (O_250,N_2980,N_2995);
or UO_251 (O_251,N_2957,N_2978);
xor UO_252 (O_252,N_2963,N_2964);
or UO_253 (O_253,N_2966,N_2980);
and UO_254 (O_254,N_2952,N_2963);
nand UO_255 (O_255,N_2966,N_2995);
or UO_256 (O_256,N_2994,N_2992);
or UO_257 (O_257,N_2962,N_2996);
and UO_258 (O_258,N_2969,N_2973);
nor UO_259 (O_259,N_2988,N_2989);
nor UO_260 (O_260,N_2960,N_2985);
nor UO_261 (O_261,N_2961,N_2984);
or UO_262 (O_262,N_2969,N_2950);
or UO_263 (O_263,N_2967,N_2991);
nor UO_264 (O_264,N_2992,N_2967);
or UO_265 (O_265,N_2962,N_2989);
nand UO_266 (O_266,N_2988,N_2975);
nor UO_267 (O_267,N_2954,N_2984);
nor UO_268 (O_268,N_2960,N_2998);
nand UO_269 (O_269,N_2963,N_2997);
or UO_270 (O_270,N_2975,N_2993);
and UO_271 (O_271,N_2985,N_2984);
or UO_272 (O_272,N_2967,N_2977);
and UO_273 (O_273,N_2954,N_2963);
xor UO_274 (O_274,N_2990,N_2961);
nand UO_275 (O_275,N_2991,N_2953);
or UO_276 (O_276,N_2979,N_2969);
nor UO_277 (O_277,N_2976,N_2993);
and UO_278 (O_278,N_2997,N_2973);
and UO_279 (O_279,N_2955,N_2989);
and UO_280 (O_280,N_2995,N_2963);
and UO_281 (O_281,N_2951,N_2995);
nand UO_282 (O_282,N_2991,N_2961);
nor UO_283 (O_283,N_2993,N_2959);
and UO_284 (O_284,N_2971,N_2960);
or UO_285 (O_285,N_2977,N_2971);
or UO_286 (O_286,N_2985,N_2968);
nor UO_287 (O_287,N_2991,N_2999);
nor UO_288 (O_288,N_2967,N_2963);
xor UO_289 (O_289,N_2997,N_2975);
xor UO_290 (O_290,N_2970,N_2987);
or UO_291 (O_291,N_2959,N_2956);
nand UO_292 (O_292,N_2963,N_2994);
or UO_293 (O_293,N_2991,N_2969);
nor UO_294 (O_294,N_2958,N_2955);
nor UO_295 (O_295,N_2995,N_2993);
nor UO_296 (O_296,N_2973,N_2989);
or UO_297 (O_297,N_2951,N_2956);
nor UO_298 (O_298,N_2987,N_2988);
nor UO_299 (O_299,N_2957,N_2960);
nor UO_300 (O_300,N_2981,N_2992);
xor UO_301 (O_301,N_2995,N_2962);
and UO_302 (O_302,N_2985,N_2969);
nand UO_303 (O_303,N_2982,N_2968);
xnor UO_304 (O_304,N_2952,N_2972);
or UO_305 (O_305,N_2975,N_2970);
and UO_306 (O_306,N_2984,N_2966);
or UO_307 (O_307,N_2979,N_2977);
nor UO_308 (O_308,N_2962,N_2956);
or UO_309 (O_309,N_2985,N_2995);
or UO_310 (O_310,N_2956,N_2979);
nor UO_311 (O_311,N_2993,N_2983);
nand UO_312 (O_312,N_2983,N_2985);
nand UO_313 (O_313,N_2989,N_2981);
and UO_314 (O_314,N_2992,N_2997);
nor UO_315 (O_315,N_2968,N_2989);
xor UO_316 (O_316,N_2969,N_2987);
or UO_317 (O_317,N_2990,N_2998);
nand UO_318 (O_318,N_2994,N_2952);
and UO_319 (O_319,N_2994,N_2972);
xor UO_320 (O_320,N_2976,N_2965);
or UO_321 (O_321,N_2955,N_2993);
and UO_322 (O_322,N_2953,N_2993);
and UO_323 (O_323,N_2994,N_2973);
or UO_324 (O_324,N_2966,N_2968);
or UO_325 (O_325,N_2954,N_2979);
nand UO_326 (O_326,N_2994,N_2965);
nor UO_327 (O_327,N_2982,N_2973);
and UO_328 (O_328,N_2988,N_2955);
nor UO_329 (O_329,N_2968,N_2960);
nor UO_330 (O_330,N_2977,N_2997);
nand UO_331 (O_331,N_2980,N_2959);
nor UO_332 (O_332,N_2983,N_2974);
or UO_333 (O_333,N_2989,N_2992);
or UO_334 (O_334,N_2974,N_2982);
nor UO_335 (O_335,N_2968,N_2961);
nor UO_336 (O_336,N_2961,N_2978);
and UO_337 (O_337,N_2977,N_2961);
nand UO_338 (O_338,N_2995,N_2959);
nand UO_339 (O_339,N_2973,N_2965);
and UO_340 (O_340,N_2992,N_2959);
xnor UO_341 (O_341,N_2972,N_2951);
and UO_342 (O_342,N_2965,N_2962);
nand UO_343 (O_343,N_2995,N_2979);
xnor UO_344 (O_344,N_2973,N_2987);
nand UO_345 (O_345,N_2991,N_2972);
nand UO_346 (O_346,N_2998,N_2953);
or UO_347 (O_347,N_2994,N_2962);
and UO_348 (O_348,N_2966,N_2983);
nand UO_349 (O_349,N_2960,N_2999);
xor UO_350 (O_350,N_2970,N_2961);
or UO_351 (O_351,N_2951,N_2957);
nor UO_352 (O_352,N_2963,N_2990);
and UO_353 (O_353,N_2992,N_2996);
nand UO_354 (O_354,N_2990,N_2994);
nor UO_355 (O_355,N_2985,N_2988);
and UO_356 (O_356,N_2980,N_2987);
nand UO_357 (O_357,N_2958,N_2976);
and UO_358 (O_358,N_2969,N_2957);
nor UO_359 (O_359,N_2955,N_2957);
and UO_360 (O_360,N_2958,N_2964);
nand UO_361 (O_361,N_2959,N_2964);
xor UO_362 (O_362,N_2964,N_2983);
xor UO_363 (O_363,N_2987,N_2989);
nor UO_364 (O_364,N_2978,N_2968);
nor UO_365 (O_365,N_2990,N_2986);
nor UO_366 (O_366,N_2998,N_2955);
or UO_367 (O_367,N_2997,N_2955);
xor UO_368 (O_368,N_2958,N_2999);
nand UO_369 (O_369,N_2987,N_2950);
xnor UO_370 (O_370,N_2950,N_2962);
nand UO_371 (O_371,N_2988,N_2971);
nor UO_372 (O_372,N_2989,N_2974);
and UO_373 (O_373,N_2969,N_2951);
nand UO_374 (O_374,N_2962,N_2979);
nand UO_375 (O_375,N_2970,N_2989);
and UO_376 (O_376,N_2976,N_2986);
nor UO_377 (O_377,N_2996,N_2986);
nor UO_378 (O_378,N_2964,N_2965);
nand UO_379 (O_379,N_2997,N_2960);
or UO_380 (O_380,N_2979,N_2990);
xnor UO_381 (O_381,N_2980,N_2967);
nand UO_382 (O_382,N_2960,N_2988);
nor UO_383 (O_383,N_2954,N_2959);
or UO_384 (O_384,N_2962,N_2990);
and UO_385 (O_385,N_2997,N_2951);
nor UO_386 (O_386,N_2988,N_2950);
nor UO_387 (O_387,N_2965,N_2967);
or UO_388 (O_388,N_2963,N_2960);
xor UO_389 (O_389,N_2992,N_2987);
nand UO_390 (O_390,N_2991,N_2977);
or UO_391 (O_391,N_2976,N_2995);
nor UO_392 (O_392,N_2969,N_2971);
xnor UO_393 (O_393,N_2983,N_2978);
and UO_394 (O_394,N_2972,N_2968);
or UO_395 (O_395,N_2969,N_2962);
and UO_396 (O_396,N_2962,N_2957);
and UO_397 (O_397,N_2979,N_2953);
nor UO_398 (O_398,N_2984,N_2993);
nor UO_399 (O_399,N_2954,N_2998);
xnor UO_400 (O_400,N_2987,N_2954);
nor UO_401 (O_401,N_2954,N_2964);
nand UO_402 (O_402,N_2969,N_2988);
nand UO_403 (O_403,N_2991,N_2952);
or UO_404 (O_404,N_2998,N_2951);
and UO_405 (O_405,N_2992,N_2971);
and UO_406 (O_406,N_2999,N_2978);
xnor UO_407 (O_407,N_2957,N_2977);
nand UO_408 (O_408,N_2967,N_2950);
and UO_409 (O_409,N_2989,N_2959);
and UO_410 (O_410,N_2964,N_2995);
nor UO_411 (O_411,N_2961,N_2989);
nor UO_412 (O_412,N_2963,N_2984);
nor UO_413 (O_413,N_2990,N_2989);
and UO_414 (O_414,N_2965,N_2951);
xor UO_415 (O_415,N_2990,N_2967);
nor UO_416 (O_416,N_2986,N_2960);
and UO_417 (O_417,N_2966,N_2987);
or UO_418 (O_418,N_2981,N_2952);
nand UO_419 (O_419,N_2951,N_2981);
nor UO_420 (O_420,N_2971,N_2974);
and UO_421 (O_421,N_2975,N_2995);
nor UO_422 (O_422,N_2963,N_2950);
nor UO_423 (O_423,N_2976,N_2982);
or UO_424 (O_424,N_2971,N_2970);
nor UO_425 (O_425,N_2962,N_2970);
or UO_426 (O_426,N_2958,N_2994);
or UO_427 (O_427,N_2982,N_2963);
or UO_428 (O_428,N_2959,N_2967);
xnor UO_429 (O_429,N_2950,N_2972);
and UO_430 (O_430,N_2973,N_2991);
nor UO_431 (O_431,N_2977,N_2951);
nor UO_432 (O_432,N_2956,N_2966);
nand UO_433 (O_433,N_2990,N_2996);
and UO_434 (O_434,N_2986,N_2985);
nor UO_435 (O_435,N_2990,N_2978);
or UO_436 (O_436,N_2982,N_2984);
or UO_437 (O_437,N_2983,N_2995);
xnor UO_438 (O_438,N_2980,N_2989);
and UO_439 (O_439,N_2984,N_2987);
nand UO_440 (O_440,N_2967,N_2961);
nor UO_441 (O_441,N_2981,N_2954);
nand UO_442 (O_442,N_2961,N_2985);
xnor UO_443 (O_443,N_2989,N_2952);
and UO_444 (O_444,N_2964,N_2982);
and UO_445 (O_445,N_2985,N_2966);
and UO_446 (O_446,N_2957,N_2950);
or UO_447 (O_447,N_2952,N_2966);
nor UO_448 (O_448,N_2967,N_2978);
nand UO_449 (O_449,N_2989,N_2967);
and UO_450 (O_450,N_2987,N_2972);
nand UO_451 (O_451,N_2960,N_2975);
or UO_452 (O_452,N_2972,N_2999);
nor UO_453 (O_453,N_2995,N_2969);
or UO_454 (O_454,N_2970,N_2994);
or UO_455 (O_455,N_2965,N_2969);
nand UO_456 (O_456,N_2990,N_2953);
nor UO_457 (O_457,N_2972,N_2967);
or UO_458 (O_458,N_2978,N_2984);
nand UO_459 (O_459,N_2959,N_2961);
or UO_460 (O_460,N_2991,N_2997);
and UO_461 (O_461,N_2955,N_2970);
and UO_462 (O_462,N_2981,N_2950);
and UO_463 (O_463,N_2953,N_2994);
or UO_464 (O_464,N_2976,N_2964);
and UO_465 (O_465,N_2956,N_2984);
nand UO_466 (O_466,N_2966,N_2971);
nor UO_467 (O_467,N_2950,N_2978);
and UO_468 (O_468,N_2970,N_2973);
xor UO_469 (O_469,N_2997,N_2998);
and UO_470 (O_470,N_2994,N_2981);
and UO_471 (O_471,N_2982,N_2958);
xor UO_472 (O_472,N_2973,N_2968);
xnor UO_473 (O_473,N_2997,N_2962);
xor UO_474 (O_474,N_2980,N_2958);
xor UO_475 (O_475,N_2950,N_2965);
nand UO_476 (O_476,N_2996,N_2965);
nor UO_477 (O_477,N_2979,N_2982);
nand UO_478 (O_478,N_2976,N_2991);
xnor UO_479 (O_479,N_2994,N_2975);
xor UO_480 (O_480,N_2995,N_2957);
and UO_481 (O_481,N_2976,N_2956);
nor UO_482 (O_482,N_2972,N_2983);
or UO_483 (O_483,N_2981,N_2985);
or UO_484 (O_484,N_2976,N_2977);
nand UO_485 (O_485,N_2986,N_2952);
or UO_486 (O_486,N_2988,N_2951);
and UO_487 (O_487,N_2974,N_2992);
nand UO_488 (O_488,N_2987,N_2995);
xor UO_489 (O_489,N_2991,N_2993);
xor UO_490 (O_490,N_2999,N_2992);
nand UO_491 (O_491,N_2998,N_2957);
or UO_492 (O_492,N_2999,N_2984);
nand UO_493 (O_493,N_2980,N_2979);
nand UO_494 (O_494,N_2955,N_2950);
or UO_495 (O_495,N_2960,N_2958);
and UO_496 (O_496,N_2971,N_2983);
xnor UO_497 (O_497,N_2952,N_2954);
nand UO_498 (O_498,N_2977,N_2974);
and UO_499 (O_499,N_2984,N_2972);
endmodule