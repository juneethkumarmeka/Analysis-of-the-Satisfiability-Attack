module basic_500_3000_500_3_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_341,In_470);
or U1 (N_1,In_374,In_131);
xor U2 (N_2,In_132,In_334);
and U3 (N_3,In_199,In_256);
nor U4 (N_4,In_177,In_323);
or U5 (N_5,In_178,In_349);
and U6 (N_6,In_93,In_104);
nor U7 (N_7,In_432,In_33);
nand U8 (N_8,In_152,In_15);
nand U9 (N_9,In_148,In_480);
nor U10 (N_10,In_51,In_316);
xnor U11 (N_11,In_386,In_494);
or U12 (N_12,In_207,In_7);
xnor U13 (N_13,In_41,In_422);
nor U14 (N_14,In_263,In_21);
nor U15 (N_15,In_311,In_390);
and U16 (N_16,In_72,In_388);
nand U17 (N_17,In_373,In_195);
and U18 (N_18,In_279,In_300);
nor U19 (N_19,In_85,In_429);
and U20 (N_20,In_380,In_428);
xnor U21 (N_21,In_3,In_483);
xnor U22 (N_22,In_205,In_450);
and U23 (N_23,In_100,In_83);
xnor U24 (N_24,In_184,In_162);
nand U25 (N_25,In_427,In_4);
nand U26 (N_26,In_324,In_92);
nand U27 (N_27,In_435,In_319);
xnor U28 (N_28,In_317,In_116);
or U29 (N_29,In_475,In_262);
nand U30 (N_30,In_20,In_16);
nand U31 (N_31,In_457,In_473);
or U32 (N_32,In_322,In_98);
or U33 (N_33,In_117,In_232);
nand U34 (N_34,In_168,In_102);
nor U35 (N_35,In_347,In_387);
or U36 (N_36,In_74,In_155);
nand U37 (N_37,In_46,In_19);
xnor U38 (N_38,In_165,In_124);
nor U39 (N_39,In_249,In_411);
nor U40 (N_40,In_180,In_325);
nor U41 (N_41,In_298,In_56);
and U42 (N_42,In_440,In_101);
and U43 (N_43,In_42,In_35);
or U44 (N_44,In_136,In_237);
nor U45 (N_45,In_448,In_273);
and U46 (N_46,In_71,In_488);
nor U47 (N_47,In_143,In_357);
and U48 (N_48,In_14,In_350);
nor U49 (N_49,In_467,In_406);
xnor U50 (N_50,In_153,In_458);
nand U51 (N_51,In_326,In_496);
and U52 (N_52,In_245,In_287);
nand U53 (N_53,In_377,In_80);
or U54 (N_54,In_268,In_353);
nand U55 (N_55,In_487,In_306);
or U56 (N_56,In_416,In_340);
or U57 (N_57,In_454,In_354);
nand U58 (N_58,In_461,In_108);
nand U59 (N_59,In_186,In_352);
nor U60 (N_60,In_425,In_295);
or U61 (N_61,In_211,In_369);
and U62 (N_62,In_399,In_360);
nand U63 (N_63,In_90,In_27);
or U64 (N_64,In_40,In_275);
and U65 (N_65,In_361,In_243);
and U66 (N_66,In_172,In_410);
nand U67 (N_67,In_413,In_459);
and U68 (N_68,In_289,In_217);
and U69 (N_69,In_52,In_121);
nor U70 (N_70,In_368,In_370);
nor U71 (N_71,In_79,In_156);
xor U72 (N_72,In_414,In_401);
nor U73 (N_73,In_105,In_299);
or U74 (N_74,In_261,In_106);
or U75 (N_75,In_490,In_478);
and U76 (N_76,In_333,In_332);
xor U77 (N_77,In_320,In_392);
nand U78 (N_78,In_179,In_315);
xor U79 (N_79,In_331,In_48);
nand U80 (N_80,In_5,In_53);
nand U81 (N_81,In_460,In_69);
xnor U82 (N_82,In_145,In_75);
or U83 (N_83,In_118,In_222);
or U84 (N_84,In_173,In_38);
nor U85 (N_85,In_498,In_88);
nor U86 (N_86,In_359,In_11);
nand U87 (N_87,In_305,In_127);
or U88 (N_88,In_215,In_336);
nand U89 (N_89,In_321,In_81);
nor U90 (N_90,In_492,In_433);
nand U91 (N_91,In_125,In_286);
xor U92 (N_92,In_238,In_327);
nor U93 (N_93,In_398,In_246);
nand U94 (N_94,In_170,In_96);
nor U95 (N_95,In_407,In_120);
nand U96 (N_96,In_194,In_472);
or U97 (N_97,In_240,In_45);
and U98 (N_98,In_111,In_54);
nand U99 (N_99,In_267,In_351);
or U100 (N_100,In_229,In_201);
or U101 (N_101,In_66,In_329);
or U102 (N_102,In_95,In_364);
and U103 (N_103,In_122,In_154);
or U104 (N_104,In_394,In_474);
or U105 (N_105,In_420,In_452);
and U106 (N_106,In_218,In_157);
or U107 (N_107,In_250,In_200);
nand U108 (N_108,In_231,In_216);
or U109 (N_109,In_59,In_50);
or U110 (N_110,In_109,In_130);
nor U111 (N_111,In_346,In_70);
nand U112 (N_112,In_419,In_26);
and U113 (N_113,In_139,In_495);
and U114 (N_114,In_424,In_451);
and U115 (N_115,In_444,In_77);
nor U116 (N_116,In_241,In_174);
or U117 (N_117,In_313,In_277);
or U118 (N_118,In_185,In_146);
and U119 (N_119,In_337,In_383);
nor U120 (N_120,In_375,In_129);
and U121 (N_121,In_36,In_303);
nor U122 (N_122,In_192,In_363);
and U123 (N_123,In_187,In_61);
and U124 (N_124,In_438,In_292);
and U125 (N_125,In_34,In_288);
nand U126 (N_126,In_9,In_396);
nor U127 (N_127,In_455,In_119);
or U128 (N_128,In_482,In_198);
nor U129 (N_129,In_31,In_82);
nor U130 (N_130,In_191,In_114);
and U131 (N_131,In_22,In_115);
nand U132 (N_132,In_356,In_468);
and U133 (N_133,In_190,In_138);
and U134 (N_134,In_437,In_389);
xor U135 (N_135,In_23,In_29);
nand U136 (N_136,In_339,In_28);
nand U137 (N_137,In_338,In_134);
nand U138 (N_138,In_196,In_447);
nor U139 (N_139,In_208,In_110);
nor U140 (N_140,In_381,In_436);
nand U141 (N_141,In_293,In_342);
and U142 (N_142,In_248,In_160);
or U143 (N_143,In_404,In_376);
xor U144 (N_144,In_466,In_149);
nand U145 (N_145,In_44,In_228);
and U146 (N_146,In_255,In_158);
or U147 (N_147,In_465,In_214);
and U148 (N_148,In_37,In_169);
nand U149 (N_149,In_304,In_135);
or U150 (N_150,In_309,In_89);
nand U151 (N_151,In_391,In_280);
xor U152 (N_152,In_113,In_78);
or U153 (N_153,In_441,In_123);
nor U154 (N_154,In_290,In_234);
or U155 (N_155,In_203,In_202);
nor U156 (N_156,In_8,In_285);
and U157 (N_157,In_239,In_126);
nand U158 (N_158,In_445,In_302);
and U159 (N_159,In_348,In_18);
nor U160 (N_160,In_282,In_133);
nand U161 (N_161,In_439,In_251);
nor U162 (N_162,In_378,In_67);
or U163 (N_163,In_272,In_367);
nor U164 (N_164,In_224,In_371);
or U165 (N_165,In_366,In_330);
and U166 (N_166,In_225,In_264);
nand U167 (N_167,In_84,In_39);
xor U168 (N_168,In_87,In_63);
nor U169 (N_169,In_230,In_385);
and U170 (N_170,In_462,In_400);
nor U171 (N_171,In_212,In_463);
and U172 (N_172,In_164,In_242);
nand U173 (N_173,In_395,In_477);
and U174 (N_174,In_297,In_365);
nand U175 (N_175,In_144,In_171);
nand U176 (N_176,In_484,In_12);
or U177 (N_177,In_479,In_210);
or U178 (N_178,In_247,In_13);
nand U179 (N_179,In_57,In_274);
or U180 (N_180,In_25,In_2);
or U181 (N_181,In_499,In_30);
or U182 (N_182,In_76,In_476);
nor U183 (N_183,In_308,In_58);
xor U184 (N_184,In_204,In_403);
xnor U185 (N_185,In_393,In_65);
nand U186 (N_186,In_271,In_464);
or U187 (N_187,In_449,In_252);
nand U188 (N_188,In_163,In_276);
nand U189 (N_189,In_379,In_235);
nand U190 (N_190,In_497,In_259);
and U191 (N_191,In_423,In_91);
nand U192 (N_192,In_345,In_426);
nand U193 (N_193,In_183,In_60);
xor U194 (N_194,In_412,In_97);
and U195 (N_195,In_107,In_32);
or U196 (N_196,In_193,In_206);
nand U197 (N_197,In_372,In_0);
nand U198 (N_198,In_254,In_141);
and U199 (N_199,In_49,In_291);
nor U200 (N_200,In_446,In_397);
nand U201 (N_201,In_226,In_128);
or U202 (N_202,In_434,In_481);
or U203 (N_203,In_94,In_167);
and U204 (N_204,In_142,In_453);
and U205 (N_205,In_213,In_1);
or U206 (N_206,In_197,In_418);
or U207 (N_207,In_335,In_258);
nor U208 (N_208,In_415,In_266);
or U209 (N_209,In_312,In_485);
nand U210 (N_210,In_278,In_281);
and U211 (N_211,In_318,In_344);
nor U212 (N_212,In_188,In_219);
nand U213 (N_213,In_17,In_62);
and U214 (N_214,In_233,In_159);
and U215 (N_215,In_10,In_469);
nor U216 (N_216,In_175,In_431);
nor U217 (N_217,In_310,In_112);
or U218 (N_218,In_384,In_417);
nand U219 (N_219,In_236,In_284);
nand U220 (N_220,In_283,In_68);
nand U221 (N_221,In_221,In_176);
and U222 (N_222,In_189,In_301);
and U223 (N_223,In_55,In_296);
and U224 (N_224,In_421,In_489);
nand U225 (N_225,In_64,In_103);
and U226 (N_226,In_181,In_150);
nand U227 (N_227,In_294,In_151);
and U228 (N_228,In_355,In_430);
and U229 (N_229,In_314,In_140);
and U230 (N_230,In_257,In_402);
nor U231 (N_231,In_307,In_409);
and U232 (N_232,In_47,In_161);
or U233 (N_233,In_6,In_73);
nand U234 (N_234,In_24,In_358);
and U235 (N_235,In_270,In_269);
and U236 (N_236,In_443,In_220);
nor U237 (N_237,In_166,In_471);
and U238 (N_238,In_405,In_265);
nand U239 (N_239,In_343,In_362);
nor U240 (N_240,In_408,In_182);
nor U241 (N_241,In_260,In_137);
nor U242 (N_242,In_86,In_442);
nor U243 (N_243,In_486,In_209);
or U244 (N_244,In_99,In_223);
nor U245 (N_245,In_227,In_244);
or U246 (N_246,In_253,In_493);
and U247 (N_247,In_456,In_43);
nor U248 (N_248,In_147,In_328);
or U249 (N_249,In_382,In_491);
nand U250 (N_250,In_79,In_353);
nand U251 (N_251,In_188,In_353);
or U252 (N_252,In_4,In_173);
and U253 (N_253,In_124,In_317);
nand U254 (N_254,In_170,In_42);
or U255 (N_255,In_296,In_285);
and U256 (N_256,In_102,In_327);
nand U257 (N_257,In_167,In_47);
nand U258 (N_258,In_135,In_357);
xnor U259 (N_259,In_74,In_205);
nor U260 (N_260,In_412,In_21);
or U261 (N_261,In_380,In_442);
and U262 (N_262,In_328,In_437);
and U263 (N_263,In_336,In_273);
and U264 (N_264,In_420,In_130);
nor U265 (N_265,In_228,In_321);
and U266 (N_266,In_235,In_221);
nand U267 (N_267,In_167,In_87);
or U268 (N_268,In_336,In_368);
nand U269 (N_269,In_173,In_58);
and U270 (N_270,In_242,In_376);
and U271 (N_271,In_41,In_114);
xnor U272 (N_272,In_438,In_70);
xnor U273 (N_273,In_332,In_52);
or U274 (N_274,In_37,In_468);
nand U275 (N_275,In_223,In_426);
or U276 (N_276,In_381,In_201);
nor U277 (N_277,In_307,In_48);
nor U278 (N_278,In_393,In_236);
nand U279 (N_279,In_383,In_281);
or U280 (N_280,In_101,In_180);
nor U281 (N_281,In_291,In_2);
nor U282 (N_282,In_228,In_155);
xor U283 (N_283,In_381,In_407);
and U284 (N_284,In_68,In_429);
xor U285 (N_285,In_262,In_202);
xnor U286 (N_286,In_349,In_434);
or U287 (N_287,In_116,In_341);
and U288 (N_288,In_392,In_383);
and U289 (N_289,In_11,In_320);
nand U290 (N_290,In_395,In_380);
nand U291 (N_291,In_200,In_203);
nand U292 (N_292,In_461,In_49);
nand U293 (N_293,In_86,In_110);
nor U294 (N_294,In_112,In_106);
nand U295 (N_295,In_440,In_73);
nand U296 (N_296,In_341,In_227);
and U297 (N_297,In_56,In_381);
nand U298 (N_298,In_302,In_146);
nand U299 (N_299,In_124,In_401);
nand U300 (N_300,In_328,In_360);
and U301 (N_301,In_353,In_481);
nand U302 (N_302,In_306,In_131);
xnor U303 (N_303,In_261,In_322);
or U304 (N_304,In_453,In_432);
or U305 (N_305,In_294,In_218);
or U306 (N_306,In_207,In_46);
xor U307 (N_307,In_441,In_68);
and U308 (N_308,In_471,In_276);
and U309 (N_309,In_489,In_419);
and U310 (N_310,In_411,In_378);
nand U311 (N_311,In_102,In_455);
nor U312 (N_312,In_35,In_242);
nand U313 (N_313,In_399,In_327);
nor U314 (N_314,In_294,In_63);
nand U315 (N_315,In_251,In_487);
and U316 (N_316,In_238,In_141);
nand U317 (N_317,In_384,In_305);
nor U318 (N_318,In_495,In_24);
xor U319 (N_319,In_356,In_277);
nor U320 (N_320,In_368,In_376);
nor U321 (N_321,In_483,In_422);
nor U322 (N_322,In_381,In_58);
nor U323 (N_323,In_318,In_32);
nand U324 (N_324,In_382,In_44);
or U325 (N_325,In_445,In_357);
nand U326 (N_326,In_62,In_230);
nand U327 (N_327,In_418,In_149);
nor U328 (N_328,In_136,In_119);
nand U329 (N_329,In_340,In_8);
xor U330 (N_330,In_132,In_497);
or U331 (N_331,In_114,In_76);
or U332 (N_332,In_301,In_182);
nor U333 (N_333,In_303,In_170);
nand U334 (N_334,In_42,In_131);
or U335 (N_335,In_74,In_499);
nor U336 (N_336,In_18,In_173);
and U337 (N_337,In_482,In_76);
and U338 (N_338,In_120,In_105);
and U339 (N_339,In_328,In_76);
or U340 (N_340,In_141,In_27);
nand U341 (N_341,In_68,In_407);
nor U342 (N_342,In_282,In_35);
nor U343 (N_343,In_81,In_392);
xor U344 (N_344,In_130,In_475);
and U345 (N_345,In_438,In_419);
and U346 (N_346,In_273,In_338);
xnor U347 (N_347,In_144,In_346);
nor U348 (N_348,In_105,In_8);
or U349 (N_349,In_376,In_296);
nand U350 (N_350,In_100,In_336);
or U351 (N_351,In_426,In_30);
nor U352 (N_352,In_249,In_430);
xnor U353 (N_353,In_33,In_486);
or U354 (N_354,In_386,In_474);
or U355 (N_355,In_327,In_340);
xnor U356 (N_356,In_388,In_446);
or U357 (N_357,In_412,In_354);
or U358 (N_358,In_220,In_59);
and U359 (N_359,In_499,In_43);
xor U360 (N_360,In_48,In_308);
and U361 (N_361,In_80,In_6);
or U362 (N_362,In_429,In_417);
or U363 (N_363,In_383,In_294);
or U364 (N_364,In_304,In_198);
and U365 (N_365,In_375,In_90);
and U366 (N_366,In_436,In_374);
or U367 (N_367,In_240,In_259);
and U368 (N_368,In_39,In_359);
xnor U369 (N_369,In_157,In_282);
or U370 (N_370,In_142,In_381);
nand U371 (N_371,In_309,In_12);
nor U372 (N_372,In_426,In_227);
nand U373 (N_373,In_307,In_277);
or U374 (N_374,In_332,In_79);
or U375 (N_375,In_161,In_365);
nand U376 (N_376,In_382,In_310);
or U377 (N_377,In_251,In_82);
nand U378 (N_378,In_426,In_207);
nand U379 (N_379,In_30,In_393);
nand U380 (N_380,In_253,In_381);
or U381 (N_381,In_239,In_19);
nand U382 (N_382,In_202,In_369);
nand U383 (N_383,In_220,In_188);
xnor U384 (N_384,In_360,In_131);
and U385 (N_385,In_269,In_24);
nand U386 (N_386,In_169,In_306);
nor U387 (N_387,In_83,In_216);
nand U388 (N_388,In_266,In_109);
or U389 (N_389,In_239,In_438);
or U390 (N_390,In_26,In_205);
and U391 (N_391,In_407,In_88);
or U392 (N_392,In_2,In_399);
nor U393 (N_393,In_99,In_74);
and U394 (N_394,In_251,In_156);
nor U395 (N_395,In_67,In_458);
nand U396 (N_396,In_132,In_236);
nor U397 (N_397,In_122,In_269);
nor U398 (N_398,In_272,In_185);
or U399 (N_399,In_316,In_213);
or U400 (N_400,In_348,In_145);
or U401 (N_401,In_332,In_166);
or U402 (N_402,In_210,In_365);
or U403 (N_403,In_395,In_203);
nand U404 (N_404,In_101,In_244);
nor U405 (N_405,In_10,In_381);
and U406 (N_406,In_11,In_291);
nor U407 (N_407,In_289,In_484);
or U408 (N_408,In_102,In_385);
and U409 (N_409,In_248,In_66);
or U410 (N_410,In_243,In_293);
nor U411 (N_411,In_415,In_349);
or U412 (N_412,In_41,In_370);
nor U413 (N_413,In_404,In_354);
xnor U414 (N_414,In_246,In_67);
nand U415 (N_415,In_416,In_401);
or U416 (N_416,In_313,In_194);
or U417 (N_417,In_196,In_171);
or U418 (N_418,In_340,In_34);
or U419 (N_419,In_19,In_108);
xor U420 (N_420,In_65,In_459);
nor U421 (N_421,In_62,In_200);
or U422 (N_422,In_447,In_491);
nand U423 (N_423,In_42,In_378);
and U424 (N_424,In_299,In_49);
or U425 (N_425,In_238,In_445);
nand U426 (N_426,In_102,In_187);
nand U427 (N_427,In_401,In_489);
nor U428 (N_428,In_117,In_366);
nor U429 (N_429,In_99,In_39);
or U430 (N_430,In_174,In_93);
nor U431 (N_431,In_257,In_6);
nor U432 (N_432,In_297,In_50);
nand U433 (N_433,In_217,In_8);
nand U434 (N_434,In_347,In_416);
nand U435 (N_435,In_376,In_231);
and U436 (N_436,In_10,In_458);
or U437 (N_437,In_197,In_336);
nand U438 (N_438,In_297,In_111);
nor U439 (N_439,In_455,In_483);
and U440 (N_440,In_446,In_381);
xor U441 (N_441,In_91,In_140);
nor U442 (N_442,In_426,In_463);
or U443 (N_443,In_81,In_452);
and U444 (N_444,In_302,In_185);
or U445 (N_445,In_444,In_320);
nor U446 (N_446,In_233,In_444);
xnor U447 (N_447,In_191,In_416);
or U448 (N_448,In_21,In_265);
nor U449 (N_449,In_325,In_133);
and U450 (N_450,In_32,In_154);
and U451 (N_451,In_324,In_272);
and U452 (N_452,In_154,In_446);
nand U453 (N_453,In_470,In_107);
nor U454 (N_454,In_124,In_223);
nand U455 (N_455,In_134,In_314);
and U456 (N_456,In_340,In_404);
nor U457 (N_457,In_192,In_441);
nor U458 (N_458,In_44,In_229);
or U459 (N_459,In_267,In_478);
and U460 (N_460,In_444,In_368);
and U461 (N_461,In_15,In_345);
and U462 (N_462,In_31,In_469);
nand U463 (N_463,In_79,In_292);
or U464 (N_464,In_387,In_369);
nor U465 (N_465,In_326,In_262);
nor U466 (N_466,In_12,In_352);
and U467 (N_467,In_196,In_133);
and U468 (N_468,In_498,In_481);
and U469 (N_469,In_446,In_344);
nand U470 (N_470,In_319,In_84);
and U471 (N_471,In_110,In_452);
nand U472 (N_472,In_164,In_179);
nand U473 (N_473,In_169,In_90);
nor U474 (N_474,In_180,In_141);
or U475 (N_475,In_337,In_223);
or U476 (N_476,In_453,In_411);
nand U477 (N_477,In_256,In_132);
nor U478 (N_478,In_86,In_81);
nand U479 (N_479,In_183,In_423);
nor U480 (N_480,In_299,In_83);
nor U481 (N_481,In_3,In_240);
and U482 (N_482,In_268,In_177);
nand U483 (N_483,In_476,In_159);
and U484 (N_484,In_398,In_193);
or U485 (N_485,In_158,In_162);
nand U486 (N_486,In_148,In_291);
nor U487 (N_487,In_88,In_206);
and U488 (N_488,In_21,In_475);
nor U489 (N_489,In_341,In_456);
or U490 (N_490,In_156,In_194);
or U491 (N_491,In_110,In_269);
nor U492 (N_492,In_375,In_207);
nor U493 (N_493,In_210,In_187);
nand U494 (N_494,In_202,In_58);
xnor U495 (N_495,In_26,In_374);
nor U496 (N_496,In_110,In_384);
nor U497 (N_497,In_162,In_279);
or U498 (N_498,In_292,In_484);
or U499 (N_499,In_55,In_95);
nor U500 (N_500,In_141,In_211);
and U501 (N_501,In_454,In_112);
or U502 (N_502,In_443,In_242);
and U503 (N_503,In_362,In_241);
nor U504 (N_504,In_184,In_285);
and U505 (N_505,In_323,In_480);
nand U506 (N_506,In_281,In_171);
nand U507 (N_507,In_414,In_264);
or U508 (N_508,In_166,In_417);
nor U509 (N_509,In_367,In_120);
nor U510 (N_510,In_321,In_419);
and U511 (N_511,In_303,In_239);
nor U512 (N_512,In_217,In_130);
nor U513 (N_513,In_270,In_169);
nor U514 (N_514,In_105,In_491);
and U515 (N_515,In_9,In_96);
and U516 (N_516,In_0,In_282);
nor U517 (N_517,In_48,In_67);
nand U518 (N_518,In_80,In_48);
and U519 (N_519,In_337,In_481);
nor U520 (N_520,In_483,In_133);
xor U521 (N_521,In_278,In_445);
or U522 (N_522,In_292,In_10);
and U523 (N_523,In_234,In_327);
nor U524 (N_524,In_127,In_313);
nor U525 (N_525,In_40,In_205);
nand U526 (N_526,In_330,In_352);
nor U527 (N_527,In_7,In_251);
and U528 (N_528,In_219,In_361);
or U529 (N_529,In_267,In_74);
xor U530 (N_530,In_19,In_448);
nor U531 (N_531,In_166,In_127);
and U532 (N_532,In_394,In_364);
nand U533 (N_533,In_33,In_266);
nand U534 (N_534,In_315,In_289);
and U535 (N_535,In_326,In_389);
nor U536 (N_536,In_142,In_286);
and U537 (N_537,In_129,In_228);
nand U538 (N_538,In_161,In_342);
nor U539 (N_539,In_485,In_309);
and U540 (N_540,In_477,In_434);
nor U541 (N_541,In_35,In_100);
or U542 (N_542,In_36,In_185);
nand U543 (N_543,In_332,In_187);
nor U544 (N_544,In_383,In_452);
and U545 (N_545,In_184,In_397);
or U546 (N_546,In_294,In_105);
or U547 (N_547,In_182,In_329);
nor U548 (N_548,In_194,In_44);
and U549 (N_549,In_192,In_278);
nand U550 (N_550,In_70,In_382);
nand U551 (N_551,In_116,In_320);
xor U552 (N_552,In_356,In_53);
nor U553 (N_553,In_196,In_69);
or U554 (N_554,In_34,In_313);
and U555 (N_555,In_205,In_469);
and U556 (N_556,In_223,In_168);
nor U557 (N_557,In_258,In_117);
nand U558 (N_558,In_375,In_262);
nand U559 (N_559,In_1,In_147);
nor U560 (N_560,In_112,In_442);
or U561 (N_561,In_490,In_213);
nor U562 (N_562,In_148,In_283);
nand U563 (N_563,In_286,In_452);
and U564 (N_564,In_416,In_202);
and U565 (N_565,In_429,In_269);
or U566 (N_566,In_456,In_106);
and U567 (N_567,In_425,In_190);
nand U568 (N_568,In_204,In_30);
xnor U569 (N_569,In_349,In_330);
nand U570 (N_570,In_310,In_477);
nand U571 (N_571,In_50,In_148);
nand U572 (N_572,In_495,In_367);
xnor U573 (N_573,In_224,In_368);
nand U574 (N_574,In_353,In_465);
nor U575 (N_575,In_167,In_456);
nand U576 (N_576,In_2,In_494);
and U577 (N_577,In_392,In_473);
or U578 (N_578,In_72,In_128);
nor U579 (N_579,In_456,In_84);
or U580 (N_580,In_371,In_148);
or U581 (N_581,In_101,In_194);
or U582 (N_582,In_348,In_301);
nand U583 (N_583,In_249,In_36);
nor U584 (N_584,In_54,In_30);
xnor U585 (N_585,In_394,In_483);
nand U586 (N_586,In_279,In_294);
and U587 (N_587,In_278,In_274);
nand U588 (N_588,In_275,In_236);
nor U589 (N_589,In_415,In_462);
or U590 (N_590,In_191,In_403);
nor U591 (N_591,In_316,In_77);
nand U592 (N_592,In_224,In_92);
or U593 (N_593,In_213,In_325);
nor U594 (N_594,In_437,In_1);
or U595 (N_595,In_0,In_137);
nand U596 (N_596,In_479,In_444);
xor U597 (N_597,In_70,In_394);
or U598 (N_598,In_468,In_329);
or U599 (N_599,In_121,In_392);
and U600 (N_600,In_218,In_85);
nor U601 (N_601,In_87,In_435);
nor U602 (N_602,In_123,In_146);
nand U603 (N_603,In_442,In_66);
nor U604 (N_604,In_257,In_322);
nand U605 (N_605,In_107,In_229);
xnor U606 (N_606,In_493,In_404);
nor U607 (N_607,In_343,In_390);
or U608 (N_608,In_118,In_306);
nand U609 (N_609,In_54,In_302);
nor U610 (N_610,In_306,In_254);
or U611 (N_611,In_396,In_272);
and U612 (N_612,In_121,In_40);
or U613 (N_613,In_477,In_256);
and U614 (N_614,In_251,In_486);
or U615 (N_615,In_397,In_70);
nor U616 (N_616,In_456,In_424);
and U617 (N_617,In_377,In_407);
nand U618 (N_618,In_37,In_327);
or U619 (N_619,In_262,In_89);
nor U620 (N_620,In_72,In_487);
nor U621 (N_621,In_438,In_40);
nor U622 (N_622,In_494,In_306);
nand U623 (N_623,In_21,In_353);
nand U624 (N_624,In_299,In_420);
nor U625 (N_625,In_140,In_84);
nor U626 (N_626,In_297,In_428);
nand U627 (N_627,In_305,In_265);
nand U628 (N_628,In_4,In_37);
or U629 (N_629,In_142,In_166);
xor U630 (N_630,In_211,In_174);
or U631 (N_631,In_155,In_270);
xnor U632 (N_632,In_78,In_192);
and U633 (N_633,In_184,In_54);
nor U634 (N_634,In_244,In_28);
nor U635 (N_635,In_299,In_116);
xor U636 (N_636,In_286,In_199);
xnor U637 (N_637,In_461,In_481);
nand U638 (N_638,In_377,In_43);
nor U639 (N_639,In_422,In_266);
nand U640 (N_640,In_374,In_279);
nand U641 (N_641,In_160,In_341);
nand U642 (N_642,In_172,In_48);
and U643 (N_643,In_313,In_347);
nand U644 (N_644,In_344,In_414);
xor U645 (N_645,In_70,In_493);
and U646 (N_646,In_228,In_471);
nand U647 (N_647,In_87,In_64);
nand U648 (N_648,In_336,In_177);
and U649 (N_649,In_213,In_347);
nand U650 (N_650,In_120,In_9);
or U651 (N_651,In_449,In_156);
nand U652 (N_652,In_319,In_67);
nand U653 (N_653,In_315,In_203);
xor U654 (N_654,In_322,In_89);
nor U655 (N_655,In_320,In_297);
nor U656 (N_656,In_305,In_190);
nand U657 (N_657,In_374,In_420);
and U658 (N_658,In_250,In_430);
and U659 (N_659,In_311,In_183);
xnor U660 (N_660,In_250,In_427);
and U661 (N_661,In_105,In_11);
nor U662 (N_662,In_71,In_456);
nor U663 (N_663,In_467,In_495);
nand U664 (N_664,In_69,In_435);
xnor U665 (N_665,In_292,In_329);
nor U666 (N_666,In_282,In_190);
nand U667 (N_667,In_92,In_72);
xnor U668 (N_668,In_255,In_405);
and U669 (N_669,In_428,In_280);
or U670 (N_670,In_167,In_266);
nor U671 (N_671,In_298,In_55);
and U672 (N_672,In_115,In_149);
nor U673 (N_673,In_217,In_112);
xnor U674 (N_674,In_296,In_167);
and U675 (N_675,In_32,In_183);
or U676 (N_676,In_178,In_84);
or U677 (N_677,In_250,In_390);
nand U678 (N_678,In_293,In_109);
nand U679 (N_679,In_219,In_259);
xnor U680 (N_680,In_37,In_256);
and U681 (N_681,In_95,In_398);
or U682 (N_682,In_40,In_8);
and U683 (N_683,In_130,In_333);
xnor U684 (N_684,In_431,In_316);
or U685 (N_685,In_318,In_268);
or U686 (N_686,In_343,In_301);
xnor U687 (N_687,In_175,In_372);
nand U688 (N_688,In_137,In_55);
or U689 (N_689,In_39,In_18);
nor U690 (N_690,In_439,In_466);
or U691 (N_691,In_429,In_290);
and U692 (N_692,In_50,In_468);
and U693 (N_693,In_476,In_67);
or U694 (N_694,In_100,In_394);
nor U695 (N_695,In_238,In_173);
and U696 (N_696,In_415,In_369);
or U697 (N_697,In_299,In_479);
or U698 (N_698,In_106,In_373);
and U699 (N_699,In_225,In_250);
or U700 (N_700,In_12,In_232);
nor U701 (N_701,In_346,In_401);
xor U702 (N_702,In_81,In_67);
and U703 (N_703,In_83,In_223);
and U704 (N_704,In_120,In_487);
xor U705 (N_705,In_64,In_212);
and U706 (N_706,In_346,In_284);
or U707 (N_707,In_448,In_70);
and U708 (N_708,In_166,In_277);
or U709 (N_709,In_424,In_461);
nor U710 (N_710,In_497,In_402);
or U711 (N_711,In_305,In_221);
nand U712 (N_712,In_204,In_378);
and U713 (N_713,In_74,In_31);
nand U714 (N_714,In_408,In_104);
xor U715 (N_715,In_292,In_485);
nand U716 (N_716,In_386,In_183);
nor U717 (N_717,In_248,In_284);
and U718 (N_718,In_24,In_403);
and U719 (N_719,In_353,In_367);
nand U720 (N_720,In_228,In_235);
nand U721 (N_721,In_351,In_371);
or U722 (N_722,In_281,In_114);
nor U723 (N_723,In_412,In_147);
xor U724 (N_724,In_288,In_317);
nand U725 (N_725,In_229,In_186);
and U726 (N_726,In_170,In_76);
and U727 (N_727,In_154,In_461);
nand U728 (N_728,In_203,In_458);
nor U729 (N_729,In_475,In_344);
and U730 (N_730,In_197,In_163);
and U731 (N_731,In_251,In_212);
nor U732 (N_732,In_472,In_301);
nand U733 (N_733,In_93,In_319);
nor U734 (N_734,In_275,In_297);
nand U735 (N_735,In_363,In_179);
and U736 (N_736,In_325,In_360);
nor U737 (N_737,In_188,In_269);
nor U738 (N_738,In_436,In_304);
nor U739 (N_739,In_69,In_373);
or U740 (N_740,In_333,In_0);
nand U741 (N_741,In_427,In_356);
or U742 (N_742,In_85,In_117);
xnor U743 (N_743,In_370,In_171);
nand U744 (N_744,In_159,In_134);
nor U745 (N_745,In_239,In_153);
and U746 (N_746,In_327,In_359);
nor U747 (N_747,In_448,In_35);
or U748 (N_748,In_382,In_289);
nand U749 (N_749,In_221,In_427);
and U750 (N_750,In_230,In_23);
nand U751 (N_751,In_231,In_85);
nor U752 (N_752,In_316,In_146);
nand U753 (N_753,In_313,In_461);
or U754 (N_754,In_449,In_351);
and U755 (N_755,In_270,In_432);
nand U756 (N_756,In_244,In_258);
and U757 (N_757,In_461,In_0);
nor U758 (N_758,In_246,In_7);
xor U759 (N_759,In_424,In_13);
nand U760 (N_760,In_27,In_125);
or U761 (N_761,In_395,In_183);
nand U762 (N_762,In_164,In_387);
nand U763 (N_763,In_212,In_153);
or U764 (N_764,In_276,In_463);
and U765 (N_765,In_165,In_253);
nand U766 (N_766,In_303,In_159);
or U767 (N_767,In_108,In_24);
nor U768 (N_768,In_117,In_107);
nand U769 (N_769,In_214,In_145);
xnor U770 (N_770,In_473,In_266);
nand U771 (N_771,In_448,In_438);
nand U772 (N_772,In_258,In_421);
nor U773 (N_773,In_380,In_401);
or U774 (N_774,In_50,In_368);
nand U775 (N_775,In_305,In_462);
or U776 (N_776,In_118,In_391);
or U777 (N_777,In_283,In_211);
nor U778 (N_778,In_158,In_224);
nand U779 (N_779,In_445,In_154);
and U780 (N_780,In_403,In_46);
xnor U781 (N_781,In_32,In_339);
and U782 (N_782,In_366,In_107);
or U783 (N_783,In_325,In_49);
nor U784 (N_784,In_64,In_358);
or U785 (N_785,In_304,In_379);
or U786 (N_786,In_51,In_117);
and U787 (N_787,In_158,In_394);
nor U788 (N_788,In_86,In_56);
and U789 (N_789,In_50,In_404);
nand U790 (N_790,In_159,In_61);
nand U791 (N_791,In_77,In_272);
and U792 (N_792,In_493,In_283);
nor U793 (N_793,In_31,In_450);
and U794 (N_794,In_158,In_175);
nor U795 (N_795,In_165,In_464);
nor U796 (N_796,In_109,In_121);
nand U797 (N_797,In_179,In_469);
and U798 (N_798,In_208,In_99);
and U799 (N_799,In_56,In_469);
nand U800 (N_800,In_318,In_59);
or U801 (N_801,In_139,In_44);
xor U802 (N_802,In_198,In_277);
nor U803 (N_803,In_30,In_101);
or U804 (N_804,In_138,In_21);
xor U805 (N_805,In_278,In_263);
nor U806 (N_806,In_61,In_194);
and U807 (N_807,In_373,In_177);
nor U808 (N_808,In_330,In_285);
nor U809 (N_809,In_27,In_17);
and U810 (N_810,In_293,In_287);
or U811 (N_811,In_197,In_476);
nand U812 (N_812,In_55,In_184);
nand U813 (N_813,In_76,In_150);
and U814 (N_814,In_20,In_87);
and U815 (N_815,In_462,In_87);
and U816 (N_816,In_430,In_33);
or U817 (N_817,In_271,In_98);
or U818 (N_818,In_111,In_494);
and U819 (N_819,In_494,In_428);
nor U820 (N_820,In_265,In_225);
xor U821 (N_821,In_382,In_161);
or U822 (N_822,In_498,In_398);
and U823 (N_823,In_176,In_410);
nor U824 (N_824,In_13,In_155);
nand U825 (N_825,In_294,In_20);
nand U826 (N_826,In_376,In_164);
nor U827 (N_827,In_180,In_443);
nand U828 (N_828,In_487,In_166);
and U829 (N_829,In_49,In_307);
nor U830 (N_830,In_147,In_150);
nor U831 (N_831,In_241,In_336);
and U832 (N_832,In_198,In_278);
or U833 (N_833,In_470,In_239);
xor U834 (N_834,In_460,In_304);
nand U835 (N_835,In_239,In_430);
nor U836 (N_836,In_470,In_57);
nor U837 (N_837,In_274,In_374);
or U838 (N_838,In_479,In_366);
nand U839 (N_839,In_51,In_269);
nor U840 (N_840,In_405,In_435);
and U841 (N_841,In_34,In_393);
and U842 (N_842,In_240,In_14);
nand U843 (N_843,In_420,In_144);
nand U844 (N_844,In_103,In_241);
or U845 (N_845,In_123,In_21);
nand U846 (N_846,In_87,In_406);
or U847 (N_847,In_248,In_152);
xor U848 (N_848,In_110,In_194);
and U849 (N_849,In_135,In_285);
or U850 (N_850,In_461,In_342);
and U851 (N_851,In_354,In_344);
nor U852 (N_852,In_191,In_492);
and U853 (N_853,In_75,In_442);
nand U854 (N_854,In_449,In_304);
nand U855 (N_855,In_112,In_487);
and U856 (N_856,In_182,In_152);
nand U857 (N_857,In_107,In_213);
and U858 (N_858,In_30,In_308);
nand U859 (N_859,In_470,In_2);
nor U860 (N_860,In_428,In_218);
or U861 (N_861,In_418,In_356);
and U862 (N_862,In_212,In_12);
nand U863 (N_863,In_361,In_410);
xnor U864 (N_864,In_473,In_143);
and U865 (N_865,In_201,In_287);
xor U866 (N_866,In_469,In_347);
and U867 (N_867,In_138,In_356);
nand U868 (N_868,In_412,In_405);
and U869 (N_869,In_330,In_84);
nor U870 (N_870,In_350,In_43);
or U871 (N_871,In_390,In_451);
nand U872 (N_872,In_361,In_453);
nand U873 (N_873,In_6,In_131);
nand U874 (N_874,In_98,In_334);
nand U875 (N_875,In_243,In_206);
nand U876 (N_876,In_335,In_13);
nand U877 (N_877,In_105,In_192);
or U878 (N_878,In_325,In_469);
and U879 (N_879,In_66,In_314);
nand U880 (N_880,In_20,In_327);
and U881 (N_881,In_52,In_126);
nor U882 (N_882,In_183,In_51);
nor U883 (N_883,In_0,In_256);
or U884 (N_884,In_2,In_75);
nor U885 (N_885,In_8,In_270);
or U886 (N_886,In_161,In_115);
xor U887 (N_887,In_184,In_37);
or U888 (N_888,In_16,In_217);
or U889 (N_889,In_220,In_178);
and U890 (N_890,In_380,In_129);
nor U891 (N_891,In_72,In_353);
nand U892 (N_892,In_323,In_33);
nor U893 (N_893,In_117,In_340);
or U894 (N_894,In_180,In_257);
xor U895 (N_895,In_230,In_116);
and U896 (N_896,In_408,In_357);
nand U897 (N_897,In_319,In_30);
nor U898 (N_898,In_304,In_319);
nor U899 (N_899,In_244,In_353);
and U900 (N_900,In_224,In_497);
and U901 (N_901,In_405,In_428);
nor U902 (N_902,In_468,In_159);
nor U903 (N_903,In_392,In_480);
or U904 (N_904,In_27,In_432);
nor U905 (N_905,In_2,In_271);
xnor U906 (N_906,In_214,In_243);
nand U907 (N_907,In_436,In_145);
nand U908 (N_908,In_183,In_1);
and U909 (N_909,In_377,In_354);
nor U910 (N_910,In_466,In_308);
and U911 (N_911,In_77,In_93);
nand U912 (N_912,In_37,In_118);
nand U913 (N_913,In_116,In_112);
or U914 (N_914,In_100,In_248);
and U915 (N_915,In_11,In_171);
nand U916 (N_916,In_76,In_262);
or U917 (N_917,In_174,In_182);
and U918 (N_918,In_267,In_147);
nand U919 (N_919,In_117,In_134);
or U920 (N_920,In_408,In_199);
xor U921 (N_921,In_370,In_174);
nand U922 (N_922,In_437,In_172);
and U923 (N_923,In_183,In_439);
nand U924 (N_924,In_280,In_380);
or U925 (N_925,In_483,In_416);
and U926 (N_926,In_304,In_450);
nor U927 (N_927,In_238,In_429);
nand U928 (N_928,In_345,In_376);
or U929 (N_929,In_29,In_419);
nand U930 (N_930,In_439,In_144);
and U931 (N_931,In_468,In_253);
and U932 (N_932,In_159,In_0);
and U933 (N_933,In_364,In_57);
xnor U934 (N_934,In_167,In_68);
nor U935 (N_935,In_216,In_305);
nand U936 (N_936,In_322,In_90);
or U937 (N_937,In_393,In_387);
nand U938 (N_938,In_120,In_472);
and U939 (N_939,In_150,In_75);
nor U940 (N_940,In_59,In_113);
xor U941 (N_941,In_66,In_414);
or U942 (N_942,In_287,In_363);
or U943 (N_943,In_318,In_357);
nor U944 (N_944,In_50,In_410);
or U945 (N_945,In_312,In_145);
and U946 (N_946,In_115,In_478);
and U947 (N_947,In_2,In_258);
nor U948 (N_948,In_90,In_405);
nand U949 (N_949,In_151,In_161);
and U950 (N_950,In_206,In_178);
or U951 (N_951,In_470,In_268);
nor U952 (N_952,In_202,In_167);
nor U953 (N_953,In_328,In_58);
nand U954 (N_954,In_425,In_396);
nor U955 (N_955,In_71,In_388);
and U956 (N_956,In_206,In_449);
or U957 (N_957,In_358,In_399);
nand U958 (N_958,In_328,In_292);
nand U959 (N_959,In_65,In_125);
nor U960 (N_960,In_443,In_59);
xnor U961 (N_961,In_457,In_170);
or U962 (N_962,In_251,In_55);
and U963 (N_963,In_388,In_422);
nor U964 (N_964,In_295,In_26);
nor U965 (N_965,In_63,In_12);
nor U966 (N_966,In_302,In_206);
and U967 (N_967,In_129,In_349);
nand U968 (N_968,In_487,In_420);
and U969 (N_969,In_113,In_249);
and U970 (N_970,In_53,In_123);
nand U971 (N_971,In_44,In_188);
or U972 (N_972,In_84,In_60);
nor U973 (N_973,In_80,In_479);
nor U974 (N_974,In_395,In_406);
nor U975 (N_975,In_155,In_14);
nor U976 (N_976,In_273,In_112);
nand U977 (N_977,In_423,In_372);
nand U978 (N_978,In_112,In_455);
nand U979 (N_979,In_112,In_221);
and U980 (N_980,In_317,In_0);
and U981 (N_981,In_44,In_12);
nand U982 (N_982,In_99,In_479);
or U983 (N_983,In_137,In_439);
or U984 (N_984,In_54,In_135);
nand U985 (N_985,In_30,In_455);
and U986 (N_986,In_360,In_274);
xor U987 (N_987,In_367,In_107);
or U988 (N_988,In_62,In_238);
nor U989 (N_989,In_294,In_449);
or U990 (N_990,In_183,In_121);
and U991 (N_991,In_365,In_70);
or U992 (N_992,In_253,In_201);
and U993 (N_993,In_422,In_2);
nor U994 (N_994,In_462,In_178);
nand U995 (N_995,In_34,In_359);
nand U996 (N_996,In_43,In_76);
nor U997 (N_997,In_412,In_195);
nand U998 (N_998,In_464,In_198);
nand U999 (N_999,In_463,In_20);
nand U1000 (N_1000,N_299,N_32);
nor U1001 (N_1001,N_545,N_276);
xor U1002 (N_1002,N_747,N_919);
nor U1003 (N_1003,N_673,N_870);
nand U1004 (N_1004,N_755,N_185);
nor U1005 (N_1005,N_238,N_865);
nor U1006 (N_1006,N_547,N_611);
or U1007 (N_1007,N_245,N_842);
nor U1008 (N_1008,N_597,N_173);
nand U1009 (N_1009,N_588,N_441);
xnor U1010 (N_1010,N_53,N_168);
nor U1011 (N_1011,N_888,N_419);
nand U1012 (N_1012,N_570,N_620);
nand U1013 (N_1013,N_212,N_183);
nor U1014 (N_1014,N_150,N_180);
or U1015 (N_1015,N_445,N_88);
or U1016 (N_1016,N_830,N_996);
nand U1017 (N_1017,N_681,N_408);
nand U1018 (N_1018,N_801,N_469);
nor U1019 (N_1019,N_78,N_444);
and U1020 (N_1020,N_915,N_770);
nand U1021 (N_1021,N_128,N_568);
nand U1022 (N_1022,N_590,N_468);
nand U1023 (N_1023,N_7,N_343);
xnor U1024 (N_1024,N_694,N_113);
and U1025 (N_1025,N_320,N_159);
and U1026 (N_1026,N_223,N_943);
nand U1027 (N_1027,N_407,N_310);
and U1028 (N_1028,N_574,N_227);
nand U1029 (N_1029,N_354,N_540);
or U1030 (N_1030,N_610,N_867);
nand U1031 (N_1031,N_431,N_455);
nor U1032 (N_1032,N_246,N_237);
and U1033 (N_1033,N_108,N_411);
and U1034 (N_1034,N_330,N_765);
nor U1035 (N_1035,N_432,N_121);
xor U1036 (N_1036,N_255,N_43);
nand U1037 (N_1037,N_756,N_767);
or U1038 (N_1038,N_862,N_93);
nand U1039 (N_1039,N_69,N_195);
nor U1040 (N_1040,N_924,N_460);
and U1041 (N_1041,N_598,N_509);
xor U1042 (N_1042,N_373,N_880);
nor U1043 (N_1043,N_855,N_951);
and U1044 (N_1044,N_548,N_571);
and U1045 (N_1045,N_662,N_562);
nand U1046 (N_1046,N_627,N_278);
nor U1047 (N_1047,N_58,N_512);
xor U1048 (N_1048,N_91,N_231);
nand U1049 (N_1049,N_940,N_931);
or U1050 (N_1050,N_146,N_771);
nand U1051 (N_1051,N_304,N_690);
nand U1052 (N_1052,N_820,N_563);
or U1053 (N_1053,N_504,N_351);
nand U1054 (N_1054,N_17,N_873);
or U1055 (N_1055,N_24,N_942);
nand U1056 (N_1056,N_401,N_267);
nor U1057 (N_1057,N_934,N_955);
or U1058 (N_1058,N_632,N_306);
and U1059 (N_1059,N_470,N_394);
nand U1060 (N_1060,N_658,N_575);
and U1061 (N_1061,N_380,N_983);
and U1062 (N_1062,N_77,N_753);
or U1063 (N_1063,N_702,N_657);
or U1064 (N_1064,N_626,N_19);
nor U1065 (N_1065,N_695,N_560);
nor U1066 (N_1066,N_221,N_669);
and U1067 (N_1067,N_925,N_435);
and U1068 (N_1068,N_250,N_894);
or U1069 (N_1069,N_184,N_135);
and U1070 (N_1070,N_123,N_856);
or U1071 (N_1071,N_112,N_608);
nor U1072 (N_1072,N_181,N_734);
or U1073 (N_1073,N_583,N_663);
nor U1074 (N_1074,N_697,N_833);
or U1075 (N_1075,N_286,N_655);
and U1076 (N_1076,N_349,N_956);
nand U1077 (N_1077,N_61,N_243);
xor U1078 (N_1078,N_328,N_47);
nand U1079 (N_1079,N_13,N_745);
or U1080 (N_1080,N_599,N_258);
nor U1081 (N_1081,N_985,N_100);
nand U1082 (N_1082,N_175,N_740);
or U1083 (N_1083,N_216,N_605);
or U1084 (N_1084,N_288,N_840);
or U1085 (N_1085,N_283,N_201);
nand U1086 (N_1086,N_806,N_21);
or U1087 (N_1087,N_240,N_946);
or U1088 (N_1088,N_927,N_234);
nand U1089 (N_1089,N_777,N_538);
or U1090 (N_1090,N_284,N_155);
nand U1091 (N_1091,N_164,N_696);
or U1092 (N_1092,N_406,N_333);
nand U1093 (N_1093,N_139,N_828);
nor U1094 (N_1094,N_198,N_478);
and U1095 (N_1095,N_327,N_45);
and U1096 (N_1096,N_837,N_645);
and U1097 (N_1097,N_998,N_390);
or U1098 (N_1098,N_481,N_425);
nand U1099 (N_1099,N_322,N_641);
nand U1100 (N_1100,N_975,N_253);
and U1101 (N_1101,N_50,N_60);
nand U1102 (N_1102,N_784,N_5);
xor U1103 (N_1103,N_735,N_868);
or U1104 (N_1104,N_718,N_825);
or U1105 (N_1105,N_324,N_26);
nand U1106 (N_1106,N_79,N_271);
nand U1107 (N_1107,N_810,N_773);
nor U1108 (N_1108,N_875,N_864);
nand U1109 (N_1109,N_721,N_437);
nor U1110 (N_1110,N_300,N_666);
and U1111 (N_1111,N_118,N_623);
xor U1112 (N_1112,N_775,N_652);
xor U1113 (N_1113,N_904,N_171);
and U1114 (N_1114,N_746,N_778);
nor U1115 (N_1115,N_410,N_215);
nor U1116 (N_1116,N_947,N_766);
or U1117 (N_1117,N_485,N_901);
nand U1118 (N_1118,N_821,N_417);
or U1119 (N_1119,N_903,N_169);
or U1120 (N_1120,N_642,N_990);
nand U1121 (N_1121,N_358,N_591);
and U1122 (N_1122,N_664,N_161);
and U1123 (N_1123,N_680,N_687);
nand U1124 (N_1124,N_964,N_369);
or U1125 (N_1125,N_787,N_704);
nor U1126 (N_1126,N_495,N_715);
or U1127 (N_1127,N_22,N_367);
nor U1128 (N_1128,N_222,N_440);
nand U1129 (N_1129,N_365,N_827);
nor U1130 (N_1130,N_206,N_189);
nand U1131 (N_1131,N_675,N_414);
nor U1132 (N_1132,N_792,N_405);
nand U1133 (N_1133,N_854,N_984);
and U1134 (N_1134,N_334,N_534);
and U1135 (N_1135,N_116,N_395);
nor U1136 (N_1136,N_292,N_488);
and U1137 (N_1137,N_689,N_815);
nand U1138 (N_1138,N_883,N_152);
or U1139 (N_1139,N_683,N_637);
and U1140 (N_1140,N_147,N_295);
xor U1141 (N_1141,N_686,N_226);
or U1142 (N_1142,N_758,N_316);
nand U1143 (N_1143,N_779,N_839);
nor U1144 (N_1144,N_363,N_531);
nand U1145 (N_1145,N_433,N_582);
or U1146 (N_1146,N_151,N_41);
nor U1147 (N_1147,N_507,N_217);
nor U1148 (N_1148,N_166,N_404);
and U1149 (N_1149,N_877,N_370);
and U1150 (N_1150,N_525,N_630);
or U1151 (N_1151,N_353,N_550);
or U1152 (N_1152,N_829,N_672);
nor U1153 (N_1153,N_760,N_602);
and U1154 (N_1154,N_502,N_661);
nor U1155 (N_1155,N_907,N_714);
or U1156 (N_1156,N_705,N_336);
or U1157 (N_1157,N_466,N_92);
nand U1158 (N_1158,N_144,N_447);
or U1159 (N_1159,N_517,N_520);
and U1160 (N_1160,N_415,N_515);
nor U1161 (N_1161,N_887,N_224);
nand U1162 (N_1162,N_893,N_257);
and U1163 (N_1163,N_233,N_140);
xnor U1164 (N_1164,N_634,N_852);
nor U1165 (N_1165,N_954,N_667);
nand U1166 (N_1166,N_178,N_961);
xnor U1167 (N_1167,N_581,N_285);
and U1168 (N_1168,N_94,N_134);
or U1169 (N_1169,N_935,N_885);
nor U1170 (N_1170,N_589,N_754);
nand U1171 (N_1171,N_997,N_945);
xor U1172 (N_1172,N_796,N_501);
nor U1173 (N_1173,N_731,N_305);
xor U1174 (N_1174,N_480,N_307);
nand U1175 (N_1175,N_37,N_220);
or U1176 (N_1176,N_219,N_311);
nor U1177 (N_1177,N_120,N_677);
nor U1178 (N_1178,N_302,N_791);
or U1179 (N_1179,N_90,N_699);
or U1180 (N_1180,N_622,N_969);
nand U1181 (N_1181,N_55,N_89);
nand U1182 (N_1182,N_209,N_912);
xnor U1183 (N_1183,N_500,N_229);
or U1184 (N_1184,N_341,N_473);
and U1185 (N_1185,N_160,N_103);
and U1186 (N_1186,N_38,N_863);
or U1187 (N_1187,N_314,N_194);
or U1188 (N_1188,N_162,N_177);
and U1189 (N_1189,N_966,N_429);
nand U1190 (N_1190,N_950,N_54);
nand U1191 (N_1191,N_318,N_321);
and U1192 (N_1192,N_709,N_111);
nor U1193 (N_1193,N_889,N_952);
or U1194 (N_1194,N_392,N_992);
or U1195 (N_1195,N_688,N_190);
and U1196 (N_1196,N_807,N_35);
nand U1197 (N_1197,N_200,N_968);
nor U1198 (N_1198,N_399,N_741);
xnor U1199 (N_1199,N_953,N_649);
nor U1200 (N_1200,N_154,N_930);
xnor U1201 (N_1201,N_595,N_813);
nand U1202 (N_1202,N_671,N_529);
nor U1203 (N_1203,N_388,N_980);
or U1204 (N_1204,N_565,N_542);
xor U1205 (N_1205,N_848,N_838);
and U1206 (N_1206,N_640,N_732);
nand U1207 (N_1207,N_557,N_616);
or U1208 (N_1208,N_274,N_808);
nand U1209 (N_1209,N_567,N_115);
and U1210 (N_1210,N_340,N_498);
nand U1211 (N_1211,N_674,N_174);
nor U1212 (N_1212,N_668,N_654);
xor U1213 (N_1213,N_513,N_514);
and U1214 (N_1214,N_890,N_691);
and U1215 (N_1215,N_277,N_119);
nand U1216 (N_1216,N_923,N_594);
nor U1217 (N_1217,N_149,N_895);
or U1218 (N_1218,N_317,N_851);
or U1219 (N_1219,N_420,N_619);
nand U1220 (N_1220,N_938,N_326);
nand U1221 (N_1221,N_412,N_802);
and U1222 (N_1222,N_249,N_993);
and U1223 (N_1223,N_323,N_772);
or U1224 (N_1224,N_857,N_580);
nor U1225 (N_1225,N_254,N_725);
nor U1226 (N_1226,N_98,N_823);
nor U1227 (N_1227,N_464,N_339);
xor U1228 (N_1228,N_973,N_869);
xor U1229 (N_1229,N_726,N_604);
nand U1230 (N_1230,N_315,N_16);
or U1231 (N_1231,N_376,N_920);
nand U1232 (N_1232,N_561,N_296);
nor U1233 (N_1233,N_700,N_211);
nor U1234 (N_1234,N_126,N_102);
nand U1235 (N_1235,N_66,N_86);
nand U1236 (N_1236,N_493,N_264);
nor U1237 (N_1237,N_426,N_629);
or U1238 (N_1238,N_290,N_107);
and U1239 (N_1239,N_83,N_362);
nor U1240 (N_1240,N_374,N_519);
or U1241 (N_1241,N_761,N_578);
nor U1242 (N_1242,N_818,N_465);
nor U1243 (N_1243,N_165,N_142);
or U1244 (N_1244,N_527,N_449);
and U1245 (N_1245,N_566,N_572);
and U1246 (N_1246,N_87,N_360);
nand U1247 (N_1247,N_532,N_577);
or U1248 (N_1248,N_303,N_609);
nor U1249 (N_1249,N_708,N_651);
or U1250 (N_1250,N_335,N_163);
and U1251 (N_1251,N_462,N_479);
nor U1252 (N_1252,N_443,N_716);
nand U1253 (N_1253,N_280,N_1);
nor U1254 (N_1254,N_707,N_576);
xnor U1255 (N_1255,N_783,N_703);
nor U1256 (N_1256,N_876,N_832);
and U1257 (N_1257,N_505,N_272);
nand U1258 (N_1258,N_615,N_941);
nor U1259 (N_1259,N_881,N_742);
or U1260 (N_1260,N_722,N_592);
nand U1261 (N_1261,N_110,N_95);
nor U1262 (N_1262,N_559,N_467);
nand U1263 (N_1263,N_338,N_396);
xnor U1264 (N_1264,N_970,N_918);
nor U1265 (N_1265,N_387,N_819);
nor U1266 (N_1266,N_247,N_207);
nand U1267 (N_1267,N_23,N_143);
nor U1268 (N_1268,N_988,N_2);
nand U1269 (N_1269,N_319,N_618);
nor U1270 (N_1270,N_347,N_730);
nor U1271 (N_1271,N_82,N_739);
nor U1272 (N_1272,N_603,N_960);
xnor U1273 (N_1273,N_738,N_191);
or U1274 (N_1274,N_477,N_372);
and U1275 (N_1275,N_416,N_70);
or U1276 (N_1276,N_510,N_593);
or U1277 (N_1277,N_73,N_446);
or U1278 (N_1278,N_11,N_29);
nor U1279 (N_1279,N_101,N_685);
xor U1280 (N_1280,N_712,N_452);
nand U1281 (N_1281,N_418,N_643);
and U1282 (N_1282,N_656,N_384);
nor U1283 (N_1283,N_346,N_68);
nand U1284 (N_1284,N_910,N_345);
and U1285 (N_1285,N_210,N_496);
and U1286 (N_1286,N_137,N_724);
and U1287 (N_1287,N_541,N_635);
xnor U1288 (N_1288,N_197,N_921);
nor U1289 (N_1289,N_85,N_293);
or U1290 (N_1290,N_15,N_621);
nand U1291 (N_1291,N_628,N_971);
nor U1292 (N_1292,N_743,N_994);
and U1293 (N_1293,N_483,N_170);
nor U1294 (N_1294,N_400,N_853);
and U1295 (N_1295,N_0,N_794);
nand U1296 (N_1296,N_719,N_403);
nand U1297 (N_1297,N_81,N_138);
and U1298 (N_1298,N_882,N_733);
nand U1299 (N_1299,N_793,N_203);
or U1300 (N_1300,N_650,N_48);
or U1301 (N_1301,N_64,N_804);
and U1302 (N_1302,N_235,N_49);
and U1303 (N_1303,N_554,N_402);
or U1304 (N_1304,N_987,N_965);
nand U1305 (N_1305,N_701,N_74);
nor U1306 (N_1306,N_386,N_551);
xor U1307 (N_1307,N_156,N_494);
or U1308 (N_1308,N_31,N_461);
or U1309 (N_1309,N_125,N_543);
nand U1310 (N_1310,N_585,N_57);
and U1311 (N_1311,N_913,N_356);
nor U1312 (N_1312,N_361,N_944);
xor U1313 (N_1313,N_282,N_273);
or U1314 (N_1314,N_790,N_752);
or U1315 (N_1315,N_814,N_976);
or U1316 (N_1316,N_368,N_244);
or U1317 (N_1317,N_241,N_978);
or U1318 (N_1318,N_167,N_312);
nor U1319 (N_1319,N_36,N_230);
xor U1320 (N_1320,N_906,N_805);
or U1321 (N_1321,N_706,N_744);
or U1322 (N_1322,N_14,N_298);
nor U1323 (N_1323,N_65,N_601);
nand U1324 (N_1324,N_242,N_377);
nor U1325 (N_1325,N_803,N_892);
nor U1326 (N_1326,N_768,N_157);
nand U1327 (N_1327,N_788,N_798);
nand U1328 (N_1328,N_871,N_639);
xnor U1329 (N_1329,N_252,N_558);
or U1330 (N_1330,N_555,N_63);
and U1331 (N_1331,N_59,N_448);
xnor U1332 (N_1332,N_104,N_928);
xor U1333 (N_1333,N_526,N_533);
nor U1334 (N_1334,N_693,N_482);
nor U1335 (N_1335,N_393,N_644);
xor U1336 (N_1336,N_625,N_858);
or U1337 (N_1337,N_192,N_549);
and U1338 (N_1338,N_294,N_332);
or U1339 (N_1339,N_350,N_845);
nor U1340 (N_1340,N_624,N_122);
or U1341 (N_1341,N_51,N_937);
or U1342 (N_1342,N_381,N_759);
xnor U1343 (N_1343,N_442,N_989);
nor U1344 (N_1344,N_397,N_780);
and U1345 (N_1345,N_636,N_325);
nand U1346 (N_1346,N_434,N_430);
nor U1347 (N_1347,N_676,N_389);
nand U1348 (N_1348,N_902,N_967);
nor U1349 (N_1349,N_487,N_9);
nor U1350 (N_1350,N_879,N_471);
and U1351 (N_1351,N_995,N_348);
or U1352 (N_1352,N_186,N_398);
or U1353 (N_1353,N_457,N_522);
or U1354 (N_1354,N_385,N_866);
nand U1355 (N_1355,N_309,N_539);
and U1356 (N_1356,N_962,N_898);
xnor U1357 (N_1357,N_922,N_463);
and U1358 (N_1358,N_188,N_260);
nand U1359 (N_1359,N_109,N_287);
and U1360 (N_1360,N_884,N_492);
and U1361 (N_1361,N_484,N_256);
and U1362 (N_1362,N_56,N_251);
nor U1363 (N_1363,N_281,N_289);
or U1364 (N_1364,N_3,N_979);
or U1365 (N_1365,N_957,N_782);
or U1366 (N_1366,N_800,N_337);
or U1367 (N_1367,N_236,N_556);
or U1368 (N_1368,N_891,N_844);
or U1369 (N_1369,N_489,N_225);
nor U1370 (N_1370,N_516,N_30);
or U1371 (N_1371,N_422,N_552);
nand U1372 (N_1372,N_949,N_698);
nor U1373 (N_1373,N_6,N_817);
xor U1374 (N_1374,N_932,N_886);
or U1375 (N_1375,N_342,N_785);
nor U1376 (N_1376,N_97,N_456);
or U1377 (N_1377,N_76,N_208);
xnor U1378 (N_1378,N_275,N_391);
or U1379 (N_1379,N_750,N_503);
xor U1380 (N_1380,N_917,N_375);
xnor U1381 (N_1381,N_914,N_359);
xor U1382 (N_1382,N_564,N_508);
nor U1383 (N_1383,N_291,N_105);
xnor U1384 (N_1384,N_999,N_33);
and U1385 (N_1385,N_972,N_148);
and U1386 (N_1386,N_261,N_355);
and U1387 (N_1387,N_158,N_799);
nor U1388 (N_1388,N_849,N_737);
xor U1389 (N_1389,N_647,N_682);
nor U1390 (N_1390,N_897,N_214);
and U1391 (N_1391,N_860,N_182);
and U1392 (N_1392,N_20,N_717);
nor U1393 (N_1393,N_262,N_4);
and U1394 (N_1394,N_631,N_723);
and U1395 (N_1395,N_265,N_606);
nand U1396 (N_1396,N_939,N_176);
or U1397 (N_1397,N_313,N_301);
or U1398 (N_1398,N_711,N_269);
or U1399 (N_1399,N_179,N_963);
nor U1400 (N_1400,N_239,N_297);
or U1401 (N_1401,N_809,N_266);
and U1402 (N_1402,N_684,N_789);
and U1403 (N_1403,N_982,N_10);
nand U1404 (N_1404,N_836,N_268);
nand U1405 (N_1405,N_352,N_607);
or U1406 (N_1406,N_44,N_172);
and U1407 (N_1407,N_653,N_232);
nand U1408 (N_1408,N_659,N_308);
or U1409 (N_1409,N_600,N_378);
nand U1410 (N_1410,N_861,N_117);
and U1411 (N_1411,N_553,N_46);
and U1412 (N_1412,N_454,N_846);
and U1413 (N_1413,N_587,N_748);
or U1414 (N_1414,N_841,N_366);
nand U1415 (N_1415,N_364,N_8);
nand U1416 (N_1416,N_991,N_331);
and U1417 (N_1417,N_491,N_911);
or U1418 (N_1418,N_75,N_436);
or U1419 (N_1419,N_874,N_106);
nor U1420 (N_1420,N_133,N_130);
nand U1421 (N_1421,N_579,N_458);
nor U1422 (N_1422,N_728,N_27);
nor U1423 (N_1423,N_424,N_679);
nand U1424 (N_1424,N_569,N_218);
and U1425 (N_1425,N_831,N_763);
nand U1426 (N_1426,N_926,N_129);
nor U1427 (N_1427,N_646,N_213);
xnor U1428 (N_1428,N_136,N_421);
and U1429 (N_1429,N_25,N_909);
and U1430 (N_1430,N_34,N_933);
and U1431 (N_1431,N_506,N_228);
nand U1432 (N_1432,N_713,N_528);
and U1433 (N_1433,N_834,N_499);
nor U1434 (N_1434,N_781,N_535);
and U1435 (N_1435,N_678,N_518);
nand U1436 (N_1436,N_450,N_524);
nor U1437 (N_1437,N_28,N_40);
or U1438 (N_1438,N_259,N_476);
nand U1439 (N_1439,N_382,N_977);
nor U1440 (N_1440,N_80,N_99);
xor U1441 (N_1441,N_586,N_379);
and U1442 (N_1442,N_475,N_371);
nand U1443 (N_1443,N_472,N_497);
and U1444 (N_1444,N_757,N_824);
nor U1445 (N_1445,N_929,N_795);
nand U1446 (N_1446,N_199,N_96);
nor U1447 (N_1447,N_835,N_665);
and U1448 (N_1448,N_537,N_67);
xnor U1449 (N_1449,N_764,N_762);
or U1450 (N_1450,N_132,N_248);
and U1451 (N_1451,N_797,N_145);
xor U1452 (N_1452,N_948,N_986);
nand U1453 (N_1453,N_124,N_279);
nor U1454 (N_1454,N_459,N_329);
nor U1455 (N_1455,N_202,N_383);
xor U1456 (N_1456,N_769,N_523);
and U1457 (N_1457,N_816,N_18);
or U1458 (N_1458,N_729,N_521);
xor U1459 (N_1459,N_114,N_899);
or U1460 (N_1460,N_613,N_859);
nor U1461 (N_1461,N_614,N_905);
nand U1462 (N_1462,N_596,N_52);
or U1463 (N_1463,N_900,N_638);
nand U1464 (N_1464,N_878,N_413);
and U1465 (N_1465,N_749,N_826);
nand U1466 (N_1466,N_774,N_617);
nand U1467 (N_1467,N_720,N_822);
nand U1468 (N_1468,N_62,N_959);
nor U1469 (N_1469,N_205,N_544);
nand U1470 (N_1470,N_270,N_71);
and U1471 (N_1471,N_12,N_847);
and U1472 (N_1472,N_439,N_127);
and U1473 (N_1473,N_786,N_428);
nand U1474 (N_1474,N_670,N_423);
and U1475 (N_1475,N_196,N_981);
nand U1476 (N_1476,N_736,N_850);
nor U1477 (N_1477,N_427,N_263);
or U1478 (N_1478,N_39,N_958);
and U1479 (N_1479,N_872,N_490);
nor U1480 (N_1480,N_936,N_153);
and U1481 (N_1481,N_344,N_974);
xnor U1482 (N_1482,N_710,N_511);
and U1483 (N_1483,N_474,N_573);
or U1484 (N_1484,N_751,N_584);
nor U1485 (N_1485,N_811,N_84);
nor U1486 (N_1486,N_727,N_486);
nor U1487 (N_1487,N_916,N_42);
xor U1488 (N_1488,N_546,N_692);
and U1489 (N_1489,N_187,N_451);
or U1490 (N_1490,N_776,N_633);
nor U1491 (N_1491,N_843,N_812);
xor U1492 (N_1492,N_72,N_612);
or U1493 (N_1493,N_536,N_453);
nor U1494 (N_1494,N_357,N_660);
nand U1495 (N_1495,N_908,N_131);
nor U1496 (N_1496,N_530,N_896);
xnor U1497 (N_1497,N_648,N_204);
nor U1498 (N_1498,N_438,N_193);
nand U1499 (N_1499,N_409,N_141);
or U1500 (N_1500,N_575,N_985);
nor U1501 (N_1501,N_672,N_781);
nor U1502 (N_1502,N_884,N_404);
and U1503 (N_1503,N_255,N_176);
and U1504 (N_1504,N_755,N_827);
nand U1505 (N_1505,N_257,N_425);
nand U1506 (N_1506,N_930,N_151);
or U1507 (N_1507,N_884,N_834);
and U1508 (N_1508,N_181,N_942);
nand U1509 (N_1509,N_625,N_712);
and U1510 (N_1510,N_538,N_818);
nor U1511 (N_1511,N_950,N_428);
nor U1512 (N_1512,N_596,N_133);
or U1513 (N_1513,N_468,N_419);
nor U1514 (N_1514,N_176,N_333);
and U1515 (N_1515,N_405,N_180);
nand U1516 (N_1516,N_481,N_141);
or U1517 (N_1517,N_281,N_203);
nand U1518 (N_1518,N_536,N_274);
or U1519 (N_1519,N_538,N_634);
xor U1520 (N_1520,N_390,N_979);
and U1521 (N_1521,N_85,N_372);
nor U1522 (N_1522,N_207,N_527);
and U1523 (N_1523,N_301,N_277);
or U1524 (N_1524,N_386,N_130);
nor U1525 (N_1525,N_776,N_248);
nand U1526 (N_1526,N_747,N_262);
or U1527 (N_1527,N_169,N_112);
nor U1528 (N_1528,N_608,N_246);
nand U1529 (N_1529,N_622,N_44);
or U1530 (N_1530,N_740,N_566);
and U1531 (N_1531,N_247,N_841);
or U1532 (N_1532,N_900,N_77);
nand U1533 (N_1533,N_139,N_572);
and U1534 (N_1534,N_508,N_151);
xor U1535 (N_1535,N_657,N_881);
nand U1536 (N_1536,N_847,N_910);
xnor U1537 (N_1537,N_713,N_649);
and U1538 (N_1538,N_22,N_655);
nor U1539 (N_1539,N_922,N_661);
and U1540 (N_1540,N_355,N_131);
nor U1541 (N_1541,N_802,N_780);
and U1542 (N_1542,N_267,N_632);
or U1543 (N_1543,N_256,N_440);
nand U1544 (N_1544,N_765,N_184);
or U1545 (N_1545,N_280,N_437);
nand U1546 (N_1546,N_485,N_465);
nor U1547 (N_1547,N_700,N_62);
xnor U1548 (N_1548,N_661,N_429);
nor U1549 (N_1549,N_584,N_826);
or U1550 (N_1550,N_645,N_164);
nand U1551 (N_1551,N_784,N_590);
and U1552 (N_1552,N_879,N_758);
or U1553 (N_1553,N_297,N_424);
and U1554 (N_1554,N_531,N_823);
nor U1555 (N_1555,N_333,N_820);
nand U1556 (N_1556,N_560,N_104);
and U1557 (N_1557,N_17,N_439);
nand U1558 (N_1558,N_377,N_711);
or U1559 (N_1559,N_40,N_259);
nor U1560 (N_1560,N_611,N_847);
or U1561 (N_1561,N_148,N_783);
and U1562 (N_1562,N_235,N_69);
nor U1563 (N_1563,N_667,N_20);
and U1564 (N_1564,N_630,N_645);
nand U1565 (N_1565,N_984,N_880);
nand U1566 (N_1566,N_41,N_357);
nor U1567 (N_1567,N_500,N_14);
nand U1568 (N_1568,N_647,N_412);
nand U1569 (N_1569,N_833,N_278);
xnor U1570 (N_1570,N_642,N_358);
and U1571 (N_1571,N_348,N_972);
or U1572 (N_1572,N_405,N_298);
and U1573 (N_1573,N_276,N_530);
nor U1574 (N_1574,N_402,N_678);
nor U1575 (N_1575,N_124,N_539);
or U1576 (N_1576,N_662,N_693);
and U1577 (N_1577,N_293,N_594);
and U1578 (N_1578,N_715,N_868);
nand U1579 (N_1579,N_989,N_262);
nor U1580 (N_1580,N_644,N_188);
nor U1581 (N_1581,N_286,N_358);
nand U1582 (N_1582,N_55,N_980);
or U1583 (N_1583,N_366,N_971);
or U1584 (N_1584,N_400,N_739);
and U1585 (N_1585,N_821,N_603);
or U1586 (N_1586,N_856,N_282);
nand U1587 (N_1587,N_269,N_330);
xor U1588 (N_1588,N_461,N_590);
nor U1589 (N_1589,N_315,N_671);
nand U1590 (N_1590,N_977,N_628);
and U1591 (N_1591,N_919,N_164);
nor U1592 (N_1592,N_60,N_353);
xnor U1593 (N_1593,N_556,N_225);
nand U1594 (N_1594,N_911,N_634);
or U1595 (N_1595,N_479,N_32);
nor U1596 (N_1596,N_767,N_528);
nor U1597 (N_1597,N_607,N_879);
nor U1598 (N_1598,N_357,N_399);
nor U1599 (N_1599,N_117,N_362);
or U1600 (N_1600,N_130,N_708);
or U1601 (N_1601,N_662,N_61);
xnor U1602 (N_1602,N_541,N_803);
and U1603 (N_1603,N_588,N_309);
nand U1604 (N_1604,N_717,N_151);
nor U1605 (N_1605,N_252,N_739);
xnor U1606 (N_1606,N_815,N_999);
or U1607 (N_1607,N_34,N_84);
xnor U1608 (N_1608,N_974,N_168);
and U1609 (N_1609,N_610,N_98);
or U1610 (N_1610,N_488,N_297);
or U1611 (N_1611,N_66,N_961);
and U1612 (N_1612,N_780,N_476);
and U1613 (N_1613,N_530,N_841);
or U1614 (N_1614,N_663,N_158);
nand U1615 (N_1615,N_208,N_810);
nor U1616 (N_1616,N_558,N_967);
xnor U1617 (N_1617,N_965,N_671);
or U1618 (N_1618,N_159,N_181);
nand U1619 (N_1619,N_796,N_672);
nor U1620 (N_1620,N_694,N_376);
xor U1621 (N_1621,N_362,N_34);
or U1622 (N_1622,N_398,N_389);
nor U1623 (N_1623,N_703,N_857);
nand U1624 (N_1624,N_265,N_288);
xnor U1625 (N_1625,N_820,N_957);
or U1626 (N_1626,N_673,N_24);
xor U1627 (N_1627,N_728,N_20);
or U1628 (N_1628,N_559,N_802);
xnor U1629 (N_1629,N_886,N_896);
nand U1630 (N_1630,N_94,N_32);
and U1631 (N_1631,N_291,N_67);
xor U1632 (N_1632,N_585,N_130);
nand U1633 (N_1633,N_54,N_145);
and U1634 (N_1634,N_690,N_343);
nor U1635 (N_1635,N_361,N_766);
nor U1636 (N_1636,N_725,N_157);
or U1637 (N_1637,N_730,N_414);
nand U1638 (N_1638,N_21,N_580);
nor U1639 (N_1639,N_109,N_100);
and U1640 (N_1640,N_876,N_325);
xor U1641 (N_1641,N_505,N_292);
or U1642 (N_1642,N_746,N_484);
and U1643 (N_1643,N_226,N_492);
nor U1644 (N_1644,N_495,N_986);
xnor U1645 (N_1645,N_338,N_317);
nand U1646 (N_1646,N_956,N_319);
or U1647 (N_1647,N_731,N_93);
or U1648 (N_1648,N_976,N_712);
and U1649 (N_1649,N_9,N_223);
nor U1650 (N_1650,N_339,N_986);
nand U1651 (N_1651,N_304,N_626);
nor U1652 (N_1652,N_636,N_830);
or U1653 (N_1653,N_964,N_397);
nand U1654 (N_1654,N_936,N_73);
nor U1655 (N_1655,N_389,N_559);
nand U1656 (N_1656,N_414,N_715);
nand U1657 (N_1657,N_281,N_46);
and U1658 (N_1658,N_265,N_541);
nand U1659 (N_1659,N_392,N_933);
or U1660 (N_1660,N_792,N_972);
and U1661 (N_1661,N_127,N_106);
nand U1662 (N_1662,N_42,N_607);
or U1663 (N_1663,N_167,N_318);
and U1664 (N_1664,N_758,N_933);
nand U1665 (N_1665,N_411,N_473);
xnor U1666 (N_1666,N_637,N_179);
and U1667 (N_1667,N_195,N_425);
nor U1668 (N_1668,N_800,N_931);
or U1669 (N_1669,N_633,N_22);
or U1670 (N_1670,N_626,N_878);
nand U1671 (N_1671,N_930,N_16);
and U1672 (N_1672,N_17,N_714);
and U1673 (N_1673,N_328,N_915);
and U1674 (N_1674,N_119,N_683);
and U1675 (N_1675,N_399,N_57);
and U1676 (N_1676,N_982,N_576);
nor U1677 (N_1677,N_301,N_860);
nor U1678 (N_1678,N_593,N_8);
xor U1679 (N_1679,N_69,N_164);
xor U1680 (N_1680,N_111,N_162);
or U1681 (N_1681,N_660,N_769);
nand U1682 (N_1682,N_73,N_329);
xor U1683 (N_1683,N_295,N_893);
nor U1684 (N_1684,N_73,N_393);
nand U1685 (N_1685,N_761,N_289);
nand U1686 (N_1686,N_626,N_288);
and U1687 (N_1687,N_832,N_105);
or U1688 (N_1688,N_765,N_743);
nand U1689 (N_1689,N_392,N_454);
or U1690 (N_1690,N_824,N_336);
nand U1691 (N_1691,N_78,N_559);
nor U1692 (N_1692,N_259,N_925);
xnor U1693 (N_1693,N_32,N_454);
and U1694 (N_1694,N_750,N_786);
and U1695 (N_1695,N_690,N_437);
or U1696 (N_1696,N_98,N_781);
and U1697 (N_1697,N_699,N_943);
and U1698 (N_1698,N_686,N_390);
nand U1699 (N_1699,N_427,N_640);
or U1700 (N_1700,N_669,N_93);
nor U1701 (N_1701,N_546,N_54);
or U1702 (N_1702,N_5,N_531);
nor U1703 (N_1703,N_845,N_952);
nor U1704 (N_1704,N_780,N_924);
or U1705 (N_1705,N_464,N_250);
xor U1706 (N_1706,N_842,N_523);
nand U1707 (N_1707,N_128,N_461);
or U1708 (N_1708,N_253,N_556);
or U1709 (N_1709,N_183,N_951);
and U1710 (N_1710,N_58,N_232);
and U1711 (N_1711,N_740,N_819);
and U1712 (N_1712,N_182,N_219);
or U1713 (N_1713,N_420,N_691);
or U1714 (N_1714,N_142,N_632);
or U1715 (N_1715,N_284,N_256);
and U1716 (N_1716,N_618,N_385);
xnor U1717 (N_1717,N_640,N_475);
and U1718 (N_1718,N_925,N_13);
xor U1719 (N_1719,N_522,N_362);
nor U1720 (N_1720,N_834,N_964);
or U1721 (N_1721,N_683,N_561);
nand U1722 (N_1722,N_61,N_676);
nor U1723 (N_1723,N_460,N_469);
nand U1724 (N_1724,N_503,N_574);
nor U1725 (N_1725,N_568,N_660);
nand U1726 (N_1726,N_88,N_316);
nor U1727 (N_1727,N_611,N_860);
nor U1728 (N_1728,N_324,N_50);
nand U1729 (N_1729,N_288,N_270);
nor U1730 (N_1730,N_205,N_677);
nand U1731 (N_1731,N_26,N_58);
nand U1732 (N_1732,N_964,N_615);
xnor U1733 (N_1733,N_297,N_277);
nand U1734 (N_1734,N_991,N_747);
and U1735 (N_1735,N_590,N_178);
and U1736 (N_1736,N_699,N_401);
and U1737 (N_1737,N_346,N_948);
nand U1738 (N_1738,N_31,N_149);
nor U1739 (N_1739,N_762,N_883);
or U1740 (N_1740,N_818,N_977);
nor U1741 (N_1741,N_909,N_446);
or U1742 (N_1742,N_817,N_10);
and U1743 (N_1743,N_480,N_639);
and U1744 (N_1744,N_209,N_42);
nor U1745 (N_1745,N_320,N_6);
nor U1746 (N_1746,N_430,N_812);
nor U1747 (N_1747,N_861,N_926);
nor U1748 (N_1748,N_691,N_901);
nand U1749 (N_1749,N_982,N_63);
or U1750 (N_1750,N_47,N_193);
and U1751 (N_1751,N_15,N_265);
nand U1752 (N_1752,N_122,N_217);
nand U1753 (N_1753,N_124,N_875);
nand U1754 (N_1754,N_292,N_269);
nor U1755 (N_1755,N_764,N_635);
or U1756 (N_1756,N_661,N_281);
or U1757 (N_1757,N_983,N_313);
xnor U1758 (N_1758,N_198,N_821);
nand U1759 (N_1759,N_363,N_453);
nand U1760 (N_1760,N_505,N_217);
nor U1761 (N_1761,N_565,N_804);
nor U1762 (N_1762,N_384,N_220);
xor U1763 (N_1763,N_443,N_593);
or U1764 (N_1764,N_426,N_686);
and U1765 (N_1765,N_863,N_325);
xor U1766 (N_1766,N_582,N_490);
nor U1767 (N_1767,N_763,N_534);
nor U1768 (N_1768,N_687,N_748);
or U1769 (N_1769,N_643,N_789);
or U1770 (N_1770,N_320,N_740);
nand U1771 (N_1771,N_112,N_735);
and U1772 (N_1772,N_254,N_589);
or U1773 (N_1773,N_106,N_267);
nor U1774 (N_1774,N_370,N_606);
nor U1775 (N_1775,N_439,N_235);
or U1776 (N_1776,N_648,N_170);
nand U1777 (N_1777,N_895,N_177);
nand U1778 (N_1778,N_840,N_121);
and U1779 (N_1779,N_687,N_946);
or U1780 (N_1780,N_355,N_141);
and U1781 (N_1781,N_602,N_865);
or U1782 (N_1782,N_362,N_703);
xnor U1783 (N_1783,N_645,N_708);
nand U1784 (N_1784,N_547,N_485);
and U1785 (N_1785,N_769,N_702);
and U1786 (N_1786,N_535,N_735);
or U1787 (N_1787,N_293,N_558);
nor U1788 (N_1788,N_576,N_809);
nor U1789 (N_1789,N_76,N_260);
nand U1790 (N_1790,N_10,N_116);
or U1791 (N_1791,N_16,N_64);
and U1792 (N_1792,N_982,N_850);
or U1793 (N_1793,N_413,N_275);
xnor U1794 (N_1794,N_437,N_317);
and U1795 (N_1795,N_17,N_973);
and U1796 (N_1796,N_338,N_42);
and U1797 (N_1797,N_84,N_71);
or U1798 (N_1798,N_900,N_551);
or U1799 (N_1799,N_425,N_4);
and U1800 (N_1800,N_536,N_510);
xnor U1801 (N_1801,N_474,N_95);
or U1802 (N_1802,N_521,N_882);
nor U1803 (N_1803,N_767,N_770);
and U1804 (N_1804,N_245,N_458);
nand U1805 (N_1805,N_542,N_514);
nand U1806 (N_1806,N_271,N_637);
nand U1807 (N_1807,N_342,N_672);
and U1808 (N_1808,N_507,N_37);
xor U1809 (N_1809,N_136,N_915);
and U1810 (N_1810,N_824,N_212);
nand U1811 (N_1811,N_265,N_760);
and U1812 (N_1812,N_879,N_394);
nor U1813 (N_1813,N_124,N_270);
xnor U1814 (N_1814,N_762,N_322);
nor U1815 (N_1815,N_671,N_947);
and U1816 (N_1816,N_669,N_69);
nor U1817 (N_1817,N_106,N_27);
and U1818 (N_1818,N_743,N_717);
nand U1819 (N_1819,N_127,N_368);
and U1820 (N_1820,N_600,N_672);
nor U1821 (N_1821,N_604,N_392);
nand U1822 (N_1822,N_476,N_490);
and U1823 (N_1823,N_793,N_194);
nor U1824 (N_1824,N_979,N_927);
or U1825 (N_1825,N_208,N_343);
or U1826 (N_1826,N_559,N_932);
and U1827 (N_1827,N_497,N_815);
nand U1828 (N_1828,N_961,N_394);
nor U1829 (N_1829,N_750,N_541);
nor U1830 (N_1830,N_496,N_50);
nor U1831 (N_1831,N_554,N_685);
or U1832 (N_1832,N_517,N_879);
nand U1833 (N_1833,N_743,N_312);
and U1834 (N_1834,N_947,N_97);
and U1835 (N_1835,N_581,N_256);
or U1836 (N_1836,N_396,N_114);
or U1837 (N_1837,N_555,N_602);
or U1838 (N_1838,N_340,N_485);
xor U1839 (N_1839,N_640,N_464);
and U1840 (N_1840,N_644,N_360);
nand U1841 (N_1841,N_907,N_237);
or U1842 (N_1842,N_698,N_980);
or U1843 (N_1843,N_219,N_262);
or U1844 (N_1844,N_180,N_752);
nand U1845 (N_1845,N_177,N_967);
nand U1846 (N_1846,N_228,N_387);
and U1847 (N_1847,N_709,N_839);
nand U1848 (N_1848,N_969,N_638);
nand U1849 (N_1849,N_939,N_767);
or U1850 (N_1850,N_371,N_206);
or U1851 (N_1851,N_195,N_468);
nand U1852 (N_1852,N_389,N_34);
and U1853 (N_1853,N_308,N_319);
and U1854 (N_1854,N_656,N_702);
and U1855 (N_1855,N_368,N_148);
xor U1856 (N_1856,N_754,N_845);
and U1857 (N_1857,N_82,N_149);
nand U1858 (N_1858,N_948,N_229);
nand U1859 (N_1859,N_240,N_791);
nor U1860 (N_1860,N_687,N_843);
and U1861 (N_1861,N_412,N_48);
and U1862 (N_1862,N_747,N_749);
and U1863 (N_1863,N_653,N_217);
and U1864 (N_1864,N_313,N_235);
nand U1865 (N_1865,N_609,N_43);
nand U1866 (N_1866,N_57,N_188);
and U1867 (N_1867,N_602,N_279);
and U1868 (N_1868,N_576,N_371);
and U1869 (N_1869,N_839,N_954);
or U1870 (N_1870,N_602,N_52);
and U1871 (N_1871,N_676,N_574);
xor U1872 (N_1872,N_877,N_414);
and U1873 (N_1873,N_782,N_323);
and U1874 (N_1874,N_285,N_257);
nand U1875 (N_1875,N_136,N_274);
and U1876 (N_1876,N_675,N_496);
or U1877 (N_1877,N_617,N_341);
nor U1878 (N_1878,N_103,N_986);
xor U1879 (N_1879,N_564,N_791);
and U1880 (N_1880,N_604,N_949);
or U1881 (N_1881,N_21,N_574);
xor U1882 (N_1882,N_199,N_291);
or U1883 (N_1883,N_513,N_630);
nor U1884 (N_1884,N_165,N_389);
nor U1885 (N_1885,N_193,N_768);
or U1886 (N_1886,N_713,N_410);
or U1887 (N_1887,N_271,N_830);
or U1888 (N_1888,N_713,N_706);
nand U1889 (N_1889,N_93,N_205);
nand U1890 (N_1890,N_153,N_19);
xor U1891 (N_1891,N_992,N_100);
nand U1892 (N_1892,N_65,N_228);
or U1893 (N_1893,N_782,N_332);
and U1894 (N_1894,N_452,N_656);
nor U1895 (N_1895,N_707,N_657);
nand U1896 (N_1896,N_676,N_917);
nand U1897 (N_1897,N_910,N_309);
nand U1898 (N_1898,N_411,N_620);
nand U1899 (N_1899,N_898,N_857);
and U1900 (N_1900,N_266,N_319);
nor U1901 (N_1901,N_668,N_328);
nor U1902 (N_1902,N_76,N_810);
nand U1903 (N_1903,N_999,N_136);
nand U1904 (N_1904,N_665,N_185);
or U1905 (N_1905,N_567,N_908);
or U1906 (N_1906,N_898,N_164);
nor U1907 (N_1907,N_460,N_235);
xor U1908 (N_1908,N_209,N_190);
xnor U1909 (N_1909,N_673,N_406);
nor U1910 (N_1910,N_961,N_25);
nor U1911 (N_1911,N_719,N_836);
nand U1912 (N_1912,N_216,N_946);
xnor U1913 (N_1913,N_989,N_309);
and U1914 (N_1914,N_305,N_13);
and U1915 (N_1915,N_485,N_687);
nand U1916 (N_1916,N_825,N_403);
nand U1917 (N_1917,N_323,N_451);
nand U1918 (N_1918,N_627,N_568);
nor U1919 (N_1919,N_849,N_779);
nand U1920 (N_1920,N_208,N_146);
nor U1921 (N_1921,N_137,N_242);
or U1922 (N_1922,N_439,N_993);
nor U1923 (N_1923,N_307,N_16);
nor U1924 (N_1924,N_306,N_500);
and U1925 (N_1925,N_132,N_329);
or U1926 (N_1926,N_816,N_308);
or U1927 (N_1927,N_896,N_263);
nor U1928 (N_1928,N_524,N_609);
and U1929 (N_1929,N_251,N_276);
nand U1930 (N_1930,N_172,N_821);
nand U1931 (N_1931,N_503,N_231);
and U1932 (N_1932,N_196,N_895);
nor U1933 (N_1933,N_234,N_178);
nand U1934 (N_1934,N_419,N_4);
nand U1935 (N_1935,N_673,N_468);
nor U1936 (N_1936,N_7,N_486);
or U1937 (N_1937,N_654,N_542);
or U1938 (N_1938,N_736,N_763);
nand U1939 (N_1939,N_876,N_234);
and U1940 (N_1940,N_949,N_121);
and U1941 (N_1941,N_858,N_594);
and U1942 (N_1942,N_408,N_104);
xor U1943 (N_1943,N_218,N_773);
nand U1944 (N_1944,N_198,N_305);
and U1945 (N_1945,N_996,N_919);
and U1946 (N_1946,N_574,N_859);
or U1947 (N_1947,N_817,N_695);
nor U1948 (N_1948,N_530,N_984);
xnor U1949 (N_1949,N_90,N_802);
xnor U1950 (N_1950,N_411,N_409);
and U1951 (N_1951,N_19,N_387);
nand U1952 (N_1952,N_922,N_946);
nand U1953 (N_1953,N_161,N_139);
nor U1954 (N_1954,N_333,N_750);
nand U1955 (N_1955,N_508,N_943);
nand U1956 (N_1956,N_570,N_902);
nor U1957 (N_1957,N_30,N_87);
and U1958 (N_1958,N_576,N_92);
nand U1959 (N_1959,N_832,N_135);
or U1960 (N_1960,N_47,N_494);
and U1961 (N_1961,N_27,N_593);
and U1962 (N_1962,N_962,N_696);
nor U1963 (N_1963,N_202,N_881);
and U1964 (N_1964,N_90,N_327);
nand U1965 (N_1965,N_728,N_876);
nor U1966 (N_1966,N_166,N_653);
nor U1967 (N_1967,N_418,N_508);
or U1968 (N_1968,N_37,N_760);
xor U1969 (N_1969,N_590,N_803);
or U1970 (N_1970,N_759,N_168);
or U1971 (N_1971,N_38,N_87);
nand U1972 (N_1972,N_851,N_627);
and U1973 (N_1973,N_211,N_137);
nor U1974 (N_1974,N_31,N_278);
xor U1975 (N_1975,N_433,N_548);
nor U1976 (N_1976,N_334,N_464);
or U1977 (N_1977,N_96,N_502);
nor U1978 (N_1978,N_238,N_799);
or U1979 (N_1979,N_722,N_718);
and U1980 (N_1980,N_322,N_442);
or U1981 (N_1981,N_55,N_436);
or U1982 (N_1982,N_631,N_202);
and U1983 (N_1983,N_761,N_523);
nor U1984 (N_1984,N_903,N_577);
nor U1985 (N_1985,N_415,N_528);
or U1986 (N_1986,N_85,N_369);
nand U1987 (N_1987,N_882,N_299);
nand U1988 (N_1988,N_494,N_941);
nor U1989 (N_1989,N_603,N_902);
or U1990 (N_1990,N_214,N_793);
nor U1991 (N_1991,N_718,N_147);
nor U1992 (N_1992,N_329,N_251);
xnor U1993 (N_1993,N_177,N_730);
and U1994 (N_1994,N_837,N_259);
and U1995 (N_1995,N_715,N_278);
nor U1996 (N_1996,N_345,N_172);
or U1997 (N_1997,N_235,N_738);
and U1998 (N_1998,N_318,N_951);
xor U1999 (N_1999,N_152,N_32);
xor U2000 (N_2000,N_1452,N_1767);
nand U2001 (N_2001,N_1589,N_1210);
nor U2002 (N_2002,N_1110,N_1167);
and U2003 (N_2003,N_1851,N_1896);
nand U2004 (N_2004,N_1638,N_1438);
and U2005 (N_2005,N_1398,N_1789);
or U2006 (N_2006,N_1235,N_1935);
and U2007 (N_2007,N_1250,N_1297);
or U2008 (N_2008,N_1051,N_1525);
and U2009 (N_2009,N_1987,N_1082);
xor U2010 (N_2010,N_1641,N_1468);
or U2011 (N_2011,N_1678,N_1300);
and U2012 (N_2012,N_1883,N_1008);
xnor U2013 (N_2013,N_1724,N_1961);
nand U2014 (N_2014,N_1196,N_1958);
and U2015 (N_2015,N_1255,N_1295);
and U2016 (N_2016,N_1891,N_1424);
and U2017 (N_2017,N_1249,N_1937);
nand U2018 (N_2018,N_1572,N_1323);
nor U2019 (N_2019,N_1462,N_1842);
or U2020 (N_2020,N_1565,N_1666);
nand U2021 (N_2021,N_1338,N_1748);
xor U2022 (N_2022,N_1366,N_1068);
or U2023 (N_2023,N_1928,N_1893);
and U2024 (N_2024,N_1882,N_1072);
or U2025 (N_2025,N_1770,N_1529);
xor U2026 (N_2026,N_1546,N_1077);
nand U2027 (N_2027,N_1561,N_1618);
xor U2028 (N_2028,N_1450,N_1147);
and U2029 (N_2029,N_1417,N_1706);
nand U2030 (N_2030,N_1263,N_1870);
or U2031 (N_2031,N_1444,N_1014);
xor U2032 (N_2032,N_1824,N_1888);
nor U2033 (N_2033,N_1391,N_1363);
nor U2034 (N_2034,N_1804,N_1091);
nand U2035 (N_2035,N_1631,N_1408);
nand U2036 (N_2036,N_1203,N_1562);
xor U2037 (N_2037,N_1066,N_1412);
or U2038 (N_2038,N_1244,N_1763);
nor U2039 (N_2039,N_1791,N_1909);
and U2040 (N_2040,N_1624,N_1907);
nor U2041 (N_2041,N_1714,N_1950);
nor U2042 (N_2042,N_1115,N_1173);
and U2043 (N_2043,N_1028,N_1459);
or U2044 (N_2044,N_1164,N_1880);
or U2045 (N_2045,N_1220,N_1813);
nand U2046 (N_2046,N_1350,N_1771);
or U2047 (N_2047,N_1858,N_1513);
or U2048 (N_2048,N_1689,N_1116);
xor U2049 (N_2049,N_1522,N_1319);
or U2050 (N_2050,N_1490,N_1687);
and U2051 (N_2051,N_1286,N_1154);
nand U2052 (N_2052,N_1537,N_1416);
nand U2053 (N_2053,N_1247,N_1948);
and U2054 (N_2054,N_1698,N_1699);
nand U2055 (N_2055,N_1984,N_1818);
xnor U2056 (N_2056,N_1360,N_1336);
or U2057 (N_2057,N_1700,N_1908);
or U2058 (N_2058,N_1314,N_1060);
xnor U2059 (N_2059,N_1308,N_1176);
and U2060 (N_2060,N_1169,N_1180);
xor U2061 (N_2061,N_1160,N_1540);
xor U2062 (N_2062,N_1711,N_1633);
or U2063 (N_2063,N_1015,N_1113);
nand U2064 (N_2064,N_1423,N_1253);
nor U2065 (N_2065,N_1185,N_1703);
and U2066 (N_2066,N_1017,N_1020);
nor U2067 (N_2067,N_1402,N_1753);
xnor U2068 (N_2068,N_1397,N_1257);
nor U2069 (N_2069,N_1647,N_1362);
xnor U2070 (N_2070,N_1534,N_1520);
and U2071 (N_2071,N_1476,N_1707);
or U2072 (N_2072,N_1079,N_1764);
or U2073 (N_2073,N_1282,N_1493);
nand U2074 (N_2074,N_1514,N_1799);
nand U2075 (N_2075,N_1299,N_1857);
and U2076 (N_2076,N_1309,N_1337);
and U2077 (N_2077,N_1980,N_1849);
xnor U2078 (N_2078,N_1903,N_1382);
or U2079 (N_2079,N_1663,N_1577);
and U2080 (N_2080,N_1328,N_1347);
nand U2081 (N_2081,N_1936,N_1492);
xnor U2082 (N_2082,N_1171,N_1820);
and U2083 (N_2083,N_1766,N_1061);
nor U2084 (N_2084,N_1685,N_1795);
nor U2085 (N_2085,N_1786,N_1458);
and U2086 (N_2086,N_1701,N_1652);
or U2087 (N_2087,N_1730,N_1104);
xor U2088 (N_2088,N_1127,N_1548);
or U2089 (N_2089,N_1415,N_1528);
nand U2090 (N_2090,N_1039,N_1358);
nor U2091 (N_2091,N_1944,N_1611);
nor U2092 (N_2092,N_1425,N_1453);
nand U2093 (N_2093,N_1403,N_1228);
nand U2094 (N_2094,N_1670,N_1628);
or U2095 (N_2095,N_1926,N_1022);
nand U2096 (N_2096,N_1165,N_1946);
nand U2097 (N_2097,N_1722,N_1088);
nor U2098 (N_2098,N_1034,N_1930);
or U2099 (N_2099,N_1662,N_1951);
or U2100 (N_2100,N_1594,N_1479);
or U2101 (N_2101,N_1997,N_1801);
nor U2102 (N_2102,N_1217,N_1457);
or U2103 (N_2103,N_1590,N_1636);
and U2104 (N_2104,N_1311,N_1828);
and U2105 (N_2105,N_1592,N_1863);
nand U2106 (N_2106,N_1427,N_1233);
nor U2107 (N_2107,N_1218,N_1639);
nor U2108 (N_2108,N_1879,N_1083);
and U2109 (N_2109,N_1443,N_1952);
nand U2110 (N_2110,N_1899,N_1616);
or U2111 (N_2111,N_1836,N_1188);
xor U2112 (N_2112,N_1288,N_1107);
nor U2113 (N_2113,N_1274,N_1601);
xor U2114 (N_2114,N_1277,N_1759);
nor U2115 (N_2115,N_1121,N_1195);
nand U2116 (N_2116,N_1062,N_1105);
xor U2117 (N_2117,N_1686,N_1809);
and U2118 (N_2118,N_1521,N_1779);
and U2119 (N_2119,N_1845,N_1569);
nand U2120 (N_2120,N_1152,N_1024);
or U2121 (N_2121,N_1640,N_1667);
or U2122 (N_2122,N_1758,N_1378);
and U2123 (N_2123,N_1339,N_1271);
nand U2124 (N_2124,N_1838,N_1793);
and U2125 (N_2125,N_1568,N_1124);
or U2126 (N_2126,N_1627,N_1011);
nor U2127 (N_2127,N_1619,N_1234);
or U2128 (N_2128,N_1591,N_1733);
or U2129 (N_2129,N_1489,N_1209);
or U2130 (N_2130,N_1006,N_1298);
or U2131 (N_2131,N_1966,N_1989);
and U2132 (N_2132,N_1207,N_1414);
nor U2133 (N_2133,N_1029,N_1697);
or U2134 (N_2134,N_1861,N_1585);
xor U2135 (N_2135,N_1158,N_1302);
or U2136 (N_2136,N_1003,N_1656);
nand U2137 (N_2137,N_1995,N_1413);
nor U2138 (N_2138,N_1099,N_1676);
xor U2139 (N_2139,N_1731,N_1649);
or U2140 (N_2140,N_1692,N_1632);
xor U2141 (N_2141,N_1500,N_1435);
nand U2142 (N_2142,N_1322,N_1637);
or U2143 (N_2143,N_1582,N_1241);
nor U2144 (N_2144,N_1943,N_1816);
nor U2145 (N_2145,N_1872,N_1688);
nand U2146 (N_2146,N_1198,N_1103);
or U2147 (N_2147,N_1449,N_1517);
nor U2148 (N_2148,N_1071,N_1031);
nand U2149 (N_2149,N_1967,N_1232);
nand U2150 (N_2150,N_1651,N_1693);
nor U2151 (N_2151,N_1368,N_1716);
xnor U2152 (N_2152,N_1823,N_1137);
nand U2153 (N_2153,N_1392,N_1702);
and U2154 (N_2154,N_1192,N_1102);
or U2155 (N_2155,N_1538,N_1467);
and U2156 (N_2156,N_1310,N_1998);
and U2157 (N_2157,N_1197,N_1254);
xnor U2158 (N_2158,N_1615,N_1214);
nor U2159 (N_2159,N_1996,N_1830);
nor U2160 (N_2160,N_1655,N_1016);
nand U2161 (N_2161,N_1134,N_1959);
nor U2162 (N_2162,N_1136,N_1133);
or U2163 (N_2163,N_1132,N_1484);
and U2164 (N_2164,N_1372,N_1078);
and U2165 (N_2165,N_1376,N_1434);
or U2166 (N_2166,N_1150,N_1629);
and U2167 (N_2167,N_1149,N_1622);
nor U2168 (N_2168,N_1259,N_1222);
nor U2169 (N_2169,N_1783,N_1400);
or U2170 (N_2170,N_1564,N_1992);
or U2171 (N_2171,N_1523,N_1626);
nand U2172 (N_2172,N_1977,N_1225);
and U2173 (N_2173,N_1963,N_1613);
nor U2174 (N_2174,N_1272,N_1972);
and U2175 (N_2175,N_1905,N_1511);
nand U2176 (N_2176,N_1991,N_1574);
and U2177 (N_2177,N_1867,N_1335);
or U2178 (N_2178,N_1499,N_1200);
and U2179 (N_2179,N_1042,N_1802);
xor U2180 (N_2180,N_1915,N_1329);
or U2181 (N_2181,N_1478,N_1119);
and U2182 (N_2182,N_1605,N_1608);
nand U2183 (N_2183,N_1181,N_1874);
and U2184 (N_2184,N_1917,N_1087);
or U2185 (N_2185,N_1202,N_1588);
nand U2186 (N_2186,N_1974,N_1541);
nor U2187 (N_2187,N_1226,N_1877);
xor U2188 (N_2188,N_1032,N_1566);
and U2189 (N_2189,N_1054,N_1118);
nand U2190 (N_2190,N_1757,N_1983);
nor U2191 (N_2191,N_1151,N_1446);
and U2192 (N_2192,N_1349,N_1834);
and U2193 (N_2193,N_1558,N_1922);
nor U2194 (N_2194,N_1644,N_1826);
or U2195 (N_2195,N_1839,N_1000);
and U2196 (N_2196,N_1238,N_1433);
nand U2197 (N_2197,N_1447,N_1620);
nor U2198 (N_2198,N_1355,N_1545);
nor U2199 (N_2199,N_1533,N_1193);
xor U2200 (N_2200,N_1418,N_1837);
nand U2201 (N_2201,N_1596,N_1211);
nor U2202 (N_2202,N_1623,N_1025);
nand U2203 (N_2203,N_1796,N_1178);
or U2204 (N_2204,N_1868,N_1325);
xnor U2205 (N_2205,N_1825,N_1781);
or U2206 (N_2206,N_1661,N_1442);
or U2207 (N_2207,N_1223,N_1841);
or U2208 (N_2208,N_1906,N_1954);
or U2209 (N_2209,N_1156,N_1956);
nor U2210 (N_2210,N_1890,N_1046);
and U2211 (N_2211,N_1064,N_1108);
nand U2212 (N_2212,N_1516,N_1138);
or U2213 (N_2213,N_1166,N_1307);
or U2214 (N_2214,N_1395,N_1659);
nor U2215 (N_2215,N_1246,N_1634);
nor U2216 (N_2216,N_1455,N_1503);
xor U2217 (N_2217,N_1897,N_1862);
and U2218 (N_2218,N_1660,N_1848);
or U2219 (N_2219,N_1096,N_1001);
and U2220 (N_2220,N_1161,N_1055);
and U2221 (N_2221,N_1947,N_1811);
or U2222 (N_2222,N_1267,N_1440);
nand U2223 (N_2223,N_1201,N_1735);
or U2224 (N_2224,N_1021,N_1215);
nand U2225 (N_2225,N_1852,N_1399);
and U2226 (N_2226,N_1101,N_1070);
nand U2227 (N_2227,N_1155,N_1406);
xnor U2228 (N_2228,N_1923,N_1509);
nand U2229 (N_2229,N_1798,N_1162);
and U2230 (N_2230,N_1048,N_1273);
nand U2231 (N_2231,N_1788,N_1186);
nor U2232 (N_2232,N_1038,N_1894);
or U2233 (N_2233,N_1456,N_1065);
nand U2234 (N_2234,N_1206,N_1284);
nand U2235 (N_2235,N_1812,N_1885);
or U2236 (N_2236,N_1919,N_1373);
and U2237 (N_2237,N_1320,N_1982);
or U2238 (N_2238,N_1609,N_1607);
nand U2239 (N_2239,N_1940,N_1387);
and U2240 (N_2240,N_1343,N_1751);
nand U2241 (N_2241,N_1142,N_1856);
and U2242 (N_2242,N_1831,N_1289);
nand U2243 (N_2243,N_1496,N_1231);
and U2244 (N_2244,N_1199,N_1695);
nor U2245 (N_2245,N_1432,N_1669);
or U2246 (N_2246,N_1621,N_1542);
and U2247 (N_2247,N_1240,N_1985);
nor U2248 (N_2248,N_1614,N_1850);
nor U2249 (N_2249,N_1381,N_1643);
or U2250 (N_2250,N_1004,N_1552);
nor U2251 (N_2251,N_1750,N_1109);
or U2252 (N_2252,N_1385,N_1469);
or U2253 (N_2253,N_1912,N_1603);
nand U2254 (N_2254,N_1465,N_1098);
or U2255 (N_2255,N_1769,N_1033);
or U2256 (N_2256,N_1510,N_1043);
nand U2257 (N_2257,N_1865,N_1507);
nand U2258 (N_2258,N_1315,N_1248);
nand U2259 (N_2259,N_1817,N_1921);
nand U2260 (N_2260,N_1990,N_1237);
nand U2261 (N_2261,N_1664,N_1597);
nor U2262 (N_2262,N_1407,N_1679);
or U2263 (N_2263,N_1287,N_1712);
nor U2264 (N_2264,N_1183,N_1860);
nand U2265 (N_2265,N_1778,N_1829);
and U2266 (N_2266,N_1074,N_1041);
and U2267 (N_2267,N_1575,N_1964);
nand U2268 (N_2268,N_1057,N_1846);
nor U2269 (N_2269,N_1544,N_1131);
nor U2270 (N_2270,N_1044,N_1324);
and U2271 (N_2271,N_1729,N_1971);
or U2272 (N_2272,N_1683,N_1719);
xnor U2273 (N_2273,N_1291,N_1117);
nand U2274 (N_2274,N_1734,N_1986);
or U2275 (N_2275,N_1718,N_1901);
and U2276 (N_2276,N_1389,N_1306);
nand U2277 (N_2277,N_1938,N_1721);
xnor U2278 (N_2278,N_1081,N_1819);
and U2279 (N_2279,N_1059,N_1326);
or U2280 (N_2280,N_1097,N_1827);
xor U2281 (N_2281,N_1035,N_1682);
nor U2282 (N_2282,N_1550,N_1085);
nand U2283 (N_2283,N_1204,N_1473);
or U2284 (N_2284,N_1554,N_1120);
or U2285 (N_2285,N_1563,N_1285);
nand U2286 (N_2286,N_1945,N_1053);
nor U2287 (N_2287,N_1739,N_1673);
nor U2288 (N_2288,N_1371,N_1895);
nand U2289 (N_2289,N_1526,N_1942);
and U2290 (N_2290,N_1969,N_1230);
xnor U2291 (N_2291,N_1774,N_1191);
or U2292 (N_2292,N_1163,N_1129);
nand U2293 (N_2293,N_1581,N_1095);
and U2294 (N_2294,N_1010,N_1316);
nand U2295 (N_2295,N_1790,N_1080);
nor U2296 (N_2296,N_1738,N_1321);
or U2297 (N_2297,N_1612,N_1784);
and U2298 (N_2298,N_1369,N_1881);
or U2299 (N_2299,N_1005,N_1258);
nor U2300 (N_2300,N_1747,N_1727);
nand U2301 (N_2301,N_1367,N_1797);
or U2302 (N_2302,N_1461,N_1847);
or U2303 (N_2303,N_1380,N_1216);
nand U2304 (N_2304,N_1092,N_1345);
nor U2305 (N_2305,N_1761,N_1106);
xor U2306 (N_2306,N_1835,N_1939);
nor U2307 (N_2307,N_1815,N_1884);
nand U2308 (N_2308,N_1675,N_1579);
nor U2309 (N_2309,N_1949,N_1153);
nor U2310 (N_2310,N_1063,N_1236);
nor U2311 (N_2311,N_1892,N_1803);
or U2312 (N_2312,N_1026,N_1765);
or U2313 (N_2313,N_1045,N_1981);
and U2314 (N_2314,N_1187,N_1960);
nand U2315 (N_2315,N_1471,N_1278);
nand U2316 (N_2316,N_1436,N_1294);
nand U2317 (N_2317,N_1123,N_1914);
and U2318 (N_2318,N_1141,N_1713);
nand U2319 (N_2319,N_1340,N_1007);
nand U2320 (N_2320,N_1419,N_1642);
nand U2321 (N_2321,N_1076,N_1970);
nor U2322 (N_2322,N_1130,N_1913);
or U2323 (N_2323,N_1037,N_1595);
nor U2324 (N_2324,N_1576,N_1227);
or U2325 (N_2325,N_1741,N_1318);
nand U2326 (N_2326,N_1768,N_1012);
and U2327 (N_2327,N_1968,N_1409);
and U2328 (N_2328,N_1018,N_1090);
and U2329 (N_2329,N_1772,N_1674);
nand U2330 (N_2330,N_1610,N_1242);
or U2331 (N_2331,N_1933,N_1920);
nand U2332 (N_2332,N_1704,N_1512);
nand U2333 (N_2333,N_1354,N_1067);
nor U2334 (N_2334,N_1725,N_1744);
nor U2335 (N_2335,N_1353,N_1497);
nand U2336 (N_2336,N_1428,N_1317);
and U2337 (N_2337,N_1212,N_1668);
and U2338 (N_2338,N_1957,N_1876);
nor U2339 (N_2339,N_1501,N_1807);
nor U2340 (N_2340,N_1690,N_1331);
nor U2341 (N_2341,N_1515,N_1832);
nor U2342 (N_2342,N_1357,N_1737);
nand U2343 (N_2343,N_1777,N_1988);
or U2344 (N_2344,N_1539,N_1889);
nor U2345 (N_2345,N_1978,N_1245);
and U2346 (N_2346,N_1488,N_1265);
nand U2347 (N_2347,N_1785,N_1506);
and U2348 (N_2348,N_1364,N_1710);
and U2349 (N_2349,N_1556,N_1973);
and U2350 (N_2350,N_1114,N_1543);
or U2351 (N_2351,N_1487,N_1527);
nand U2352 (N_2352,N_1962,N_1535);
and U2353 (N_2353,N_1805,N_1224);
nor U2354 (N_2354,N_1720,N_1184);
xnor U2355 (N_2355,N_1334,N_1491);
and U2356 (N_2356,N_1266,N_1717);
or U2357 (N_2357,N_1694,N_1886);
or U2358 (N_2358,N_1139,N_1208);
and U2359 (N_2359,N_1089,N_1756);
and U2360 (N_2360,N_1775,N_1975);
or U2361 (N_2361,N_1430,N_1654);
nand U2362 (N_2362,N_1833,N_1342);
or U2363 (N_2363,N_1445,N_1047);
nand U2364 (N_2364,N_1177,N_1587);
or U2365 (N_2365,N_1536,N_1604);
xnor U2366 (N_2366,N_1390,N_1279);
nor U2367 (N_2367,N_1146,N_1027);
or U2368 (N_2368,N_1386,N_1330);
and U2369 (N_2369,N_1709,N_1058);
and U2370 (N_2370,N_1810,N_1270);
and U2371 (N_2371,N_1296,N_1094);
nor U2372 (N_2372,N_1175,N_1221);
nand U2373 (N_2373,N_1929,N_1480);
nor U2374 (N_2374,N_1481,N_1084);
and U2375 (N_2375,N_1658,N_1736);
or U2376 (N_2376,N_1927,N_1470);
or U2377 (N_2377,N_1135,N_1429);
and U2378 (N_2378,N_1293,N_1505);
xnor U2379 (N_2379,N_1742,N_1843);
nor U2380 (N_2380,N_1555,N_1050);
nand U2381 (N_2381,N_1916,N_1023);
xor U2382 (N_2382,N_1549,N_1030);
and U2383 (N_2383,N_1593,N_1586);
nor U2384 (N_2384,N_1840,N_1268);
nor U2385 (N_2385,N_1979,N_1451);
nor U2386 (N_2386,N_1281,N_1560);
and U2387 (N_2387,N_1910,N_1822);
xor U2388 (N_2388,N_1229,N_1143);
nand U2389 (N_2389,N_1474,N_1280);
and U2390 (N_2390,N_1365,N_1994);
nor U2391 (N_2391,N_1439,N_1168);
or U2392 (N_2392,N_1645,N_1696);
xor U2393 (N_2393,N_1276,N_1782);
and U2394 (N_2394,N_1976,N_1049);
and U2395 (N_2395,N_1745,N_1332);
and U2396 (N_2396,N_1580,N_1194);
or U2397 (N_2397,N_1498,N_1352);
nor U2398 (N_2398,N_1404,N_1924);
nand U2399 (N_2399,N_1559,N_1866);
or U2400 (N_2400,N_1377,N_1052);
nand U2401 (N_2401,N_1448,N_1174);
nand U2402 (N_2402,N_1292,N_1383);
nor U2403 (N_2403,N_1570,N_1477);
or U2404 (N_2404,N_1379,N_1553);
and U2405 (N_2405,N_1953,N_1431);
or U2406 (N_2406,N_1441,N_1172);
nand U2407 (N_2407,N_1728,N_1219);
nor U2408 (N_2408,N_1261,N_1873);
nand U2409 (N_2409,N_1752,N_1530);
nor U2410 (N_2410,N_1684,N_1557);
or U2411 (N_2411,N_1086,N_1691);
nor U2412 (N_2412,N_1584,N_1705);
nor U2413 (N_2413,N_1344,N_1532);
and U2414 (N_2414,N_1904,N_1726);
nor U2415 (N_2415,N_1374,N_1567);
or U2416 (N_2416,N_1900,N_1653);
xnor U2417 (N_2417,N_1732,N_1275);
and U2418 (N_2418,N_1902,N_1665);
xnor U2419 (N_2419,N_1190,N_1494);
and U2420 (N_2420,N_1454,N_1421);
or U2421 (N_2421,N_1672,N_1925);
or U2422 (N_2422,N_1128,N_1122);
or U2423 (N_2423,N_1313,N_1878);
nor U2424 (N_2424,N_1918,N_1760);
or U2425 (N_2425,N_1504,N_1426);
nand U2426 (N_2426,N_1482,N_1305);
nand U2427 (N_2427,N_1875,N_1126);
nand U2428 (N_2428,N_1073,N_1844);
and U2429 (N_2429,N_1495,N_1547);
and U2430 (N_2430,N_1485,N_1303);
and U2431 (N_2431,N_1359,N_1009);
or U2432 (N_2432,N_1213,N_1475);
nor U2433 (N_2433,N_1159,N_1410);
xnor U2434 (N_2434,N_1650,N_1677);
and U2435 (N_2435,N_1384,N_1551);
nor U2436 (N_2436,N_1502,N_1599);
or U2437 (N_2437,N_1486,N_1871);
nor U2438 (N_2438,N_1394,N_1932);
xnor U2439 (N_2439,N_1787,N_1304);
and U2440 (N_2440,N_1754,N_1993);
nand U2441 (N_2441,N_1112,N_1657);
and U2442 (N_2442,N_1483,N_1859);
xnor U2443 (N_2443,N_1625,N_1646);
and U2444 (N_2444,N_1260,N_1341);
nor U2445 (N_2445,N_1312,N_1911);
or U2446 (N_2446,N_1361,N_1965);
or U2447 (N_2447,N_1598,N_1356);
nor U2448 (N_2448,N_1671,N_1941);
and U2449 (N_2449,N_1808,N_1405);
nor U2450 (N_2450,N_1648,N_1463);
nor U2451 (N_2451,N_1100,N_1411);
nor U2452 (N_2452,N_1144,N_1472);
nor U2453 (N_2453,N_1617,N_1148);
nor U2454 (N_2454,N_1571,N_1125);
nor U2455 (N_2455,N_1170,N_1999);
nand U2456 (N_2456,N_1140,N_1370);
nand U2457 (N_2457,N_1855,N_1346);
nor U2458 (N_2458,N_1762,N_1388);
nor U2459 (N_2459,N_1955,N_1794);
nor U2460 (N_2460,N_1780,N_1743);
nand U2461 (N_2461,N_1853,N_1821);
or U2462 (N_2462,N_1040,N_1531);
xor U2463 (N_2463,N_1854,N_1814);
xor U2464 (N_2464,N_1252,N_1864);
or U2465 (N_2465,N_1635,N_1898);
or U2466 (N_2466,N_1508,N_1262);
nand U2467 (N_2467,N_1348,N_1182);
nor U2468 (N_2468,N_1327,N_1887);
nand U2469 (N_2469,N_1420,N_1396);
nor U2470 (N_2470,N_1746,N_1019);
nand U2471 (N_2471,N_1422,N_1630);
nor U2472 (N_2472,N_1239,N_1931);
and U2473 (N_2473,N_1740,N_1519);
and U2474 (N_2474,N_1606,N_1934);
and U2475 (N_2475,N_1157,N_1179);
nand U2476 (N_2476,N_1792,N_1573);
nor U2477 (N_2477,N_1680,N_1806);
and U2478 (N_2478,N_1351,N_1600);
xnor U2479 (N_2479,N_1401,N_1708);
and U2480 (N_2480,N_1393,N_1460);
nor U2481 (N_2481,N_1723,N_1583);
or U2482 (N_2482,N_1264,N_1464);
xnor U2483 (N_2483,N_1075,N_1333);
nand U2484 (N_2484,N_1301,N_1145);
nand U2485 (N_2485,N_1755,N_1243);
nand U2486 (N_2486,N_1256,N_1093);
and U2487 (N_2487,N_1111,N_1283);
xnor U2488 (N_2488,N_1800,N_1205);
and U2489 (N_2489,N_1251,N_1466);
and U2490 (N_2490,N_1869,N_1002);
or U2491 (N_2491,N_1749,N_1290);
or U2492 (N_2492,N_1036,N_1681);
and U2493 (N_2493,N_1776,N_1069);
nor U2494 (N_2494,N_1189,N_1524);
nand U2495 (N_2495,N_1269,N_1056);
nor U2496 (N_2496,N_1518,N_1602);
and U2497 (N_2497,N_1578,N_1013);
nand U2498 (N_2498,N_1715,N_1773);
nor U2499 (N_2499,N_1375,N_1437);
nor U2500 (N_2500,N_1241,N_1248);
xor U2501 (N_2501,N_1033,N_1530);
or U2502 (N_2502,N_1310,N_1113);
and U2503 (N_2503,N_1098,N_1870);
nor U2504 (N_2504,N_1415,N_1661);
nor U2505 (N_2505,N_1410,N_1422);
nor U2506 (N_2506,N_1491,N_1134);
nand U2507 (N_2507,N_1648,N_1482);
nand U2508 (N_2508,N_1577,N_1652);
and U2509 (N_2509,N_1017,N_1480);
nor U2510 (N_2510,N_1121,N_1446);
and U2511 (N_2511,N_1887,N_1854);
xor U2512 (N_2512,N_1958,N_1891);
nor U2513 (N_2513,N_1165,N_1384);
nand U2514 (N_2514,N_1757,N_1813);
or U2515 (N_2515,N_1675,N_1649);
or U2516 (N_2516,N_1418,N_1683);
nand U2517 (N_2517,N_1032,N_1940);
nand U2518 (N_2518,N_1893,N_1428);
and U2519 (N_2519,N_1287,N_1114);
nand U2520 (N_2520,N_1246,N_1601);
and U2521 (N_2521,N_1550,N_1291);
and U2522 (N_2522,N_1953,N_1130);
or U2523 (N_2523,N_1658,N_1663);
nor U2524 (N_2524,N_1158,N_1053);
and U2525 (N_2525,N_1192,N_1466);
and U2526 (N_2526,N_1491,N_1054);
xor U2527 (N_2527,N_1835,N_1457);
or U2528 (N_2528,N_1545,N_1223);
or U2529 (N_2529,N_1557,N_1354);
nor U2530 (N_2530,N_1030,N_1429);
xnor U2531 (N_2531,N_1503,N_1771);
or U2532 (N_2532,N_1788,N_1682);
nor U2533 (N_2533,N_1277,N_1823);
and U2534 (N_2534,N_1239,N_1091);
and U2535 (N_2535,N_1967,N_1954);
or U2536 (N_2536,N_1526,N_1965);
and U2537 (N_2537,N_1504,N_1199);
nand U2538 (N_2538,N_1091,N_1853);
xor U2539 (N_2539,N_1428,N_1000);
nor U2540 (N_2540,N_1058,N_1071);
xnor U2541 (N_2541,N_1665,N_1686);
or U2542 (N_2542,N_1150,N_1831);
nor U2543 (N_2543,N_1756,N_1107);
nand U2544 (N_2544,N_1999,N_1034);
and U2545 (N_2545,N_1651,N_1209);
or U2546 (N_2546,N_1824,N_1796);
nor U2547 (N_2547,N_1613,N_1480);
and U2548 (N_2548,N_1534,N_1239);
or U2549 (N_2549,N_1702,N_1495);
nand U2550 (N_2550,N_1591,N_1047);
or U2551 (N_2551,N_1631,N_1729);
nor U2552 (N_2552,N_1255,N_1927);
nand U2553 (N_2553,N_1688,N_1105);
or U2554 (N_2554,N_1272,N_1112);
xor U2555 (N_2555,N_1827,N_1786);
or U2556 (N_2556,N_1720,N_1612);
nand U2557 (N_2557,N_1499,N_1780);
nand U2558 (N_2558,N_1384,N_1884);
and U2559 (N_2559,N_1799,N_1196);
and U2560 (N_2560,N_1670,N_1034);
or U2561 (N_2561,N_1130,N_1438);
nor U2562 (N_2562,N_1573,N_1323);
and U2563 (N_2563,N_1009,N_1979);
nand U2564 (N_2564,N_1895,N_1767);
and U2565 (N_2565,N_1931,N_1826);
nor U2566 (N_2566,N_1015,N_1185);
nor U2567 (N_2567,N_1921,N_1854);
and U2568 (N_2568,N_1705,N_1042);
and U2569 (N_2569,N_1124,N_1225);
or U2570 (N_2570,N_1024,N_1179);
or U2571 (N_2571,N_1885,N_1575);
or U2572 (N_2572,N_1463,N_1200);
and U2573 (N_2573,N_1865,N_1784);
nand U2574 (N_2574,N_1424,N_1474);
xnor U2575 (N_2575,N_1642,N_1309);
xor U2576 (N_2576,N_1362,N_1396);
xor U2577 (N_2577,N_1217,N_1652);
nor U2578 (N_2578,N_1123,N_1275);
or U2579 (N_2579,N_1720,N_1923);
nand U2580 (N_2580,N_1266,N_1991);
nand U2581 (N_2581,N_1741,N_1864);
xnor U2582 (N_2582,N_1995,N_1750);
and U2583 (N_2583,N_1322,N_1931);
or U2584 (N_2584,N_1689,N_1351);
xor U2585 (N_2585,N_1653,N_1901);
nand U2586 (N_2586,N_1195,N_1271);
nor U2587 (N_2587,N_1237,N_1302);
nor U2588 (N_2588,N_1923,N_1155);
nor U2589 (N_2589,N_1495,N_1621);
xor U2590 (N_2590,N_1830,N_1032);
and U2591 (N_2591,N_1415,N_1772);
or U2592 (N_2592,N_1058,N_1781);
nor U2593 (N_2593,N_1386,N_1369);
and U2594 (N_2594,N_1973,N_1853);
nand U2595 (N_2595,N_1410,N_1564);
nand U2596 (N_2596,N_1325,N_1292);
or U2597 (N_2597,N_1928,N_1626);
xor U2598 (N_2598,N_1543,N_1546);
and U2599 (N_2599,N_1501,N_1753);
nor U2600 (N_2600,N_1670,N_1161);
xnor U2601 (N_2601,N_1366,N_1774);
nor U2602 (N_2602,N_1161,N_1825);
nand U2603 (N_2603,N_1954,N_1692);
nand U2604 (N_2604,N_1207,N_1020);
nor U2605 (N_2605,N_1058,N_1496);
nor U2606 (N_2606,N_1668,N_1395);
or U2607 (N_2607,N_1058,N_1117);
xnor U2608 (N_2608,N_1745,N_1818);
nor U2609 (N_2609,N_1825,N_1872);
xnor U2610 (N_2610,N_1634,N_1465);
or U2611 (N_2611,N_1722,N_1561);
or U2612 (N_2612,N_1550,N_1053);
nand U2613 (N_2613,N_1369,N_1479);
nand U2614 (N_2614,N_1402,N_1973);
xnor U2615 (N_2615,N_1113,N_1293);
and U2616 (N_2616,N_1242,N_1992);
or U2617 (N_2617,N_1979,N_1273);
xor U2618 (N_2618,N_1662,N_1258);
nand U2619 (N_2619,N_1017,N_1343);
and U2620 (N_2620,N_1549,N_1080);
nor U2621 (N_2621,N_1700,N_1266);
and U2622 (N_2622,N_1390,N_1812);
or U2623 (N_2623,N_1455,N_1211);
nand U2624 (N_2624,N_1037,N_1629);
nor U2625 (N_2625,N_1995,N_1118);
or U2626 (N_2626,N_1768,N_1750);
and U2627 (N_2627,N_1095,N_1612);
and U2628 (N_2628,N_1698,N_1920);
nand U2629 (N_2629,N_1670,N_1607);
or U2630 (N_2630,N_1965,N_1533);
and U2631 (N_2631,N_1014,N_1081);
nand U2632 (N_2632,N_1249,N_1165);
and U2633 (N_2633,N_1679,N_1288);
and U2634 (N_2634,N_1471,N_1630);
nor U2635 (N_2635,N_1440,N_1914);
nand U2636 (N_2636,N_1108,N_1055);
and U2637 (N_2637,N_1907,N_1850);
xnor U2638 (N_2638,N_1403,N_1825);
or U2639 (N_2639,N_1033,N_1670);
nand U2640 (N_2640,N_1615,N_1216);
and U2641 (N_2641,N_1266,N_1417);
or U2642 (N_2642,N_1510,N_1127);
or U2643 (N_2643,N_1921,N_1771);
nor U2644 (N_2644,N_1444,N_1010);
nand U2645 (N_2645,N_1497,N_1052);
or U2646 (N_2646,N_1999,N_1444);
and U2647 (N_2647,N_1716,N_1334);
nand U2648 (N_2648,N_1606,N_1246);
or U2649 (N_2649,N_1523,N_1724);
nand U2650 (N_2650,N_1579,N_1992);
nand U2651 (N_2651,N_1366,N_1378);
nand U2652 (N_2652,N_1001,N_1865);
or U2653 (N_2653,N_1070,N_1029);
nand U2654 (N_2654,N_1403,N_1348);
nor U2655 (N_2655,N_1336,N_1914);
and U2656 (N_2656,N_1327,N_1077);
and U2657 (N_2657,N_1237,N_1882);
nor U2658 (N_2658,N_1878,N_1458);
nor U2659 (N_2659,N_1496,N_1115);
or U2660 (N_2660,N_1405,N_1143);
or U2661 (N_2661,N_1577,N_1969);
nor U2662 (N_2662,N_1234,N_1635);
or U2663 (N_2663,N_1335,N_1953);
and U2664 (N_2664,N_1955,N_1539);
nand U2665 (N_2665,N_1674,N_1324);
nor U2666 (N_2666,N_1326,N_1701);
nor U2667 (N_2667,N_1218,N_1778);
nand U2668 (N_2668,N_1847,N_1487);
xnor U2669 (N_2669,N_1825,N_1527);
nor U2670 (N_2670,N_1039,N_1335);
nor U2671 (N_2671,N_1711,N_1203);
nand U2672 (N_2672,N_1491,N_1833);
and U2673 (N_2673,N_1151,N_1178);
or U2674 (N_2674,N_1724,N_1619);
nor U2675 (N_2675,N_1046,N_1731);
and U2676 (N_2676,N_1257,N_1538);
and U2677 (N_2677,N_1650,N_1081);
or U2678 (N_2678,N_1602,N_1202);
nor U2679 (N_2679,N_1804,N_1177);
nor U2680 (N_2680,N_1747,N_1917);
nand U2681 (N_2681,N_1635,N_1349);
or U2682 (N_2682,N_1683,N_1235);
and U2683 (N_2683,N_1112,N_1976);
and U2684 (N_2684,N_1495,N_1529);
nand U2685 (N_2685,N_1933,N_1935);
or U2686 (N_2686,N_1549,N_1965);
xor U2687 (N_2687,N_1576,N_1545);
nand U2688 (N_2688,N_1525,N_1643);
or U2689 (N_2689,N_1511,N_1183);
or U2690 (N_2690,N_1805,N_1863);
nor U2691 (N_2691,N_1142,N_1361);
nor U2692 (N_2692,N_1581,N_1335);
nand U2693 (N_2693,N_1254,N_1422);
or U2694 (N_2694,N_1653,N_1152);
or U2695 (N_2695,N_1759,N_1145);
or U2696 (N_2696,N_1513,N_1289);
nor U2697 (N_2697,N_1796,N_1671);
xnor U2698 (N_2698,N_1903,N_1789);
and U2699 (N_2699,N_1476,N_1376);
and U2700 (N_2700,N_1038,N_1759);
or U2701 (N_2701,N_1318,N_1883);
nand U2702 (N_2702,N_1653,N_1581);
or U2703 (N_2703,N_1891,N_1107);
and U2704 (N_2704,N_1968,N_1619);
nand U2705 (N_2705,N_1201,N_1115);
nand U2706 (N_2706,N_1552,N_1885);
nor U2707 (N_2707,N_1200,N_1427);
nand U2708 (N_2708,N_1041,N_1753);
and U2709 (N_2709,N_1842,N_1226);
or U2710 (N_2710,N_1610,N_1091);
nor U2711 (N_2711,N_1029,N_1417);
nand U2712 (N_2712,N_1061,N_1436);
or U2713 (N_2713,N_1962,N_1304);
nor U2714 (N_2714,N_1952,N_1440);
and U2715 (N_2715,N_1852,N_1510);
or U2716 (N_2716,N_1036,N_1712);
nand U2717 (N_2717,N_1736,N_1259);
xnor U2718 (N_2718,N_1911,N_1338);
or U2719 (N_2719,N_1330,N_1283);
and U2720 (N_2720,N_1137,N_1329);
and U2721 (N_2721,N_1987,N_1357);
nor U2722 (N_2722,N_1522,N_1602);
and U2723 (N_2723,N_1502,N_1711);
or U2724 (N_2724,N_1357,N_1666);
nand U2725 (N_2725,N_1003,N_1872);
and U2726 (N_2726,N_1124,N_1276);
xnor U2727 (N_2727,N_1326,N_1474);
nor U2728 (N_2728,N_1318,N_1256);
or U2729 (N_2729,N_1705,N_1842);
or U2730 (N_2730,N_1017,N_1461);
nor U2731 (N_2731,N_1225,N_1617);
nand U2732 (N_2732,N_1896,N_1755);
nor U2733 (N_2733,N_1441,N_1459);
nand U2734 (N_2734,N_1603,N_1960);
and U2735 (N_2735,N_1545,N_1755);
or U2736 (N_2736,N_1645,N_1098);
or U2737 (N_2737,N_1058,N_1556);
nor U2738 (N_2738,N_1999,N_1524);
xor U2739 (N_2739,N_1600,N_1561);
and U2740 (N_2740,N_1830,N_1314);
or U2741 (N_2741,N_1952,N_1428);
and U2742 (N_2742,N_1298,N_1945);
and U2743 (N_2743,N_1223,N_1661);
nor U2744 (N_2744,N_1872,N_1557);
nand U2745 (N_2745,N_1453,N_1648);
or U2746 (N_2746,N_1213,N_1279);
and U2747 (N_2747,N_1913,N_1570);
or U2748 (N_2748,N_1411,N_1626);
xnor U2749 (N_2749,N_1759,N_1402);
xor U2750 (N_2750,N_1368,N_1173);
or U2751 (N_2751,N_1686,N_1775);
xor U2752 (N_2752,N_1818,N_1391);
xnor U2753 (N_2753,N_1471,N_1350);
or U2754 (N_2754,N_1648,N_1965);
nor U2755 (N_2755,N_1438,N_1343);
or U2756 (N_2756,N_1232,N_1746);
and U2757 (N_2757,N_1463,N_1939);
nand U2758 (N_2758,N_1281,N_1131);
nand U2759 (N_2759,N_1969,N_1290);
xnor U2760 (N_2760,N_1655,N_1707);
and U2761 (N_2761,N_1491,N_1411);
and U2762 (N_2762,N_1873,N_1346);
or U2763 (N_2763,N_1631,N_1751);
xnor U2764 (N_2764,N_1840,N_1185);
nor U2765 (N_2765,N_1546,N_1929);
nor U2766 (N_2766,N_1515,N_1761);
nand U2767 (N_2767,N_1766,N_1175);
nor U2768 (N_2768,N_1413,N_1615);
nor U2769 (N_2769,N_1354,N_1075);
nand U2770 (N_2770,N_1248,N_1593);
and U2771 (N_2771,N_1364,N_1346);
or U2772 (N_2772,N_1521,N_1283);
nand U2773 (N_2773,N_1697,N_1401);
nor U2774 (N_2774,N_1669,N_1925);
nand U2775 (N_2775,N_1427,N_1118);
or U2776 (N_2776,N_1217,N_1720);
or U2777 (N_2777,N_1561,N_1092);
or U2778 (N_2778,N_1063,N_1124);
or U2779 (N_2779,N_1097,N_1817);
nor U2780 (N_2780,N_1403,N_1382);
nand U2781 (N_2781,N_1444,N_1729);
nand U2782 (N_2782,N_1393,N_1201);
and U2783 (N_2783,N_1803,N_1752);
and U2784 (N_2784,N_1511,N_1222);
and U2785 (N_2785,N_1245,N_1263);
or U2786 (N_2786,N_1373,N_1638);
nor U2787 (N_2787,N_1158,N_1598);
nand U2788 (N_2788,N_1772,N_1462);
nand U2789 (N_2789,N_1679,N_1757);
and U2790 (N_2790,N_1047,N_1927);
nand U2791 (N_2791,N_1468,N_1345);
and U2792 (N_2792,N_1170,N_1512);
nand U2793 (N_2793,N_1203,N_1801);
nor U2794 (N_2794,N_1154,N_1580);
nor U2795 (N_2795,N_1794,N_1264);
nor U2796 (N_2796,N_1607,N_1311);
and U2797 (N_2797,N_1175,N_1882);
nor U2798 (N_2798,N_1606,N_1928);
nor U2799 (N_2799,N_1007,N_1532);
xnor U2800 (N_2800,N_1562,N_1028);
and U2801 (N_2801,N_1014,N_1962);
or U2802 (N_2802,N_1129,N_1858);
and U2803 (N_2803,N_1881,N_1987);
nand U2804 (N_2804,N_1717,N_1815);
xnor U2805 (N_2805,N_1570,N_1755);
nand U2806 (N_2806,N_1161,N_1909);
nand U2807 (N_2807,N_1495,N_1653);
nand U2808 (N_2808,N_1725,N_1805);
and U2809 (N_2809,N_1696,N_1608);
nand U2810 (N_2810,N_1973,N_1348);
and U2811 (N_2811,N_1927,N_1174);
or U2812 (N_2812,N_1272,N_1663);
nand U2813 (N_2813,N_1207,N_1052);
or U2814 (N_2814,N_1365,N_1640);
or U2815 (N_2815,N_1399,N_1864);
nor U2816 (N_2816,N_1455,N_1861);
and U2817 (N_2817,N_1046,N_1588);
and U2818 (N_2818,N_1764,N_1375);
nor U2819 (N_2819,N_1519,N_1318);
nor U2820 (N_2820,N_1300,N_1692);
or U2821 (N_2821,N_1192,N_1620);
nor U2822 (N_2822,N_1471,N_1419);
or U2823 (N_2823,N_1004,N_1484);
and U2824 (N_2824,N_1399,N_1854);
xor U2825 (N_2825,N_1645,N_1665);
and U2826 (N_2826,N_1674,N_1407);
and U2827 (N_2827,N_1356,N_1114);
and U2828 (N_2828,N_1181,N_1945);
nor U2829 (N_2829,N_1040,N_1157);
or U2830 (N_2830,N_1015,N_1849);
nand U2831 (N_2831,N_1248,N_1855);
nor U2832 (N_2832,N_1176,N_1751);
nand U2833 (N_2833,N_1312,N_1462);
and U2834 (N_2834,N_1162,N_1097);
or U2835 (N_2835,N_1420,N_1970);
nand U2836 (N_2836,N_1637,N_1818);
or U2837 (N_2837,N_1204,N_1822);
nand U2838 (N_2838,N_1694,N_1471);
and U2839 (N_2839,N_1466,N_1203);
nor U2840 (N_2840,N_1002,N_1738);
or U2841 (N_2841,N_1358,N_1080);
and U2842 (N_2842,N_1407,N_1628);
or U2843 (N_2843,N_1718,N_1977);
and U2844 (N_2844,N_1149,N_1033);
or U2845 (N_2845,N_1016,N_1454);
or U2846 (N_2846,N_1557,N_1341);
nand U2847 (N_2847,N_1212,N_1218);
and U2848 (N_2848,N_1044,N_1649);
xnor U2849 (N_2849,N_1704,N_1347);
nand U2850 (N_2850,N_1276,N_1248);
xnor U2851 (N_2851,N_1877,N_1959);
nor U2852 (N_2852,N_1795,N_1374);
or U2853 (N_2853,N_1581,N_1741);
and U2854 (N_2854,N_1229,N_1157);
xor U2855 (N_2855,N_1406,N_1393);
nand U2856 (N_2856,N_1804,N_1097);
nor U2857 (N_2857,N_1793,N_1862);
nand U2858 (N_2858,N_1557,N_1036);
nor U2859 (N_2859,N_1539,N_1502);
or U2860 (N_2860,N_1910,N_1767);
or U2861 (N_2861,N_1132,N_1066);
and U2862 (N_2862,N_1230,N_1777);
nor U2863 (N_2863,N_1530,N_1426);
nor U2864 (N_2864,N_1386,N_1524);
and U2865 (N_2865,N_1413,N_1099);
and U2866 (N_2866,N_1213,N_1227);
nand U2867 (N_2867,N_1090,N_1803);
or U2868 (N_2868,N_1842,N_1506);
nor U2869 (N_2869,N_1944,N_1269);
nor U2870 (N_2870,N_1921,N_1850);
nand U2871 (N_2871,N_1356,N_1314);
or U2872 (N_2872,N_1109,N_1785);
nor U2873 (N_2873,N_1867,N_1090);
and U2874 (N_2874,N_1289,N_1288);
xnor U2875 (N_2875,N_1723,N_1479);
nor U2876 (N_2876,N_1721,N_1998);
nand U2877 (N_2877,N_1578,N_1746);
nor U2878 (N_2878,N_1082,N_1419);
or U2879 (N_2879,N_1134,N_1487);
xor U2880 (N_2880,N_1408,N_1836);
nand U2881 (N_2881,N_1721,N_1010);
or U2882 (N_2882,N_1295,N_1983);
and U2883 (N_2883,N_1450,N_1258);
or U2884 (N_2884,N_1802,N_1504);
nand U2885 (N_2885,N_1869,N_1138);
xnor U2886 (N_2886,N_1210,N_1796);
xor U2887 (N_2887,N_1432,N_1789);
nor U2888 (N_2888,N_1758,N_1109);
and U2889 (N_2889,N_1230,N_1885);
nand U2890 (N_2890,N_1760,N_1647);
and U2891 (N_2891,N_1139,N_1520);
nor U2892 (N_2892,N_1355,N_1207);
nand U2893 (N_2893,N_1368,N_1269);
nor U2894 (N_2894,N_1048,N_1889);
and U2895 (N_2895,N_1195,N_1831);
and U2896 (N_2896,N_1471,N_1947);
or U2897 (N_2897,N_1059,N_1835);
or U2898 (N_2898,N_1844,N_1811);
and U2899 (N_2899,N_1908,N_1396);
or U2900 (N_2900,N_1447,N_1384);
nand U2901 (N_2901,N_1378,N_1792);
or U2902 (N_2902,N_1177,N_1365);
and U2903 (N_2903,N_1461,N_1456);
nand U2904 (N_2904,N_1049,N_1024);
nand U2905 (N_2905,N_1175,N_1271);
or U2906 (N_2906,N_1025,N_1001);
xnor U2907 (N_2907,N_1547,N_1774);
nand U2908 (N_2908,N_1546,N_1374);
and U2909 (N_2909,N_1574,N_1485);
nand U2910 (N_2910,N_1940,N_1517);
xnor U2911 (N_2911,N_1714,N_1077);
nor U2912 (N_2912,N_1533,N_1937);
and U2913 (N_2913,N_1700,N_1679);
and U2914 (N_2914,N_1316,N_1161);
nand U2915 (N_2915,N_1003,N_1084);
xor U2916 (N_2916,N_1217,N_1855);
and U2917 (N_2917,N_1607,N_1391);
or U2918 (N_2918,N_1015,N_1574);
and U2919 (N_2919,N_1817,N_1906);
and U2920 (N_2920,N_1461,N_1865);
and U2921 (N_2921,N_1379,N_1490);
and U2922 (N_2922,N_1394,N_1922);
or U2923 (N_2923,N_1503,N_1658);
nand U2924 (N_2924,N_1140,N_1570);
and U2925 (N_2925,N_1160,N_1019);
nor U2926 (N_2926,N_1989,N_1973);
or U2927 (N_2927,N_1076,N_1730);
xnor U2928 (N_2928,N_1237,N_1732);
nand U2929 (N_2929,N_1428,N_1918);
nand U2930 (N_2930,N_1842,N_1071);
and U2931 (N_2931,N_1293,N_1182);
nand U2932 (N_2932,N_1154,N_1917);
nor U2933 (N_2933,N_1376,N_1976);
nand U2934 (N_2934,N_1585,N_1205);
or U2935 (N_2935,N_1953,N_1633);
or U2936 (N_2936,N_1763,N_1411);
or U2937 (N_2937,N_1048,N_1697);
xnor U2938 (N_2938,N_1651,N_1486);
xor U2939 (N_2939,N_1407,N_1369);
nor U2940 (N_2940,N_1522,N_1690);
nor U2941 (N_2941,N_1884,N_1810);
nand U2942 (N_2942,N_1423,N_1661);
or U2943 (N_2943,N_1303,N_1121);
nand U2944 (N_2944,N_1478,N_1437);
and U2945 (N_2945,N_1853,N_1544);
and U2946 (N_2946,N_1597,N_1499);
nand U2947 (N_2947,N_1109,N_1059);
nand U2948 (N_2948,N_1149,N_1309);
and U2949 (N_2949,N_1042,N_1568);
nand U2950 (N_2950,N_1291,N_1860);
and U2951 (N_2951,N_1863,N_1012);
nor U2952 (N_2952,N_1496,N_1483);
nor U2953 (N_2953,N_1040,N_1788);
or U2954 (N_2954,N_1464,N_1709);
nor U2955 (N_2955,N_1755,N_1821);
nand U2956 (N_2956,N_1702,N_1435);
or U2957 (N_2957,N_1396,N_1771);
nor U2958 (N_2958,N_1271,N_1067);
xor U2959 (N_2959,N_1477,N_1164);
and U2960 (N_2960,N_1389,N_1466);
nand U2961 (N_2961,N_1518,N_1121);
nand U2962 (N_2962,N_1179,N_1793);
xor U2963 (N_2963,N_1220,N_1473);
nor U2964 (N_2964,N_1259,N_1750);
or U2965 (N_2965,N_1953,N_1267);
nor U2966 (N_2966,N_1591,N_1068);
xnor U2967 (N_2967,N_1877,N_1723);
and U2968 (N_2968,N_1893,N_1240);
nor U2969 (N_2969,N_1656,N_1497);
xnor U2970 (N_2970,N_1128,N_1746);
nand U2971 (N_2971,N_1461,N_1934);
nand U2972 (N_2972,N_1890,N_1815);
or U2973 (N_2973,N_1462,N_1183);
nor U2974 (N_2974,N_1045,N_1790);
or U2975 (N_2975,N_1233,N_1892);
xnor U2976 (N_2976,N_1637,N_1575);
nand U2977 (N_2977,N_1027,N_1562);
or U2978 (N_2978,N_1985,N_1682);
or U2979 (N_2979,N_1149,N_1841);
or U2980 (N_2980,N_1964,N_1056);
nor U2981 (N_2981,N_1917,N_1935);
and U2982 (N_2982,N_1918,N_1267);
and U2983 (N_2983,N_1316,N_1934);
xnor U2984 (N_2984,N_1180,N_1640);
xnor U2985 (N_2985,N_1594,N_1005);
and U2986 (N_2986,N_1162,N_1828);
nand U2987 (N_2987,N_1704,N_1281);
nand U2988 (N_2988,N_1853,N_1401);
nor U2989 (N_2989,N_1993,N_1209);
nor U2990 (N_2990,N_1415,N_1582);
nor U2991 (N_2991,N_1834,N_1035);
and U2992 (N_2992,N_1165,N_1829);
and U2993 (N_2993,N_1038,N_1031);
nor U2994 (N_2994,N_1153,N_1874);
nor U2995 (N_2995,N_1868,N_1566);
xor U2996 (N_2996,N_1532,N_1778);
nand U2997 (N_2997,N_1023,N_1540);
and U2998 (N_2998,N_1458,N_1008);
or U2999 (N_2999,N_1362,N_1948);
nor UO_0 (O_0,N_2051,N_2345);
and UO_1 (O_1,N_2480,N_2990);
nor UO_2 (O_2,N_2607,N_2939);
xnor UO_3 (O_3,N_2694,N_2123);
nor UO_4 (O_4,N_2011,N_2549);
and UO_5 (O_5,N_2100,N_2054);
nor UO_6 (O_6,N_2908,N_2073);
or UO_7 (O_7,N_2926,N_2696);
and UO_8 (O_8,N_2435,N_2035);
xnor UO_9 (O_9,N_2765,N_2910);
and UO_10 (O_10,N_2555,N_2064);
and UO_11 (O_11,N_2677,N_2157);
and UO_12 (O_12,N_2037,N_2657);
or UO_13 (O_13,N_2308,N_2568);
nor UO_14 (O_14,N_2986,N_2211);
nand UO_15 (O_15,N_2843,N_2659);
and UO_16 (O_16,N_2961,N_2286);
nor UO_17 (O_17,N_2400,N_2270);
or UO_18 (O_18,N_2040,N_2902);
and UO_19 (O_19,N_2953,N_2228);
and UO_20 (O_20,N_2869,N_2274);
and UO_21 (O_21,N_2213,N_2331);
or UO_22 (O_22,N_2871,N_2716);
nand UO_23 (O_23,N_2505,N_2605);
nor UO_24 (O_24,N_2097,N_2641);
and UO_25 (O_25,N_2614,N_2457);
nor UO_26 (O_26,N_2976,N_2998);
and UO_27 (O_27,N_2580,N_2341);
nand UO_28 (O_28,N_2850,N_2978);
nor UO_29 (O_29,N_2380,N_2662);
or UO_30 (O_30,N_2646,N_2179);
or UO_31 (O_31,N_2323,N_2918);
xor UO_32 (O_32,N_2676,N_2470);
nor UO_33 (O_33,N_2015,N_2279);
or UO_34 (O_34,N_2152,N_2726);
nand UO_35 (O_35,N_2068,N_2429);
and UO_36 (O_36,N_2298,N_2132);
nor UO_37 (O_37,N_2236,N_2810);
nand UO_38 (O_38,N_2455,N_2388);
nor UO_39 (O_39,N_2326,N_2249);
and UO_40 (O_40,N_2940,N_2729);
or UO_41 (O_41,N_2027,N_2129);
or UO_42 (O_42,N_2030,N_2122);
nand UO_43 (O_43,N_2565,N_2645);
nor UO_44 (O_44,N_2526,N_2651);
or UO_45 (O_45,N_2250,N_2784);
nand UO_46 (O_46,N_2453,N_2300);
and UO_47 (O_47,N_2629,N_2672);
nand UO_48 (O_48,N_2410,N_2234);
nand UO_49 (O_49,N_2118,N_2924);
nand UO_50 (O_50,N_2823,N_2570);
xor UO_51 (O_51,N_2116,N_2596);
nor UO_52 (O_52,N_2535,N_2194);
nor UO_53 (O_53,N_2377,N_2255);
xnor UO_54 (O_54,N_2691,N_2876);
or UO_55 (O_55,N_2577,N_2114);
or UO_56 (O_56,N_2099,N_2635);
and UO_57 (O_57,N_2833,N_2995);
or UO_58 (O_58,N_2412,N_2170);
xnor UO_59 (O_59,N_2649,N_2959);
xor UO_60 (O_60,N_2973,N_2550);
and UO_61 (O_61,N_2531,N_2151);
and UO_62 (O_62,N_2057,N_2022);
nor UO_63 (O_63,N_2688,N_2751);
nor UO_64 (O_64,N_2439,N_2746);
or UO_65 (O_65,N_2778,N_2463);
nor UO_66 (O_66,N_2163,N_2386);
or UO_67 (O_67,N_2897,N_2942);
and UO_68 (O_68,N_2533,N_2311);
nand UO_69 (O_69,N_2357,N_2725);
and UO_70 (O_70,N_2822,N_2447);
and UO_71 (O_71,N_2898,N_2825);
nand UO_72 (O_72,N_2665,N_2985);
or UO_73 (O_73,N_2623,N_2306);
and UO_74 (O_74,N_2759,N_2436);
nand UO_75 (O_75,N_2102,N_2322);
nand UO_76 (O_76,N_2144,N_2711);
and UO_77 (O_77,N_2090,N_2553);
nor UO_78 (O_78,N_2143,N_2736);
nand UO_79 (O_79,N_2133,N_2834);
and UO_80 (O_80,N_2445,N_2950);
or UO_81 (O_81,N_2372,N_2797);
nor UO_82 (O_82,N_2437,N_2220);
nand UO_83 (O_83,N_2256,N_2328);
or UO_84 (O_84,N_2595,N_2363);
or UO_85 (O_85,N_2957,N_2342);
xnor UO_86 (O_86,N_2544,N_2055);
and UO_87 (O_87,N_2227,N_2415);
and UO_88 (O_88,N_2232,N_2919);
xnor UO_89 (O_89,N_2408,N_2799);
or UO_90 (O_90,N_2273,N_2999);
or UO_91 (O_91,N_2171,N_2356);
xor UO_92 (O_92,N_2317,N_2233);
xnor UO_93 (O_93,N_2224,N_2793);
or UO_94 (O_94,N_2977,N_2126);
nor UO_95 (O_95,N_2534,N_2110);
xor UO_96 (O_96,N_2837,N_2839);
and UO_97 (O_97,N_2589,N_2085);
nor UO_98 (O_98,N_2643,N_2492);
nor UO_99 (O_99,N_2530,N_2347);
nor UO_100 (O_100,N_2310,N_2841);
and UO_101 (O_101,N_2218,N_2974);
nor UO_102 (O_102,N_2134,N_2146);
xor UO_103 (O_103,N_2174,N_2744);
or UO_104 (O_104,N_2047,N_2222);
xor UO_105 (O_105,N_2597,N_2087);
and UO_106 (O_106,N_2283,N_2703);
and UO_107 (O_107,N_2755,N_2259);
nand UO_108 (O_108,N_2483,N_2873);
nor UO_109 (O_109,N_2714,N_2655);
nor UO_110 (O_110,N_2512,N_2658);
or UO_111 (O_111,N_2241,N_2208);
and UO_112 (O_112,N_2066,N_2251);
nand UO_113 (O_113,N_2007,N_2774);
xor UO_114 (O_114,N_2588,N_2147);
and UO_115 (O_115,N_2325,N_2804);
nand UO_116 (O_116,N_2954,N_2185);
xnor UO_117 (O_117,N_2316,N_2896);
or UO_118 (O_118,N_2290,N_2014);
and UO_119 (O_119,N_2851,N_2814);
or UO_120 (O_120,N_2956,N_2993);
nand UO_121 (O_121,N_2466,N_2141);
xnor UO_122 (O_122,N_2656,N_2121);
xor UO_123 (O_123,N_2769,N_2689);
nand UO_124 (O_124,N_2359,N_2642);
nor UO_125 (O_125,N_2315,N_2382);
and UO_126 (O_126,N_2667,N_2265);
and UO_127 (O_127,N_2478,N_2237);
or UO_128 (O_128,N_2089,N_2023);
or UO_129 (O_129,N_2187,N_2422);
and UO_130 (O_130,N_2739,N_2970);
nand UO_131 (O_131,N_2829,N_2922);
nand UO_132 (O_132,N_2601,N_2581);
or UO_133 (O_133,N_2852,N_2708);
or UO_134 (O_134,N_2749,N_2038);
or UO_135 (O_135,N_2285,N_2197);
nor UO_136 (O_136,N_2547,N_2883);
or UO_137 (O_137,N_2375,N_2604);
nor UO_138 (O_138,N_2067,N_2154);
and UO_139 (O_139,N_2488,N_2301);
nand UO_140 (O_140,N_2448,N_2442);
or UO_141 (O_141,N_2859,N_2603);
and UO_142 (O_142,N_2562,N_2836);
xor UO_143 (O_143,N_2812,N_2551);
or UO_144 (O_144,N_2167,N_2028);
nor UO_145 (O_145,N_2210,N_2881);
nor UO_146 (O_146,N_2907,N_2862);
nor UO_147 (O_147,N_2292,N_2299);
or UO_148 (O_148,N_2631,N_2206);
or UO_149 (O_149,N_2679,N_2148);
and UO_150 (O_150,N_2639,N_2606);
nand UO_151 (O_151,N_2518,N_2039);
and UO_152 (O_152,N_2390,N_2107);
nand UO_153 (O_153,N_2928,N_2021);
or UO_154 (O_154,N_2405,N_2465);
nand UO_155 (O_155,N_2093,N_2888);
xor UO_156 (O_156,N_2891,N_2666);
xnor UO_157 (O_157,N_2202,N_2450);
xnor UO_158 (O_158,N_2282,N_2225);
nand UO_159 (O_159,N_2594,N_2846);
nor UO_160 (O_160,N_2710,N_2702);
nor UO_161 (O_161,N_2756,N_2712);
nor UO_162 (O_162,N_2190,N_2675);
or UO_163 (O_163,N_2901,N_2625);
or UO_164 (O_164,N_2360,N_2955);
and UO_165 (O_165,N_2303,N_2351);
or UO_166 (O_166,N_2767,N_2540);
nand UO_167 (O_167,N_2403,N_2223);
and UO_168 (O_168,N_2262,N_2006);
nand UO_169 (O_169,N_2293,N_2280);
and UO_170 (O_170,N_2748,N_2046);
nand UO_171 (O_171,N_2766,N_2002);
or UO_172 (O_172,N_2681,N_2169);
nand UO_173 (O_173,N_2644,N_2117);
or UO_174 (O_174,N_2515,N_2692);
nor UO_175 (O_175,N_2567,N_2307);
or UO_176 (O_176,N_2199,N_2352);
nor UO_177 (O_177,N_2091,N_2525);
or UO_178 (O_178,N_2608,N_2140);
nand UO_179 (O_179,N_2468,N_2387);
and UO_180 (O_180,N_2879,N_2272);
nand UO_181 (O_181,N_2018,N_2821);
and UO_182 (O_182,N_2212,N_2680);
nand UO_183 (O_183,N_2886,N_2240);
nand UO_184 (O_184,N_2997,N_2699);
and UO_185 (O_185,N_2162,N_2695);
xnor UO_186 (O_186,N_2800,N_2678);
and UO_187 (O_187,N_2640,N_2059);
xnor UO_188 (O_188,N_2034,N_2269);
nand UO_189 (O_189,N_2231,N_2032);
nand UO_190 (O_190,N_2776,N_2747);
xnor UO_191 (O_191,N_2494,N_2284);
and UO_192 (O_192,N_2854,N_2795);
and UO_193 (O_193,N_2706,N_2404);
nand UO_194 (O_194,N_2557,N_2916);
or UO_195 (O_195,N_2149,N_2215);
or UO_196 (O_196,N_2556,N_2069);
xnor UO_197 (O_197,N_2626,N_2192);
xor UO_198 (O_198,N_2586,N_2796);
or UO_199 (O_199,N_2109,N_2105);
nor UO_200 (O_200,N_2934,N_2186);
and UO_201 (O_201,N_2337,N_2816);
or UO_202 (O_202,N_2757,N_2430);
and UO_203 (O_203,N_2566,N_2630);
and UO_204 (O_204,N_2569,N_2892);
or UO_205 (O_205,N_2458,N_2717);
xnor UO_206 (O_206,N_2025,N_2078);
or UO_207 (O_207,N_2261,N_2461);
and UO_208 (O_208,N_2616,N_2583);
nor UO_209 (O_209,N_2044,N_2219);
nand UO_210 (O_210,N_2083,N_2361);
or UO_211 (O_211,N_2754,N_2740);
nor UO_212 (O_212,N_2930,N_2611);
or UO_213 (O_213,N_2967,N_2938);
nor UO_214 (O_214,N_2684,N_2558);
xor UO_215 (O_215,N_2277,N_2925);
xnor UO_216 (O_216,N_2783,N_2988);
xor UO_217 (O_217,N_2019,N_2546);
nor UO_218 (O_218,N_2663,N_2071);
xor UO_219 (O_219,N_2529,N_2313);
or UO_220 (O_220,N_2155,N_2895);
nand UO_221 (O_221,N_2243,N_2336);
and UO_222 (O_222,N_2522,N_2456);
and UO_223 (O_223,N_2992,N_2130);
nor UO_224 (O_224,N_2203,N_2932);
nor UO_225 (O_225,N_2153,N_2402);
or UO_226 (O_226,N_2004,N_2254);
nand UO_227 (O_227,N_2951,N_2943);
and UO_228 (O_228,N_2819,N_2613);
nor UO_229 (O_229,N_2861,N_2731);
and UO_230 (O_230,N_2654,N_2701);
or UO_231 (O_231,N_2773,N_2407);
nand UO_232 (O_232,N_2082,N_2787);
nand UO_233 (O_233,N_2500,N_2917);
nand UO_234 (O_234,N_2444,N_2176);
or UO_235 (O_235,N_2443,N_2532);
and UO_236 (O_236,N_2131,N_2718);
and UO_237 (O_237,N_2183,N_2878);
nor UO_238 (O_238,N_2933,N_2395);
and UO_239 (O_239,N_2523,N_2010);
xnor UO_240 (O_240,N_2180,N_2079);
xor UO_241 (O_241,N_2333,N_2669);
or UO_242 (O_242,N_2741,N_2428);
xor UO_243 (O_243,N_2258,N_2609);
nand UO_244 (O_244,N_2983,N_2191);
and UO_245 (O_245,N_2204,N_2968);
nor UO_246 (O_246,N_2245,N_2520);
nor UO_247 (O_247,N_2574,N_2966);
nor UO_248 (O_248,N_2929,N_2324);
nor UO_249 (O_249,N_2513,N_2158);
nand UO_250 (O_250,N_2894,N_2673);
nand UO_251 (O_251,N_2622,N_2801);
and UO_252 (O_252,N_2314,N_2009);
nand UO_253 (O_253,N_2592,N_2882);
nor UO_254 (O_254,N_2159,N_2947);
nand UO_255 (O_255,N_2866,N_2497);
or UO_256 (O_256,N_2392,N_2971);
nand UO_257 (O_257,N_2792,N_2393);
or UO_258 (O_258,N_2289,N_2752);
or UO_259 (O_259,N_2438,N_2538);
nor UO_260 (O_260,N_2136,N_2914);
nor UO_261 (O_261,N_2660,N_2949);
xnor UO_262 (O_262,N_2828,N_2340);
nand UO_263 (O_263,N_2031,N_2856);
or UO_264 (O_264,N_2409,N_2786);
and UO_265 (O_265,N_2981,N_2214);
nor UO_266 (O_266,N_2824,N_2573);
and UO_267 (O_267,N_2931,N_2175);
nor UO_268 (O_268,N_2509,N_2086);
xor UO_269 (O_269,N_2033,N_2052);
nor UO_270 (O_270,N_2503,N_2150);
and UO_271 (O_271,N_2420,N_2771);
nor UO_272 (O_272,N_2166,N_2817);
and UO_273 (O_273,N_2474,N_2276);
and UO_274 (O_274,N_2991,N_2802);
and UO_275 (O_275,N_2036,N_2617);
nor UO_276 (O_276,N_2698,N_2471);
and UO_277 (O_277,N_2397,N_2473);
and UO_278 (O_278,N_2857,N_2807);
nor UO_279 (O_279,N_2849,N_2264);
nand UO_280 (O_280,N_2411,N_2058);
xnor UO_281 (O_281,N_2832,N_2571);
xor UO_282 (O_282,N_2432,N_2738);
nand UO_283 (O_283,N_2541,N_2135);
or UO_284 (O_284,N_2378,N_2593);
nor UO_285 (O_285,N_2330,N_2575);
nand UO_286 (O_286,N_2760,N_2049);
and UO_287 (O_287,N_2063,N_2329);
or UO_288 (O_288,N_2106,N_2872);
and UO_289 (O_289,N_2788,N_2413);
or UO_290 (O_290,N_2207,N_2275);
or UO_291 (O_291,N_2870,N_2244);
or UO_292 (O_292,N_2785,N_2564);
nor UO_293 (O_293,N_2733,N_2373);
or UO_294 (O_294,N_2521,N_2743);
nor UO_295 (O_295,N_2440,N_2537);
or UO_296 (O_296,N_2138,N_2634);
xnor UO_297 (O_297,N_2904,N_2479);
or UO_298 (O_298,N_2962,N_2887);
or UO_299 (O_299,N_2094,N_2552);
nand UO_300 (O_300,N_2399,N_2923);
and UO_301 (O_301,N_2686,N_2772);
or UO_302 (O_302,N_2745,N_2120);
xnor UO_303 (O_303,N_2029,N_2198);
and UO_304 (O_304,N_2113,N_2524);
and UO_305 (O_305,N_2043,N_2469);
nand UO_306 (O_306,N_2374,N_2041);
or UO_307 (O_307,N_2065,N_2000);
nand UO_308 (O_308,N_2221,N_2768);
or UO_309 (O_309,N_2103,N_2385);
xnor UO_310 (O_310,N_2628,N_2668);
or UO_311 (O_311,N_2391,N_2514);
xor UO_312 (O_312,N_2900,N_2598);
nor UO_313 (O_313,N_2338,N_2875);
and UO_314 (O_314,N_2863,N_2506);
xor UO_315 (O_315,N_2181,N_2636);
nand UO_316 (O_316,N_2358,N_2905);
and UO_317 (O_317,N_2848,N_2724);
or UO_318 (O_318,N_2346,N_2257);
nand UO_319 (O_319,N_2952,N_2794);
and UO_320 (O_320,N_2779,N_2101);
and UO_321 (O_321,N_2753,N_2906);
nand UO_322 (O_322,N_2650,N_2016);
or UO_323 (O_323,N_2946,N_2913);
nor UO_324 (O_324,N_2050,N_2344);
nor UO_325 (O_325,N_2890,N_2582);
nor UO_326 (O_326,N_2209,N_2098);
nand UO_327 (O_327,N_2061,N_2156);
nand UO_328 (O_328,N_2633,N_2507);
nand UO_329 (O_329,N_2481,N_2160);
and UO_330 (O_330,N_2076,N_2734);
and UO_331 (O_331,N_2173,N_2618);
nor UO_332 (O_332,N_2305,N_2108);
nand UO_333 (O_333,N_2818,N_2498);
nor UO_334 (O_334,N_2591,N_2587);
or UO_335 (O_335,N_2462,N_2704);
nand UO_336 (O_336,N_2543,N_2811);
nor UO_337 (O_337,N_2637,N_2687);
or UO_338 (O_338,N_2268,N_2735);
nand UO_339 (O_339,N_2188,N_2349);
or UO_340 (O_340,N_2172,N_2798);
nor UO_341 (O_341,N_2831,N_2366);
nand UO_342 (O_342,N_2889,N_2343);
and UO_343 (O_343,N_2433,N_2217);
nand UO_344 (O_344,N_2454,N_2809);
nor UO_345 (O_345,N_2353,N_2425);
xnor UO_346 (O_346,N_2542,N_2253);
or UO_347 (O_347,N_2563,N_2003);
and UO_348 (O_348,N_2496,N_2072);
nand UO_349 (O_349,N_2075,N_2246);
or UO_350 (O_350,N_2674,N_2899);
nor UO_351 (O_351,N_2088,N_2077);
xor UO_352 (O_352,N_2376,N_2539);
nand UO_353 (O_353,N_2782,N_2791);
and UO_354 (O_354,N_2302,N_2417);
nand UO_355 (O_355,N_2813,N_2528);
or UO_356 (O_356,N_2062,N_2394);
nor UO_357 (O_357,N_2423,N_2354);
or UO_358 (O_358,N_2780,N_2384);
nor UO_359 (O_359,N_2722,N_2612);
or UO_360 (O_360,N_2042,N_2012);
nor UO_361 (O_361,N_2431,N_2196);
and UO_362 (O_362,N_2424,N_2226);
nand UO_363 (O_363,N_2024,N_2267);
or UO_364 (O_364,N_2383,N_2559);
nand UO_365 (O_365,N_2972,N_2291);
and UO_366 (O_366,N_2288,N_2948);
and UO_367 (O_367,N_2996,N_2719);
or UO_368 (O_368,N_2017,N_2826);
nor UO_369 (O_369,N_2477,N_2536);
and UO_370 (O_370,N_2620,N_2578);
and UO_371 (O_371,N_2936,N_2332);
and UO_372 (O_372,N_2652,N_2781);
or UO_373 (O_373,N_2920,N_2247);
or UO_374 (O_374,N_2287,N_2242);
and UO_375 (O_375,N_2619,N_2309);
nor UO_376 (O_376,N_2294,N_2545);
and UO_377 (O_377,N_2980,N_2119);
and UO_378 (O_378,N_2661,N_2452);
xor UO_379 (O_379,N_2727,N_2963);
nand UO_380 (O_380,N_2260,N_2168);
nor UO_381 (O_381,N_2517,N_2381);
nor UO_382 (O_382,N_2446,N_2266);
nor UO_383 (O_383,N_2490,N_2252);
or UO_384 (O_384,N_2624,N_2111);
nor UO_385 (O_385,N_2115,N_2127);
xor UO_386 (O_386,N_2868,N_2867);
nand UO_387 (O_387,N_2576,N_2790);
nand UO_388 (O_388,N_2070,N_2053);
and UO_389 (O_389,N_2648,N_2295);
and UO_390 (O_390,N_2838,N_2421);
and UO_391 (O_391,N_2216,N_2835);
nand UO_392 (O_392,N_2321,N_2464);
nor UO_393 (O_393,N_2501,N_2697);
or UO_394 (O_394,N_2026,N_2911);
and UO_395 (O_395,N_2860,N_2632);
nand UO_396 (O_396,N_2020,N_2775);
and UO_397 (O_397,N_2484,N_2885);
or UO_398 (O_398,N_2485,N_2742);
and UO_399 (O_399,N_2355,N_2161);
nand UO_400 (O_400,N_2806,N_2845);
xor UO_401 (O_401,N_2820,N_2827);
nand UO_402 (O_402,N_2713,N_2401);
nand UO_403 (O_403,N_2434,N_2994);
or UO_404 (O_404,N_2128,N_2682);
nand UO_405 (O_405,N_2627,N_2960);
or UO_406 (O_406,N_2369,N_2671);
nand UO_407 (O_407,N_2737,N_2426);
xnor UO_408 (O_408,N_2855,N_2884);
and UO_409 (O_409,N_2145,N_2847);
nor UO_410 (O_410,N_2789,N_2815);
and UO_411 (O_411,N_2935,N_2193);
nand UO_412 (O_412,N_2396,N_2693);
and UO_413 (O_413,N_2449,N_2367);
or UO_414 (O_414,N_2205,N_2230);
or UO_415 (O_415,N_2865,N_2398);
nor UO_416 (O_416,N_2761,N_2304);
nor UO_417 (O_417,N_2511,N_2200);
and UO_418 (O_418,N_2074,N_2296);
or UO_419 (O_419,N_2527,N_2189);
nand UO_420 (O_420,N_2615,N_2486);
and UO_421 (O_421,N_2728,N_2475);
nand UO_422 (O_422,N_2750,N_2427);
or UO_423 (O_423,N_2664,N_2965);
nor UO_424 (O_424,N_2104,N_2418);
and UO_425 (O_425,N_2502,N_2958);
xor UO_426 (O_426,N_2278,N_2610);
or UO_427 (O_427,N_2182,N_2915);
nor UO_428 (O_428,N_2647,N_2001);
and UO_429 (O_429,N_2912,N_2600);
and UO_430 (O_430,N_2080,N_2602);
nor UO_431 (O_431,N_2487,N_2139);
and UO_432 (O_432,N_2989,N_2137);
nand UO_433 (O_433,N_2803,N_2459);
and UO_434 (O_434,N_2909,N_2008);
and UO_435 (O_435,N_2638,N_2519);
xnor UO_436 (O_436,N_2764,N_2084);
or UO_437 (O_437,N_2334,N_2584);
xor UO_438 (O_438,N_2414,N_2653);
nor UO_439 (O_439,N_2945,N_2335);
nor UO_440 (O_440,N_2092,N_2045);
or UO_441 (O_441,N_2201,N_2560);
or UO_442 (O_442,N_2864,N_2964);
nand UO_443 (O_443,N_2777,N_2482);
and UO_444 (O_444,N_2489,N_2112);
nor UO_445 (O_445,N_2880,N_2239);
nand UO_446 (O_446,N_2318,N_2312);
and UO_447 (O_447,N_2081,N_2561);
and UO_448 (O_448,N_2893,N_2048);
nor UO_449 (O_449,N_2248,N_2339);
nor UO_450 (O_450,N_2723,N_2969);
nor UO_451 (O_451,N_2927,N_2830);
nand UO_452 (O_452,N_2491,N_2142);
nor UO_453 (O_453,N_2984,N_2683);
xnor UO_454 (O_454,N_2235,N_2472);
nand UO_455 (O_455,N_2721,N_2709);
or UO_456 (O_456,N_2362,N_2164);
nand UO_457 (O_457,N_2516,N_2348);
nor UO_458 (O_458,N_2364,N_2579);
and UO_459 (O_459,N_2095,N_2937);
nand UO_460 (O_460,N_2805,N_2184);
and UO_461 (O_461,N_2368,N_2554);
nor UO_462 (O_462,N_2125,N_2715);
nor UO_463 (O_463,N_2370,N_2499);
or UO_464 (O_464,N_2379,N_2700);
nand UO_465 (O_465,N_2979,N_2013);
and UO_466 (O_466,N_2510,N_2297);
xor UO_467 (O_467,N_2982,N_2124);
nor UO_468 (O_468,N_2389,N_2758);
or UO_469 (O_469,N_2921,N_2441);
and UO_470 (O_470,N_2874,N_2165);
or UO_471 (O_471,N_2263,N_2685);
and UO_472 (O_472,N_2281,N_2858);
and UO_473 (O_473,N_2493,N_2005);
or UO_474 (O_474,N_2096,N_2451);
nor UO_475 (O_475,N_2320,N_2178);
nor UO_476 (O_476,N_2975,N_2732);
nand UO_477 (O_477,N_2350,N_2271);
xor UO_478 (O_478,N_2720,N_2460);
or UO_479 (O_479,N_2707,N_2195);
nor UO_480 (O_480,N_2504,N_2416);
or UO_481 (O_481,N_2056,N_2808);
or UO_482 (O_482,N_2670,N_2903);
or UO_483 (O_483,N_2763,N_2941);
or UO_484 (O_484,N_2476,N_2842);
xor UO_485 (O_485,N_2730,N_2987);
nor UO_486 (O_486,N_2590,N_2319);
nor UO_487 (O_487,N_2585,N_2548);
nand UO_488 (O_488,N_2762,N_2406);
and UO_489 (O_489,N_2177,N_2770);
and UO_490 (O_490,N_2690,N_2705);
or UO_491 (O_491,N_2508,N_2599);
nand UO_492 (O_492,N_2844,N_2621);
and UO_493 (O_493,N_2229,N_2944);
or UO_494 (O_494,N_2853,N_2495);
or UO_495 (O_495,N_2327,N_2840);
and UO_496 (O_496,N_2419,N_2365);
or UO_497 (O_497,N_2877,N_2060);
nand UO_498 (O_498,N_2467,N_2572);
and UO_499 (O_499,N_2371,N_2238);
endmodule