module basic_500_3000_500_6_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_89,In_219);
or U1 (N_1,In_128,In_134);
or U2 (N_2,In_409,In_77);
or U3 (N_3,In_343,In_179);
nor U4 (N_4,In_490,In_416);
or U5 (N_5,In_55,In_363);
or U6 (N_6,In_370,In_160);
xor U7 (N_7,In_58,In_329);
nor U8 (N_8,In_262,In_478);
and U9 (N_9,In_441,In_492);
nand U10 (N_10,In_308,In_342);
nor U11 (N_11,In_309,In_136);
nand U12 (N_12,In_265,In_210);
nand U13 (N_13,In_222,In_93);
nor U14 (N_14,In_379,In_479);
and U15 (N_15,In_291,In_203);
and U16 (N_16,In_372,In_458);
xnor U17 (N_17,In_350,In_72);
or U18 (N_18,In_383,In_239);
or U19 (N_19,In_75,In_378);
nand U20 (N_20,In_74,In_231);
nand U21 (N_21,In_420,In_322);
nor U22 (N_22,In_86,In_387);
or U23 (N_23,In_155,In_169);
and U24 (N_24,In_389,In_116);
nand U25 (N_25,In_402,In_170);
nand U26 (N_26,In_401,In_137);
or U27 (N_27,In_192,In_76);
nand U28 (N_28,In_419,In_284);
nor U29 (N_29,In_319,In_288);
or U30 (N_30,In_277,In_23);
nor U31 (N_31,In_359,In_330);
and U32 (N_32,In_424,In_158);
nor U33 (N_33,In_421,In_323);
or U34 (N_34,In_146,In_19);
and U35 (N_35,In_122,In_166);
and U36 (N_36,In_295,In_235);
and U37 (N_37,In_272,In_446);
nor U38 (N_38,In_285,In_392);
nor U39 (N_39,In_448,In_127);
and U40 (N_40,In_119,In_242);
nor U41 (N_41,In_199,In_292);
or U42 (N_42,In_436,In_17);
nor U43 (N_43,In_324,In_220);
or U44 (N_44,In_394,In_261);
nand U45 (N_45,In_167,In_123);
nor U46 (N_46,In_404,In_298);
nand U47 (N_47,In_150,In_37);
nor U48 (N_48,In_42,In_488);
or U49 (N_49,In_108,In_70);
or U50 (N_50,In_278,In_29);
and U51 (N_51,In_484,In_443);
or U52 (N_52,In_321,In_354);
nor U53 (N_53,In_230,In_18);
nor U54 (N_54,In_112,In_467);
or U55 (N_55,In_398,In_346);
nor U56 (N_56,In_105,In_333);
and U57 (N_57,In_302,In_24);
nand U58 (N_58,In_294,In_53);
nor U59 (N_59,In_460,In_51);
and U60 (N_60,In_229,In_491);
xor U61 (N_61,In_362,In_264);
nor U62 (N_62,In_84,In_426);
nand U63 (N_63,In_205,In_463);
and U64 (N_64,In_190,In_52);
nor U65 (N_65,In_133,In_87);
nor U66 (N_66,In_139,In_297);
or U67 (N_67,In_412,In_117);
and U68 (N_68,In_109,In_14);
xor U69 (N_69,In_400,In_258);
nor U70 (N_70,In_151,In_188);
xor U71 (N_71,In_369,In_431);
xor U72 (N_72,In_198,In_396);
nor U73 (N_73,In_191,In_260);
and U74 (N_74,In_341,In_252);
xor U75 (N_75,In_444,In_9);
or U76 (N_76,In_279,In_131);
nor U77 (N_77,In_227,In_32);
nand U78 (N_78,In_493,In_355);
nand U79 (N_79,In_358,In_481);
xnor U80 (N_80,In_327,In_245);
and U81 (N_81,In_480,In_223);
or U82 (N_82,In_339,In_111);
xnor U83 (N_83,In_263,In_445);
nand U84 (N_84,In_451,In_73);
nand U85 (N_85,In_499,In_33);
nor U86 (N_86,In_225,In_152);
and U87 (N_87,In_442,In_215);
or U88 (N_88,In_187,In_120);
or U89 (N_89,In_345,In_254);
xnor U90 (N_90,In_386,In_332);
nand U91 (N_91,In_54,In_38);
nand U92 (N_92,In_410,In_382);
or U93 (N_93,In_331,In_20);
and U94 (N_94,In_209,In_453);
nand U95 (N_95,In_224,In_440);
or U96 (N_96,In_197,In_124);
or U97 (N_97,In_142,In_79);
or U98 (N_98,In_381,In_282);
nor U99 (N_99,In_59,In_154);
nor U100 (N_100,In_41,In_96);
nor U101 (N_101,In_161,In_301);
nor U102 (N_102,In_312,In_476);
nand U103 (N_103,In_184,In_30);
nand U104 (N_104,In_320,In_328);
nor U105 (N_105,In_256,In_100);
nand U106 (N_106,In_449,In_408);
nor U107 (N_107,In_240,In_290);
nor U108 (N_108,In_65,In_374);
nor U109 (N_109,In_45,In_496);
and U110 (N_110,In_39,In_438);
nor U111 (N_111,In_360,In_454);
and U112 (N_112,In_44,In_99);
or U113 (N_113,In_405,In_300);
nor U114 (N_114,In_106,In_34);
and U115 (N_115,In_450,In_182);
nor U116 (N_116,In_201,In_94);
and U117 (N_117,In_35,In_406);
and U118 (N_118,In_218,In_418);
xnor U119 (N_119,In_248,In_266);
nor U120 (N_120,In_395,In_174);
or U121 (N_121,In_207,In_299);
nor U122 (N_122,In_121,In_101);
nor U123 (N_123,In_21,In_125);
or U124 (N_124,In_439,In_306);
nor U125 (N_125,In_283,In_233);
nand U126 (N_126,In_64,In_16);
nand U127 (N_127,In_457,In_415);
nand U128 (N_128,In_271,In_376);
and U129 (N_129,In_67,In_391);
nor U130 (N_130,In_384,In_307);
or U131 (N_131,In_335,In_472);
xnor U132 (N_132,In_1,In_114);
or U133 (N_133,In_465,In_255);
nand U134 (N_134,In_81,In_62);
xor U135 (N_135,In_364,In_243);
nor U136 (N_136,In_238,In_474);
nor U137 (N_137,In_115,In_336);
or U138 (N_138,In_165,In_303);
xor U139 (N_139,In_138,In_482);
and U140 (N_140,In_148,In_25);
nand U141 (N_141,In_82,In_206);
nor U142 (N_142,In_36,In_311);
nand U143 (N_143,In_429,In_173);
nand U144 (N_144,In_456,In_390);
nand U145 (N_145,In_226,In_293);
nand U146 (N_146,In_305,In_68);
and U147 (N_147,In_175,In_3);
and U148 (N_148,In_494,In_90);
and U149 (N_149,In_437,In_334);
nand U150 (N_150,In_428,In_462);
nand U151 (N_151,In_126,In_353);
and U152 (N_152,In_434,In_13);
nand U153 (N_153,In_464,In_236);
nand U154 (N_154,In_221,In_407);
nand U155 (N_155,In_97,In_489);
nor U156 (N_156,In_10,In_194);
xor U157 (N_157,In_399,In_373);
nor U158 (N_158,In_27,In_276);
nor U159 (N_159,In_352,In_183);
xor U160 (N_160,In_71,In_447);
xor U161 (N_161,In_251,In_275);
and U162 (N_162,In_403,In_417);
or U163 (N_163,In_193,In_459);
nand U164 (N_164,In_286,In_473);
xnor U165 (N_165,In_104,In_157);
and U166 (N_166,In_316,In_241);
and U167 (N_167,In_56,In_356);
nor U168 (N_168,In_469,In_107);
nor U169 (N_169,In_162,In_228);
nor U170 (N_170,In_274,In_287);
nand U171 (N_171,In_200,In_31);
nor U172 (N_172,In_347,In_171);
or U173 (N_173,In_326,In_344);
or U174 (N_174,In_185,In_348);
and U175 (N_175,In_313,In_164);
nor U176 (N_176,In_69,In_366);
nand U177 (N_177,In_430,In_6);
or U178 (N_178,In_61,In_377);
or U179 (N_179,In_361,In_181);
nand U180 (N_180,In_317,In_246);
or U181 (N_181,In_296,In_318);
nor U182 (N_182,In_273,In_135);
and U183 (N_183,In_98,In_118);
and U184 (N_184,In_83,In_351);
or U185 (N_185,In_43,In_85);
and U186 (N_186,In_140,In_195);
nand U187 (N_187,In_466,In_48);
or U188 (N_188,In_189,In_211);
or U189 (N_189,In_314,In_393);
nor U190 (N_190,In_145,In_397);
nor U191 (N_191,In_47,In_132);
nand U192 (N_192,In_92,In_470);
nor U193 (N_193,In_214,In_337);
nor U194 (N_194,In_80,In_15);
and U195 (N_195,In_7,In_249);
nand U196 (N_196,In_423,In_253);
nand U197 (N_197,In_113,In_259);
nor U198 (N_198,In_267,In_497);
nor U199 (N_199,In_176,In_186);
and U200 (N_200,In_22,In_78);
xor U201 (N_201,In_60,In_422);
and U202 (N_202,In_2,In_427);
xnor U203 (N_203,In_365,In_216);
nand U204 (N_204,In_88,In_204);
or U205 (N_205,In_141,In_483);
xnor U206 (N_206,In_433,In_178);
nand U207 (N_207,In_367,In_163);
or U208 (N_208,In_237,In_232);
nand U209 (N_209,In_315,In_310);
nor U210 (N_210,In_495,In_468);
or U211 (N_211,In_143,In_177);
xnor U212 (N_212,In_63,In_349);
or U213 (N_213,In_234,In_172);
or U214 (N_214,In_461,In_66);
nand U215 (N_215,In_357,In_385);
xnor U216 (N_216,In_50,In_477);
nor U217 (N_217,In_486,In_244);
nor U218 (N_218,In_338,In_11);
and U219 (N_219,In_435,In_180);
and U220 (N_220,In_270,In_487);
and U221 (N_221,In_485,In_8);
or U222 (N_222,In_103,In_281);
nor U223 (N_223,In_208,In_91);
and U224 (N_224,In_95,In_153);
nor U225 (N_225,In_168,In_250);
or U226 (N_226,In_257,In_325);
and U227 (N_227,In_452,In_110);
and U228 (N_228,In_471,In_388);
nor U229 (N_229,In_475,In_217);
and U230 (N_230,In_413,In_130);
and U231 (N_231,In_46,In_149);
nand U232 (N_232,In_455,In_156);
nand U233 (N_233,In_371,In_432);
xor U234 (N_234,In_380,In_414);
nand U235 (N_235,In_268,In_5);
nand U236 (N_236,In_102,In_28);
xor U237 (N_237,In_40,In_498);
xor U238 (N_238,In_247,In_411);
and U239 (N_239,In_368,In_26);
nor U240 (N_240,In_269,In_159);
and U241 (N_241,In_202,In_289);
and U242 (N_242,In_212,In_0);
and U243 (N_243,In_213,In_375);
and U244 (N_244,In_340,In_4);
nor U245 (N_245,In_425,In_147);
xor U246 (N_246,In_304,In_49);
xor U247 (N_247,In_280,In_144);
xnor U248 (N_248,In_12,In_129);
nor U249 (N_249,In_196,In_57);
or U250 (N_250,In_348,In_202);
nand U251 (N_251,In_420,In_253);
or U252 (N_252,In_35,In_172);
and U253 (N_253,In_237,In_179);
nor U254 (N_254,In_140,In_183);
nand U255 (N_255,In_345,In_170);
and U256 (N_256,In_356,In_335);
xor U257 (N_257,In_176,In_315);
nand U258 (N_258,In_214,In_420);
nand U259 (N_259,In_45,In_146);
nand U260 (N_260,In_375,In_338);
nor U261 (N_261,In_33,In_114);
nor U262 (N_262,In_458,In_325);
xnor U263 (N_263,In_121,In_63);
and U264 (N_264,In_220,In_159);
or U265 (N_265,In_170,In_369);
nand U266 (N_266,In_402,In_87);
xor U267 (N_267,In_88,In_271);
and U268 (N_268,In_38,In_276);
nor U269 (N_269,In_99,In_399);
xnor U270 (N_270,In_57,In_490);
nor U271 (N_271,In_106,In_24);
and U272 (N_272,In_176,In_362);
and U273 (N_273,In_457,In_472);
and U274 (N_274,In_88,In_58);
and U275 (N_275,In_492,In_72);
or U276 (N_276,In_35,In_228);
nand U277 (N_277,In_44,In_481);
nand U278 (N_278,In_34,In_288);
nor U279 (N_279,In_363,In_482);
or U280 (N_280,In_455,In_443);
or U281 (N_281,In_338,In_332);
xnor U282 (N_282,In_327,In_277);
xor U283 (N_283,In_487,In_124);
nor U284 (N_284,In_116,In_378);
nor U285 (N_285,In_104,In_492);
or U286 (N_286,In_67,In_279);
or U287 (N_287,In_247,In_466);
or U288 (N_288,In_107,In_446);
nor U289 (N_289,In_413,In_180);
nor U290 (N_290,In_130,In_235);
and U291 (N_291,In_7,In_247);
and U292 (N_292,In_434,In_455);
nor U293 (N_293,In_241,In_462);
or U294 (N_294,In_483,In_24);
or U295 (N_295,In_422,In_319);
xor U296 (N_296,In_281,In_47);
nor U297 (N_297,In_303,In_400);
nand U298 (N_298,In_209,In_99);
nand U299 (N_299,In_297,In_459);
nor U300 (N_300,In_456,In_190);
nor U301 (N_301,In_404,In_148);
and U302 (N_302,In_32,In_35);
xnor U303 (N_303,In_223,In_485);
and U304 (N_304,In_423,In_205);
xnor U305 (N_305,In_116,In_223);
and U306 (N_306,In_301,In_381);
nor U307 (N_307,In_177,In_428);
or U308 (N_308,In_388,In_400);
nor U309 (N_309,In_454,In_447);
and U310 (N_310,In_33,In_474);
nor U311 (N_311,In_98,In_261);
nor U312 (N_312,In_401,In_435);
nand U313 (N_313,In_361,In_119);
and U314 (N_314,In_460,In_201);
nand U315 (N_315,In_451,In_208);
nor U316 (N_316,In_474,In_389);
or U317 (N_317,In_205,In_227);
or U318 (N_318,In_382,In_173);
nor U319 (N_319,In_35,In_443);
and U320 (N_320,In_455,In_220);
or U321 (N_321,In_19,In_498);
or U322 (N_322,In_105,In_106);
nor U323 (N_323,In_493,In_332);
and U324 (N_324,In_105,In_423);
xor U325 (N_325,In_450,In_274);
xnor U326 (N_326,In_319,In_483);
xor U327 (N_327,In_257,In_53);
xor U328 (N_328,In_188,In_309);
nand U329 (N_329,In_72,In_353);
and U330 (N_330,In_343,In_334);
and U331 (N_331,In_331,In_296);
xor U332 (N_332,In_277,In_14);
nand U333 (N_333,In_359,In_127);
nor U334 (N_334,In_64,In_383);
or U335 (N_335,In_271,In_35);
or U336 (N_336,In_455,In_301);
nand U337 (N_337,In_239,In_149);
or U338 (N_338,In_34,In_322);
and U339 (N_339,In_390,In_348);
or U340 (N_340,In_462,In_423);
and U341 (N_341,In_324,In_144);
and U342 (N_342,In_155,In_493);
nor U343 (N_343,In_130,In_18);
nor U344 (N_344,In_456,In_152);
or U345 (N_345,In_428,In_397);
and U346 (N_346,In_258,In_177);
and U347 (N_347,In_158,In_429);
nor U348 (N_348,In_74,In_101);
and U349 (N_349,In_346,In_77);
or U350 (N_350,In_487,In_423);
xor U351 (N_351,In_342,In_444);
or U352 (N_352,In_438,In_496);
nand U353 (N_353,In_153,In_16);
nand U354 (N_354,In_288,In_327);
nor U355 (N_355,In_306,In_20);
nor U356 (N_356,In_484,In_200);
nor U357 (N_357,In_1,In_275);
and U358 (N_358,In_416,In_491);
xnor U359 (N_359,In_487,In_317);
nand U360 (N_360,In_28,In_158);
nand U361 (N_361,In_308,In_144);
and U362 (N_362,In_408,In_359);
and U363 (N_363,In_24,In_70);
xor U364 (N_364,In_110,In_303);
nor U365 (N_365,In_35,In_154);
or U366 (N_366,In_166,In_425);
xnor U367 (N_367,In_406,In_336);
xor U368 (N_368,In_376,In_439);
nor U369 (N_369,In_454,In_314);
xor U370 (N_370,In_468,In_459);
and U371 (N_371,In_452,In_97);
or U372 (N_372,In_404,In_26);
xnor U373 (N_373,In_156,In_118);
nand U374 (N_374,In_497,In_17);
nand U375 (N_375,In_89,In_168);
and U376 (N_376,In_123,In_378);
nand U377 (N_377,In_189,In_42);
or U378 (N_378,In_181,In_90);
nand U379 (N_379,In_243,In_493);
nand U380 (N_380,In_339,In_44);
nor U381 (N_381,In_167,In_341);
nand U382 (N_382,In_122,In_79);
xnor U383 (N_383,In_179,In_418);
nor U384 (N_384,In_56,In_220);
nand U385 (N_385,In_459,In_165);
and U386 (N_386,In_252,In_478);
and U387 (N_387,In_63,In_453);
nor U388 (N_388,In_55,In_4);
nand U389 (N_389,In_162,In_342);
nand U390 (N_390,In_327,In_316);
xor U391 (N_391,In_215,In_431);
nand U392 (N_392,In_188,In_49);
or U393 (N_393,In_296,In_451);
or U394 (N_394,In_340,In_293);
nand U395 (N_395,In_293,In_311);
and U396 (N_396,In_334,In_57);
nor U397 (N_397,In_137,In_287);
or U398 (N_398,In_29,In_429);
nand U399 (N_399,In_288,In_486);
xor U400 (N_400,In_63,In_254);
or U401 (N_401,In_440,In_142);
and U402 (N_402,In_418,In_97);
nor U403 (N_403,In_437,In_92);
or U404 (N_404,In_222,In_64);
xnor U405 (N_405,In_303,In_447);
nor U406 (N_406,In_103,In_400);
nor U407 (N_407,In_162,In_245);
xor U408 (N_408,In_20,In_141);
nor U409 (N_409,In_429,In_208);
or U410 (N_410,In_89,In_231);
and U411 (N_411,In_267,In_181);
nand U412 (N_412,In_407,In_428);
nor U413 (N_413,In_179,In_59);
nor U414 (N_414,In_180,In_386);
and U415 (N_415,In_245,In_239);
nand U416 (N_416,In_481,In_390);
and U417 (N_417,In_302,In_445);
nor U418 (N_418,In_297,In_386);
xnor U419 (N_419,In_452,In_223);
nand U420 (N_420,In_205,In_57);
nor U421 (N_421,In_220,In_416);
nand U422 (N_422,In_465,In_267);
nand U423 (N_423,In_190,In_95);
nor U424 (N_424,In_424,In_360);
or U425 (N_425,In_470,In_34);
and U426 (N_426,In_36,In_113);
or U427 (N_427,In_264,In_405);
or U428 (N_428,In_214,In_73);
and U429 (N_429,In_70,In_8);
nand U430 (N_430,In_218,In_326);
or U431 (N_431,In_119,In_372);
or U432 (N_432,In_319,In_304);
and U433 (N_433,In_86,In_228);
and U434 (N_434,In_304,In_72);
nand U435 (N_435,In_72,In_12);
xor U436 (N_436,In_447,In_163);
nand U437 (N_437,In_55,In_347);
or U438 (N_438,In_62,In_34);
and U439 (N_439,In_25,In_196);
nand U440 (N_440,In_159,In_65);
nand U441 (N_441,In_422,In_280);
and U442 (N_442,In_210,In_104);
xor U443 (N_443,In_297,In_404);
nand U444 (N_444,In_72,In_298);
and U445 (N_445,In_410,In_428);
nand U446 (N_446,In_432,In_240);
nor U447 (N_447,In_242,In_296);
nand U448 (N_448,In_210,In_410);
nor U449 (N_449,In_107,In_65);
nor U450 (N_450,In_76,In_79);
nor U451 (N_451,In_161,In_66);
nand U452 (N_452,In_52,In_411);
and U453 (N_453,In_374,In_407);
or U454 (N_454,In_138,In_187);
xnor U455 (N_455,In_308,In_253);
nor U456 (N_456,In_6,In_148);
nor U457 (N_457,In_104,In_141);
and U458 (N_458,In_27,In_17);
and U459 (N_459,In_454,In_436);
nor U460 (N_460,In_301,In_406);
nor U461 (N_461,In_124,In_457);
or U462 (N_462,In_161,In_130);
nor U463 (N_463,In_392,In_72);
and U464 (N_464,In_379,In_390);
or U465 (N_465,In_82,In_64);
nand U466 (N_466,In_5,In_499);
and U467 (N_467,In_400,In_232);
nor U468 (N_468,In_4,In_53);
nand U469 (N_469,In_403,In_162);
nor U470 (N_470,In_242,In_496);
xnor U471 (N_471,In_340,In_438);
xnor U472 (N_472,In_65,In_36);
nand U473 (N_473,In_344,In_306);
nor U474 (N_474,In_373,In_352);
or U475 (N_475,In_225,In_367);
xnor U476 (N_476,In_374,In_19);
or U477 (N_477,In_388,In_408);
nor U478 (N_478,In_284,In_321);
xnor U479 (N_479,In_274,In_215);
and U480 (N_480,In_57,In_55);
and U481 (N_481,In_370,In_80);
and U482 (N_482,In_70,In_260);
nor U483 (N_483,In_261,In_142);
xor U484 (N_484,In_45,In_429);
nor U485 (N_485,In_429,In_481);
or U486 (N_486,In_125,In_235);
or U487 (N_487,In_45,In_6);
or U488 (N_488,In_485,In_203);
nor U489 (N_489,In_120,In_115);
nand U490 (N_490,In_79,In_342);
nor U491 (N_491,In_44,In_194);
or U492 (N_492,In_42,In_352);
or U493 (N_493,In_36,In_150);
or U494 (N_494,In_362,In_169);
or U495 (N_495,In_135,In_299);
nand U496 (N_496,In_370,In_48);
and U497 (N_497,In_212,In_437);
nand U498 (N_498,In_401,In_394);
or U499 (N_499,In_74,In_108);
nand U500 (N_500,N_350,N_13);
or U501 (N_501,N_311,N_246);
xor U502 (N_502,N_136,N_194);
nand U503 (N_503,N_11,N_305);
nor U504 (N_504,N_145,N_54);
and U505 (N_505,N_129,N_81);
or U506 (N_506,N_21,N_118);
xor U507 (N_507,N_167,N_53);
or U508 (N_508,N_113,N_349);
nor U509 (N_509,N_317,N_230);
nand U510 (N_510,N_201,N_451);
nor U511 (N_511,N_278,N_128);
or U512 (N_512,N_7,N_20);
nor U513 (N_513,N_430,N_452);
xnor U514 (N_514,N_231,N_390);
xnor U515 (N_515,N_368,N_449);
nand U516 (N_516,N_237,N_431);
nor U517 (N_517,N_57,N_394);
xnor U518 (N_518,N_405,N_312);
nor U519 (N_519,N_208,N_438);
and U520 (N_520,N_325,N_76);
and U521 (N_521,N_8,N_27);
and U522 (N_522,N_106,N_183);
and U523 (N_523,N_226,N_144);
nand U524 (N_524,N_26,N_332);
or U525 (N_525,N_467,N_135);
nor U526 (N_526,N_143,N_112);
xor U527 (N_527,N_435,N_49);
nand U528 (N_528,N_108,N_425);
xor U529 (N_529,N_371,N_424);
nand U530 (N_530,N_139,N_292);
nand U531 (N_531,N_197,N_468);
nor U532 (N_532,N_473,N_364);
and U533 (N_533,N_427,N_491);
nor U534 (N_534,N_119,N_179);
xnor U535 (N_535,N_454,N_33);
xnor U536 (N_536,N_458,N_482);
nand U537 (N_537,N_63,N_34);
nor U538 (N_538,N_416,N_360);
nor U539 (N_539,N_132,N_382);
and U540 (N_540,N_293,N_289);
xnor U541 (N_541,N_62,N_156);
nor U542 (N_542,N_363,N_61);
xnor U543 (N_543,N_304,N_28);
nor U544 (N_544,N_362,N_302);
nor U545 (N_545,N_433,N_29);
or U546 (N_546,N_429,N_374);
nand U547 (N_547,N_399,N_376);
and U548 (N_548,N_264,N_184);
nor U549 (N_549,N_267,N_19);
or U550 (N_550,N_72,N_242);
nor U551 (N_551,N_367,N_0);
nand U552 (N_552,N_164,N_155);
nand U553 (N_553,N_379,N_271);
nor U554 (N_554,N_48,N_206);
nor U555 (N_555,N_496,N_97);
or U556 (N_556,N_265,N_36);
nor U557 (N_557,N_121,N_393);
and U558 (N_558,N_186,N_225);
nor U559 (N_559,N_444,N_150);
or U560 (N_560,N_263,N_219);
and U561 (N_561,N_494,N_77);
xnor U562 (N_562,N_377,N_455);
or U563 (N_563,N_181,N_120);
nand U564 (N_564,N_295,N_35);
or U565 (N_565,N_497,N_16);
or U566 (N_566,N_440,N_100);
or U567 (N_567,N_46,N_196);
or U568 (N_568,N_98,N_207);
nand U569 (N_569,N_60,N_443);
xnor U570 (N_570,N_114,N_241);
and U571 (N_571,N_366,N_474);
xor U572 (N_572,N_352,N_32);
nor U573 (N_573,N_169,N_274);
or U574 (N_574,N_470,N_127);
nor U575 (N_575,N_273,N_204);
xor U576 (N_576,N_175,N_9);
and U577 (N_577,N_116,N_96);
and U578 (N_578,N_495,N_462);
nor U579 (N_579,N_174,N_224);
or U580 (N_580,N_222,N_492);
or U581 (N_581,N_414,N_213);
or U582 (N_582,N_401,N_463);
or U583 (N_583,N_10,N_154);
nand U584 (N_584,N_249,N_244);
nand U585 (N_585,N_437,N_280);
nor U586 (N_586,N_99,N_199);
nor U587 (N_587,N_30,N_66);
and U588 (N_588,N_67,N_422);
and U589 (N_589,N_456,N_191);
or U590 (N_590,N_110,N_303);
nor U591 (N_591,N_369,N_408);
and U592 (N_592,N_333,N_160);
and U593 (N_593,N_447,N_464);
nand U594 (N_594,N_402,N_283);
or U595 (N_595,N_126,N_45);
nor U596 (N_596,N_43,N_445);
or U597 (N_597,N_300,N_409);
nor U598 (N_598,N_499,N_287);
xnor U599 (N_599,N_162,N_227);
and U600 (N_600,N_381,N_288);
or U601 (N_601,N_205,N_94);
or U602 (N_602,N_466,N_326);
nor U603 (N_603,N_338,N_58);
nor U604 (N_604,N_17,N_220);
or U605 (N_605,N_80,N_89);
and U606 (N_606,N_484,N_346);
and U607 (N_607,N_39,N_163);
nand U608 (N_608,N_248,N_56);
nand U609 (N_609,N_55,N_442);
and U610 (N_610,N_477,N_211);
and U611 (N_611,N_365,N_165);
and U612 (N_612,N_309,N_375);
nor U613 (N_613,N_420,N_12);
or U614 (N_614,N_90,N_488);
and U615 (N_615,N_232,N_103);
and U616 (N_616,N_318,N_487);
or U617 (N_617,N_315,N_261);
and U618 (N_618,N_342,N_256);
nand U619 (N_619,N_134,N_307);
nand U620 (N_620,N_417,N_239);
or U621 (N_621,N_290,N_324);
xor U622 (N_622,N_200,N_257);
and U623 (N_623,N_101,N_221);
nor U624 (N_624,N_299,N_141);
nand U625 (N_625,N_328,N_182);
nand U626 (N_626,N_339,N_275);
and U627 (N_627,N_353,N_210);
nor U628 (N_628,N_107,N_124);
and U629 (N_629,N_44,N_2);
nand U630 (N_630,N_460,N_347);
nor U631 (N_631,N_493,N_250);
or U632 (N_632,N_387,N_6);
nor U633 (N_633,N_459,N_461);
nand U634 (N_634,N_457,N_262);
or U635 (N_635,N_193,N_345);
or U636 (N_636,N_386,N_198);
xor U637 (N_637,N_469,N_380);
and U638 (N_638,N_260,N_296);
or U639 (N_639,N_188,N_178);
nand U640 (N_640,N_212,N_410);
xnor U641 (N_641,N_321,N_281);
nor U642 (N_642,N_272,N_319);
or U643 (N_643,N_301,N_70);
and U644 (N_644,N_68,N_370);
nand U645 (N_645,N_18,N_322);
nand U646 (N_646,N_395,N_356);
xor U647 (N_647,N_490,N_88);
or U648 (N_648,N_138,N_357);
and U649 (N_649,N_413,N_412);
nor U650 (N_650,N_330,N_146);
and U651 (N_651,N_258,N_323);
or U652 (N_652,N_453,N_209);
nor U653 (N_653,N_252,N_75);
or U654 (N_654,N_329,N_373);
and U655 (N_655,N_93,N_117);
xnor U656 (N_656,N_172,N_343);
or U657 (N_657,N_157,N_64);
and U658 (N_658,N_400,N_40);
nor U659 (N_659,N_1,N_109);
nor U660 (N_660,N_245,N_51);
and U661 (N_661,N_270,N_78);
and U662 (N_662,N_125,N_192);
or U663 (N_663,N_254,N_170);
nand U664 (N_664,N_446,N_483);
xnor U665 (N_665,N_269,N_355);
and U666 (N_666,N_471,N_359);
and U667 (N_667,N_4,N_91);
nor U668 (N_668,N_348,N_149);
nor U669 (N_669,N_69,N_202);
xnor U670 (N_670,N_71,N_398);
nor U671 (N_671,N_485,N_74);
and U672 (N_672,N_147,N_441);
or U673 (N_673,N_354,N_277);
nor U674 (N_674,N_276,N_223);
and U675 (N_675,N_418,N_87);
nor U676 (N_676,N_185,N_187);
nand U677 (N_677,N_31,N_358);
or U678 (N_678,N_336,N_426);
or U679 (N_679,N_50,N_498);
xnor U680 (N_680,N_285,N_25);
and U681 (N_681,N_153,N_234);
nor U682 (N_682,N_140,N_22);
and U683 (N_683,N_23,N_421);
nand U684 (N_684,N_298,N_279);
or U685 (N_685,N_41,N_84);
or U686 (N_686,N_308,N_392);
and U687 (N_687,N_314,N_238);
nand U688 (N_688,N_284,N_331);
or U689 (N_689,N_351,N_450);
nor U690 (N_690,N_52,N_14);
and U691 (N_691,N_137,N_478);
xor U692 (N_692,N_176,N_428);
or U693 (N_693,N_361,N_85);
nor U694 (N_694,N_148,N_215);
nor U695 (N_695,N_228,N_122);
nor U696 (N_696,N_73,N_102);
and U697 (N_697,N_251,N_216);
and U698 (N_698,N_475,N_105);
nor U699 (N_699,N_189,N_439);
or U700 (N_700,N_436,N_235);
xor U701 (N_701,N_217,N_166);
and U702 (N_702,N_297,N_286);
and U703 (N_703,N_344,N_253);
or U704 (N_704,N_233,N_95);
nor U705 (N_705,N_486,N_65);
and U706 (N_706,N_79,N_152);
nor U707 (N_707,N_465,N_266);
nor U708 (N_708,N_268,N_24);
and U709 (N_709,N_218,N_229);
or U710 (N_710,N_173,N_479);
nor U711 (N_711,N_161,N_131);
or U712 (N_712,N_489,N_294);
or U713 (N_713,N_236,N_142);
and U714 (N_714,N_5,N_282);
or U715 (N_715,N_203,N_334);
and U716 (N_716,N_391,N_115);
or U717 (N_717,N_190,N_397);
nor U718 (N_718,N_327,N_396);
nor U719 (N_719,N_385,N_151);
nor U720 (N_720,N_123,N_480);
and U721 (N_721,N_337,N_177);
nand U722 (N_722,N_419,N_259);
xor U723 (N_723,N_404,N_37);
nand U724 (N_724,N_86,N_384);
nor U725 (N_725,N_3,N_407);
nor U726 (N_726,N_341,N_195);
or U727 (N_727,N_472,N_434);
nand U728 (N_728,N_180,N_158);
nor U729 (N_729,N_378,N_240);
nand U730 (N_730,N_15,N_306);
and U731 (N_731,N_432,N_423);
or U732 (N_732,N_316,N_130);
and U733 (N_733,N_372,N_92);
or U734 (N_734,N_383,N_168);
nor U735 (N_735,N_403,N_111);
nand U736 (N_736,N_38,N_159);
nor U737 (N_737,N_104,N_415);
nor U738 (N_738,N_389,N_171);
and U739 (N_739,N_255,N_247);
and U740 (N_740,N_42,N_411);
or U741 (N_741,N_406,N_82);
or U742 (N_742,N_388,N_59);
and U743 (N_743,N_448,N_133);
xnor U744 (N_744,N_83,N_214);
nand U745 (N_745,N_243,N_310);
or U746 (N_746,N_313,N_320);
or U747 (N_747,N_291,N_47);
or U748 (N_748,N_335,N_340);
and U749 (N_749,N_476,N_481);
nor U750 (N_750,N_253,N_210);
and U751 (N_751,N_327,N_74);
and U752 (N_752,N_239,N_66);
and U753 (N_753,N_364,N_48);
nor U754 (N_754,N_331,N_199);
or U755 (N_755,N_285,N_31);
nor U756 (N_756,N_268,N_333);
nand U757 (N_757,N_263,N_296);
nand U758 (N_758,N_460,N_326);
nand U759 (N_759,N_301,N_336);
or U760 (N_760,N_188,N_95);
xnor U761 (N_761,N_9,N_286);
or U762 (N_762,N_413,N_36);
nor U763 (N_763,N_348,N_261);
xnor U764 (N_764,N_211,N_471);
and U765 (N_765,N_307,N_184);
nand U766 (N_766,N_461,N_494);
and U767 (N_767,N_304,N_185);
or U768 (N_768,N_389,N_109);
xor U769 (N_769,N_22,N_220);
nand U770 (N_770,N_70,N_186);
nand U771 (N_771,N_58,N_373);
xor U772 (N_772,N_145,N_383);
or U773 (N_773,N_143,N_199);
nor U774 (N_774,N_153,N_135);
nand U775 (N_775,N_270,N_126);
nand U776 (N_776,N_72,N_12);
nor U777 (N_777,N_197,N_426);
and U778 (N_778,N_379,N_328);
and U779 (N_779,N_279,N_239);
or U780 (N_780,N_308,N_460);
nand U781 (N_781,N_65,N_214);
and U782 (N_782,N_39,N_114);
and U783 (N_783,N_415,N_430);
and U784 (N_784,N_147,N_244);
and U785 (N_785,N_243,N_406);
nand U786 (N_786,N_406,N_449);
or U787 (N_787,N_305,N_460);
or U788 (N_788,N_310,N_73);
xor U789 (N_789,N_236,N_343);
nor U790 (N_790,N_355,N_284);
and U791 (N_791,N_278,N_333);
and U792 (N_792,N_210,N_169);
nand U793 (N_793,N_271,N_227);
or U794 (N_794,N_463,N_123);
and U795 (N_795,N_211,N_438);
or U796 (N_796,N_469,N_219);
nor U797 (N_797,N_217,N_207);
nor U798 (N_798,N_241,N_210);
and U799 (N_799,N_122,N_404);
nor U800 (N_800,N_283,N_177);
and U801 (N_801,N_16,N_289);
and U802 (N_802,N_366,N_82);
or U803 (N_803,N_216,N_114);
nand U804 (N_804,N_68,N_362);
or U805 (N_805,N_316,N_126);
and U806 (N_806,N_420,N_448);
xor U807 (N_807,N_16,N_189);
or U808 (N_808,N_435,N_175);
or U809 (N_809,N_364,N_209);
nand U810 (N_810,N_481,N_175);
xor U811 (N_811,N_44,N_220);
nand U812 (N_812,N_2,N_403);
or U813 (N_813,N_472,N_180);
and U814 (N_814,N_383,N_475);
or U815 (N_815,N_411,N_18);
and U816 (N_816,N_172,N_80);
nand U817 (N_817,N_348,N_269);
and U818 (N_818,N_327,N_325);
or U819 (N_819,N_282,N_310);
nand U820 (N_820,N_35,N_296);
xnor U821 (N_821,N_83,N_169);
nor U822 (N_822,N_315,N_437);
nand U823 (N_823,N_475,N_367);
nand U824 (N_824,N_321,N_141);
and U825 (N_825,N_392,N_429);
nand U826 (N_826,N_215,N_483);
or U827 (N_827,N_304,N_84);
nand U828 (N_828,N_135,N_186);
and U829 (N_829,N_89,N_56);
nand U830 (N_830,N_143,N_436);
xnor U831 (N_831,N_135,N_447);
or U832 (N_832,N_394,N_334);
or U833 (N_833,N_320,N_120);
nor U834 (N_834,N_284,N_247);
nand U835 (N_835,N_133,N_279);
nor U836 (N_836,N_325,N_98);
nand U837 (N_837,N_186,N_419);
nor U838 (N_838,N_359,N_27);
and U839 (N_839,N_60,N_34);
nand U840 (N_840,N_328,N_50);
nor U841 (N_841,N_235,N_28);
xor U842 (N_842,N_214,N_197);
and U843 (N_843,N_408,N_212);
xnor U844 (N_844,N_9,N_323);
nor U845 (N_845,N_443,N_63);
or U846 (N_846,N_82,N_39);
and U847 (N_847,N_40,N_425);
and U848 (N_848,N_144,N_56);
nand U849 (N_849,N_76,N_215);
nor U850 (N_850,N_23,N_395);
and U851 (N_851,N_392,N_52);
and U852 (N_852,N_240,N_434);
nor U853 (N_853,N_197,N_219);
nand U854 (N_854,N_82,N_360);
nor U855 (N_855,N_33,N_194);
nand U856 (N_856,N_253,N_48);
xor U857 (N_857,N_58,N_119);
and U858 (N_858,N_438,N_165);
or U859 (N_859,N_371,N_311);
and U860 (N_860,N_3,N_389);
and U861 (N_861,N_389,N_43);
and U862 (N_862,N_121,N_250);
xor U863 (N_863,N_478,N_327);
and U864 (N_864,N_425,N_232);
or U865 (N_865,N_428,N_441);
or U866 (N_866,N_294,N_337);
nor U867 (N_867,N_423,N_87);
nand U868 (N_868,N_320,N_81);
xnor U869 (N_869,N_210,N_20);
nor U870 (N_870,N_99,N_124);
and U871 (N_871,N_441,N_41);
nand U872 (N_872,N_344,N_14);
xor U873 (N_873,N_75,N_78);
and U874 (N_874,N_88,N_269);
and U875 (N_875,N_21,N_278);
nor U876 (N_876,N_100,N_217);
xor U877 (N_877,N_217,N_444);
xor U878 (N_878,N_83,N_420);
and U879 (N_879,N_470,N_294);
nor U880 (N_880,N_68,N_387);
or U881 (N_881,N_349,N_125);
nand U882 (N_882,N_373,N_285);
or U883 (N_883,N_402,N_386);
or U884 (N_884,N_433,N_214);
nand U885 (N_885,N_189,N_224);
nor U886 (N_886,N_402,N_186);
and U887 (N_887,N_343,N_156);
xor U888 (N_888,N_132,N_399);
nor U889 (N_889,N_428,N_23);
and U890 (N_890,N_355,N_452);
or U891 (N_891,N_20,N_143);
and U892 (N_892,N_332,N_360);
nor U893 (N_893,N_172,N_489);
or U894 (N_894,N_324,N_140);
nand U895 (N_895,N_92,N_12);
nand U896 (N_896,N_415,N_270);
or U897 (N_897,N_391,N_394);
nor U898 (N_898,N_387,N_499);
nor U899 (N_899,N_62,N_199);
xor U900 (N_900,N_416,N_181);
nand U901 (N_901,N_52,N_396);
nor U902 (N_902,N_22,N_217);
nand U903 (N_903,N_386,N_442);
and U904 (N_904,N_392,N_163);
nor U905 (N_905,N_1,N_493);
nor U906 (N_906,N_477,N_480);
nor U907 (N_907,N_470,N_25);
xnor U908 (N_908,N_9,N_70);
nor U909 (N_909,N_197,N_211);
and U910 (N_910,N_2,N_381);
nor U911 (N_911,N_177,N_40);
nor U912 (N_912,N_271,N_300);
and U913 (N_913,N_460,N_424);
nand U914 (N_914,N_333,N_64);
xor U915 (N_915,N_121,N_101);
nor U916 (N_916,N_349,N_26);
and U917 (N_917,N_41,N_326);
or U918 (N_918,N_450,N_354);
xnor U919 (N_919,N_295,N_101);
xnor U920 (N_920,N_263,N_25);
or U921 (N_921,N_474,N_228);
nor U922 (N_922,N_355,N_343);
nor U923 (N_923,N_315,N_173);
xor U924 (N_924,N_21,N_98);
nor U925 (N_925,N_444,N_157);
or U926 (N_926,N_442,N_74);
and U927 (N_927,N_41,N_164);
nor U928 (N_928,N_32,N_280);
or U929 (N_929,N_187,N_11);
xor U930 (N_930,N_200,N_430);
nor U931 (N_931,N_35,N_313);
nor U932 (N_932,N_378,N_451);
and U933 (N_933,N_399,N_145);
or U934 (N_934,N_301,N_451);
and U935 (N_935,N_217,N_383);
nand U936 (N_936,N_367,N_350);
or U937 (N_937,N_369,N_231);
xor U938 (N_938,N_158,N_350);
nand U939 (N_939,N_176,N_326);
and U940 (N_940,N_133,N_56);
nand U941 (N_941,N_13,N_344);
or U942 (N_942,N_133,N_467);
nand U943 (N_943,N_18,N_29);
nand U944 (N_944,N_150,N_164);
and U945 (N_945,N_314,N_289);
or U946 (N_946,N_266,N_172);
or U947 (N_947,N_424,N_122);
nand U948 (N_948,N_488,N_25);
or U949 (N_949,N_1,N_119);
nand U950 (N_950,N_148,N_223);
nand U951 (N_951,N_38,N_85);
or U952 (N_952,N_373,N_19);
or U953 (N_953,N_80,N_17);
and U954 (N_954,N_285,N_170);
and U955 (N_955,N_238,N_417);
or U956 (N_956,N_98,N_315);
nand U957 (N_957,N_370,N_496);
nand U958 (N_958,N_331,N_201);
and U959 (N_959,N_483,N_36);
and U960 (N_960,N_134,N_258);
nor U961 (N_961,N_320,N_94);
and U962 (N_962,N_64,N_16);
or U963 (N_963,N_120,N_35);
nand U964 (N_964,N_308,N_391);
xor U965 (N_965,N_173,N_374);
nand U966 (N_966,N_76,N_488);
nand U967 (N_967,N_458,N_25);
nand U968 (N_968,N_325,N_491);
xnor U969 (N_969,N_140,N_11);
and U970 (N_970,N_248,N_285);
and U971 (N_971,N_269,N_178);
nor U972 (N_972,N_299,N_275);
nand U973 (N_973,N_362,N_107);
and U974 (N_974,N_425,N_160);
or U975 (N_975,N_205,N_106);
and U976 (N_976,N_232,N_188);
nand U977 (N_977,N_62,N_439);
nand U978 (N_978,N_411,N_22);
nand U979 (N_979,N_79,N_204);
nor U980 (N_980,N_32,N_1);
nand U981 (N_981,N_202,N_31);
nor U982 (N_982,N_270,N_260);
and U983 (N_983,N_222,N_351);
and U984 (N_984,N_482,N_239);
or U985 (N_985,N_113,N_398);
nand U986 (N_986,N_216,N_125);
or U987 (N_987,N_9,N_48);
nand U988 (N_988,N_234,N_302);
or U989 (N_989,N_411,N_249);
nand U990 (N_990,N_386,N_155);
and U991 (N_991,N_171,N_369);
or U992 (N_992,N_259,N_199);
nand U993 (N_993,N_11,N_194);
and U994 (N_994,N_286,N_361);
or U995 (N_995,N_251,N_209);
nand U996 (N_996,N_64,N_464);
nor U997 (N_997,N_278,N_258);
or U998 (N_998,N_466,N_229);
and U999 (N_999,N_384,N_39);
or U1000 (N_1000,N_833,N_964);
xnor U1001 (N_1001,N_751,N_911);
or U1002 (N_1002,N_693,N_558);
xor U1003 (N_1003,N_812,N_729);
xnor U1004 (N_1004,N_761,N_805);
or U1005 (N_1005,N_528,N_999);
or U1006 (N_1006,N_508,N_672);
and U1007 (N_1007,N_828,N_983);
nor U1008 (N_1008,N_872,N_897);
nor U1009 (N_1009,N_647,N_668);
nor U1010 (N_1010,N_832,N_803);
nand U1011 (N_1011,N_825,N_847);
nor U1012 (N_1012,N_859,N_741);
nor U1013 (N_1013,N_598,N_992);
nor U1014 (N_1014,N_656,N_666);
nor U1015 (N_1015,N_703,N_652);
xnor U1016 (N_1016,N_762,N_695);
nand U1017 (N_1017,N_869,N_745);
and U1018 (N_1018,N_605,N_600);
or U1019 (N_1019,N_694,N_994);
nand U1020 (N_1020,N_644,N_720);
nand U1021 (N_1021,N_798,N_754);
nand U1022 (N_1022,N_519,N_628);
or U1023 (N_1023,N_548,N_629);
or U1024 (N_1024,N_535,N_568);
nor U1025 (N_1025,N_549,N_737);
or U1026 (N_1026,N_986,N_640);
and U1027 (N_1027,N_526,N_830);
nor U1028 (N_1028,N_939,N_697);
xor U1029 (N_1029,N_739,N_961);
nand U1030 (N_1030,N_619,N_804);
nor U1031 (N_1031,N_837,N_881);
nor U1032 (N_1032,N_532,N_716);
and U1033 (N_1033,N_602,N_854);
nor U1034 (N_1034,N_722,N_910);
or U1035 (N_1035,N_544,N_546);
xnor U1036 (N_1036,N_844,N_721);
nor U1037 (N_1037,N_815,N_930);
nor U1038 (N_1038,N_587,N_740);
and U1039 (N_1039,N_642,N_915);
nor U1040 (N_1040,N_505,N_514);
nor U1041 (N_1041,N_507,N_823);
nand U1042 (N_1042,N_891,N_503);
nor U1043 (N_1043,N_521,N_743);
nand U1044 (N_1044,N_905,N_809);
nor U1045 (N_1045,N_578,N_843);
and U1046 (N_1046,N_931,N_554);
nor U1047 (N_1047,N_635,N_683);
nand U1048 (N_1048,N_923,N_597);
or U1049 (N_1049,N_820,N_615);
nor U1050 (N_1050,N_664,N_900);
nor U1051 (N_1051,N_632,N_922);
nor U1052 (N_1052,N_902,N_772);
and U1053 (N_1053,N_614,N_572);
nor U1054 (N_1054,N_726,N_529);
or U1055 (N_1055,N_790,N_565);
or U1056 (N_1056,N_858,N_935);
nand U1057 (N_1057,N_955,N_840);
nor U1058 (N_1058,N_715,N_564);
nand U1059 (N_1059,N_993,N_914);
and U1060 (N_1060,N_696,N_878);
or U1061 (N_1061,N_756,N_516);
nor U1062 (N_1062,N_945,N_776);
nand U1063 (N_1063,N_953,N_541);
or U1064 (N_1064,N_971,N_995);
and U1065 (N_1065,N_792,N_620);
and U1066 (N_1066,N_661,N_609);
and U1067 (N_1067,N_785,N_967);
nand U1068 (N_1068,N_796,N_731);
nor U1069 (N_1069,N_511,N_969);
nand U1070 (N_1070,N_977,N_612);
nand U1071 (N_1071,N_706,N_944);
and U1072 (N_1072,N_637,N_690);
nand U1073 (N_1073,N_960,N_876);
and U1074 (N_1074,N_545,N_929);
or U1075 (N_1075,N_894,N_829);
and U1076 (N_1076,N_870,N_566);
nor U1077 (N_1077,N_807,N_898);
or U1078 (N_1078,N_691,N_571);
nor U1079 (N_1079,N_752,N_538);
or U1080 (N_1080,N_657,N_822);
nand U1081 (N_1081,N_727,N_592);
nor U1082 (N_1082,N_608,N_603);
and U1083 (N_1083,N_787,N_821);
and U1084 (N_1084,N_692,N_595);
or U1085 (N_1085,N_708,N_579);
and U1086 (N_1086,N_799,N_968);
or U1087 (N_1087,N_801,N_938);
xnor U1088 (N_1088,N_730,N_641);
nor U1089 (N_1089,N_895,N_636);
and U1090 (N_1090,N_951,N_996);
nand U1091 (N_1091,N_634,N_979);
and U1092 (N_1092,N_921,N_622);
nor U1093 (N_1093,N_523,N_723);
or U1094 (N_1094,N_845,N_838);
nor U1095 (N_1095,N_537,N_633);
and U1096 (N_1096,N_728,N_972);
nand U1097 (N_1097,N_610,N_757);
xnor U1098 (N_1098,N_784,N_937);
nand U1099 (N_1099,N_989,N_501);
nand U1100 (N_1100,N_700,N_686);
nand U1101 (N_1101,N_886,N_848);
nand U1102 (N_1102,N_601,N_574);
nand U1103 (N_1103,N_880,N_827);
and U1104 (N_1104,N_839,N_724);
and U1105 (N_1105,N_525,N_788);
and U1106 (N_1106,N_940,N_981);
or U1107 (N_1107,N_725,N_570);
and U1108 (N_1108,N_714,N_534);
or U1109 (N_1109,N_689,N_750);
and U1110 (N_1110,N_717,N_956);
nor U1111 (N_1111,N_674,N_860);
xor U1112 (N_1112,N_709,N_638);
xor U1113 (N_1113,N_861,N_543);
nand U1114 (N_1114,N_681,N_651);
nand U1115 (N_1115,N_950,N_959);
nor U1116 (N_1116,N_780,N_875);
nand U1117 (N_1117,N_718,N_679);
nor U1118 (N_1118,N_824,N_753);
or U1119 (N_1119,N_888,N_583);
nand U1120 (N_1120,N_517,N_766);
nor U1121 (N_1121,N_997,N_621);
nor U1122 (N_1122,N_903,N_687);
and U1123 (N_1123,N_678,N_575);
nor U1124 (N_1124,N_626,N_966);
nand U1125 (N_1125,N_536,N_819);
nor U1126 (N_1126,N_863,N_871);
nor U1127 (N_1127,N_589,N_639);
nand U1128 (N_1128,N_506,N_925);
nand U1129 (N_1129,N_795,N_794);
and U1130 (N_1130,N_735,N_867);
nor U1131 (N_1131,N_596,N_588);
and U1132 (N_1132,N_857,N_849);
and U1133 (N_1133,N_947,N_648);
or U1134 (N_1134,N_982,N_623);
nor U1135 (N_1135,N_707,N_527);
xor U1136 (N_1136,N_758,N_625);
and U1137 (N_1137,N_530,N_711);
and U1138 (N_1138,N_818,N_613);
or U1139 (N_1139,N_698,N_942);
or U1140 (N_1140,N_941,N_893);
and U1141 (N_1141,N_577,N_561);
and U1142 (N_1142,N_631,N_531);
or U1143 (N_1143,N_771,N_786);
xor U1144 (N_1144,N_800,N_851);
and U1145 (N_1145,N_599,N_813);
or U1146 (N_1146,N_581,N_755);
xnor U1147 (N_1147,N_684,N_590);
nand U1148 (N_1148,N_909,N_917);
or U1149 (N_1149,N_591,N_585);
nor U1150 (N_1150,N_913,N_932);
and U1151 (N_1151,N_701,N_747);
nand U1152 (N_1152,N_665,N_865);
and U1153 (N_1153,N_943,N_883);
xor U1154 (N_1154,N_510,N_949);
and U1155 (N_1155,N_770,N_593);
nor U1156 (N_1156,N_797,N_767);
nor U1157 (N_1157,N_744,N_948);
nand U1158 (N_1158,N_906,N_984);
nor U1159 (N_1159,N_892,N_582);
nor U1160 (N_1160,N_879,N_524);
or U1161 (N_1161,N_663,N_733);
nand U1162 (N_1162,N_630,N_952);
nor U1163 (N_1163,N_826,N_896);
nand U1164 (N_1164,N_963,N_560);
and U1165 (N_1165,N_936,N_974);
or U1166 (N_1166,N_580,N_901);
nor U1167 (N_1167,N_653,N_811);
or U1168 (N_1168,N_862,N_885);
nand U1169 (N_1169,N_985,N_978);
nand U1170 (N_1170,N_904,N_688);
nand U1171 (N_1171,N_810,N_778);
and U1172 (N_1172,N_748,N_781);
nor U1173 (N_1173,N_779,N_873);
and U1174 (N_1174,N_675,N_556);
nand U1175 (N_1175,N_899,N_624);
or U1176 (N_1176,N_889,N_533);
nor U1177 (N_1177,N_775,N_611);
or U1178 (N_1178,N_562,N_842);
nand U1179 (N_1179,N_831,N_970);
xnor U1180 (N_1180,N_954,N_669);
and U1181 (N_1181,N_557,N_606);
or U1182 (N_1182,N_908,N_710);
nor U1183 (N_1183,N_789,N_515);
or U1184 (N_1184,N_573,N_987);
or U1185 (N_1185,N_607,N_890);
nor U1186 (N_1186,N_887,N_783);
nor U1187 (N_1187,N_504,N_973);
nand U1188 (N_1188,N_976,N_736);
nor U1189 (N_1189,N_868,N_927);
xnor U1190 (N_1190,N_685,N_918);
and U1191 (N_1191,N_509,N_671);
nor U1192 (N_1192,N_836,N_576);
and U1193 (N_1193,N_522,N_884);
xor U1194 (N_1194,N_975,N_616);
or U1195 (N_1195,N_667,N_907);
and U1196 (N_1196,N_777,N_513);
nand U1197 (N_1197,N_808,N_802);
nor U1198 (N_1198,N_542,N_817);
or U1199 (N_1199,N_850,N_742);
and U1200 (N_1200,N_699,N_957);
nand U1201 (N_1201,N_806,N_933);
nor U1202 (N_1202,N_760,N_550);
xnor U1203 (N_1203,N_877,N_732);
and U1204 (N_1204,N_655,N_856);
nor U1205 (N_1205,N_928,N_500);
nor U1206 (N_1206,N_540,N_846);
and U1207 (N_1207,N_924,N_852);
nand U1208 (N_1208,N_712,N_926);
and U1209 (N_1209,N_874,N_835);
and U1210 (N_1210,N_604,N_853);
or U1211 (N_1211,N_773,N_547);
nand U1212 (N_1212,N_518,N_763);
or U1213 (N_1213,N_654,N_991);
or U1214 (N_1214,N_965,N_676);
or U1215 (N_1215,N_841,N_774);
nor U1216 (N_1216,N_934,N_919);
and U1217 (N_1217,N_662,N_555);
or U1218 (N_1218,N_650,N_920);
and U1219 (N_1219,N_791,N_746);
and U1220 (N_1220,N_704,N_834);
nand U1221 (N_1221,N_946,N_670);
or U1222 (N_1222,N_512,N_677);
nor U1223 (N_1223,N_764,N_793);
nand U1224 (N_1224,N_866,N_990);
and U1225 (N_1225,N_586,N_962);
nand U1226 (N_1226,N_882,N_864);
and U1227 (N_1227,N_682,N_980);
and U1228 (N_1228,N_649,N_551);
nand U1229 (N_1229,N_594,N_584);
or U1230 (N_1230,N_645,N_643);
and U1231 (N_1231,N_816,N_618);
or U1232 (N_1232,N_738,N_659);
nand U1233 (N_1233,N_988,N_719);
nor U1234 (N_1234,N_559,N_660);
or U1235 (N_1235,N_855,N_627);
or U1236 (N_1236,N_673,N_680);
or U1237 (N_1237,N_563,N_814);
nand U1238 (N_1238,N_912,N_553);
and U1239 (N_1239,N_520,N_759);
nand U1240 (N_1240,N_782,N_552);
or U1241 (N_1241,N_658,N_765);
and U1242 (N_1242,N_646,N_768);
and U1243 (N_1243,N_569,N_705);
and U1244 (N_1244,N_916,N_567);
or U1245 (N_1245,N_998,N_539);
and U1246 (N_1246,N_502,N_749);
or U1247 (N_1247,N_617,N_702);
nand U1248 (N_1248,N_734,N_713);
and U1249 (N_1249,N_769,N_958);
and U1250 (N_1250,N_651,N_909);
nand U1251 (N_1251,N_802,N_748);
nor U1252 (N_1252,N_657,N_879);
nand U1253 (N_1253,N_567,N_686);
and U1254 (N_1254,N_896,N_602);
and U1255 (N_1255,N_825,N_738);
and U1256 (N_1256,N_603,N_652);
nor U1257 (N_1257,N_536,N_929);
nor U1258 (N_1258,N_629,N_994);
nand U1259 (N_1259,N_844,N_872);
and U1260 (N_1260,N_846,N_958);
or U1261 (N_1261,N_863,N_677);
xor U1262 (N_1262,N_909,N_826);
and U1263 (N_1263,N_752,N_601);
and U1264 (N_1264,N_590,N_880);
nand U1265 (N_1265,N_682,N_714);
and U1266 (N_1266,N_598,N_887);
and U1267 (N_1267,N_689,N_830);
xnor U1268 (N_1268,N_582,N_526);
or U1269 (N_1269,N_899,N_626);
and U1270 (N_1270,N_929,N_919);
nand U1271 (N_1271,N_675,N_964);
nand U1272 (N_1272,N_534,N_679);
nor U1273 (N_1273,N_987,N_645);
xnor U1274 (N_1274,N_986,N_739);
nor U1275 (N_1275,N_559,N_971);
xnor U1276 (N_1276,N_552,N_509);
or U1277 (N_1277,N_708,N_653);
and U1278 (N_1278,N_884,N_663);
nand U1279 (N_1279,N_566,N_625);
nand U1280 (N_1280,N_903,N_902);
and U1281 (N_1281,N_934,N_799);
nor U1282 (N_1282,N_762,N_738);
and U1283 (N_1283,N_986,N_661);
or U1284 (N_1284,N_975,N_946);
nor U1285 (N_1285,N_937,N_567);
and U1286 (N_1286,N_923,N_721);
xor U1287 (N_1287,N_736,N_839);
or U1288 (N_1288,N_559,N_508);
nand U1289 (N_1289,N_972,N_907);
nor U1290 (N_1290,N_522,N_945);
or U1291 (N_1291,N_520,N_884);
or U1292 (N_1292,N_542,N_561);
nor U1293 (N_1293,N_772,N_722);
or U1294 (N_1294,N_869,N_633);
nor U1295 (N_1295,N_674,N_878);
or U1296 (N_1296,N_828,N_553);
nor U1297 (N_1297,N_613,N_616);
and U1298 (N_1298,N_568,N_704);
nand U1299 (N_1299,N_847,N_679);
xnor U1300 (N_1300,N_531,N_953);
nor U1301 (N_1301,N_829,N_670);
and U1302 (N_1302,N_831,N_699);
nor U1303 (N_1303,N_571,N_595);
nor U1304 (N_1304,N_508,N_523);
or U1305 (N_1305,N_582,N_899);
nor U1306 (N_1306,N_988,N_554);
and U1307 (N_1307,N_761,N_669);
and U1308 (N_1308,N_916,N_881);
or U1309 (N_1309,N_792,N_574);
and U1310 (N_1310,N_874,N_644);
xor U1311 (N_1311,N_510,N_537);
nor U1312 (N_1312,N_905,N_524);
xor U1313 (N_1313,N_990,N_855);
and U1314 (N_1314,N_577,N_648);
nand U1315 (N_1315,N_923,N_866);
nor U1316 (N_1316,N_757,N_574);
and U1317 (N_1317,N_557,N_915);
xor U1318 (N_1318,N_529,N_843);
or U1319 (N_1319,N_811,N_595);
nand U1320 (N_1320,N_691,N_633);
or U1321 (N_1321,N_986,N_614);
nand U1322 (N_1322,N_829,N_671);
nor U1323 (N_1323,N_577,N_797);
or U1324 (N_1324,N_680,N_685);
nor U1325 (N_1325,N_922,N_507);
nand U1326 (N_1326,N_595,N_793);
xnor U1327 (N_1327,N_799,N_816);
nor U1328 (N_1328,N_733,N_721);
and U1329 (N_1329,N_935,N_818);
nand U1330 (N_1330,N_775,N_854);
or U1331 (N_1331,N_954,N_526);
or U1332 (N_1332,N_873,N_663);
and U1333 (N_1333,N_837,N_717);
or U1334 (N_1334,N_635,N_593);
or U1335 (N_1335,N_624,N_820);
nand U1336 (N_1336,N_521,N_826);
nor U1337 (N_1337,N_639,N_597);
and U1338 (N_1338,N_821,N_538);
and U1339 (N_1339,N_857,N_528);
nor U1340 (N_1340,N_986,N_655);
nand U1341 (N_1341,N_663,N_896);
and U1342 (N_1342,N_978,N_826);
nand U1343 (N_1343,N_830,N_549);
or U1344 (N_1344,N_505,N_789);
xnor U1345 (N_1345,N_776,N_979);
and U1346 (N_1346,N_579,N_603);
nand U1347 (N_1347,N_500,N_617);
nand U1348 (N_1348,N_781,N_514);
and U1349 (N_1349,N_615,N_562);
nand U1350 (N_1350,N_966,N_853);
nand U1351 (N_1351,N_977,N_937);
and U1352 (N_1352,N_593,N_993);
or U1353 (N_1353,N_794,N_503);
nand U1354 (N_1354,N_583,N_769);
nor U1355 (N_1355,N_774,N_778);
nand U1356 (N_1356,N_788,N_507);
xnor U1357 (N_1357,N_723,N_847);
and U1358 (N_1358,N_666,N_808);
or U1359 (N_1359,N_632,N_577);
nor U1360 (N_1360,N_603,N_961);
xor U1361 (N_1361,N_809,N_587);
nor U1362 (N_1362,N_846,N_891);
nand U1363 (N_1363,N_986,N_674);
nand U1364 (N_1364,N_536,N_526);
nor U1365 (N_1365,N_900,N_813);
and U1366 (N_1366,N_688,N_863);
and U1367 (N_1367,N_635,N_975);
nand U1368 (N_1368,N_991,N_912);
nand U1369 (N_1369,N_514,N_756);
and U1370 (N_1370,N_649,N_981);
nor U1371 (N_1371,N_751,N_935);
nor U1372 (N_1372,N_561,N_754);
or U1373 (N_1373,N_875,N_651);
nand U1374 (N_1374,N_940,N_870);
and U1375 (N_1375,N_792,N_922);
and U1376 (N_1376,N_886,N_881);
nor U1377 (N_1377,N_716,N_836);
and U1378 (N_1378,N_860,N_904);
and U1379 (N_1379,N_786,N_717);
xnor U1380 (N_1380,N_562,N_619);
nand U1381 (N_1381,N_814,N_977);
nor U1382 (N_1382,N_913,N_521);
or U1383 (N_1383,N_711,N_814);
and U1384 (N_1384,N_758,N_563);
and U1385 (N_1385,N_685,N_582);
and U1386 (N_1386,N_876,N_617);
nor U1387 (N_1387,N_817,N_841);
nor U1388 (N_1388,N_851,N_815);
and U1389 (N_1389,N_919,N_598);
or U1390 (N_1390,N_981,N_619);
and U1391 (N_1391,N_727,N_588);
and U1392 (N_1392,N_630,N_956);
or U1393 (N_1393,N_507,N_723);
and U1394 (N_1394,N_994,N_911);
nand U1395 (N_1395,N_821,N_686);
nor U1396 (N_1396,N_951,N_624);
nand U1397 (N_1397,N_903,N_811);
and U1398 (N_1398,N_881,N_742);
and U1399 (N_1399,N_692,N_857);
nand U1400 (N_1400,N_556,N_788);
nand U1401 (N_1401,N_559,N_792);
nand U1402 (N_1402,N_632,N_946);
nor U1403 (N_1403,N_866,N_780);
and U1404 (N_1404,N_522,N_739);
nand U1405 (N_1405,N_709,N_946);
or U1406 (N_1406,N_705,N_596);
or U1407 (N_1407,N_581,N_650);
nand U1408 (N_1408,N_509,N_787);
nand U1409 (N_1409,N_684,N_987);
xor U1410 (N_1410,N_820,N_501);
and U1411 (N_1411,N_766,N_803);
nor U1412 (N_1412,N_956,N_796);
nand U1413 (N_1413,N_740,N_742);
and U1414 (N_1414,N_539,N_644);
nand U1415 (N_1415,N_765,N_803);
nor U1416 (N_1416,N_616,N_598);
nor U1417 (N_1417,N_692,N_693);
nand U1418 (N_1418,N_918,N_911);
or U1419 (N_1419,N_694,N_632);
or U1420 (N_1420,N_940,N_919);
or U1421 (N_1421,N_853,N_907);
xor U1422 (N_1422,N_517,N_638);
nand U1423 (N_1423,N_934,N_680);
nand U1424 (N_1424,N_732,N_723);
and U1425 (N_1425,N_994,N_659);
or U1426 (N_1426,N_605,N_759);
nor U1427 (N_1427,N_681,N_973);
or U1428 (N_1428,N_763,N_680);
nand U1429 (N_1429,N_551,N_661);
xor U1430 (N_1430,N_729,N_886);
and U1431 (N_1431,N_635,N_562);
nor U1432 (N_1432,N_906,N_760);
nor U1433 (N_1433,N_858,N_857);
nor U1434 (N_1434,N_603,N_638);
nand U1435 (N_1435,N_789,N_698);
or U1436 (N_1436,N_614,N_778);
xor U1437 (N_1437,N_869,N_880);
or U1438 (N_1438,N_630,N_537);
nor U1439 (N_1439,N_556,N_787);
or U1440 (N_1440,N_911,N_739);
nor U1441 (N_1441,N_558,N_670);
and U1442 (N_1442,N_971,N_951);
nor U1443 (N_1443,N_835,N_830);
or U1444 (N_1444,N_804,N_920);
nand U1445 (N_1445,N_775,N_804);
nor U1446 (N_1446,N_531,N_576);
or U1447 (N_1447,N_504,N_668);
nand U1448 (N_1448,N_592,N_701);
xnor U1449 (N_1449,N_672,N_728);
or U1450 (N_1450,N_993,N_851);
and U1451 (N_1451,N_549,N_532);
and U1452 (N_1452,N_858,N_956);
xor U1453 (N_1453,N_863,N_948);
and U1454 (N_1454,N_810,N_987);
and U1455 (N_1455,N_780,N_759);
nor U1456 (N_1456,N_801,N_612);
nor U1457 (N_1457,N_635,N_830);
nand U1458 (N_1458,N_928,N_898);
or U1459 (N_1459,N_870,N_840);
and U1460 (N_1460,N_846,N_595);
nor U1461 (N_1461,N_853,N_825);
nor U1462 (N_1462,N_703,N_902);
or U1463 (N_1463,N_650,N_543);
or U1464 (N_1464,N_725,N_777);
and U1465 (N_1465,N_693,N_839);
nor U1466 (N_1466,N_767,N_788);
nand U1467 (N_1467,N_591,N_803);
nor U1468 (N_1468,N_561,N_924);
nand U1469 (N_1469,N_808,N_521);
nand U1470 (N_1470,N_585,N_996);
nor U1471 (N_1471,N_780,N_856);
or U1472 (N_1472,N_523,N_560);
nand U1473 (N_1473,N_921,N_668);
and U1474 (N_1474,N_903,N_805);
xor U1475 (N_1475,N_782,N_911);
and U1476 (N_1476,N_628,N_825);
or U1477 (N_1477,N_862,N_673);
nor U1478 (N_1478,N_620,N_986);
or U1479 (N_1479,N_814,N_922);
xnor U1480 (N_1480,N_815,N_671);
or U1481 (N_1481,N_726,N_573);
and U1482 (N_1482,N_893,N_534);
nor U1483 (N_1483,N_919,N_699);
nand U1484 (N_1484,N_535,N_517);
and U1485 (N_1485,N_826,N_533);
nor U1486 (N_1486,N_701,N_575);
or U1487 (N_1487,N_701,N_550);
xnor U1488 (N_1488,N_949,N_962);
nand U1489 (N_1489,N_829,N_822);
nor U1490 (N_1490,N_593,N_821);
nor U1491 (N_1491,N_765,N_584);
nor U1492 (N_1492,N_973,N_869);
nor U1493 (N_1493,N_709,N_854);
xor U1494 (N_1494,N_861,N_538);
xor U1495 (N_1495,N_711,N_939);
nand U1496 (N_1496,N_771,N_655);
xor U1497 (N_1497,N_865,N_896);
xor U1498 (N_1498,N_940,N_972);
and U1499 (N_1499,N_775,N_666);
xnor U1500 (N_1500,N_1461,N_1184);
xnor U1501 (N_1501,N_1013,N_1023);
or U1502 (N_1502,N_1346,N_1279);
nand U1503 (N_1503,N_1098,N_1322);
nor U1504 (N_1504,N_1062,N_1429);
nor U1505 (N_1505,N_1196,N_1448);
nand U1506 (N_1506,N_1263,N_1056);
or U1507 (N_1507,N_1016,N_1412);
xor U1508 (N_1508,N_1038,N_1345);
nand U1509 (N_1509,N_1291,N_1180);
and U1510 (N_1510,N_1402,N_1252);
xnor U1511 (N_1511,N_1024,N_1383);
nand U1512 (N_1512,N_1048,N_1108);
and U1513 (N_1513,N_1266,N_1189);
or U1514 (N_1514,N_1361,N_1101);
nand U1515 (N_1515,N_1002,N_1115);
nand U1516 (N_1516,N_1157,N_1372);
or U1517 (N_1517,N_1264,N_1432);
and U1518 (N_1518,N_1274,N_1401);
or U1519 (N_1519,N_1281,N_1214);
or U1520 (N_1520,N_1090,N_1276);
xor U1521 (N_1521,N_1210,N_1234);
nand U1522 (N_1522,N_1193,N_1363);
and U1523 (N_1523,N_1467,N_1083);
nand U1524 (N_1524,N_1220,N_1445);
or U1525 (N_1525,N_1319,N_1035);
nand U1526 (N_1526,N_1265,N_1208);
nand U1527 (N_1527,N_1040,N_1139);
xnor U1528 (N_1528,N_1007,N_1162);
nor U1529 (N_1529,N_1267,N_1046);
nor U1530 (N_1530,N_1073,N_1029);
or U1531 (N_1531,N_1063,N_1354);
or U1532 (N_1532,N_1405,N_1457);
nor U1533 (N_1533,N_1443,N_1143);
nor U1534 (N_1534,N_1380,N_1369);
and U1535 (N_1535,N_1427,N_1191);
and U1536 (N_1536,N_1112,N_1333);
and U1537 (N_1537,N_1364,N_1285);
xor U1538 (N_1538,N_1399,N_1065);
nor U1539 (N_1539,N_1250,N_1034);
nand U1540 (N_1540,N_1070,N_1392);
nor U1541 (N_1541,N_1223,N_1147);
nand U1542 (N_1542,N_1419,N_1166);
nand U1543 (N_1543,N_1275,N_1391);
xor U1544 (N_1544,N_1168,N_1347);
and U1545 (N_1545,N_1489,N_1312);
or U1546 (N_1546,N_1407,N_1353);
nor U1547 (N_1547,N_1069,N_1351);
and U1548 (N_1548,N_1087,N_1130);
nor U1549 (N_1549,N_1449,N_1175);
nor U1550 (N_1550,N_1413,N_1375);
and U1551 (N_1551,N_1182,N_1349);
xnor U1552 (N_1552,N_1122,N_1378);
nand U1553 (N_1553,N_1177,N_1207);
and U1554 (N_1554,N_1174,N_1339);
and U1555 (N_1555,N_1044,N_1459);
nor U1556 (N_1556,N_1227,N_1258);
or U1557 (N_1557,N_1136,N_1014);
nand U1558 (N_1558,N_1054,N_1160);
or U1559 (N_1559,N_1309,N_1140);
nand U1560 (N_1560,N_1079,N_1424);
or U1561 (N_1561,N_1368,N_1039);
nor U1562 (N_1562,N_1032,N_1071);
xor U1563 (N_1563,N_1067,N_1204);
or U1564 (N_1564,N_1451,N_1493);
and U1565 (N_1565,N_1420,N_1474);
nand U1566 (N_1566,N_1326,N_1441);
nor U1567 (N_1567,N_1386,N_1117);
xor U1568 (N_1568,N_1228,N_1327);
nor U1569 (N_1569,N_1211,N_1433);
xnor U1570 (N_1570,N_1479,N_1010);
nor U1571 (N_1571,N_1439,N_1161);
or U1572 (N_1572,N_1213,N_1141);
nor U1573 (N_1573,N_1450,N_1226);
nor U1574 (N_1574,N_1400,N_1476);
nor U1575 (N_1575,N_1356,N_1464);
or U1576 (N_1576,N_1195,N_1303);
nand U1577 (N_1577,N_1201,N_1317);
nor U1578 (N_1578,N_1338,N_1165);
or U1579 (N_1579,N_1164,N_1418);
nand U1580 (N_1580,N_1109,N_1167);
nand U1581 (N_1581,N_1481,N_1491);
or U1582 (N_1582,N_1005,N_1240);
and U1583 (N_1583,N_1337,N_1239);
nor U1584 (N_1584,N_1145,N_1494);
or U1585 (N_1585,N_1415,N_1422);
nor U1586 (N_1586,N_1251,N_1492);
and U1587 (N_1587,N_1119,N_1404);
nor U1588 (N_1588,N_1416,N_1301);
and U1589 (N_1589,N_1288,N_1088);
and U1590 (N_1590,N_1248,N_1273);
and U1591 (N_1591,N_1430,N_1409);
nor U1592 (N_1592,N_1472,N_1019);
or U1593 (N_1593,N_1357,N_1370);
xnor U1594 (N_1594,N_1172,N_1314);
or U1595 (N_1595,N_1390,N_1020);
or U1596 (N_1596,N_1254,N_1395);
nor U1597 (N_1597,N_1095,N_1229);
or U1598 (N_1598,N_1100,N_1015);
xnor U1599 (N_1599,N_1114,N_1125);
nand U1600 (N_1600,N_1231,N_1280);
and U1601 (N_1601,N_1307,N_1225);
nand U1602 (N_1602,N_1324,N_1061);
nor U1603 (N_1603,N_1183,N_1053);
xnor U1604 (N_1604,N_1484,N_1096);
or U1605 (N_1605,N_1209,N_1064);
nor U1606 (N_1606,N_1304,N_1490);
nor U1607 (N_1607,N_1192,N_1411);
nand U1608 (N_1608,N_1149,N_1150);
and U1609 (N_1609,N_1477,N_1076);
nor U1610 (N_1610,N_1004,N_1128);
nand U1611 (N_1611,N_1253,N_1442);
nand U1612 (N_1612,N_1387,N_1131);
nor U1613 (N_1613,N_1287,N_1292);
or U1614 (N_1614,N_1107,N_1340);
nor U1615 (N_1615,N_1097,N_1217);
nor U1616 (N_1616,N_1495,N_1296);
nand U1617 (N_1617,N_1270,N_1367);
nand U1618 (N_1618,N_1126,N_1052);
nand U1619 (N_1619,N_1268,N_1092);
xor U1620 (N_1620,N_1142,N_1233);
xor U1621 (N_1621,N_1066,N_1278);
nand U1622 (N_1622,N_1417,N_1022);
nand U1623 (N_1623,N_1403,N_1148);
or U1624 (N_1624,N_1435,N_1480);
nand U1625 (N_1625,N_1408,N_1085);
nor U1626 (N_1626,N_1041,N_1178);
or U1627 (N_1627,N_1124,N_1074);
nor U1628 (N_1628,N_1179,N_1200);
and U1629 (N_1629,N_1028,N_1487);
nand U1630 (N_1630,N_1241,N_1205);
or U1631 (N_1631,N_1075,N_1256);
nor U1632 (N_1632,N_1336,N_1138);
and U1633 (N_1633,N_1255,N_1155);
nor U1634 (N_1634,N_1452,N_1365);
nand U1635 (N_1635,N_1104,N_1198);
and U1636 (N_1636,N_1121,N_1488);
and U1637 (N_1637,N_1244,N_1388);
nand U1638 (N_1638,N_1271,N_1018);
nor U1639 (N_1639,N_1300,N_1468);
nor U1640 (N_1640,N_1453,N_1078);
nor U1641 (N_1641,N_1436,N_1421);
nor U1642 (N_1642,N_1043,N_1379);
xor U1643 (N_1643,N_1352,N_1091);
nand U1644 (N_1644,N_1219,N_1371);
and U1645 (N_1645,N_1000,N_1077);
and U1646 (N_1646,N_1084,N_1325);
nand U1647 (N_1647,N_1158,N_1058);
nor U1648 (N_1648,N_1156,N_1003);
nand U1649 (N_1649,N_1470,N_1146);
or U1650 (N_1650,N_1169,N_1006);
xnor U1651 (N_1651,N_1110,N_1106);
xnor U1652 (N_1652,N_1320,N_1343);
xor U1653 (N_1653,N_1134,N_1245);
xor U1654 (N_1654,N_1235,N_1102);
and U1655 (N_1655,N_1099,N_1033);
nand U1656 (N_1656,N_1358,N_1008);
or U1657 (N_1657,N_1050,N_1215);
and U1658 (N_1658,N_1080,N_1308);
or U1659 (N_1659,N_1259,N_1036);
and U1660 (N_1660,N_1290,N_1042);
nand U1661 (N_1661,N_1414,N_1261);
nor U1662 (N_1662,N_1344,N_1426);
nor U1663 (N_1663,N_1373,N_1382);
or U1664 (N_1664,N_1133,N_1456);
nor U1665 (N_1665,N_1446,N_1103);
nor U1666 (N_1666,N_1009,N_1318);
and U1667 (N_1667,N_1305,N_1362);
and U1668 (N_1668,N_1473,N_1483);
or U1669 (N_1669,N_1293,N_1111);
nand U1670 (N_1670,N_1499,N_1163);
and U1671 (N_1671,N_1315,N_1428);
xor U1672 (N_1672,N_1068,N_1331);
or U1673 (N_1673,N_1355,N_1321);
nand U1674 (N_1674,N_1306,N_1469);
or U1675 (N_1675,N_1072,N_1334);
or U1676 (N_1676,N_1247,N_1249);
nor U1677 (N_1677,N_1152,N_1463);
xor U1678 (N_1678,N_1299,N_1012);
and U1679 (N_1679,N_1001,N_1438);
or U1680 (N_1680,N_1218,N_1094);
and U1681 (N_1681,N_1113,N_1176);
and U1682 (N_1682,N_1366,N_1237);
and U1683 (N_1683,N_1082,N_1316);
or U1684 (N_1684,N_1011,N_1203);
or U1685 (N_1685,N_1377,N_1478);
nand U1686 (N_1686,N_1423,N_1458);
nor U1687 (N_1687,N_1289,N_1030);
and U1688 (N_1688,N_1159,N_1129);
nand U1689 (N_1689,N_1410,N_1455);
or U1690 (N_1690,N_1295,N_1381);
or U1691 (N_1691,N_1135,N_1238);
nand U1692 (N_1692,N_1144,N_1328);
and U1693 (N_1693,N_1132,N_1021);
nand U1694 (N_1694,N_1485,N_1482);
nor U1695 (N_1695,N_1497,N_1462);
nor U1696 (N_1696,N_1181,N_1398);
or U1697 (N_1697,N_1359,N_1335);
or U1698 (N_1698,N_1310,N_1434);
nor U1699 (N_1699,N_1116,N_1425);
nand U1700 (N_1700,N_1466,N_1173);
nor U1701 (N_1701,N_1447,N_1123);
or U1702 (N_1702,N_1086,N_1031);
nand U1703 (N_1703,N_1389,N_1055);
or U1704 (N_1704,N_1329,N_1486);
nor U1705 (N_1705,N_1170,N_1236);
and U1706 (N_1706,N_1199,N_1047);
nor U1707 (N_1707,N_1385,N_1297);
nand U1708 (N_1708,N_1360,N_1027);
and U1709 (N_1709,N_1242,N_1342);
nand U1710 (N_1710,N_1194,N_1396);
nor U1711 (N_1711,N_1460,N_1206);
nand U1712 (N_1712,N_1257,N_1118);
or U1713 (N_1713,N_1049,N_1465);
nor U1714 (N_1714,N_1394,N_1026);
or U1715 (N_1715,N_1286,N_1393);
nand U1716 (N_1716,N_1283,N_1397);
nand U1717 (N_1717,N_1186,N_1475);
or U1718 (N_1718,N_1332,N_1187);
or U1719 (N_1719,N_1025,N_1348);
or U1720 (N_1720,N_1224,N_1269);
nand U1721 (N_1721,N_1137,N_1212);
or U1722 (N_1722,N_1017,N_1243);
xnor U1723 (N_1723,N_1057,N_1089);
or U1724 (N_1724,N_1093,N_1037);
nor U1725 (N_1725,N_1302,N_1051);
or U1726 (N_1726,N_1221,N_1471);
xor U1727 (N_1727,N_1496,N_1277);
nand U1728 (N_1728,N_1330,N_1153);
nand U1729 (N_1729,N_1127,N_1350);
or U1730 (N_1730,N_1384,N_1298);
xnor U1731 (N_1731,N_1341,N_1222);
nor U1732 (N_1732,N_1059,N_1045);
or U1733 (N_1733,N_1431,N_1376);
or U1734 (N_1734,N_1081,N_1313);
nor U1735 (N_1735,N_1246,N_1120);
and U1736 (N_1736,N_1154,N_1202);
nand U1737 (N_1737,N_1188,N_1272);
and U1738 (N_1738,N_1311,N_1284);
or U1739 (N_1739,N_1444,N_1406);
or U1740 (N_1740,N_1282,N_1216);
nor U1741 (N_1741,N_1151,N_1171);
or U1742 (N_1742,N_1440,N_1323);
nor U1743 (N_1743,N_1498,N_1294);
nor U1744 (N_1744,N_1105,N_1232);
nor U1745 (N_1745,N_1060,N_1262);
and U1746 (N_1746,N_1197,N_1190);
or U1747 (N_1747,N_1437,N_1374);
nand U1748 (N_1748,N_1260,N_1230);
nand U1749 (N_1749,N_1185,N_1454);
nand U1750 (N_1750,N_1148,N_1249);
and U1751 (N_1751,N_1151,N_1150);
or U1752 (N_1752,N_1169,N_1352);
and U1753 (N_1753,N_1143,N_1402);
nand U1754 (N_1754,N_1262,N_1068);
xor U1755 (N_1755,N_1437,N_1338);
nand U1756 (N_1756,N_1372,N_1243);
and U1757 (N_1757,N_1272,N_1057);
nor U1758 (N_1758,N_1423,N_1171);
or U1759 (N_1759,N_1225,N_1081);
xor U1760 (N_1760,N_1226,N_1147);
or U1761 (N_1761,N_1020,N_1251);
and U1762 (N_1762,N_1233,N_1093);
and U1763 (N_1763,N_1167,N_1397);
or U1764 (N_1764,N_1201,N_1342);
nand U1765 (N_1765,N_1088,N_1350);
nor U1766 (N_1766,N_1440,N_1369);
nor U1767 (N_1767,N_1091,N_1258);
or U1768 (N_1768,N_1020,N_1209);
xnor U1769 (N_1769,N_1037,N_1090);
nand U1770 (N_1770,N_1253,N_1139);
nor U1771 (N_1771,N_1077,N_1037);
nor U1772 (N_1772,N_1361,N_1049);
nand U1773 (N_1773,N_1372,N_1491);
nand U1774 (N_1774,N_1043,N_1212);
and U1775 (N_1775,N_1255,N_1005);
nand U1776 (N_1776,N_1228,N_1091);
or U1777 (N_1777,N_1218,N_1482);
and U1778 (N_1778,N_1419,N_1232);
nand U1779 (N_1779,N_1425,N_1466);
nor U1780 (N_1780,N_1108,N_1047);
nor U1781 (N_1781,N_1459,N_1418);
and U1782 (N_1782,N_1288,N_1320);
or U1783 (N_1783,N_1171,N_1085);
and U1784 (N_1784,N_1026,N_1292);
and U1785 (N_1785,N_1220,N_1363);
nor U1786 (N_1786,N_1050,N_1052);
nor U1787 (N_1787,N_1338,N_1118);
or U1788 (N_1788,N_1129,N_1349);
and U1789 (N_1789,N_1325,N_1267);
nand U1790 (N_1790,N_1041,N_1122);
nand U1791 (N_1791,N_1470,N_1104);
or U1792 (N_1792,N_1125,N_1211);
nand U1793 (N_1793,N_1068,N_1066);
or U1794 (N_1794,N_1352,N_1089);
or U1795 (N_1795,N_1242,N_1229);
and U1796 (N_1796,N_1425,N_1364);
nor U1797 (N_1797,N_1059,N_1171);
xnor U1798 (N_1798,N_1465,N_1498);
nor U1799 (N_1799,N_1030,N_1215);
and U1800 (N_1800,N_1404,N_1474);
xnor U1801 (N_1801,N_1094,N_1353);
or U1802 (N_1802,N_1019,N_1014);
xnor U1803 (N_1803,N_1378,N_1071);
or U1804 (N_1804,N_1381,N_1253);
nand U1805 (N_1805,N_1363,N_1093);
nand U1806 (N_1806,N_1166,N_1470);
and U1807 (N_1807,N_1034,N_1343);
or U1808 (N_1808,N_1168,N_1071);
and U1809 (N_1809,N_1415,N_1098);
nor U1810 (N_1810,N_1438,N_1269);
or U1811 (N_1811,N_1053,N_1395);
and U1812 (N_1812,N_1156,N_1345);
nor U1813 (N_1813,N_1201,N_1202);
nand U1814 (N_1814,N_1175,N_1227);
and U1815 (N_1815,N_1299,N_1047);
nand U1816 (N_1816,N_1204,N_1472);
nor U1817 (N_1817,N_1385,N_1331);
nand U1818 (N_1818,N_1215,N_1104);
or U1819 (N_1819,N_1380,N_1461);
nor U1820 (N_1820,N_1497,N_1417);
nor U1821 (N_1821,N_1110,N_1368);
nand U1822 (N_1822,N_1391,N_1340);
nor U1823 (N_1823,N_1321,N_1173);
or U1824 (N_1824,N_1106,N_1465);
nor U1825 (N_1825,N_1167,N_1103);
nand U1826 (N_1826,N_1413,N_1122);
nand U1827 (N_1827,N_1122,N_1190);
or U1828 (N_1828,N_1011,N_1180);
nor U1829 (N_1829,N_1088,N_1179);
nor U1830 (N_1830,N_1100,N_1185);
or U1831 (N_1831,N_1237,N_1045);
nor U1832 (N_1832,N_1410,N_1407);
nand U1833 (N_1833,N_1059,N_1486);
nand U1834 (N_1834,N_1240,N_1081);
nand U1835 (N_1835,N_1365,N_1324);
nand U1836 (N_1836,N_1196,N_1471);
nor U1837 (N_1837,N_1383,N_1374);
nand U1838 (N_1838,N_1259,N_1488);
nor U1839 (N_1839,N_1239,N_1256);
or U1840 (N_1840,N_1426,N_1153);
xor U1841 (N_1841,N_1389,N_1483);
xnor U1842 (N_1842,N_1286,N_1475);
and U1843 (N_1843,N_1435,N_1210);
nand U1844 (N_1844,N_1258,N_1327);
or U1845 (N_1845,N_1011,N_1434);
xnor U1846 (N_1846,N_1234,N_1199);
or U1847 (N_1847,N_1418,N_1015);
nand U1848 (N_1848,N_1450,N_1214);
nand U1849 (N_1849,N_1236,N_1386);
and U1850 (N_1850,N_1408,N_1478);
nand U1851 (N_1851,N_1056,N_1271);
and U1852 (N_1852,N_1081,N_1254);
and U1853 (N_1853,N_1379,N_1128);
or U1854 (N_1854,N_1389,N_1069);
nand U1855 (N_1855,N_1484,N_1068);
xnor U1856 (N_1856,N_1340,N_1077);
nor U1857 (N_1857,N_1070,N_1063);
and U1858 (N_1858,N_1401,N_1209);
nor U1859 (N_1859,N_1426,N_1238);
and U1860 (N_1860,N_1468,N_1302);
and U1861 (N_1861,N_1194,N_1405);
or U1862 (N_1862,N_1487,N_1050);
and U1863 (N_1863,N_1117,N_1426);
nor U1864 (N_1864,N_1078,N_1236);
nand U1865 (N_1865,N_1026,N_1452);
nor U1866 (N_1866,N_1083,N_1481);
nor U1867 (N_1867,N_1062,N_1268);
or U1868 (N_1868,N_1203,N_1042);
nand U1869 (N_1869,N_1105,N_1137);
nor U1870 (N_1870,N_1135,N_1274);
nor U1871 (N_1871,N_1319,N_1363);
nor U1872 (N_1872,N_1432,N_1258);
nor U1873 (N_1873,N_1339,N_1384);
nand U1874 (N_1874,N_1386,N_1406);
or U1875 (N_1875,N_1031,N_1023);
nor U1876 (N_1876,N_1256,N_1446);
and U1877 (N_1877,N_1068,N_1435);
xnor U1878 (N_1878,N_1168,N_1118);
nand U1879 (N_1879,N_1471,N_1213);
or U1880 (N_1880,N_1411,N_1216);
and U1881 (N_1881,N_1423,N_1018);
xnor U1882 (N_1882,N_1094,N_1492);
and U1883 (N_1883,N_1322,N_1080);
nor U1884 (N_1884,N_1043,N_1163);
nand U1885 (N_1885,N_1223,N_1321);
and U1886 (N_1886,N_1273,N_1403);
and U1887 (N_1887,N_1365,N_1278);
and U1888 (N_1888,N_1249,N_1404);
xnor U1889 (N_1889,N_1194,N_1480);
nor U1890 (N_1890,N_1302,N_1248);
nand U1891 (N_1891,N_1006,N_1313);
and U1892 (N_1892,N_1060,N_1077);
nor U1893 (N_1893,N_1052,N_1448);
xnor U1894 (N_1894,N_1103,N_1398);
nor U1895 (N_1895,N_1060,N_1395);
nand U1896 (N_1896,N_1167,N_1123);
nand U1897 (N_1897,N_1453,N_1257);
nand U1898 (N_1898,N_1021,N_1430);
nor U1899 (N_1899,N_1479,N_1065);
and U1900 (N_1900,N_1349,N_1097);
nand U1901 (N_1901,N_1324,N_1008);
or U1902 (N_1902,N_1183,N_1042);
nor U1903 (N_1903,N_1112,N_1329);
nor U1904 (N_1904,N_1411,N_1488);
xnor U1905 (N_1905,N_1421,N_1015);
or U1906 (N_1906,N_1114,N_1081);
nor U1907 (N_1907,N_1104,N_1484);
and U1908 (N_1908,N_1061,N_1311);
and U1909 (N_1909,N_1265,N_1458);
xnor U1910 (N_1910,N_1373,N_1350);
nor U1911 (N_1911,N_1471,N_1455);
and U1912 (N_1912,N_1105,N_1498);
xor U1913 (N_1913,N_1406,N_1373);
nor U1914 (N_1914,N_1049,N_1084);
and U1915 (N_1915,N_1242,N_1467);
nand U1916 (N_1916,N_1213,N_1203);
or U1917 (N_1917,N_1291,N_1063);
or U1918 (N_1918,N_1179,N_1432);
and U1919 (N_1919,N_1104,N_1363);
or U1920 (N_1920,N_1426,N_1273);
and U1921 (N_1921,N_1256,N_1194);
nor U1922 (N_1922,N_1061,N_1466);
and U1923 (N_1923,N_1105,N_1196);
nand U1924 (N_1924,N_1223,N_1195);
or U1925 (N_1925,N_1445,N_1235);
and U1926 (N_1926,N_1054,N_1407);
or U1927 (N_1927,N_1471,N_1314);
xor U1928 (N_1928,N_1448,N_1132);
or U1929 (N_1929,N_1122,N_1193);
xor U1930 (N_1930,N_1425,N_1306);
nor U1931 (N_1931,N_1062,N_1227);
nand U1932 (N_1932,N_1439,N_1347);
or U1933 (N_1933,N_1217,N_1468);
xor U1934 (N_1934,N_1494,N_1128);
and U1935 (N_1935,N_1044,N_1310);
and U1936 (N_1936,N_1365,N_1176);
and U1937 (N_1937,N_1017,N_1029);
nand U1938 (N_1938,N_1019,N_1398);
and U1939 (N_1939,N_1188,N_1254);
xor U1940 (N_1940,N_1376,N_1065);
and U1941 (N_1941,N_1174,N_1442);
nor U1942 (N_1942,N_1223,N_1404);
or U1943 (N_1943,N_1204,N_1353);
xor U1944 (N_1944,N_1135,N_1029);
nand U1945 (N_1945,N_1053,N_1134);
nor U1946 (N_1946,N_1080,N_1366);
or U1947 (N_1947,N_1212,N_1342);
and U1948 (N_1948,N_1301,N_1474);
xnor U1949 (N_1949,N_1147,N_1325);
or U1950 (N_1950,N_1024,N_1239);
nand U1951 (N_1951,N_1429,N_1266);
or U1952 (N_1952,N_1280,N_1098);
nand U1953 (N_1953,N_1059,N_1129);
nand U1954 (N_1954,N_1097,N_1024);
and U1955 (N_1955,N_1175,N_1334);
nor U1956 (N_1956,N_1479,N_1300);
nor U1957 (N_1957,N_1307,N_1359);
and U1958 (N_1958,N_1463,N_1044);
nor U1959 (N_1959,N_1077,N_1231);
nor U1960 (N_1960,N_1295,N_1146);
nor U1961 (N_1961,N_1370,N_1462);
nor U1962 (N_1962,N_1225,N_1222);
nand U1963 (N_1963,N_1161,N_1212);
or U1964 (N_1964,N_1434,N_1361);
nand U1965 (N_1965,N_1253,N_1152);
and U1966 (N_1966,N_1080,N_1140);
or U1967 (N_1967,N_1319,N_1111);
and U1968 (N_1968,N_1086,N_1273);
and U1969 (N_1969,N_1115,N_1025);
and U1970 (N_1970,N_1066,N_1276);
and U1971 (N_1971,N_1253,N_1407);
or U1972 (N_1972,N_1465,N_1368);
nor U1973 (N_1973,N_1391,N_1186);
or U1974 (N_1974,N_1397,N_1241);
nand U1975 (N_1975,N_1137,N_1196);
or U1976 (N_1976,N_1390,N_1238);
nand U1977 (N_1977,N_1200,N_1496);
or U1978 (N_1978,N_1173,N_1255);
or U1979 (N_1979,N_1092,N_1279);
nand U1980 (N_1980,N_1010,N_1148);
nor U1981 (N_1981,N_1097,N_1493);
nand U1982 (N_1982,N_1304,N_1395);
and U1983 (N_1983,N_1268,N_1409);
or U1984 (N_1984,N_1182,N_1097);
xor U1985 (N_1985,N_1023,N_1337);
nand U1986 (N_1986,N_1270,N_1285);
nand U1987 (N_1987,N_1246,N_1386);
and U1988 (N_1988,N_1481,N_1029);
or U1989 (N_1989,N_1456,N_1476);
nor U1990 (N_1990,N_1170,N_1367);
xnor U1991 (N_1991,N_1096,N_1045);
nand U1992 (N_1992,N_1161,N_1226);
and U1993 (N_1993,N_1049,N_1331);
nor U1994 (N_1994,N_1338,N_1431);
nand U1995 (N_1995,N_1131,N_1045);
nor U1996 (N_1996,N_1253,N_1136);
nand U1997 (N_1997,N_1180,N_1117);
nand U1998 (N_1998,N_1308,N_1289);
nor U1999 (N_1999,N_1118,N_1228);
and U2000 (N_2000,N_1719,N_1533);
or U2001 (N_2001,N_1895,N_1590);
xor U2002 (N_2002,N_1647,N_1918);
and U2003 (N_2003,N_1829,N_1663);
nand U2004 (N_2004,N_1718,N_1591);
and U2005 (N_2005,N_1735,N_1826);
xnor U2006 (N_2006,N_1701,N_1926);
nor U2007 (N_2007,N_1705,N_1618);
nand U2008 (N_2008,N_1970,N_1715);
nand U2009 (N_2009,N_1742,N_1616);
and U2010 (N_2010,N_1642,N_1751);
nor U2011 (N_2011,N_1984,N_1631);
or U2012 (N_2012,N_1502,N_1620);
and U2013 (N_2013,N_1939,N_1828);
nand U2014 (N_2014,N_1649,N_1587);
nor U2015 (N_2015,N_1670,N_1571);
nor U2016 (N_2016,N_1917,N_1517);
nor U2017 (N_2017,N_1688,N_1986);
nor U2018 (N_2018,N_1854,N_1777);
nand U2019 (N_2019,N_1695,N_1860);
nand U2020 (N_2020,N_1504,N_1801);
and U2021 (N_2021,N_1583,N_1798);
and U2022 (N_2022,N_1942,N_1633);
nor U2023 (N_2023,N_1867,N_1919);
or U2024 (N_2024,N_1744,N_1646);
and U2025 (N_2025,N_1935,N_1645);
and U2026 (N_2026,N_1865,N_1762);
nor U2027 (N_2027,N_1643,N_1885);
nand U2028 (N_2028,N_1786,N_1545);
or U2029 (N_2029,N_1617,N_1793);
nand U2030 (N_2030,N_1522,N_1627);
and U2031 (N_2031,N_1577,N_1914);
and U2032 (N_2032,N_1888,N_1958);
and U2033 (N_2033,N_1745,N_1960);
nand U2034 (N_2034,N_1671,N_1792);
and U2035 (N_2035,N_1559,N_1610);
or U2036 (N_2036,N_1845,N_1848);
nand U2037 (N_2037,N_1922,N_1526);
nand U2038 (N_2038,N_1874,N_1853);
nor U2039 (N_2039,N_1740,N_1902);
nand U2040 (N_2040,N_1799,N_1700);
nand U2041 (N_2041,N_1875,N_1609);
nor U2042 (N_2042,N_1730,N_1698);
and U2043 (N_2043,N_1586,N_1843);
nand U2044 (N_2044,N_1995,N_1597);
and U2045 (N_2045,N_1772,N_1655);
nand U2046 (N_2046,N_1666,N_1964);
and U2047 (N_2047,N_1598,N_1934);
nand U2048 (N_2048,N_1953,N_1669);
nor U2049 (N_2049,N_1501,N_1524);
or U2050 (N_2050,N_1624,N_1813);
or U2051 (N_2051,N_1551,N_1720);
and U2052 (N_2052,N_1972,N_1776);
or U2053 (N_2053,N_1835,N_1509);
nor U2054 (N_2054,N_1552,N_1523);
xor U2055 (N_2055,N_1987,N_1863);
nand U2056 (N_2056,N_1607,N_1614);
xor U2057 (N_2057,N_1553,N_1831);
or U2058 (N_2058,N_1768,N_1941);
nor U2059 (N_2059,N_1911,N_1521);
or U2060 (N_2060,N_1750,N_1894);
and U2061 (N_2061,N_1588,N_1980);
and U2062 (N_2062,N_1778,N_1870);
nor U2063 (N_2063,N_1806,N_1928);
and U2064 (N_2064,N_1938,N_1932);
nand U2065 (N_2065,N_1575,N_1573);
nor U2066 (N_2066,N_1612,N_1743);
nor U2067 (N_2067,N_1710,N_1839);
xnor U2068 (N_2068,N_1991,N_1908);
and U2069 (N_2069,N_1725,N_1561);
or U2070 (N_2070,N_1804,N_1548);
nand U2071 (N_2071,N_1693,N_1846);
or U2072 (N_2072,N_1965,N_1789);
and U2073 (N_2073,N_1513,N_1613);
nand U2074 (N_2074,N_1738,N_1542);
and U2075 (N_2075,N_1653,N_1999);
nand U2076 (N_2076,N_1662,N_1530);
nor U2077 (N_2077,N_1706,N_1654);
and U2078 (N_2078,N_1825,N_1833);
or U2079 (N_2079,N_1503,N_1759);
and U2080 (N_2080,N_1716,N_1659);
and U2081 (N_2081,N_1557,N_1989);
nand U2082 (N_2082,N_1956,N_1723);
or U2083 (N_2083,N_1520,N_1899);
or U2084 (N_2084,N_1676,N_1873);
or U2085 (N_2085,N_1684,N_1581);
and U2086 (N_2086,N_1621,N_1982);
or U2087 (N_2087,N_1973,N_1712);
or U2088 (N_2088,N_1976,N_1962);
or U2089 (N_2089,N_1511,N_1940);
nor U2090 (N_2090,N_1808,N_1775);
nand U2091 (N_2091,N_1830,N_1696);
nand U2092 (N_2092,N_1741,N_1651);
nand U2093 (N_2093,N_1834,N_1556);
nand U2094 (N_2094,N_1547,N_1594);
and U2095 (N_2095,N_1803,N_1605);
nor U2096 (N_2096,N_1838,N_1981);
xor U2097 (N_2097,N_1998,N_1978);
and U2098 (N_2098,N_1851,N_1944);
and U2099 (N_2099,N_1857,N_1729);
nand U2100 (N_2100,N_1925,N_1817);
or U2101 (N_2101,N_1985,N_1996);
and U2102 (N_2102,N_1563,N_1736);
nor U2103 (N_2103,N_1576,N_1818);
nor U2104 (N_2104,N_1945,N_1589);
or U2105 (N_2105,N_1936,N_1623);
and U2106 (N_2106,N_1816,N_1634);
nand U2107 (N_2107,N_1680,N_1897);
and U2108 (N_2108,N_1949,N_1758);
xnor U2109 (N_2109,N_1858,N_1527);
and U2110 (N_2110,N_1794,N_1564);
nor U2111 (N_2111,N_1667,N_1550);
and U2112 (N_2112,N_1844,N_1505);
and U2113 (N_2113,N_1983,N_1820);
and U2114 (N_2114,N_1852,N_1567);
and U2115 (N_2115,N_1677,N_1931);
or U2116 (N_2116,N_1795,N_1988);
or U2117 (N_2117,N_1579,N_1927);
and U2118 (N_2118,N_1619,N_1841);
xor U2119 (N_2119,N_1967,N_1892);
or U2120 (N_2120,N_1748,N_1539);
nand U2121 (N_2121,N_1746,N_1779);
and U2122 (N_2122,N_1689,N_1668);
and U2123 (N_2123,N_1770,N_1657);
and U2124 (N_2124,N_1585,N_1815);
or U2125 (N_2125,N_1648,N_1900);
and U2126 (N_2126,N_1990,N_1787);
nor U2127 (N_2127,N_1946,N_1603);
nand U2128 (N_2128,N_1728,N_1554);
nand U2129 (N_2129,N_1652,N_1752);
nand U2130 (N_2130,N_1724,N_1969);
nor U2131 (N_2131,N_1537,N_1568);
nand U2132 (N_2132,N_1904,N_1578);
nor U2133 (N_2133,N_1766,N_1531);
and U2134 (N_2134,N_1907,N_1697);
nand U2135 (N_2135,N_1910,N_1555);
or U2136 (N_2136,N_1516,N_1544);
nand U2137 (N_2137,N_1824,N_1797);
or U2138 (N_2138,N_1543,N_1704);
or U2139 (N_2139,N_1993,N_1593);
or U2140 (N_2140,N_1933,N_1749);
nand U2141 (N_2141,N_1665,N_1507);
nor U2142 (N_2142,N_1673,N_1856);
or U2143 (N_2143,N_1699,N_1672);
and U2144 (N_2144,N_1687,N_1951);
nand U2145 (N_2145,N_1832,N_1639);
and U2146 (N_2146,N_1790,N_1562);
nor U2147 (N_2147,N_1959,N_1821);
or U2148 (N_2148,N_1781,N_1681);
and U2149 (N_2149,N_1862,N_1887);
or U2150 (N_2150,N_1871,N_1678);
nor U2151 (N_2151,N_1761,N_1727);
nand U2152 (N_2152,N_1869,N_1850);
nand U2153 (N_2153,N_1827,N_1957);
or U2154 (N_2154,N_1717,N_1558);
and U2155 (N_2155,N_1753,N_1739);
nand U2156 (N_2156,N_1569,N_1685);
xor U2157 (N_2157,N_1664,N_1915);
or U2158 (N_2158,N_1943,N_1847);
or U2159 (N_2159,N_1506,N_1679);
nor U2160 (N_2160,N_1811,N_1763);
nor U2161 (N_2161,N_1783,N_1675);
nand U2162 (N_2162,N_1515,N_1754);
and U2163 (N_2163,N_1930,N_1683);
xnor U2164 (N_2164,N_1747,N_1877);
nor U2165 (N_2165,N_1708,N_1785);
or U2166 (N_2166,N_1864,N_1534);
xor U2167 (N_2167,N_1884,N_1629);
or U2168 (N_2168,N_1674,N_1961);
nor U2169 (N_2169,N_1963,N_1582);
nand U2170 (N_2170,N_1882,N_1809);
and U2171 (N_2171,N_1630,N_1637);
and U2172 (N_2172,N_1774,N_1810);
and U2173 (N_2173,N_1912,N_1656);
nand U2174 (N_2174,N_1510,N_1968);
nand U2175 (N_2175,N_1903,N_1733);
nor U2176 (N_2176,N_1948,N_1508);
xnor U2177 (N_2177,N_1822,N_1535);
xor U2178 (N_2178,N_1755,N_1604);
xor U2179 (N_2179,N_1950,N_1566);
and U2180 (N_2180,N_1714,N_1625);
nand U2181 (N_2181,N_1893,N_1641);
nor U2182 (N_2182,N_1694,N_1879);
nand U2183 (N_2183,N_1861,N_1606);
nand U2184 (N_2184,N_1722,N_1840);
xor U2185 (N_2185,N_1916,N_1890);
or U2186 (N_2186,N_1823,N_1901);
nor U2187 (N_2187,N_1560,N_1691);
nor U2188 (N_2188,N_1954,N_1898);
nand U2189 (N_2189,N_1732,N_1686);
and U2190 (N_2190,N_1601,N_1765);
and U2191 (N_2191,N_1549,N_1541);
nand U2192 (N_2192,N_1713,N_1532);
nor U2193 (N_2193,N_1731,N_1711);
and U2194 (N_2194,N_1837,N_1660);
or U2195 (N_2195,N_1615,N_1784);
xnor U2196 (N_2196,N_1635,N_1528);
nand U2197 (N_2197,N_1538,N_1971);
or U2198 (N_2198,N_1878,N_1709);
or U2199 (N_2199,N_1909,N_1525);
xor U2200 (N_2200,N_1977,N_1905);
nand U2201 (N_2201,N_1611,N_1819);
or U2202 (N_2202,N_1979,N_1836);
or U2203 (N_2203,N_1771,N_1737);
nand U2204 (N_2204,N_1580,N_1896);
or U2205 (N_2205,N_1868,N_1937);
xnor U2206 (N_2206,N_1921,N_1807);
nor U2207 (N_2207,N_1572,N_1906);
or U2208 (N_2208,N_1628,N_1632);
and U2209 (N_2209,N_1756,N_1880);
xnor U2210 (N_2210,N_1920,N_1883);
nand U2211 (N_2211,N_1859,N_1760);
and U2212 (N_2212,N_1592,N_1872);
nor U2213 (N_2213,N_1891,N_1800);
and U2214 (N_2214,N_1682,N_1600);
nor U2215 (N_2215,N_1726,N_1791);
nor U2216 (N_2216,N_1805,N_1626);
or U2217 (N_2217,N_1570,N_1529);
nor U2218 (N_2218,N_1757,N_1886);
or U2219 (N_2219,N_1952,N_1638);
nand U2220 (N_2220,N_1947,N_1866);
xor U2221 (N_2221,N_1929,N_1661);
and U2222 (N_2222,N_1644,N_1975);
nor U2223 (N_2223,N_1734,N_1849);
and U2224 (N_2224,N_1769,N_1565);
nand U2225 (N_2225,N_1913,N_1518);
or U2226 (N_2226,N_1650,N_1796);
and U2227 (N_2227,N_1764,N_1636);
nand U2228 (N_2228,N_1596,N_1546);
nor U2229 (N_2229,N_1519,N_1812);
nand U2230 (N_2230,N_1889,N_1584);
or U2231 (N_2231,N_1640,N_1622);
xor U2232 (N_2232,N_1992,N_1788);
or U2233 (N_2233,N_1599,N_1842);
nand U2234 (N_2234,N_1924,N_1876);
xor U2235 (N_2235,N_1690,N_1923);
nand U2236 (N_2236,N_1782,N_1574);
or U2237 (N_2237,N_1608,N_1721);
or U2238 (N_2238,N_1692,N_1997);
and U2239 (N_2239,N_1780,N_1702);
or U2240 (N_2240,N_1540,N_1994);
nor U2241 (N_2241,N_1966,N_1955);
nor U2242 (N_2242,N_1881,N_1814);
nand U2243 (N_2243,N_1767,N_1602);
and U2244 (N_2244,N_1500,N_1974);
xnor U2245 (N_2245,N_1707,N_1595);
and U2246 (N_2246,N_1773,N_1802);
and U2247 (N_2247,N_1514,N_1658);
nor U2248 (N_2248,N_1536,N_1855);
nand U2249 (N_2249,N_1703,N_1512);
nor U2250 (N_2250,N_1781,N_1638);
or U2251 (N_2251,N_1798,N_1914);
xor U2252 (N_2252,N_1565,N_1590);
nor U2253 (N_2253,N_1905,N_1806);
nand U2254 (N_2254,N_1838,N_1523);
or U2255 (N_2255,N_1704,N_1808);
nor U2256 (N_2256,N_1753,N_1617);
nor U2257 (N_2257,N_1989,N_1556);
and U2258 (N_2258,N_1744,N_1633);
nor U2259 (N_2259,N_1933,N_1634);
nor U2260 (N_2260,N_1674,N_1617);
xor U2261 (N_2261,N_1943,N_1556);
xnor U2262 (N_2262,N_1735,N_1675);
and U2263 (N_2263,N_1519,N_1605);
nand U2264 (N_2264,N_1987,N_1632);
xor U2265 (N_2265,N_1593,N_1781);
xnor U2266 (N_2266,N_1724,N_1659);
or U2267 (N_2267,N_1506,N_1936);
or U2268 (N_2268,N_1811,N_1659);
nand U2269 (N_2269,N_1972,N_1628);
or U2270 (N_2270,N_1744,N_1990);
and U2271 (N_2271,N_1723,N_1760);
nor U2272 (N_2272,N_1737,N_1534);
xor U2273 (N_2273,N_1963,N_1552);
nand U2274 (N_2274,N_1973,N_1577);
and U2275 (N_2275,N_1774,N_1726);
nand U2276 (N_2276,N_1856,N_1950);
nor U2277 (N_2277,N_1611,N_1501);
or U2278 (N_2278,N_1640,N_1521);
nand U2279 (N_2279,N_1608,N_1966);
or U2280 (N_2280,N_1935,N_1585);
or U2281 (N_2281,N_1775,N_1550);
nand U2282 (N_2282,N_1851,N_1975);
and U2283 (N_2283,N_1753,N_1807);
or U2284 (N_2284,N_1888,N_1570);
nor U2285 (N_2285,N_1783,N_1609);
or U2286 (N_2286,N_1760,N_1731);
nor U2287 (N_2287,N_1901,N_1566);
or U2288 (N_2288,N_1819,N_1635);
nor U2289 (N_2289,N_1531,N_1508);
and U2290 (N_2290,N_1928,N_1603);
nand U2291 (N_2291,N_1856,N_1976);
and U2292 (N_2292,N_1822,N_1999);
and U2293 (N_2293,N_1856,N_1798);
nor U2294 (N_2294,N_1867,N_1687);
xnor U2295 (N_2295,N_1927,N_1774);
nand U2296 (N_2296,N_1846,N_1974);
nor U2297 (N_2297,N_1558,N_1764);
nand U2298 (N_2298,N_1967,N_1551);
or U2299 (N_2299,N_1579,N_1987);
nand U2300 (N_2300,N_1955,N_1912);
nand U2301 (N_2301,N_1664,N_1546);
xor U2302 (N_2302,N_1935,N_1701);
nand U2303 (N_2303,N_1989,N_1968);
nor U2304 (N_2304,N_1567,N_1858);
nand U2305 (N_2305,N_1909,N_1540);
nand U2306 (N_2306,N_1945,N_1725);
and U2307 (N_2307,N_1557,N_1721);
or U2308 (N_2308,N_1649,N_1828);
nand U2309 (N_2309,N_1576,N_1843);
nor U2310 (N_2310,N_1933,N_1842);
nor U2311 (N_2311,N_1832,N_1958);
and U2312 (N_2312,N_1697,N_1555);
or U2313 (N_2313,N_1878,N_1566);
or U2314 (N_2314,N_1801,N_1522);
and U2315 (N_2315,N_1651,N_1798);
xor U2316 (N_2316,N_1818,N_1853);
and U2317 (N_2317,N_1928,N_1934);
nand U2318 (N_2318,N_1969,N_1892);
and U2319 (N_2319,N_1958,N_1917);
nand U2320 (N_2320,N_1586,N_1888);
and U2321 (N_2321,N_1504,N_1500);
nand U2322 (N_2322,N_1979,N_1724);
and U2323 (N_2323,N_1713,N_1552);
or U2324 (N_2324,N_1978,N_1719);
and U2325 (N_2325,N_1603,N_1656);
or U2326 (N_2326,N_1722,N_1809);
nand U2327 (N_2327,N_1601,N_1988);
and U2328 (N_2328,N_1513,N_1834);
and U2329 (N_2329,N_1732,N_1932);
xor U2330 (N_2330,N_1545,N_1775);
nand U2331 (N_2331,N_1580,N_1853);
xnor U2332 (N_2332,N_1949,N_1660);
xor U2333 (N_2333,N_1697,N_1562);
nor U2334 (N_2334,N_1676,N_1723);
nor U2335 (N_2335,N_1971,N_1681);
nor U2336 (N_2336,N_1971,N_1731);
or U2337 (N_2337,N_1688,N_1844);
nand U2338 (N_2338,N_1706,N_1808);
or U2339 (N_2339,N_1698,N_1965);
nand U2340 (N_2340,N_1893,N_1590);
or U2341 (N_2341,N_1830,N_1536);
nand U2342 (N_2342,N_1759,N_1908);
and U2343 (N_2343,N_1566,N_1734);
nor U2344 (N_2344,N_1604,N_1672);
or U2345 (N_2345,N_1723,N_1524);
nand U2346 (N_2346,N_1771,N_1544);
xnor U2347 (N_2347,N_1516,N_1641);
nor U2348 (N_2348,N_1730,N_1922);
or U2349 (N_2349,N_1880,N_1927);
nor U2350 (N_2350,N_1862,N_1936);
nor U2351 (N_2351,N_1975,N_1780);
or U2352 (N_2352,N_1660,N_1621);
nand U2353 (N_2353,N_1653,N_1529);
or U2354 (N_2354,N_1744,N_1985);
nor U2355 (N_2355,N_1908,N_1976);
nand U2356 (N_2356,N_1917,N_1526);
xnor U2357 (N_2357,N_1724,N_1997);
nor U2358 (N_2358,N_1948,N_1815);
xor U2359 (N_2359,N_1785,N_1613);
nand U2360 (N_2360,N_1525,N_1743);
nor U2361 (N_2361,N_1608,N_1942);
xnor U2362 (N_2362,N_1509,N_1722);
or U2363 (N_2363,N_1575,N_1987);
or U2364 (N_2364,N_1517,N_1683);
nor U2365 (N_2365,N_1770,N_1636);
and U2366 (N_2366,N_1598,N_1605);
or U2367 (N_2367,N_1921,N_1874);
nor U2368 (N_2368,N_1844,N_1735);
nor U2369 (N_2369,N_1505,N_1661);
or U2370 (N_2370,N_1769,N_1949);
or U2371 (N_2371,N_1989,N_1967);
xor U2372 (N_2372,N_1784,N_1516);
and U2373 (N_2373,N_1764,N_1883);
or U2374 (N_2374,N_1800,N_1607);
or U2375 (N_2375,N_1887,N_1952);
xnor U2376 (N_2376,N_1701,N_1662);
nor U2377 (N_2377,N_1517,N_1718);
nor U2378 (N_2378,N_1919,N_1620);
nand U2379 (N_2379,N_1822,N_1750);
nor U2380 (N_2380,N_1764,N_1921);
xor U2381 (N_2381,N_1985,N_1888);
or U2382 (N_2382,N_1943,N_1625);
and U2383 (N_2383,N_1857,N_1676);
nor U2384 (N_2384,N_1741,N_1641);
or U2385 (N_2385,N_1928,N_1598);
or U2386 (N_2386,N_1957,N_1744);
and U2387 (N_2387,N_1899,N_1668);
and U2388 (N_2388,N_1923,N_1654);
and U2389 (N_2389,N_1558,N_1756);
or U2390 (N_2390,N_1823,N_1687);
or U2391 (N_2391,N_1608,N_1565);
nor U2392 (N_2392,N_1515,N_1758);
nor U2393 (N_2393,N_1900,N_1977);
nor U2394 (N_2394,N_1727,N_1965);
or U2395 (N_2395,N_1527,N_1565);
and U2396 (N_2396,N_1690,N_1888);
nor U2397 (N_2397,N_1791,N_1543);
or U2398 (N_2398,N_1645,N_1806);
xor U2399 (N_2399,N_1973,N_1588);
nor U2400 (N_2400,N_1652,N_1591);
nor U2401 (N_2401,N_1957,N_1749);
xor U2402 (N_2402,N_1753,N_1741);
xnor U2403 (N_2403,N_1635,N_1597);
or U2404 (N_2404,N_1643,N_1965);
nor U2405 (N_2405,N_1811,N_1884);
and U2406 (N_2406,N_1931,N_1792);
and U2407 (N_2407,N_1668,N_1620);
or U2408 (N_2408,N_1546,N_1954);
xor U2409 (N_2409,N_1926,N_1513);
nor U2410 (N_2410,N_1829,N_1511);
or U2411 (N_2411,N_1606,N_1864);
nor U2412 (N_2412,N_1751,N_1580);
nor U2413 (N_2413,N_1703,N_1811);
nor U2414 (N_2414,N_1606,N_1601);
or U2415 (N_2415,N_1915,N_1716);
or U2416 (N_2416,N_1775,N_1976);
xnor U2417 (N_2417,N_1712,N_1637);
nand U2418 (N_2418,N_1971,N_1582);
and U2419 (N_2419,N_1903,N_1781);
and U2420 (N_2420,N_1566,N_1654);
and U2421 (N_2421,N_1893,N_1817);
nor U2422 (N_2422,N_1710,N_1802);
nor U2423 (N_2423,N_1519,N_1598);
nor U2424 (N_2424,N_1551,N_1819);
and U2425 (N_2425,N_1687,N_1733);
nand U2426 (N_2426,N_1723,N_1935);
or U2427 (N_2427,N_1634,N_1554);
or U2428 (N_2428,N_1841,N_1618);
nor U2429 (N_2429,N_1514,N_1969);
or U2430 (N_2430,N_1958,N_1997);
and U2431 (N_2431,N_1529,N_1760);
or U2432 (N_2432,N_1771,N_1822);
nand U2433 (N_2433,N_1959,N_1738);
or U2434 (N_2434,N_1884,N_1646);
nand U2435 (N_2435,N_1909,N_1889);
nor U2436 (N_2436,N_1967,N_1738);
or U2437 (N_2437,N_1614,N_1783);
or U2438 (N_2438,N_1511,N_1964);
and U2439 (N_2439,N_1620,N_1603);
nand U2440 (N_2440,N_1899,N_1504);
nand U2441 (N_2441,N_1610,N_1964);
nand U2442 (N_2442,N_1626,N_1955);
and U2443 (N_2443,N_1596,N_1741);
and U2444 (N_2444,N_1642,N_1590);
and U2445 (N_2445,N_1764,N_1847);
nand U2446 (N_2446,N_1531,N_1717);
nand U2447 (N_2447,N_1938,N_1521);
xor U2448 (N_2448,N_1626,N_1716);
or U2449 (N_2449,N_1849,N_1954);
and U2450 (N_2450,N_1866,N_1561);
xnor U2451 (N_2451,N_1706,N_1957);
or U2452 (N_2452,N_1639,N_1528);
and U2453 (N_2453,N_1950,N_1714);
xnor U2454 (N_2454,N_1582,N_1680);
nor U2455 (N_2455,N_1923,N_1999);
xor U2456 (N_2456,N_1561,N_1879);
and U2457 (N_2457,N_1588,N_1638);
xor U2458 (N_2458,N_1621,N_1932);
and U2459 (N_2459,N_1801,N_1502);
and U2460 (N_2460,N_1929,N_1530);
or U2461 (N_2461,N_1709,N_1571);
or U2462 (N_2462,N_1750,N_1780);
and U2463 (N_2463,N_1509,N_1595);
nor U2464 (N_2464,N_1914,N_1658);
nor U2465 (N_2465,N_1938,N_1961);
or U2466 (N_2466,N_1999,N_1525);
or U2467 (N_2467,N_1991,N_1602);
nand U2468 (N_2468,N_1502,N_1657);
and U2469 (N_2469,N_1652,N_1695);
and U2470 (N_2470,N_1952,N_1589);
and U2471 (N_2471,N_1759,N_1603);
nor U2472 (N_2472,N_1588,N_1832);
nand U2473 (N_2473,N_1647,N_1766);
nor U2474 (N_2474,N_1661,N_1906);
xnor U2475 (N_2475,N_1767,N_1986);
nor U2476 (N_2476,N_1710,N_1963);
nor U2477 (N_2477,N_1771,N_1538);
or U2478 (N_2478,N_1919,N_1836);
or U2479 (N_2479,N_1626,N_1771);
or U2480 (N_2480,N_1907,N_1532);
xor U2481 (N_2481,N_1948,N_1740);
nor U2482 (N_2482,N_1975,N_1863);
and U2483 (N_2483,N_1559,N_1699);
nand U2484 (N_2484,N_1696,N_1545);
nor U2485 (N_2485,N_1782,N_1656);
nand U2486 (N_2486,N_1648,N_1612);
or U2487 (N_2487,N_1542,N_1587);
nand U2488 (N_2488,N_1651,N_1818);
and U2489 (N_2489,N_1803,N_1814);
or U2490 (N_2490,N_1985,N_1603);
nor U2491 (N_2491,N_1940,N_1996);
or U2492 (N_2492,N_1749,N_1687);
and U2493 (N_2493,N_1615,N_1533);
nand U2494 (N_2494,N_1607,N_1636);
nor U2495 (N_2495,N_1546,N_1914);
and U2496 (N_2496,N_1865,N_1635);
nor U2497 (N_2497,N_1771,N_1752);
nor U2498 (N_2498,N_1920,N_1787);
or U2499 (N_2499,N_1678,N_1675);
and U2500 (N_2500,N_2490,N_2400);
or U2501 (N_2501,N_2079,N_2371);
and U2502 (N_2502,N_2018,N_2238);
nand U2503 (N_2503,N_2463,N_2289);
nor U2504 (N_2504,N_2432,N_2270);
nand U2505 (N_2505,N_2235,N_2358);
nor U2506 (N_2506,N_2337,N_2007);
nor U2507 (N_2507,N_2058,N_2187);
and U2508 (N_2508,N_2468,N_2327);
nand U2509 (N_2509,N_2478,N_2475);
or U2510 (N_2510,N_2210,N_2294);
nand U2511 (N_2511,N_2341,N_2301);
nand U2512 (N_2512,N_2039,N_2375);
and U2513 (N_2513,N_2143,N_2183);
nand U2514 (N_2514,N_2394,N_2448);
or U2515 (N_2515,N_2022,N_2196);
nor U2516 (N_2516,N_2125,N_2258);
nor U2517 (N_2517,N_2250,N_2055);
or U2518 (N_2518,N_2174,N_2360);
nand U2519 (N_2519,N_2180,N_2488);
nor U2520 (N_2520,N_2128,N_2090);
and U2521 (N_2521,N_2267,N_2252);
nand U2522 (N_2522,N_2446,N_2229);
or U2523 (N_2523,N_2461,N_2160);
nand U2524 (N_2524,N_2356,N_2362);
or U2525 (N_2525,N_2081,N_2111);
or U2526 (N_2526,N_2037,N_2479);
nand U2527 (N_2527,N_2170,N_2156);
or U2528 (N_2528,N_2257,N_2395);
or U2529 (N_2529,N_2094,N_2197);
nor U2530 (N_2530,N_2287,N_2189);
xor U2531 (N_2531,N_2036,N_2265);
or U2532 (N_2532,N_2142,N_2054);
or U2533 (N_2533,N_2398,N_2165);
nor U2534 (N_2534,N_2012,N_2135);
or U2535 (N_2535,N_2099,N_2422);
nor U2536 (N_2536,N_2164,N_2199);
nor U2537 (N_2537,N_2304,N_2239);
nor U2538 (N_2538,N_2254,N_2122);
nand U2539 (N_2539,N_2149,N_2323);
and U2540 (N_2540,N_2025,N_2438);
xor U2541 (N_2541,N_2086,N_2065);
xnor U2542 (N_2542,N_2224,N_2480);
and U2543 (N_2543,N_2218,N_2179);
nor U2544 (N_2544,N_2038,N_2083);
nor U2545 (N_2545,N_2487,N_2281);
nor U2546 (N_2546,N_2013,N_2373);
and U2547 (N_2547,N_2017,N_2279);
nand U2548 (N_2548,N_2391,N_2310);
nand U2549 (N_2549,N_2009,N_2466);
or U2550 (N_2550,N_2280,N_2469);
or U2551 (N_2551,N_2060,N_2137);
and U2552 (N_2552,N_2455,N_2228);
nand U2553 (N_2553,N_2417,N_2109);
xnor U2554 (N_2554,N_2473,N_2464);
nor U2555 (N_2555,N_2155,N_2350);
nand U2556 (N_2556,N_2100,N_2130);
nand U2557 (N_2557,N_2406,N_2368);
nand U2558 (N_2558,N_2144,N_2117);
nand U2559 (N_2559,N_2256,N_2393);
or U2560 (N_2560,N_2316,N_2233);
nand U2561 (N_2561,N_2451,N_2336);
and U2562 (N_2562,N_2127,N_2011);
nor U2563 (N_2563,N_2452,N_2282);
nor U2564 (N_2564,N_2416,N_2383);
or U2565 (N_2565,N_2484,N_2205);
nor U2566 (N_2566,N_2177,N_2061);
nor U2567 (N_2567,N_2277,N_2253);
and U2568 (N_2568,N_2425,N_2110);
xnor U2569 (N_2569,N_2440,N_2107);
and U2570 (N_2570,N_2001,N_2420);
nor U2571 (N_2571,N_2049,N_2274);
nor U2572 (N_2572,N_2048,N_2077);
or U2573 (N_2573,N_2296,N_2275);
and U2574 (N_2574,N_2412,N_2331);
or U2575 (N_2575,N_2016,N_2088);
xnor U2576 (N_2576,N_2115,N_2151);
and U2577 (N_2577,N_2119,N_2000);
nor U2578 (N_2578,N_2105,N_2476);
nor U2579 (N_2579,N_2114,N_2098);
and U2580 (N_2580,N_2486,N_2171);
and U2581 (N_2581,N_2159,N_2329);
or U2582 (N_2582,N_2147,N_2133);
nor U2583 (N_2583,N_2184,N_2194);
nor U2584 (N_2584,N_2146,N_2450);
nor U2585 (N_2585,N_2093,N_2046);
and U2586 (N_2586,N_2070,N_2351);
nand U2587 (N_2587,N_2365,N_2315);
nand U2588 (N_2588,N_2053,N_2186);
nand U2589 (N_2589,N_2374,N_2328);
or U2590 (N_2590,N_2101,N_2421);
or U2591 (N_2591,N_2414,N_2104);
nor U2592 (N_2592,N_2231,N_2401);
nor U2593 (N_2593,N_2206,N_2349);
and U2594 (N_2594,N_2169,N_2405);
nand U2595 (N_2595,N_2008,N_2162);
or U2596 (N_2596,N_2424,N_2284);
or U2597 (N_2597,N_2116,N_2106);
or U2598 (N_2598,N_2069,N_2261);
and U2599 (N_2599,N_2278,N_2215);
nand U2600 (N_2600,N_2091,N_2260);
nand U2601 (N_2601,N_2345,N_2191);
and U2602 (N_2602,N_2392,N_2047);
nand U2603 (N_2603,N_2407,N_2439);
and U2604 (N_2604,N_2458,N_2010);
and U2605 (N_2605,N_2491,N_2321);
xnor U2606 (N_2606,N_2176,N_2259);
xor U2607 (N_2607,N_2057,N_2029);
nand U2608 (N_2608,N_2302,N_2471);
nor U2609 (N_2609,N_2353,N_2059);
and U2610 (N_2610,N_2166,N_2474);
xnor U2611 (N_2611,N_2234,N_2410);
and U2612 (N_2612,N_2467,N_2385);
xor U2613 (N_2613,N_2326,N_2409);
and U2614 (N_2614,N_2330,N_2207);
nor U2615 (N_2615,N_2482,N_2141);
nand U2616 (N_2616,N_2499,N_2245);
or U2617 (N_2617,N_2071,N_2064);
nor U2618 (N_2618,N_2121,N_2495);
xor U2619 (N_2619,N_2472,N_2002);
nor U2620 (N_2620,N_2300,N_2095);
nor U2621 (N_2621,N_2370,N_2102);
xor U2622 (N_2622,N_2092,N_2271);
nor U2623 (N_2623,N_2023,N_2050);
nand U2624 (N_2624,N_2209,N_2340);
nor U2625 (N_2625,N_2158,N_2028);
xor U2626 (N_2626,N_2042,N_2223);
nand U2627 (N_2627,N_2457,N_2359);
xor U2628 (N_2628,N_2402,N_2444);
and U2629 (N_2629,N_2066,N_2443);
or U2630 (N_2630,N_2434,N_2283);
xnor U2631 (N_2631,N_2247,N_2449);
xor U2632 (N_2632,N_2033,N_2355);
nand U2633 (N_2633,N_2150,N_2306);
or U2634 (N_2634,N_2230,N_2322);
xor U2635 (N_2635,N_2273,N_2226);
nand U2636 (N_2636,N_2136,N_2052);
or U2637 (N_2637,N_2388,N_2041);
nand U2638 (N_2638,N_2390,N_2411);
nand U2639 (N_2639,N_2242,N_2477);
nor U2640 (N_2640,N_2335,N_2295);
nor U2641 (N_2641,N_2297,N_2404);
and U2642 (N_2642,N_2222,N_2132);
nand U2643 (N_2643,N_2369,N_2276);
nor U2644 (N_2644,N_2292,N_2485);
or U2645 (N_2645,N_2334,N_2056);
nand U2646 (N_2646,N_2386,N_2173);
and U2647 (N_2647,N_2080,N_2481);
and U2648 (N_2648,N_2408,N_2266);
or U2649 (N_2649,N_2318,N_2342);
nand U2650 (N_2650,N_2427,N_2379);
or U2651 (N_2651,N_2442,N_2040);
or U2652 (N_2652,N_2441,N_2377);
nand U2653 (N_2653,N_2465,N_2225);
nor U2654 (N_2654,N_2437,N_2154);
and U2655 (N_2655,N_2131,N_2163);
xnor U2656 (N_2656,N_2399,N_2435);
or U2657 (N_2657,N_2241,N_2268);
and U2658 (N_2658,N_2493,N_2462);
and U2659 (N_2659,N_2456,N_2195);
nand U2660 (N_2660,N_2181,N_2324);
nor U2661 (N_2661,N_2338,N_2354);
or U2662 (N_2662,N_2303,N_2497);
and U2663 (N_2663,N_2243,N_2138);
nand U2664 (N_2664,N_2494,N_2293);
nor U2665 (N_2665,N_2062,N_2063);
nor U2666 (N_2666,N_2445,N_2248);
nand U2667 (N_2667,N_2212,N_2214);
nor U2668 (N_2668,N_2015,N_2286);
and U2669 (N_2669,N_2262,N_2249);
nor U2670 (N_2670,N_2357,N_2019);
nand U2671 (N_2671,N_2403,N_2044);
or U2672 (N_2672,N_2367,N_2307);
nand U2673 (N_2673,N_2034,N_2032);
and U2674 (N_2674,N_2237,N_2182);
nor U2675 (N_2675,N_2496,N_2285);
or U2676 (N_2676,N_2072,N_2087);
nor U2677 (N_2677,N_2382,N_2024);
and U2678 (N_2678,N_2004,N_2255);
nor U2679 (N_2679,N_2168,N_2067);
nand U2680 (N_2680,N_2103,N_2026);
and U2681 (N_2681,N_2118,N_2112);
nor U2682 (N_2682,N_2352,N_2298);
xor U2683 (N_2683,N_2263,N_2175);
nor U2684 (N_2684,N_2498,N_2120);
xnor U2685 (N_2685,N_2188,N_2311);
and U2686 (N_2686,N_2244,N_2030);
nand U2687 (N_2687,N_2363,N_2314);
or U2688 (N_2688,N_2246,N_2430);
and U2689 (N_2689,N_2227,N_2193);
nor U2690 (N_2690,N_2460,N_2021);
nand U2691 (N_2691,N_2006,N_2167);
or U2692 (N_2692,N_2074,N_2423);
or U2693 (N_2693,N_2178,N_2236);
and U2694 (N_2694,N_2433,N_2202);
or U2695 (N_2695,N_2190,N_2346);
nand U2696 (N_2696,N_2126,N_2251);
and U2697 (N_2697,N_2387,N_2113);
nand U2698 (N_2698,N_2372,N_2208);
nand U2699 (N_2699,N_2313,N_2076);
nor U2700 (N_2700,N_2459,N_2108);
and U2701 (N_2701,N_2361,N_2453);
xor U2702 (N_2702,N_2145,N_2198);
nand U2703 (N_2703,N_2211,N_2389);
xnor U2704 (N_2704,N_2419,N_2157);
and U2705 (N_2705,N_2454,N_2045);
nor U2706 (N_2706,N_2123,N_2380);
or U2707 (N_2707,N_2172,N_2470);
and U2708 (N_2708,N_2429,N_2290);
nor U2709 (N_2709,N_2082,N_2068);
xnor U2710 (N_2710,N_2384,N_2129);
nand U2711 (N_2711,N_2483,N_2027);
nor U2712 (N_2712,N_2291,N_2161);
nand U2713 (N_2713,N_2005,N_2348);
nor U2714 (N_2714,N_2192,N_2381);
nand U2715 (N_2715,N_2085,N_2139);
nand U2716 (N_2716,N_2232,N_2084);
and U2717 (N_2717,N_2343,N_2221);
or U2718 (N_2718,N_2344,N_2319);
or U2719 (N_2719,N_2204,N_2378);
or U2720 (N_2720,N_2134,N_2185);
and U2721 (N_2721,N_2317,N_2031);
and U2722 (N_2722,N_2020,N_2299);
nand U2723 (N_2723,N_2272,N_2124);
and U2724 (N_2724,N_2320,N_2153);
nand U2725 (N_2725,N_2152,N_2431);
and U2726 (N_2726,N_2305,N_2075);
and U2727 (N_2727,N_2413,N_2489);
xnor U2728 (N_2728,N_2428,N_2217);
xor U2729 (N_2729,N_2325,N_2097);
or U2730 (N_2730,N_2269,N_2312);
and U2731 (N_2731,N_2418,N_2366);
or U2732 (N_2732,N_2347,N_2014);
nor U2733 (N_2733,N_2043,N_2240);
xnor U2734 (N_2734,N_2308,N_2333);
and U2735 (N_2735,N_2309,N_2213);
nand U2736 (N_2736,N_2426,N_2436);
nand U2737 (N_2737,N_2264,N_2339);
and U2738 (N_2738,N_2200,N_2203);
and U2739 (N_2739,N_2220,N_2148);
nand U2740 (N_2740,N_2003,N_2332);
or U2741 (N_2741,N_2216,N_2089);
xor U2742 (N_2742,N_2397,N_2415);
xor U2743 (N_2743,N_2376,N_2078);
nand U2744 (N_2744,N_2364,N_2396);
nand U2745 (N_2745,N_2140,N_2035);
xnor U2746 (N_2746,N_2096,N_2447);
nor U2747 (N_2747,N_2073,N_2492);
nand U2748 (N_2748,N_2219,N_2201);
nand U2749 (N_2749,N_2288,N_2051);
and U2750 (N_2750,N_2145,N_2420);
nand U2751 (N_2751,N_2248,N_2044);
nor U2752 (N_2752,N_2224,N_2119);
nor U2753 (N_2753,N_2101,N_2371);
or U2754 (N_2754,N_2297,N_2339);
or U2755 (N_2755,N_2048,N_2116);
or U2756 (N_2756,N_2284,N_2477);
or U2757 (N_2757,N_2306,N_2281);
nand U2758 (N_2758,N_2136,N_2054);
nor U2759 (N_2759,N_2293,N_2180);
nor U2760 (N_2760,N_2060,N_2361);
xnor U2761 (N_2761,N_2406,N_2090);
nor U2762 (N_2762,N_2374,N_2383);
or U2763 (N_2763,N_2488,N_2469);
or U2764 (N_2764,N_2007,N_2408);
nor U2765 (N_2765,N_2059,N_2335);
nor U2766 (N_2766,N_2026,N_2291);
nor U2767 (N_2767,N_2263,N_2126);
nor U2768 (N_2768,N_2144,N_2409);
and U2769 (N_2769,N_2373,N_2398);
and U2770 (N_2770,N_2187,N_2386);
nand U2771 (N_2771,N_2143,N_2320);
and U2772 (N_2772,N_2341,N_2234);
and U2773 (N_2773,N_2106,N_2416);
nor U2774 (N_2774,N_2382,N_2139);
nand U2775 (N_2775,N_2431,N_2161);
or U2776 (N_2776,N_2103,N_2273);
nor U2777 (N_2777,N_2346,N_2229);
nor U2778 (N_2778,N_2064,N_2469);
nand U2779 (N_2779,N_2497,N_2294);
xnor U2780 (N_2780,N_2494,N_2137);
nand U2781 (N_2781,N_2424,N_2085);
nor U2782 (N_2782,N_2352,N_2274);
nor U2783 (N_2783,N_2308,N_2343);
nand U2784 (N_2784,N_2402,N_2497);
and U2785 (N_2785,N_2192,N_2258);
nand U2786 (N_2786,N_2457,N_2267);
nand U2787 (N_2787,N_2362,N_2051);
or U2788 (N_2788,N_2380,N_2133);
xnor U2789 (N_2789,N_2484,N_2476);
or U2790 (N_2790,N_2116,N_2045);
nand U2791 (N_2791,N_2430,N_2389);
or U2792 (N_2792,N_2087,N_2357);
or U2793 (N_2793,N_2036,N_2458);
and U2794 (N_2794,N_2293,N_2370);
nor U2795 (N_2795,N_2163,N_2237);
nand U2796 (N_2796,N_2351,N_2168);
and U2797 (N_2797,N_2357,N_2222);
nor U2798 (N_2798,N_2107,N_2315);
and U2799 (N_2799,N_2361,N_2006);
or U2800 (N_2800,N_2115,N_2288);
nor U2801 (N_2801,N_2169,N_2047);
nor U2802 (N_2802,N_2377,N_2273);
nor U2803 (N_2803,N_2110,N_2001);
or U2804 (N_2804,N_2011,N_2136);
nor U2805 (N_2805,N_2067,N_2466);
nor U2806 (N_2806,N_2119,N_2106);
and U2807 (N_2807,N_2433,N_2495);
or U2808 (N_2808,N_2330,N_2205);
nor U2809 (N_2809,N_2339,N_2160);
nor U2810 (N_2810,N_2435,N_2142);
nor U2811 (N_2811,N_2453,N_2157);
or U2812 (N_2812,N_2177,N_2484);
nor U2813 (N_2813,N_2476,N_2470);
nor U2814 (N_2814,N_2443,N_2171);
and U2815 (N_2815,N_2116,N_2071);
nand U2816 (N_2816,N_2070,N_2422);
nand U2817 (N_2817,N_2025,N_2340);
nor U2818 (N_2818,N_2143,N_2157);
or U2819 (N_2819,N_2119,N_2170);
or U2820 (N_2820,N_2383,N_2492);
and U2821 (N_2821,N_2282,N_2044);
or U2822 (N_2822,N_2150,N_2017);
or U2823 (N_2823,N_2166,N_2203);
nor U2824 (N_2824,N_2131,N_2169);
or U2825 (N_2825,N_2024,N_2265);
nor U2826 (N_2826,N_2077,N_2012);
or U2827 (N_2827,N_2360,N_2235);
xnor U2828 (N_2828,N_2376,N_2035);
nand U2829 (N_2829,N_2450,N_2441);
or U2830 (N_2830,N_2483,N_2458);
and U2831 (N_2831,N_2139,N_2410);
or U2832 (N_2832,N_2425,N_2467);
nor U2833 (N_2833,N_2381,N_2055);
or U2834 (N_2834,N_2432,N_2148);
nand U2835 (N_2835,N_2047,N_2241);
nand U2836 (N_2836,N_2005,N_2139);
and U2837 (N_2837,N_2268,N_2105);
nor U2838 (N_2838,N_2140,N_2233);
nor U2839 (N_2839,N_2109,N_2279);
nand U2840 (N_2840,N_2136,N_2357);
and U2841 (N_2841,N_2435,N_2059);
nand U2842 (N_2842,N_2010,N_2367);
nand U2843 (N_2843,N_2065,N_2261);
and U2844 (N_2844,N_2195,N_2233);
and U2845 (N_2845,N_2285,N_2336);
and U2846 (N_2846,N_2310,N_2404);
or U2847 (N_2847,N_2088,N_2477);
or U2848 (N_2848,N_2456,N_2197);
and U2849 (N_2849,N_2407,N_2062);
nand U2850 (N_2850,N_2095,N_2001);
xor U2851 (N_2851,N_2249,N_2411);
and U2852 (N_2852,N_2372,N_2285);
nand U2853 (N_2853,N_2144,N_2251);
nand U2854 (N_2854,N_2415,N_2055);
nor U2855 (N_2855,N_2439,N_2272);
nand U2856 (N_2856,N_2411,N_2156);
nor U2857 (N_2857,N_2132,N_2320);
nor U2858 (N_2858,N_2097,N_2078);
xnor U2859 (N_2859,N_2023,N_2293);
nand U2860 (N_2860,N_2037,N_2053);
nor U2861 (N_2861,N_2295,N_2177);
nor U2862 (N_2862,N_2314,N_2162);
or U2863 (N_2863,N_2459,N_2045);
and U2864 (N_2864,N_2310,N_2238);
xor U2865 (N_2865,N_2249,N_2271);
and U2866 (N_2866,N_2329,N_2040);
nor U2867 (N_2867,N_2283,N_2498);
or U2868 (N_2868,N_2088,N_2039);
and U2869 (N_2869,N_2242,N_2133);
or U2870 (N_2870,N_2116,N_2118);
nor U2871 (N_2871,N_2453,N_2414);
nand U2872 (N_2872,N_2095,N_2141);
nand U2873 (N_2873,N_2466,N_2228);
or U2874 (N_2874,N_2451,N_2253);
nor U2875 (N_2875,N_2445,N_2334);
or U2876 (N_2876,N_2195,N_2144);
nor U2877 (N_2877,N_2026,N_2302);
and U2878 (N_2878,N_2288,N_2272);
and U2879 (N_2879,N_2327,N_2314);
and U2880 (N_2880,N_2299,N_2022);
or U2881 (N_2881,N_2087,N_2410);
or U2882 (N_2882,N_2440,N_2279);
or U2883 (N_2883,N_2468,N_2046);
nand U2884 (N_2884,N_2185,N_2443);
and U2885 (N_2885,N_2194,N_2412);
nor U2886 (N_2886,N_2167,N_2043);
xnor U2887 (N_2887,N_2066,N_2213);
nand U2888 (N_2888,N_2345,N_2153);
or U2889 (N_2889,N_2192,N_2459);
or U2890 (N_2890,N_2111,N_2440);
or U2891 (N_2891,N_2352,N_2241);
and U2892 (N_2892,N_2103,N_2202);
nor U2893 (N_2893,N_2272,N_2097);
and U2894 (N_2894,N_2040,N_2072);
nand U2895 (N_2895,N_2191,N_2422);
or U2896 (N_2896,N_2229,N_2284);
nand U2897 (N_2897,N_2057,N_2459);
and U2898 (N_2898,N_2295,N_2031);
and U2899 (N_2899,N_2060,N_2192);
or U2900 (N_2900,N_2070,N_2287);
xnor U2901 (N_2901,N_2000,N_2488);
or U2902 (N_2902,N_2426,N_2392);
or U2903 (N_2903,N_2359,N_2408);
nor U2904 (N_2904,N_2210,N_2401);
nor U2905 (N_2905,N_2238,N_2228);
nand U2906 (N_2906,N_2278,N_2463);
or U2907 (N_2907,N_2080,N_2419);
nor U2908 (N_2908,N_2325,N_2442);
nor U2909 (N_2909,N_2414,N_2034);
nor U2910 (N_2910,N_2327,N_2284);
nor U2911 (N_2911,N_2340,N_2208);
and U2912 (N_2912,N_2060,N_2127);
or U2913 (N_2913,N_2295,N_2433);
nor U2914 (N_2914,N_2074,N_2214);
nor U2915 (N_2915,N_2498,N_2465);
or U2916 (N_2916,N_2234,N_2414);
and U2917 (N_2917,N_2389,N_2320);
and U2918 (N_2918,N_2007,N_2310);
and U2919 (N_2919,N_2416,N_2422);
or U2920 (N_2920,N_2210,N_2344);
and U2921 (N_2921,N_2366,N_2245);
and U2922 (N_2922,N_2423,N_2015);
nor U2923 (N_2923,N_2382,N_2287);
or U2924 (N_2924,N_2171,N_2063);
or U2925 (N_2925,N_2002,N_2036);
and U2926 (N_2926,N_2007,N_2042);
or U2927 (N_2927,N_2468,N_2182);
nor U2928 (N_2928,N_2297,N_2370);
or U2929 (N_2929,N_2262,N_2363);
or U2930 (N_2930,N_2030,N_2044);
or U2931 (N_2931,N_2407,N_2441);
nor U2932 (N_2932,N_2301,N_2435);
nor U2933 (N_2933,N_2357,N_2145);
xnor U2934 (N_2934,N_2495,N_2139);
nand U2935 (N_2935,N_2154,N_2415);
nor U2936 (N_2936,N_2156,N_2225);
nand U2937 (N_2937,N_2169,N_2343);
nand U2938 (N_2938,N_2104,N_2379);
or U2939 (N_2939,N_2047,N_2466);
nor U2940 (N_2940,N_2128,N_2351);
nor U2941 (N_2941,N_2071,N_2267);
or U2942 (N_2942,N_2067,N_2110);
or U2943 (N_2943,N_2359,N_2002);
and U2944 (N_2944,N_2418,N_2328);
or U2945 (N_2945,N_2079,N_2297);
nor U2946 (N_2946,N_2226,N_2132);
and U2947 (N_2947,N_2381,N_2136);
or U2948 (N_2948,N_2266,N_2491);
xor U2949 (N_2949,N_2447,N_2292);
and U2950 (N_2950,N_2291,N_2261);
and U2951 (N_2951,N_2365,N_2279);
xor U2952 (N_2952,N_2173,N_2322);
and U2953 (N_2953,N_2098,N_2491);
nand U2954 (N_2954,N_2235,N_2314);
nand U2955 (N_2955,N_2057,N_2103);
and U2956 (N_2956,N_2192,N_2035);
and U2957 (N_2957,N_2468,N_2139);
nand U2958 (N_2958,N_2279,N_2415);
xor U2959 (N_2959,N_2069,N_2363);
or U2960 (N_2960,N_2287,N_2338);
nor U2961 (N_2961,N_2424,N_2287);
nor U2962 (N_2962,N_2440,N_2026);
nand U2963 (N_2963,N_2403,N_2487);
or U2964 (N_2964,N_2219,N_2410);
nor U2965 (N_2965,N_2169,N_2261);
nand U2966 (N_2966,N_2088,N_2328);
nor U2967 (N_2967,N_2432,N_2397);
nand U2968 (N_2968,N_2343,N_2028);
and U2969 (N_2969,N_2002,N_2372);
nand U2970 (N_2970,N_2426,N_2265);
or U2971 (N_2971,N_2366,N_2385);
or U2972 (N_2972,N_2372,N_2156);
or U2973 (N_2973,N_2042,N_2240);
and U2974 (N_2974,N_2340,N_2292);
nand U2975 (N_2975,N_2289,N_2358);
nor U2976 (N_2976,N_2258,N_2318);
or U2977 (N_2977,N_2363,N_2270);
or U2978 (N_2978,N_2268,N_2447);
and U2979 (N_2979,N_2387,N_2467);
and U2980 (N_2980,N_2162,N_2201);
xor U2981 (N_2981,N_2476,N_2339);
and U2982 (N_2982,N_2241,N_2025);
nor U2983 (N_2983,N_2194,N_2328);
and U2984 (N_2984,N_2355,N_2479);
nand U2985 (N_2985,N_2455,N_2304);
or U2986 (N_2986,N_2308,N_2489);
and U2987 (N_2987,N_2418,N_2488);
and U2988 (N_2988,N_2171,N_2290);
and U2989 (N_2989,N_2245,N_2045);
nor U2990 (N_2990,N_2445,N_2132);
or U2991 (N_2991,N_2159,N_2317);
or U2992 (N_2992,N_2470,N_2056);
or U2993 (N_2993,N_2051,N_2005);
xnor U2994 (N_2994,N_2341,N_2003);
or U2995 (N_2995,N_2064,N_2100);
nand U2996 (N_2996,N_2276,N_2054);
and U2997 (N_2997,N_2332,N_2475);
or U2998 (N_2998,N_2160,N_2272);
nor U2999 (N_2999,N_2366,N_2365);
or UO_0 (O_0,N_2891,N_2669);
nand UO_1 (O_1,N_2503,N_2772);
or UO_2 (O_2,N_2856,N_2925);
nand UO_3 (O_3,N_2823,N_2853);
nand UO_4 (O_4,N_2639,N_2935);
and UO_5 (O_5,N_2657,N_2865);
and UO_6 (O_6,N_2918,N_2501);
and UO_7 (O_7,N_2697,N_2919);
and UO_8 (O_8,N_2912,N_2846);
and UO_9 (O_9,N_2554,N_2628);
and UO_10 (O_10,N_2577,N_2949);
nand UO_11 (O_11,N_2871,N_2708);
nand UO_12 (O_12,N_2933,N_2505);
and UO_13 (O_13,N_2551,N_2597);
nand UO_14 (O_14,N_2567,N_2666);
or UO_15 (O_15,N_2979,N_2981);
and UO_16 (O_16,N_2841,N_2616);
and UO_17 (O_17,N_2924,N_2637);
nor UO_18 (O_18,N_2952,N_2508);
or UO_19 (O_19,N_2517,N_2582);
nand UO_20 (O_20,N_2620,N_2768);
or UO_21 (O_21,N_2928,N_2660);
nor UO_22 (O_22,N_2513,N_2754);
nor UO_23 (O_23,N_2834,N_2529);
or UO_24 (O_24,N_2855,N_2808);
nand UO_25 (O_25,N_2920,N_2926);
and UO_26 (O_26,N_2690,N_2795);
nor UO_27 (O_27,N_2654,N_2804);
or UO_28 (O_28,N_2817,N_2715);
nand UO_29 (O_29,N_2632,N_2990);
nand UO_30 (O_30,N_2993,N_2664);
or UO_31 (O_31,N_2889,N_2614);
nand UO_32 (O_32,N_2872,N_2782);
and UO_33 (O_33,N_2904,N_2914);
and UO_34 (O_34,N_2803,N_2605);
nor UO_35 (O_35,N_2759,N_2913);
and UO_36 (O_36,N_2923,N_2946);
nor UO_37 (O_37,N_2948,N_2543);
nand UO_38 (O_38,N_2764,N_2672);
nand UO_39 (O_39,N_2676,N_2552);
nand UO_40 (O_40,N_2835,N_2570);
nand UO_41 (O_41,N_2504,N_2910);
nand UO_42 (O_42,N_2659,N_2929);
nor UO_43 (O_43,N_2864,N_2774);
nor UO_44 (O_44,N_2721,N_2623);
nand UO_45 (O_45,N_2731,N_2518);
or UO_46 (O_46,N_2645,N_2566);
nand UO_47 (O_47,N_2944,N_2862);
nand UO_48 (O_48,N_2511,N_2894);
nor UO_49 (O_49,N_2514,N_2562);
nand UO_50 (O_50,N_2932,N_2820);
nor UO_51 (O_51,N_2942,N_2585);
or UO_52 (O_52,N_2601,N_2879);
or UO_53 (O_53,N_2773,N_2814);
nand UO_54 (O_54,N_2793,N_2712);
nor UO_55 (O_55,N_2502,N_2594);
and UO_56 (O_56,N_2674,N_2553);
and UO_57 (O_57,N_2578,N_2580);
nand UO_58 (O_58,N_2825,N_2983);
nor UO_59 (O_59,N_2828,N_2705);
or UO_60 (O_60,N_2618,N_2515);
or UO_61 (O_61,N_2767,N_2533);
nor UO_62 (O_62,N_2652,N_2550);
or UO_63 (O_63,N_2987,N_2701);
and UO_64 (O_64,N_2982,N_2727);
nand UO_65 (O_65,N_2742,N_2922);
nor UO_66 (O_66,N_2573,N_2905);
and UO_67 (O_67,N_2936,N_2863);
xor UO_68 (O_68,N_2854,N_2678);
xor UO_69 (O_69,N_2583,N_2723);
nand UO_70 (O_70,N_2592,N_2916);
nor UO_71 (O_71,N_2525,N_2794);
nor UO_72 (O_72,N_2538,N_2873);
nor UO_73 (O_73,N_2574,N_2930);
or UO_74 (O_74,N_2500,N_2753);
xor UO_75 (O_75,N_2867,N_2702);
nand UO_76 (O_76,N_2693,N_2746);
or UO_77 (O_77,N_2670,N_2845);
and UO_78 (O_78,N_2745,N_2899);
or UO_79 (O_79,N_2810,N_2530);
nand UO_80 (O_80,N_2756,N_2851);
or UO_81 (O_81,N_2575,N_2945);
nor UO_82 (O_82,N_2978,N_2868);
nor UO_83 (O_83,N_2897,N_2760);
and UO_84 (O_84,N_2941,N_2587);
or UO_85 (O_85,N_2939,N_2622);
nand UO_86 (O_86,N_2586,N_2655);
xor UO_87 (O_87,N_2943,N_2569);
or UO_88 (O_88,N_2765,N_2895);
nand UO_89 (O_89,N_2734,N_2624);
and UO_90 (O_90,N_2732,N_2581);
nand UO_91 (O_91,N_2847,N_2984);
nor UO_92 (O_92,N_2850,N_2758);
nor UO_93 (O_93,N_2947,N_2726);
and UO_94 (O_94,N_2736,N_2679);
and UO_95 (O_95,N_2537,N_2681);
nand UO_96 (O_96,N_2821,N_2805);
nand UO_97 (O_97,N_2859,N_2596);
and UO_98 (O_98,N_2740,N_2520);
or UO_99 (O_99,N_2829,N_2707);
or UO_100 (O_100,N_2516,N_2642);
and UO_101 (O_101,N_2792,N_2519);
and UO_102 (O_102,N_2507,N_2974);
nand UO_103 (O_103,N_2668,N_2547);
xnor UO_104 (O_104,N_2940,N_2600);
nor UO_105 (O_105,N_2752,N_2838);
nor UO_106 (O_106,N_2630,N_2634);
and UO_107 (O_107,N_2836,N_2966);
and UO_108 (O_108,N_2991,N_2662);
and UO_109 (O_109,N_2650,N_2741);
nor UO_110 (O_110,N_2606,N_2813);
nand UO_111 (O_111,N_2776,N_2555);
nand UO_112 (O_112,N_2536,N_2961);
nand UO_113 (O_113,N_2761,N_2667);
xnor UO_114 (O_114,N_2878,N_2688);
and UO_115 (O_115,N_2684,N_2921);
nor UO_116 (O_116,N_2743,N_2785);
and UO_117 (O_117,N_2779,N_2653);
or UO_118 (O_118,N_2692,N_2787);
nand UO_119 (O_119,N_2700,N_2778);
and UO_120 (O_120,N_2711,N_2901);
nand UO_121 (O_121,N_2874,N_2967);
or UO_122 (O_122,N_2777,N_2870);
and UO_123 (O_123,N_2506,N_2512);
nand UO_124 (O_124,N_2848,N_2802);
or UO_125 (O_125,N_2527,N_2571);
nand UO_126 (O_126,N_2563,N_2877);
xnor UO_127 (O_127,N_2903,N_2717);
or UO_128 (O_128,N_2747,N_2739);
nor UO_129 (O_129,N_2771,N_2539);
and UO_130 (O_130,N_2975,N_2576);
nor UO_131 (O_131,N_2833,N_2584);
nand UO_132 (O_132,N_2781,N_2720);
nand UO_133 (O_133,N_2883,N_2589);
nand UO_134 (O_134,N_2950,N_2718);
nor UO_135 (O_135,N_2695,N_2648);
nand UO_136 (O_136,N_2959,N_2911);
and UO_137 (O_137,N_2775,N_2909);
and UO_138 (O_138,N_2748,N_2619);
or UO_139 (O_139,N_2977,N_2938);
nand UO_140 (O_140,N_2880,N_2963);
nor UO_141 (O_141,N_2900,N_2931);
nor UO_142 (O_142,N_2699,N_2524);
nor UO_143 (O_143,N_2615,N_2541);
or UO_144 (O_144,N_2893,N_2633);
or UO_145 (O_145,N_2881,N_2969);
nor UO_146 (O_146,N_2790,N_2783);
nor UO_147 (O_147,N_2647,N_2682);
or UO_148 (O_148,N_2651,N_2696);
and UO_149 (O_149,N_2858,N_2561);
nand UO_150 (O_150,N_2857,N_2534);
and UO_151 (O_151,N_2824,N_2994);
nor UO_152 (O_152,N_2876,N_2509);
or UO_153 (O_153,N_2598,N_2751);
or UO_154 (O_154,N_2789,N_2557);
xor UO_155 (O_155,N_2641,N_2980);
nor UO_156 (O_156,N_2698,N_2714);
and UO_157 (O_157,N_2907,N_2556);
nor UO_158 (O_158,N_2716,N_2780);
or UO_159 (O_159,N_2593,N_2843);
nand UO_160 (O_160,N_2730,N_2646);
nand UO_161 (O_161,N_2750,N_2784);
or UO_162 (O_162,N_2869,N_2663);
nand UO_163 (O_163,N_2788,N_2704);
and UO_164 (O_164,N_2523,N_2591);
and UO_165 (O_165,N_2687,N_2812);
and UO_166 (O_166,N_2713,N_2999);
nor UO_167 (O_167,N_2542,N_2724);
nor UO_168 (O_168,N_2613,N_2840);
and UO_169 (O_169,N_2837,N_2989);
xor UO_170 (O_170,N_2629,N_2861);
or UO_171 (O_171,N_2689,N_2860);
and UO_172 (O_172,N_2522,N_2995);
or UO_173 (O_173,N_2649,N_2827);
or UO_174 (O_174,N_2839,N_2766);
or UO_175 (O_175,N_2602,N_2565);
nor UO_176 (O_176,N_2954,N_2965);
nor UO_177 (O_177,N_2611,N_2559);
nor UO_178 (O_178,N_2971,N_2510);
nor UO_179 (O_179,N_2703,N_2934);
or UO_180 (O_180,N_2535,N_2960);
or UO_181 (O_181,N_2807,N_2882);
nand UO_182 (O_182,N_2770,N_2769);
or UO_183 (O_183,N_2819,N_2590);
and UO_184 (O_184,N_2737,N_2560);
xor UO_185 (O_185,N_2733,N_2626);
xor UO_186 (O_186,N_2545,N_2709);
xnor UO_187 (O_187,N_2548,N_2744);
or UO_188 (O_188,N_2675,N_2603);
nand UO_189 (O_189,N_2830,N_2607);
nor UO_190 (O_190,N_2927,N_2612);
and UO_191 (O_191,N_2621,N_2985);
and UO_192 (O_192,N_2604,N_2627);
nand UO_193 (O_193,N_2722,N_2844);
and UO_194 (O_194,N_2806,N_2656);
or UO_195 (O_195,N_2735,N_2998);
nor UO_196 (O_196,N_2885,N_2568);
and UO_197 (O_197,N_2908,N_2917);
nor UO_198 (O_198,N_2818,N_2617);
nor UO_199 (O_199,N_2797,N_2992);
nand UO_200 (O_200,N_2738,N_2786);
xor UO_201 (O_201,N_2884,N_2898);
nor UO_202 (O_202,N_2997,N_2609);
nor UO_203 (O_203,N_2686,N_2671);
or UO_204 (O_204,N_2588,N_2638);
nor UO_205 (O_205,N_2896,N_2799);
or UO_206 (O_206,N_2968,N_2953);
or UO_207 (O_207,N_2729,N_2986);
nor UO_208 (O_208,N_2532,N_2832);
nand UO_209 (O_209,N_2852,N_2892);
and UO_210 (O_210,N_2831,N_2719);
and UO_211 (O_211,N_2757,N_2599);
or UO_212 (O_212,N_2544,N_2866);
nor UO_213 (O_213,N_2643,N_2680);
nor UO_214 (O_214,N_2610,N_2763);
or UO_215 (O_215,N_2755,N_2800);
and UO_216 (O_216,N_2677,N_2890);
or UO_217 (O_217,N_2826,N_2887);
and UO_218 (O_218,N_2996,N_2528);
nor UO_219 (O_219,N_2673,N_2875);
xnor UO_220 (O_220,N_2956,N_2970);
nand UO_221 (O_221,N_2796,N_2962);
nand UO_222 (O_222,N_2915,N_2976);
nor UO_223 (O_223,N_2640,N_2725);
xnor UO_224 (O_224,N_2951,N_2636);
and UO_225 (O_225,N_2749,N_2955);
nor UO_226 (O_226,N_2728,N_2809);
nand UO_227 (O_227,N_2815,N_2710);
or UO_228 (O_228,N_2762,N_2540);
nand UO_229 (O_229,N_2625,N_2683);
nand UO_230 (O_230,N_2631,N_2888);
or UO_231 (O_231,N_2958,N_2849);
xnor UO_232 (O_232,N_2665,N_2801);
and UO_233 (O_233,N_2886,N_2579);
and UO_234 (O_234,N_2546,N_2572);
and UO_235 (O_235,N_2791,N_2558);
or UO_236 (O_236,N_2521,N_2564);
nor UO_237 (O_237,N_2658,N_2906);
xnor UO_238 (O_238,N_2691,N_2595);
nor UO_239 (O_239,N_2644,N_2811);
nor UO_240 (O_240,N_2988,N_2608);
or UO_241 (O_241,N_2902,N_2635);
or UO_242 (O_242,N_2549,N_2685);
or UO_243 (O_243,N_2816,N_2822);
or UO_244 (O_244,N_2694,N_2526);
or UO_245 (O_245,N_2973,N_2531);
nor UO_246 (O_246,N_2706,N_2972);
nor UO_247 (O_247,N_2842,N_2937);
and UO_248 (O_248,N_2964,N_2661);
xor UO_249 (O_249,N_2798,N_2957);
nand UO_250 (O_250,N_2648,N_2508);
nand UO_251 (O_251,N_2590,N_2897);
and UO_252 (O_252,N_2832,N_2786);
or UO_253 (O_253,N_2579,N_2530);
nand UO_254 (O_254,N_2610,N_2801);
nand UO_255 (O_255,N_2869,N_2659);
or UO_256 (O_256,N_2503,N_2872);
xnor UO_257 (O_257,N_2706,N_2584);
and UO_258 (O_258,N_2941,N_2627);
or UO_259 (O_259,N_2532,N_2779);
or UO_260 (O_260,N_2962,N_2968);
nor UO_261 (O_261,N_2803,N_2691);
nor UO_262 (O_262,N_2768,N_2735);
or UO_263 (O_263,N_2673,N_2766);
nand UO_264 (O_264,N_2736,N_2535);
nand UO_265 (O_265,N_2648,N_2520);
or UO_266 (O_266,N_2988,N_2654);
nor UO_267 (O_267,N_2864,N_2638);
nand UO_268 (O_268,N_2562,N_2808);
or UO_269 (O_269,N_2567,N_2704);
nand UO_270 (O_270,N_2782,N_2589);
nor UO_271 (O_271,N_2518,N_2632);
and UO_272 (O_272,N_2755,N_2896);
or UO_273 (O_273,N_2742,N_2635);
or UO_274 (O_274,N_2865,N_2569);
or UO_275 (O_275,N_2745,N_2739);
or UO_276 (O_276,N_2699,N_2893);
nand UO_277 (O_277,N_2527,N_2656);
xnor UO_278 (O_278,N_2626,N_2753);
nand UO_279 (O_279,N_2952,N_2996);
and UO_280 (O_280,N_2910,N_2840);
nand UO_281 (O_281,N_2817,N_2881);
xor UO_282 (O_282,N_2621,N_2710);
xnor UO_283 (O_283,N_2603,N_2998);
nor UO_284 (O_284,N_2504,N_2854);
nor UO_285 (O_285,N_2856,N_2523);
and UO_286 (O_286,N_2922,N_2510);
nand UO_287 (O_287,N_2676,N_2519);
nand UO_288 (O_288,N_2529,N_2672);
nor UO_289 (O_289,N_2534,N_2564);
and UO_290 (O_290,N_2695,N_2575);
or UO_291 (O_291,N_2545,N_2663);
or UO_292 (O_292,N_2582,N_2719);
nor UO_293 (O_293,N_2912,N_2820);
nand UO_294 (O_294,N_2982,N_2935);
or UO_295 (O_295,N_2811,N_2979);
nand UO_296 (O_296,N_2704,N_2650);
or UO_297 (O_297,N_2982,N_2527);
nand UO_298 (O_298,N_2540,N_2621);
nand UO_299 (O_299,N_2621,N_2973);
nand UO_300 (O_300,N_2945,N_2804);
nand UO_301 (O_301,N_2911,N_2790);
nor UO_302 (O_302,N_2969,N_2680);
or UO_303 (O_303,N_2560,N_2618);
and UO_304 (O_304,N_2794,N_2933);
nand UO_305 (O_305,N_2893,N_2874);
and UO_306 (O_306,N_2689,N_2755);
xor UO_307 (O_307,N_2501,N_2897);
or UO_308 (O_308,N_2986,N_2645);
nor UO_309 (O_309,N_2870,N_2917);
nand UO_310 (O_310,N_2894,N_2936);
or UO_311 (O_311,N_2632,N_2757);
xnor UO_312 (O_312,N_2512,N_2763);
nor UO_313 (O_313,N_2709,N_2651);
nor UO_314 (O_314,N_2875,N_2723);
nand UO_315 (O_315,N_2861,N_2551);
or UO_316 (O_316,N_2917,N_2705);
and UO_317 (O_317,N_2665,N_2817);
nor UO_318 (O_318,N_2932,N_2578);
nand UO_319 (O_319,N_2979,N_2730);
nand UO_320 (O_320,N_2832,N_2610);
nor UO_321 (O_321,N_2568,N_2817);
or UO_322 (O_322,N_2705,N_2631);
or UO_323 (O_323,N_2972,N_2989);
or UO_324 (O_324,N_2882,N_2938);
or UO_325 (O_325,N_2821,N_2681);
nor UO_326 (O_326,N_2625,N_2920);
nor UO_327 (O_327,N_2910,N_2828);
or UO_328 (O_328,N_2598,N_2587);
nor UO_329 (O_329,N_2521,N_2666);
xnor UO_330 (O_330,N_2734,N_2928);
nand UO_331 (O_331,N_2541,N_2703);
or UO_332 (O_332,N_2790,N_2885);
and UO_333 (O_333,N_2847,N_2852);
nor UO_334 (O_334,N_2710,N_2930);
nor UO_335 (O_335,N_2751,N_2971);
nand UO_336 (O_336,N_2501,N_2514);
nor UO_337 (O_337,N_2609,N_2644);
nand UO_338 (O_338,N_2514,N_2737);
or UO_339 (O_339,N_2613,N_2890);
nand UO_340 (O_340,N_2741,N_2958);
xnor UO_341 (O_341,N_2901,N_2967);
and UO_342 (O_342,N_2873,N_2976);
and UO_343 (O_343,N_2848,N_2775);
and UO_344 (O_344,N_2511,N_2663);
or UO_345 (O_345,N_2933,N_2911);
nor UO_346 (O_346,N_2500,N_2501);
nor UO_347 (O_347,N_2503,N_2943);
nor UO_348 (O_348,N_2646,N_2839);
and UO_349 (O_349,N_2999,N_2851);
nor UO_350 (O_350,N_2922,N_2638);
and UO_351 (O_351,N_2583,N_2852);
nor UO_352 (O_352,N_2748,N_2849);
nand UO_353 (O_353,N_2994,N_2512);
xnor UO_354 (O_354,N_2982,N_2876);
nand UO_355 (O_355,N_2732,N_2628);
xnor UO_356 (O_356,N_2658,N_2699);
xor UO_357 (O_357,N_2833,N_2527);
nor UO_358 (O_358,N_2534,N_2854);
and UO_359 (O_359,N_2580,N_2943);
nand UO_360 (O_360,N_2795,N_2661);
nor UO_361 (O_361,N_2810,N_2662);
nand UO_362 (O_362,N_2736,N_2558);
nor UO_363 (O_363,N_2825,N_2950);
xor UO_364 (O_364,N_2680,N_2754);
or UO_365 (O_365,N_2686,N_2635);
nand UO_366 (O_366,N_2854,N_2677);
or UO_367 (O_367,N_2959,N_2723);
and UO_368 (O_368,N_2812,N_2645);
nand UO_369 (O_369,N_2806,N_2515);
xor UO_370 (O_370,N_2792,N_2970);
nor UO_371 (O_371,N_2949,N_2715);
xnor UO_372 (O_372,N_2804,N_2573);
and UO_373 (O_373,N_2908,N_2767);
nand UO_374 (O_374,N_2991,N_2811);
and UO_375 (O_375,N_2533,N_2911);
or UO_376 (O_376,N_2597,N_2811);
nand UO_377 (O_377,N_2888,N_2575);
and UO_378 (O_378,N_2760,N_2646);
and UO_379 (O_379,N_2710,N_2970);
nor UO_380 (O_380,N_2608,N_2545);
or UO_381 (O_381,N_2818,N_2804);
xnor UO_382 (O_382,N_2937,N_2871);
and UO_383 (O_383,N_2632,N_2861);
xor UO_384 (O_384,N_2631,N_2763);
nand UO_385 (O_385,N_2734,N_2504);
or UO_386 (O_386,N_2960,N_2784);
nor UO_387 (O_387,N_2771,N_2651);
nor UO_388 (O_388,N_2864,N_2812);
nor UO_389 (O_389,N_2880,N_2647);
nor UO_390 (O_390,N_2506,N_2707);
and UO_391 (O_391,N_2902,N_2615);
or UO_392 (O_392,N_2816,N_2945);
nor UO_393 (O_393,N_2961,N_2582);
nor UO_394 (O_394,N_2601,N_2553);
nand UO_395 (O_395,N_2595,N_2534);
and UO_396 (O_396,N_2875,N_2976);
nand UO_397 (O_397,N_2855,N_2520);
nor UO_398 (O_398,N_2618,N_2947);
nor UO_399 (O_399,N_2655,N_2709);
or UO_400 (O_400,N_2809,N_2993);
and UO_401 (O_401,N_2852,N_2760);
and UO_402 (O_402,N_2651,N_2853);
nor UO_403 (O_403,N_2627,N_2730);
xnor UO_404 (O_404,N_2532,N_2986);
or UO_405 (O_405,N_2668,N_2726);
or UO_406 (O_406,N_2997,N_2922);
nor UO_407 (O_407,N_2996,N_2634);
nor UO_408 (O_408,N_2518,N_2502);
or UO_409 (O_409,N_2928,N_2763);
and UO_410 (O_410,N_2526,N_2763);
nand UO_411 (O_411,N_2671,N_2814);
nand UO_412 (O_412,N_2732,N_2688);
nand UO_413 (O_413,N_2680,N_2668);
nor UO_414 (O_414,N_2822,N_2551);
and UO_415 (O_415,N_2546,N_2788);
nor UO_416 (O_416,N_2545,N_2778);
and UO_417 (O_417,N_2788,N_2685);
xor UO_418 (O_418,N_2894,N_2786);
and UO_419 (O_419,N_2600,N_2868);
and UO_420 (O_420,N_2637,N_2583);
and UO_421 (O_421,N_2976,N_2679);
and UO_422 (O_422,N_2520,N_2847);
nor UO_423 (O_423,N_2736,N_2775);
xnor UO_424 (O_424,N_2803,N_2616);
nor UO_425 (O_425,N_2939,N_2575);
nand UO_426 (O_426,N_2674,N_2899);
nand UO_427 (O_427,N_2567,N_2565);
nor UO_428 (O_428,N_2948,N_2681);
nor UO_429 (O_429,N_2954,N_2755);
nand UO_430 (O_430,N_2961,N_2677);
and UO_431 (O_431,N_2722,N_2995);
xnor UO_432 (O_432,N_2885,N_2800);
nand UO_433 (O_433,N_2584,N_2807);
or UO_434 (O_434,N_2909,N_2768);
nand UO_435 (O_435,N_2651,N_2560);
or UO_436 (O_436,N_2550,N_2784);
nor UO_437 (O_437,N_2922,N_2728);
nor UO_438 (O_438,N_2646,N_2999);
nor UO_439 (O_439,N_2564,N_2648);
nor UO_440 (O_440,N_2588,N_2789);
nand UO_441 (O_441,N_2980,N_2820);
and UO_442 (O_442,N_2788,N_2859);
nand UO_443 (O_443,N_2579,N_2937);
nor UO_444 (O_444,N_2892,N_2734);
nand UO_445 (O_445,N_2578,N_2631);
or UO_446 (O_446,N_2527,N_2645);
or UO_447 (O_447,N_2721,N_2764);
xor UO_448 (O_448,N_2884,N_2593);
nand UO_449 (O_449,N_2816,N_2594);
nor UO_450 (O_450,N_2677,N_2761);
nor UO_451 (O_451,N_2508,N_2821);
xor UO_452 (O_452,N_2553,N_2903);
and UO_453 (O_453,N_2974,N_2988);
or UO_454 (O_454,N_2702,N_2969);
or UO_455 (O_455,N_2894,N_2647);
and UO_456 (O_456,N_2724,N_2784);
nor UO_457 (O_457,N_2813,N_2944);
nand UO_458 (O_458,N_2675,N_2870);
nand UO_459 (O_459,N_2832,N_2920);
or UO_460 (O_460,N_2812,N_2851);
nor UO_461 (O_461,N_2607,N_2753);
or UO_462 (O_462,N_2875,N_2755);
or UO_463 (O_463,N_2826,N_2928);
and UO_464 (O_464,N_2711,N_2746);
or UO_465 (O_465,N_2804,N_2781);
nor UO_466 (O_466,N_2790,N_2592);
or UO_467 (O_467,N_2652,N_2635);
nor UO_468 (O_468,N_2974,N_2625);
or UO_469 (O_469,N_2715,N_2672);
or UO_470 (O_470,N_2770,N_2994);
nor UO_471 (O_471,N_2658,N_2563);
nand UO_472 (O_472,N_2882,N_2744);
or UO_473 (O_473,N_2542,N_2889);
xnor UO_474 (O_474,N_2648,N_2888);
nor UO_475 (O_475,N_2917,N_2702);
or UO_476 (O_476,N_2910,N_2608);
and UO_477 (O_477,N_2898,N_2946);
and UO_478 (O_478,N_2695,N_2869);
and UO_479 (O_479,N_2787,N_2793);
or UO_480 (O_480,N_2510,N_2683);
or UO_481 (O_481,N_2815,N_2980);
or UO_482 (O_482,N_2686,N_2539);
xnor UO_483 (O_483,N_2670,N_2956);
xor UO_484 (O_484,N_2900,N_2841);
nor UO_485 (O_485,N_2801,N_2536);
nor UO_486 (O_486,N_2903,N_2693);
nor UO_487 (O_487,N_2711,N_2958);
xor UO_488 (O_488,N_2932,N_2583);
or UO_489 (O_489,N_2931,N_2974);
and UO_490 (O_490,N_2922,N_2932);
or UO_491 (O_491,N_2565,N_2912);
and UO_492 (O_492,N_2542,N_2779);
and UO_493 (O_493,N_2952,N_2809);
and UO_494 (O_494,N_2975,N_2672);
nand UO_495 (O_495,N_2695,N_2522);
and UO_496 (O_496,N_2975,N_2649);
and UO_497 (O_497,N_2505,N_2899);
or UO_498 (O_498,N_2551,N_2855);
nand UO_499 (O_499,N_2577,N_2880);
endmodule