module basic_1500_15000_2000_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_843,In_1389);
or U1 (N_1,In_66,In_513);
xnor U2 (N_2,In_914,In_262);
nand U3 (N_3,In_952,In_304);
xnor U4 (N_4,In_1145,In_1489);
xor U5 (N_5,In_554,In_283);
and U6 (N_6,In_49,In_422);
nor U7 (N_7,In_617,In_606);
xnor U8 (N_8,In_217,In_3);
nor U9 (N_9,In_1157,In_418);
nor U10 (N_10,In_867,In_499);
nor U11 (N_11,In_726,In_1116);
nor U12 (N_12,In_447,In_662);
or U13 (N_13,In_641,In_430);
xor U14 (N_14,In_980,In_1235);
nand U15 (N_15,In_1233,In_132);
and U16 (N_16,In_1449,In_1068);
nor U17 (N_17,In_1009,In_734);
or U18 (N_18,In_74,In_586);
xor U19 (N_19,In_460,In_114);
nor U20 (N_20,In_77,In_524);
or U21 (N_21,In_1448,In_1273);
and U22 (N_22,In_1276,In_280);
or U23 (N_23,In_152,In_674);
xnor U24 (N_24,In_932,In_511);
or U25 (N_25,In_935,In_317);
or U26 (N_26,In_992,In_667);
and U27 (N_27,In_311,In_895);
xnor U28 (N_28,In_1360,In_465);
nor U29 (N_29,In_1099,In_1209);
nor U30 (N_30,In_1158,In_119);
xnor U31 (N_31,In_1049,In_1117);
nand U32 (N_32,In_1460,In_1071);
or U33 (N_33,In_1372,In_94);
nand U34 (N_34,In_1057,In_1179);
or U35 (N_35,In_487,In_368);
nor U36 (N_36,In_1282,In_1459);
nor U37 (N_37,In_602,In_695);
nor U38 (N_38,In_815,In_358);
xor U39 (N_39,In_302,In_1180);
xnor U40 (N_40,In_1348,In_1087);
or U41 (N_41,In_782,In_906);
and U42 (N_42,In_321,In_716);
nand U43 (N_43,In_1487,In_637);
nand U44 (N_44,In_970,In_400);
nor U45 (N_45,In_593,In_338);
nand U46 (N_46,In_16,In_922);
nor U47 (N_47,In_854,In_37);
xor U48 (N_48,In_1485,In_1030);
xor U49 (N_49,In_620,In_207);
and U50 (N_50,In_616,In_1012);
or U51 (N_51,In_1352,In_708);
or U52 (N_52,In_439,In_290);
nor U53 (N_53,In_610,In_937);
or U54 (N_54,In_296,In_1318);
and U55 (N_55,In_174,In_976);
nand U56 (N_56,In_975,In_1440);
nor U57 (N_57,In_799,In_911);
or U58 (N_58,In_113,In_1369);
and U59 (N_59,In_256,In_828);
and U60 (N_60,In_1398,In_1134);
or U61 (N_61,In_1194,In_719);
xnor U62 (N_62,In_44,In_2);
nor U63 (N_63,In_746,In_688);
and U64 (N_64,In_489,In_1256);
nor U65 (N_65,In_864,In_1047);
xnor U66 (N_66,In_785,In_1111);
or U67 (N_67,In_608,In_502);
xnor U68 (N_68,In_90,In_60);
xor U69 (N_69,In_219,In_443);
nand U70 (N_70,In_1102,In_1085);
xor U71 (N_71,In_1106,In_107);
or U72 (N_72,In_1455,In_731);
xor U73 (N_73,In_23,In_160);
nor U74 (N_74,In_1472,In_1008);
xnor U75 (N_75,In_1045,In_446);
nor U76 (N_76,In_196,In_176);
and U77 (N_77,In_229,In_1149);
nand U78 (N_78,In_1065,In_1141);
nor U79 (N_79,In_794,In_310);
nor U80 (N_80,In_102,In_93);
nor U81 (N_81,In_798,In_936);
xnor U82 (N_82,In_1488,In_1379);
or U83 (N_83,In_8,In_562);
and U84 (N_84,In_53,In_215);
and U85 (N_85,In_1078,In_241);
nor U86 (N_86,In_1481,In_1224);
nor U87 (N_87,In_352,In_238);
nand U88 (N_88,In_1468,In_636);
xor U89 (N_89,In_792,In_747);
nor U90 (N_90,In_1197,In_1254);
xnor U91 (N_91,In_1132,In_36);
xnor U92 (N_92,In_1280,In_1413);
nand U93 (N_93,In_530,In_182);
xnor U94 (N_94,In_1129,In_823);
or U95 (N_95,In_694,In_12);
nand U96 (N_96,In_703,In_1174);
xor U97 (N_97,In_301,In_812);
nor U98 (N_98,In_783,In_1173);
xnor U99 (N_99,In_300,In_224);
nor U100 (N_100,In_879,In_62);
nor U101 (N_101,In_998,In_904);
or U102 (N_102,In_1059,In_1013);
xnor U103 (N_103,In_1015,In_1275);
and U104 (N_104,In_1362,In_813);
or U105 (N_105,In_950,In_1407);
nor U106 (N_106,In_425,In_983);
xnor U107 (N_107,In_947,In_1090);
and U108 (N_108,In_409,In_924);
nor U109 (N_109,In_1014,In_190);
nor U110 (N_110,In_1063,In_1107);
nor U111 (N_111,In_1255,In_779);
or U112 (N_112,In_379,In_270);
and U113 (N_113,In_827,In_1269);
xor U114 (N_114,In_1246,In_591);
and U115 (N_115,In_1385,In_381);
and U116 (N_116,In_434,In_816);
nor U117 (N_117,In_202,In_1412);
nor U118 (N_118,In_145,In_265);
nor U119 (N_119,In_717,In_367);
xnor U120 (N_120,In_35,In_137);
or U121 (N_121,In_462,In_665);
and U122 (N_122,In_917,In_449);
or U123 (N_123,In_455,In_578);
nand U124 (N_124,In_13,In_1387);
and U125 (N_125,In_1365,In_656);
and U126 (N_126,In_1397,In_1312);
or U127 (N_127,In_220,In_40);
nand U128 (N_128,In_755,In_941);
xor U129 (N_129,In_161,In_1354);
and U130 (N_130,In_691,In_912);
and U131 (N_131,In_255,In_32);
or U132 (N_132,In_250,In_68);
and U133 (N_133,In_353,In_108);
or U134 (N_134,In_1370,In_309);
nand U135 (N_135,In_336,In_715);
or U136 (N_136,In_705,In_390);
or U137 (N_137,In_488,In_1230);
nor U138 (N_138,In_450,In_401);
or U139 (N_139,In_659,In_239);
xor U140 (N_140,In_1147,In_738);
nand U141 (N_141,In_866,In_825);
xor U142 (N_142,In_1183,In_550);
and U143 (N_143,In_273,In_557);
or U144 (N_144,In_635,In_166);
xor U145 (N_145,In_1093,In_1004);
and U146 (N_146,In_1108,In_902);
xor U147 (N_147,In_672,In_123);
and U148 (N_148,In_954,In_526);
and U149 (N_149,In_706,In_1429);
nand U150 (N_150,In_320,In_6);
nand U151 (N_151,In_1154,In_42);
xnor U152 (N_152,In_218,In_873);
nor U153 (N_153,In_351,In_582);
xnor U154 (N_154,In_382,In_870);
nand U155 (N_155,In_1120,In_246);
xor U156 (N_156,In_39,In_1044);
and U157 (N_157,In_673,In_851);
or U158 (N_158,In_216,In_1214);
xor U159 (N_159,In_185,In_201);
nand U160 (N_160,In_1084,In_677);
xnor U161 (N_161,In_426,In_574);
and U162 (N_162,In_1279,In_329);
nor U163 (N_163,In_1374,In_745);
and U164 (N_164,In_743,In_288);
nor U165 (N_165,In_589,In_1346);
and U166 (N_166,In_516,In_881);
xor U167 (N_167,In_527,In_496);
and U168 (N_168,In_1188,In_803);
nor U169 (N_169,In_1446,In_1064);
and U170 (N_170,In_1094,In_1458);
xor U171 (N_171,In_634,In_159);
or U172 (N_172,In_1396,In_433);
xor U173 (N_173,In_188,In_1143);
xor U174 (N_174,In_1278,In_1035);
xnor U175 (N_175,In_929,In_1327);
xnor U176 (N_176,In_1416,In_1046);
nor U177 (N_177,In_1293,In_212);
nor U178 (N_178,In_1190,In_438);
nand U179 (N_179,In_1479,In_233);
and U180 (N_180,In_981,In_21);
nand U181 (N_181,In_1220,In_445);
xor U182 (N_182,In_1038,In_1142);
or U183 (N_183,In_164,In_1097);
nand U184 (N_184,In_1131,In_323);
nand U185 (N_185,In_31,In_46);
xor U186 (N_186,In_1028,In_626);
or U187 (N_187,In_555,In_1210);
or U188 (N_188,In_649,In_1140);
xor U189 (N_189,In_1155,In_109);
or U190 (N_190,In_393,In_821);
or U191 (N_191,In_862,In_966);
nor U192 (N_192,In_1123,In_1218);
and U193 (N_193,In_824,In_135);
nor U194 (N_194,In_331,In_1466);
or U195 (N_195,In_1480,In_1029);
xnor U196 (N_196,In_529,In_1283);
nor U197 (N_197,In_597,In_1494);
nor U198 (N_198,In_934,In_964);
nand U199 (N_199,In_236,In_1050);
nand U200 (N_200,In_1041,In_886);
and U201 (N_201,In_14,In_1442);
nor U202 (N_202,In_538,In_1286);
and U203 (N_203,In_279,In_880);
and U204 (N_204,In_507,In_153);
nand U205 (N_205,In_1005,In_22);
and U206 (N_206,In_1320,In_274);
or U207 (N_207,In_1053,In_1338);
or U208 (N_208,In_208,In_1033);
nand U209 (N_209,In_410,In_1323);
xor U210 (N_210,In_809,In_1020);
and U211 (N_211,In_149,In_454);
and U212 (N_212,In_1062,In_1016);
and U213 (N_213,In_729,In_25);
nand U214 (N_214,In_24,In_305);
and U215 (N_215,In_429,In_903);
and U216 (N_216,In_1456,In_139);
nand U217 (N_217,In_742,In_1290);
xnor U218 (N_218,In_820,In_572);
xnor U219 (N_219,In_633,In_1427);
nor U220 (N_220,In_1184,In_627);
nor U221 (N_221,In_986,In_131);
xor U222 (N_222,In_1211,In_909);
xor U223 (N_223,In_1137,In_702);
and U224 (N_224,In_211,In_566);
or U225 (N_225,In_1072,In_293);
xnor U226 (N_226,In_1253,In_1);
and U227 (N_227,In_1039,In_615);
or U228 (N_228,In_276,In_1037);
xnor U229 (N_229,In_1195,In_775);
nand U230 (N_230,In_192,In_451);
and U231 (N_231,In_592,In_722);
or U232 (N_232,In_272,In_1417);
nor U233 (N_233,In_1115,In_1225);
and U234 (N_234,In_1263,In_774);
xor U235 (N_235,In_596,In_711);
or U236 (N_236,In_800,In_267);
nand U237 (N_237,In_181,In_1426);
or U238 (N_238,In_1003,In_652);
or U239 (N_239,In_389,In_85);
nor U240 (N_240,In_503,In_413);
or U241 (N_241,In_19,In_15);
and U242 (N_242,In_1169,In_786);
xor U243 (N_243,In_1322,In_1146);
nor U244 (N_244,In_243,In_961);
nor U245 (N_245,In_173,In_347);
and U246 (N_246,In_318,In_271);
xor U247 (N_247,In_1393,In_1150);
xor U248 (N_248,In_1223,In_669);
nor U249 (N_249,In_34,In_965);
and U250 (N_250,In_1351,In_350);
or U251 (N_251,In_653,In_392);
xnor U252 (N_252,In_570,In_284);
and U253 (N_253,In_312,In_832);
nand U254 (N_254,In_260,In_790);
nor U255 (N_255,In_630,In_1478);
or U256 (N_256,In_638,In_1101);
xor U257 (N_257,In_1333,In_234);
nand U258 (N_258,In_97,In_639);
or U259 (N_259,In_737,In_709);
nand U260 (N_260,In_1465,In_713);
nor U261 (N_261,In_1181,In_104);
nor U262 (N_262,In_479,In_1042);
or U263 (N_263,In_660,In_957);
nand U264 (N_264,In_889,In_209);
xor U265 (N_265,In_1395,In_788);
nor U266 (N_266,In_343,In_1274);
nor U267 (N_267,In_18,In_1432);
or U268 (N_268,In_83,In_1475);
or U269 (N_269,In_707,In_896);
xor U270 (N_270,In_79,In_1198);
and U271 (N_271,In_757,In_951);
and U272 (N_272,In_958,In_5);
and U273 (N_273,In_804,In_1285);
xnor U274 (N_274,In_333,In_927);
nand U275 (N_275,In_1419,In_404);
and U276 (N_276,In_1031,In_1000);
and U277 (N_277,In_826,In_1259);
nand U278 (N_278,In_834,In_391);
nand U279 (N_279,In_990,In_278);
nand U280 (N_280,In_1227,In_850);
nor U281 (N_281,In_509,In_644);
nand U282 (N_282,In_187,In_933);
xnor U283 (N_283,In_661,In_1368);
nand U284 (N_284,In_1249,In_960);
or U285 (N_285,In_206,In_837);
or U286 (N_286,In_232,In_563);
and U287 (N_287,In_900,In_363);
nand U288 (N_288,In_697,In_1110);
or U289 (N_289,In_165,In_65);
xor U290 (N_290,In_1388,In_741);
xnor U291 (N_291,In_1423,In_1328);
or U292 (N_292,In_890,In_931);
xor U293 (N_293,In_1367,In_340);
and U294 (N_294,In_1136,In_700);
xnor U295 (N_295,In_191,In_1067);
or U296 (N_296,In_122,In_655);
or U297 (N_297,In_106,In_67);
nand U298 (N_298,In_33,In_1392);
nor U299 (N_299,In_567,In_643);
and U300 (N_300,In_648,In_763);
and U301 (N_301,In_628,In_100);
nor U302 (N_302,In_723,In_150);
and U303 (N_303,In_1234,In_584);
xor U304 (N_304,In_282,In_1382);
xor U305 (N_305,In_84,In_721);
nor U306 (N_306,In_956,In_991);
nand U307 (N_307,In_683,In_1277);
xor U308 (N_308,In_268,In_461);
xor U309 (N_309,In_865,In_1499);
nor U310 (N_310,In_500,In_1221);
and U311 (N_311,In_186,In_407);
nor U312 (N_312,In_134,In_1390);
nor U313 (N_313,In_601,In_136);
nor U314 (N_314,In_1289,In_1216);
xnor U315 (N_315,In_1469,In_1495);
nor U316 (N_316,In_226,In_997);
and U317 (N_317,In_1163,In_1100);
or U318 (N_318,In_1332,In_497);
xor U319 (N_319,In_1118,In_1433);
and U320 (N_320,In_614,In_651);
nor U321 (N_321,In_30,In_1018);
xnor U322 (N_322,In_1152,In_611);
or U323 (N_323,In_1228,In_378);
xnor U324 (N_324,In_1311,In_882);
nor U325 (N_325,In_442,In_1353);
nand U326 (N_326,In_807,In_725);
or U327 (N_327,In_814,In_1470);
and U328 (N_328,In_1447,In_115);
nor U329 (N_329,In_547,In_7);
nor U330 (N_330,In_427,In_887);
nor U331 (N_331,In_183,In_859);
nand U332 (N_332,In_348,In_248);
nand U333 (N_333,In_607,In_402);
and U334 (N_334,In_222,In_728);
nor U335 (N_335,In_979,In_495);
and U336 (N_336,In_386,In_536);
nand U337 (N_337,In_1261,In_1051);
nor U338 (N_338,In_1402,In_642);
and U339 (N_339,In_228,In_1358);
and U340 (N_340,In_1187,In_1193);
or U341 (N_341,In_805,In_1026);
nor U342 (N_342,In_1420,In_1222);
or U343 (N_343,In_953,In_988);
xor U344 (N_344,In_1303,In_1342);
and U345 (N_345,In_1340,In_1341);
xnor U346 (N_346,In_1307,In_1060);
and U347 (N_347,In_55,In_146);
or U348 (N_348,In_277,In_1196);
and U349 (N_349,In_128,In_80);
or U350 (N_350,In_629,In_1347);
xnor U351 (N_351,In_43,In_978);
and U352 (N_352,In_1355,In_844);
xor U353 (N_353,In_847,In_898);
and U354 (N_354,In_269,In_172);
nand U355 (N_355,In_1213,In_754);
xnor U356 (N_356,In_907,In_1032);
or U357 (N_357,In_385,In_925);
nand U358 (N_358,In_942,In_82);
nand U359 (N_359,In_412,In_585);
nor U360 (N_360,In_1010,In_421);
or U361 (N_361,In_605,In_680);
xnor U362 (N_362,In_405,In_1329);
nor U363 (N_363,In_1125,In_327);
nand U364 (N_364,In_1498,In_314);
nor U365 (N_365,In_341,In_797);
xor U366 (N_366,In_517,In_275);
nand U367 (N_367,In_1076,In_142);
nor U368 (N_368,In_480,In_993);
xnor U369 (N_369,In_1264,In_1299);
or U370 (N_370,In_435,In_789);
xor U371 (N_371,In_198,In_518);
xor U372 (N_372,In_1250,In_1444);
nand U373 (N_373,In_486,In_116);
and U374 (N_374,In_818,In_1287);
or U375 (N_375,In_1052,In_913);
nor U376 (N_376,In_1156,In_289);
nand U377 (N_377,In_681,In_622);
xor U378 (N_378,In_1260,In_1166);
nor U379 (N_379,In_227,In_1086);
or U380 (N_380,In_1422,In_242);
or U381 (N_381,In_1452,In_765);
xor U382 (N_382,In_504,In_1241);
and U383 (N_383,In_1266,In_169);
and U384 (N_384,In_437,In_817);
or U385 (N_385,In_1454,In_415);
nor U386 (N_386,In_1079,In_263);
xor U387 (N_387,In_682,In_1436);
and U388 (N_388,In_1048,In_962);
xor U389 (N_389,In_1404,In_292);
and U390 (N_390,In_1400,In_984);
or U391 (N_391,In_780,In_1077);
nand U392 (N_392,In_72,In_1191);
nor U393 (N_393,In_808,In_1199);
and U394 (N_394,In_1339,In_751);
nor U395 (N_395,In_945,In_1135);
and U396 (N_396,In_1284,In_1151);
nand U397 (N_397,In_893,In_1128);
xnor U398 (N_398,In_535,In_1036);
and U399 (N_399,In_1343,In_50);
nand U400 (N_400,In_147,In_1414);
and U401 (N_401,In_604,In_974);
or U402 (N_402,In_47,In_1002);
nor U403 (N_403,In_89,In_230);
nor U404 (N_404,In_1424,In_490);
or U405 (N_405,In_756,In_158);
xnor U406 (N_406,In_842,In_10);
nand U407 (N_407,In_213,In_760);
xnor U408 (N_408,In_995,In_463);
nor U409 (N_409,In_266,In_918);
xnor U410 (N_410,In_1095,In_1127);
xor U411 (N_411,In_1080,In_926);
nand U412 (N_412,In_654,In_739);
or U413 (N_413,In_1081,In_1105);
or U414 (N_414,In_118,In_735);
nor U415 (N_415,In_1484,In_474);
or U416 (N_416,In_38,In_1177);
and U417 (N_417,In_297,In_1324);
or U418 (N_418,In_326,In_251);
and U419 (N_419,In_441,In_456);
and U420 (N_420,In_261,In_822);
nor U421 (N_421,In_424,In_714);
nor U422 (N_422,In_491,In_1055);
xnor U423 (N_423,In_671,In_973);
xor U424 (N_424,In_98,In_334);
xnor U425 (N_425,In_151,In_1408);
xor U426 (N_426,In_157,In_853);
and U427 (N_427,In_156,In_1298);
or U428 (N_428,In_354,In_1314);
and U429 (N_429,In_464,In_793);
xor U430 (N_430,In_1435,In_534);
xnor U431 (N_431,In_704,In_915);
and U432 (N_432,In_346,In_595);
xnor U433 (N_433,In_1207,In_1386);
nor U434 (N_434,In_1439,In_919);
or U435 (N_435,In_811,In_71);
xnor U436 (N_436,In_1356,In_27);
and U437 (N_437,In_184,In_1394);
or U438 (N_438,In_1297,In_26);
or U439 (N_439,In_770,In_259);
xnor U440 (N_440,In_1212,In_1109);
nand U441 (N_441,In_1215,In_571);
or U442 (N_442,In_41,In_1237);
nand U443 (N_443,In_1295,In_776);
xnor U444 (N_444,In_189,In_399);
xor U445 (N_445,In_1231,In_819);
nand U446 (N_446,In_366,In_1204);
xnor U447 (N_447,In_1334,In_525);
or U448 (N_448,In_170,In_883);
and U449 (N_449,In_481,In_78);
or U450 (N_450,In_796,In_514);
and U451 (N_451,In_420,In_91);
or U452 (N_452,In_657,In_891);
xnor U453 (N_453,In_1301,In_1477);
xnor U454 (N_454,In_1138,In_663);
xor U455 (N_455,In_720,In_1066);
nor U456 (N_456,In_568,In_699);
xnor U457 (N_457,In_237,In_1305);
and U458 (N_458,In_1258,In_52);
or U459 (N_459,In_1153,In_632);
nand U460 (N_460,In_920,In_428);
nand U461 (N_461,In_784,In_1482);
and U462 (N_462,In_732,In_339);
nor U463 (N_463,In_787,In_901);
nand U464 (N_464,In_1162,In_193);
xor U465 (N_465,In_876,In_383);
xor U466 (N_466,In_360,In_687);
or U467 (N_467,In_1054,In_1126);
or U468 (N_468,In_897,In_1267);
nand U469 (N_469,In_101,In_996);
nor U470 (N_470,In_330,In_129);
xnor U471 (N_471,In_1164,In_575);
and U472 (N_472,In_1226,In_308);
nor U473 (N_473,In_1088,In_838);
xnor U474 (N_474,In_125,In_344);
or U475 (N_475,In_1464,In_1243);
or U476 (N_476,In_1103,In_594);
nand U477 (N_477,In_791,In_1406);
or U478 (N_478,In_1121,In_552);
nand U479 (N_479,In_117,In_744);
or U480 (N_480,In_580,In_1361);
nand U481 (N_481,In_795,In_1300);
and U482 (N_482,In_1434,In_845);
and U483 (N_483,In_1428,In_247);
nor U484 (N_484,In_1325,In_885);
and U485 (N_485,In_86,In_625);
nor U486 (N_486,In_930,In_264);
or U487 (N_487,In_328,In_1089);
xor U488 (N_488,In_528,In_194);
or U489 (N_489,In_1350,In_940);
nor U490 (N_490,In_221,In_45);
or U491 (N_491,In_878,In_1070);
nand U492 (N_492,In_1421,In_863);
nand U493 (N_493,In_781,In_299);
or U494 (N_494,In_658,In_103);
nor U495 (N_495,In_387,In_1457);
or U496 (N_496,In_1359,In_749);
and U497 (N_497,In_81,In_857);
nor U498 (N_498,In_1474,In_1168);
nand U499 (N_499,In_88,In_899);
nand U500 (N_500,In_361,In_718);
nor U501 (N_501,In_179,In_1251);
nand U502 (N_502,In_494,In_285);
or U503 (N_503,In_510,In_1306);
xor U504 (N_504,In_1270,In_337);
xor U505 (N_505,In_515,In_650);
and U506 (N_506,In_1083,In_969);
and U507 (N_507,In_698,In_963);
nand U508 (N_508,In_971,In_143);
nor U509 (N_509,In_417,In_1319);
nand U510 (N_510,In_1040,In_752);
nand U511 (N_511,In_1262,In_645);
nand U512 (N_512,In_921,In_1373);
nand U513 (N_513,In_1486,In_985);
nor U514 (N_514,In_856,In_397);
nor U515 (N_515,In_1271,In_1219);
or U516 (N_516,In_1244,In_1161);
or U517 (N_517,In_619,In_1252);
nand U518 (N_518,In_1330,In_1165);
nor U519 (N_519,In_852,In_1114);
nor U520 (N_520,In_1203,In_1208);
nor U521 (N_521,In_598,In_1410);
xor U522 (N_522,In_316,In_768);
nand U523 (N_523,In_908,In_609);
xnor U524 (N_524,In_223,In_1383);
or U525 (N_525,In_453,In_967);
and U526 (N_526,In_148,In_56);
and U527 (N_527,In_693,In_748);
nor U528 (N_528,In_668,In_493);
or U529 (N_529,In_1441,In_127);
or U530 (N_530,In_1331,In_1113);
xor U531 (N_531,In_110,In_551);
xnor U532 (N_532,In_533,In_664);
and U533 (N_533,In_1043,In_1399);
nand U534 (N_534,In_1461,In_1122);
nor U535 (N_535,In_1056,In_512);
or U536 (N_536,In_476,In_431);
or U537 (N_537,In_730,In_543);
or U538 (N_538,In_600,In_440);
and U539 (N_539,In_767,In_1206);
and U540 (N_540,In_419,In_355);
xnor U541 (N_541,In_1337,In_623);
or U542 (N_542,In_1317,In_1091);
nor U543 (N_543,In_231,In_1415);
nor U544 (N_544,In_1366,In_678);
xor U545 (N_545,In_1058,In_923);
nand U546 (N_546,In_613,In_686);
and U547 (N_547,In_670,In_894);
nor U548 (N_548,In_1061,In_621);
or U549 (N_549,In_1493,In_306);
nor U550 (N_550,In_1418,In_590);
xor U551 (N_551,In_506,In_51);
or U552 (N_552,In_468,In_532);
xor U553 (N_553,In_1192,In_452);
nand U554 (N_554,In_542,In_830);
and U555 (N_555,In_1160,In_1451);
xor U556 (N_556,In_520,In_712);
xor U557 (N_557,In_565,In_294);
xor U558 (N_558,In_549,In_1467);
nand U559 (N_559,In_96,In_764);
nand U560 (N_560,In_121,In_618);
xor U561 (N_561,In_910,In_939);
xor U562 (N_562,In_1315,In_1349);
xnor U563 (N_563,In_210,In_1133);
xor U564 (N_564,In_587,In_1471);
or U565 (N_565,In_1391,In_777);
and U566 (N_566,In_281,In_214);
or U567 (N_567,In_999,In_531);
or U568 (N_568,In_1291,In_1294);
xor U569 (N_569,In_1335,In_384);
nand U570 (N_570,In_1492,In_171);
or U571 (N_571,In_1232,In_802);
nand U572 (N_572,In_313,In_1130);
nand U573 (N_573,In_140,In_1357);
nand U574 (N_574,In_195,In_335);
nand U575 (N_575,In_154,In_349);
xnor U576 (N_576,In_325,In_180);
xnor U577 (N_577,In_810,In_943);
or U578 (N_578,In_324,In_1119);
nand U579 (N_579,In_560,In_205);
and U580 (N_580,In_869,In_1247);
and U581 (N_581,In_388,In_949);
nor U582 (N_582,In_432,In_1496);
xor U583 (N_583,In_1017,In_380);
and U584 (N_584,In_394,In_75);
nor U585 (N_585,In_801,In_291);
nand U586 (N_586,In_254,In_249);
and U587 (N_587,In_884,In_959);
or U588 (N_588,In_545,In_319);
nor U589 (N_589,In_1376,In_1069);
nor U590 (N_590,In_1186,In_403);
nand U591 (N_591,In_17,In_11);
or U592 (N_592,In_357,In_73);
nor U593 (N_593,In_416,In_467);
or U594 (N_594,In_1443,In_640);
xor U595 (N_595,In_588,In_1364);
nand U596 (N_596,In_477,In_307);
nor U597 (N_597,In_1167,In_778);
or U598 (N_598,In_1363,In_396);
nor U599 (N_599,In_736,In_583);
or U600 (N_600,In_54,In_938);
nor U601 (N_601,In_286,In_144);
xnor U602 (N_602,In_240,In_773);
or U603 (N_603,In_1075,In_168);
and U604 (N_604,In_1281,In_1490);
xor U605 (N_605,In_989,In_1265);
xnor U606 (N_606,In_1437,In_581);
nor U607 (N_607,In_200,In_1124);
nand U608 (N_608,In_133,In_561);
or U609 (N_609,In_177,In_868);
xnor U610 (N_610,In_521,In_1409);
nand U611 (N_611,In_1384,In_1021);
nand U612 (N_612,In_666,In_492);
nand U613 (N_613,In_905,In_1380);
and U614 (N_614,In_599,In_1430);
nand U615 (N_615,In_1345,In_835);
nand U616 (N_616,In_994,In_733);
or U617 (N_617,In_579,In_1463);
and U618 (N_618,In_70,In_4);
nand U619 (N_619,In_759,In_806);
or U620 (N_620,In_1139,In_544);
xnor U621 (N_621,In_564,In_1175);
or U622 (N_622,In_690,In_369);
and U623 (N_623,In_423,In_505);
or U624 (N_624,In_1316,In_356);
and U625 (N_625,In_345,In_855);
or U626 (N_626,In_235,In_861);
or U627 (N_627,In_1185,In_1112);
and U628 (N_628,In_840,In_631);
or U629 (N_629,In_1182,In_458);
nand U630 (N_630,In_1309,In_484);
nor U631 (N_631,In_1483,In_1022);
and U632 (N_632,In_603,In_162);
or U633 (N_633,In_436,In_1476);
or U634 (N_634,In_875,In_849);
xnor U635 (N_635,In_28,In_871);
and U636 (N_636,In_374,In_473);
and U637 (N_637,In_522,In_398);
nor U638 (N_638,In_692,In_1082);
or U639 (N_639,In_647,In_848);
nor U640 (N_640,In_470,In_1148);
or U641 (N_641,In_676,In_498);
xnor U642 (N_642,In_414,In_111);
and U643 (N_643,In_155,In_1024);
nand U644 (N_644,In_1006,In_408);
or U645 (N_645,In_395,In_1159);
or U646 (N_646,In_375,In_1098);
xnor U647 (N_647,In_519,In_76);
or U648 (N_648,In_0,In_1497);
or U649 (N_649,In_577,In_612);
or U650 (N_650,In_761,In_1288);
nor U651 (N_651,In_57,In_540);
or U652 (N_652,In_1092,In_411);
nand U653 (N_653,In_459,In_1378);
nor U654 (N_654,In_1248,In_1313);
xnor U655 (N_655,In_9,In_750);
nand U656 (N_656,In_359,In_689);
or U657 (N_657,In_204,In_95);
nor U658 (N_658,In_982,In_1034);
nor U659 (N_659,In_332,In_1171);
and U660 (N_660,In_29,In_472);
xor U661 (N_661,In_948,In_298);
or U662 (N_662,In_888,In_701);
xor U663 (N_663,In_322,In_1292);
nand U664 (N_664,In_1217,In_203);
and U665 (N_665,In_1176,In_244);
nand U666 (N_666,In_696,In_1011);
nor U667 (N_667,In_1445,In_1242);
xor U668 (N_668,In_548,In_1375);
nand U669 (N_669,In_1491,In_829);
nor U670 (N_670,In_252,In_1336);
nor U671 (N_671,In_727,In_944);
or U672 (N_672,In_365,In_372);
or U673 (N_673,In_1240,In_1205);
or U674 (N_674,In_872,In_541);
xnor U675 (N_675,In_928,In_1438);
and U676 (N_676,In_556,In_1001);
nand U677 (N_677,In_126,In_376);
nor U678 (N_678,In_362,In_968);
nor U679 (N_679,In_1025,In_406);
nor U680 (N_680,In_771,In_972);
or U681 (N_681,In_977,In_1201);
xor U682 (N_682,In_485,In_253);
and U683 (N_683,In_1104,In_831);
and U684 (N_684,In_1200,In_1073);
or U685 (N_685,In_1074,In_466);
or U686 (N_686,In_546,In_1189);
and U687 (N_687,In_1304,In_874);
or U688 (N_688,In_471,In_537);
nor U689 (N_689,In_877,In_679);
nand U690 (N_690,In_245,In_1411);
xnor U691 (N_691,In_1178,In_1096);
nand U692 (N_692,In_342,In_63);
or U693 (N_693,In_836,In_370);
or U694 (N_694,In_1453,In_955);
or U695 (N_695,In_576,In_1462);
or U696 (N_696,In_710,In_772);
xor U697 (N_697,In_685,In_1236);
nor U698 (N_698,In_1019,In_448);
nor U699 (N_699,In_120,In_1450);
nand U700 (N_700,In_841,In_1268);
and U701 (N_701,In_105,In_99);
and U702 (N_702,In_199,In_558);
nand U703 (N_703,In_178,In_858);
nand U704 (N_704,In_373,In_124);
nor U705 (N_705,In_20,In_946);
nor U706 (N_706,In_469,In_1308);
and U707 (N_707,In_1257,In_675);
nand U708 (N_708,In_303,In_475);
xnor U709 (N_709,In_1023,In_1027);
and U710 (N_710,In_839,In_916);
nand U711 (N_711,In_1377,In_1425);
xnor U712 (N_712,In_523,In_573);
nand U713 (N_713,In_87,In_501);
nor U714 (N_714,In_762,In_483);
or U715 (N_715,In_92,In_1296);
and U716 (N_716,In_846,In_48);
or U717 (N_717,In_1403,In_724);
or U718 (N_718,In_1321,In_1172);
xor U719 (N_719,In_758,In_559);
and U720 (N_720,In_1381,In_1310);
xor U721 (N_721,In_892,In_163);
and U722 (N_722,In_766,In_138);
nor U723 (N_723,In_646,In_1239);
and U724 (N_724,In_197,In_508);
nor U725 (N_725,In_1431,In_58);
or U726 (N_726,In_257,In_1202);
nand U727 (N_727,In_1007,In_69);
nor U728 (N_728,In_258,In_1401);
xnor U729 (N_729,In_1326,In_1144);
xor U730 (N_730,In_1473,In_1170);
xnor U731 (N_731,In_753,In_769);
xnor U732 (N_732,In_141,In_1405);
nand U733 (N_733,In_569,In_684);
or U734 (N_734,In_1344,In_287);
nor U735 (N_735,In_61,In_364);
nor U736 (N_736,In_833,In_478);
or U737 (N_737,In_59,In_112);
xnor U738 (N_738,In_64,In_539);
xor U739 (N_739,In_315,In_377);
or U740 (N_740,In_987,In_860);
and U741 (N_741,In_624,In_167);
and U742 (N_742,In_553,In_740);
or U743 (N_743,In_1302,In_1371);
xnor U744 (N_744,In_1272,In_457);
and U745 (N_745,In_1238,In_444);
xnor U746 (N_746,In_295,In_175);
nor U747 (N_747,In_130,In_1245);
or U748 (N_748,In_482,In_1229);
nand U749 (N_749,In_225,In_371);
nor U750 (N_750,In_620,In_937);
and U751 (N_751,In_1171,In_555);
or U752 (N_752,In_1365,In_585);
nand U753 (N_753,In_988,In_541);
xor U754 (N_754,In_1408,In_632);
xnor U755 (N_755,In_793,In_1238);
nand U756 (N_756,In_1024,In_563);
nand U757 (N_757,In_991,In_445);
nand U758 (N_758,In_583,In_164);
nand U759 (N_759,In_721,In_385);
nand U760 (N_760,In_892,In_975);
nand U761 (N_761,In_1000,In_1180);
and U762 (N_762,In_296,In_484);
and U763 (N_763,In_1100,In_747);
xor U764 (N_764,In_668,In_593);
nand U765 (N_765,In_1426,In_1271);
or U766 (N_766,In_889,In_785);
xnor U767 (N_767,In_826,In_559);
nor U768 (N_768,In_1001,In_204);
or U769 (N_769,In_283,In_901);
nor U770 (N_770,In_1194,In_592);
xnor U771 (N_771,In_1284,In_133);
and U772 (N_772,In_383,In_803);
or U773 (N_773,In_1009,In_1493);
nor U774 (N_774,In_429,In_1033);
and U775 (N_775,In_116,In_984);
and U776 (N_776,In_1304,In_91);
nor U777 (N_777,In_1478,In_52);
nand U778 (N_778,In_1041,In_1390);
nor U779 (N_779,In_379,In_247);
xor U780 (N_780,In_169,In_170);
or U781 (N_781,In_999,In_1084);
nor U782 (N_782,In_565,In_665);
nor U783 (N_783,In_1330,In_1350);
xor U784 (N_784,In_824,In_1352);
or U785 (N_785,In_1336,In_59);
nand U786 (N_786,In_909,In_616);
and U787 (N_787,In_863,In_1486);
and U788 (N_788,In_538,In_1038);
xnor U789 (N_789,In_1498,In_542);
or U790 (N_790,In_1250,In_38);
or U791 (N_791,In_699,In_896);
and U792 (N_792,In_985,In_967);
xor U793 (N_793,In_1117,In_1017);
nor U794 (N_794,In_774,In_837);
xnor U795 (N_795,In_783,In_1308);
nand U796 (N_796,In_171,In_1379);
or U797 (N_797,In_219,In_802);
nand U798 (N_798,In_727,In_1402);
xor U799 (N_799,In_543,In_382);
nand U800 (N_800,In_183,In_1205);
xnor U801 (N_801,In_989,In_876);
or U802 (N_802,In_581,In_180);
or U803 (N_803,In_853,In_567);
nand U804 (N_804,In_42,In_170);
and U805 (N_805,In_1462,In_233);
nor U806 (N_806,In_510,In_988);
nor U807 (N_807,In_541,In_924);
nor U808 (N_808,In_1092,In_771);
or U809 (N_809,In_1493,In_1405);
or U810 (N_810,In_1459,In_300);
and U811 (N_811,In_31,In_1304);
nand U812 (N_812,In_984,In_1116);
nor U813 (N_813,In_212,In_509);
xor U814 (N_814,In_672,In_232);
nor U815 (N_815,In_829,In_1412);
xor U816 (N_816,In_45,In_674);
or U817 (N_817,In_998,In_793);
nor U818 (N_818,In_779,In_1393);
xor U819 (N_819,In_1496,In_947);
nor U820 (N_820,In_805,In_944);
nand U821 (N_821,In_401,In_791);
xor U822 (N_822,In_604,In_732);
and U823 (N_823,In_34,In_1444);
nor U824 (N_824,In_1142,In_515);
nor U825 (N_825,In_130,In_328);
and U826 (N_826,In_917,In_1105);
xor U827 (N_827,In_448,In_679);
xor U828 (N_828,In_934,In_513);
or U829 (N_829,In_328,In_860);
nor U830 (N_830,In_1331,In_571);
or U831 (N_831,In_223,In_968);
and U832 (N_832,In_809,In_1336);
xnor U833 (N_833,In_580,In_85);
or U834 (N_834,In_311,In_1038);
xnor U835 (N_835,In_664,In_162);
or U836 (N_836,In_674,In_538);
or U837 (N_837,In_1223,In_830);
nor U838 (N_838,In_864,In_1097);
and U839 (N_839,In_142,In_869);
or U840 (N_840,In_637,In_679);
nand U841 (N_841,In_371,In_766);
nor U842 (N_842,In_476,In_1279);
or U843 (N_843,In_111,In_313);
xnor U844 (N_844,In_735,In_1088);
or U845 (N_845,In_587,In_1258);
and U846 (N_846,In_1349,In_340);
nor U847 (N_847,In_755,In_526);
or U848 (N_848,In_527,In_194);
nand U849 (N_849,In_1271,In_1477);
nor U850 (N_850,In_1387,In_1009);
nand U851 (N_851,In_1196,In_1281);
nand U852 (N_852,In_1387,In_193);
and U853 (N_853,In_460,In_922);
and U854 (N_854,In_1023,In_391);
or U855 (N_855,In_483,In_1349);
nor U856 (N_856,In_1471,In_1176);
nand U857 (N_857,In_143,In_674);
and U858 (N_858,In_1312,In_1226);
or U859 (N_859,In_164,In_354);
nor U860 (N_860,In_1209,In_16);
xnor U861 (N_861,In_75,In_827);
and U862 (N_862,In_1084,In_1479);
nor U863 (N_863,In_894,In_527);
and U864 (N_864,In_1450,In_1477);
and U865 (N_865,In_1406,In_834);
or U866 (N_866,In_288,In_564);
nor U867 (N_867,In_1015,In_609);
and U868 (N_868,In_935,In_418);
nor U869 (N_869,In_747,In_83);
xor U870 (N_870,In_1304,In_182);
xnor U871 (N_871,In_1062,In_1233);
nor U872 (N_872,In_1231,In_1264);
nand U873 (N_873,In_1056,In_911);
nand U874 (N_874,In_1004,In_661);
or U875 (N_875,In_1095,In_964);
and U876 (N_876,In_796,In_582);
xnor U877 (N_877,In_1157,In_943);
and U878 (N_878,In_1131,In_283);
and U879 (N_879,In_251,In_635);
and U880 (N_880,In_1201,In_972);
and U881 (N_881,In_547,In_773);
nor U882 (N_882,In_756,In_792);
xor U883 (N_883,In_518,In_975);
xor U884 (N_884,In_540,In_925);
or U885 (N_885,In_506,In_931);
or U886 (N_886,In_1185,In_451);
and U887 (N_887,In_890,In_992);
or U888 (N_888,In_1065,In_1205);
nor U889 (N_889,In_1176,In_1161);
nand U890 (N_890,In_1067,In_593);
xor U891 (N_891,In_399,In_1216);
xnor U892 (N_892,In_104,In_1063);
nor U893 (N_893,In_168,In_244);
nor U894 (N_894,In_415,In_426);
or U895 (N_895,In_963,In_569);
or U896 (N_896,In_1343,In_58);
or U897 (N_897,In_695,In_436);
xor U898 (N_898,In_494,In_500);
nand U899 (N_899,In_654,In_51);
nor U900 (N_900,In_56,In_763);
or U901 (N_901,In_468,In_1109);
or U902 (N_902,In_1248,In_878);
or U903 (N_903,In_1082,In_1214);
xnor U904 (N_904,In_926,In_83);
or U905 (N_905,In_781,In_649);
nand U906 (N_906,In_833,In_1141);
xnor U907 (N_907,In_911,In_929);
xnor U908 (N_908,In_288,In_829);
nand U909 (N_909,In_1137,In_208);
nand U910 (N_910,In_1424,In_318);
or U911 (N_911,In_878,In_1234);
nor U912 (N_912,In_1469,In_894);
xnor U913 (N_913,In_203,In_1178);
nand U914 (N_914,In_1020,In_78);
xor U915 (N_915,In_1012,In_1192);
or U916 (N_916,In_75,In_1347);
and U917 (N_917,In_1367,In_79);
xnor U918 (N_918,In_489,In_598);
xnor U919 (N_919,In_1319,In_569);
xor U920 (N_920,In_209,In_284);
nand U921 (N_921,In_550,In_1282);
and U922 (N_922,In_133,In_1490);
or U923 (N_923,In_210,In_828);
nor U924 (N_924,In_1212,In_1204);
xor U925 (N_925,In_788,In_643);
nor U926 (N_926,In_178,In_1109);
or U927 (N_927,In_1470,In_1145);
and U928 (N_928,In_159,In_835);
or U929 (N_929,In_99,In_218);
or U930 (N_930,In_1170,In_291);
nor U931 (N_931,In_329,In_604);
and U932 (N_932,In_1009,In_802);
or U933 (N_933,In_1098,In_1259);
nor U934 (N_934,In_335,In_922);
or U935 (N_935,In_758,In_775);
xnor U936 (N_936,In_520,In_828);
xnor U937 (N_937,In_48,In_412);
or U938 (N_938,In_1308,In_972);
nand U939 (N_939,In_1167,In_103);
or U940 (N_940,In_284,In_806);
or U941 (N_941,In_622,In_94);
nor U942 (N_942,In_268,In_1234);
nor U943 (N_943,In_525,In_1205);
and U944 (N_944,In_297,In_314);
nand U945 (N_945,In_1497,In_196);
nand U946 (N_946,In_32,In_1443);
nand U947 (N_947,In_443,In_129);
or U948 (N_948,In_698,In_288);
nand U949 (N_949,In_1059,In_436);
nor U950 (N_950,In_852,In_874);
nand U951 (N_951,In_495,In_1276);
xnor U952 (N_952,In_535,In_579);
and U953 (N_953,In_1388,In_987);
nor U954 (N_954,In_630,In_1179);
or U955 (N_955,In_454,In_1139);
and U956 (N_956,In_810,In_742);
or U957 (N_957,In_1126,In_1369);
nand U958 (N_958,In_706,In_1472);
and U959 (N_959,In_1436,In_1123);
and U960 (N_960,In_286,In_717);
or U961 (N_961,In_336,In_199);
nor U962 (N_962,In_169,In_112);
or U963 (N_963,In_1084,In_453);
xor U964 (N_964,In_752,In_1172);
nand U965 (N_965,In_826,In_1477);
and U966 (N_966,In_982,In_1352);
nand U967 (N_967,In_713,In_1261);
xor U968 (N_968,In_281,In_55);
or U969 (N_969,In_1337,In_267);
nor U970 (N_970,In_349,In_1153);
xor U971 (N_971,In_107,In_10);
nand U972 (N_972,In_844,In_474);
nor U973 (N_973,In_500,In_723);
nor U974 (N_974,In_867,In_1304);
or U975 (N_975,In_1457,In_941);
xnor U976 (N_976,In_1385,In_977);
nor U977 (N_977,In_517,In_1230);
nand U978 (N_978,In_591,In_788);
nand U979 (N_979,In_1193,In_72);
xnor U980 (N_980,In_371,In_75);
xnor U981 (N_981,In_612,In_1485);
and U982 (N_982,In_478,In_618);
and U983 (N_983,In_815,In_1081);
and U984 (N_984,In_918,In_614);
and U985 (N_985,In_1368,In_364);
or U986 (N_986,In_106,In_288);
or U987 (N_987,In_685,In_30);
nor U988 (N_988,In_55,In_223);
or U989 (N_989,In_908,In_575);
nand U990 (N_990,In_1408,In_355);
or U991 (N_991,In_1211,In_1059);
xnor U992 (N_992,In_174,In_950);
nand U993 (N_993,In_1396,In_714);
nor U994 (N_994,In_301,In_1107);
xnor U995 (N_995,In_620,In_240);
nor U996 (N_996,In_833,In_1075);
and U997 (N_997,In_272,In_292);
and U998 (N_998,In_364,In_843);
or U999 (N_999,In_561,In_322);
xor U1000 (N_1000,In_448,In_445);
and U1001 (N_1001,In_1394,In_314);
nor U1002 (N_1002,In_734,In_1443);
or U1003 (N_1003,In_366,In_1041);
nand U1004 (N_1004,In_335,In_699);
nor U1005 (N_1005,In_550,In_1171);
or U1006 (N_1006,In_768,In_1366);
and U1007 (N_1007,In_446,In_874);
or U1008 (N_1008,In_711,In_393);
and U1009 (N_1009,In_970,In_1381);
nand U1010 (N_1010,In_307,In_1041);
nand U1011 (N_1011,In_184,In_1337);
nor U1012 (N_1012,In_1085,In_1048);
nand U1013 (N_1013,In_283,In_1423);
xnor U1014 (N_1014,In_706,In_260);
and U1015 (N_1015,In_793,In_1063);
xnor U1016 (N_1016,In_23,In_614);
nand U1017 (N_1017,In_705,In_1398);
xnor U1018 (N_1018,In_574,In_1444);
nand U1019 (N_1019,In_590,In_1101);
or U1020 (N_1020,In_364,In_1283);
and U1021 (N_1021,In_970,In_1170);
nor U1022 (N_1022,In_932,In_563);
or U1023 (N_1023,In_0,In_328);
and U1024 (N_1024,In_1153,In_1380);
xnor U1025 (N_1025,In_807,In_409);
nand U1026 (N_1026,In_76,In_730);
nand U1027 (N_1027,In_907,In_219);
nand U1028 (N_1028,In_441,In_1474);
nand U1029 (N_1029,In_699,In_809);
nor U1030 (N_1030,In_438,In_1391);
or U1031 (N_1031,In_332,In_1301);
or U1032 (N_1032,In_401,In_1388);
and U1033 (N_1033,In_755,In_1160);
nand U1034 (N_1034,In_393,In_63);
nand U1035 (N_1035,In_380,In_178);
and U1036 (N_1036,In_1309,In_988);
xor U1037 (N_1037,In_1018,In_1226);
and U1038 (N_1038,In_1200,In_70);
and U1039 (N_1039,In_1162,In_1406);
nor U1040 (N_1040,In_53,In_1332);
or U1041 (N_1041,In_140,In_1322);
or U1042 (N_1042,In_705,In_918);
or U1043 (N_1043,In_887,In_377);
xnor U1044 (N_1044,In_750,In_848);
nor U1045 (N_1045,In_710,In_1020);
and U1046 (N_1046,In_516,In_980);
nor U1047 (N_1047,In_1337,In_105);
nor U1048 (N_1048,In_691,In_444);
or U1049 (N_1049,In_1265,In_1433);
nor U1050 (N_1050,In_3,In_106);
xnor U1051 (N_1051,In_1252,In_923);
and U1052 (N_1052,In_538,In_442);
or U1053 (N_1053,In_17,In_234);
xor U1054 (N_1054,In_33,In_799);
nand U1055 (N_1055,In_736,In_1343);
nor U1056 (N_1056,In_411,In_1321);
nand U1057 (N_1057,In_1451,In_513);
xor U1058 (N_1058,In_132,In_928);
and U1059 (N_1059,In_238,In_255);
or U1060 (N_1060,In_378,In_1045);
or U1061 (N_1061,In_1098,In_875);
nand U1062 (N_1062,In_1291,In_1346);
and U1063 (N_1063,In_750,In_357);
xor U1064 (N_1064,In_1296,In_1105);
nor U1065 (N_1065,In_101,In_1295);
or U1066 (N_1066,In_568,In_579);
xnor U1067 (N_1067,In_382,In_560);
nand U1068 (N_1068,In_271,In_743);
or U1069 (N_1069,In_856,In_1263);
and U1070 (N_1070,In_211,In_450);
and U1071 (N_1071,In_1356,In_111);
and U1072 (N_1072,In_859,In_1206);
or U1073 (N_1073,In_592,In_1465);
or U1074 (N_1074,In_837,In_1403);
or U1075 (N_1075,In_741,In_933);
xor U1076 (N_1076,In_789,In_1499);
and U1077 (N_1077,In_841,In_1415);
and U1078 (N_1078,In_247,In_529);
xnor U1079 (N_1079,In_802,In_857);
nand U1080 (N_1080,In_216,In_710);
and U1081 (N_1081,In_333,In_552);
nor U1082 (N_1082,In_833,In_773);
nor U1083 (N_1083,In_811,In_607);
xnor U1084 (N_1084,In_201,In_1096);
xnor U1085 (N_1085,In_1000,In_571);
and U1086 (N_1086,In_545,In_672);
nand U1087 (N_1087,In_375,In_1406);
nor U1088 (N_1088,In_316,In_823);
and U1089 (N_1089,In_397,In_1315);
xor U1090 (N_1090,In_1313,In_527);
nand U1091 (N_1091,In_83,In_208);
xor U1092 (N_1092,In_1213,In_584);
xor U1093 (N_1093,In_1238,In_871);
nand U1094 (N_1094,In_540,In_986);
xor U1095 (N_1095,In_14,In_313);
xor U1096 (N_1096,In_633,In_250);
xnor U1097 (N_1097,In_745,In_890);
and U1098 (N_1098,In_1113,In_590);
and U1099 (N_1099,In_913,In_873);
or U1100 (N_1100,In_122,In_447);
nand U1101 (N_1101,In_1063,In_759);
xnor U1102 (N_1102,In_21,In_723);
nor U1103 (N_1103,In_379,In_1351);
or U1104 (N_1104,In_857,In_391);
or U1105 (N_1105,In_1162,In_953);
and U1106 (N_1106,In_533,In_851);
nor U1107 (N_1107,In_1333,In_439);
or U1108 (N_1108,In_1132,In_1204);
and U1109 (N_1109,In_1424,In_803);
nand U1110 (N_1110,In_665,In_1090);
xnor U1111 (N_1111,In_1131,In_590);
and U1112 (N_1112,In_80,In_831);
nor U1113 (N_1113,In_1349,In_1415);
or U1114 (N_1114,In_20,In_835);
or U1115 (N_1115,In_1392,In_114);
or U1116 (N_1116,In_1224,In_704);
or U1117 (N_1117,In_0,In_810);
xor U1118 (N_1118,In_1217,In_534);
or U1119 (N_1119,In_1013,In_1185);
or U1120 (N_1120,In_946,In_834);
xor U1121 (N_1121,In_514,In_1204);
nand U1122 (N_1122,In_482,In_757);
xor U1123 (N_1123,In_1129,In_937);
or U1124 (N_1124,In_193,In_442);
nor U1125 (N_1125,In_274,In_1049);
and U1126 (N_1126,In_492,In_1455);
and U1127 (N_1127,In_1477,In_246);
and U1128 (N_1128,In_1067,In_1260);
xor U1129 (N_1129,In_1271,In_143);
and U1130 (N_1130,In_354,In_871);
nand U1131 (N_1131,In_1254,In_641);
nand U1132 (N_1132,In_131,In_1331);
xnor U1133 (N_1133,In_503,In_115);
and U1134 (N_1134,In_576,In_1037);
nor U1135 (N_1135,In_629,In_690);
nand U1136 (N_1136,In_691,In_19);
nor U1137 (N_1137,In_140,In_578);
or U1138 (N_1138,In_837,In_1136);
xor U1139 (N_1139,In_277,In_14);
nor U1140 (N_1140,In_1274,In_258);
nor U1141 (N_1141,In_72,In_1156);
xor U1142 (N_1142,In_1415,In_373);
and U1143 (N_1143,In_386,In_813);
xnor U1144 (N_1144,In_1197,In_391);
nand U1145 (N_1145,In_1481,In_1312);
and U1146 (N_1146,In_768,In_445);
xor U1147 (N_1147,In_461,In_1485);
nand U1148 (N_1148,In_180,In_727);
and U1149 (N_1149,In_106,In_591);
nand U1150 (N_1150,In_975,In_942);
or U1151 (N_1151,In_119,In_511);
xor U1152 (N_1152,In_151,In_1223);
xor U1153 (N_1153,In_267,In_91);
xor U1154 (N_1154,In_619,In_552);
nor U1155 (N_1155,In_1176,In_127);
xnor U1156 (N_1156,In_737,In_1255);
nor U1157 (N_1157,In_388,In_1118);
nor U1158 (N_1158,In_92,In_203);
xor U1159 (N_1159,In_1448,In_34);
xor U1160 (N_1160,In_335,In_717);
nand U1161 (N_1161,In_860,In_1240);
nor U1162 (N_1162,In_425,In_783);
or U1163 (N_1163,In_779,In_219);
or U1164 (N_1164,In_1317,In_562);
nand U1165 (N_1165,In_1451,In_447);
nor U1166 (N_1166,In_888,In_459);
or U1167 (N_1167,In_728,In_303);
or U1168 (N_1168,In_175,In_1421);
nor U1169 (N_1169,In_52,In_1044);
nor U1170 (N_1170,In_897,In_1032);
nor U1171 (N_1171,In_1337,In_204);
xnor U1172 (N_1172,In_1181,In_142);
nand U1173 (N_1173,In_413,In_748);
nand U1174 (N_1174,In_1171,In_1440);
and U1175 (N_1175,In_1490,In_839);
nor U1176 (N_1176,In_149,In_691);
nor U1177 (N_1177,In_536,In_2);
or U1178 (N_1178,In_7,In_658);
nand U1179 (N_1179,In_488,In_426);
xnor U1180 (N_1180,In_202,In_960);
xnor U1181 (N_1181,In_869,In_99);
nor U1182 (N_1182,In_467,In_199);
nor U1183 (N_1183,In_1252,In_846);
or U1184 (N_1184,In_1379,In_986);
nor U1185 (N_1185,In_1276,In_523);
nor U1186 (N_1186,In_877,In_653);
nor U1187 (N_1187,In_856,In_149);
or U1188 (N_1188,In_1379,In_221);
xor U1189 (N_1189,In_1411,In_1210);
or U1190 (N_1190,In_717,In_217);
xnor U1191 (N_1191,In_1036,In_1254);
or U1192 (N_1192,In_975,In_106);
nand U1193 (N_1193,In_554,In_1208);
and U1194 (N_1194,In_107,In_1336);
or U1195 (N_1195,In_811,In_491);
nor U1196 (N_1196,In_159,In_860);
or U1197 (N_1197,In_1393,In_877);
nand U1198 (N_1198,In_50,In_1106);
and U1199 (N_1199,In_426,In_401);
or U1200 (N_1200,In_1477,In_1250);
and U1201 (N_1201,In_146,In_405);
nor U1202 (N_1202,In_622,In_867);
xnor U1203 (N_1203,In_1449,In_663);
or U1204 (N_1204,In_1279,In_1337);
and U1205 (N_1205,In_13,In_362);
nor U1206 (N_1206,In_582,In_554);
nand U1207 (N_1207,In_1352,In_1150);
and U1208 (N_1208,In_1062,In_18);
and U1209 (N_1209,In_1337,In_610);
and U1210 (N_1210,In_1139,In_810);
nand U1211 (N_1211,In_477,In_526);
xnor U1212 (N_1212,In_1126,In_320);
and U1213 (N_1213,In_1387,In_711);
and U1214 (N_1214,In_425,In_942);
and U1215 (N_1215,In_617,In_713);
or U1216 (N_1216,In_1391,In_1327);
nor U1217 (N_1217,In_1440,In_805);
nand U1218 (N_1218,In_1285,In_1199);
xnor U1219 (N_1219,In_253,In_387);
and U1220 (N_1220,In_965,In_500);
xor U1221 (N_1221,In_666,In_586);
or U1222 (N_1222,In_454,In_360);
and U1223 (N_1223,In_1120,In_517);
nor U1224 (N_1224,In_1056,In_789);
nand U1225 (N_1225,In_176,In_118);
xor U1226 (N_1226,In_762,In_439);
xor U1227 (N_1227,In_898,In_282);
xor U1228 (N_1228,In_312,In_1493);
xor U1229 (N_1229,In_1120,In_465);
or U1230 (N_1230,In_1254,In_997);
nor U1231 (N_1231,In_887,In_1012);
or U1232 (N_1232,In_642,In_395);
and U1233 (N_1233,In_934,In_130);
nand U1234 (N_1234,In_1145,In_1455);
nand U1235 (N_1235,In_1343,In_919);
or U1236 (N_1236,In_143,In_742);
xnor U1237 (N_1237,In_747,In_1120);
or U1238 (N_1238,In_27,In_852);
nor U1239 (N_1239,In_1420,In_1237);
or U1240 (N_1240,In_952,In_478);
nand U1241 (N_1241,In_891,In_236);
nor U1242 (N_1242,In_1326,In_1377);
nand U1243 (N_1243,In_1420,In_90);
xor U1244 (N_1244,In_866,In_1296);
and U1245 (N_1245,In_132,In_1140);
and U1246 (N_1246,In_1004,In_343);
xor U1247 (N_1247,In_1170,In_782);
nor U1248 (N_1248,In_1352,In_1302);
nand U1249 (N_1249,In_1194,In_980);
nor U1250 (N_1250,In_523,In_136);
nand U1251 (N_1251,In_1178,In_763);
xor U1252 (N_1252,In_1163,In_1202);
nand U1253 (N_1253,In_452,In_1411);
or U1254 (N_1254,In_385,In_436);
nand U1255 (N_1255,In_613,In_385);
or U1256 (N_1256,In_1193,In_578);
xnor U1257 (N_1257,In_147,In_1242);
nor U1258 (N_1258,In_1326,In_72);
xor U1259 (N_1259,In_227,In_551);
and U1260 (N_1260,In_1062,In_1286);
and U1261 (N_1261,In_895,In_1227);
nor U1262 (N_1262,In_622,In_1119);
or U1263 (N_1263,In_231,In_349);
nand U1264 (N_1264,In_83,In_557);
nor U1265 (N_1265,In_1032,In_440);
or U1266 (N_1266,In_1343,In_193);
nand U1267 (N_1267,In_1220,In_700);
or U1268 (N_1268,In_212,In_1246);
nand U1269 (N_1269,In_379,In_988);
xnor U1270 (N_1270,In_247,In_398);
or U1271 (N_1271,In_315,In_12);
and U1272 (N_1272,In_1399,In_57);
nor U1273 (N_1273,In_1357,In_566);
xnor U1274 (N_1274,In_394,In_520);
and U1275 (N_1275,In_488,In_568);
nand U1276 (N_1276,In_645,In_746);
and U1277 (N_1277,In_26,In_1200);
nand U1278 (N_1278,In_997,In_1207);
or U1279 (N_1279,In_162,In_791);
and U1280 (N_1280,In_439,In_413);
and U1281 (N_1281,In_848,In_668);
nand U1282 (N_1282,In_209,In_447);
and U1283 (N_1283,In_579,In_684);
or U1284 (N_1284,In_828,In_1318);
nor U1285 (N_1285,In_485,In_761);
xnor U1286 (N_1286,In_848,In_1480);
xor U1287 (N_1287,In_820,In_622);
nand U1288 (N_1288,In_1305,In_1093);
nand U1289 (N_1289,In_859,In_504);
xnor U1290 (N_1290,In_77,In_931);
xor U1291 (N_1291,In_1056,In_1372);
or U1292 (N_1292,In_825,In_708);
nand U1293 (N_1293,In_172,In_1052);
or U1294 (N_1294,In_760,In_1297);
nor U1295 (N_1295,In_391,In_1438);
nor U1296 (N_1296,In_897,In_416);
and U1297 (N_1297,In_1398,In_595);
nor U1298 (N_1298,In_438,In_1087);
and U1299 (N_1299,In_1312,In_1005);
or U1300 (N_1300,In_579,In_1029);
nor U1301 (N_1301,In_896,In_653);
nand U1302 (N_1302,In_271,In_804);
nand U1303 (N_1303,In_1230,In_1342);
nand U1304 (N_1304,In_1172,In_1230);
or U1305 (N_1305,In_757,In_1096);
or U1306 (N_1306,In_964,In_1192);
or U1307 (N_1307,In_138,In_914);
nor U1308 (N_1308,In_1005,In_1282);
xnor U1309 (N_1309,In_647,In_146);
nor U1310 (N_1310,In_1264,In_119);
or U1311 (N_1311,In_1103,In_599);
or U1312 (N_1312,In_217,In_1370);
nor U1313 (N_1313,In_1131,In_878);
or U1314 (N_1314,In_365,In_376);
xnor U1315 (N_1315,In_271,In_1443);
and U1316 (N_1316,In_1196,In_166);
and U1317 (N_1317,In_1446,In_612);
nor U1318 (N_1318,In_643,In_1305);
and U1319 (N_1319,In_201,In_1392);
and U1320 (N_1320,In_671,In_602);
xnor U1321 (N_1321,In_1279,In_77);
or U1322 (N_1322,In_287,In_761);
nand U1323 (N_1323,In_949,In_557);
or U1324 (N_1324,In_244,In_287);
and U1325 (N_1325,In_1401,In_1013);
nand U1326 (N_1326,In_717,In_1413);
xnor U1327 (N_1327,In_516,In_491);
or U1328 (N_1328,In_863,In_248);
and U1329 (N_1329,In_730,In_529);
nor U1330 (N_1330,In_1061,In_268);
and U1331 (N_1331,In_1055,In_1414);
nor U1332 (N_1332,In_502,In_66);
or U1333 (N_1333,In_17,In_790);
xnor U1334 (N_1334,In_970,In_976);
or U1335 (N_1335,In_777,In_836);
nand U1336 (N_1336,In_937,In_680);
and U1337 (N_1337,In_229,In_664);
nor U1338 (N_1338,In_168,In_600);
nor U1339 (N_1339,In_461,In_526);
xnor U1340 (N_1340,In_642,In_265);
nor U1341 (N_1341,In_226,In_276);
and U1342 (N_1342,In_1035,In_606);
or U1343 (N_1343,In_1164,In_924);
xor U1344 (N_1344,In_1133,In_17);
and U1345 (N_1345,In_90,In_1301);
xor U1346 (N_1346,In_1451,In_517);
or U1347 (N_1347,In_399,In_1050);
and U1348 (N_1348,In_1335,In_202);
nor U1349 (N_1349,In_768,In_1260);
nand U1350 (N_1350,In_670,In_1417);
nand U1351 (N_1351,In_856,In_815);
xor U1352 (N_1352,In_77,In_230);
or U1353 (N_1353,In_330,In_1101);
xnor U1354 (N_1354,In_10,In_449);
and U1355 (N_1355,In_1015,In_749);
and U1356 (N_1356,In_140,In_173);
nor U1357 (N_1357,In_1384,In_950);
and U1358 (N_1358,In_476,In_1308);
nor U1359 (N_1359,In_403,In_1050);
and U1360 (N_1360,In_1320,In_400);
nor U1361 (N_1361,In_33,In_1172);
nand U1362 (N_1362,In_513,In_1491);
nor U1363 (N_1363,In_1456,In_1203);
and U1364 (N_1364,In_699,In_291);
nand U1365 (N_1365,In_1403,In_570);
xor U1366 (N_1366,In_1253,In_703);
xor U1367 (N_1367,In_96,In_146);
xnor U1368 (N_1368,In_444,In_180);
xnor U1369 (N_1369,In_10,In_1134);
or U1370 (N_1370,In_332,In_1003);
and U1371 (N_1371,In_1481,In_1375);
and U1372 (N_1372,In_1432,In_667);
xnor U1373 (N_1373,In_638,In_1239);
nor U1374 (N_1374,In_463,In_183);
nor U1375 (N_1375,In_107,In_1310);
nor U1376 (N_1376,In_692,In_1362);
or U1377 (N_1377,In_249,In_294);
xnor U1378 (N_1378,In_537,In_757);
nor U1379 (N_1379,In_402,In_560);
nand U1380 (N_1380,In_233,In_104);
xnor U1381 (N_1381,In_789,In_1457);
or U1382 (N_1382,In_40,In_746);
or U1383 (N_1383,In_557,In_1408);
nor U1384 (N_1384,In_1235,In_1351);
nor U1385 (N_1385,In_336,In_394);
and U1386 (N_1386,In_1000,In_1431);
nor U1387 (N_1387,In_154,In_1413);
or U1388 (N_1388,In_33,In_186);
nor U1389 (N_1389,In_673,In_1454);
or U1390 (N_1390,In_1446,In_76);
and U1391 (N_1391,In_518,In_1095);
nor U1392 (N_1392,In_866,In_802);
xor U1393 (N_1393,In_817,In_911);
or U1394 (N_1394,In_180,In_207);
or U1395 (N_1395,In_62,In_362);
nand U1396 (N_1396,In_1276,In_1390);
and U1397 (N_1397,In_1146,In_1162);
nand U1398 (N_1398,In_353,In_645);
nand U1399 (N_1399,In_30,In_1434);
or U1400 (N_1400,In_1444,In_282);
nand U1401 (N_1401,In_842,In_477);
nand U1402 (N_1402,In_977,In_1426);
and U1403 (N_1403,In_310,In_1385);
and U1404 (N_1404,In_137,In_518);
or U1405 (N_1405,In_86,In_844);
nor U1406 (N_1406,In_1326,In_21);
and U1407 (N_1407,In_289,In_1079);
and U1408 (N_1408,In_571,In_138);
nand U1409 (N_1409,In_1485,In_1291);
or U1410 (N_1410,In_192,In_916);
nor U1411 (N_1411,In_1207,In_865);
xor U1412 (N_1412,In_598,In_26);
or U1413 (N_1413,In_410,In_166);
and U1414 (N_1414,In_787,In_1233);
nor U1415 (N_1415,In_1247,In_194);
and U1416 (N_1416,In_741,In_764);
xnor U1417 (N_1417,In_416,In_1186);
xor U1418 (N_1418,In_1104,In_331);
nor U1419 (N_1419,In_319,In_866);
or U1420 (N_1420,In_330,In_298);
or U1421 (N_1421,In_1033,In_871);
nand U1422 (N_1422,In_633,In_1307);
nand U1423 (N_1423,In_507,In_396);
or U1424 (N_1424,In_203,In_344);
and U1425 (N_1425,In_994,In_1184);
or U1426 (N_1426,In_278,In_247);
or U1427 (N_1427,In_1256,In_1102);
nand U1428 (N_1428,In_395,In_1175);
nor U1429 (N_1429,In_867,In_789);
or U1430 (N_1430,In_1129,In_239);
or U1431 (N_1431,In_884,In_1025);
or U1432 (N_1432,In_959,In_987);
nor U1433 (N_1433,In_921,In_988);
and U1434 (N_1434,In_1424,In_403);
nor U1435 (N_1435,In_357,In_925);
and U1436 (N_1436,In_909,In_141);
xor U1437 (N_1437,In_468,In_1373);
nand U1438 (N_1438,In_230,In_1165);
nor U1439 (N_1439,In_393,In_1367);
nand U1440 (N_1440,In_415,In_1354);
nor U1441 (N_1441,In_1263,In_7);
nand U1442 (N_1442,In_125,In_549);
nand U1443 (N_1443,In_334,In_1496);
nand U1444 (N_1444,In_619,In_396);
nand U1445 (N_1445,In_1446,In_738);
nand U1446 (N_1446,In_189,In_954);
or U1447 (N_1447,In_1031,In_1313);
xnor U1448 (N_1448,In_1204,In_1247);
xnor U1449 (N_1449,In_176,In_1436);
and U1450 (N_1450,In_1140,In_586);
xnor U1451 (N_1451,In_726,In_1318);
or U1452 (N_1452,In_1318,In_1490);
nand U1453 (N_1453,In_1478,In_692);
nor U1454 (N_1454,In_1085,In_104);
nor U1455 (N_1455,In_118,In_1196);
and U1456 (N_1456,In_926,In_868);
nand U1457 (N_1457,In_1045,In_699);
xor U1458 (N_1458,In_615,In_514);
or U1459 (N_1459,In_894,In_1226);
or U1460 (N_1460,In_1329,In_1397);
and U1461 (N_1461,In_434,In_314);
xnor U1462 (N_1462,In_374,In_895);
nor U1463 (N_1463,In_78,In_818);
xnor U1464 (N_1464,In_811,In_1398);
and U1465 (N_1465,In_1498,In_780);
or U1466 (N_1466,In_119,In_265);
nand U1467 (N_1467,In_1022,In_478);
xnor U1468 (N_1468,In_166,In_90);
nand U1469 (N_1469,In_14,In_1014);
nand U1470 (N_1470,In_1235,In_682);
xor U1471 (N_1471,In_603,In_852);
xnor U1472 (N_1472,In_334,In_921);
nor U1473 (N_1473,In_556,In_1296);
xor U1474 (N_1474,In_369,In_3);
xor U1475 (N_1475,In_390,In_307);
nand U1476 (N_1476,In_1348,In_646);
nor U1477 (N_1477,In_442,In_1339);
xor U1478 (N_1478,In_638,In_471);
xnor U1479 (N_1479,In_1235,In_299);
xnor U1480 (N_1480,In_964,In_533);
and U1481 (N_1481,In_788,In_627);
nor U1482 (N_1482,In_785,In_928);
nor U1483 (N_1483,In_489,In_58);
xor U1484 (N_1484,In_105,In_309);
or U1485 (N_1485,In_1195,In_992);
nor U1486 (N_1486,In_1483,In_931);
xnor U1487 (N_1487,In_1364,In_288);
and U1488 (N_1488,In_979,In_88);
or U1489 (N_1489,In_652,In_54);
nand U1490 (N_1490,In_559,In_323);
and U1491 (N_1491,In_1387,In_169);
xnor U1492 (N_1492,In_583,In_1347);
xnor U1493 (N_1493,In_671,In_633);
nand U1494 (N_1494,In_249,In_241);
nand U1495 (N_1495,In_569,In_957);
nor U1496 (N_1496,In_643,In_848);
nand U1497 (N_1497,In_1262,In_1192);
or U1498 (N_1498,In_83,In_1288);
nor U1499 (N_1499,In_766,In_784);
xor U1500 (N_1500,N_792,N_740);
nor U1501 (N_1501,N_1027,N_374);
nor U1502 (N_1502,N_1187,N_858);
xor U1503 (N_1503,N_818,N_447);
and U1504 (N_1504,N_1390,N_90);
nand U1505 (N_1505,N_822,N_640);
xor U1506 (N_1506,N_1226,N_1266);
and U1507 (N_1507,N_796,N_1100);
or U1508 (N_1508,N_1475,N_1158);
xnor U1509 (N_1509,N_264,N_1119);
xnor U1510 (N_1510,N_1261,N_377);
nand U1511 (N_1511,N_450,N_1265);
xnor U1512 (N_1512,N_61,N_632);
nand U1513 (N_1513,N_314,N_357);
xor U1514 (N_1514,N_203,N_1301);
xnor U1515 (N_1515,N_1327,N_252);
or U1516 (N_1516,N_139,N_1026);
and U1517 (N_1517,N_616,N_948);
nor U1518 (N_1518,N_1370,N_920);
xnor U1519 (N_1519,N_267,N_835);
xnor U1520 (N_1520,N_407,N_915);
nand U1521 (N_1521,N_1238,N_1395);
and U1522 (N_1522,N_1016,N_83);
or U1523 (N_1523,N_1409,N_806);
nand U1524 (N_1524,N_70,N_378);
nor U1525 (N_1525,N_927,N_1448);
xnor U1526 (N_1526,N_899,N_1352);
or U1527 (N_1527,N_958,N_843);
and U1528 (N_1528,N_1242,N_1224);
nand U1529 (N_1529,N_0,N_1249);
nor U1530 (N_1530,N_313,N_1223);
xor U1531 (N_1531,N_700,N_355);
nor U1532 (N_1532,N_112,N_74);
xor U1533 (N_1533,N_986,N_1112);
nor U1534 (N_1534,N_1302,N_260);
and U1535 (N_1535,N_541,N_1392);
xor U1536 (N_1536,N_1099,N_1414);
xnor U1537 (N_1537,N_1366,N_922);
xor U1538 (N_1538,N_1332,N_1058);
and U1539 (N_1539,N_1123,N_1313);
xnor U1540 (N_1540,N_790,N_1470);
nand U1541 (N_1541,N_215,N_837);
nand U1542 (N_1542,N_815,N_857);
nand U1543 (N_1543,N_552,N_869);
nand U1544 (N_1544,N_530,N_103);
or U1545 (N_1545,N_914,N_610);
xnor U1546 (N_1546,N_570,N_380);
and U1547 (N_1547,N_393,N_285);
nor U1548 (N_1548,N_1021,N_697);
and U1549 (N_1549,N_84,N_1008);
nand U1550 (N_1550,N_344,N_743);
nor U1551 (N_1551,N_46,N_636);
xor U1552 (N_1552,N_1157,N_852);
nand U1553 (N_1553,N_269,N_68);
nor U1554 (N_1554,N_1499,N_472);
nand U1555 (N_1555,N_1193,N_1437);
xor U1556 (N_1556,N_134,N_578);
or U1557 (N_1557,N_404,N_4);
xor U1558 (N_1558,N_270,N_412);
nor U1559 (N_1559,N_1346,N_1329);
nor U1560 (N_1560,N_435,N_508);
nor U1561 (N_1561,N_575,N_902);
xnor U1562 (N_1562,N_1270,N_1036);
nor U1563 (N_1563,N_545,N_1046);
nand U1564 (N_1564,N_710,N_746);
and U1565 (N_1565,N_750,N_691);
nor U1566 (N_1566,N_672,N_606);
nor U1567 (N_1567,N_918,N_943);
or U1568 (N_1568,N_135,N_1479);
or U1569 (N_1569,N_1154,N_434);
or U1570 (N_1570,N_906,N_1280);
and U1571 (N_1571,N_438,N_542);
and U1572 (N_1572,N_1048,N_1330);
nor U1573 (N_1573,N_133,N_81);
nand U1574 (N_1574,N_224,N_1398);
or U1575 (N_1575,N_753,N_1375);
xnor U1576 (N_1576,N_535,N_1296);
nand U1577 (N_1577,N_905,N_1387);
and U1578 (N_1578,N_779,N_887);
nand U1579 (N_1579,N_167,N_589);
nand U1580 (N_1580,N_1439,N_851);
nor U1581 (N_1581,N_395,N_860);
or U1582 (N_1582,N_536,N_396);
nor U1583 (N_1583,N_680,N_1424);
or U1584 (N_1584,N_1294,N_97);
xor U1585 (N_1585,N_565,N_834);
nand U1586 (N_1586,N_1004,N_946);
xnor U1587 (N_1587,N_480,N_1304);
or U1588 (N_1588,N_644,N_349);
nor U1589 (N_1589,N_350,N_894);
nor U1590 (N_1590,N_443,N_1369);
nor U1591 (N_1591,N_312,N_641);
and U1592 (N_1592,N_853,N_253);
nor U1593 (N_1593,N_1068,N_701);
and U1594 (N_1594,N_26,N_772);
xor U1595 (N_1595,N_343,N_86);
nor U1596 (N_1596,N_1441,N_7);
nand U1597 (N_1597,N_1221,N_392);
nor U1598 (N_1598,N_1396,N_1140);
nor U1599 (N_1599,N_159,N_1305);
nor U1600 (N_1600,N_24,N_1397);
nor U1601 (N_1601,N_984,N_829);
and U1602 (N_1602,N_1477,N_1417);
and U1603 (N_1603,N_1324,N_1188);
nand U1604 (N_1604,N_603,N_954);
nor U1605 (N_1605,N_328,N_96);
nand U1606 (N_1606,N_573,N_247);
xor U1607 (N_1607,N_874,N_330);
and U1608 (N_1608,N_1174,N_1380);
and U1609 (N_1609,N_271,N_297);
nand U1610 (N_1610,N_85,N_153);
or U1611 (N_1611,N_1148,N_141);
xor U1612 (N_1612,N_1049,N_891);
xor U1613 (N_1613,N_645,N_635);
xnor U1614 (N_1614,N_888,N_1385);
xor U1615 (N_1615,N_960,N_816);
xor U1616 (N_1616,N_1117,N_1394);
or U1617 (N_1617,N_382,N_953);
nor U1618 (N_1618,N_1128,N_992);
nand U1619 (N_1619,N_1368,N_12);
xor U1620 (N_1620,N_165,N_1338);
and U1621 (N_1621,N_388,N_1285);
or U1622 (N_1622,N_1271,N_411);
nor U1623 (N_1623,N_939,N_1045);
xnor U1624 (N_1624,N_912,N_1126);
nand U1625 (N_1625,N_130,N_1497);
nor U1626 (N_1626,N_705,N_1198);
xor U1627 (N_1627,N_65,N_93);
or U1628 (N_1628,N_774,N_830);
nor U1629 (N_1629,N_819,N_1015);
nand U1630 (N_1630,N_582,N_1062);
nor U1631 (N_1631,N_662,N_403);
nand U1632 (N_1632,N_1156,N_1463);
nand U1633 (N_1633,N_773,N_1020);
xnor U1634 (N_1634,N_1443,N_136);
nand U1635 (N_1635,N_223,N_122);
or U1636 (N_1636,N_1011,N_677);
xor U1637 (N_1637,N_21,N_166);
and U1638 (N_1638,N_1044,N_1371);
nand U1639 (N_1639,N_770,N_526);
and U1640 (N_1640,N_1064,N_272);
xnor U1641 (N_1641,N_544,N_651);
and U1642 (N_1642,N_1006,N_277);
nand U1643 (N_1643,N_1209,N_352);
xnor U1644 (N_1644,N_1031,N_696);
xnor U1645 (N_1645,N_311,N_1225);
nand U1646 (N_1646,N_1430,N_967);
or U1647 (N_1647,N_1365,N_771);
nor U1648 (N_1648,N_690,N_319);
nand U1649 (N_1649,N_703,N_1466);
or U1650 (N_1650,N_336,N_512);
nand U1651 (N_1651,N_455,N_415);
nor U1652 (N_1652,N_793,N_409);
nor U1653 (N_1653,N_1127,N_975);
and U1654 (N_1654,N_346,N_502);
nand U1655 (N_1655,N_279,N_34);
nand U1656 (N_1656,N_1235,N_600);
nand U1657 (N_1657,N_685,N_278);
or U1658 (N_1658,N_591,N_1061);
and U1659 (N_1659,N_1095,N_687);
nor U1660 (N_1660,N_187,N_384);
or U1661 (N_1661,N_622,N_893);
and U1662 (N_1662,N_1267,N_298);
or U1663 (N_1663,N_1388,N_1149);
and U1664 (N_1664,N_451,N_1491);
and U1665 (N_1665,N_440,N_257);
nor U1666 (N_1666,N_156,N_1292);
and U1667 (N_1667,N_33,N_569);
xor U1668 (N_1668,N_1022,N_219);
xnor U1669 (N_1669,N_515,N_1216);
xnor U1670 (N_1670,N_307,N_588);
nor U1671 (N_1671,N_94,N_716);
xor U1672 (N_1672,N_1108,N_1070);
nand U1673 (N_1673,N_1336,N_332);
nand U1674 (N_1674,N_143,N_1263);
xor U1675 (N_1675,N_1075,N_9);
xor U1676 (N_1676,N_491,N_522);
or U1677 (N_1677,N_627,N_1239);
nand U1678 (N_1678,N_1217,N_1245);
nand U1679 (N_1679,N_410,N_1166);
and U1680 (N_1680,N_1040,N_1350);
and U1681 (N_1681,N_699,N_500);
and U1682 (N_1682,N_423,N_1106);
nor U1683 (N_1683,N_52,N_1401);
nor U1684 (N_1684,N_454,N_164);
nand U1685 (N_1685,N_549,N_855);
nand U1686 (N_1686,N_1384,N_574);
nand U1687 (N_1687,N_1186,N_1);
and U1688 (N_1688,N_1115,N_638);
or U1689 (N_1689,N_712,N_125);
nand U1690 (N_1690,N_1143,N_1323);
or U1691 (N_1691,N_748,N_580);
nand U1692 (N_1692,N_1078,N_901);
nor U1693 (N_1693,N_754,N_1257);
xnor U1694 (N_1694,N_1185,N_1234);
nor U1695 (N_1695,N_1339,N_251);
nor U1696 (N_1696,N_1110,N_266);
or U1697 (N_1697,N_209,N_431);
xnor U1698 (N_1698,N_683,N_528);
nand U1699 (N_1699,N_559,N_840);
or U1700 (N_1700,N_496,N_1103);
or U1701 (N_1701,N_1118,N_157);
nor U1702 (N_1702,N_318,N_1152);
or U1703 (N_1703,N_262,N_624);
or U1704 (N_1704,N_182,N_405);
and U1705 (N_1705,N_1273,N_1449);
nor U1706 (N_1706,N_1207,N_904);
nor U1707 (N_1707,N_487,N_206);
nor U1708 (N_1708,N_788,N_1383);
xnor U1709 (N_1709,N_809,N_493);
nand U1710 (N_1710,N_78,N_1467);
nand U1711 (N_1711,N_720,N_227);
nand U1712 (N_1712,N_465,N_1403);
xnor U1713 (N_1713,N_1101,N_733);
nand U1714 (N_1714,N_129,N_947);
nor U1715 (N_1715,N_1317,N_482);
nand U1716 (N_1716,N_463,N_196);
and U1717 (N_1717,N_873,N_230);
nand U1718 (N_1718,N_814,N_55);
and U1719 (N_1719,N_637,N_492);
and U1720 (N_1720,N_16,N_876);
nand U1721 (N_1721,N_1136,N_198);
nand U1722 (N_1722,N_999,N_1476);
and U1723 (N_1723,N_471,N_1325);
and U1724 (N_1724,N_205,N_657);
nor U1725 (N_1725,N_604,N_1051);
or U1726 (N_1726,N_646,N_885);
and U1727 (N_1727,N_1113,N_969);
or U1728 (N_1728,N_306,N_137);
nor U1729 (N_1729,N_989,N_1462);
or U1730 (N_1730,N_1460,N_1408);
and U1731 (N_1731,N_120,N_79);
xnor U1732 (N_1732,N_1130,N_1013);
or U1733 (N_1733,N_803,N_1129);
or U1734 (N_1734,N_76,N_427);
xnor U1735 (N_1735,N_674,N_1256);
or U1736 (N_1736,N_1247,N_254);
nor U1737 (N_1737,N_861,N_188);
nor U1738 (N_1738,N_654,N_501);
and U1739 (N_1739,N_1423,N_725);
xor U1740 (N_1740,N_1125,N_89);
nand U1741 (N_1741,N_414,N_397);
nor U1742 (N_1742,N_351,N_560);
and U1743 (N_1743,N_163,N_1452);
nand U1744 (N_1744,N_1167,N_1486);
nand U1745 (N_1745,N_111,N_1233);
and U1746 (N_1746,N_190,N_671);
xor U1747 (N_1747,N_1243,N_147);
nor U1748 (N_1748,N_590,N_1047);
and U1749 (N_1749,N_579,N_903);
xor U1750 (N_1750,N_1295,N_1244);
nand U1751 (N_1751,N_113,N_634);
xnor U1752 (N_1752,N_218,N_221);
and U1753 (N_1753,N_320,N_1083);
xor U1754 (N_1754,N_1057,N_577);
and U1755 (N_1755,N_974,N_1073);
xor U1756 (N_1756,N_174,N_1309);
xor U1757 (N_1757,N_1354,N_1429);
and U1758 (N_1758,N_1144,N_42);
or U1759 (N_1759,N_1298,N_211);
xnor U1760 (N_1760,N_1411,N_1469);
and U1761 (N_1761,N_963,N_1105);
or U1762 (N_1762,N_759,N_738);
nand U1763 (N_1763,N_115,N_785);
nor U1764 (N_1764,N_280,N_323);
and U1765 (N_1765,N_875,N_381);
or U1766 (N_1766,N_1168,N_356);
nor U1767 (N_1767,N_1382,N_399);
and U1768 (N_1768,N_919,N_1192);
xnor U1769 (N_1769,N_1372,N_132);
xnor U1770 (N_1770,N_1311,N_178);
xor U1771 (N_1771,N_365,N_694);
or U1772 (N_1772,N_1010,N_370);
xnor U1773 (N_1773,N_114,N_879);
and U1774 (N_1774,N_1229,N_1341);
nand U1775 (N_1775,N_1089,N_1321);
and U1776 (N_1776,N_444,N_765);
nand U1777 (N_1777,N_527,N_688);
nor U1778 (N_1778,N_1150,N_826);
xnor U1779 (N_1779,N_1173,N_232);
and U1780 (N_1780,N_239,N_742);
or U1781 (N_1781,N_878,N_109);
and U1782 (N_1782,N_630,N_308);
and U1783 (N_1783,N_1310,N_1287);
nand U1784 (N_1784,N_1155,N_1445);
xor U1785 (N_1785,N_1056,N_1237);
nand U1786 (N_1786,N_564,N_171);
nor U1787 (N_1787,N_185,N_123);
xnor U1788 (N_1788,N_341,N_398);
nand U1789 (N_1789,N_75,N_626);
nand U1790 (N_1790,N_537,N_149);
nand U1791 (N_1791,N_186,N_489);
nor U1792 (N_1792,N_841,N_666);
and U1793 (N_1793,N_889,N_1190);
and U1794 (N_1794,N_309,N_62);
or U1795 (N_1795,N_305,N_301);
nor U1796 (N_1796,N_1326,N_1059);
xor U1797 (N_1797,N_1279,N_1389);
and U1798 (N_1798,N_661,N_464);
nor U1799 (N_1799,N_1335,N_1374);
nor U1800 (N_1800,N_428,N_908);
and U1801 (N_1801,N_1351,N_1307);
or U1802 (N_1802,N_1005,N_871);
nand U1803 (N_1803,N_576,N_99);
nor U1804 (N_1804,N_776,N_757);
or U1805 (N_1805,N_48,N_821);
or U1806 (N_1806,N_1286,N_25);
xnor U1807 (N_1807,N_1253,N_1032);
xnor U1808 (N_1808,N_18,N_562);
nor U1809 (N_1809,N_926,N_595);
nand U1810 (N_1810,N_1137,N_1161);
or U1811 (N_1811,N_106,N_895);
and U1812 (N_1812,N_828,N_191);
xnor U1813 (N_1813,N_838,N_514);
nor U1814 (N_1814,N_794,N_35);
xnor U1815 (N_1815,N_1050,N_1412);
or U1816 (N_1816,N_1391,N_1222);
xor U1817 (N_1817,N_1163,N_583);
xnor U1818 (N_1818,N_1054,N_1200);
nand U1819 (N_1819,N_194,N_726);
and U1820 (N_1820,N_599,N_854);
xor U1821 (N_1821,N_1171,N_242);
or U1822 (N_1822,N_1197,N_650);
nand U1823 (N_1823,N_286,N_836);
or U1824 (N_1824,N_1175,N_928);
and U1825 (N_1825,N_824,N_965);
or U1826 (N_1826,N_59,N_1483);
nor U1827 (N_1827,N_909,N_972);
nand U1828 (N_1828,N_1450,N_364);
and U1829 (N_1829,N_1357,N_1342);
and U1830 (N_1830,N_56,N_6);
nand U1831 (N_1831,N_181,N_789);
nor U1832 (N_1832,N_767,N_2);
and U1833 (N_1833,N_1146,N_248);
and U1834 (N_1834,N_353,N_87);
nand U1835 (N_1835,N_390,N_467);
xnor U1836 (N_1836,N_800,N_1160);
and U1837 (N_1837,N_1415,N_670);
or U1838 (N_1838,N_1306,N_424);
or U1839 (N_1839,N_1276,N_47);
nand U1840 (N_1840,N_347,N_1043);
nor U1841 (N_1841,N_184,N_760);
xnor U1842 (N_1842,N_1347,N_929);
xnor U1843 (N_1843,N_1145,N_931);
or U1844 (N_1844,N_294,N_587);
nor U1845 (N_1845,N_686,N_892);
nor U1846 (N_1846,N_619,N_468);
or U1847 (N_1847,N_786,N_222);
xnor U1848 (N_1848,N_168,N_37);
and U1849 (N_1849,N_1480,N_1184);
and U1850 (N_1850,N_192,N_140);
xor U1851 (N_1851,N_932,N_41);
or U1852 (N_1852,N_921,N_1381);
nor U1853 (N_1853,N_717,N_421);
and U1854 (N_1854,N_100,N_32);
and U1855 (N_1855,N_387,N_1053);
or U1856 (N_1856,N_935,N_801);
and U1857 (N_1857,N_1183,N_146);
and U1858 (N_1858,N_862,N_386);
and U1859 (N_1859,N_101,N_193);
xnor U1860 (N_1860,N_1172,N_1202);
nor U1861 (N_1861,N_1199,N_1104);
or U1862 (N_1862,N_1189,N_202);
and U1863 (N_1863,N_1422,N_29);
nand U1864 (N_1864,N_367,N_210);
xnor U1865 (N_1865,N_755,N_14);
nand U1866 (N_1866,N_758,N_1495);
nand U1867 (N_1867,N_1181,N_1260);
nor U1868 (N_1868,N_849,N_473);
xnor U1869 (N_1869,N_708,N_27);
and U1870 (N_1870,N_1453,N_448);
or U1871 (N_1871,N_615,N_172);
nand U1872 (N_1872,N_238,N_968);
nor U1873 (N_1873,N_783,N_499);
nand U1874 (N_1874,N_970,N_293);
nor U1875 (N_1875,N_413,N_507);
and U1876 (N_1876,N_805,N_807);
nor U1877 (N_1877,N_631,N_1107);
or U1878 (N_1878,N_551,N_1231);
nor U1879 (N_1879,N_916,N_1410);
xnor U1880 (N_1880,N_1139,N_811);
or U1881 (N_1881,N_1488,N_756);
or U1882 (N_1882,N_1009,N_739);
and U1883 (N_1883,N_459,N_486);
nand U1884 (N_1884,N_848,N_1334);
and U1885 (N_1885,N_127,N_1359);
nand U1886 (N_1886,N_92,N_724);
nor U1887 (N_1887,N_23,N_1428);
nand U1888 (N_1888,N_30,N_1314);
xnor U1889 (N_1889,N_886,N_847);
or U1890 (N_1890,N_998,N_383);
and U1891 (N_1891,N_38,N_1251);
nor U1892 (N_1892,N_1281,N_1211);
nor U1893 (N_1893,N_1293,N_354);
nor U1894 (N_1894,N_1399,N_333);
and U1895 (N_1895,N_317,N_1033);
nand U1896 (N_1896,N_1496,N_548);
or U1897 (N_1897,N_337,N_1079);
nor U1898 (N_1898,N_728,N_1364);
and U1899 (N_1899,N_245,N_69);
and U1900 (N_1900,N_371,N_633);
and U1901 (N_1901,N_400,N_812);
or U1902 (N_1902,N_102,N_613);
nand U1903 (N_1903,N_98,N_1065);
nor U1904 (N_1904,N_1085,N_360);
xor U1905 (N_1905,N_817,N_1164);
and U1906 (N_1906,N_721,N_258);
nor U1907 (N_1907,N_745,N_532);
xor U1908 (N_1908,N_1120,N_1252);
nor U1909 (N_1909,N_689,N_476);
nand U1910 (N_1910,N_1210,N_518);
and U1911 (N_1911,N_1438,N_204);
nor U1912 (N_1912,N_53,N_593);
nand U1913 (N_1913,N_618,N_433);
and U1914 (N_1914,N_160,N_326);
nor U1915 (N_1915,N_458,N_108);
nand U1916 (N_1916,N_540,N_1030);
or U1917 (N_1917,N_1241,N_1378);
nor U1918 (N_1918,N_881,N_1456);
nor U1919 (N_1919,N_497,N_533);
nor U1920 (N_1920,N_1254,N_1418);
and U1921 (N_1921,N_1344,N_520);
and U1922 (N_1922,N_1096,N_469);
nand U1923 (N_1923,N_804,N_596);
nor U1924 (N_1924,N_1023,N_1176);
nand U1925 (N_1925,N_1447,N_625);
or U1926 (N_1926,N_639,N_555);
nand U1927 (N_1927,N_1179,N_45);
or U1928 (N_1928,N_1494,N_1191);
nor U1929 (N_1929,N_1109,N_585);
and U1930 (N_1930,N_732,N_1343);
nor U1931 (N_1931,N_597,N_667);
nor U1932 (N_1932,N_722,N_303);
nor U1933 (N_1933,N_179,N_231);
and U1934 (N_1934,N_503,N_1220);
nor U1935 (N_1935,N_1312,N_981);
or U1936 (N_1936,N_1291,N_1203);
and U1937 (N_1937,N_1299,N_531);
and U1938 (N_1938,N_292,N_617);
nand U1939 (N_1939,N_605,N_510);
nand U1940 (N_1940,N_620,N_1024);
nor U1941 (N_1941,N_516,N_1262);
xor U1942 (N_1942,N_1018,N_1482);
nand U1943 (N_1943,N_1228,N_1213);
xor U1944 (N_1944,N_449,N_1000);
nand U1945 (N_1945,N_787,N_276);
nand U1946 (N_1946,N_1297,N_870);
nor U1947 (N_1947,N_734,N_268);
nand U1948 (N_1948,N_1416,N_1170);
nor U1949 (N_1949,N_832,N_925);
nand U1950 (N_1950,N_1012,N_950);
xor U1951 (N_1951,N_13,N_170);
and U1952 (N_1952,N_978,N_509);
xnor U1953 (N_1953,N_942,N_1404);
and U1954 (N_1954,N_1320,N_799);
and U1955 (N_1955,N_695,N_898);
nand U1956 (N_1956,N_128,N_1355);
xor U1957 (N_1957,N_775,N_979);
xnor U1958 (N_1958,N_877,N_1250);
nor U1959 (N_1959,N_119,N_692);
xor U1960 (N_1960,N_63,N_539);
or U1961 (N_1961,N_665,N_19);
or U1962 (N_1962,N_723,N_362);
nor U1963 (N_1963,N_825,N_521);
nor U1964 (N_1964,N_976,N_850);
nor U1965 (N_1965,N_1218,N_495);
nor U1966 (N_1966,N_11,N_259);
nand U1967 (N_1967,N_629,N_288);
xor U1968 (N_1968,N_1331,N_938);
or U1969 (N_1969,N_1069,N_543);
nand U1970 (N_1970,N_910,N_1084);
nor U1971 (N_1971,N_116,N_917);
or U1972 (N_1972,N_95,N_1215);
and U1973 (N_1973,N_934,N_795);
xnor U1974 (N_1974,N_684,N_173);
nor U1975 (N_1975,N_735,N_820);
and U1976 (N_1976,N_940,N_110);
and U1977 (N_1977,N_791,N_913);
nand U1978 (N_1978,N_475,N_249);
xnor U1979 (N_1979,N_681,N_964);
or U1980 (N_1980,N_142,N_310);
xnor U1981 (N_1981,N_1284,N_813);
nor U1982 (N_1982,N_890,N_479);
and U1983 (N_1983,N_933,N_300);
xor U1984 (N_1984,N_244,N_704);
or U1985 (N_1985,N_553,N_338);
nor U1986 (N_1986,N_563,N_1132);
or U1987 (N_1987,N_1093,N_810);
or U1988 (N_1988,N_608,N_162);
nor U1989 (N_1989,N_993,N_82);
nor U1990 (N_1990,N_3,N_1498);
or U1991 (N_1991,N_43,N_1001);
nor U1992 (N_1992,N_481,N_766);
and U1993 (N_1993,N_679,N_762);
and U1994 (N_1994,N_212,N_1091);
and U1995 (N_1995,N_868,N_763);
xnor U1996 (N_1996,N_175,N_1067);
nand U1997 (N_1997,N_295,N_331);
and U1998 (N_1998,N_611,N_764);
or U1999 (N_1999,N_997,N_180);
and U2000 (N_2000,N_1162,N_1360);
nand U2001 (N_2001,N_643,N_287);
nand U2002 (N_2002,N_1072,N_1255);
nor U2003 (N_2003,N_675,N_777);
or U2004 (N_2004,N_1092,N_358);
and U2005 (N_2005,N_1426,N_1328);
nor U2006 (N_2006,N_867,N_144);
xor U2007 (N_2007,N_1315,N_124);
nand U2008 (N_2008,N_477,N_649);
nand U2009 (N_2009,N_261,N_1124);
or U2010 (N_2010,N_145,N_1345);
nand U2011 (N_2011,N_334,N_235);
xor U2012 (N_2012,N_1377,N_982);
and U2013 (N_2013,N_1153,N_839);
xnor U2014 (N_2014,N_1159,N_1451);
nand U2015 (N_2015,N_461,N_731);
or U2016 (N_2016,N_158,N_462);
xnor U2017 (N_2017,N_250,N_402);
nor U2018 (N_2018,N_490,N_1212);
or U2019 (N_2019,N_1055,N_216);
nor U2020 (N_2020,N_1319,N_214);
or U2021 (N_2021,N_911,N_1077);
xnor U2022 (N_2022,N_148,N_1379);
or U2023 (N_2023,N_1481,N_417);
nand U2024 (N_2024,N_1102,N_1454);
nor U2025 (N_2025,N_1035,N_1131);
nor U2026 (N_2026,N_1300,N_602);
nor U2027 (N_2027,N_1178,N_833);
or U2028 (N_2028,N_513,N_488);
and U2029 (N_2029,N_237,N_1182);
nor U2030 (N_2030,N_430,N_780);
xnor U2031 (N_2031,N_154,N_859);
nor U2032 (N_2032,N_391,N_550);
nor U2033 (N_2033,N_1436,N_752);
xor U2034 (N_2034,N_1074,N_1425);
xnor U2035 (N_2035,N_863,N_883);
and U2036 (N_2036,N_315,N_827);
nand U2037 (N_2037,N_1444,N_1002);
xor U2038 (N_2038,N_1419,N_1007);
or U2039 (N_2039,N_547,N_483);
or U2040 (N_2040,N_105,N_1081);
nand U2041 (N_2041,N_1034,N_1490);
nand U2042 (N_2042,N_389,N_453);
xor U2043 (N_2043,N_844,N_557);
xor U2044 (N_2044,N_1090,N_842);
and U2045 (N_2045,N_872,N_1082);
or U2046 (N_2046,N_1468,N_478);
or U2047 (N_2047,N_1165,N_951);
and U2048 (N_2048,N_736,N_846);
nand U2049 (N_2049,N_189,N_1386);
xnor U2050 (N_2050,N_40,N_990);
nor U2051 (N_2051,N_39,N_664);
nand U2052 (N_2052,N_1028,N_882);
xor U2053 (N_2053,N_296,N_676);
nor U2054 (N_2054,N_363,N_1017);
and U2055 (N_2055,N_1141,N_1308);
nor U2056 (N_2056,N_718,N_1269);
nand U2057 (N_2057,N_1455,N_1037);
or U2058 (N_2058,N_1041,N_944);
nand U2059 (N_2059,N_668,N_1484);
or U2060 (N_2060,N_22,N_275);
and U2061 (N_2061,N_316,N_64);
nand U2062 (N_2062,N_1373,N_880);
and U2063 (N_2063,N_959,N_706);
nand U2064 (N_2064,N_797,N_379);
and U2065 (N_2065,N_1289,N_71);
nand U2066 (N_2066,N_937,N_802);
nand U2067 (N_2067,N_856,N_1349);
nand U2068 (N_2068,N_554,N_1489);
nand U2069 (N_2069,N_66,N_1290);
nor U2070 (N_2070,N_601,N_714);
xnor U2071 (N_2071,N_1134,N_556);
nand U2072 (N_2072,N_366,N_282);
nand U2073 (N_2073,N_523,N_781);
nor U2074 (N_2074,N_983,N_442);
or U2075 (N_2075,N_1240,N_1358);
and U2076 (N_2076,N_682,N_1406);
xnor U2077 (N_2077,N_329,N_67);
xor U2078 (N_2078,N_1098,N_121);
nor U2079 (N_2079,N_971,N_729);
or U2080 (N_2080,N_208,N_586);
nand U2081 (N_2081,N_138,N_1362);
or U2082 (N_2082,N_1052,N_1232);
xnor U2083 (N_2083,N_1086,N_1393);
or U2084 (N_2084,N_741,N_348);
nor U2085 (N_2085,N_1446,N_15);
nor U2086 (N_2086,N_1039,N_213);
and U2087 (N_2087,N_678,N_1236);
or U2088 (N_2088,N_519,N_719);
nand U2089 (N_2089,N_506,N_660);
nor U2090 (N_2090,N_456,N_1303);
xor U2091 (N_2091,N_290,N_155);
xnor U2092 (N_2092,N_655,N_299);
nor U2093 (N_2093,N_1087,N_1195);
or U2094 (N_2094,N_54,N_923);
or U2095 (N_2095,N_768,N_1025);
xor U2096 (N_2096,N_1433,N_325);
nand U2097 (N_2097,N_1367,N_698);
xor U2098 (N_2098,N_995,N_1478);
xor U2099 (N_2099,N_368,N_1427);
xnor U2100 (N_2100,N_5,N_17);
xnor U2101 (N_2101,N_1201,N_1461);
nor U2102 (N_2102,N_446,N_737);
nor U2103 (N_2103,N_1413,N_1019);
nor U2104 (N_2104,N_1487,N_474);
nand U2105 (N_2105,N_1431,N_274);
nor U2106 (N_2106,N_1122,N_996);
nand U2107 (N_2107,N_217,N_1402);
xnor U2108 (N_2108,N_594,N_1151);
nor U2109 (N_2109,N_321,N_709);
or U2110 (N_2110,N_1097,N_335);
and U2111 (N_2111,N_973,N_1088);
or U2112 (N_2112,N_652,N_1288);
and U2113 (N_2113,N_302,N_470);
nor U2114 (N_2114,N_907,N_289);
and U2115 (N_2115,N_1038,N_255);
nor U2116 (N_2116,N_420,N_663);
and U2117 (N_2117,N_1356,N_416);
or U2118 (N_2118,N_1485,N_88);
nor U2119 (N_2119,N_429,N_612);
and U2120 (N_2120,N_241,N_361);
and U2121 (N_2121,N_426,N_195);
or U2122 (N_2122,N_1363,N_1434);
nand U2123 (N_2123,N_1348,N_930);
nor U2124 (N_2124,N_169,N_1473);
nor U2125 (N_2125,N_1214,N_823);
nand U2126 (N_2126,N_1471,N_1094);
or U2127 (N_2127,N_952,N_1318);
nor U2128 (N_2128,N_897,N_584);
or U2129 (N_2129,N_263,N_236);
and U2130 (N_2130,N_1063,N_452);
and U2131 (N_2131,N_1435,N_77);
nor U2132 (N_2132,N_376,N_49);
or U2133 (N_2133,N_432,N_505);
nor U2134 (N_2134,N_1080,N_751);
nand U2135 (N_2135,N_524,N_339);
and U2136 (N_2136,N_8,N_1420);
or U2137 (N_2137,N_558,N_57);
xor U2138 (N_2138,N_504,N_1440);
nand U2139 (N_2139,N_1400,N_1457);
nand U2140 (N_2140,N_1277,N_60);
nor U2141 (N_2141,N_233,N_1206);
or U2142 (N_2142,N_956,N_91);
and U2143 (N_2143,N_1283,N_900);
xnor U2144 (N_2144,N_647,N_345);
or U2145 (N_2145,N_621,N_422);
or U2146 (N_2146,N_957,N_226);
and U2147 (N_2147,N_10,N_1029);
or U2148 (N_2148,N_1066,N_962);
xnor U2149 (N_2149,N_566,N_107);
and U2150 (N_2150,N_715,N_966);
nand U2151 (N_2151,N_642,N_20);
or U2152 (N_2152,N_784,N_418);
and U2153 (N_2153,N_151,N_1258);
nor U2154 (N_2154,N_1138,N_1259);
xnor U2155 (N_2155,N_44,N_324);
and U2156 (N_2156,N_485,N_713);
nand U2157 (N_2157,N_1464,N_1268);
xor U2158 (N_2158,N_1248,N_1114);
nand U2159 (N_2159,N_778,N_707);
xnor U2160 (N_2160,N_669,N_152);
nand U2161 (N_2161,N_445,N_484);
xor U2162 (N_2162,N_1204,N_538);
nand U2163 (N_2163,N_711,N_375);
or U2164 (N_2164,N_201,N_369);
xnor U2165 (N_2165,N_702,N_340);
and U2166 (N_2166,N_749,N_866);
nor U2167 (N_2167,N_798,N_782);
nand U2168 (N_2168,N_385,N_73);
or U2169 (N_2169,N_592,N_1492);
nand U2170 (N_2170,N_1111,N_1227);
xor U2171 (N_2171,N_31,N_1474);
or U2172 (N_2172,N_1135,N_980);
xnor U2173 (N_2173,N_104,N_436);
nand U2174 (N_2174,N_529,N_598);
nor U2175 (N_2175,N_281,N_80);
nand U2176 (N_2176,N_511,N_1274);
nor U2177 (N_2177,N_936,N_36);
and U2178 (N_2178,N_150,N_177);
nor U2179 (N_2179,N_131,N_1205);
and U2180 (N_2180,N_207,N_1421);
and U2181 (N_2181,N_744,N_659);
nand U2182 (N_2182,N_1116,N_372);
and U2183 (N_2183,N_1133,N_256);
xor U2184 (N_2184,N_1472,N_991);
nand U2185 (N_2185,N_896,N_693);
nor U2186 (N_2186,N_1278,N_126);
and U2187 (N_2187,N_1142,N_322);
xor U2188 (N_2188,N_327,N_408);
xnor U2189 (N_2189,N_1340,N_246);
and U2190 (N_2190,N_28,N_534);
xor U2191 (N_2191,N_1014,N_1071);
nand U2192 (N_2192,N_425,N_1432);
nand U2193 (N_2193,N_498,N_1275);
and U2194 (N_2194,N_845,N_1337);
xor U2195 (N_2195,N_884,N_1272);
or U2196 (N_2196,N_494,N_653);
nand U2197 (N_2197,N_401,N_273);
or U2198 (N_2198,N_243,N_1230);
nor U2199 (N_2199,N_50,N_949);
nor U2200 (N_2200,N_406,N_220);
nand U2201 (N_2201,N_658,N_1076);
or U2202 (N_2202,N_769,N_614);
nand U2203 (N_2203,N_118,N_994);
or U2204 (N_2204,N_460,N_229);
nor U2205 (N_2205,N_466,N_457);
xor U2206 (N_2206,N_283,N_284);
nand U2207 (N_2207,N_240,N_1333);
or U2208 (N_2208,N_961,N_945);
nand U2209 (N_2209,N_571,N_561);
xor U2210 (N_2210,N_1376,N_865);
xnor U2211 (N_2211,N_117,N_1194);
or U2212 (N_2212,N_1147,N_941);
nor U2213 (N_2213,N_304,N_225);
or U2214 (N_2214,N_265,N_1121);
and U2215 (N_2215,N_1169,N_977);
xnor U2216 (N_2216,N_1003,N_747);
and U2217 (N_2217,N_1493,N_1177);
xnor U2218 (N_2218,N_197,N_1208);
xor U2219 (N_2219,N_831,N_1442);
xor U2220 (N_2220,N_394,N_439);
or U2221 (N_2221,N_1042,N_1246);
and U2222 (N_2222,N_517,N_1060);
nor U2223 (N_2223,N_228,N_525);
or U2224 (N_2224,N_1264,N_1219);
and U2225 (N_2225,N_291,N_581);
and U2226 (N_2226,N_628,N_987);
or U2227 (N_2227,N_607,N_727);
or U2228 (N_2228,N_1196,N_673);
and U2229 (N_2229,N_161,N_1353);
or U2230 (N_2230,N_572,N_761);
and U2231 (N_2231,N_656,N_1361);
or U2232 (N_2232,N_568,N_546);
nor U2233 (N_2233,N_623,N_988);
and U2234 (N_2234,N_183,N_1459);
xor U2235 (N_2235,N_199,N_1322);
nor U2236 (N_2236,N_1407,N_176);
or U2237 (N_2237,N_1180,N_1458);
and U2238 (N_2238,N_1282,N_567);
nand U2239 (N_2239,N_648,N_437);
nor U2240 (N_2240,N_808,N_72);
or U2241 (N_2241,N_955,N_373);
xnor U2242 (N_2242,N_200,N_1405);
and U2243 (N_2243,N_234,N_609);
nand U2244 (N_2244,N_1465,N_924);
nor U2245 (N_2245,N_51,N_359);
or U2246 (N_2246,N_985,N_864);
nor U2247 (N_2247,N_441,N_342);
nor U2248 (N_2248,N_419,N_1316);
nor U2249 (N_2249,N_58,N_730);
nand U2250 (N_2250,N_1059,N_1244);
and U2251 (N_2251,N_1227,N_1404);
and U2252 (N_2252,N_332,N_824);
nor U2253 (N_2253,N_987,N_746);
and U2254 (N_2254,N_1340,N_747);
and U2255 (N_2255,N_465,N_784);
xor U2256 (N_2256,N_649,N_424);
nand U2257 (N_2257,N_874,N_1164);
or U2258 (N_2258,N_821,N_788);
and U2259 (N_2259,N_70,N_651);
nand U2260 (N_2260,N_1021,N_15);
xor U2261 (N_2261,N_485,N_426);
nand U2262 (N_2262,N_732,N_906);
or U2263 (N_2263,N_406,N_1000);
or U2264 (N_2264,N_868,N_798);
xnor U2265 (N_2265,N_226,N_338);
xnor U2266 (N_2266,N_254,N_1313);
nand U2267 (N_2267,N_307,N_134);
nand U2268 (N_2268,N_1326,N_581);
or U2269 (N_2269,N_1425,N_947);
xor U2270 (N_2270,N_1363,N_667);
nor U2271 (N_2271,N_203,N_1407);
xnor U2272 (N_2272,N_572,N_851);
xnor U2273 (N_2273,N_104,N_639);
and U2274 (N_2274,N_760,N_1238);
or U2275 (N_2275,N_142,N_652);
xor U2276 (N_2276,N_34,N_1042);
xor U2277 (N_2277,N_268,N_990);
nor U2278 (N_2278,N_1150,N_916);
or U2279 (N_2279,N_9,N_646);
nand U2280 (N_2280,N_222,N_945);
and U2281 (N_2281,N_417,N_1048);
or U2282 (N_2282,N_166,N_953);
and U2283 (N_2283,N_646,N_127);
xor U2284 (N_2284,N_355,N_34);
and U2285 (N_2285,N_291,N_779);
xnor U2286 (N_2286,N_1338,N_553);
nand U2287 (N_2287,N_1349,N_742);
xnor U2288 (N_2288,N_1301,N_1008);
nor U2289 (N_2289,N_1136,N_674);
and U2290 (N_2290,N_451,N_1223);
xor U2291 (N_2291,N_314,N_823);
nor U2292 (N_2292,N_407,N_1037);
nor U2293 (N_2293,N_1333,N_123);
or U2294 (N_2294,N_1275,N_919);
nand U2295 (N_2295,N_291,N_1138);
nand U2296 (N_2296,N_530,N_306);
and U2297 (N_2297,N_1279,N_346);
xor U2298 (N_2298,N_119,N_589);
and U2299 (N_2299,N_319,N_1257);
and U2300 (N_2300,N_1442,N_1227);
xor U2301 (N_2301,N_1351,N_71);
and U2302 (N_2302,N_1166,N_749);
nor U2303 (N_2303,N_653,N_634);
nor U2304 (N_2304,N_1211,N_1288);
or U2305 (N_2305,N_936,N_323);
nor U2306 (N_2306,N_535,N_1110);
or U2307 (N_2307,N_112,N_1406);
or U2308 (N_2308,N_526,N_39);
xnor U2309 (N_2309,N_835,N_1169);
nand U2310 (N_2310,N_503,N_369);
xor U2311 (N_2311,N_398,N_1115);
and U2312 (N_2312,N_918,N_746);
nor U2313 (N_2313,N_231,N_1406);
xor U2314 (N_2314,N_1028,N_817);
and U2315 (N_2315,N_1291,N_798);
and U2316 (N_2316,N_244,N_781);
nor U2317 (N_2317,N_413,N_387);
and U2318 (N_2318,N_1202,N_184);
and U2319 (N_2319,N_1018,N_423);
nor U2320 (N_2320,N_1245,N_765);
and U2321 (N_2321,N_442,N_500);
and U2322 (N_2322,N_1037,N_546);
nor U2323 (N_2323,N_684,N_1221);
or U2324 (N_2324,N_690,N_559);
or U2325 (N_2325,N_931,N_1068);
xor U2326 (N_2326,N_402,N_1494);
and U2327 (N_2327,N_1038,N_408);
nand U2328 (N_2328,N_142,N_818);
nor U2329 (N_2329,N_190,N_839);
or U2330 (N_2330,N_1388,N_1134);
nand U2331 (N_2331,N_110,N_1375);
nand U2332 (N_2332,N_119,N_1208);
nor U2333 (N_2333,N_86,N_672);
or U2334 (N_2334,N_513,N_212);
xnor U2335 (N_2335,N_17,N_73);
and U2336 (N_2336,N_602,N_695);
nor U2337 (N_2337,N_850,N_275);
nand U2338 (N_2338,N_731,N_246);
nor U2339 (N_2339,N_691,N_62);
and U2340 (N_2340,N_817,N_309);
nor U2341 (N_2341,N_1172,N_617);
nand U2342 (N_2342,N_577,N_525);
xnor U2343 (N_2343,N_161,N_620);
nor U2344 (N_2344,N_1165,N_990);
and U2345 (N_2345,N_1270,N_887);
nor U2346 (N_2346,N_204,N_1302);
nand U2347 (N_2347,N_818,N_1019);
nor U2348 (N_2348,N_159,N_1173);
nand U2349 (N_2349,N_636,N_781);
or U2350 (N_2350,N_278,N_115);
nor U2351 (N_2351,N_419,N_734);
and U2352 (N_2352,N_402,N_852);
xnor U2353 (N_2353,N_1326,N_1255);
xnor U2354 (N_2354,N_1414,N_1231);
or U2355 (N_2355,N_755,N_643);
or U2356 (N_2356,N_134,N_251);
or U2357 (N_2357,N_322,N_634);
or U2358 (N_2358,N_184,N_612);
and U2359 (N_2359,N_316,N_1277);
and U2360 (N_2360,N_474,N_901);
or U2361 (N_2361,N_911,N_1090);
or U2362 (N_2362,N_664,N_1198);
xnor U2363 (N_2363,N_338,N_1425);
or U2364 (N_2364,N_621,N_1259);
and U2365 (N_2365,N_1220,N_369);
xnor U2366 (N_2366,N_1225,N_382);
nand U2367 (N_2367,N_1046,N_1254);
or U2368 (N_2368,N_285,N_607);
and U2369 (N_2369,N_176,N_786);
xor U2370 (N_2370,N_22,N_437);
or U2371 (N_2371,N_33,N_773);
xnor U2372 (N_2372,N_1204,N_145);
or U2373 (N_2373,N_1448,N_214);
or U2374 (N_2374,N_934,N_241);
nor U2375 (N_2375,N_336,N_0);
nand U2376 (N_2376,N_1290,N_1204);
and U2377 (N_2377,N_649,N_332);
or U2378 (N_2378,N_386,N_1394);
nand U2379 (N_2379,N_17,N_598);
or U2380 (N_2380,N_907,N_775);
xor U2381 (N_2381,N_1118,N_627);
or U2382 (N_2382,N_560,N_524);
or U2383 (N_2383,N_267,N_662);
and U2384 (N_2384,N_51,N_376);
and U2385 (N_2385,N_1241,N_44);
nand U2386 (N_2386,N_987,N_645);
xnor U2387 (N_2387,N_1440,N_106);
xnor U2388 (N_2388,N_562,N_324);
xnor U2389 (N_2389,N_1340,N_646);
and U2390 (N_2390,N_888,N_1248);
xor U2391 (N_2391,N_584,N_1397);
and U2392 (N_2392,N_376,N_739);
or U2393 (N_2393,N_579,N_594);
nor U2394 (N_2394,N_944,N_397);
and U2395 (N_2395,N_792,N_173);
nor U2396 (N_2396,N_1,N_1122);
or U2397 (N_2397,N_1344,N_586);
xnor U2398 (N_2398,N_681,N_42);
xor U2399 (N_2399,N_308,N_1156);
nor U2400 (N_2400,N_721,N_632);
nor U2401 (N_2401,N_1333,N_1269);
and U2402 (N_2402,N_734,N_47);
xor U2403 (N_2403,N_781,N_787);
or U2404 (N_2404,N_72,N_616);
xnor U2405 (N_2405,N_1328,N_763);
xor U2406 (N_2406,N_682,N_313);
and U2407 (N_2407,N_38,N_303);
xnor U2408 (N_2408,N_1329,N_773);
or U2409 (N_2409,N_1289,N_917);
nor U2410 (N_2410,N_1317,N_545);
or U2411 (N_2411,N_486,N_876);
nor U2412 (N_2412,N_674,N_898);
nor U2413 (N_2413,N_1196,N_502);
or U2414 (N_2414,N_320,N_979);
and U2415 (N_2415,N_1210,N_775);
and U2416 (N_2416,N_535,N_264);
or U2417 (N_2417,N_20,N_774);
or U2418 (N_2418,N_644,N_1031);
nand U2419 (N_2419,N_847,N_947);
and U2420 (N_2420,N_416,N_1407);
nor U2421 (N_2421,N_691,N_729);
xnor U2422 (N_2422,N_616,N_926);
xor U2423 (N_2423,N_34,N_44);
or U2424 (N_2424,N_510,N_332);
nor U2425 (N_2425,N_181,N_818);
and U2426 (N_2426,N_616,N_338);
or U2427 (N_2427,N_443,N_917);
or U2428 (N_2428,N_623,N_1091);
or U2429 (N_2429,N_428,N_1435);
and U2430 (N_2430,N_1282,N_1239);
and U2431 (N_2431,N_305,N_1254);
nor U2432 (N_2432,N_675,N_1316);
xnor U2433 (N_2433,N_453,N_1386);
nor U2434 (N_2434,N_1389,N_591);
or U2435 (N_2435,N_674,N_234);
xor U2436 (N_2436,N_245,N_7);
or U2437 (N_2437,N_973,N_403);
or U2438 (N_2438,N_1106,N_1214);
or U2439 (N_2439,N_1482,N_159);
or U2440 (N_2440,N_545,N_333);
nand U2441 (N_2441,N_582,N_202);
nand U2442 (N_2442,N_1203,N_921);
or U2443 (N_2443,N_1311,N_1130);
nor U2444 (N_2444,N_1110,N_298);
or U2445 (N_2445,N_1006,N_284);
nor U2446 (N_2446,N_1154,N_1105);
or U2447 (N_2447,N_682,N_367);
nor U2448 (N_2448,N_915,N_1288);
or U2449 (N_2449,N_1237,N_1340);
xor U2450 (N_2450,N_782,N_372);
xor U2451 (N_2451,N_222,N_601);
nand U2452 (N_2452,N_617,N_530);
or U2453 (N_2453,N_1030,N_705);
xor U2454 (N_2454,N_662,N_614);
or U2455 (N_2455,N_1039,N_831);
or U2456 (N_2456,N_1408,N_414);
xor U2457 (N_2457,N_1260,N_94);
xor U2458 (N_2458,N_245,N_599);
or U2459 (N_2459,N_1311,N_303);
and U2460 (N_2460,N_873,N_815);
and U2461 (N_2461,N_712,N_1381);
and U2462 (N_2462,N_461,N_610);
nand U2463 (N_2463,N_557,N_212);
or U2464 (N_2464,N_1291,N_1338);
or U2465 (N_2465,N_1256,N_1141);
and U2466 (N_2466,N_1364,N_1378);
and U2467 (N_2467,N_1386,N_1158);
nand U2468 (N_2468,N_179,N_347);
or U2469 (N_2469,N_594,N_501);
and U2470 (N_2470,N_49,N_461);
or U2471 (N_2471,N_520,N_1395);
nor U2472 (N_2472,N_780,N_1467);
nand U2473 (N_2473,N_1282,N_1305);
or U2474 (N_2474,N_913,N_1335);
xor U2475 (N_2475,N_994,N_488);
nor U2476 (N_2476,N_766,N_1206);
nor U2477 (N_2477,N_327,N_1016);
xor U2478 (N_2478,N_332,N_1386);
nand U2479 (N_2479,N_1184,N_1497);
nand U2480 (N_2480,N_519,N_399);
nor U2481 (N_2481,N_506,N_1199);
or U2482 (N_2482,N_934,N_1412);
nand U2483 (N_2483,N_1216,N_1008);
or U2484 (N_2484,N_980,N_204);
nor U2485 (N_2485,N_1440,N_28);
nor U2486 (N_2486,N_922,N_1224);
and U2487 (N_2487,N_8,N_887);
nand U2488 (N_2488,N_140,N_800);
nor U2489 (N_2489,N_970,N_1007);
nand U2490 (N_2490,N_486,N_240);
and U2491 (N_2491,N_944,N_801);
and U2492 (N_2492,N_72,N_36);
nor U2493 (N_2493,N_736,N_869);
or U2494 (N_2494,N_655,N_1123);
xor U2495 (N_2495,N_644,N_1253);
or U2496 (N_2496,N_133,N_1439);
and U2497 (N_2497,N_939,N_1309);
nand U2498 (N_2498,N_795,N_1393);
nor U2499 (N_2499,N_924,N_632);
nand U2500 (N_2500,N_570,N_572);
nand U2501 (N_2501,N_333,N_821);
nand U2502 (N_2502,N_53,N_218);
nor U2503 (N_2503,N_352,N_771);
or U2504 (N_2504,N_164,N_549);
xnor U2505 (N_2505,N_915,N_922);
nand U2506 (N_2506,N_1046,N_69);
and U2507 (N_2507,N_265,N_96);
and U2508 (N_2508,N_406,N_1405);
or U2509 (N_2509,N_69,N_1037);
and U2510 (N_2510,N_814,N_835);
nor U2511 (N_2511,N_836,N_1204);
and U2512 (N_2512,N_1485,N_281);
xnor U2513 (N_2513,N_162,N_916);
and U2514 (N_2514,N_1069,N_1153);
xor U2515 (N_2515,N_186,N_768);
or U2516 (N_2516,N_771,N_160);
or U2517 (N_2517,N_1432,N_203);
or U2518 (N_2518,N_1049,N_419);
nand U2519 (N_2519,N_461,N_617);
or U2520 (N_2520,N_238,N_464);
and U2521 (N_2521,N_1237,N_454);
nand U2522 (N_2522,N_489,N_418);
xor U2523 (N_2523,N_248,N_878);
nor U2524 (N_2524,N_610,N_459);
or U2525 (N_2525,N_981,N_968);
nor U2526 (N_2526,N_645,N_627);
nor U2527 (N_2527,N_1115,N_791);
or U2528 (N_2528,N_922,N_190);
xor U2529 (N_2529,N_31,N_10);
nor U2530 (N_2530,N_1096,N_173);
and U2531 (N_2531,N_401,N_875);
or U2532 (N_2532,N_759,N_42);
or U2533 (N_2533,N_329,N_259);
or U2534 (N_2534,N_95,N_1320);
nand U2535 (N_2535,N_1099,N_1120);
xor U2536 (N_2536,N_1448,N_855);
xor U2537 (N_2537,N_1292,N_1129);
or U2538 (N_2538,N_625,N_654);
and U2539 (N_2539,N_366,N_1290);
xnor U2540 (N_2540,N_814,N_1291);
or U2541 (N_2541,N_263,N_1225);
nor U2542 (N_2542,N_1246,N_104);
nor U2543 (N_2543,N_793,N_606);
nand U2544 (N_2544,N_1065,N_531);
nand U2545 (N_2545,N_880,N_647);
nand U2546 (N_2546,N_1307,N_1383);
and U2547 (N_2547,N_163,N_276);
nor U2548 (N_2548,N_695,N_248);
xnor U2549 (N_2549,N_1168,N_512);
or U2550 (N_2550,N_659,N_942);
xnor U2551 (N_2551,N_334,N_1264);
nand U2552 (N_2552,N_1132,N_930);
or U2553 (N_2553,N_1187,N_315);
xor U2554 (N_2554,N_1392,N_868);
nor U2555 (N_2555,N_1188,N_949);
or U2556 (N_2556,N_299,N_652);
xor U2557 (N_2557,N_992,N_1114);
or U2558 (N_2558,N_62,N_731);
nor U2559 (N_2559,N_343,N_755);
nor U2560 (N_2560,N_295,N_761);
nand U2561 (N_2561,N_1458,N_27);
or U2562 (N_2562,N_1387,N_1374);
nor U2563 (N_2563,N_257,N_1078);
nor U2564 (N_2564,N_812,N_407);
and U2565 (N_2565,N_273,N_921);
or U2566 (N_2566,N_974,N_1463);
and U2567 (N_2567,N_1373,N_1025);
nor U2568 (N_2568,N_339,N_520);
and U2569 (N_2569,N_246,N_137);
and U2570 (N_2570,N_220,N_1154);
nor U2571 (N_2571,N_650,N_667);
nor U2572 (N_2572,N_1067,N_12);
xor U2573 (N_2573,N_1463,N_478);
nor U2574 (N_2574,N_912,N_1208);
and U2575 (N_2575,N_508,N_131);
nor U2576 (N_2576,N_1150,N_196);
xor U2577 (N_2577,N_1360,N_839);
or U2578 (N_2578,N_606,N_668);
nor U2579 (N_2579,N_1395,N_1304);
or U2580 (N_2580,N_867,N_1471);
nor U2581 (N_2581,N_923,N_168);
or U2582 (N_2582,N_1300,N_418);
xor U2583 (N_2583,N_996,N_1109);
xnor U2584 (N_2584,N_826,N_1463);
or U2585 (N_2585,N_982,N_388);
xnor U2586 (N_2586,N_886,N_1203);
nor U2587 (N_2587,N_835,N_865);
or U2588 (N_2588,N_869,N_423);
nor U2589 (N_2589,N_256,N_747);
nor U2590 (N_2590,N_63,N_922);
or U2591 (N_2591,N_4,N_1325);
and U2592 (N_2592,N_625,N_1264);
nor U2593 (N_2593,N_1071,N_458);
xnor U2594 (N_2594,N_327,N_882);
nand U2595 (N_2595,N_1468,N_1019);
or U2596 (N_2596,N_256,N_746);
xor U2597 (N_2597,N_747,N_577);
xnor U2598 (N_2598,N_1207,N_396);
and U2599 (N_2599,N_619,N_1125);
nand U2600 (N_2600,N_32,N_616);
nor U2601 (N_2601,N_1084,N_5);
nand U2602 (N_2602,N_1068,N_120);
and U2603 (N_2603,N_886,N_722);
nand U2604 (N_2604,N_954,N_772);
nor U2605 (N_2605,N_1020,N_207);
and U2606 (N_2606,N_1313,N_142);
nor U2607 (N_2607,N_433,N_28);
nor U2608 (N_2608,N_649,N_951);
xnor U2609 (N_2609,N_87,N_1470);
xor U2610 (N_2610,N_1373,N_286);
xor U2611 (N_2611,N_471,N_535);
xnor U2612 (N_2612,N_307,N_659);
nor U2613 (N_2613,N_1328,N_647);
nand U2614 (N_2614,N_209,N_885);
nor U2615 (N_2615,N_1244,N_758);
or U2616 (N_2616,N_1304,N_432);
nand U2617 (N_2617,N_1253,N_1465);
and U2618 (N_2618,N_1211,N_405);
xnor U2619 (N_2619,N_789,N_676);
nand U2620 (N_2620,N_876,N_1169);
xor U2621 (N_2621,N_366,N_264);
nor U2622 (N_2622,N_513,N_962);
and U2623 (N_2623,N_678,N_404);
and U2624 (N_2624,N_231,N_1282);
and U2625 (N_2625,N_685,N_762);
xnor U2626 (N_2626,N_288,N_1138);
or U2627 (N_2627,N_780,N_127);
nand U2628 (N_2628,N_609,N_776);
xnor U2629 (N_2629,N_1273,N_21);
nor U2630 (N_2630,N_235,N_932);
or U2631 (N_2631,N_719,N_608);
and U2632 (N_2632,N_1,N_1425);
xnor U2633 (N_2633,N_160,N_1463);
nor U2634 (N_2634,N_513,N_695);
nand U2635 (N_2635,N_64,N_1307);
xor U2636 (N_2636,N_1098,N_520);
xnor U2637 (N_2637,N_519,N_1291);
and U2638 (N_2638,N_375,N_717);
and U2639 (N_2639,N_915,N_1362);
and U2640 (N_2640,N_873,N_1347);
nor U2641 (N_2641,N_967,N_1404);
xor U2642 (N_2642,N_1128,N_1292);
xnor U2643 (N_2643,N_830,N_457);
nand U2644 (N_2644,N_156,N_580);
nand U2645 (N_2645,N_1158,N_1197);
xnor U2646 (N_2646,N_507,N_555);
and U2647 (N_2647,N_109,N_1349);
and U2648 (N_2648,N_244,N_303);
nor U2649 (N_2649,N_86,N_1459);
nor U2650 (N_2650,N_1316,N_1317);
xnor U2651 (N_2651,N_1445,N_375);
xor U2652 (N_2652,N_909,N_290);
nand U2653 (N_2653,N_77,N_148);
nand U2654 (N_2654,N_866,N_1390);
nand U2655 (N_2655,N_1416,N_786);
or U2656 (N_2656,N_178,N_1299);
nor U2657 (N_2657,N_1478,N_444);
and U2658 (N_2658,N_232,N_1446);
and U2659 (N_2659,N_88,N_1179);
xnor U2660 (N_2660,N_664,N_665);
and U2661 (N_2661,N_1348,N_598);
nor U2662 (N_2662,N_859,N_1460);
nor U2663 (N_2663,N_1462,N_581);
or U2664 (N_2664,N_361,N_1178);
and U2665 (N_2665,N_514,N_1282);
nand U2666 (N_2666,N_1174,N_64);
nand U2667 (N_2667,N_753,N_734);
nand U2668 (N_2668,N_583,N_272);
xor U2669 (N_2669,N_775,N_1310);
or U2670 (N_2670,N_1412,N_833);
nand U2671 (N_2671,N_366,N_312);
xnor U2672 (N_2672,N_944,N_1026);
nand U2673 (N_2673,N_74,N_41);
xnor U2674 (N_2674,N_924,N_1212);
nand U2675 (N_2675,N_136,N_1188);
nand U2676 (N_2676,N_1406,N_1465);
and U2677 (N_2677,N_471,N_1109);
and U2678 (N_2678,N_1044,N_350);
nand U2679 (N_2679,N_571,N_250);
nand U2680 (N_2680,N_781,N_989);
and U2681 (N_2681,N_380,N_13);
nand U2682 (N_2682,N_1047,N_706);
or U2683 (N_2683,N_857,N_90);
or U2684 (N_2684,N_1319,N_1091);
nor U2685 (N_2685,N_30,N_291);
xor U2686 (N_2686,N_1093,N_1130);
nor U2687 (N_2687,N_1354,N_759);
nor U2688 (N_2688,N_600,N_640);
nor U2689 (N_2689,N_1213,N_954);
nor U2690 (N_2690,N_1373,N_79);
nor U2691 (N_2691,N_1442,N_210);
nor U2692 (N_2692,N_521,N_1091);
nand U2693 (N_2693,N_591,N_136);
nand U2694 (N_2694,N_689,N_152);
nor U2695 (N_2695,N_716,N_1377);
nor U2696 (N_2696,N_1148,N_760);
nand U2697 (N_2697,N_217,N_841);
xnor U2698 (N_2698,N_1356,N_476);
and U2699 (N_2699,N_58,N_207);
nor U2700 (N_2700,N_713,N_842);
xnor U2701 (N_2701,N_798,N_135);
and U2702 (N_2702,N_740,N_287);
and U2703 (N_2703,N_1317,N_1489);
or U2704 (N_2704,N_678,N_439);
and U2705 (N_2705,N_695,N_1148);
xnor U2706 (N_2706,N_1437,N_1248);
nor U2707 (N_2707,N_923,N_1404);
nor U2708 (N_2708,N_1177,N_1400);
nor U2709 (N_2709,N_1146,N_902);
and U2710 (N_2710,N_1181,N_332);
xnor U2711 (N_2711,N_387,N_629);
or U2712 (N_2712,N_264,N_1453);
nor U2713 (N_2713,N_1374,N_829);
or U2714 (N_2714,N_1345,N_534);
or U2715 (N_2715,N_1189,N_711);
and U2716 (N_2716,N_905,N_478);
and U2717 (N_2717,N_705,N_765);
nor U2718 (N_2718,N_1001,N_960);
nor U2719 (N_2719,N_1403,N_964);
nor U2720 (N_2720,N_445,N_955);
nand U2721 (N_2721,N_1411,N_273);
or U2722 (N_2722,N_1099,N_1382);
and U2723 (N_2723,N_1297,N_1029);
xor U2724 (N_2724,N_1115,N_238);
nand U2725 (N_2725,N_1165,N_944);
nand U2726 (N_2726,N_435,N_1147);
xnor U2727 (N_2727,N_65,N_1354);
nand U2728 (N_2728,N_1002,N_697);
and U2729 (N_2729,N_614,N_504);
nand U2730 (N_2730,N_431,N_248);
nand U2731 (N_2731,N_243,N_473);
or U2732 (N_2732,N_9,N_491);
nor U2733 (N_2733,N_42,N_959);
nor U2734 (N_2734,N_754,N_501);
and U2735 (N_2735,N_1396,N_606);
or U2736 (N_2736,N_117,N_0);
nand U2737 (N_2737,N_838,N_1246);
and U2738 (N_2738,N_1040,N_762);
or U2739 (N_2739,N_1101,N_272);
xor U2740 (N_2740,N_1445,N_1179);
or U2741 (N_2741,N_598,N_1099);
nor U2742 (N_2742,N_90,N_936);
nor U2743 (N_2743,N_784,N_162);
nand U2744 (N_2744,N_1082,N_1323);
and U2745 (N_2745,N_126,N_828);
or U2746 (N_2746,N_1227,N_1413);
nor U2747 (N_2747,N_1445,N_811);
and U2748 (N_2748,N_1062,N_387);
and U2749 (N_2749,N_1233,N_355);
or U2750 (N_2750,N_72,N_712);
or U2751 (N_2751,N_1125,N_1371);
or U2752 (N_2752,N_661,N_890);
or U2753 (N_2753,N_516,N_328);
or U2754 (N_2754,N_1059,N_1274);
nand U2755 (N_2755,N_1303,N_1290);
and U2756 (N_2756,N_702,N_1402);
nor U2757 (N_2757,N_1303,N_1309);
or U2758 (N_2758,N_1436,N_119);
xnor U2759 (N_2759,N_344,N_566);
and U2760 (N_2760,N_1172,N_264);
or U2761 (N_2761,N_1438,N_454);
and U2762 (N_2762,N_1374,N_136);
xnor U2763 (N_2763,N_1447,N_1330);
xor U2764 (N_2764,N_792,N_645);
xnor U2765 (N_2765,N_286,N_527);
xnor U2766 (N_2766,N_1094,N_348);
or U2767 (N_2767,N_869,N_661);
or U2768 (N_2768,N_991,N_215);
or U2769 (N_2769,N_1287,N_1308);
nor U2770 (N_2770,N_1064,N_1423);
xor U2771 (N_2771,N_354,N_955);
xor U2772 (N_2772,N_837,N_971);
xnor U2773 (N_2773,N_990,N_218);
nand U2774 (N_2774,N_887,N_940);
and U2775 (N_2775,N_1179,N_253);
and U2776 (N_2776,N_863,N_106);
and U2777 (N_2777,N_1309,N_191);
or U2778 (N_2778,N_169,N_977);
nand U2779 (N_2779,N_1158,N_79);
nand U2780 (N_2780,N_449,N_479);
or U2781 (N_2781,N_505,N_287);
and U2782 (N_2782,N_663,N_1279);
and U2783 (N_2783,N_1351,N_176);
and U2784 (N_2784,N_950,N_349);
or U2785 (N_2785,N_793,N_707);
and U2786 (N_2786,N_610,N_338);
or U2787 (N_2787,N_1295,N_184);
or U2788 (N_2788,N_348,N_154);
nor U2789 (N_2789,N_529,N_354);
xor U2790 (N_2790,N_48,N_228);
xor U2791 (N_2791,N_1321,N_115);
or U2792 (N_2792,N_174,N_1013);
nor U2793 (N_2793,N_441,N_507);
or U2794 (N_2794,N_257,N_1435);
nand U2795 (N_2795,N_168,N_1127);
or U2796 (N_2796,N_932,N_823);
and U2797 (N_2797,N_244,N_1269);
or U2798 (N_2798,N_1371,N_883);
or U2799 (N_2799,N_127,N_69);
nor U2800 (N_2800,N_837,N_1427);
and U2801 (N_2801,N_587,N_1177);
and U2802 (N_2802,N_824,N_108);
xor U2803 (N_2803,N_76,N_468);
or U2804 (N_2804,N_1193,N_656);
and U2805 (N_2805,N_781,N_832);
nand U2806 (N_2806,N_598,N_809);
nor U2807 (N_2807,N_1332,N_353);
or U2808 (N_2808,N_485,N_207);
xnor U2809 (N_2809,N_1420,N_494);
nand U2810 (N_2810,N_1255,N_604);
nand U2811 (N_2811,N_116,N_297);
and U2812 (N_2812,N_1398,N_1216);
xor U2813 (N_2813,N_699,N_1167);
and U2814 (N_2814,N_506,N_224);
xor U2815 (N_2815,N_24,N_1182);
xnor U2816 (N_2816,N_99,N_1180);
and U2817 (N_2817,N_1027,N_675);
or U2818 (N_2818,N_586,N_499);
or U2819 (N_2819,N_1029,N_1455);
xnor U2820 (N_2820,N_818,N_330);
xor U2821 (N_2821,N_149,N_1222);
nand U2822 (N_2822,N_755,N_1158);
and U2823 (N_2823,N_773,N_9);
nor U2824 (N_2824,N_1127,N_1089);
xnor U2825 (N_2825,N_854,N_1337);
xor U2826 (N_2826,N_483,N_1481);
nand U2827 (N_2827,N_1059,N_258);
and U2828 (N_2828,N_863,N_1133);
and U2829 (N_2829,N_719,N_76);
nor U2830 (N_2830,N_139,N_1076);
nand U2831 (N_2831,N_224,N_1001);
nand U2832 (N_2832,N_862,N_1294);
xor U2833 (N_2833,N_130,N_1097);
xnor U2834 (N_2834,N_979,N_704);
nand U2835 (N_2835,N_1471,N_560);
xor U2836 (N_2836,N_722,N_464);
nor U2837 (N_2837,N_987,N_527);
and U2838 (N_2838,N_1121,N_1367);
xnor U2839 (N_2839,N_407,N_529);
nor U2840 (N_2840,N_1377,N_821);
or U2841 (N_2841,N_48,N_1289);
nor U2842 (N_2842,N_566,N_597);
xnor U2843 (N_2843,N_1438,N_1217);
nor U2844 (N_2844,N_1325,N_896);
nor U2845 (N_2845,N_1276,N_833);
and U2846 (N_2846,N_231,N_1092);
xnor U2847 (N_2847,N_594,N_1350);
and U2848 (N_2848,N_119,N_892);
nor U2849 (N_2849,N_554,N_754);
nor U2850 (N_2850,N_771,N_1470);
xnor U2851 (N_2851,N_615,N_830);
or U2852 (N_2852,N_67,N_361);
and U2853 (N_2853,N_547,N_1160);
or U2854 (N_2854,N_665,N_1247);
nand U2855 (N_2855,N_130,N_121);
nor U2856 (N_2856,N_699,N_369);
nand U2857 (N_2857,N_719,N_1127);
nor U2858 (N_2858,N_287,N_920);
and U2859 (N_2859,N_1064,N_563);
nand U2860 (N_2860,N_275,N_918);
nand U2861 (N_2861,N_858,N_634);
or U2862 (N_2862,N_1491,N_789);
xnor U2863 (N_2863,N_192,N_1173);
xor U2864 (N_2864,N_558,N_853);
or U2865 (N_2865,N_1042,N_740);
xor U2866 (N_2866,N_529,N_1233);
and U2867 (N_2867,N_477,N_1022);
and U2868 (N_2868,N_828,N_1207);
nor U2869 (N_2869,N_1069,N_732);
nand U2870 (N_2870,N_1436,N_32);
and U2871 (N_2871,N_689,N_1211);
nor U2872 (N_2872,N_1026,N_907);
nor U2873 (N_2873,N_1392,N_922);
nand U2874 (N_2874,N_1391,N_743);
and U2875 (N_2875,N_393,N_729);
or U2876 (N_2876,N_443,N_259);
nor U2877 (N_2877,N_203,N_622);
or U2878 (N_2878,N_1412,N_583);
nand U2879 (N_2879,N_793,N_635);
and U2880 (N_2880,N_388,N_280);
nor U2881 (N_2881,N_680,N_1274);
or U2882 (N_2882,N_1204,N_845);
nor U2883 (N_2883,N_984,N_203);
nor U2884 (N_2884,N_1020,N_1241);
nand U2885 (N_2885,N_176,N_1391);
xor U2886 (N_2886,N_262,N_629);
and U2887 (N_2887,N_1197,N_1392);
and U2888 (N_2888,N_62,N_857);
xnor U2889 (N_2889,N_1354,N_273);
nand U2890 (N_2890,N_1477,N_773);
nand U2891 (N_2891,N_376,N_1375);
or U2892 (N_2892,N_159,N_1399);
and U2893 (N_2893,N_953,N_475);
and U2894 (N_2894,N_246,N_325);
nand U2895 (N_2895,N_700,N_586);
or U2896 (N_2896,N_823,N_651);
or U2897 (N_2897,N_103,N_1299);
xnor U2898 (N_2898,N_1140,N_1425);
xnor U2899 (N_2899,N_883,N_46);
and U2900 (N_2900,N_1462,N_883);
nor U2901 (N_2901,N_68,N_82);
and U2902 (N_2902,N_796,N_1370);
xnor U2903 (N_2903,N_1493,N_365);
and U2904 (N_2904,N_1028,N_1094);
or U2905 (N_2905,N_166,N_304);
nand U2906 (N_2906,N_15,N_1243);
nand U2907 (N_2907,N_853,N_896);
or U2908 (N_2908,N_403,N_1157);
nor U2909 (N_2909,N_212,N_659);
nor U2910 (N_2910,N_1117,N_859);
nand U2911 (N_2911,N_589,N_1091);
nor U2912 (N_2912,N_168,N_930);
nand U2913 (N_2913,N_285,N_114);
nor U2914 (N_2914,N_690,N_39);
and U2915 (N_2915,N_443,N_1396);
and U2916 (N_2916,N_1105,N_694);
xor U2917 (N_2917,N_1051,N_1434);
xor U2918 (N_2918,N_1211,N_1086);
and U2919 (N_2919,N_1257,N_312);
or U2920 (N_2920,N_1063,N_199);
or U2921 (N_2921,N_1204,N_1289);
xnor U2922 (N_2922,N_1490,N_332);
or U2923 (N_2923,N_267,N_62);
nand U2924 (N_2924,N_639,N_1079);
nor U2925 (N_2925,N_1253,N_1316);
xnor U2926 (N_2926,N_1215,N_490);
xnor U2927 (N_2927,N_1396,N_162);
nor U2928 (N_2928,N_458,N_1281);
and U2929 (N_2929,N_999,N_1473);
or U2930 (N_2930,N_1287,N_415);
xor U2931 (N_2931,N_166,N_548);
and U2932 (N_2932,N_552,N_382);
and U2933 (N_2933,N_1080,N_896);
and U2934 (N_2934,N_154,N_495);
and U2935 (N_2935,N_1081,N_451);
or U2936 (N_2936,N_1287,N_1167);
or U2937 (N_2937,N_1198,N_945);
nand U2938 (N_2938,N_115,N_401);
xnor U2939 (N_2939,N_162,N_44);
nand U2940 (N_2940,N_268,N_1405);
nor U2941 (N_2941,N_557,N_939);
nor U2942 (N_2942,N_1267,N_1256);
nor U2943 (N_2943,N_1375,N_408);
nor U2944 (N_2944,N_960,N_923);
or U2945 (N_2945,N_81,N_1152);
xnor U2946 (N_2946,N_334,N_909);
nand U2947 (N_2947,N_846,N_1164);
nand U2948 (N_2948,N_772,N_1268);
and U2949 (N_2949,N_177,N_325);
xor U2950 (N_2950,N_292,N_1152);
or U2951 (N_2951,N_528,N_1289);
nor U2952 (N_2952,N_1349,N_1016);
and U2953 (N_2953,N_1424,N_580);
or U2954 (N_2954,N_9,N_1467);
nand U2955 (N_2955,N_765,N_1230);
xor U2956 (N_2956,N_515,N_607);
and U2957 (N_2957,N_423,N_585);
nor U2958 (N_2958,N_1348,N_540);
nand U2959 (N_2959,N_108,N_1498);
and U2960 (N_2960,N_316,N_118);
nor U2961 (N_2961,N_8,N_1239);
nor U2962 (N_2962,N_830,N_453);
nand U2963 (N_2963,N_1000,N_884);
nand U2964 (N_2964,N_213,N_298);
nor U2965 (N_2965,N_1407,N_327);
and U2966 (N_2966,N_1044,N_63);
and U2967 (N_2967,N_141,N_58);
and U2968 (N_2968,N_368,N_277);
nor U2969 (N_2969,N_203,N_125);
nand U2970 (N_2970,N_1448,N_1490);
and U2971 (N_2971,N_1324,N_460);
xor U2972 (N_2972,N_525,N_285);
or U2973 (N_2973,N_24,N_1260);
or U2974 (N_2974,N_283,N_1192);
xnor U2975 (N_2975,N_1401,N_375);
xnor U2976 (N_2976,N_1320,N_1078);
or U2977 (N_2977,N_800,N_1395);
or U2978 (N_2978,N_839,N_921);
nand U2979 (N_2979,N_321,N_429);
nor U2980 (N_2980,N_268,N_1349);
xnor U2981 (N_2981,N_697,N_1398);
nand U2982 (N_2982,N_72,N_432);
nor U2983 (N_2983,N_1295,N_111);
xor U2984 (N_2984,N_715,N_448);
or U2985 (N_2985,N_1300,N_1090);
nor U2986 (N_2986,N_784,N_433);
xor U2987 (N_2987,N_516,N_484);
xor U2988 (N_2988,N_892,N_12);
nand U2989 (N_2989,N_203,N_386);
or U2990 (N_2990,N_1041,N_1449);
and U2991 (N_2991,N_1378,N_1474);
nor U2992 (N_2992,N_879,N_1454);
or U2993 (N_2993,N_341,N_363);
xnor U2994 (N_2994,N_1372,N_353);
xnor U2995 (N_2995,N_1490,N_431);
or U2996 (N_2996,N_1427,N_704);
nor U2997 (N_2997,N_760,N_187);
nand U2998 (N_2998,N_1338,N_651);
or U2999 (N_2999,N_237,N_860);
nand U3000 (N_3000,N_1903,N_2674);
or U3001 (N_3001,N_2549,N_2951);
or U3002 (N_3002,N_2683,N_2160);
xor U3003 (N_3003,N_2917,N_2026);
xnor U3004 (N_3004,N_2841,N_2924);
xor U3005 (N_3005,N_2719,N_2697);
nor U3006 (N_3006,N_2808,N_2000);
nand U3007 (N_3007,N_1879,N_2165);
xor U3008 (N_3008,N_2374,N_2237);
or U3009 (N_3009,N_2042,N_2502);
nand U3010 (N_3010,N_1830,N_2846);
or U3011 (N_3011,N_2937,N_2071);
and U3012 (N_3012,N_2546,N_2747);
nand U3013 (N_3013,N_2359,N_2974);
nand U3014 (N_3014,N_2452,N_1991);
xnor U3015 (N_3015,N_2327,N_2700);
and U3016 (N_3016,N_1718,N_1806);
nor U3017 (N_3017,N_2240,N_2305);
and U3018 (N_3018,N_2550,N_2539);
nor U3019 (N_3019,N_1530,N_2272);
nand U3020 (N_3020,N_1599,N_2439);
nand U3021 (N_3021,N_2140,N_2762);
nor U3022 (N_3022,N_2168,N_2708);
nor U3023 (N_3023,N_2336,N_1663);
xor U3024 (N_3024,N_2832,N_1623);
and U3025 (N_3025,N_2002,N_2801);
or U3026 (N_3026,N_2454,N_1794);
or U3027 (N_3027,N_2433,N_2823);
nand U3028 (N_3028,N_2676,N_2360);
nor U3029 (N_3029,N_1935,N_2909);
nand U3030 (N_3030,N_2227,N_2202);
or U3031 (N_3031,N_1790,N_2877);
or U3032 (N_3032,N_2701,N_2045);
nand U3033 (N_3033,N_2353,N_2512);
and U3034 (N_3034,N_1885,N_2013);
or U3035 (N_3035,N_2334,N_1643);
nor U3036 (N_3036,N_1967,N_1914);
nor U3037 (N_3037,N_2208,N_1977);
nand U3038 (N_3038,N_1818,N_2681);
nor U3039 (N_3039,N_2562,N_2725);
nand U3040 (N_3040,N_2741,N_1943);
xor U3041 (N_3041,N_2092,N_2622);
nor U3042 (N_3042,N_2956,N_2756);
nand U3043 (N_3043,N_1796,N_1963);
and U3044 (N_3044,N_2868,N_2354);
xor U3045 (N_3045,N_1805,N_2185);
or U3046 (N_3046,N_2484,N_2720);
xnor U3047 (N_3047,N_2825,N_1752);
xor U3048 (N_3048,N_2406,N_1844);
xnor U3049 (N_3049,N_2234,N_2568);
or U3050 (N_3050,N_2582,N_2992);
nand U3051 (N_3051,N_2803,N_2356);
or U3052 (N_3052,N_2181,N_2745);
nor U3053 (N_3053,N_2736,N_2890);
nand U3054 (N_3054,N_1831,N_2008);
and U3055 (N_3055,N_1978,N_2540);
xor U3056 (N_3056,N_2754,N_2102);
xnor U3057 (N_3057,N_2211,N_1961);
xor U3058 (N_3058,N_1620,N_2383);
nor U3059 (N_3059,N_2285,N_2450);
or U3060 (N_3060,N_2624,N_1832);
nand U3061 (N_3061,N_2369,N_2282);
nor U3062 (N_3062,N_2579,N_2385);
or U3063 (N_3063,N_1645,N_2099);
nor U3064 (N_3064,N_1930,N_2085);
nor U3065 (N_3065,N_2120,N_2584);
nor U3066 (N_3066,N_2842,N_2270);
and U3067 (N_3067,N_2184,N_2771);
or U3068 (N_3068,N_2203,N_2428);
xor U3069 (N_3069,N_2705,N_2031);
and U3070 (N_3070,N_2942,N_2694);
xnor U3071 (N_3071,N_1749,N_1501);
nand U3072 (N_3072,N_2124,N_2918);
nand U3073 (N_3073,N_2693,N_2769);
and U3074 (N_3074,N_2019,N_2685);
nand U3075 (N_3075,N_2036,N_1803);
or U3076 (N_3076,N_1947,N_2279);
and U3077 (N_3077,N_2254,N_2819);
nor U3078 (N_3078,N_2351,N_2511);
and U3079 (N_3079,N_1675,N_1694);
or U3080 (N_3080,N_2711,N_1756);
and U3081 (N_3081,N_2341,N_2895);
nor U3082 (N_3082,N_2446,N_2938);
nor U3083 (N_3083,N_2695,N_1625);
nor U3084 (N_3084,N_2486,N_2014);
or U3085 (N_3085,N_1804,N_1783);
or U3086 (N_3086,N_2112,N_2405);
and U3087 (N_3087,N_2618,N_2134);
or U3088 (N_3088,N_1709,N_2188);
nand U3089 (N_3089,N_2207,N_2804);
xnor U3090 (N_3090,N_1812,N_2996);
or U3091 (N_3091,N_2717,N_1556);
or U3092 (N_3092,N_2557,N_2827);
or U3093 (N_3093,N_2326,N_2167);
and U3094 (N_3094,N_2407,N_2636);
and U3095 (N_3095,N_2343,N_2492);
xor U3096 (N_3096,N_1521,N_1577);
nor U3097 (N_3097,N_1560,N_1719);
or U3098 (N_3098,N_1737,N_2962);
and U3099 (N_3099,N_1924,N_2419);
nand U3100 (N_3100,N_2422,N_2444);
nand U3101 (N_3101,N_2316,N_2111);
nor U3102 (N_3102,N_1764,N_1542);
nor U3103 (N_3103,N_1692,N_1870);
and U3104 (N_3104,N_2853,N_2905);
nor U3105 (N_3105,N_2344,N_2268);
xor U3106 (N_3106,N_2730,N_2812);
nand U3107 (N_3107,N_2100,N_1955);
nor U3108 (N_3108,N_2798,N_1860);
and U3109 (N_3109,N_2623,N_2236);
nand U3110 (N_3110,N_1527,N_2792);
and U3111 (N_3111,N_2474,N_2109);
and U3112 (N_3112,N_2456,N_1894);
nor U3113 (N_3113,N_2090,N_1544);
or U3114 (N_3114,N_2716,N_1595);
nand U3115 (N_3115,N_2519,N_2367);
nor U3116 (N_3116,N_2654,N_2097);
nand U3117 (N_3117,N_2314,N_2573);
nor U3118 (N_3118,N_2094,N_2066);
nand U3119 (N_3119,N_1918,N_2640);
and U3120 (N_3120,N_2509,N_1738);
or U3121 (N_3121,N_2258,N_2157);
xnor U3122 (N_3122,N_2763,N_2912);
nor U3123 (N_3123,N_2605,N_1964);
and U3124 (N_3124,N_1950,N_1644);
xor U3125 (N_3125,N_1791,N_2488);
xnor U3126 (N_3126,N_1518,N_1992);
and U3127 (N_3127,N_1863,N_1546);
xor U3128 (N_3128,N_2914,N_2321);
or U3129 (N_3129,N_2675,N_1776);
nor U3130 (N_3130,N_2269,N_1656);
xor U3131 (N_3131,N_2513,N_1584);
or U3132 (N_3132,N_1529,N_1676);
xor U3133 (N_3133,N_1899,N_1814);
nand U3134 (N_3134,N_2328,N_1858);
or U3135 (N_3135,N_2280,N_2752);
xor U3136 (N_3136,N_2121,N_2993);
and U3137 (N_3137,N_2323,N_2648);
and U3138 (N_3138,N_2872,N_2978);
xnor U3139 (N_3139,N_1611,N_2011);
and U3140 (N_3140,N_2880,N_2964);
xnor U3141 (N_3141,N_2970,N_2119);
xnor U3142 (N_3142,N_1695,N_2527);
or U3143 (N_3143,N_2617,N_2921);
and U3144 (N_3144,N_2899,N_2789);
nor U3145 (N_3145,N_1538,N_2418);
xnor U3146 (N_3146,N_2434,N_2136);
nor U3147 (N_3147,N_2516,N_2785);
xor U3148 (N_3148,N_2806,N_2751);
or U3149 (N_3149,N_2592,N_1979);
and U3150 (N_3150,N_2940,N_1777);
xnor U3151 (N_3151,N_2571,N_1626);
xor U3152 (N_3152,N_1674,N_2186);
nand U3153 (N_3153,N_1822,N_2977);
nor U3154 (N_3154,N_1678,N_2818);
or U3155 (N_3155,N_1745,N_2295);
nor U3156 (N_3156,N_1868,N_1946);
nor U3157 (N_3157,N_1988,N_1531);
or U3158 (N_3158,N_1802,N_2440);
nor U3159 (N_3159,N_2273,N_2765);
xnor U3160 (N_3160,N_1664,N_1909);
and U3161 (N_3161,N_2477,N_1951);
nand U3162 (N_3162,N_1701,N_2548);
or U3163 (N_3163,N_2309,N_2891);
or U3164 (N_3164,N_2146,N_2906);
or U3165 (N_3165,N_1565,N_2863);
nand U3166 (N_3166,N_2835,N_1853);
and U3167 (N_3167,N_1843,N_2426);
or U3168 (N_3168,N_2349,N_1601);
and U3169 (N_3169,N_2703,N_1887);
nand U3170 (N_3170,N_2122,N_1683);
nand U3171 (N_3171,N_2784,N_1665);
or U3172 (N_3172,N_2535,N_2723);
and U3173 (N_3173,N_2649,N_2222);
nand U3174 (N_3174,N_2224,N_2001);
xor U3175 (N_3175,N_2151,N_2850);
xnor U3176 (N_3176,N_1705,N_2604);
nor U3177 (N_3177,N_2370,N_2786);
xnor U3178 (N_3178,N_1974,N_2517);
or U3179 (N_3179,N_2294,N_2365);
nor U3180 (N_3180,N_1691,N_2619);
xnor U3181 (N_3181,N_2245,N_2402);
or U3182 (N_3182,N_2417,N_1847);
nand U3183 (N_3183,N_2554,N_1715);
or U3184 (N_3184,N_2503,N_2041);
nor U3185 (N_3185,N_2047,N_2834);
nand U3186 (N_3186,N_2318,N_2973);
xor U3187 (N_3187,N_2052,N_2174);
xnor U3188 (N_3188,N_2278,N_1765);
nor U3189 (N_3189,N_1881,N_2997);
nor U3190 (N_3190,N_2555,N_2209);
nand U3191 (N_3191,N_2559,N_2838);
and U3192 (N_3192,N_1669,N_1566);
and U3193 (N_3193,N_2199,N_2101);
xnor U3194 (N_3194,N_1913,N_2657);
or U3195 (N_3195,N_2936,N_2733);
nand U3196 (N_3196,N_1567,N_2189);
or U3197 (N_3197,N_2757,N_1515);
xnor U3198 (N_3198,N_1516,N_2532);
and U3199 (N_3199,N_2311,N_2560);
nand U3200 (N_3200,N_2088,N_1539);
and U3201 (N_3201,N_2277,N_2178);
nor U3202 (N_3202,N_1986,N_1704);
or U3203 (N_3203,N_2907,N_1864);
xnor U3204 (N_3204,N_2217,N_2156);
nor U3205 (N_3205,N_2459,N_2116);
nand U3206 (N_3206,N_1976,N_1722);
xor U3207 (N_3207,N_2462,N_2073);
and U3208 (N_3208,N_2855,N_2647);
and U3209 (N_3209,N_2445,N_2129);
nor U3210 (N_3210,N_1829,N_1528);
and U3211 (N_3211,N_2781,N_2040);
nand U3212 (N_3212,N_2656,N_2998);
and U3213 (N_3213,N_2761,N_1936);
or U3214 (N_3214,N_2377,N_2286);
nor U3215 (N_3215,N_2276,N_1609);
xor U3216 (N_3216,N_1801,N_2195);
or U3217 (N_3217,N_2176,N_2558);
or U3218 (N_3218,N_2871,N_1892);
or U3219 (N_3219,N_1916,N_1736);
nand U3220 (N_3220,N_2991,N_2496);
nor U3221 (N_3221,N_2794,N_2642);
nand U3222 (N_3222,N_1740,N_2251);
xnor U3223 (N_3223,N_2672,N_1898);
and U3224 (N_3224,N_2123,N_2275);
xor U3225 (N_3225,N_1834,N_1712);
xnor U3226 (N_3226,N_1622,N_2304);
and U3227 (N_3227,N_2067,N_2489);
xor U3228 (N_3228,N_2479,N_2255);
nand U3229 (N_3229,N_2577,N_2429);
nor U3230 (N_3230,N_2319,N_2056);
xor U3231 (N_3231,N_2373,N_2536);
xnor U3232 (N_3232,N_2587,N_1593);
xnor U3233 (N_3233,N_2722,N_2204);
or U3234 (N_3234,N_2080,N_2091);
xor U3235 (N_3235,N_2879,N_2687);
and U3236 (N_3236,N_2264,N_2634);
and U3237 (N_3237,N_1773,N_2778);
or U3238 (N_3238,N_2357,N_1841);
nor U3239 (N_3239,N_2455,N_1727);
nor U3240 (N_3240,N_2159,N_1820);
nand U3241 (N_3241,N_2468,N_2791);
and U3242 (N_3242,N_2148,N_1957);
nand U3243 (N_3243,N_2413,N_1867);
nor U3244 (N_3244,N_2049,N_2117);
nor U3245 (N_3245,N_1633,N_2198);
or U3246 (N_3246,N_1915,N_2797);
nand U3247 (N_3247,N_2478,N_2876);
and U3248 (N_3248,N_1763,N_2408);
xor U3249 (N_3249,N_2632,N_1502);
and U3250 (N_3250,N_1579,N_2796);
xnor U3251 (N_3251,N_2215,N_2155);
xnor U3252 (N_3252,N_1690,N_2788);
nor U3253 (N_3253,N_2313,N_1775);
xor U3254 (N_3254,N_2415,N_2126);
and U3255 (N_3255,N_1762,N_1889);
xor U3256 (N_3256,N_1563,N_1716);
nand U3257 (N_3257,N_2875,N_2830);
nor U3258 (N_3258,N_2025,N_1636);
nand U3259 (N_3259,N_1781,N_2263);
or U3260 (N_3260,N_1734,N_1607);
nand U3261 (N_3261,N_1631,N_2127);
nand U3262 (N_3262,N_2988,N_2661);
nand U3263 (N_3263,N_2696,N_2340);
nand U3264 (N_3264,N_2563,N_2985);
xor U3265 (N_3265,N_2086,N_1994);
xor U3266 (N_3266,N_2130,N_2153);
nor U3267 (N_3267,N_1869,N_1862);
nor U3268 (N_3268,N_2448,N_2543);
nand U3269 (N_3269,N_1982,N_2424);
or U3270 (N_3270,N_2020,N_1861);
and U3271 (N_3271,N_2487,N_1846);
and U3272 (N_3272,N_2615,N_2060);
and U3273 (N_3273,N_1667,N_1504);
or U3274 (N_3274,N_2465,N_2154);
nand U3275 (N_3275,N_2024,N_2403);
or U3276 (N_3276,N_1652,N_2858);
xnor U3277 (N_3277,N_2082,N_2766);
nor U3278 (N_3278,N_2986,N_1925);
nand U3279 (N_3279,N_1826,N_2320);
xor U3280 (N_3280,N_2069,N_2449);
and U3281 (N_3281,N_1699,N_1984);
and U3282 (N_3282,N_1702,N_2903);
or U3283 (N_3283,N_2095,N_1912);
and U3284 (N_3284,N_1904,N_1707);
xor U3285 (N_3285,N_2980,N_2057);
or U3286 (N_3286,N_2175,N_2888);
or U3287 (N_3287,N_1987,N_1875);
or U3288 (N_3288,N_1621,N_1807);
and U3289 (N_3289,N_2421,N_2162);
or U3290 (N_3290,N_2999,N_2274);
or U3291 (N_3291,N_2125,N_1996);
and U3292 (N_3292,N_2829,N_1714);
or U3293 (N_3293,N_1989,N_2528);
and U3294 (N_3294,N_1677,N_2171);
and U3295 (N_3295,N_2570,N_2566);
nor U3296 (N_3296,N_2494,N_1604);
or U3297 (N_3297,N_1723,N_1911);
or U3298 (N_3298,N_1758,N_2288);
nor U3299 (N_3299,N_1828,N_1548);
xnor U3300 (N_3300,N_2296,N_2522);
xnor U3301 (N_3301,N_2633,N_2746);
or U3302 (N_3302,N_2959,N_2594);
nor U3303 (N_3303,N_1732,N_2149);
nand U3304 (N_3304,N_1559,N_2641);
or U3305 (N_3305,N_1578,N_1617);
or U3306 (N_3306,N_1835,N_2501);
xnor U3307 (N_3307,N_2271,N_1642);
or U3308 (N_3308,N_2810,N_2505);
or U3309 (N_3309,N_2894,N_2076);
or U3310 (N_3310,N_2645,N_2910);
and U3311 (N_3311,N_2346,N_1784);
or U3312 (N_3312,N_2820,N_2362);
nand U3313 (N_3313,N_2737,N_2187);
or U3314 (N_3314,N_2780,N_2643);
nor U3315 (N_3315,N_2046,N_1511);
and U3316 (N_3316,N_1685,N_2911);
nand U3317 (N_3317,N_1517,N_2103);
or U3318 (N_3318,N_2231,N_1576);
xor U3319 (N_3319,N_1618,N_2960);
nand U3320 (N_3320,N_1825,N_2581);
nand U3321 (N_3321,N_2933,N_2824);
nand U3322 (N_3322,N_2228,N_2994);
nand U3323 (N_3323,N_2646,N_1995);
and U3324 (N_3324,N_1670,N_1613);
nand U3325 (N_3325,N_1837,N_1587);
nand U3326 (N_3326,N_2347,N_2979);
and U3327 (N_3327,N_1968,N_2726);
or U3328 (N_3328,N_1811,N_1526);
or U3329 (N_3329,N_2603,N_2787);
and U3330 (N_3330,N_1923,N_2690);
or U3331 (N_3331,N_1603,N_2238);
nand U3332 (N_3332,N_1505,N_2811);
nand U3333 (N_3333,N_2902,N_2668);
nand U3334 (N_3334,N_1981,N_1612);
nor U3335 (N_3335,N_1574,N_2691);
nand U3336 (N_3336,N_1759,N_1886);
and U3337 (N_3337,N_2401,N_2293);
xor U3338 (N_3338,N_1922,N_1525);
nor U3339 (N_3339,N_1827,N_2729);
nand U3340 (N_3340,N_1572,N_1509);
or U3341 (N_3341,N_2982,N_1666);
nor U3342 (N_3342,N_1896,N_2375);
and U3343 (N_3343,N_2414,N_1966);
and U3344 (N_3344,N_1954,N_2205);
nand U3345 (N_3345,N_2950,N_2790);
nor U3346 (N_3346,N_2467,N_1660);
and U3347 (N_3347,N_2177,N_1639);
or U3348 (N_3348,N_2699,N_2389);
xnor U3349 (N_3349,N_2283,N_1541);
nor U3350 (N_3350,N_1972,N_2055);
nor U3351 (N_3351,N_2915,N_2995);
xnor U3352 (N_3352,N_2965,N_1503);
xor U3353 (N_3353,N_2302,N_2614);
nor U3354 (N_3354,N_2022,N_1931);
xnor U3355 (N_3355,N_1562,N_2172);
nand U3356 (N_3356,N_1686,N_2009);
xor U3357 (N_3357,N_2541,N_1747);
nor U3358 (N_3358,N_2299,N_2971);
and U3359 (N_3359,N_1932,N_1585);
and U3360 (N_3360,N_2411,N_2957);
and U3361 (N_3361,N_2431,N_2702);
and U3362 (N_3362,N_2164,N_2934);
and U3363 (N_3363,N_1921,N_2706);
and U3364 (N_3364,N_2926,N_2601);
nand U3365 (N_3365,N_2348,N_1833);
xnor U3366 (N_3366,N_1985,N_2471);
nor U3367 (N_3367,N_1792,N_2453);
nand U3368 (N_3368,N_2242,N_1768);
nand U3369 (N_3369,N_2485,N_2896);
nand U3370 (N_3370,N_2983,N_1533);
nand U3371 (N_3371,N_2925,N_2021);
nand U3372 (N_3372,N_2190,N_2966);
nor U3373 (N_3373,N_2883,N_1602);
xnor U3374 (N_3374,N_2740,N_2828);
nand U3375 (N_3375,N_2335,N_2929);
or U3376 (N_3376,N_2848,N_2075);
or U3377 (N_3377,N_1933,N_1721);
or U3378 (N_3378,N_1872,N_1938);
or U3379 (N_3379,N_2096,N_1646);
or U3380 (N_3380,N_1632,N_1520);
or U3381 (N_3381,N_2144,N_2843);
and U3382 (N_3382,N_2884,N_2425);
or U3383 (N_3383,N_1682,N_2338);
or U3384 (N_3384,N_2470,N_2984);
and U3385 (N_3385,N_2170,N_1877);
xor U3386 (N_3386,N_1545,N_2518);
and U3387 (N_3387,N_2715,N_2764);
nor U3388 (N_3388,N_1651,N_1878);
xor U3389 (N_3389,N_1993,N_2243);
xor U3390 (N_3390,N_2856,N_1999);
or U3391 (N_3391,N_2589,N_2023);
and U3392 (N_3392,N_1630,N_1624);
or U3393 (N_3393,N_2138,N_1901);
nor U3394 (N_3394,N_1513,N_2423);
or U3395 (N_3395,N_2892,N_2475);
and U3396 (N_3396,N_1586,N_2194);
and U3397 (N_3397,N_2381,N_2324);
xnor U3398 (N_3398,N_1856,N_1614);
nor U3399 (N_3399,N_2358,N_2920);
xnor U3400 (N_3400,N_2259,N_2664);
and U3401 (N_3401,N_2246,N_2115);
xor U3402 (N_3402,N_1908,N_1554);
nor U3403 (N_3403,N_1596,N_2289);
xnor U3404 (N_3404,N_1766,N_2898);
or U3405 (N_3405,N_2750,N_2457);
and U3406 (N_3406,N_2773,N_1637);
nor U3407 (N_3407,N_1510,N_2072);
or U3408 (N_3408,N_1673,N_1956);
or U3409 (N_3409,N_2671,N_2844);
nand U3410 (N_3410,N_1848,N_2034);
and U3411 (N_3411,N_1998,N_2087);
nor U3412 (N_3412,N_2166,N_2552);
xnor U3413 (N_3413,N_1573,N_2523);
xnor U3414 (N_3414,N_2631,N_2900);
or U3415 (N_3415,N_1851,N_1949);
nand U3416 (N_3416,N_2616,N_2941);
nor U3417 (N_3417,N_2260,N_2840);
xor U3418 (N_3418,N_2035,N_1698);
or U3419 (N_3419,N_2760,N_1859);
or U3420 (N_3420,N_2748,N_2345);
nor U3421 (N_3421,N_2062,N_2219);
and U3422 (N_3422,N_1890,N_1882);
or U3423 (N_3423,N_1671,N_1638);
nor U3424 (N_3424,N_1919,N_2196);
xor U3425 (N_3425,N_2578,N_1742);
nand U3426 (N_3426,N_2139,N_1873);
xor U3427 (N_3427,N_2352,N_2944);
xor U3428 (N_3428,N_2968,N_1767);
xor U3429 (N_3429,N_2531,N_2989);
xor U3430 (N_3430,N_2620,N_2826);
nand U3431 (N_3431,N_2232,N_2150);
nor U3432 (N_3432,N_2753,N_1937);
or U3433 (N_3433,N_2707,N_2525);
nand U3434 (N_3434,N_2476,N_2839);
nor U3435 (N_3435,N_2145,N_2061);
nand U3436 (N_3436,N_1871,N_1580);
and U3437 (N_3437,N_1760,N_1780);
xor U3438 (N_3438,N_1703,N_2783);
or U3439 (N_3439,N_2108,N_1929);
xnor U3440 (N_3440,N_2530,N_1522);
or U3441 (N_3441,N_1590,N_2665);
or U3442 (N_3442,N_2913,N_1852);
xnor U3443 (N_3443,N_1785,N_2682);
or U3444 (N_3444,N_2028,N_2637);
and U3445 (N_3445,N_2859,N_2378);
xor U3446 (N_3446,N_2881,N_2793);
or U3447 (N_3447,N_1658,N_2849);
nor U3448 (N_3448,N_2223,N_1755);
and U3449 (N_3449,N_2831,N_1850);
or U3450 (N_3450,N_1910,N_2666);
and U3451 (N_3451,N_1819,N_2068);
nand U3452 (N_3452,N_1523,N_1569);
nand U3453 (N_3453,N_1975,N_2464);
or U3454 (N_3454,N_2256,N_2669);
xnor U3455 (N_3455,N_2469,N_2398);
nor U3456 (N_3456,N_2113,N_2010);
xor U3457 (N_3457,N_1817,N_1696);
nand U3458 (N_3458,N_2212,N_2506);
nand U3459 (N_3459,N_2498,N_1605);
xnor U3460 (N_3460,N_2776,N_2038);
nand U3461 (N_3461,N_2248,N_1739);
and U3462 (N_3462,N_1551,N_1536);
nand U3463 (N_3463,N_1519,N_1726);
and U3464 (N_3464,N_2442,N_2821);
or U3465 (N_3465,N_2089,N_1838);
or U3466 (N_3466,N_2807,N_2074);
nor U3467 (N_3467,N_1983,N_2644);
nor U3468 (N_3468,N_2460,N_2854);
nor U3469 (N_3469,N_2404,N_2585);
xor U3470 (N_3470,N_2593,N_1874);
and U3471 (N_3471,N_2441,N_1710);
xnor U3472 (N_3472,N_2325,N_2728);
nor U3473 (N_3473,N_2480,N_2714);
and U3474 (N_3474,N_2158,N_1532);
nor U3475 (N_3475,N_1697,N_2430);
or U3476 (N_3476,N_1589,N_2775);
nor U3477 (N_3477,N_2241,N_1897);
nand U3478 (N_3478,N_2809,N_1741);
nor U3479 (N_3479,N_2864,N_1700);
xnor U3480 (N_3480,N_1550,N_1926);
nand U3481 (N_3481,N_2281,N_1952);
or U3482 (N_3482,N_1907,N_2612);
and U3483 (N_3483,N_2698,N_2284);
or U3484 (N_3484,N_2333,N_1672);
and U3485 (N_3485,N_2967,N_1687);
nand U3486 (N_3486,N_1662,N_2395);
or U3487 (N_3487,N_1654,N_1627);
xor U3488 (N_3488,N_2491,N_2862);
or U3489 (N_3489,N_1680,N_2590);
or U3490 (N_3490,N_2686,N_2420);
and U3491 (N_3491,N_2192,N_2930);
and U3492 (N_3492,N_2436,N_2814);
and U3493 (N_3493,N_2043,N_2308);
or U3494 (N_3494,N_2180,N_1751);
or U3495 (N_3495,N_2315,N_2427);
nor U3496 (N_3496,N_2822,N_2226);
nand U3497 (N_3497,N_1774,N_2361);
or U3498 (N_3498,N_2638,N_1500);
xnor U3499 (N_3499,N_2322,N_1535);
nand U3500 (N_3500,N_1540,N_2081);
xor U3501 (N_3501,N_2290,N_1855);
and U3502 (N_3502,N_2572,N_2267);
xor U3503 (N_3503,N_2564,N_2412);
nor U3504 (N_3504,N_2567,N_2857);
nor U3505 (N_3505,N_1729,N_2261);
nand U3506 (N_3506,N_2107,N_2466);
xor U3507 (N_3507,N_2300,N_1895);
or U3508 (N_3508,N_1893,N_2225);
and U3509 (N_3509,N_2244,N_2504);
or U3510 (N_3510,N_1958,N_1842);
or U3511 (N_3511,N_1934,N_2845);
nor U3512 (N_3512,N_1980,N_1815);
or U3513 (N_3513,N_2213,N_2758);
nand U3514 (N_3514,N_2262,N_1772);
and U3515 (N_3515,N_2551,N_2800);
and U3516 (N_3516,N_1789,N_2287);
nand U3517 (N_3517,N_2935,N_2981);
nor U3518 (N_3518,N_1769,N_2744);
nand U3519 (N_3519,N_2229,N_2802);
nand U3520 (N_3520,N_2292,N_2779);
xor U3521 (N_3521,N_1948,N_2366);
nand U3522 (N_3522,N_1514,N_2580);
xor U3523 (N_3523,N_2093,N_2443);
xor U3524 (N_3524,N_2583,N_2774);
nand U3525 (N_3525,N_2510,N_2576);
or U3526 (N_3526,N_2538,N_1571);
or U3527 (N_3527,N_2514,N_2463);
or U3528 (N_3528,N_1608,N_2599);
nor U3529 (N_3529,N_1866,N_2027);
and U3530 (N_3530,N_2893,N_2553);
or U3531 (N_3531,N_2064,N_2376);
and U3532 (N_3532,N_2596,N_1735);
xor U3533 (N_3533,N_2922,N_2077);
xnor U3534 (N_3534,N_1941,N_1597);
or U3535 (N_3535,N_2976,N_2384);
nand U3536 (N_3536,N_2870,N_1549);
xor U3537 (N_3537,N_1706,N_2949);
nand U3538 (N_3538,N_2482,N_2128);
nand U3539 (N_3539,N_1884,N_2310);
nor U3540 (N_3540,N_2388,N_1905);
and U3541 (N_3541,N_2861,N_1557);
xnor U3542 (N_3542,N_1606,N_2731);
nor U3543 (N_3543,N_2368,N_2214);
xor U3544 (N_3544,N_2869,N_1888);
nor U3545 (N_3545,N_1581,N_1808);
or U3546 (N_3546,N_2084,N_2526);
or U3547 (N_3547,N_2597,N_1761);
xnor U3548 (N_3548,N_2257,N_1534);
nor U3549 (N_3549,N_2932,N_2183);
and U3550 (N_3550,N_2461,N_2495);
xnor U3551 (N_3551,N_1798,N_2397);
xor U3552 (N_3552,N_2692,N_2396);
nor U3553 (N_3553,N_2721,N_1973);
and U3554 (N_3554,N_2131,N_2709);
xnor U3555 (N_3555,N_2732,N_2958);
nor U3556 (N_3556,N_2312,N_2865);
and U3557 (N_3557,N_2201,N_1720);
xor U3558 (N_3558,N_2070,N_2317);
nand U3559 (N_3559,N_2847,N_2610);
or U3560 (N_3560,N_2777,N_1942);
or U3561 (N_3561,N_1600,N_2508);
nand U3562 (N_3562,N_2458,N_2249);
xor U3563 (N_3563,N_2003,N_2799);
and U3564 (N_3564,N_2927,N_2490);
xor U3565 (N_3565,N_1547,N_2602);
nor U3566 (N_3566,N_2727,N_2739);
or U3567 (N_3567,N_1634,N_2250);
nand U3568 (N_3568,N_2006,N_2106);
and U3569 (N_3569,N_2561,N_1748);
or U3570 (N_3570,N_2515,N_1659);
xor U3571 (N_3571,N_2816,N_2065);
nor U3572 (N_3572,N_1824,N_2606);
xnor U3573 (N_3573,N_2297,N_1857);
or U3574 (N_3574,N_2963,N_1797);
nand U3575 (N_3575,N_2330,N_1965);
nand U3576 (N_3576,N_1733,N_2169);
xnor U3577 (N_3577,N_2897,N_2220);
nor U3578 (N_3578,N_2887,N_2039);
xnor U3579 (N_3579,N_1969,N_2037);
nand U3580 (N_3580,N_1990,N_1920);
xor U3581 (N_3581,N_1771,N_2860);
xnor U3582 (N_3582,N_2007,N_2630);
or U3583 (N_3583,N_2306,N_2054);
xor U3584 (N_3584,N_2291,N_2749);
and U3585 (N_3585,N_2191,N_2507);
nand U3586 (N_3586,N_1615,N_2221);
nand U3587 (N_3587,N_2472,N_2364);
nor U3588 (N_3588,N_1839,N_1594);
nor U3589 (N_3589,N_2575,N_2533);
nor U3590 (N_3590,N_1786,N_2833);
or U3591 (N_3591,N_2677,N_2943);
and U3592 (N_3592,N_2613,N_2565);
nor U3593 (N_3593,N_2079,N_2782);
nor U3594 (N_3594,N_2033,N_2342);
xor U3595 (N_3595,N_2114,N_2133);
nor U3596 (N_3596,N_2147,N_1770);
nor U3597 (N_3597,N_1753,N_2626);
or U3598 (N_3598,N_2975,N_1940);
xor U3599 (N_3599,N_1821,N_2904);
and U3600 (N_3600,N_2735,N_1575);
or U3601 (N_3601,N_1582,N_2591);
and U3602 (N_3602,N_2247,N_2409);
or U3603 (N_3603,N_2952,N_1553);
xnor U3604 (N_3604,N_2537,N_1655);
xnor U3605 (N_3605,N_1653,N_2044);
nor U3606 (N_3606,N_2990,N_1854);
xnor U3607 (N_3607,N_2451,N_2083);
and U3608 (N_3608,N_2961,N_2400);
nor U3609 (N_3609,N_1507,N_2889);
xnor U3610 (N_3610,N_2650,N_2018);
nand U3611 (N_3611,N_2659,N_1778);
or U3612 (N_3612,N_1757,N_2416);
xor U3613 (N_3613,N_1959,N_2387);
or U3614 (N_3614,N_1754,N_2252);
nand U3615 (N_3615,N_2718,N_1649);
nor U3616 (N_3616,N_2394,N_2759);
nand U3617 (N_3617,N_2625,N_1684);
xnor U3618 (N_3618,N_2329,N_2500);
nor U3619 (N_3619,N_2118,N_2885);
and U3620 (N_3620,N_2742,N_2947);
xnor U3621 (N_3621,N_2350,N_1640);
xor U3622 (N_3622,N_2948,N_2684);
and U3623 (N_3623,N_1583,N_2058);
nand U3624 (N_3624,N_2704,N_2627);
xnor U3625 (N_3625,N_2547,N_2679);
or U3626 (N_3626,N_2770,N_1845);
nor U3627 (N_3627,N_1558,N_2059);
and U3628 (N_3628,N_2954,N_2946);
or U3629 (N_3629,N_2639,N_2331);
nand U3630 (N_3630,N_1588,N_2852);
xor U3631 (N_3631,N_2600,N_2689);
nand U3632 (N_3632,N_2874,N_2432);
nand U3633 (N_3633,N_1809,N_1679);
xor U3634 (N_3634,N_1688,N_1800);
or U3635 (N_3635,N_2588,N_1917);
and U3636 (N_3636,N_2051,N_2651);
or U3637 (N_3637,N_1647,N_2303);
or U3638 (N_3638,N_1788,N_2919);
or U3639 (N_3639,N_2173,N_2712);
nor U3640 (N_3640,N_2030,N_1970);
nor U3641 (N_3641,N_1944,N_2098);
xor U3642 (N_3642,N_2916,N_1725);
xnor U3643 (N_3643,N_2586,N_2521);
nand U3644 (N_3644,N_2813,N_2142);
nor U3645 (N_3645,N_2301,N_1793);
or U3646 (N_3646,N_1543,N_1997);
or U3647 (N_3647,N_2137,N_2266);
or U3648 (N_3648,N_2497,N_2265);
and U3649 (N_3649,N_2608,N_1628);
and U3650 (N_3650,N_2015,N_1876);
or U3651 (N_3651,N_1635,N_2032);
nand U3652 (N_3652,N_2078,N_1795);
and U3653 (N_3653,N_1524,N_2969);
xnor U3654 (N_3654,N_2163,N_1731);
xor U3655 (N_3655,N_2197,N_2629);
and U3656 (N_3656,N_1713,N_1953);
or U3657 (N_3657,N_1883,N_2768);
and U3658 (N_3658,N_2379,N_2483);
or U3659 (N_3659,N_2193,N_2393);
and U3660 (N_3660,N_1537,N_1902);
and U3661 (N_3661,N_2499,N_2004);
nor U3662 (N_3662,N_2218,N_1650);
nor U3663 (N_3663,N_2390,N_1648);
xor U3664 (N_3664,N_2836,N_1960);
or U3665 (N_3665,N_2928,N_2923);
or U3666 (N_3666,N_2012,N_1746);
nor U3667 (N_3667,N_1823,N_2391);
or U3668 (N_3668,N_2179,N_2901);
or U3669 (N_3669,N_2688,N_2016);
or U3670 (N_3670,N_1564,N_2569);
xnor U3671 (N_3671,N_2355,N_2529);
or U3672 (N_3672,N_2931,N_1610);
xor U3673 (N_3673,N_2447,N_2053);
and U3674 (N_3674,N_1641,N_2435);
and U3675 (N_3675,N_1939,N_2337);
nand U3676 (N_3676,N_2545,N_2945);
and U3677 (N_3677,N_2371,N_2866);
and U3678 (N_3678,N_2386,N_2382);
xnor U3679 (N_3679,N_2233,N_2410);
xor U3680 (N_3680,N_1693,N_2235);
or U3681 (N_3681,N_1708,N_1657);
xnor U3682 (N_3682,N_2152,N_2050);
nand U3683 (N_3683,N_2851,N_2135);
nor U3684 (N_3684,N_2556,N_2772);
or U3685 (N_3685,N_2953,N_1900);
and U3686 (N_3686,N_1779,N_1816);
and U3687 (N_3687,N_1661,N_2743);
xnor U3688 (N_3688,N_2598,N_2534);
nor U3689 (N_3689,N_2132,N_2363);
and U3690 (N_3690,N_2200,N_1928);
and U3691 (N_3691,N_2713,N_2473);
nor U3692 (N_3692,N_1552,N_2210);
nor U3693 (N_3693,N_2048,N_1619);
and U3694 (N_3694,N_1629,N_1787);
xnor U3695 (N_3695,N_1865,N_1962);
or U3696 (N_3696,N_2481,N_2673);
or U3697 (N_3697,N_2595,N_2230);
or U3698 (N_3698,N_2652,N_1568);
and U3699 (N_3699,N_1728,N_2574);
and U3700 (N_3700,N_1591,N_2339);
nand U3701 (N_3701,N_2939,N_2660);
or U3702 (N_3702,N_1711,N_2658);
nand U3703 (N_3703,N_2678,N_2767);
and U3704 (N_3704,N_2734,N_2886);
and U3705 (N_3705,N_2063,N_1561);
and U3706 (N_3706,N_1810,N_1717);
nand U3707 (N_3707,N_1971,N_1744);
xnor U3708 (N_3708,N_2653,N_1668);
and U3709 (N_3709,N_2621,N_2392);
xor U3710 (N_3710,N_1724,N_2524);
or U3711 (N_3711,N_2380,N_1730);
nand U3712 (N_3712,N_2206,N_2005);
and U3713 (N_3713,N_1799,N_2437);
nand U3714 (N_3714,N_1508,N_1555);
nor U3715 (N_3715,N_2662,N_2544);
nor U3716 (N_3716,N_2670,N_2972);
or U3717 (N_3717,N_2607,N_2663);
nor U3718 (N_3718,N_2609,N_1598);
nand U3719 (N_3719,N_2908,N_1616);
and U3720 (N_3720,N_1906,N_1927);
or U3721 (N_3721,N_1840,N_2161);
nor U3722 (N_3722,N_2372,N_1681);
xnor U3723 (N_3723,N_2882,N_1782);
xnor U3724 (N_3724,N_2307,N_2680);
and U3725 (N_3725,N_2867,N_2542);
or U3726 (N_3726,N_2817,N_1945);
nor U3727 (N_3727,N_2815,N_2710);
and U3728 (N_3728,N_2628,N_2332);
nand U3729 (N_3729,N_2755,N_1689);
xnor U3730 (N_3730,N_2438,N_2738);
or U3731 (N_3731,N_1750,N_2987);
xor U3732 (N_3732,N_2520,N_1592);
nor U3733 (N_3733,N_1891,N_2239);
nor U3734 (N_3734,N_2017,N_2878);
nand U3735 (N_3735,N_2655,N_2110);
and U3736 (N_3736,N_2724,N_2667);
nor U3737 (N_3737,N_1512,N_1506);
nand U3738 (N_3738,N_2635,N_1813);
and U3739 (N_3739,N_2143,N_2182);
nor U3740 (N_3740,N_2805,N_2141);
nor U3741 (N_3741,N_2611,N_2795);
nor U3742 (N_3742,N_1880,N_2029);
xor U3743 (N_3743,N_2104,N_2955);
and U3744 (N_3744,N_2837,N_1836);
nand U3745 (N_3745,N_2873,N_2399);
nand U3746 (N_3746,N_2298,N_2493);
and U3747 (N_3747,N_1849,N_2253);
or U3748 (N_3748,N_1570,N_2216);
nor U3749 (N_3749,N_1743,N_2105);
nor U3750 (N_3750,N_2618,N_2148);
and U3751 (N_3751,N_2596,N_2094);
or U3752 (N_3752,N_1642,N_2282);
and U3753 (N_3753,N_2739,N_2245);
nor U3754 (N_3754,N_2688,N_2973);
nand U3755 (N_3755,N_2658,N_1993);
nand U3756 (N_3756,N_2985,N_2941);
nand U3757 (N_3757,N_2823,N_2711);
and U3758 (N_3758,N_1825,N_2945);
and U3759 (N_3759,N_1976,N_2508);
and U3760 (N_3760,N_2074,N_2646);
nor U3761 (N_3761,N_1988,N_2449);
and U3762 (N_3762,N_2412,N_2609);
and U3763 (N_3763,N_2156,N_2514);
nor U3764 (N_3764,N_2795,N_2044);
nand U3765 (N_3765,N_1717,N_1725);
xor U3766 (N_3766,N_1845,N_1774);
nand U3767 (N_3767,N_1784,N_1971);
nor U3768 (N_3768,N_2728,N_2190);
nor U3769 (N_3769,N_2892,N_2384);
nand U3770 (N_3770,N_1583,N_1593);
nand U3771 (N_3771,N_2558,N_2021);
nand U3772 (N_3772,N_2986,N_2706);
and U3773 (N_3773,N_1996,N_2528);
and U3774 (N_3774,N_2277,N_2857);
nor U3775 (N_3775,N_1561,N_1648);
nor U3776 (N_3776,N_1919,N_1686);
nand U3777 (N_3777,N_2474,N_1974);
xor U3778 (N_3778,N_2982,N_2914);
xor U3779 (N_3779,N_1683,N_2672);
and U3780 (N_3780,N_2719,N_1933);
nand U3781 (N_3781,N_2318,N_2694);
nand U3782 (N_3782,N_1659,N_2615);
and U3783 (N_3783,N_1546,N_1962);
nor U3784 (N_3784,N_2360,N_1673);
xor U3785 (N_3785,N_2096,N_1882);
and U3786 (N_3786,N_2695,N_2392);
xor U3787 (N_3787,N_2463,N_2784);
and U3788 (N_3788,N_2111,N_2915);
and U3789 (N_3789,N_2794,N_2864);
and U3790 (N_3790,N_2364,N_1711);
nor U3791 (N_3791,N_2046,N_1654);
nor U3792 (N_3792,N_1569,N_1530);
xnor U3793 (N_3793,N_1511,N_1943);
xnor U3794 (N_3794,N_1658,N_1761);
xor U3795 (N_3795,N_2303,N_2318);
and U3796 (N_3796,N_1864,N_1861);
nor U3797 (N_3797,N_1817,N_2303);
nor U3798 (N_3798,N_2634,N_2371);
and U3799 (N_3799,N_2998,N_2515);
nand U3800 (N_3800,N_2124,N_1761);
nand U3801 (N_3801,N_1830,N_2554);
nor U3802 (N_3802,N_1559,N_2810);
nor U3803 (N_3803,N_2480,N_2609);
and U3804 (N_3804,N_1599,N_1896);
nor U3805 (N_3805,N_2051,N_2182);
nand U3806 (N_3806,N_2429,N_1941);
and U3807 (N_3807,N_2730,N_2097);
nor U3808 (N_3808,N_2765,N_1964);
xor U3809 (N_3809,N_2829,N_2937);
and U3810 (N_3810,N_1795,N_2072);
xnor U3811 (N_3811,N_2723,N_2372);
nor U3812 (N_3812,N_1557,N_2620);
nor U3813 (N_3813,N_2062,N_1964);
and U3814 (N_3814,N_1736,N_1969);
xnor U3815 (N_3815,N_2616,N_2869);
xor U3816 (N_3816,N_1608,N_2437);
or U3817 (N_3817,N_2839,N_1826);
xor U3818 (N_3818,N_2121,N_1726);
nand U3819 (N_3819,N_2920,N_1619);
and U3820 (N_3820,N_2414,N_2272);
or U3821 (N_3821,N_2575,N_2306);
nor U3822 (N_3822,N_1677,N_2864);
nor U3823 (N_3823,N_2715,N_2557);
nor U3824 (N_3824,N_1859,N_2532);
nor U3825 (N_3825,N_2419,N_1951);
and U3826 (N_3826,N_2903,N_2904);
or U3827 (N_3827,N_2367,N_1604);
nand U3828 (N_3828,N_2874,N_1530);
nand U3829 (N_3829,N_2361,N_2341);
xnor U3830 (N_3830,N_1665,N_1550);
xnor U3831 (N_3831,N_2418,N_2089);
nor U3832 (N_3832,N_1609,N_1617);
xor U3833 (N_3833,N_2912,N_1786);
and U3834 (N_3834,N_2161,N_2329);
nand U3835 (N_3835,N_2313,N_1861);
or U3836 (N_3836,N_2131,N_1515);
nand U3837 (N_3837,N_2525,N_2643);
nand U3838 (N_3838,N_1581,N_1991);
and U3839 (N_3839,N_2439,N_1512);
xor U3840 (N_3840,N_2188,N_2730);
and U3841 (N_3841,N_2351,N_1514);
and U3842 (N_3842,N_2103,N_2206);
nor U3843 (N_3843,N_2227,N_1931);
and U3844 (N_3844,N_1791,N_2273);
xnor U3845 (N_3845,N_1771,N_1776);
nor U3846 (N_3846,N_2836,N_2305);
or U3847 (N_3847,N_1527,N_1859);
nor U3848 (N_3848,N_2361,N_1783);
nand U3849 (N_3849,N_1721,N_2664);
xor U3850 (N_3850,N_1907,N_1511);
or U3851 (N_3851,N_1628,N_2558);
and U3852 (N_3852,N_1595,N_2505);
or U3853 (N_3853,N_2551,N_1552);
and U3854 (N_3854,N_2801,N_2689);
nor U3855 (N_3855,N_2401,N_1725);
nor U3856 (N_3856,N_2897,N_2778);
nor U3857 (N_3857,N_1787,N_1594);
nand U3858 (N_3858,N_1758,N_1637);
xor U3859 (N_3859,N_2391,N_1898);
nor U3860 (N_3860,N_2931,N_2465);
xor U3861 (N_3861,N_1656,N_2880);
or U3862 (N_3862,N_1559,N_1607);
nor U3863 (N_3863,N_2037,N_2540);
and U3864 (N_3864,N_2394,N_2999);
nand U3865 (N_3865,N_2656,N_2134);
nand U3866 (N_3866,N_2506,N_2159);
xnor U3867 (N_3867,N_2312,N_2962);
xnor U3868 (N_3868,N_1714,N_2826);
and U3869 (N_3869,N_2287,N_2498);
and U3870 (N_3870,N_2979,N_2969);
or U3871 (N_3871,N_1759,N_1595);
and U3872 (N_3872,N_2313,N_2948);
nor U3873 (N_3873,N_2547,N_2299);
and U3874 (N_3874,N_2089,N_2182);
or U3875 (N_3875,N_1719,N_1511);
and U3876 (N_3876,N_2617,N_2180);
or U3877 (N_3877,N_2502,N_2863);
or U3878 (N_3878,N_1995,N_2477);
and U3879 (N_3879,N_1675,N_1551);
and U3880 (N_3880,N_2215,N_1870);
or U3881 (N_3881,N_2583,N_2528);
nor U3882 (N_3882,N_2430,N_1528);
xor U3883 (N_3883,N_1621,N_2576);
or U3884 (N_3884,N_1583,N_2061);
nand U3885 (N_3885,N_2290,N_2843);
or U3886 (N_3886,N_2875,N_2611);
or U3887 (N_3887,N_2955,N_2922);
xor U3888 (N_3888,N_2483,N_1867);
and U3889 (N_3889,N_2979,N_2251);
or U3890 (N_3890,N_2805,N_1787);
nand U3891 (N_3891,N_2970,N_2407);
xor U3892 (N_3892,N_2919,N_2785);
or U3893 (N_3893,N_2188,N_2379);
nand U3894 (N_3894,N_2668,N_2003);
and U3895 (N_3895,N_2721,N_2120);
or U3896 (N_3896,N_2131,N_2608);
or U3897 (N_3897,N_2217,N_1818);
xor U3898 (N_3898,N_1827,N_1936);
nand U3899 (N_3899,N_1823,N_1683);
nand U3900 (N_3900,N_2357,N_1868);
nor U3901 (N_3901,N_2514,N_2182);
and U3902 (N_3902,N_2728,N_1752);
nor U3903 (N_3903,N_2071,N_1954);
and U3904 (N_3904,N_2186,N_2801);
nand U3905 (N_3905,N_1677,N_2161);
and U3906 (N_3906,N_2298,N_1518);
and U3907 (N_3907,N_2653,N_1998);
or U3908 (N_3908,N_1761,N_1930);
xor U3909 (N_3909,N_1719,N_2241);
nand U3910 (N_3910,N_1909,N_1553);
nor U3911 (N_3911,N_2756,N_2988);
nor U3912 (N_3912,N_1731,N_1639);
nand U3913 (N_3913,N_1875,N_2369);
xor U3914 (N_3914,N_1854,N_2175);
nand U3915 (N_3915,N_2534,N_2992);
nor U3916 (N_3916,N_2691,N_1504);
or U3917 (N_3917,N_2093,N_1556);
nor U3918 (N_3918,N_2380,N_2750);
xnor U3919 (N_3919,N_1799,N_2398);
nand U3920 (N_3920,N_2802,N_2044);
nand U3921 (N_3921,N_2071,N_1551);
or U3922 (N_3922,N_2025,N_2684);
and U3923 (N_3923,N_2037,N_2170);
xnor U3924 (N_3924,N_1839,N_2847);
or U3925 (N_3925,N_2437,N_2252);
nand U3926 (N_3926,N_2394,N_2790);
nor U3927 (N_3927,N_2782,N_2373);
or U3928 (N_3928,N_2520,N_2453);
and U3929 (N_3929,N_2807,N_2985);
or U3930 (N_3930,N_2663,N_2336);
and U3931 (N_3931,N_2829,N_2941);
nand U3932 (N_3932,N_2845,N_1635);
nor U3933 (N_3933,N_2020,N_2635);
or U3934 (N_3934,N_1542,N_2742);
and U3935 (N_3935,N_2912,N_2637);
nor U3936 (N_3936,N_2423,N_2266);
nor U3937 (N_3937,N_2305,N_1699);
and U3938 (N_3938,N_1759,N_2093);
and U3939 (N_3939,N_1646,N_2527);
nand U3940 (N_3940,N_1869,N_2509);
or U3941 (N_3941,N_2077,N_2104);
nand U3942 (N_3942,N_1648,N_2024);
and U3943 (N_3943,N_1735,N_2325);
or U3944 (N_3944,N_2838,N_2441);
or U3945 (N_3945,N_2087,N_1922);
nor U3946 (N_3946,N_2933,N_1716);
nand U3947 (N_3947,N_2036,N_2851);
xnor U3948 (N_3948,N_2430,N_2674);
xnor U3949 (N_3949,N_2183,N_2462);
or U3950 (N_3950,N_1954,N_2085);
or U3951 (N_3951,N_1563,N_1828);
xnor U3952 (N_3952,N_2493,N_2920);
nand U3953 (N_3953,N_2419,N_2043);
nand U3954 (N_3954,N_2786,N_1656);
and U3955 (N_3955,N_2836,N_2037);
or U3956 (N_3956,N_2036,N_2335);
xnor U3957 (N_3957,N_2760,N_2961);
nor U3958 (N_3958,N_1790,N_1820);
or U3959 (N_3959,N_1999,N_2956);
and U3960 (N_3960,N_2130,N_2860);
nand U3961 (N_3961,N_2746,N_2974);
nor U3962 (N_3962,N_2615,N_1820);
nand U3963 (N_3963,N_2391,N_1767);
or U3964 (N_3964,N_1999,N_1821);
nand U3965 (N_3965,N_2103,N_2748);
nor U3966 (N_3966,N_1908,N_2043);
nand U3967 (N_3967,N_2636,N_1745);
or U3968 (N_3968,N_1808,N_2545);
xnor U3969 (N_3969,N_2643,N_1965);
and U3970 (N_3970,N_2080,N_2819);
xor U3971 (N_3971,N_2412,N_1985);
nor U3972 (N_3972,N_2620,N_1919);
nor U3973 (N_3973,N_1631,N_2327);
or U3974 (N_3974,N_2525,N_2401);
xor U3975 (N_3975,N_2454,N_2628);
and U3976 (N_3976,N_2763,N_2392);
and U3977 (N_3977,N_1810,N_1557);
or U3978 (N_3978,N_2407,N_1684);
or U3979 (N_3979,N_1853,N_2862);
and U3980 (N_3980,N_1879,N_1752);
nor U3981 (N_3981,N_2750,N_1860);
and U3982 (N_3982,N_2870,N_2093);
nor U3983 (N_3983,N_2203,N_2880);
and U3984 (N_3984,N_1558,N_1565);
nand U3985 (N_3985,N_2869,N_1905);
xor U3986 (N_3986,N_2728,N_1744);
and U3987 (N_3987,N_2598,N_2511);
and U3988 (N_3988,N_1722,N_2479);
nand U3989 (N_3989,N_1921,N_1872);
and U3990 (N_3990,N_2801,N_2539);
or U3991 (N_3991,N_2630,N_2531);
nor U3992 (N_3992,N_2762,N_2282);
xnor U3993 (N_3993,N_2725,N_2196);
nor U3994 (N_3994,N_2049,N_2436);
nand U3995 (N_3995,N_2068,N_2606);
xor U3996 (N_3996,N_1959,N_1810);
nand U3997 (N_3997,N_2696,N_1788);
and U3998 (N_3998,N_1742,N_2131);
nor U3999 (N_3999,N_1926,N_2122);
nand U4000 (N_4000,N_2408,N_1675);
or U4001 (N_4001,N_2046,N_2883);
or U4002 (N_4002,N_2984,N_2729);
nand U4003 (N_4003,N_2632,N_2393);
nand U4004 (N_4004,N_1660,N_1952);
nor U4005 (N_4005,N_2871,N_2230);
and U4006 (N_4006,N_1958,N_1613);
nor U4007 (N_4007,N_1879,N_2488);
nor U4008 (N_4008,N_1647,N_2743);
or U4009 (N_4009,N_1858,N_2085);
or U4010 (N_4010,N_1936,N_2681);
xor U4011 (N_4011,N_2904,N_2063);
nor U4012 (N_4012,N_2433,N_2973);
xnor U4013 (N_4013,N_2839,N_1609);
xor U4014 (N_4014,N_2659,N_2629);
or U4015 (N_4015,N_2103,N_2000);
nor U4016 (N_4016,N_2071,N_1639);
and U4017 (N_4017,N_2224,N_2208);
or U4018 (N_4018,N_2348,N_2262);
nor U4019 (N_4019,N_1659,N_1582);
and U4020 (N_4020,N_2707,N_2225);
nor U4021 (N_4021,N_1892,N_2044);
xnor U4022 (N_4022,N_1725,N_2339);
or U4023 (N_4023,N_2034,N_1659);
nand U4024 (N_4024,N_1947,N_2510);
xnor U4025 (N_4025,N_2816,N_2760);
nor U4026 (N_4026,N_1906,N_2188);
and U4027 (N_4027,N_1642,N_2239);
nor U4028 (N_4028,N_2791,N_2500);
and U4029 (N_4029,N_1543,N_2164);
and U4030 (N_4030,N_2330,N_2879);
or U4031 (N_4031,N_2016,N_2818);
or U4032 (N_4032,N_2073,N_2687);
xnor U4033 (N_4033,N_1690,N_2977);
or U4034 (N_4034,N_2465,N_2357);
and U4035 (N_4035,N_2618,N_2169);
or U4036 (N_4036,N_1612,N_2279);
and U4037 (N_4037,N_2604,N_1758);
nand U4038 (N_4038,N_2841,N_2240);
xnor U4039 (N_4039,N_1805,N_2944);
xor U4040 (N_4040,N_1574,N_1910);
and U4041 (N_4041,N_2861,N_2006);
and U4042 (N_4042,N_2591,N_2432);
nand U4043 (N_4043,N_1849,N_2339);
or U4044 (N_4044,N_1771,N_1827);
xnor U4045 (N_4045,N_1751,N_1840);
and U4046 (N_4046,N_2557,N_1981);
or U4047 (N_4047,N_2457,N_1880);
or U4048 (N_4048,N_2639,N_2022);
nor U4049 (N_4049,N_2372,N_2850);
or U4050 (N_4050,N_2114,N_1891);
and U4051 (N_4051,N_2019,N_2897);
xnor U4052 (N_4052,N_1753,N_2941);
nor U4053 (N_4053,N_2924,N_2192);
nor U4054 (N_4054,N_2664,N_2236);
nand U4055 (N_4055,N_2189,N_2600);
nor U4056 (N_4056,N_1991,N_2089);
xnor U4057 (N_4057,N_1568,N_2241);
nand U4058 (N_4058,N_2973,N_2023);
or U4059 (N_4059,N_2624,N_1856);
or U4060 (N_4060,N_1743,N_2691);
and U4061 (N_4061,N_2662,N_2630);
nor U4062 (N_4062,N_2794,N_2554);
xnor U4063 (N_4063,N_1797,N_2650);
xnor U4064 (N_4064,N_2182,N_2215);
xor U4065 (N_4065,N_2256,N_2118);
and U4066 (N_4066,N_2646,N_2789);
nor U4067 (N_4067,N_2143,N_1826);
or U4068 (N_4068,N_2997,N_2851);
nand U4069 (N_4069,N_1642,N_2229);
nand U4070 (N_4070,N_1940,N_2257);
nor U4071 (N_4071,N_2624,N_2965);
nand U4072 (N_4072,N_2265,N_1679);
nand U4073 (N_4073,N_1880,N_2319);
nor U4074 (N_4074,N_2495,N_2755);
and U4075 (N_4075,N_2485,N_2810);
or U4076 (N_4076,N_2443,N_2261);
nand U4077 (N_4077,N_2629,N_2993);
nor U4078 (N_4078,N_2887,N_2522);
nor U4079 (N_4079,N_1751,N_1523);
or U4080 (N_4080,N_2921,N_2644);
nand U4081 (N_4081,N_1732,N_2367);
nand U4082 (N_4082,N_2350,N_2998);
xor U4083 (N_4083,N_2252,N_2278);
nand U4084 (N_4084,N_2237,N_2632);
or U4085 (N_4085,N_2293,N_2735);
xnor U4086 (N_4086,N_2425,N_2524);
nor U4087 (N_4087,N_1916,N_2072);
nor U4088 (N_4088,N_1746,N_1615);
or U4089 (N_4089,N_2909,N_2830);
nor U4090 (N_4090,N_2919,N_2180);
and U4091 (N_4091,N_1742,N_1573);
xor U4092 (N_4092,N_1730,N_2178);
nor U4093 (N_4093,N_1742,N_1634);
nand U4094 (N_4094,N_2262,N_1790);
nor U4095 (N_4095,N_1526,N_2303);
nor U4096 (N_4096,N_2976,N_2305);
and U4097 (N_4097,N_2350,N_2638);
or U4098 (N_4098,N_2662,N_1773);
xor U4099 (N_4099,N_2908,N_1516);
nor U4100 (N_4100,N_2827,N_2573);
and U4101 (N_4101,N_2246,N_1766);
nand U4102 (N_4102,N_2320,N_2911);
or U4103 (N_4103,N_1772,N_2801);
and U4104 (N_4104,N_1717,N_2601);
xnor U4105 (N_4105,N_1806,N_2821);
xor U4106 (N_4106,N_1557,N_2242);
or U4107 (N_4107,N_2566,N_2156);
nand U4108 (N_4108,N_1803,N_1678);
and U4109 (N_4109,N_1602,N_2672);
nand U4110 (N_4110,N_2665,N_2590);
xnor U4111 (N_4111,N_1755,N_1803);
or U4112 (N_4112,N_1644,N_2515);
xor U4113 (N_4113,N_2954,N_2302);
xnor U4114 (N_4114,N_2976,N_2415);
and U4115 (N_4115,N_2857,N_2574);
nor U4116 (N_4116,N_1506,N_1680);
and U4117 (N_4117,N_2411,N_2383);
nor U4118 (N_4118,N_1955,N_2654);
nor U4119 (N_4119,N_2774,N_2283);
xor U4120 (N_4120,N_2701,N_2394);
or U4121 (N_4121,N_2733,N_2841);
xnor U4122 (N_4122,N_2914,N_2284);
xor U4123 (N_4123,N_2775,N_2324);
and U4124 (N_4124,N_2007,N_1594);
nand U4125 (N_4125,N_1839,N_2713);
and U4126 (N_4126,N_2202,N_1967);
xnor U4127 (N_4127,N_2158,N_2256);
and U4128 (N_4128,N_1752,N_2945);
and U4129 (N_4129,N_2306,N_1772);
nand U4130 (N_4130,N_2899,N_1575);
and U4131 (N_4131,N_2644,N_2370);
xnor U4132 (N_4132,N_2992,N_2512);
nand U4133 (N_4133,N_1578,N_2304);
or U4134 (N_4134,N_1594,N_2693);
nand U4135 (N_4135,N_1753,N_2661);
or U4136 (N_4136,N_2357,N_2802);
nand U4137 (N_4137,N_1911,N_2296);
and U4138 (N_4138,N_2382,N_2369);
nand U4139 (N_4139,N_2272,N_2608);
xnor U4140 (N_4140,N_2923,N_2837);
or U4141 (N_4141,N_1641,N_2251);
nor U4142 (N_4142,N_2814,N_1907);
or U4143 (N_4143,N_2800,N_1532);
or U4144 (N_4144,N_2480,N_1660);
xor U4145 (N_4145,N_2531,N_2565);
xor U4146 (N_4146,N_2039,N_1626);
nand U4147 (N_4147,N_1603,N_1514);
nand U4148 (N_4148,N_2570,N_1761);
or U4149 (N_4149,N_1868,N_2467);
nor U4150 (N_4150,N_2733,N_2330);
nor U4151 (N_4151,N_2724,N_2440);
or U4152 (N_4152,N_2032,N_2628);
or U4153 (N_4153,N_2850,N_2135);
or U4154 (N_4154,N_1674,N_2326);
nand U4155 (N_4155,N_2447,N_2168);
nand U4156 (N_4156,N_1947,N_2026);
nand U4157 (N_4157,N_2988,N_2989);
nor U4158 (N_4158,N_2797,N_1854);
nor U4159 (N_4159,N_1818,N_1958);
nand U4160 (N_4160,N_2264,N_2083);
xnor U4161 (N_4161,N_2033,N_1848);
nor U4162 (N_4162,N_2775,N_2417);
nand U4163 (N_4163,N_2337,N_2374);
or U4164 (N_4164,N_1696,N_2435);
nor U4165 (N_4165,N_1749,N_1933);
xnor U4166 (N_4166,N_2718,N_1737);
nand U4167 (N_4167,N_2480,N_1516);
nor U4168 (N_4168,N_2430,N_2873);
nor U4169 (N_4169,N_2080,N_2315);
nand U4170 (N_4170,N_1696,N_2372);
nand U4171 (N_4171,N_2121,N_1824);
or U4172 (N_4172,N_1746,N_2082);
or U4173 (N_4173,N_2142,N_1892);
and U4174 (N_4174,N_2766,N_2654);
nand U4175 (N_4175,N_2156,N_2369);
xnor U4176 (N_4176,N_2709,N_1504);
nand U4177 (N_4177,N_1695,N_2544);
nand U4178 (N_4178,N_2962,N_2372);
or U4179 (N_4179,N_1524,N_1929);
nand U4180 (N_4180,N_1875,N_1610);
or U4181 (N_4181,N_1929,N_1779);
nand U4182 (N_4182,N_2841,N_1721);
xnor U4183 (N_4183,N_2720,N_2856);
or U4184 (N_4184,N_2094,N_2460);
xnor U4185 (N_4185,N_2065,N_1992);
nand U4186 (N_4186,N_2845,N_2624);
xor U4187 (N_4187,N_2893,N_1894);
and U4188 (N_4188,N_2983,N_2623);
and U4189 (N_4189,N_2208,N_1677);
and U4190 (N_4190,N_1644,N_2439);
or U4191 (N_4191,N_2171,N_1527);
or U4192 (N_4192,N_2451,N_2103);
and U4193 (N_4193,N_2082,N_2437);
nor U4194 (N_4194,N_2550,N_2152);
xnor U4195 (N_4195,N_2824,N_2216);
nand U4196 (N_4196,N_2413,N_1571);
and U4197 (N_4197,N_1883,N_2611);
or U4198 (N_4198,N_1649,N_1937);
nor U4199 (N_4199,N_1947,N_2993);
xor U4200 (N_4200,N_1827,N_2195);
or U4201 (N_4201,N_1608,N_1901);
nor U4202 (N_4202,N_1536,N_1649);
nand U4203 (N_4203,N_1860,N_2934);
nand U4204 (N_4204,N_1807,N_2927);
nor U4205 (N_4205,N_1564,N_2109);
xnor U4206 (N_4206,N_2807,N_2716);
nand U4207 (N_4207,N_1521,N_2997);
xor U4208 (N_4208,N_2856,N_2094);
and U4209 (N_4209,N_2940,N_2077);
and U4210 (N_4210,N_2699,N_2955);
nand U4211 (N_4211,N_1975,N_2041);
nand U4212 (N_4212,N_1710,N_2748);
xnor U4213 (N_4213,N_2615,N_2286);
or U4214 (N_4214,N_2928,N_1986);
nor U4215 (N_4215,N_2913,N_2927);
nor U4216 (N_4216,N_1631,N_2349);
xor U4217 (N_4217,N_1597,N_1793);
or U4218 (N_4218,N_2378,N_2599);
nand U4219 (N_4219,N_1784,N_2441);
and U4220 (N_4220,N_2040,N_2074);
nand U4221 (N_4221,N_2359,N_2010);
xor U4222 (N_4222,N_1690,N_1843);
nor U4223 (N_4223,N_2335,N_1518);
nand U4224 (N_4224,N_2589,N_2796);
or U4225 (N_4225,N_2286,N_1760);
nand U4226 (N_4226,N_2888,N_2126);
and U4227 (N_4227,N_2489,N_1685);
xor U4228 (N_4228,N_2407,N_1526);
nand U4229 (N_4229,N_2057,N_2682);
or U4230 (N_4230,N_2328,N_2507);
nand U4231 (N_4231,N_1982,N_1680);
nor U4232 (N_4232,N_2336,N_2016);
nand U4233 (N_4233,N_2624,N_2469);
nor U4234 (N_4234,N_2062,N_2474);
nor U4235 (N_4235,N_2276,N_2452);
or U4236 (N_4236,N_2350,N_2020);
and U4237 (N_4237,N_1701,N_2632);
xnor U4238 (N_4238,N_1968,N_2967);
and U4239 (N_4239,N_2680,N_2498);
nand U4240 (N_4240,N_2149,N_2250);
nand U4241 (N_4241,N_1581,N_1658);
nor U4242 (N_4242,N_2037,N_1668);
and U4243 (N_4243,N_2369,N_2786);
and U4244 (N_4244,N_2701,N_2708);
nor U4245 (N_4245,N_1813,N_1551);
nand U4246 (N_4246,N_1501,N_2708);
or U4247 (N_4247,N_2809,N_2897);
nor U4248 (N_4248,N_2728,N_2734);
or U4249 (N_4249,N_2913,N_2327);
or U4250 (N_4250,N_1763,N_2916);
or U4251 (N_4251,N_2329,N_2488);
or U4252 (N_4252,N_1651,N_2746);
xnor U4253 (N_4253,N_1505,N_1991);
nand U4254 (N_4254,N_1538,N_1533);
xnor U4255 (N_4255,N_2705,N_2804);
and U4256 (N_4256,N_1645,N_2974);
nor U4257 (N_4257,N_1930,N_2202);
nand U4258 (N_4258,N_2406,N_2700);
and U4259 (N_4259,N_2840,N_1883);
and U4260 (N_4260,N_1862,N_2283);
nor U4261 (N_4261,N_1714,N_2603);
nor U4262 (N_4262,N_2918,N_1804);
xor U4263 (N_4263,N_2162,N_1549);
or U4264 (N_4264,N_2230,N_2266);
nor U4265 (N_4265,N_1667,N_2609);
nor U4266 (N_4266,N_2087,N_1538);
or U4267 (N_4267,N_1746,N_1523);
nand U4268 (N_4268,N_1690,N_1551);
nor U4269 (N_4269,N_2380,N_2859);
nand U4270 (N_4270,N_1696,N_1673);
or U4271 (N_4271,N_2810,N_2162);
or U4272 (N_4272,N_2558,N_1880);
nand U4273 (N_4273,N_2978,N_1801);
and U4274 (N_4274,N_2763,N_2173);
and U4275 (N_4275,N_1899,N_2104);
or U4276 (N_4276,N_2474,N_1552);
and U4277 (N_4277,N_2210,N_2662);
nor U4278 (N_4278,N_1698,N_2213);
xor U4279 (N_4279,N_2814,N_2126);
nor U4280 (N_4280,N_2797,N_2479);
nor U4281 (N_4281,N_2324,N_2368);
nand U4282 (N_4282,N_1843,N_1634);
or U4283 (N_4283,N_2305,N_1714);
xor U4284 (N_4284,N_2479,N_2883);
nor U4285 (N_4285,N_1720,N_2422);
or U4286 (N_4286,N_1549,N_2494);
nor U4287 (N_4287,N_1889,N_1970);
or U4288 (N_4288,N_1564,N_2587);
nor U4289 (N_4289,N_2021,N_2213);
xnor U4290 (N_4290,N_1713,N_2977);
and U4291 (N_4291,N_2542,N_1553);
and U4292 (N_4292,N_2395,N_2682);
nor U4293 (N_4293,N_1906,N_2639);
and U4294 (N_4294,N_2460,N_1897);
nand U4295 (N_4295,N_2301,N_2405);
or U4296 (N_4296,N_2662,N_1778);
and U4297 (N_4297,N_1867,N_2759);
xnor U4298 (N_4298,N_2458,N_2870);
nor U4299 (N_4299,N_2985,N_2480);
nand U4300 (N_4300,N_2696,N_2556);
xnor U4301 (N_4301,N_2479,N_2483);
xnor U4302 (N_4302,N_1504,N_2827);
nand U4303 (N_4303,N_2180,N_2024);
nor U4304 (N_4304,N_1624,N_1597);
or U4305 (N_4305,N_2291,N_2777);
and U4306 (N_4306,N_1932,N_2226);
xor U4307 (N_4307,N_1548,N_1940);
nor U4308 (N_4308,N_2764,N_2585);
nand U4309 (N_4309,N_1864,N_2411);
xnor U4310 (N_4310,N_2013,N_2705);
nand U4311 (N_4311,N_2705,N_2089);
and U4312 (N_4312,N_2108,N_2930);
xor U4313 (N_4313,N_1730,N_2642);
nor U4314 (N_4314,N_2308,N_2883);
nand U4315 (N_4315,N_2625,N_2160);
xor U4316 (N_4316,N_1968,N_2596);
xnor U4317 (N_4317,N_1811,N_1506);
or U4318 (N_4318,N_1690,N_1610);
and U4319 (N_4319,N_2910,N_2268);
xnor U4320 (N_4320,N_2157,N_1847);
or U4321 (N_4321,N_1899,N_2372);
and U4322 (N_4322,N_2424,N_2914);
nand U4323 (N_4323,N_1882,N_1612);
nor U4324 (N_4324,N_2559,N_1586);
xor U4325 (N_4325,N_2387,N_2523);
nand U4326 (N_4326,N_2788,N_2674);
and U4327 (N_4327,N_1872,N_2118);
nor U4328 (N_4328,N_2473,N_2090);
xnor U4329 (N_4329,N_2859,N_2791);
nor U4330 (N_4330,N_1782,N_2656);
nor U4331 (N_4331,N_2180,N_1873);
nor U4332 (N_4332,N_2359,N_2867);
nand U4333 (N_4333,N_1557,N_2275);
nand U4334 (N_4334,N_1766,N_2563);
or U4335 (N_4335,N_2476,N_2473);
and U4336 (N_4336,N_1557,N_1654);
or U4337 (N_4337,N_2150,N_2026);
or U4338 (N_4338,N_2966,N_2684);
nor U4339 (N_4339,N_2238,N_2964);
nand U4340 (N_4340,N_2335,N_2168);
xor U4341 (N_4341,N_1529,N_1952);
xor U4342 (N_4342,N_2380,N_2320);
nor U4343 (N_4343,N_2303,N_1914);
xnor U4344 (N_4344,N_2368,N_1503);
xor U4345 (N_4345,N_2444,N_1692);
nand U4346 (N_4346,N_1564,N_2839);
and U4347 (N_4347,N_1817,N_1574);
nand U4348 (N_4348,N_1564,N_1867);
nand U4349 (N_4349,N_2358,N_1647);
nand U4350 (N_4350,N_2408,N_2097);
nor U4351 (N_4351,N_2420,N_2536);
nand U4352 (N_4352,N_1513,N_2402);
nor U4353 (N_4353,N_2413,N_2394);
nor U4354 (N_4354,N_2412,N_2866);
nor U4355 (N_4355,N_2696,N_2769);
nand U4356 (N_4356,N_2930,N_2439);
nand U4357 (N_4357,N_1957,N_1837);
or U4358 (N_4358,N_1632,N_2046);
nand U4359 (N_4359,N_2498,N_2517);
or U4360 (N_4360,N_1788,N_1675);
or U4361 (N_4361,N_2427,N_1604);
and U4362 (N_4362,N_2805,N_2451);
nor U4363 (N_4363,N_1939,N_1925);
xnor U4364 (N_4364,N_2014,N_1632);
nand U4365 (N_4365,N_2050,N_2878);
nor U4366 (N_4366,N_2458,N_2095);
xnor U4367 (N_4367,N_2063,N_2180);
xnor U4368 (N_4368,N_2871,N_1501);
nor U4369 (N_4369,N_2271,N_1849);
or U4370 (N_4370,N_2833,N_2061);
xnor U4371 (N_4371,N_2401,N_2267);
or U4372 (N_4372,N_2422,N_1807);
or U4373 (N_4373,N_2692,N_2616);
and U4374 (N_4374,N_2423,N_1948);
nand U4375 (N_4375,N_2500,N_2277);
or U4376 (N_4376,N_2697,N_2237);
nor U4377 (N_4377,N_1653,N_2889);
or U4378 (N_4378,N_2476,N_2328);
nand U4379 (N_4379,N_1550,N_2666);
nand U4380 (N_4380,N_2445,N_2449);
or U4381 (N_4381,N_2325,N_2099);
xor U4382 (N_4382,N_2385,N_1873);
nor U4383 (N_4383,N_2016,N_2937);
and U4384 (N_4384,N_2411,N_2481);
or U4385 (N_4385,N_1987,N_1961);
nand U4386 (N_4386,N_2665,N_2574);
nor U4387 (N_4387,N_1878,N_1947);
nand U4388 (N_4388,N_1907,N_2068);
xor U4389 (N_4389,N_1739,N_2029);
or U4390 (N_4390,N_1833,N_1548);
xor U4391 (N_4391,N_2155,N_2247);
and U4392 (N_4392,N_2488,N_1849);
or U4393 (N_4393,N_2864,N_1725);
xor U4394 (N_4394,N_1637,N_2201);
nor U4395 (N_4395,N_2868,N_2408);
or U4396 (N_4396,N_1503,N_2246);
xnor U4397 (N_4397,N_1756,N_2502);
and U4398 (N_4398,N_2001,N_2498);
nor U4399 (N_4399,N_2816,N_1722);
and U4400 (N_4400,N_1501,N_2245);
or U4401 (N_4401,N_1705,N_1852);
xnor U4402 (N_4402,N_2826,N_2375);
nand U4403 (N_4403,N_2544,N_2798);
or U4404 (N_4404,N_1830,N_2546);
nand U4405 (N_4405,N_2913,N_2175);
xor U4406 (N_4406,N_2735,N_1674);
nand U4407 (N_4407,N_2605,N_2915);
nand U4408 (N_4408,N_2920,N_1930);
or U4409 (N_4409,N_2631,N_2488);
nand U4410 (N_4410,N_2829,N_2496);
nor U4411 (N_4411,N_2695,N_2276);
or U4412 (N_4412,N_2219,N_2128);
or U4413 (N_4413,N_2570,N_2782);
nand U4414 (N_4414,N_1778,N_2911);
xor U4415 (N_4415,N_2524,N_2914);
nand U4416 (N_4416,N_2561,N_1816);
or U4417 (N_4417,N_2645,N_2439);
and U4418 (N_4418,N_2388,N_1668);
xor U4419 (N_4419,N_2278,N_2409);
xor U4420 (N_4420,N_1686,N_2149);
or U4421 (N_4421,N_2162,N_1504);
nand U4422 (N_4422,N_2245,N_1950);
or U4423 (N_4423,N_2398,N_2356);
nor U4424 (N_4424,N_1749,N_2191);
xor U4425 (N_4425,N_2674,N_2245);
nand U4426 (N_4426,N_2556,N_2866);
nor U4427 (N_4427,N_1580,N_2324);
nor U4428 (N_4428,N_2954,N_2204);
xnor U4429 (N_4429,N_1758,N_2125);
or U4430 (N_4430,N_2224,N_2181);
and U4431 (N_4431,N_2076,N_1693);
nor U4432 (N_4432,N_2272,N_1899);
or U4433 (N_4433,N_1922,N_1774);
nand U4434 (N_4434,N_1790,N_1910);
nand U4435 (N_4435,N_1949,N_2451);
nand U4436 (N_4436,N_2908,N_1998);
or U4437 (N_4437,N_2030,N_2720);
or U4438 (N_4438,N_1908,N_2330);
nand U4439 (N_4439,N_1901,N_2208);
nor U4440 (N_4440,N_2478,N_2596);
or U4441 (N_4441,N_1695,N_2121);
nor U4442 (N_4442,N_1506,N_2874);
and U4443 (N_4443,N_2394,N_2120);
and U4444 (N_4444,N_2047,N_2417);
nor U4445 (N_4445,N_2868,N_2066);
nor U4446 (N_4446,N_2483,N_2901);
and U4447 (N_4447,N_2128,N_1866);
xnor U4448 (N_4448,N_2938,N_2893);
nand U4449 (N_4449,N_2358,N_1880);
and U4450 (N_4450,N_2650,N_2409);
or U4451 (N_4451,N_2789,N_1588);
nor U4452 (N_4452,N_2696,N_2540);
nand U4453 (N_4453,N_2331,N_2109);
or U4454 (N_4454,N_2722,N_1930);
nor U4455 (N_4455,N_2702,N_2478);
nand U4456 (N_4456,N_1831,N_1877);
nand U4457 (N_4457,N_2147,N_2842);
or U4458 (N_4458,N_1534,N_1821);
nand U4459 (N_4459,N_2260,N_2490);
nor U4460 (N_4460,N_2882,N_2059);
xnor U4461 (N_4461,N_1994,N_2309);
and U4462 (N_4462,N_2549,N_2527);
xor U4463 (N_4463,N_1681,N_2597);
nand U4464 (N_4464,N_2045,N_1866);
xnor U4465 (N_4465,N_1919,N_2779);
nand U4466 (N_4466,N_2438,N_1661);
xor U4467 (N_4467,N_2198,N_1749);
or U4468 (N_4468,N_1642,N_2301);
nand U4469 (N_4469,N_2092,N_1721);
or U4470 (N_4470,N_2805,N_1536);
nand U4471 (N_4471,N_1729,N_2915);
nand U4472 (N_4472,N_2934,N_1777);
xnor U4473 (N_4473,N_2668,N_2357);
nor U4474 (N_4474,N_2407,N_1708);
nor U4475 (N_4475,N_1934,N_1885);
and U4476 (N_4476,N_2982,N_2424);
nand U4477 (N_4477,N_2099,N_1608);
or U4478 (N_4478,N_2405,N_1572);
nand U4479 (N_4479,N_1837,N_2509);
nand U4480 (N_4480,N_1595,N_2659);
nand U4481 (N_4481,N_2096,N_2652);
nor U4482 (N_4482,N_2418,N_2465);
nor U4483 (N_4483,N_1638,N_2841);
or U4484 (N_4484,N_2375,N_2782);
or U4485 (N_4485,N_1908,N_1581);
and U4486 (N_4486,N_2544,N_1938);
or U4487 (N_4487,N_1784,N_2977);
and U4488 (N_4488,N_1819,N_2297);
nand U4489 (N_4489,N_2347,N_1964);
or U4490 (N_4490,N_2787,N_2760);
nand U4491 (N_4491,N_2255,N_2262);
and U4492 (N_4492,N_2050,N_1593);
nor U4493 (N_4493,N_2811,N_2564);
nand U4494 (N_4494,N_2611,N_2160);
or U4495 (N_4495,N_2565,N_2361);
or U4496 (N_4496,N_2252,N_2064);
and U4497 (N_4497,N_2946,N_2064);
nor U4498 (N_4498,N_2650,N_1951);
or U4499 (N_4499,N_1921,N_2054);
nand U4500 (N_4500,N_4064,N_3706);
xnor U4501 (N_4501,N_4248,N_3562);
or U4502 (N_4502,N_3202,N_4134);
xnor U4503 (N_4503,N_3187,N_3621);
nor U4504 (N_4504,N_4012,N_3399);
xor U4505 (N_4505,N_3849,N_3191);
nor U4506 (N_4506,N_3766,N_3939);
xnor U4507 (N_4507,N_3943,N_3027);
or U4508 (N_4508,N_4094,N_3079);
xnor U4509 (N_4509,N_3244,N_3790);
or U4510 (N_4510,N_3061,N_3959);
nor U4511 (N_4511,N_3686,N_3398);
nand U4512 (N_4512,N_3291,N_3070);
nand U4513 (N_4513,N_4379,N_4242);
xnor U4514 (N_4514,N_4418,N_4149);
nand U4515 (N_4515,N_4068,N_3835);
xnor U4516 (N_4516,N_4048,N_3991);
nor U4517 (N_4517,N_3372,N_3629);
xor U4518 (N_4518,N_4090,N_3103);
xor U4519 (N_4519,N_3317,N_3687);
nand U4520 (N_4520,N_3446,N_4320);
nor U4521 (N_4521,N_3014,N_4361);
and U4522 (N_4522,N_3853,N_3262);
and U4523 (N_4523,N_3247,N_3513);
xnor U4524 (N_4524,N_3593,N_3985);
or U4525 (N_4525,N_3293,N_3421);
xor U4526 (N_4526,N_3833,N_3370);
xnor U4527 (N_4527,N_4011,N_3213);
xnor U4528 (N_4528,N_3577,N_4436);
or U4529 (N_4529,N_4474,N_3888);
nand U4530 (N_4530,N_3277,N_3723);
xor U4531 (N_4531,N_4319,N_4328);
nand U4532 (N_4532,N_4194,N_3366);
nand U4533 (N_4533,N_3565,N_3970);
xor U4534 (N_4534,N_3796,N_4443);
nand U4535 (N_4535,N_3854,N_3894);
and U4536 (N_4536,N_3900,N_3307);
xnor U4537 (N_4537,N_4218,N_3615);
or U4538 (N_4538,N_3937,N_3818);
xor U4539 (N_4539,N_3042,N_3223);
nor U4540 (N_4540,N_3949,N_3329);
xor U4541 (N_4541,N_3024,N_3148);
or U4542 (N_4542,N_3510,N_3531);
nor U4543 (N_4543,N_3073,N_4386);
nand U4544 (N_4544,N_3331,N_3804);
xor U4545 (N_4545,N_3207,N_4482);
xor U4546 (N_4546,N_3282,N_3936);
or U4547 (N_4547,N_3311,N_3769);
xnor U4548 (N_4548,N_3603,N_4397);
or U4549 (N_4549,N_3000,N_3381);
xor U4550 (N_4550,N_4465,N_3994);
nor U4551 (N_4551,N_3914,N_4112);
nand U4552 (N_4552,N_3590,N_3816);
nand U4553 (N_4553,N_3437,N_4026);
xor U4554 (N_4554,N_3261,N_4055);
xnor U4555 (N_4555,N_4051,N_4305);
and U4556 (N_4556,N_3647,N_3623);
and U4557 (N_4557,N_3895,N_3805);
xnor U4558 (N_4558,N_3258,N_3239);
and U4559 (N_4559,N_4342,N_3685);
xnor U4560 (N_4560,N_3928,N_4128);
and U4561 (N_4561,N_4229,N_4143);
and U4562 (N_4562,N_3459,N_3434);
xor U4563 (N_4563,N_3691,N_3762);
or U4564 (N_4564,N_4494,N_4476);
and U4565 (N_4565,N_3431,N_3375);
and U4566 (N_4566,N_3419,N_3741);
nor U4567 (N_4567,N_3166,N_3747);
nand U4568 (N_4568,N_3916,N_3338);
or U4569 (N_4569,N_4122,N_3897);
nor U4570 (N_4570,N_4306,N_3442);
nand U4571 (N_4571,N_3496,N_3764);
nand U4572 (N_4572,N_4266,N_4419);
xnor U4573 (N_4573,N_3783,N_3554);
and U4574 (N_4574,N_3905,N_4299);
xnor U4575 (N_4575,N_4261,N_3140);
nor U4576 (N_4576,N_3463,N_4017);
and U4577 (N_4577,N_3144,N_4363);
and U4578 (N_4578,N_3093,N_4167);
nor U4579 (N_4579,N_3389,N_3773);
nand U4580 (N_4580,N_4072,N_3280);
xnor U4581 (N_4581,N_3142,N_4303);
or U4582 (N_4582,N_3618,N_4097);
nor U4583 (N_4583,N_3569,N_3659);
and U4584 (N_4584,N_3848,N_3713);
xor U4585 (N_4585,N_3504,N_3004);
and U4586 (N_4586,N_3979,N_4276);
and U4587 (N_4587,N_3988,N_3272);
and U4588 (N_4588,N_3230,N_3392);
or U4589 (N_4589,N_3344,N_4224);
and U4590 (N_4590,N_3581,N_3602);
nand U4591 (N_4591,N_4080,N_3776);
nor U4592 (N_4592,N_3246,N_3479);
nor U4593 (N_4593,N_3234,N_3677);
or U4594 (N_4594,N_4425,N_3081);
and U4595 (N_4595,N_3164,N_3981);
or U4596 (N_4596,N_3114,N_3923);
and U4597 (N_4597,N_3591,N_3715);
and U4598 (N_4598,N_3248,N_3967);
and U4599 (N_4599,N_4413,N_3826);
nand U4600 (N_4600,N_3688,N_3975);
and U4601 (N_4601,N_4415,N_4073);
or U4602 (N_4602,N_4344,N_3394);
and U4603 (N_4603,N_3101,N_3057);
or U4604 (N_4604,N_4434,N_4357);
nand U4605 (N_4605,N_4467,N_3236);
xnor U4606 (N_4606,N_4478,N_3913);
nand U4607 (N_4607,N_3034,N_3544);
nor U4608 (N_4608,N_3535,N_4354);
or U4609 (N_4609,N_4005,N_4001);
nand U4610 (N_4610,N_4211,N_3794);
and U4611 (N_4611,N_3995,N_3782);
nor U4612 (N_4612,N_3726,N_3342);
xnor U4613 (N_4613,N_4416,N_4286);
and U4614 (N_4614,N_4041,N_3182);
nand U4615 (N_4615,N_3346,N_3099);
or U4616 (N_4616,N_3767,N_3567);
xnor U4617 (N_4617,N_3238,N_4377);
nand U4618 (N_4618,N_3638,N_3092);
nand U4619 (N_4619,N_3443,N_3786);
and U4620 (N_4620,N_4222,N_4235);
and U4621 (N_4621,N_3732,N_3210);
or U4622 (N_4622,N_3200,N_4269);
and U4623 (N_4623,N_3058,N_4157);
nor U4624 (N_4624,N_3157,N_3502);
xnor U4625 (N_4625,N_3118,N_3596);
or U4626 (N_4626,N_4083,N_3938);
or U4627 (N_4627,N_3199,N_3422);
xnor U4628 (N_4628,N_3522,N_3139);
nor U4629 (N_4629,N_3226,N_3951);
nor U4630 (N_4630,N_4085,N_3185);
and U4631 (N_4631,N_3473,N_3644);
xor U4632 (N_4632,N_3495,N_4495);
nand U4633 (N_4633,N_4454,N_4390);
nand U4634 (N_4634,N_3214,N_3992);
nand U4635 (N_4635,N_4160,N_4069);
nand U4636 (N_4636,N_3054,N_3974);
or U4637 (N_4637,N_4039,N_4233);
nand U4638 (N_4638,N_3456,N_3254);
and U4639 (N_4639,N_3115,N_3879);
nor U4640 (N_4640,N_4100,N_3430);
nor U4641 (N_4641,N_3983,N_3286);
and U4642 (N_4642,N_3952,N_3874);
nand U4643 (N_4643,N_3806,N_3085);
nor U4644 (N_4644,N_3126,N_4408);
nand U4645 (N_4645,N_3450,N_4325);
nand U4646 (N_4646,N_3256,N_4023);
nor U4647 (N_4647,N_4278,N_3306);
nor U4648 (N_4648,N_3511,N_4115);
and U4649 (N_4649,N_3128,N_3961);
nor U4650 (N_4650,N_3362,N_3401);
nand U4651 (N_4651,N_3650,N_3597);
xor U4652 (N_4652,N_3505,N_4384);
nor U4653 (N_4653,N_4183,N_4322);
xnor U4654 (N_4654,N_4053,N_3160);
nand U4655 (N_4655,N_4368,N_4430);
xnor U4656 (N_4656,N_3781,N_3812);
xnor U4657 (N_4657,N_4030,N_4163);
xnor U4658 (N_4658,N_3984,N_3083);
xor U4659 (N_4659,N_4166,N_3919);
nor U4660 (N_4660,N_3670,N_3449);
or U4661 (N_4661,N_3801,N_3009);
nor U4662 (N_4662,N_3302,N_3924);
nor U4663 (N_4663,N_4290,N_3725);
nand U4664 (N_4664,N_3964,N_3557);
or U4665 (N_4665,N_3673,N_4236);
nand U4666 (N_4666,N_3067,N_3015);
xnor U4667 (N_4667,N_4140,N_3233);
xnor U4668 (N_4668,N_3156,N_3656);
nand U4669 (N_4669,N_3893,N_4404);
nor U4670 (N_4670,N_3588,N_3270);
or U4671 (N_4671,N_4479,N_3066);
or U4672 (N_4672,N_3339,N_3183);
nand U4673 (N_4673,N_4161,N_4417);
nand U4674 (N_4674,N_3595,N_4285);
and U4675 (N_4675,N_4054,N_4293);
or U4676 (N_4676,N_4282,N_3123);
or U4677 (N_4677,N_3111,N_3386);
xor U4678 (N_4678,N_3509,N_4096);
nor U4679 (N_4679,N_3840,N_4182);
nor U4680 (N_4680,N_3468,N_4451);
or U4681 (N_4681,N_3538,N_3636);
nand U4682 (N_4682,N_3356,N_4447);
nand U4683 (N_4683,N_4395,N_3359);
nor U4684 (N_4684,N_3100,N_3284);
nand U4685 (N_4685,N_3521,N_3477);
xnor U4686 (N_4686,N_3935,N_3530);
and U4687 (N_4687,N_3860,N_4153);
and U4688 (N_4688,N_4027,N_3989);
xnor U4689 (N_4689,N_4437,N_4444);
nor U4690 (N_4690,N_4156,N_4273);
nor U4691 (N_4691,N_4152,N_3627);
and U4692 (N_4692,N_4237,N_3669);
nand U4693 (N_4693,N_3318,N_4093);
or U4694 (N_4694,N_4216,N_3822);
and U4695 (N_4695,N_3872,N_4065);
xor U4696 (N_4696,N_3520,N_4170);
or U4697 (N_4697,N_4297,N_3471);
or U4698 (N_4698,N_3195,N_3945);
or U4699 (N_4699,N_4389,N_4412);
nor U4700 (N_4700,N_3586,N_3391);
nor U4701 (N_4701,N_3635,N_3696);
or U4702 (N_4702,N_4117,N_4088);
nor U4703 (N_4703,N_3850,N_4374);
or U4704 (N_4704,N_3060,N_4061);
nor U4705 (N_4705,N_4022,N_3580);
and U4706 (N_4706,N_3499,N_4459);
or U4707 (N_4707,N_3445,N_3416);
or U4708 (N_4708,N_3163,N_4378);
nand U4709 (N_4709,N_4142,N_3149);
nor U4710 (N_4710,N_3841,N_3962);
or U4711 (N_4711,N_4025,N_4199);
and U4712 (N_4712,N_3043,N_4330);
nor U4713 (N_4713,N_3006,N_3420);
or U4714 (N_4714,N_3205,N_3097);
xor U4715 (N_4715,N_3326,N_4365);
xnor U4716 (N_4716,N_3825,N_3551);
xor U4717 (N_4717,N_3710,N_3536);
nor U4718 (N_4718,N_4456,N_3954);
nor U4719 (N_4719,N_3579,N_3718);
nand U4720 (N_4720,N_3982,N_3216);
xor U4721 (N_4721,N_3201,N_4168);
nand U4722 (N_4722,N_4099,N_3347);
nand U4723 (N_4723,N_3168,N_4340);
nor U4724 (N_4724,N_3411,N_3241);
nor U4725 (N_4725,N_4207,N_3613);
and U4726 (N_4726,N_4174,N_4289);
or U4727 (N_4727,N_4021,N_4145);
nand U4728 (N_4728,N_4388,N_4105);
nor U4729 (N_4729,N_3907,N_3929);
xnor U4730 (N_4730,N_4079,N_3720);
or U4731 (N_4731,N_3451,N_3151);
or U4732 (N_4732,N_3396,N_4359);
nand U4733 (N_4733,N_4280,N_4497);
nor U4734 (N_4734,N_3646,N_3374);
or U4735 (N_4735,N_3039,N_3751);
or U4736 (N_4736,N_3815,N_3921);
or U4737 (N_4737,N_4438,N_4150);
and U4738 (N_4738,N_3512,N_3315);
xnor U4739 (N_4739,N_4204,N_4159);
nor U4740 (N_4740,N_3357,N_3566);
nand U4741 (N_4741,N_4274,N_3665);
nand U4742 (N_4742,N_4126,N_4243);
and U4743 (N_4743,N_4087,N_4268);
xnor U4744 (N_4744,N_3748,N_4104);
or U4745 (N_4745,N_3859,N_3999);
nand U4746 (N_4746,N_4110,N_3458);
and U4747 (N_4747,N_3648,N_3768);
or U4748 (N_4748,N_3441,N_3727);
nand U4749 (N_4749,N_3683,N_3178);
xnor U4750 (N_4750,N_4037,N_3915);
nor U4751 (N_4751,N_3017,N_3548);
nand U4752 (N_4752,N_3948,N_3036);
nor U4753 (N_4753,N_3448,N_3264);
or U4754 (N_4754,N_3425,N_4406);
xor U4755 (N_4755,N_4256,N_3209);
and U4756 (N_4756,N_3532,N_4349);
and U4757 (N_4757,N_3145,N_3162);
nand U4758 (N_4758,N_4129,N_3436);
nand U4759 (N_4759,N_3795,N_3129);
and U4760 (N_4760,N_3652,N_3528);
or U4761 (N_4761,N_3255,N_3486);
nor U4762 (N_4762,N_4433,N_3570);
and U4763 (N_4763,N_3604,N_3744);
or U4764 (N_4764,N_3367,N_3224);
or U4765 (N_4765,N_4071,N_3953);
nor U4766 (N_4766,N_3404,N_4116);
xnor U4767 (N_4767,N_3865,N_4314);
nor U4768 (N_4768,N_4018,N_3784);
nand U4769 (N_4769,N_3384,N_3563);
and U4770 (N_4770,N_3671,N_3432);
and U4771 (N_4771,N_4492,N_4114);
or U4772 (N_4772,N_3467,N_3552);
nor U4773 (N_4773,N_3814,N_4082);
nor U4774 (N_4774,N_3492,N_3464);
and U4775 (N_4775,N_4288,N_3716);
and U4776 (N_4776,N_4351,N_4189);
xnor U4777 (N_4777,N_3639,N_4309);
and U4778 (N_4778,N_4202,N_3881);
xor U4779 (N_4779,N_3925,N_3809);
and U4780 (N_4780,N_4227,N_3104);
nand U4781 (N_4781,N_4475,N_3122);
nand U4782 (N_4782,N_3909,N_4154);
xnor U4783 (N_4783,N_3288,N_3908);
or U4784 (N_4784,N_3082,N_3676);
xor U4785 (N_4785,N_4184,N_3250);
nand U4786 (N_4786,N_3827,N_3189);
nor U4787 (N_4787,N_3780,N_3480);
and U4788 (N_4788,N_4032,N_3271);
xnor U4789 (N_4789,N_4074,N_4164);
nand U4790 (N_4790,N_4486,N_3173);
or U4791 (N_4791,N_4367,N_3294);
and U4792 (N_4792,N_4015,N_3197);
and U4793 (N_4793,N_3007,N_4151);
nand U4794 (N_4794,N_3630,N_3931);
nand U4795 (N_4795,N_3598,N_3235);
xor U4796 (N_4796,N_3211,N_3987);
and U4797 (N_4797,N_3086,N_4132);
xnor U4798 (N_4798,N_3774,N_3911);
and U4799 (N_4799,N_4135,N_3488);
or U4800 (N_4800,N_3033,N_3300);
xnor U4801 (N_4801,N_3472,N_3730);
xnor U4802 (N_4802,N_4366,N_4180);
or U4803 (N_4803,N_3503,N_3312);
and U4804 (N_4804,N_3887,N_3228);
and U4805 (N_4805,N_3065,N_4327);
and U4806 (N_4806,N_3153,N_4369);
nand U4807 (N_4807,N_3864,N_4162);
xnor U4808 (N_4808,N_3240,N_3143);
xnor U4809 (N_4809,N_4356,N_3429);
or U4810 (N_4810,N_3475,N_3666);
xor U4811 (N_4811,N_3966,N_4258);
and U4812 (N_4812,N_3899,N_3029);
or U4813 (N_4813,N_3765,N_3056);
nand U4814 (N_4814,N_3252,N_4217);
and U4815 (N_4815,N_3942,N_3851);
nor U4816 (N_4816,N_4337,N_3680);
nand U4817 (N_4817,N_4040,N_3986);
or U4818 (N_4818,N_3047,N_4343);
or U4819 (N_4819,N_3243,N_3158);
and U4820 (N_4820,N_3839,N_3515);
xnor U4821 (N_4821,N_3799,N_3349);
xor U4822 (N_4822,N_4047,N_4178);
nand U4823 (N_4823,N_3048,N_4453);
and U4824 (N_4824,N_3117,N_4181);
or U4825 (N_4825,N_3316,N_4480);
and U4826 (N_4826,N_3365,N_4370);
xor U4827 (N_4827,N_4341,N_3251);
nor U4828 (N_4828,N_3090,N_4197);
or U4829 (N_4829,N_3525,N_4446);
nor U4830 (N_4830,N_3692,N_3491);
nor U4831 (N_4831,N_4423,N_4491);
xor U4832 (N_4832,N_4392,N_3757);
nand U4833 (N_4833,N_4414,N_3275);
nor U4834 (N_4834,N_4426,N_3049);
xnor U4835 (N_4835,N_4372,N_4277);
nor U4836 (N_4836,N_3550,N_3655);
xor U4837 (N_4837,N_3700,N_4429);
xor U4838 (N_4838,N_3704,N_4008);
and U4839 (N_4839,N_4002,N_3778);
nor U4840 (N_4840,N_3354,N_4043);
and U4841 (N_4841,N_3703,N_3611);
nand U4842 (N_4842,N_3754,N_3119);
or U4843 (N_4843,N_3478,N_3867);
nor U4844 (N_4844,N_3672,N_3605);
nor U4845 (N_4845,N_3011,N_3824);
or U4846 (N_4846,N_4028,N_3559);
nand U4847 (N_4847,N_3423,N_4111);
nand U4848 (N_4848,N_3435,N_3977);
and U4849 (N_4849,N_3958,N_3089);
or U4850 (N_4850,N_4488,N_3461);
or U4851 (N_4851,N_4308,N_3273);
or U4852 (N_4852,N_3549,N_3797);
xor U4853 (N_4853,N_3956,N_4226);
and U4854 (N_4854,N_3622,N_4493);
and U4855 (N_4855,N_4057,N_3946);
nor U4856 (N_4856,N_3320,N_3413);
and U4857 (N_4857,N_4472,N_4452);
nor U4858 (N_4858,N_3279,N_3679);
and U4859 (N_4859,N_4432,N_4448);
and U4860 (N_4860,N_3973,N_3555);
xor U4861 (N_4861,N_3681,N_3044);
nor U4862 (N_4862,N_3147,N_3188);
or U4863 (N_4863,N_4391,N_4399);
nor U4864 (N_4864,N_3689,N_3321);
xor U4865 (N_4865,N_4228,N_3771);
nor U4866 (N_4866,N_3912,N_3539);
nand U4867 (N_4867,N_3310,N_3607);
or U4868 (N_4868,N_3519,N_3287);
nand U4869 (N_4869,N_3524,N_3657);
xnor U4870 (N_4870,N_4352,N_3990);
or U4871 (N_4871,N_3625,N_4420);
nor U4872 (N_4872,N_3482,N_4136);
or U4873 (N_4873,N_3847,N_3740);
or U4874 (N_4874,N_3508,N_3245);
nor U4875 (N_4875,N_3745,N_4209);
nand U4876 (N_4876,N_4148,N_3332);
nor U4877 (N_4877,N_3364,N_3926);
and U4878 (N_4878,N_4307,N_3858);
and U4879 (N_4879,N_3308,N_3896);
nor U4880 (N_4880,N_3020,N_3628);
xnor U4881 (N_4881,N_4323,N_4364);
nor U4882 (N_4882,N_3976,N_4067);
and U4883 (N_4883,N_3106,N_4106);
xor U4884 (N_4884,N_3701,N_3828);
xor U4885 (N_4885,N_4254,N_3439);
xor U4886 (N_4886,N_4208,N_3968);
nand U4887 (N_4887,N_3032,N_3965);
xnor U4888 (N_4888,N_3172,N_3113);
xnor U4889 (N_4889,N_4007,N_4063);
nor U4890 (N_4890,N_4230,N_3871);
and U4891 (N_4891,N_4095,N_3587);
or U4892 (N_4892,N_3882,N_3832);
nand U4893 (N_4893,N_3335,N_4312);
nand U4894 (N_4894,N_3699,N_4487);
nor U4895 (N_4895,N_3843,N_3204);
and U4896 (N_4896,N_4101,N_3388);
nand U4897 (N_4897,N_4133,N_3534);
nand U4898 (N_4898,N_3176,N_3064);
or U4899 (N_4899,N_3373,N_3770);
nor U4900 (N_4900,N_4205,N_3772);
nand U4901 (N_4901,N_3878,N_3087);
xnor U4902 (N_4902,N_4201,N_3167);
nor U4903 (N_4903,N_3418,N_4144);
and U4904 (N_4904,N_3120,N_3444);
and U4905 (N_4905,N_4020,N_3409);
nand U4906 (N_4906,N_3787,N_4455);
nor U4907 (N_4907,N_4084,N_3884);
and U4908 (N_4908,N_4121,N_4427);
nand U4909 (N_4909,N_3325,N_3171);
and U4910 (N_4910,N_3417,N_3829);
nand U4911 (N_4911,N_4335,N_4260);
or U4912 (N_4912,N_3634,N_3074);
and U4913 (N_4913,N_3289,N_4287);
nor U4914 (N_4914,N_3452,N_4300);
xor U4915 (N_4915,N_3141,N_4270);
and U4916 (N_4916,N_3885,N_3363);
nor U4917 (N_4917,N_3266,N_4212);
nor U4918 (N_4918,N_4463,N_3855);
and U4919 (N_4919,N_3008,N_4283);
xnor U4920 (N_4920,N_3376,N_4203);
xnor U4921 (N_4921,N_4033,N_4234);
nand U4922 (N_4922,N_3576,N_3476);
or U4923 (N_4923,N_3572,N_3013);
xnor U4924 (N_4924,N_4498,N_4405);
or U4925 (N_4925,N_3010,N_3721);
or U4926 (N_4926,N_3174,N_3415);
xor U4927 (N_4927,N_3717,N_3866);
and U4928 (N_4928,N_3756,N_3078);
and U4929 (N_4929,N_3620,N_3337);
and U4930 (N_4930,N_3760,N_3127);
xnor U4931 (N_4931,N_3807,N_4141);
nand U4932 (N_4932,N_3574,N_4272);
xor U4933 (N_4933,N_3170,N_3695);
xnor U4934 (N_4934,N_4158,N_3379);
xor U4935 (N_4935,N_3132,N_3664);
nand U4936 (N_4936,N_4172,N_3800);
nor U4937 (N_4937,N_3177,N_3369);
xnor U4938 (N_4938,N_3138,N_3775);
nor U4939 (N_4939,N_4336,N_4462);
xnor U4940 (N_4940,N_4257,N_3594);
nor U4941 (N_4941,N_3406,N_3021);
xor U4942 (N_4942,N_4460,N_3296);
nor U4943 (N_4943,N_4241,N_4137);
nand U4944 (N_4944,N_3212,N_3257);
nand U4945 (N_4945,N_3403,N_3668);
or U4946 (N_4946,N_4296,N_4029);
xor U4947 (N_4947,N_4038,N_3722);
and U4948 (N_4948,N_3660,N_3405);
xor U4949 (N_4949,N_4059,N_3940);
xor U4950 (N_4950,N_4102,N_3324);
xor U4951 (N_4951,N_3454,N_3427);
nand U4952 (N_4952,N_4469,N_3457);
xor U4953 (N_4953,N_3996,N_3334);
and U4954 (N_4954,N_3408,N_3002);
and U4955 (N_4955,N_3410,N_4188);
nor U4956 (N_4956,N_3601,N_3742);
or U4957 (N_4957,N_3514,N_3393);
and U4958 (N_4958,N_3016,N_3096);
or U4959 (N_4959,N_3259,N_3050);
nand U4960 (N_4960,N_3616,N_3932);
nor U4961 (N_4961,N_4334,N_3281);
or U4962 (N_4962,N_3729,N_3875);
or U4963 (N_4963,N_4169,N_3371);
nand U4964 (N_4964,N_3221,N_3906);
and U4965 (N_4965,N_3584,N_4333);
and U4966 (N_4966,N_4393,N_4396);
or U4967 (N_4967,N_3861,N_4317);
or U4968 (N_4968,N_3035,N_3077);
or U4969 (N_4969,N_4206,N_3026);
nor U4970 (N_4970,N_3645,N_3803);
and U4971 (N_4971,N_3705,N_3165);
and U4972 (N_4972,N_4440,N_3998);
and U4973 (N_4973,N_3438,N_3877);
or U4974 (N_4974,N_4484,N_4249);
nor U4975 (N_4975,N_3819,N_4318);
nor U4976 (N_4976,N_3619,N_3215);
or U4977 (N_4977,N_3870,N_3440);
and U4978 (N_4978,N_4191,N_3462);
nor U4979 (N_4979,N_3301,N_3222);
and U4980 (N_4980,N_4441,N_3278);
or U4981 (N_4981,N_3135,N_4424);
nor U4982 (N_4982,N_3031,N_3972);
nand U4983 (N_4983,N_3059,N_3022);
nand U4984 (N_4984,N_3537,N_3390);
xor U4985 (N_4985,N_4014,N_3734);
nor U4986 (N_4986,N_4131,N_4113);
nand U4987 (N_4987,N_3930,N_3507);
nand U4988 (N_4988,N_4375,N_3319);
xnor U4989 (N_4989,N_3738,N_3227);
nor U4990 (N_4990,N_3746,N_3624);
or U4991 (N_4991,N_3269,N_3845);
nand U4992 (N_4992,N_4232,N_4003);
and U4993 (N_4993,N_3380,N_4401);
nor U4994 (N_4994,N_3052,N_4139);
nand U4995 (N_4995,N_4091,N_3978);
or U4996 (N_4996,N_3265,N_4383);
nand U4997 (N_4997,N_3218,N_3005);
nor U4998 (N_4998,N_3109,N_4109);
or U4999 (N_4999,N_3190,N_3553);
nand U5000 (N_5000,N_3133,N_3838);
and U5001 (N_5001,N_4400,N_4062);
nand U5002 (N_5002,N_3051,N_3283);
xor U5003 (N_5003,N_3322,N_3600);
and U5004 (N_5004,N_3728,N_3526);
and U5005 (N_5005,N_3546,N_4155);
nand U5006 (N_5006,N_4267,N_3733);
xnor U5007 (N_5007,N_3455,N_3368);
nor U5008 (N_5008,N_3348,N_3798);
nand U5009 (N_5009,N_4060,N_3927);
nand U5010 (N_5010,N_4264,N_4445);
and U5011 (N_5011,N_3116,N_3071);
and U5012 (N_5012,N_4442,N_4004);
xor U5013 (N_5013,N_3836,N_3080);
or U5014 (N_5014,N_4165,N_3934);
nand U5015 (N_5015,N_4049,N_3651);
xor U5016 (N_5016,N_3599,N_4086);
xnor U5017 (N_5017,N_3025,N_3180);
nor U5018 (N_5018,N_4213,N_3159);
and U5019 (N_5019,N_4496,N_3062);
or U5020 (N_5020,N_3161,N_3817);
and U5021 (N_5021,N_3285,N_3957);
nand U5022 (N_5022,N_3229,N_3353);
xor U5023 (N_5023,N_3395,N_3309);
nor U5024 (N_5024,N_3299,N_3217);
xor U5025 (N_5025,N_3274,N_3038);
and U5026 (N_5026,N_3340,N_3950);
or U5027 (N_5027,N_3447,N_4190);
nor U5028 (N_5028,N_3573,N_3753);
nor U5029 (N_5029,N_3714,N_3360);
and U5030 (N_5030,N_4292,N_3540);
and U5031 (N_5031,N_4016,N_3328);
and U5032 (N_5032,N_4031,N_3608);
xor U5033 (N_5033,N_4173,N_4410);
nand U5034 (N_5034,N_3575,N_3323);
xnor U5035 (N_5035,N_4045,N_3184);
nor U5036 (N_5036,N_4176,N_3175);
and U5037 (N_5037,N_3955,N_4120);
and U5038 (N_5038,N_3793,N_3045);
or U5039 (N_5039,N_3003,N_3527);
and U5040 (N_5040,N_4470,N_4119);
and U5041 (N_5041,N_4238,N_3313);
nand U5042 (N_5042,N_4489,N_3752);
or U5043 (N_5043,N_4245,N_4078);
nand U5044 (N_5044,N_3763,N_3698);
or U5045 (N_5045,N_4407,N_3856);
nand U5046 (N_5046,N_3568,N_3345);
xor U5047 (N_5047,N_3124,N_3397);
or U5048 (N_5048,N_3903,N_3028);
xnor U5049 (N_5049,N_4179,N_3831);
nand U5050 (N_5050,N_3892,N_3674);
or U5051 (N_5051,N_4473,N_3820);
and U5052 (N_5052,N_3529,N_3152);
nor U5053 (N_5053,N_3469,N_3470);
xor U5054 (N_5054,N_3880,N_3969);
and U5055 (N_5055,N_3412,N_4066);
nor U5056 (N_5056,N_3154,N_3193);
nand U5057 (N_5057,N_4353,N_3290);
or U5058 (N_5058,N_3823,N_4411);
and U5059 (N_5059,N_4193,N_3414);
nand U5060 (N_5060,N_4124,N_3474);
nor U5061 (N_5061,N_3206,N_3571);
and U5062 (N_5062,N_4477,N_4376);
nand U5063 (N_5063,N_3361,N_3902);
xnor U5064 (N_5064,N_3697,N_4373);
and U5065 (N_5065,N_4221,N_4275);
and U5066 (N_5066,N_4439,N_4219);
or U5067 (N_5067,N_4409,N_3917);
nor U5068 (N_5068,N_4302,N_3098);
xnor U5069 (N_5069,N_3702,N_4471);
nand U5070 (N_5070,N_3019,N_4313);
nand U5071 (N_5071,N_3707,N_4316);
xor U5072 (N_5072,N_3219,N_3383);
xnor U5073 (N_5073,N_3351,N_3237);
xor U5074 (N_5074,N_4326,N_3102);
and U5075 (N_5075,N_4259,N_3869);
and U5076 (N_5076,N_3327,N_3517);
or U5077 (N_5077,N_4225,N_3134);
or U5078 (N_5078,N_3336,N_3500);
or U5079 (N_5079,N_3933,N_3684);
or U5080 (N_5080,N_3131,N_3493);
and U5081 (N_5081,N_3426,N_3993);
nand U5082 (N_5082,N_3709,N_3155);
nor U5083 (N_5083,N_3378,N_3494);
xnor U5084 (N_5084,N_4294,N_3297);
nand U5085 (N_5085,N_3352,N_3641);
and U5086 (N_5086,N_3001,N_3084);
nand U5087 (N_5087,N_3407,N_3343);
or U5088 (N_5088,N_3263,N_3095);
nor U5089 (N_5089,N_4187,N_3750);
or U5090 (N_5090,N_4329,N_4428);
and U5091 (N_5091,N_4394,N_4358);
or U5092 (N_5092,N_4009,N_3711);
and U5093 (N_5093,N_3759,N_4291);
and U5094 (N_5094,N_4077,N_3292);
and U5095 (N_5095,N_4092,N_4252);
or U5096 (N_5096,N_4019,N_4422);
nor U5097 (N_5097,N_3811,N_3506);
nand U5098 (N_5098,N_4362,N_3901);
nor U5099 (N_5099,N_3041,N_4147);
and U5100 (N_5100,N_3108,N_3481);
and U5101 (N_5101,N_4089,N_3886);
and U5102 (N_5102,N_3944,N_4196);
nand U5103 (N_5103,N_3545,N_3941);
xor U5104 (N_5104,N_3487,N_3658);
nand U5105 (N_5105,N_3424,N_4271);
nor U5106 (N_5106,N_3792,N_4046);
nor U5107 (N_5107,N_4118,N_3739);
xnor U5108 (N_5108,N_3076,N_4464);
xor U5109 (N_5109,N_3873,N_3068);
xor U5110 (N_5110,N_3072,N_4371);
or U5111 (N_5111,N_3125,N_3146);
or U5112 (N_5112,N_4075,N_3400);
or U5113 (N_5113,N_3889,N_3791);
and U5114 (N_5114,N_3558,N_4251);
or U5115 (N_5115,N_3678,N_3136);
nand U5116 (N_5116,N_4355,N_3891);
or U5117 (N_5117,N_4103,N_3643);
nand U5118 (N_5118,N_4081,N_3963);
nand U5119 (N_5119,N_3305,N_3761);
nor U5120 (N_5120,N_3382,N_3631);
or U5121 (N_5121,N_3063,N_3260);
nand U5122 (N_5122,N_3564,N_3377);
nand U5123 (N_5123,N_4177,N_3040);
or U5124 (N_5124,N_3708,N_3533);
nand U5125 (N_5125,N_3560,N_3249);
and U5126 (N_5126,N_3834,N_3225);
and U5127 (N_5127,N_3314,N_4403);
or U5128 (N_5128,N_3821,N_4450);
or U5129 (N_5129,N_3466,N_4056);
or U5130 (N_5130,N_3330,N_3654);
and U5131 (N_5131,N_3743,N_3661);
and U5132 (N_5132,N_4130,N_4311);
xor U5133 (N_5133,N_3069,N_3107);
nor U5134 (N_5134,N_4315,N_3186);
xor U5135 (N_5135,N_3585,N_3662);
or U5136 (N_5136,N_3682,N_4058);
nor U5137 (N_5137,N_3387,N_3497);
and U5138 (N_5138,N_3541,N_3298);
nand U5139 (N_5139,N_3304,N_4381);
nor U5140 (N_5140,N_3295,N_3920);
nand U5141 (N_5141,N_4138,N_4398);
or U5142 (N_5142,N_3460,N_3606);
or U5143 (N_5143,N_3578,N_3355);
or U5144 (N_5144,N_4006,N_3789);
or U5145 (N_5145,N_4402,N_3485);
and U5146 (N_5146,N_3501,N_3582);
nor U5147 (N_5147,N_3971,N_3542);
or U5148 (N_5148,N_4431,N_3918);
nand U5149 (N_5149,N_4332,N_3137);
nor U5150 (N_5150,N_4490,N_4380);
and U5151 (N_5151,N_3633,N_3150);
xnor U5152 (N_5152,N_4263,N_3737);
nand U5153 (N_5153,N_3614,N_3023);
nand U5154 (N_5154,N_4024,N_4466);
nand U5155 (N_5155,N_3053,N_3253);
xor U5156 (N_5156,N_4215,N_3121);
nor U5157 (N_5157,N_4098,N_4345);
and U5158 (N_5158,N_4265,N_4347);
nand U5159 (N_5159,N_3960,N_3890);
or U5160 (N_5160,N_4339,N_4247);
nand U5161 (N_5161,N_3863,N_4304);
nand U5162 (N_5162,N_3922,N_4050);
or U5163 (N_5163,N_3402,N_3980);
or U5164 (N_5164,N_4298,N_3523);
and U5165 (N_5165,N_4295,N_3663);
and U5166 (N_5166,N_3724,N_4310);
nand U5167 (N_5167,N_4146,N_3232);
or U5168 (N_5168,N_4036,N_4192);
nor U5169 (N_5169,N_3637,N_4125);
nand U5170 (N_5170,N_3862,N_3198);
nor U5171 (N_5171,N_3267,N_4253);
xor U5172 (N_5172,N_4485,N_4240);
xor U5173 (N_5173,N_3842,N_4175);
nor U5174 (N_5174,N_3358,N_3012);
nor U5175 (N_5175,N_4035,N_3758);
and U5176 (N_5176,N_4499,N_4239);
or U5177 (N_5177,N_3675,N_3736);
nand U5178 (N_5178,N_4284,N_3231);
or U5179 (N_5179,N_3868,N_3626);
xnor U5180 (N_5180,N_3130,N_3112);
and U5181 (N_5181,N_4223,N_4070);
and U5182 (N_5182,N_4250,N_3208);
xnor U5183 (N_5183,N_3779,N_3876);
or U5184 (N_5184,N_3303,N_3904);
xnor U5185 (N_5185,N_4281,N_3883);
and U5186 (N_5186,N_3777,N_4052);
xnor U5187 (N_5187,N_4468,N_3690);
and U5188 (N_5188,N_4198,N_4244);
or U5189 (N_5189,N_4186,N_3749);
nor U5190 (N_5190,N_3813,N_3592);
nand U5191 (N_5191,N_4220,N_4458);
or U5192 (N_5192,N_3220,N_4481);
or U5193 (N_5193,N_3810,N_3242);
nand U5194 (N_5194,N_3612,N_3852);
nor U5195 (N_5195,N_4461,N_3997);
xnor U5196 (N_5196,N_3755,N_4000);
and U5197 (N_5197,N_3518,N_3632);
and U5198 (N_5198,N_3640,N_4185);
nor U5199 (N_5199,N_4200,N_4449);
nand U5200 (N_5200,N_4107,N_3785);
nor U5201 (N_5201,N_4123,N_3694);
xor U5202 (N_5202,N_3341,N_4044);
nand U5203 (N_5203,N_4385,N_4457);
or U5204 (N_5204,N_3898,N_4034);
nor U5205 (N_5205,N_3037,N_3385);
nand U5206 (N_5206,N_3428,N_3731);
nor U5207 (N_5207,N_3583,N_4210);
xnor U5208 (N_5208,N_3489,N_4483);
or U5209 (N_5209,N_4076,N_4387);
or U5210 (N_5210,N_4324,N_3617);
xnor U5211 (N_5211,N_4338,N_3030);
nand U5212 (N_5212,N_3091,N_3846);
nand U5213 (N_5213,N_3653,N_3808);
or U5214 (N_5214,N_4042,N_4421);
or U5215 (N_5215,N_4331,N_4382);
nor U5216 (N_5216,N_4246,N_4279);
and U5217 (N_5217,N_3333,N_3350);
and U5218 (N_5218,N_4346,N_3276);
and U5219 (N_5219,N_3837,N_3194);
nand U5220 (N_5220,N_3543,N_3649);
nand U5221 (N_5221,N_3094,N_3516);
nor U5222 (N_5222,N_3910,N_4348);
nor U5223 (N_5223,N_3018,N_3667);
xnor U5224 (N_5224,N_3105,N_4231);
nand U5225 (N_5225,N_3268,N_3196);
and U5226 (N_5226,N_3192,N_3498);
and U5227 (N_5227,N_4360,N_3203);
nor U5228 (N_5228,N_3719,N_3735);
and U5229 (N_5229,N_4321,N_4127);
and U5230 (N_5230,N_4435,N_3561);
or U5231 (N_5231,N_4108,N_3075);
nor U5232 (N_5232,N_3556,N_3169);
and U5233 (N_5233,N_3490,N_3547);
nor U5234 (N_5234,N_3642,N_3046);
nand U5235 (N_5235,N_3857,N_3484);
nand U5236 (N_5236,N_3465,N_3589);
xor U5237 (N_5237,N_4350,N_3788);
xnor U5238 (N_5238,N_3802,N_4255);
and U5239 (N_5239,N_3609,N_4010);
xor U5240 (N_5240,N_4262,N_3055);
nand U5241 (N_5241,N_4171,N_3088);
nor U5242 (N_5242,N_4301,N_3453);
xnor U5243 (N_5243,N_3693,N_4013);
nand U5244 (N_5244,N_3844,N_4214);
nand U5245 (N_5245,N_3179,N_3947);
xor U5246 (N_5246,N_4195,N_3830);
xor U5247 (N_5247,N_3610,N_3433);
nor U5248 (N_5248,N_3483,N_3110);
nor U5249 (N_5249,N_3712,N_3181);
nand U5250 (N_5250,N_3608,N_4244);
nor U5251 (N_5251,N_3450,N_3919);
and U5252 (N_5252,N_3798,N_3170);
nand U5253 (N_5253,N_4424,N_3345);
nand U5254 (N_5254,N_3459,N_4230);
nand U5255 (N_5255,N_4416,N_3589);
or U5256 (N_5256,N_3937,N_3995);
nand U5257 (N_5257,N_3756,N_3092);
or U5258 (N_5258,N_3587,N_3789);
nor U5259 (N_5259,N_3312,N_4359);
nor U5260 (N_5260,N_3541,N_3493);
or U5261 (N_5261,N_3352,N_4235);
nor U5262 (N_5262,N_3109,N_3735);
nand U5263 (N_5263,N_3284,N_4103);
nor U5264 (N_5264,N_3491,N_4199);
and U5265 (N_5265,N_3236,N_4011);
nor U5266 (N_5266,N_3031,N_3633);
nor U5267 (N_5267,N_4202,N_3689);
xnor U5268 (N_5268,N_4216,N_3813);
or U5269 (N_5269,N_4493,N_4210);
or U5270 (N_5270,N_3183,N_3671);
nor U5271 (N_5271,N_3217,N_3735);
xnor U5272 (N_5272,N_3024,N_4242);
and U5273 (N_5273,N_3180,N_4484);
and U5274 (N_5274,N_3571,N_3216);
xor U5275 (N_5275,N_4469,N_3720);
xnor U5276 (N_5276,N_3232,N_4233);
xnor U5277 (N_5277,N_3662,N_4094);
and U5278 (N_5278,N_3682,N_3052);
nand U5279 (N_5279,N_3925,N_3868);
nor U5280 (N_5280,N_3423,N_4128);
nand U5281 (N_5281,N_4462,N_3781);
nand U5282 (N_5282,N_3486,N_4223);
and U5283 (N_5283,N_4151,N_3652);
nor U5284 (N_5284,N_3552,N_3879);
xnor U5285 (N_5285,N_4364,N_3112);
and U5286 (N_5286,N_3754,N_3451);
and U5287 (N_5287,N_4235,N_3201);
nand U5288 (N_5288,N_3955,N_3806);
xor U5289 (N_5289,N_3813,N_3181);
nand U5290 (N_5290,N_4483,N_3697);
xor U5291 (N_5291,N_4140,N_3767);
or U5292 (N_5292,N_3745,N_3514);
or U5293 (N_5293,N_3313,N_3497);
or U5294 (N_5294,N_3448,N_4157);
nand U5295 (N_5295,N_4230,N_3447);
or U5296 (N_5296,N_4485,N_3754);
and U5297 (N_5297,N_4251,N_3180);
nor U5298 (N_5298,N_3839,N_3489);
nand U5299 (N_5299,N_3081,N_3107);
and U5300 (N_5300,N_3970,N_3755);
nor U5301 (N_5301,N_4219,N_4098);
xnor U5302 (N_5302,N_3956,N_4164);
and U5303 (N_5303,N_3085,N_3075);
nor U5304 (N_5304,N_3438,N_3756);
and U5305 (N_5305,N_3927,N_4355);
xnor U5306 (N_5306,N_4057,N_3225);
nand U5307 (N_5307,N_3804,N_4179);
nand U5308 (N_5308,N_3097,N_3609);
xnor U5309 (N_5309,N_3400,N_3079);
or U5310 (N_5310,N_3989,N_3717);
nand U5311 (N_5311,N_4216,N_4172);
xor U5312 (N_5312,N_4124,N_3440);
xor U5313 (N_5313,N_3652,N_4216);
or U5314 (N_5314,N_4351,N_3858);
and U5315 (N_5315,N_4068,N_3377);
or U5316 (N_5316,N_3885,N_3399);
nand U5317 (N_5317,N_3324,N_3958);
xnor U5318 (N_5318,N_4012,N_3598);
nor U5319 (N_5319,N_4333,N_3346);
and U5320 (N_5320,N_3301,N_3882);
xor U5321 (N_5321,N_3918,N_3842);
nand U5322 (N_5322,N_3936,N_3521);
nand U5323 (N_5323,N_3046,N_3970);
nand U5324 (N_5324,N_4117,N_4258);
nand U5325 (N_5325,N_3160,N_3177);
or U5326 (N_5326,N_4245,N_3134);
nand U5327 (N_5327,N_3319,N_3996);
nand U5328 (N_5328,N_3497,N_3784);
nor U5329 (N_5329,N_3109,N_3741);
or U5330 (N_5330,N_3062,N_3346);
or U5331 (N_5331,N_4447,N_4177);
nand U5332 (N_5332,N_4479,N_3118);
and U5333 (N_5333,N_3808,N_3020);
xnor U5334 (N_5334,N_4116,N_4252);
xnor U5335 (N_5335,N_3698,N_3393);
or U5336 (N_5336,N_3806,N_4218);
nand U5337 (N_5337,N_3545,N_3514);
or U5338 (N_5338,N_3263,N_3861);
and U5339 (N_5339,N_4318,N_4227);
or U5340 (N_5340,N_3603,N_3399);
xnor U5341 (N_5341,N_3961,N_3782);
nor U5342 (N_5342,N_3714,N_3107);
or U5343 (N_5343,N_3910,N_3862);
nand U5344 (N_5344,N_3764,N_4259);
and U5345 (N_5345,N_3689,N_3997);
nand U5346 (N_5346,N_3092,N_4362);
or U5347 (N_5347,N_4475,N_4085);
nand U5348 (N_5348,N_3173,N_3771);
xor U5349 (N_5349,N_4461,N_3606);
nor U5350 (N_5350,N_3343,N_3427);
nand U5351 (N_5351,N_3185,N_3159);
nor U5352 (N_5352,N_4295,N_3521);
xnor U5353 (N_5353,N_3651,N_4377);
nand U5354 (N_5354,N_3998,N_4124);
nor U5355 (N_5355,N_3889,N_3136);
nor U5356 (N_5356,N_3200,N_4109);
nand U5357 (N_5357,N_4421,N_3790);
nor U5358 (N_5358,N_3049,N_3874);
or U5359 (N_5359,N_3346,N_4274);
xor U5360 (N_5360,N_4167,N_3734);
nand U5361 (N_5361,N_3540,N_3217);
nand U5362 (N_5362,N_4181,N_3929);
or U5363 (N_5363,N_4396,N_3198);
nor U5364 (N_5364,N_3244,N_3497);
nand U5365 (N_5365,N_3869,N_3503);
or U5366 (N_5366,N_3711,N_4388);
or U5367 (N_5367,N_3901,N_3291);
nor U5368 (N_5368,N_3379,N_3659);
or U5369 (N_5369,N_3581,N_3362);
nor U5370 (N_5370,N_3791,N_4134);
and U5371 (N_5371,N_3126,N_3719);
nor U5372 (N_5372,N_3503,N_4081);
and U5373 (N_5373,N_4397,N_3937);
nand U5374 (N_5374,N_3033,N_4360);
xnor U5375 (N_5375,N_3631,N_3351);
xor U5376 (N_5376,N_4168,N_3687);
and U5377 (N_5377,N_4130,N_3839);
xor U5378 (N_5378,N_4403,N_3240);
or U5379 (N_5379,N_3249,N_3297);
or U5380 (N_5380,N_4100,N_3888);
and U5381 (N_5381,N_4476,N_4317);
nor U5382 (N_5382,N_4208,N_3514);
nor U5383 (N_5383,N_4148,N_3704);
nand U5384 (N_5384,N_3006,N_3193);
and U5385 (N_5385,N_4440,N_3630);
xnor U5386 (N_5386,N_3051,N_3440);
nor U5387 (N_5387,N_3708,N_3895);
nor U5388 (N_5388,N_3836,N_3993);
and U5389 (N_5389,N_3436,N_4270);
or U5390 (N_5390,N_3828,N_4266);
xnor U5391 (N_5391,N_3334,N_4271);
xnor U5392 (N_5392,N_4484,N_3800);
nor U5393 (N_5393,N_4188,N_3003);
and U5394 (N_5394,N_4455,N_3113);
or U5395 (N_5395,N_3669,N_3274);
or U5396 (N_5396,N_3925,N_3964);
or U5397 (N_5397,N_3669,N_4402);
or U5398 (N_5398,N_4196,N_3337);
nor U5399 (N_5399,N_3768,N_4231);
or U5400 (N_5400,N_3608,N_3439);
nand U5401 (N_5401,N_3192,N_3427);
xor U5402 (N_5402,N_4398,N_3261);
and U5403 (N_5403,N_3126,N_4293);
nor U5404 (N_5404,N_3611,N_3623);
and U5405 (N_5405,N_3632,N_3253);
and U5406 (N_5406,N_4158,N_3744);
and U5407 (N_5407,N_4204,N_3056);
nor U5408 (N_5408,N_3738,N_3400);
nor U5409 (N_5409,N_3811,N_3714);
or U5410 (N_5410,N_3093,N_4065);
nor U5411 (N_5411,N_4084,N_4183);
xor U5412 (N_5412,N_3001,N_3810);
xor U5413 (N_5413,N_3908,N_4182);
nor U5414 (N_5414,N_3860,N_3552);
xnor U5415 (N_5415,N_3710,N_3670);
and U5416 (N_5416,N_4324,N_3827);
and U5417 (N_5417,N_3942,N_4320);
and U5418 (N_5418,N_3954,N_4412);
xor U5419 (N_5419,N_3279,N_3163);
nand U5420 (N_5420,N_4065,N_4411);
xnor U5421 (N_5421,N_4232,N_4486);
and U5422 (N_5422,N_3903,N_3296);
nand U5423 (N_5423,N_3343,N_3256);
nand U5424 (N_5424,N_4209,N_3619);
and U5425 (N_5425,N_3509,N_3064);
and U5426 (N_5426,N_3913,N_3133);
nor U5427 (N_5427,N_4084,N_3671);
nand U5428 (N_5428,N_4081,N_4117);
xor U5429 (N_5429,N_3489,N_3239);
nor U5430 (N_5430,N_4148,N_3141);
nor U5431 (N_5431,N_3741,N_3343);
xnor U5432 (N_5432,N_3799,N_4214);
nand U5433 (N_5433,N_4232,N_3534);
nor U5434 (N_5434,N_3535,N_3507);
xor U5435 (N_5435,N_4137,N_3051);
and U5436 (N_5436,N_4179,N_3641);
or U5437 (N_5437,N_3718,N_4128);
or U5438 (N_5438,N_3446,N_3810);
xnor U5439 (N_5439,N_3215,N_4453);
xnor U5440 (N_5440,N_3254,N_3273);
and U5441 (N_5441,N_4387,N_3856);
nor U5442 (N_5442,N_3265,N_3622);
and U5443 (N_5443,N_3323,N_3867);
or U5444 (N_5444,N_3232,N_3833);
or U5445 (N_5445,N_3055,N_3368);
or U5446 (N_5446,N_4166,N_4338);
xnor U5447 (N_5447,N_4439,N_4375);
and U5448 (N_5448,N_3640,N_3047);
xnor U5449 (N_5449,N_3669,N_3700);
nand U5450 (N_5450,N_4058,N_4228);
and U5451 (N_5451,N_3314,N_3905);
or U5452 (N_5452,N_3010,N_3215);
and U5453 (N_5453,N_4023,N_4315);
nand U5454 (N_5454,N_4265,N_3500);
or U5455 (N_5455,N_4189,N_3353);
or U5456 (N_5456,N_4284,N_4294);
or U5457 (N_5457,N_4284,N_3228);
xor U5458 (N_5458,N_3473,N_3725);
or U5459 (N_5459,N_3281,N_4359);
nor U5460 (N_5460,N_3355,N_3600);
or U5461 (N_5461,N_3673,N_4259);
xnor U5462 (N_5462,N_3363,N_3441);
xor U5463 (N_5463,N_3293,N_3114);
and U5464 (N_5464,N_3617,N_3689);
and U5465 (N_5465,N_4427,N_4128);
xnor U5466 (N_5466,N_3111,N_4088);
or U5467 (N_5467,N_3498,N_4017);
nand U5468 (N_5468,N_4015,N_3691);
nand U5469 (N_5469,N_4253,N_3538);
nor U5470 (N_5470,N_3859,N_4312);
or U5471 (N_5471,N_3080,N_3682);
nand U5472 (N_5472,N_3474,N_4064);
nand U5473 (N_5473,N_3447,N_3185);
nor U5474 (N_5474,N_3572,N_4235);
or U5475 (N_5475,N_3858,N_4229);
xor U5476 (N_5476,N_4425,N_3350);
xnor U5477 (N_5477,N_3823,N_4225);
nand U5478 (N_5478,N_3596,N_3515);
and U5479 (N_5479,N_3473,N_4348);
nand U5480 (N_5480,N_3621,N_4058);
nand U5481 (N_5481,N_3305,N_3677);
nand U5482 (N_5482,N_3938,N_3728);
nor U5483 (N_5483,N_3792,N_3926);
or U5484 (N_5484,N_3857,N_3793);
nor U5485 (N_5485,N_4165,N_4008);
or U5486 (N_5486,N_3982,N_3046);
and U5487 (N_5487,N_4387,N_3269);
xnor U5488 (N_5488,N_4338,N_4134);
nor U5489 (N_5489,N_3054,N_4303);
or U5490 (N_5490,N_4296,N_3408);
nor U5491 (N_5491,N_4480,N_3738);
and U5492 (N_5492,N_3319,N_3231);
and U5493 (N_5493,N_3980,N_3434);
and U5494 (N_5494,N_3319,N_3649);
nand U5495 (N_5495,N_4172,N_3640);
nor U5496 (N_5496,N_3761,N_3157);
nor U5497 (N_5497,N_4459,N_3609);
nand U5498 (N_5498,N_3732,N_4209);
and U5499 (N_5499,N_4002,N_3518);
nand U5500 (N_5500,N_3269,N_3316);
and U5501 (N_5501,N_4378,N_3205);
nand U5502 (N_5502,N_4328,N_4456);
or U5503 (N_5503,N_4410,N_4142);
xor U5504 (N_5504,N_3932,N_4158);
and U5505 (N_5505,N_3899,N_4349);
xor U5506 (N_5506,N_4203,N_3832);
nor U5507 (N_5507,N_3797,N_3496);
xor U5508 (N_5508,N_3051,N_3204);
xnor U5509 (N_5509,N_4324,N_3035);
or U5510 (N_5510,N_4475,N_3912);
or U5511 (N_5511,N_3643,N_3368);
or U5512 (N_5512,N_3603,N_3730);
nand U5513 (N_5513,N_4332,N_3750);
xor U5514 (N_5514,N_4096,N_3281);
xor U5515 (N_5515,N_3633,N_4453);
and U5516 (N_5516,N_4314,N_4078);
nand U5517 (N_5517,N_3605,N_3565);
and U5518 (N_5518,N_3578,N_4221);
nand U5519 (N_5519,N_3762,N_4480);
xnor U5520 (N_5520,N_4489,N_4215);
and U5521 (N_5521,N_4451,N_3707);
nor U5522 (N_5522,N_3904,N_4385);
nand U5523 (N_5523,N_3154,N_3578);
nor U5524 (N_5524,N_3845,N_3692);
nand U5525 (N_5525,N_4182,N_3082);
nor U5526 (N_5526,N_3574,N_3991);
xor U5527 (N_5527,N_4229,N_3188);
nand U5528 (N_5528,N_4051,N_3514);
nor U5529 (N_5529,N_3113,N_3390);
nor U5530 (N_5530,N_4473,N_4352);
xnor U5531 (N_5531,N_4487,N_4177);
and U5532 (N_5532,N_3719,N_4282);
nor U5533 (N_5533,N_3842,N_3088);
xnor U5534 (N_5534,N_3135,N_3418);
xor U5535 (N_5535,N_4198,N_3454);
nand U5536 (N_5536,N_3256,N_3861);
and U5537 (N_5537,N_4003,N_4114);
nor U5538 (N_5538,N_4371,N_3634);
nand U5539 (N_5539,N_3770,N_3411);
nand U5540 (N_5540,N_4101,N_4450);
xor U5541 (N_5541,N_4066,N_3101);
nand U5542 (N_5542,N_3979,N_3556);
nor U5543 (N_5543,N_4007,N_4156);
or U5544 (N_5544,N_3577,N_3155);
xor U5545 (N_5545,N_4057,N_3724);
nand U5546 (N_5546,N_4334,N_3682);
and U5547 (N_5547,N_3342,N_3002);
nor U5548 (N_5548,N_4480,N_4384);
xor U5549 (N_5549,N_4231,N_3978);
xor U5550 (N_5550,N_3043,N_3523);
nand U5551 (N_5551,N_4061,N_3940);
or U5552 (N_5552,N_4120,N_4085);
and U5553 (N_5553,N_3254,N_3034);
nand U5554 (N_5554,N_4425,N_4051);
xor U5555 (N_5555,N_4063,N_4201);
and U5556 (N_5556,N_4000,N_3730);
xor U5557 (N_5557,N_4020,N_4237);
nand U5558 (N_5558,N_4213,N_3524);
or U5559 (N_5559,N_4026,N_4364);
nand U5560 (N_5560,N_3177,N_4184);
xnor U5561 (N_5561,N_3222,N_3421);
nor U5562 (N_5562,N_4223,N_3589);
nor U5563 (N_5563,N_3498,N_4377);
and U5564 (N_5564,N_4100,N_4240);
or U5565 (N_5565,N_3108,N_3148);
and U5566 (N_5566,N_4164,N_3606);
xor U5567 (N_5567,N_3816,N_4366);
and U5568 (N_5568,N_4142,N_4121);
and U5569 (N_5569,N_3481,N_3642);
or U5570 (N_5570,N_3653,N_3915);
and U5571 (N_5571,N_3165,N_3586);
xnor U5572 (N_5572,N_3410,N_3763);
and U5573 (N_5573,N_4230,N_3346);
and U5574 (N_5574,N_4269,N_4391);
nor U5575 (N_5575,N_4212,N_3541);
nand U5576 (N_5576,N_4243,N_4072);
nand U5577 (N_5577,N_4019,N_3187);
or U5578 (N_5578,N_4319,N_3583);
and U5579 (N_5579,N_3853,N_3226);
xor U5580 (N_5580,N_4138,N_3866);
or U5581 (N_5581,N_3333,N_3133);
or U5582 (N_5582,N_3865,N_4184);
and U5583 (N_5583,N_4018,N_3807);
and U5584 (N_5584,N_3024,N_3400);
or U5585 (N_5585,N_3140,N_4102);
xor U5586 (N_5586,N_4312,N_4411);
or U5587 (N_5587,N_4364,N_4129);
and U5588 (N_5588,N_4406,N_4110);
xnor U5589 (N_5589,N_4210,N_3001);
nand U5590 (N_5590,N_3552,N_4177);
nor U5591 (N_5591,N_4006,N_4402);
and U5592 (N_5592,N_4146,N_4092);
xnor U5593 (N_5593,N_3423,N_3380);
nand U5594 (N_5594,N_4428,N_3207);
and U5595 (N_5595,N_4449,N_3439);
or U5596 (N_5596,N_3446,N_4211);
and U5597 (N_5597,N_3345,N_3770);
nor U5598 (N_5598,N_3434,N_3859);
and U5599 (N_5599,N_4141,N_3042);
nor U5600 (N_5600,N_3912,N_3109);
and U5601 (N_5601,N_3173,N_3562);
and U5602 (N_5602,N_4266,N_4024);
nor U5603 (N_5603,N_3943,N_3924);
nand U5604 (N_5604,N_4001,N_3339);
nor U5605 (N_5605,N_4243,N_3834);
nand U5606 (N_5606,N_3757,N_3599);
xor U5607 (N_5607,N_3887,N_3169);
nor U5608 (N_5608,N_4074,N_3637);
and U5609 (N_5609,N_4423,N_3237);
nand U5610 (N_5610,N_4395,N_3296);
nand U5611 (N_5611,N_3123,N_3547);
xor U5612 (N_5612,N_3615,N_3948);
nor U5613 (N_5613,N_4467,N_3256);
and U5614 (N_5614,N_4078,N_4387);
xor U5615 (N_5615,N_4420,N_3861);
or U5616 (N_5616,N_4342,N_3500);
and U5617 (N_5617,N_4097,N_3269);
xnor U5618 (N_5618,N_4121,N_3416);
xor U5619 (N_5619,N_3197,N_3325);
xor U5620 (N_5620,N_3753,N_4413);
xor U5621 (N_5621,N_3533,N_3313);
nor U5622 (N_5622,N_3392,N_3896);
and U5623 (N_5623,N_3431,N_3653);
or U5624 (N_5624,N_3778,N_4127);
or U5625 (N_5625,N_3612,N_3125);
xnor U5626 (N_5626,N_4147,N_4408);
or U5627 (N_5627,N_4115,N_3091);
nand U5628 (N_5628,N_3934,N_3770);
nor U5629 (N_5629,N_3830,N_3275);
and U5630 (N_5630,N_3971,N_4478);
or U5631 (N_5631,N_4194,N_3498);
nand U5632 (N_5632,N_3612,N_4446);
nand U5633 (N_5633,N_3618,N_4445);
xor U5634 (N_5634,N_3426,N_4474);
xor U5635 (N_5635,N_4249,N_4110);
nand U5636 (N_5636,N_4205,N_3718);
xor U5637 (N_5637,N_3212,N_4066);
or U5638 (N_5638,N_3350,N_3762);
nor U5639 (N_5639,N_4333,N_3545);
and U5640 (N_5640,N_4413,N_3989);
and U5641 (N_5641,N_3795,N_3756);
nand U5642 (N_5642,N_3106,N_3277);
or U5643 (N_5643,N_3621,N_3454);
nor U5644 (N_5644,N_3099,N_3801);
and U5645 (N_5645,N_3944,N_4082);
nand U5646 (N_5646,N_3075,N_3291);
and U5647 (N_5647,N_3462,N_4035);
and U5648 (N_5648,N_4323,N_4460);
or U5649 (N_5649,N_3778,N_3928);
or U5650 (N_5650,N_4426,N_4085);
nand U5651 (N_5651,N_4013,N_4304);
or U5652 (N_5652,N_4025,N_3170);
and U5653 (N_5653,N_3295,N_3649);
or U5654 (N_5654,N_3503,N_3417);
nand U5655 (N_5655,N_3769,N_4457);
or U5656 (N_5656,N_4472,N_3208);
nor U5657 (N_5657,N_3225,N_4036);
or U5658 (N_5658,N_3568,N_3081);
or U5659 (N_5659,N_4316,N_3405);
nand U5660 (N_5660,N_4490,N_4002);
nand U5661 (N_5661,N_3530,N_4288);
and U5662 (N_5662,N_4050,N_4479);
nand U5663 (N_5663,N_3986,N_3890);
nor U5664 (N_5664,N_4306,N_3695);
and U5665 (N_5665,N_3063,N_3990);
xnor U5666 (N_5666,N_4279,N_4172);
nor U5667 (N_5667,N_4461,N_4430);
xor U5668 (N_5668,N_3714,N_3927);
nor U5669 (N_5669,N_3895,N_4401);
nand U5670 (N_5670,N_4358,N_4386);
and U5671 (N_5671,N_3840,N_3915);
nor U5672 (N_5672,N_4178,N_3113);
nand U5673 (N_5673,N_3161,N_3793);
nand U5674 (N_5674,N_4411,N_3176);
nor U5675 (N_5675,N_3715,N_3879);
nand U5676 (N_5676,N_3617,N_4109);
nand U5677 (N_5677,N_3898,N_3758);
nand U5678 (N_5678,N_3016,N_4456);
and U5679 (N_5679,N_4457,N_4270);
nand U5680 (N_5680,N_4029,N_4470);
or U5681 (N_5681,N_3700,N_3930);
and U5682 (N_5682,N_3266,N_3558);
and U5683 (N_5683,N_3222,N_3080);
or U5684 (N_5684,N_3983,N_3637);
xor U5685 (N_5685,N_3823,N_3052);
nand U5686 (N_5686,N_4475,N_4352);
nand U5687 (N_5687,N_3136,N_3899);
or U5688 (N_5688,N_4282,N_3537);
and U5689 (N_5689,N_3264,N_4347);
xor U5690 (N_5690,N_3481,N_3878);
xnor U5691 (N_5691,N_4201,N_4485);
and U5692 (N_5692,N_3598,N_3710);
or U5693 (N_5693,N_3193,N_3663);
nand U5694 (N_5694,N_3140,N_4033);
xor U5695 (N_5695,N_4438,N_4488);
and U5696 (N_5696,N_3612,N_3205);
nand U5697 (N_5697,N_4001,N_4201);
nand U5698 (N_5698,N_3775,N_4367);
nor U5699 (N_5699,N_3846,N_3781);
xnor U5700 (N_5700,N_3522,N_3462);
and U5701 (N_5701,N_3758,N_3818);
and U5702 (N_5702,N_3591,N_4239);
xnor U5703 (N_5703,N_3621,N_4344);
or U5704 (N_5704,N_4463,N_4119);
nand U5705 (N_5705,N_3939,N_4190);
or U5706 (N_5706,N_4165,N_3205);
xor U5707 (N_5707,N_3921,N_4252);
xnor U5708 (N_5708,N_4137,N_3989);
nand U5709 (N_5709,N_3430,N_3326);
or U5710 (N_5710,N_4327,N_3061);
nor U5711 (N_5711,N_3321,N_4449);
nand U5712 (N_5712,N_4172,N_4255);
and U5713 (N_5713,N_3828,N_3619);
and U5714 (N_5714,N_3484,N_4458);
and U5715 (N_5715,N_4375,N_3763);
nor U5716 (N_5716,N_4050,N_3357);
or U5717 (N_5717,N_4138,N_4006);
xor U5718 (N_5718,N_4197,N_4399);
nand U5719 (N_5719,N_4000,N_3205);
or U5720 (N_5720,N_4273,N_3595);
or U5721 (N_5721,N_3325,N_3952);
and U5722 (N_5722,N_3421,N_3961);
and U5723 (N_5723,N_3782,N_4044);
nand U5724 (N_5724,N_3861,N_3175);
and U5725 (N_5725,N_3704,N_4258);
nor U5726 (N_5726,N_3392,N_4131);
xor U5727 (N_5727,N_4091,N_3402);
nor U5728 (N_5728,N_3993,N_3727);
xnor U5729 (N_5729,N_3968,N_4468);
xor U5730 (N_5730,N_3728,N_4218);
xnor U5731 (N_5731,N_3301,N_3849);
nor U5732 (N_5732,N_4160,N_4322);
nand U5733 (N_5733,N_3363,N_3806);
xor U5734 (N_5734,N_3479,N_3651);
xor U5735 (N_5735,N_3149,N_3573);
nand U5736 (N_5736,N_4080,N_4305);
xor U5737 (N_5737,N_4188,N_4127);
and U5738 (N_5738,N_4407,N_3988);
nand U5739 (N_5739,N_3389,N_4466);
nand U5740 (N_5740,N_3607,N_4157);
nand U5741 (N_5741,N_3704,N_3148);
and U5742 (N_5742,N_3573,N_3584);
nand U5743 (N_5743,N_3972,N_3009);
nand U5744 (N_5744,N_3897,N_4443);
or U5745 (N_5745,N_3160,N_3109);
nand U5746 (N_5746,N_4259,N_3559);
nor U5747 (N_5747,N_3739,N_3309);
or U5748 (N_5748,N_3343,N_3250);
nand U5749 (N_5749,N_3517,N_3538);
xor U5750 (N_5750,N_3226,N_3664);
or U5751 (N_5751,N_4434,N_3322);
or U5752 (N_5752,N_4459,N_3511);
nor U5753 (N_5753,N_3895,N_4059);
or U5754 (N_5754,N_3813,N_3070);
xor U5755 (N_5755,N_4283,N_4462);
and U5756 (N_5756,N_3098,N_4431);
nand U5757 (N_5757,N_3289,N_3796);
nand U5758 (N_5758,N_3540,N_4457);
and U5759 (N_5759,N_3714,N_4439);
nor U5760 (N_5760,N_3117,N_3180);
nor U5761 (N_5761,N_4368,N_3651);
nand U5762 (N_5762,N_3810,N_3872);
xnor U5763 (N_5763,N_3225,N_3004);
nand U5764 (N_5764,N_3498,N_4185);
xor U5765 (N_5765,N_3420,N_3104);
nand U5766 (N_5766,N_4424,N_3786);
nand U5767 (N_5767,N_3049,N_3608);
nor U5768 (N_5768,N_3511,N_4038);
xor U5769 (N_5769,N_3745,N_3183);
xnor U5770 (N_5770,N_4249,N_4159);
and U5771 (N_5771,N_3663,N_3830);
or U5772 (N_5772,N_3632,N_4377);
or U5773 (N_5773,N_4446,N_3231);
or U5774 (N_5774,N_4231,N_3433);
nand U5775 (N_5775,N_3888,N_3211);
or U5776 (N_5776,N_3410,N_3607);
or U5777 (N_5777,N_4467,N_4043);
xor U5778 (N_5778,N_3462,N_3145);
or U5779 (N_5779,N_3348,N_4298);
or U5780 (N_5780,N_3858,N_3237);
or U5781 (N_5781,N_3971,N_3653);
nor U5782 (N_5782,N_3942,N_3312);
nor U5783 (N_5783,N_4033,N_3744);
nor U5784 (N_5784,N_3459,N_3305);
or U5785 (N_5785,N_3250,N_4135);
and U5786 (N_5786,N_3945,N_4259);
or U5787 (N_5787,N_3156,N_3878);
and U5788 (N_5788,N_3248,N_3509);
nor U5789 (N_5789,N_3414,N_3184);
nor U5790 (N_5790,N_4006,N_3214);
nor U5791 (N_5791,N_3981,N_3339);
nand U5792 (N_5792,N_3759,N_4066);
and U5793 (N_5793,N_3485,N_3371);
xor U5794 (N_5794,N_3140,N_3266);
nand U5795 (N_5795,N_3410,N_3529);
nand U5796 (N_5796,N_4166,N_3190);
or U5797 (N_5797,N_4326,N_3004);
or U5798 (N_5798,N_4288,N_4083);
and U5799 (N_5799,N_3958,N_3260);
nor U5800 (N_5800,N_3877,N_3340);
or U5801 (N_5801,N_3804,N_4039);
or U5802 (N_5802,N_3999,N_4009);
nand U5803 (N_5803,N_3588,N_4371);
xnor U5804 (N_5804,N_3600,N_4375);
xnor U5805 (N_5805,N_3529,N_3173);
and U5806 (N_5806,N_4301,N_3784);
or U5807 (N_5807,N_4333,N_3668);
nand U5808 (N_5808,N_4098,N_3845);
and U5809 (N_5809,N_3673,N_3500);
or U5810 (N_5810,N_4309,N_3413);
and U5811 (N_5811,N_3585,N_3129);
nand U5812 (N_5812,N_3384,N_4062);
or U5813 (N_5813,N_4114,N_3982);
xor U5814 (N_5814,N_3437,N_3587);
and U5815 (N_5815,N_4228,N_3273);
nor U5816 (N_5816,N_4140,N_3224);
and U5817 (N_5817,N_3037,N_4476);
and U5818 (N_5818,N_3907,N_4308);
and U5819 (N_5819,N_4318,N_3119);
nor U5820 (N_5820,N_3301,N_3675);
nor U5821 (N_5821,N_3361,N_3354);
or U5822 (N_5822,N_3938,N_3284);
and U5823 (N_5823,N_3400,N_3499);
and U5824 (N_5824,N_4220,N_4449);
nand U5825 (N_5825,N_3895,N_4254);
or U5826 (N_5826,N_4173,N_3561);
nor U5827 (N_5827,N_3418,N_3861);
or U5828 (N_5828,N_3090,N_3654);
nand U5829 (N_5829,N_3989,N_3628);
xor U5830 (N_5830,N_4386,N_3256);
nand U5831 (N_5831,N_4279,N_3626);
nand U5832 (N_5832,N_3867,N_3319);
nand U5833 (N_5833,N_3076,N_3815);
nand U5834 (N_5834,N_3715,N_3765);
and U5835 (N_5835,N_3754,N_4219);
and U5836 (N_5836,N_3769,N_3165);
nor U5837 (N_5837,N_4377,N_3818);
and U5838 (N_5838,N_3141,N_3278);
xnor U5839 (N_5839,N_3611,N_3999);
or U5840 (N_5840,N_3131,N_4302);
nor U5841 (N_5841,N_3539,N_3767);
nor U5842 (N_5842,N_3964,N_3695);
nand U5843 (N_5843,N_3303,N_3718);
or U5844 (N_5844,N_4341,N_4407);
nand U5845 (N_5845,N_3926,N_3864);
xor U5846 (N_5846,N_3456,N_4345);
or U5847 (N_5847,N_4215,N_3262);
nand U5848 (N_5848,N_3027,N_3389);
nand U5849 (N_5849,N_3536,N_3092);
or U5850 (N_5850,N_3477,N_3481);
nor U5851 (N_5851,N_3721,N_3521);
xnor U5852 (N_5852,N_3382,N_3760);
or U5853 (N_5853,N_4312,N_4027);
nor U5854 (N_5854,N_3092,N_4437);
xor U5855 (N_5855,N_4070,N_4224);
and U5856 (N_5856,N_4419,N_4290);
nor U5857 (N_5857,N_3198,N_3071);
and U5858 (N_5858,N_3415,N_3562);
or U5859 (N_5859,N_4268,N_3514);
and U5860 (N_5860,N_3900,N_3683);
and U5861 (N_5861,N_3049,N_4260);
nand U5862 (N_5862,N_4052,N_3631);
xnor U5863 (N_5863,N_4439,N_3485);
xor U5864 (N_5864,N_3616,N_4458);
and U5865 (N_5865,N_4177,N_3999);
nor U5866 (N_5866,N_3628,N_3019);
nand U5867 (N_5867,N_3801,N_3224);
or U5868 (N_5868,N_3320,N_4088);
xnor U5869 (N_5869,N_3499,N_4186);
and U5870 (N_5870,N_4244,N_3443);
xor U5871 (N_5871,N_3945,N_4359);
nand U5872 (N_5872,N_3596,N_3723);
nor U5873 (N_5873,N_4020,N_3121);
or U5874 (N_5874,N_4301,N_3542);
and U5875 (N_5875,N_4460,N_4300);
nor U5876 (N_5876,N_3011,N_4201);
or U5877 (N_5877,N_3714,N_3605);
nand U5878 (N_5878,N_3451,N_3829);
or U5879 (N_5879,N_4065,N_3671);
or U5880 (N_5880,N_4307,N_3839);
nand U5881 (N_5881,N_3957,N_4241);
and U5882 (N_5882,N_3270,N_3279);
xor U5883 (N_5883,N_4065,N_3342);
nand U5884 (N_5884,N_3236,N_3710);
and U5885 (N_5885,N_3040,N_4250);
and U5886 (N_5886,N_3582,N_3153);
and U5887 (N_5887,N_3123,N_3936);
nand U5888 (N_5888,N_3533,N_3241);
or U5889 (N_5889,N_4010,N_3580);
xnor U5890 (N_5890,N_3629,N_4154);
nand U5891 (N_5891,N_3484,N_3217);
or U5892 (N_5892,N_3306,N_4080);
xnor U5893 (N_5893,N_3736,N_3536);
or U5894 (N_5894,N_3298,N_3135);
and U5895 (N_5895,N_4415,N_4233);
and U5896 (N_5896,N_3630,N_3563);
or U5897 (N_5897,N_3154,N_3493);
and U5898 (N_5898,N_3035,N_4029);
xor U5899 (N_5899,N_3942,N_3529);
nor U5900 (N_5900,N_4106,N_3471);
nor U5901 (N_5901,N_3360,N_4207);
nor U5902 (N_5902,N_4309,N_3757);
nor U5903 (N_5903,N_3812,N_3135);
nand U5904 (N_5904,N_4295,N_3127);
or U5905 (N_5905,N_4281,N_3131);
or U5906 (N_5906,N_3388,N_3531);
xnor U5907 (N_5907,N_3178,N_4397);
xnor U5908 (N_5908,N_3016,N_3185);
or U5909 (N_5909,N_3822,N_3364);
or U5910 (N_5910,N_4025,N_4406);
or U5911 (N_5911,N_3118,N_4381);
nor U5912 (N_5912,N_4059,N_3781);
or U5913 (N_5913,N_3806,N_3552);
nand U5914 (N_5914,N_3211,N_3889);
and U5915 (N_5915,N_3617,N_3451);
nand U5916 (N_5916,N_3531,N_3448);
and U5917 (N_5917,N_3955,N_3253);
nand U5918 (N_5918,N_4312,N_3171);
and U5919 (N_5919,N_4235,N_4156);
xor U5920 (N_5920,N_3566,N_3040);
xnor U5921 (N_5921,N_3366,N_3287);
xnor U5922 (N_5922,N_3708,N_3021);
xor U5923 (N_5923,N_4290,N_3239);
and U5924 (N_5924,N_4342,N_3613);
and U5925 (N_5925,N_3298,N_3525);
nand U5926 (N_5926,N_3721,N_3093);
nand U5927 (N_5927,N_3580,N_4047);
nor U5928 (N_5928,N_3606,N_4368);
or U5929 (N_5929,N_3352,N_3645);
xnor U5930 (N_5930,N_3533,N_3849);
or U5931 (N_5931,N_3765,N_3210);
nand U5932 (N_5932,N_4071,N_3842);
nand U5933 (N_5933,N_3634,N_3861);
xnor U5934 (N_5934,N_3476,N_3126);
nor U5935 (N_5935,N_3314,N_3345);
xnor U5936 (N_5936,N_3627,N_3908);
xor U5937 (N_5937,N_4023,N_3550);
xnor U5938 (N_5938,N_4171,N_4229);
nor U5939 (N_5939,N_3522,N_4435);
or U5940 (N_5940,N_3952,N_4224);
xnor U5941 (N_5941,N_4102,N_3192);
or U5942 (N_5942,N_3893,N_3972);
nand U5943 (N_5943,N_3047,N_3514);
and U5944 (N_5944,N_4476,N_3165);
or U5945 (N_5945,N_3459,N_3509);
and U5946 (N_5946,N_3190,N_3396);
nor U5947 (N_5947,N_3286,N_4425);
and U5948 (N_5948,N_3780,N_4053);
nor U5949 (N_5949,N_3272,N_3782);
and U5950 (N_5950,N_3880,N_3894);
nor U5951 (N_5951,N_3206,N_3195);
or U5952 (N_5952,N_3489,N_4461);
and U5953 (N_5953,N_3504,N_4086);
nand U5954 (N_5954,N_4055,N_3836);
nand U5955 (N_5955,N_4402,N_4034);
and U5956 (N_5956,N_4107,N_3615);
nor U5957 (N_5957,N_3503,N_3547);
and U5958 (N_5958,N_3182,N_4006);
nor U5959 (N_5959,N_3300,N_3301);
or U5960 (N_5960,N_3355,N_4419);
xnor U5961 (N_5961,N_3429,N_4107);
nand U5962 (N_5962,N_4260,N_3918);
and U5963 (N_5963,N_3870,N_3261);
nor U5964 (N_5964,N_3311,N_4414);
or U5965 (N_5965,N_3597,N_4072);
or U5966 (N_5966,N_3231,N_4014);
nand U5967 (N_5967,N_4020,N_3600);
or U5968 (N_5968,N_3592,N_3437);
nor U5969 (N_5969,N_3732,N_4283);
nand U5970 (N_5970,N_3666,N_4414);
and U5971 (N_5971,N_3524,N_3516);
nor U5972 (N_5972,N_3567,N_3139);
and U5973 (N_5973,N_3484,N_3819);
nor U5974 (N_5974,N_3575,N_4297);
and U5975 (N_5975,N_3795,N_3648);
nor U5976 (N_5976,N_3491,N_3774);
or U5977 (N_5977,N_3567,N_4302);
nor U5978 (N_5978,N_3966,N_3746);
nand U5979 (N_5979,N_3642,N_3654);
nor U5980 (N_5980,N_4179,N_4408);
nand U5981 (N_5981,N_4019,N_3367);
nor U5982 (N_5982,N_3276,N_3793);
and U5983 (N_5983,N_4327,N_3986);
and U5984 (N_5984,N_3585,N_4214);
xnor U5985 (N_5985,N_3074,N_3524);
and U5986 (N_5986,N_4234,N_3518);
nand U5987 (N_5987,N_3535,N_4467);
nor U5988 (N_5988,N_3438,N_3232);
nor U5989 (N_5989,N_3182,N_3932);
and U5990 (N_5990,N_3524,N_3134);
xnor U5991 (N_5991,N_4160,N_3743);
nor U5992 (N_5992,N_3762,N_4191);
xor U5993 (N_5993,N_3069,N_4133);
or U5994 (N_5994,N_4028,N_3576);
or U5995 (N_5995,N_3230,N_4256);
and U5996 (N_5996,N_4163,N_4427);
nand U5997 (N_5997,N_3536,N_4469);
or U5998 (N_5998,N_4465,N_3285);
or U5999 (N_5999,N_3892,N_3284);
or U6000 (N_6000,N_5407,N_5097);
xnor U6001 (N_6001,N_4970,N_4826);
nand U6002 (N_6002,N_5490,N_5600);
xnor U6003 (N_6003,N_5044,N_5760);
nand U6004 (N_6004,N_5919,N_5526);
and U6005 (N_6005,N_5889,N_4751);
nand U6006 (N_6006,N_4976,N_5505);
nand U6007 (N_6007,N_5682,N_5509);
xnor U6008 (N_6008,N_4821,N_5788);
xnor U6009 (N_6009,N_5506,N_4775);
and U6010 (N_6010,N_5213,N_5110);
xor U6011 (N_6011,N_4778,N_5549);
nand U6012 (N_6012,N_5137,N_5848);
nand U6013 (N_6013,N_4990,N_5601);
nand U6014 (N_6014,N_5071,N_5843);
and U6015 (N_6015,N_4756,N_5963);
and U6016 (N_6016,N_5274,N_5058);
xor U6017 (N_6017,N_5775,N_5145);
xor U6018 (N_6018,N_4637,N_5756);
or U6019 (N_6019,N_5221,N_5098);
or U6020 (N_6020,N_5479,N_5380);
or U6021 (N_6021,N_5295,N_4586);
xnor U6022 (N_6022,N_5829,N_5844);
or U6023 (N_6023,N_5878,N_5012);
xor U6024 (N_6024,N_5348,N_5866);
nor U6025 (N_6025,N_5925,N_5203);
nand U6026 (N_6026,N_5504,N_4791);
xor U6027 (N_6027,N_4937,N_5861);
and U6028 (N_6028,N_4793,N_5054);
or U6029 (N_6029,N_4918,N_5056);
nand U6030 (N_6030,N_5622,N_4707);
nor U6031 (N_6031,N_4571,N_4521);
or U6032 (N_6032,N_5460,N_4881);
xor U6033 (N_6033,N_5793,N_5214);
and U6034 (N_6034,N_5238,N_5027);
and U6035 (N_6035,N_5146,N_5670);
and U6036 (N_6036,N_5800,N_4520);
and U6037 (N_6037,N_5372,N_4538);
xnor U6038 (N_6038,N_5961,N_4753);
and U6039 (N_6039,N_4574,N_5086);
or U6040 (N_6040,N_4942,N_5336);
or U6041 (N_6041,N_5088,N_5651);
nand U6042 (N_6042,N_5650,N_5183);
xor U6043 (N_6043,N_4642,N_4506);
nand U6044 (N_6044,N_5576,N_4687);
or U6045 (N_6045,N_5677,N_4540);
nand U6046 (N_6046,N_4924,N_4670);
or U6047 (N_6047,N_4995,N_4633);
and U6048 (N_6048,N_5035,N_5293);
and U6049 (N_6049,N_5053,N_4974);
nor U6050 (N_6050,N_5799,N_5022);
or U6051 (N_6051,N_5117,N_5939);
nand U6052 (N_6052,N_5227,N_4711);
nor U6053 (N_6053,N_5684,N_4964);
nor U6054 (N_6054,N_4525,N_4700);
xor U6055 (N_6055,N_5329,N_5637);
and U6056 (N_6056,N_5968,N_5915);
and U6057 (N_6057,N_4729,N_5817);
nor U6058 (N_6058,N_5313,N_5176);
nand U6059 (N_6059,N_5438,N_4664);
and U6060 (N_6060,N_5898,N_4721);
and U6061 (N_6061,N_5778,N_5278);
nand U6062 (N_6062,N_5201,N_5825);
nand U6063 (N_6063,N_5165,N_5363);
xor U6064 (N_6064,N_5218,N_5748);
nand U6065 (N_6065,N_4734,N_5624);
xor U6066 (N_6066,N_5900,N_4725);
and U6067 (N_6067,N_5444,N_4871);
or U6068 (N_6068,N_4983,N_4578);
nand U6069 (N_6069,N_5710,N_4740);
nand U6070 (N_6070,N_5141,N_5580);
xor U6071 (N_6071,N_5230,N_5541);
nand U6072 (N_6072,N_5254,N_5833);
nand U6073 (N_6073,N_5072,N_4519);
nor U6074 (N_6074,N_5808,N_4653);
nor U6075 (N_6075,N_5286,N_4545);
and U6076 (N_6076,N_5699,N_5036);
and U6077 (N_6077,N_5926,N_4602);
xor U6078 (N_6078,N_5887,N_5522);
xnor U6079 (N_6079,N_5729,N_5311);
and U6080 (N_6080,N_5773,N_5248);
or U6081 (N_6081,N_5790,N_5066);
nand U6082 (N_6082,N_5344,N_5273);
nor U6083 (N_6083,N_5596,N_4855);
xnor U6084 (N_6084,N_5802,N_4548);
xnor U6085 (N_6085,N_5152,N_5157);
and U6086 (N_6086,N_5255,N_5743);
nand U6087 (N_6087,N_4730,N_4912);
or U6088 (N_6088,N_5378,N_4661);
nand U6089 (N_6089,N_5160,N_5753);
and U6090 (N_6090,N_5211,N_4958);
nor U6091 (N_6091,N_5256,N_5392);
nor U6092 (N_6092,N_4773,N_4659);
xor U6093 (N_6093,N_5482,N_5394);
xnor U6094 (N_6094,N_5084,N_5060);
nand U6095 (N_6095,N_5660,N_5385);
nand U6096 (N_6096,N_4557,N_5477);
nand U6097 (N_6097,N_5289,N_5276);
nor U6098 (N_6098,N_4712,N_4630);
and U6099 (N_6099,N_5193,N_4706);
or U6100 (N_6100,N_5496,N_5706);
xnor U6101 (N_6101,N_5062,N_5987);
nor U6102 (N_6102,N_5630,N_4731);
xor U6103 (N_6103,N_4910,N_5581);
nor U6104 (N_6104,N_5198,N_4819);
xor U6105 (N_6105,N_4652,N_4722);
nand U6106 (N_6106,N_5636,N_5920);
xnor U6107 (N_6107,N_4627,N_5190);
or U6108 (N_6108,N_5408,N_5991);
nor U6109 (N_6109,N_5972,N_5319);
xnor U6110 (N_6110,N_5184,N_5483);
and U6111 (N_6111,N_4530,N_5965);
nor U6112 (N_6112,N_5280,N_4579);
or U6113 (N_6113,N_4542,N_5030);
nor U6114 (N_6114,N_5954,N_5481);
xor U6115 (N_6115,N_5130,N_5820);
nor U6116 (N_6116,N_5649,N_4795);
and U6117 (N_6117,N_5026,N_5958);
and U6118 (N_6118,N_5924,N_5434);
and U6119 (N_6119,N_5390,N_5654);
nand U6120 (N_6120,N_5494,N_5261);
nor U6121 (N_6121,N_5129,N_5700);
or U6122 (N_6122,N_5976,N_5400);
and U6123 (N_6123,N_4555,N_5017);
nor U6124 (N_6124,N_5818,N_5448);
or U6125 (N_6125,N_5167,N_5163);
and U6126 (N_6126,N_4922,N_4864);
nand U6127 (N_6127,N_5688,N_5181);
nand U6128 (N_6128,N_5376,N_5462);
and U6129 (N_6129,N_5065,N_4893);
xor U6130 (N_6130,N_5069,N_5565);
and U6131 (N_6131,N_4556,N_5153);
or U6132 (N_6132,N_5902,N_5795);
nand U6133 (N_6133,N_5139,N_5288);
or U6134 (N_6134,N_4758,N_4547);
or U6135 (N_6135,N_5510,N_4903);
nor U6136 (N_6136,N_5405,N_5171);
or U6137 (N_6137,N_4897,N_4858);
nor U6138 (N_6138,N_5388,N_5421);
xnor U6139 (N_6139,N_5502,N_5708);
or U6140 (N_6140,N_5352,N_5142);
and U6141 (N_6141,N_5767,N_4854);
nor U6142 (N_6142,N_4639,N_4656);
xnor U6143 (N_6143,N_5912,N_5696);
xnor U6144 (N_6144,N_4619,N_4752);
nor U6145 (N_6145,N_5657,N_5331);
nor U6146 (N_6146,N_5094,N_4662);
or U6147 (N_6147,N_4772,N_5493);
nand U6148 (N_6148,N_5173,N_5822);
xnor U6149 (N_6149,N_5233,N_5835);
or U6150 (N_6150,N_4714,N_5740);
nor U6151 (N_6151,N_5321,N_5028);
xnor U6152 (N_6152,N_4895,N_5055);
and U6153 (N_6153,N_4965,N_4529);
or U6154 (N_6154,N_5643,N_5409);
xnor U6155 (N_6155,N_4747,N_5914);
and U6156 (N_6156,N_5564,N_4663);
nand U6157 (N_6157,N_5521,N_5019);
nor U6158 (N_6158,N_5356,N_5269);
or U6159 (N_6159,N_4553,N_5868);
nand U6160 (N_6160,N_5373,N_5268);
xor U6161 (N_6161,N_4516,N_5678);
xnor U6162 (N_6162,N_4833,N_5135);
nor U6163 (N_6163,N_5906,N_4634);
and U6164 (N_6164,N_5192,N_5178);
xor U6165 (N_6165,N_5897,N_4870);
nor U6166 (N_6166,N_5189,N_5783);
or U6167 (N_6167,N_5847,N_5572);
or U6168 (N_6168,N_5892,N_4562);
xnor U6169 (N_6169,N_4941,N_5705);
xor U6170 (N_6170,N_4945,N_4597);
and U6171 (N_6171,N_4523,N_4640);
or U6172 (N_6172,N_5259,N_4809);
or U6173 (N_6173,N_4514,N_5585);
or U6174 (N_6174,N_5366,N_4899);
nand U6175 (N_6175,N_5383,N_5341);
nor U6176 (N_6176,N_5535,N_5147);
nand U6177 (N_6177,N_4763,N_5821);
nand U6178 (N_6178,N_5416,N_5266);
or U6179 (N_6179,N_4617,N_5798);
or U6180 (N_6180,N_4693,N_5318);
nand U6181 (N_6181,N_5575,N_5492);
and U6182 (N_6182,N_4594,N_4901);
nand U6183 (N_6183,N_5909,N_5674);
nand U6184 (N_6184,N_4649,N_5172);
xnor U6185 (N_6185,N_5507,N_4936);
nand U6186 (N_6186,N_5780,N_5944);
and U6187 (N_6187,N_5874,N_5838);
nor U6188 (N_6188,N_5765,N_5827);
nand U6189 (N_6189,N_5002,N_4510);
nand U6190 (N_6190,N_5540,N_5953);
nor U6191 (N_6191,N_5673,N_5881);
xor U6192 (N_6192,N_4882,N_4616);
nor U6193 (N_6193,N_5258,N_5653);
or U6194 (N_6194,N_5853,N_4559);
xnor U6195 (N_6195,N_5328,N_5916);
xnor U6196 (N_6196,N_4509,N_4842);
or U6197 (N_6197,N_5947,N_5134);
or U6198 (N_6198,N_4607,N_5360);
nand U6199 (N_6199,N_5374,N_4788);
nand U6200 (N_6200,N_5888,N_5831);
or U6201 (N_6201,N_4609,N_4979);
nor U6202 (N_6202,N_5896,N_5246);
xor U6203 (N_6203,N_4807,N_5536);
nand U6204 (N_6204,N_5327,N_5402);
or U6205 (N_6205,N_5981,N_5464);
nand U6206 (N_6206,N_5964,N_5665);
or U6207 (N_6207,N_4839,N_5162);
nor U6208 (N_6208,N_5647,N_5950);
or U6209 (N_6209,N_4632,N_4651);
nand U6210 (N_6210,N_4697,N_4950);
nor U6211 (N_6211,N_5292,N_4641);
nor U6212 (N_6212,N_5792,N_5128);
or U6213 (N_6213,N_5949,N_5784);
nand U6214 (N_6214,N_5320,N_5260);
xor U6215 (N_6215,N_5752,N_4907);
xor U6216 (N_6216,N_5675,N_5197);
and U6217 (N_6217,N_4787,N_5852);
nor U6218 (N_6218,N_4611,N_4623);
nor U6219 (N_6219,N_5113,N_4977);
or U6220 (N_6220,N_5850,N_5543);
and U6221 (N_6221,N_4690,N_5468);
or U6222 (N_6222,N_5412,N_5733);
or U6223 (N_6223,N_5597,N_5542);
or U6224 (N_6224,N_5486,N_5895);
or U6225 (N_6225,N_5701,N_5984);
nand U6226 (N_6226,N_4624,N_5307);
or U6227 (N_6227,N_5904,N_4532);
xor U6228 (N_6228,N_4513,N_5774);
or U6229 (N_6229,N_5805,N_4911);
and U6230 (N_6230,N_5309,N_5697);
nor U6231 (N_6231,N_5736,N_5771);
xnor U6232 (N_6232,N_5484,N_5302);
xor U6233 (N_6233,N_5689,N_5877);
xor U6234 (N_6234,N_5208,N_5668);
xor U6235 (N_6235,N_5865,N_5317);
and U6236 (N_6236,N_4863,N_4531);
xnor U6237 (N_6237,N_4940,N_4832);
nand U6238 (N_6238,N_4962,N_5119);
nand U6239 (N_6239,N_4985,N_5435);
and U6240 (N_6240,N_4955,N_5742);
and U6241 (N_6241,N_5980,N_5957);
and U6242 (N_6242,N_4635,N_5620);
nand U6243 (N_6243,N_4935,N_5207);
nand U6244 (N_6244,N_5174,N_5384);
nor U6245 (N_6245,N_5975,N_5960);
and U6246 (N_6246,N_5283,N_4789);
xor U6247 (N_6247,N_4800,N_4761);
nand U6248 (N_6248,N_5641,N_5796);
xor U6249 (N_6249,N_4544,N_5245);
and U6250 (N_6250,N_5081,N_5794);
nor U6251 (N_6251,N_5867,N_5277);
nand U6252 (N_6252,N_5096,N_5015);
nor U6253 (N_6253,N_5310,N_5104);
nor U6254 (N_6254,N_4733,N_5143);
nor U6255 (N_6255,N_4908,N_4563);
and U6256 (N_6256,N_4518,N_5691);
or U6257 (N_6257,N_4992,N_5854);
xnor U6258 (N_6258,N_5661,N_5672);
or U6259 (N_6259,N_5862,N_5358);
or U6260 (N_6260,N_4837,N_4949);
xnor U6261 (N_6261,N_4710,N_5154);
or U6262 (N_6262,N_5476,N_5680);
and U6263 (N_6263,N_5325,N_5429);
nor U6264 (N_6264,N_4917,N_5052);
nor U6265 (N_6265,N_5525,N_5681);
or U6266 (N_6266,N_5403,N_4524);
nor U6267 (N_6267,N_5669,N_5959);
nor U6268 (N_6268,N_4628,N_4896);
nor U6269 (N_6269,N_5048,N_5629);
nor U6270 (N_6270,N_5290,N_5879);
xor U6271 (N_6271,N_5815,N_5621);
and U6272 (N_6272,N_5244,N_4914);
nor U6273 (N_6273,N_4696,N_5921);
nor U6274 (N_6274,N_5334,N_4862);
nor U6275 (N_6275,N_5241,N_5910);
and U6276 (N_6276,N_5042,N_5010);
and U6277 (N_6277,N_5711,N_4890);
or U6278 (N_6278,N_5609,N_4673);
and U6279 (N_6279,N_5095,N_5574);
and U6280 (N_6280,N_4764,N_5612);
and U6281 (N_6281,N_4680,N_5397);
nand U6282 (N_6282,N_4980,N_5432);
xor U6283 (N_6283,N_5884,N_5466);
nand U6284 (N_6284,N_5614,N_5876);
xor U6285 (N_6285,N_5075,N_5547);
or U6286 (N_6286,N_4873,N_4589);
or U6287 (N_6287,N_5553,N_4677);
nand U6288 (N_6288,N_5410,N_5658);
and U6289 (N_6289,N_5131,N_5698);
nor U6290 (N_6290,N_4646,N_5508);
xnor U6291 (N_6291,N_4679,N_5801);
nor U6292 (N_6292,N_5299,N_4600);
and U6293 (N_6293,N_5446,N_5004);
and U6294 (N_6294,N_5573,N_5431);
or U6295 (N_6295,N_5518,N_5423);
or U6296 (N_6296,N_4591,N_5676);
nor U6297 (N_6297,N_4806,N_4767);
xnor U6298 (N_6298,N_4885,N_5108);
and U6299 (N_6299,N_5727,N_5140);
or U6300 (N_6300,N_5685,N_5365);
and U6301 (N_6301,N_4834,N_5419);
or U6302 (N_6302,N_5625,N_4618);
nand U6303 (N_6303,N_5436,N_5107);
nor U6304 (N_6304,N_5883,N_5538);
nor U6305 (N_6305,N_5014,N_5100);
and U6306 (N_6306,N_4565,N_4500);
nor U6307 (N_6307,N_5369,N_5996);
and U6308 (N_6308,N_5023,N_4554);
nor U6309 (N_6309,N_4657,N_4526);
nor U6310 (N_6310,N_5164,N_5196);
nor U6311 (N_6311,N_4913,N_4952);
and U6312 (N_6312,N_4969,N_5463);
xor U6313 (N_6313,N_4626,N_5322);
and U6314 (N_6314,N_5770,N_5594);
or U6315 (N_6315,N_5869,N_5426);
or U6316 (N_6316,N_5552,N_4879);
nand U6317 (N_6317,N_5159,N_5039);
nand U6318 (N_6318,N_5782,N_5282);
and U6319 (N_6319,N_4934,N_5206);
nand U6320 (N_6320,N_5840,N_4999);
and U6321 (N_6321,N_5300,N_5512);
nand U6322 (N_6322,N_5746,N_4860);
nand U6323 (N_6323,N_5080,N_5942);
nor U6324 (N_6324,N_4822,N_5008);
and U6325 (N_6325,N_4735,N_5450);
xor U6326 (N_6326,N_5662,N_5702);
or U6327 (N_6327,N_5082,N_5841);
and U6328 (N_6328,N_4743,N_5237);
nor U6329 (N_6329,N_5533,N_4570);
and U6330 (N_6330,N_5461,N_4757);
nand U6331 (N_6331,N_5452,N_5166);
and U6332 (N_6332,N_5123,N_5537);
and U6333 (N_6333,N_4701,N_5554);
nand U6334 (N_6334,N_5901,N_5393);
and U6335 (N_6335,N_5929,N_5265);
or U6336 (N_6336,N_4984,N_5779);
xnor U6337 (N_6337,N_4675,N_5205);
and U6338 (N_6338,N_4539,N_4943);
or U6339 (N_6339,N_5640,N_4843);
and U6340 (N_6340,N_5875,N_5938);
xor U6341 (N_6341,N_4550,N_5769);
xnor U6342 (N_6342,N_5546,N_5655);
xnor U6343 (N_6343,N_5242,N_4801);
xor U6344 (N_6344,N_5279,N_5132);
or U6345 (N_6345,N_5997,N_5441);
xnor U6346 (N_6346,N_5990,N_4904);
nand U6347 (N_6347,N_4527,N_5489);
nor U6348 (N_6348,N_5839,N_4674);
or U6349 (N_6349,N_5962,N_4861);
xnor U6350 (N_6350,N_5120,N_5927);
nor U6351 (N_6351,N_5731,N_5891);
nand U6352 (N_6352,N_5047,N_5351);
or U6353 (N_6353,N_5870,N_5009);
and U6354 (N_6354,N_5642,N_5556);
xnor U6355 (N_6355,N_5578,N_5557);
or U6356 (N_6356,N_5064,N_5011);
xnor U6357 (N_6357,N_5362,N_4515);
or U6358 (N_6358,N_5515,N_5830);
and U6359 (N_6359,N_4869,N_5523);
xor U6360 (N_6360,N_5224,N_5005);
or U6361 (N_6361,N_5528,N_5584);
nor U6362 (N_6362,N_5846,N_5755);
or U6363 (N_6363,N_5871,N_5487);
nor U6364 (N_6364,N_5730,N_5966);
xor U6365 (N_6365,N_5298,N_4840);
nor U6366 (N_6366,N_5355,N_4776);
xor U6367 (N_6367,N_5340,N_5079);
nand U6368 (N_6368,N_5312,N_5186);
and U6369 (N_6369,N_5738,N_4944);
or U6370 (N_6370,N_5301,N_4568);
or U6371 (N_6371,N_5326,N_5606);
nand U6372 (N_6372,N_4902,N_4853);
or U6373 (N_6373,N_5091,N_4771);
nand U6374 (N_6374,N_5040,N_5456);
and U6375 (N_6375,N_5024,N_4750);
or U6376 (N_6376,N_5855,N_5018);
xor U6377 (N_6377,N_5229,N_5591);
or U6378 (N_6378,N_4878,N_5762);
and U6379 (N_6379,N_5045,N_5102);
and U6380 (N_6380,N_4888,N_4723);
nor U6381 (N_6381,N_4541,N_5499);
and U6382 (N_6382,N_5583,N_4717);
nand U6383 (N_6383,N_5656,N_5586);
xnor U6384 (N_6384,N_5994,N_5948);
nand U6385 (N_6385,N_5937,N_4599);
nor U6386 (N_6386,N_5338,N_5034);
or U6387 (N_6387,N_5766,N_4921);
nand U6388 (N_6388,N_5475,N_4780);
and U6389 (N_6389,N_5979,N_4558);
nand U6390 (N_6390,N_5714,N_4580);
or U6391 (N_6391,N_4808,N_4972);
and U6392 (N_6392,N_5013,N_5225);
or U6393 (N_6393,N_4577,N_4713);
nor U6394 (N_6394,N_5988,N_4794);
nand U6395 (N_6395,N_5168,N_4835);
xnor U6396 (N_6396,N_4830,N_5202);
or U6397 (N_6397,N_4762,N_5411);
xnor U6398 (N_6398,N_4749,N_5038);
nor U6399 (N_6399,N_5945,N_5719);
nand U6400 (N_6400,N_5592,N_5741);
xor U6401 (N_6401,N_5032,N_4954);
or U6402 (N_6402,N_5716,N_5566);
nor U6403 (N_6403,N_5396,N_4682);
and U6404 (N_6404,N_5111,N_5764);
nand U6405 (N_6405,N_5634,N_5604);
xor U6406 (N_6406,N_5695,N_5222);
nand U6407 (N_6407,N_5382,N_4810);
or U6408 (N_6408,N_4552,N_4884);
nor U6409 (N_6409,N_5381,N_4647);
and U6410 (N_6410,N_4508,N_5112);
nor U6411 (N_6411,N_4987,N_5458);
nor U6412 (N_6412,N_5003,N_5739);
nor U6413 (N_6413,N_5077,N_5995);
xor U6414 (N_6414,N_5342,N_5063);
nor U6415 (N_6415,N_4708,N_5404);
xor U6416 (N_6416,N_4569,N_5316);
or U6417 (N_6417,N_4929,N_5519);
nand U6418 (N_6418,N_4537,N_5037);
xor U6419 (N_6419,N_5704,N_5933);
and U6420 (N_6420,N_5617,N_5343);
nor U6421 (N_6421,N_4695,N_4953);
nand U6422 (N_6422,N_5607,N_5074);
nand U6423 (N_6423,N_5033,N_4946);
nor U6424 (N_6424,N_5723,N_5886);
and U6425 (N_6425,N_5652,N_4991);
and U6426 (N_6426,N_4636,N_5715);
or U6427 (N_6427,N_4817,N_5370);
nand U6428 (N_6428,N_5083,N_5956);
xor U6429 (N_6429,N_4745,N_5467);
nor U6430 (N_6430,N_5819,N_4989);
nor U6431 (N_6431,N_5804,N_5663);
nor U6432 (N_6432,N_5415,N_5406);
or U6433 (N_6433,N_5199,N_4926);
nand U6434 (N_6434,N_4575,N_4973);
and U6435 (N_6435,N_5598,N_5215);
or U6436 (N_6436,N_4678,N_4755);
nand U6437 (N_6437,N_5337,N_5267);
or U6438 (N_6438,N_4507,N_4968);
or U6439 (N_6439,N_4736,N_5579);
xor U6440 (N_6440,N_5474,N_5666);
and U6441 (N_6441,N_5735,N_4669);
nand U6442 (N_6442,N_5534,N_4981);
xor U6443 (N_6443,N_5918,N_4692);
nor U6444 (N_6444,N_5158,N_4686);
and U6445 (N_6445,N_5932,N_5428);
and U6446 (N_6446,N_4535,N_5099);
nor U6447 (N_6447,N_5967,N_4536);
nor U6448 (N_6448,N_5430,N_5357);
nand U6449 (N_6449,N_5480,N_4933);
and U6450 (N_6450,N_4573,N_5750);
xor U6451 (N_6451,N_5532,N_5387);
or U6452 (N_6452,N_4802,N_5973);
and U6453 (N_6453,N_5398,N_5568);
or U6454 (N_6454,N_5367,N_4815);
and U6455 (N_6455,N_5281,N_5679);
or U6456 (N_6456,N_4742,N_5720);
and U6457 (N_6457,N_5223,N_5085);
nand U6458 (N_6458,N_5455,N_4596);
nand U6459 (N_6459,N_4741,N_4567);
or U6460 (N_6460,N_4820,N_5757);
xor U6461 (N_6461,N_5257,N_5982);
and U6462 (N_6462,N_5737,N_5619);
nor U6463 (N_6463,N_4765,N_4846);
nand U6464 (N_6464,N_4716,N_5262);
and U6465 (N_6465,N_4608,N_4847);
or U6466 (N_6466,N_5150,N_4916);
nand U6467 (N_6467,N_5386,N_4585);
and U6468 (N_6468,N_5763,N_4622);
or U6469 (N_6469,N_4898,N_5781);
nor U6470 (N_6470,N_5577,N_4528);
nor U6471 (N_6471,N_5529,N_5882);
and U6472 (N_6472,N_5031,N_4798);
xnor U6473 (N_6473,N_5115,N_4786);
and U6474 (N_6474,N_5250,N_5728);
nor U6475 (N_6475,N_4923,N_5986);
nand U6476 (N_6476,N_4759,N_5144);
nor U6477 (N_6477,N_5845,N_5864);
nand U6478 (N_6478,N_5503,N_5422);
and U6479 (N_6479,N_5616,N_4848);
nand U6480 (N_6480,N_5116,N_5747);
or U6481 (N_6481,N_5324,N_4930);
nor U6482 (N_6482,N_4782,N_4703);
nand U6483 (N_6483,N_4705,N_4702);
nor U6484 (N_6484,N_5628,N_4856);
and U6485 (N_6485,N_5391,N_5787);
or U6486 (N_6486,N_4849,N_4698);
or U6487 (N_6487,N_5558,N_5093);
and U6488 (N_6488,N_5051,N_4685);
and U6489 (N_6489,N_5118,N_5236);
nand U6490 (N_6490,N_4841,N_5969);
nand U6491 (N_6491,N_4645,N_4738);
nand U6492 (N_6492,N_4792,N_4522);
nor U6493 (N_6493,N_5562,N_5797);
or U6494 (N_6494,N_4828,N_4625);
or U6495 (N_6495,N_5126,N_5703);
xor U6496 (N_6496,N_4845,N_5648);
and U6497 (N_6497,N_5814,N_5353);
and U6498 (N_6498,N_4605,N_5734);
nand U6499 (N_6499,N_5722,N_4996);
and U6500 (N_6500,N_4770,N_5109);
nor U6501 (N_6501,N_5090,N_5513);
nand U6502 (N_6502,N_5122,N_5041);
nor U6503 (N_6503,N_5133,N_5977);
nor U6504 (N_6504,N_4694,N_4939);
nor U6505 (N_6505,N_5270,N_5985);
nor U6506 (N_6506,N_5550,N_5989);
or U6507 (N_6507,N_4865,N_5936);
nor U6508 (N_6508,N_5156,N_5922);
and U6509 (N_6509,N_5243,N_4718);
nor U6510 (N_6510,N_5885,N_4603);
xor U6511 (N_6511,N_5182,N_4561);
xor U6512 (N_6512,N_5006,N_4927);
xor U6513 (N_6513,N_5751,N_4672);
and U6514 (N_6514,N_4604,N_4666);
or U6515 (N_6515,N_5789,N_5350);
xnor U6516 (N_6516,N_4804,N_5314);
or U6517 (N_6517,N_5453,N_4774);
nor U6518 (N_6518,N_4872,N_5725);
nor U6519 (N_6519,N_4683,N_5025);
and U6520 (N_6520,N_5893,N_4688);
nor U6521 (N_6521,N_5191,N_4610);
nand U6522 (N_6522,N_4850,N_4709);
nand U6523 (N_6523,N_4963,N_5683);
nand U6524 (N_6524,N_5440,N_5179);
xnor U6525 (N_6525,N_5447,N_5046);
nor U6526 (N_6526,N_4947,N_5124);
and U6527 (N_6527,N_5602,N_5613);
and U6528 (N_6528,N_4823,N_4503);
nand U6529 (N_6529,N_4781,N_4876);
or U6530 (N_6530,N_4986,N_5371);
xor U6531 (N_6531,N_5151,N_5007);
or U6532 (N_6532,N_4601,N_5127);
nand U6533 (N_6533,N_5836,N_5170);
and U6534 (N_6534,N_5138,N_5823);
nor U6535 (N_6535,N_5076,N_5761);
nor U6536 (N_6536,N_5608,N_5457);
nand U6537 (N_6537,N_4874,N_5527);
and U6538 (N_6538,N_5828,N_4704);
and U6539 (N_6539,N_5917,N_5232);
xor U6540 (N_6540,N_5219,N_4566);
xnor U6541 (N_6541,N_5050,N_4951);
nor U6542 (N_6542,N_5349,N_4960);
nor U6543 (N_6543,N_5333,N_4689);
and U6544 (N_6544,N_4564,N_4825);
xor U6545 (N_6545,N_5745,N_5812);
nand U6546 (N_6546,N_4582,N_5627);
nand U6547 (N_6547,N_5087,N_5029);
and U6548 (N_6548,N_5899,N_5347);
or U6549 (N_6549,N_5443,N_5114);
nor U6550 (N_6550,N_5291,N_5101);
xnor U6551 (N_6551,N_5425,N_5449);
nand U6552 (N_6552,N_5073,N_5417);
nand U6553 (N_6553,N_5346,N_4612);
and U6554 (N_6554,N_4614,N_4581);
xor U6555 (N_6555,N_5303,N_4915);
nand U6556 (N_6556,N_4658,N_5520);
nand U6557 (N_6557,N_4517,N_4920);
nand U6558 (N_6558,N_5495,N_4760);
and U6559 (N_6559,N_4615,N_4665);
nand U6560 (N_6560,N_5717,N_5940);
nand U6561 (N_6561,N_4576,N_5809);
and U6562 (N_6562,N_5618,N_4928);
and U6563 (N_6563,N_4889,N_5105);
nand U6564 (N_6564,N_5599,N_5418);
nand U6565 (N_6565,N_5234,N_5645);
or U6566 (N_6566,N_4644,N_5686);
nand U6567 (N_6567,N_5437,N_4906);
nor U6568 (N_6568,N_4957,N_5485);
nand U6569 (N_6569,N_5498,N_4720);
or U6570 (N_6570,N_4737,N_5555);
or U6571 (N_6571,N_5859,N_5626);
xnor U6572 (N_6572,N_5264,N_5587);
nand U6573 (N_6573,N_5377,N_4512);
and U6574 (N_6574,N_5180,N_5070);
and U6575 (N_6575,N_5834,N_4971);
xor U6576 (N_6576,N_5539,N_4588);
nor U6577 (N_6577,N_5049,N_5610);
and U6578 (N_6578,N_5530,N_5561);
and U6579 (N_6579,N_5754,N_4875);
nor U6580 (N_6580,N_5471,N_4650);
xor U6581 (N_6581,N_5451,N_5590);
xor U6582 (N_6582,N_5813,N_5807);
nor U6583 (N_6583,N_5284,N_5928);
and U6584 (N_6584,N_4892,N_5473);
xor U6585 (N_6585,N_4719,N_5239);
and U6586 (N_6586,N_5424,N_5379);
and U6587 (N_6587,N_5414,N_5571);
xor U6588 (N_6588,N_5667,N_5777);
xnor U6589 (N_6589,N_5306,N_5955);
xor U6590 (N_6590,N_4909,N_5188);
nand U6591 (N_6591,N_5217,N_4859);
nand U6592 (N_6592,N_5588,N_5941);
or U6593 (N_6593,N_5671,N_4549);
or U6594 (N_6594,N_5433,N_5545);
xnor U6595 (N_6595,N_4877,N_4744);
nor U6596 (N_6596,N_5323,N_4966);
nor U6597 (N_6597,N_4867,N_4654);
nand U6598 (N_6598,N_5469,N_5297);
or U6599 (N_6599,N_5803,N_5000);
and U6600 (N_6600,N_5786,N_5332);
or U6601 (N_6601,N_4595,N_5768);
nor U6602 (N_6602,N_5272,N_5155);
or U6603 (N_6603,N_4797,N_5478);
nand U6604 (N_6604,N_4959,N_5253);
nand U6605 (N_6605,N_4868,N_5531);
or U6606 (N_6606,N_5161,N_5632);
nor U6607 (N_6607,N_5413,N_4546);
nand U6608 (N_6608,N_5908,N_4938);
or U6609 (N_6609,N_4655,N_4784);
nand U6610 (N_6610,N_5212,N_5849);
nor U6611 (N_6611,N_5659,N_4667);
nor U6612 (N_6612,N_5330,N_5569);
and U6613 (N_6613,N_4572,N_4852);
xor U6614 (N_6614,N_4732,N_5078);
xnor U6615 (N_6615,N_4919,N_5718);
and U6616 (N_6616,N_5514,N_5304);
nand U6617 (N_6617,N_4883,N_5175);
nor U6618 (N_6618,N_5951,N_5603);
and U6619 (N_6619,N_5842,N_5375);
or U6620 (N_6620,N_5427,N_5806);
xnor U6621 (N_6621,N_5200,N_4501);
nor U6622 (N_6622,N_5732,N_4746);
nand U6623 (N_6623,N_4631,N_5235);
or U6624 (N_6624,N_5744,N_5148);
nor U6625 (N_6625,N_5511,N_5501);
or U6626 (N_6626,N_4894,N_5559);
nor U6627 (N_6627,N_5001,N_4590);
nand U6628 (N_6628,N_5856,N_5952);
nand U6629 (N_6629,N_5121,N_5315);
and U6630 (N_6630,N_5860,N_4768);
xnor U6631 (N_6631,N_5210,N_5707);
xor U6632 (N_6632,N_5894,N_5858);
xnor U6633 (N_6633,N_5308,N_4584);
xor U6634 (N_6634,N_5389,N_5043);
and U6635 (N_6635,N_5560,N_5401);
nor U6636 (N_6636,N_4956,N_5709);
nand U6637 (N_6637,N_5974,N_5354);
nand U6638 (N_6638,N_4997,N_4812);
nand U6639 (N_6639,N_5470,N_4988);
and U6640 (N_6640,N_5694,N_5983);
nand U6641 (N_6641,N_4866,N_5826);
xnor U6642 (N_6642,N_4887,N_4671);
or U6643 (N_6643,N_5067,N_5923);
xnor U6644 (N_6644,N_4816,N_5517);
or U6645 (N_6645,N_4668,N_4754);
nor U6646 (N_6646,N_5271,N_5693);
or U6647 (N_6647,N_5690,N_5726);
and U6648 (N_6648,N_4724,N_5816);
and U6649 (N_6649,N_5791,N_4629);
or U6650 (N_6650,N_5016,N_4790);
xor U6651 (N_6651,N_5339,N_5399);
nand U6652 (N_6652,N_5247,N_5582);
xnor U6653 (N_6653,N_5943,N_5935);
nor U6654 (N_6654,N_5911,N_5776);
and U6655 (N_6655,N_4814,N_5646);
nor U6656 (N_6656,N_5611,N_5296);
xnor U6657 (N_6657,N_4728,N_4994);
or U6658 (N_6658,N_5863,N_5231);
xnor U6659 (N_6659,N_4857,N_4905);
and U6660 (N_6660,N_5345,N_5497);
and U6661 (N_6661,N_5251,N_5516);
and U6662 (N_6662,N_4727,N_5305);
or U6663 (N_6663,N_4831,N_4769);
xnor U6664 (N_6664,N_4766,N_5759);
and U6665 (N_6665,N_5638,N_5240);
xor U6666 (N_6666,N_4993,N_5459);
and U6667 (N_6667,N_4504,N_4886);
xnor U6668 (N_6668,N_5364,N_5992);
xor U6669 (N_6669,N_5092,N_4785);
nor U6670 (N_6670,N_5195,N_5335);
nor U6671 (N_6671,N_5905,N_4505);
and U6672 (N_6672,N_5103,N_5713);
nand U6673 (N_6673,N_5615,N_5758);
nor U6674 (N_6674,N_5136,N_5832);
nor U6675 (N_6675,N_5998,N_5946);
or U6676 (N_6676,N_4583,N_5395);
xnor U6677 (N_6677,N_4880,N_4511);
nand U6678 (N_6678,N_5810,N_5491);
and U6679 (N_6679,N_5724,N_5811);
nand U6680 (N_6680,N_5913,N_4813);
or U6681 (N_6681,N_5824,N_5020);
or U6682 (N_6682,N_5488,N_4593);
or U6683 (N_6683,N_4621,N_4598);
nor U6684 (N_6684,N_5177,N_5228);
xor U6685 (N_6685,N_5837,N_5068);
and U6686 (N_6686,N_4592,N_5772);
and U6687 (N_6687,N_4978,N_5567);
nand U6688 (N_6688,N_5285,N_4699);
xor U6689 (N_6689,N_5359,N_4799);
nand U6690 (N_6690,N_5687,N_4534);
and U6691 (N_6691,N_4533,N_4502);
xor U6692 (N_6692,N_5785,N_4551);
or U6693 (N_6693,N_5500,N_4684);
or U6694 (N_6694,N_5420,N_5216);
xor U6695 (N_6695,N_5106,N_5692);
nand U6696 (N_6696,N_5442,N_5851);
or U6697 (N_6697,N_5368,N_5721);
or U6698 (N_6698,N_5623,N_4811);
or U6699 (N_6699,N_5149,N_5551);
nand U6700 (N_6700,N_4998,N_4982);
nor U6701 (N_6701,N_5194,N_4587);
xor U6702 (N_6702,N_4676,N_5059);
nor U6703 (N_6703,N_5249,N_5089);
or U6704 (N_6704,N_4648,N_4805);
nand U6705 (N_6705,N_4925,N_5209);
nand U6706 (N_6706,N_5749,N_5057);
xor U6707 (N_6707,N_5544,N_5263);
xnor U6708 (N_6708,N_5880,N_4967);
nor U6709 (N_6709,N_5187,N_4660);
and U6710 (N_6710,N_4961,N_5226);
and U6711 (N_6711,N_5361,N_5712);
xor U6712 (N_6712,N_5633,N_5563);
and U6713 (N_6713,N_5639,N_5445);
or U6714 (N_6714,N_4638,N_5857);
nand U6715 (N_6715,N_5570,N_5169);
and U6716 (N_6716,N_5472,N_4779);
nor U6717 (N_6717,N_4975,N_4836);
and U6718 (N_6718,N_4739,N_5635);
and U6719 (N_6719,N_4691,N_5275);
nand U6720 (N_6720,N_5125,N_5978);
nand U6721 (N_6721,N_4803,N_4783);
xor U6722 (N_6722,N_4715,N_5061);
nor U6723 (N_6723,N_4932,N_5548);
nand U6724 (N_6724,N_4829,N_5465);
xor U6725 (N_6725,N_4681,N_5993);
nor U6726 (N_6726,N_4543,N_5930);
nand U6727 (N_6727,N_4620,N_5931);
nor U6728 (N_6728,N_5454,N_4606);
or U6729 (N_6729,N_4900,N_4931);
nand U6730 (N_6730,N_5907,N_4824);
xnor U6731 (N_6731,N_5439,N_4948);
or U6732 (N_6732,N_4891,N_4777);
or U6733 (N_6733,N_5644,N_4827);
xor U6734 (N_6734,N_5294,N_4748);
or U6735 (N_6735,N_5185,N_4726);
nor U6736 (N_6736,N_5220,N_5873);
nand U6737 (N_6737,N_4796,N_5524);
nand U6738 (N_6738,N_5872,N_5934);
and U6739 (N_6739,N_4838,N_4851);
or U6740 (N_6740,N_4613,N_5595);
or U6741 (N_6741,N_5204,N_5593);
and U6742 (N_6742,N_5664,N_5589);
and U6743 (N_6743,N_5287,N_5970);
or U6744 (N_6744,N_4560,N_4643);
xnor U6745 (N_6745,N_4818,N_4844);
nand U6746 (N_6746,N_5252,N_5631);
nor U6747 (N_6747,N_5021,N_5903);
nand U6748 (N_6748,N_5999,N_5605);
nor U6749 (N_6749,N_5890,N_5971);
xnor U6750 (N_6750,N_4520,N_5352);
xnor U6751 (N_6751,N_4921,N_4655);
nand U6752 (N_6752,N_4756,N_4814);
or U6753 (N_6753,N_5256,N_5243);
nand U6754 (N_6754,N_5148,N_5307);
xnor U6755 (N_6755,N_4698,N_4915);
or U6756 (N_6756,N_5532,N_5052);
xor U6757 (N_6757,N_5202,N_4733);
nand U6758 (N_6758,N_5881,N_4544);
and U6759 (N_6759,N_5529,N_5661);
nand U6760 (N_6760,N_5841,N_4541);
and U6761 (N_6761,N_5916,N_5670);
xnor U6762 (N_6762,N_4532,N_4660);
or U6763 (N_6763,N_4972,N_5018);
xnor U6764 (N_6764,N_5815,N_5275);
or U6765 (N_6765,N_5933,N_5977);
and U6766 (N_6766,N_5190,N_4502);
and U6767 (N_6767,N_5336,N_5280);
nor U6768 (N_6768,N_5671,N_5568);
xor U6769 (N_6769,N_4687,N_4634);
xor U6770 (N_6770,N_5086,N_5566);
or U6771 (N_6771,N_5147,N_4719);
nor U6772 (N_6772,N_5326,N_5073);
nor U6773 (N_6773,N_5045,N_5779);
xor U6774 (N_6774,N_5687,N_4854);
or U6775 (N_6775,N_5019,N_5520);
xnor U6776 (N_6776,N_4951,N_5266);
xnor U6777 (N_6777,N_5624,N_4818);
xnor U6778 (N_6778,N_5957,N_5211);
nand U6779 (N_6779,N_4614,N_5787);
nor U6780 (N_6780,N_5697,N_4817);
or U6781 (N_6781,N_5952,N_4756);
nand U6782 (N_6782,N_4502,N_4962);
nand U6783 (N_6783,N_4676,N_5984);
nand U6784 (N_6784,N_4971,N_4638);
or U6785 (N_6785,N_4993,N_5330);
nor U6786 (N_6786,N_5195,N_5296);
nor U6787 (N_6787,N_5527,N_5493);
or U6788 (N_6788,N_5390,N_4838);
or U6789 (N_6789,N_5025,N_5709);
xor U6790 (N_6790,N_4953,N_5387);
and U6791 (N_6791,N_5842,N_4627);
or U6792 (N_6792,N_4595,N_4714);
or U6793 (N_6793,N_5024,N_4610);
nor U6794 (N_6794,N_4839,N_5526);
and U6795 (N_6795,N_5584,N_5668);
nand U6796 (N_6796,N_4510,N_5086);
xor U6797 (N_6797,N_4600,N_4651);
and U6798 (N_6798,N_4952,N_5110);
and U6799 (N_6799,N_4852,N_5972);
xnor U6800 (N_6800,N_5908,N_5500);
and U6801 (N_6801,N_5885,N_4951);
or U6802 (N_6802,N_4730,N_5150);
nor U6803 (N_6803,N_5915,N_5640);
or U6804 (N_6804,N_4806,N_5567);
xnor U6805 (N_6805,N_5366,N_5159);
nand U6806 (N_6806,N_4821,N_5585);
and U6807 (N_6807,N_5556,N_5739);
nand U6808 (N_6808,N_4559,N_4761);
nor U6809 (N_6809,N_5155,N_5806);
xor U6810 (N_6810,N_5987,N_5589);
nand U6811 (N_6811,N_5276,N_4668);
and U6812 (N_6812,N_5238,N_5440);
nor U6813 (N_6813,N_5185,N_5601);
xor U6814 (N_6814,N_5825,N_5114);
and U6815 (N_6815,N_5118,N_4534);
or U6816 (N_6816,N_5222,N_4712);
nand U6817 (N_6817,N_5767,N_5740);
nor U6818 (N_6818,N_5710,N_5538);
nand U6819 (N_6819,N_5701,N_5840);
nand U6820 (N_6820,N_5746,N_4969);
and U6821 (N_6821,N_5440,N_5787);
nand U6822 (N_6822,N_5121,N_5650);
and U6823 (N_6823,N_4949,N_5247);
nor U6824 (N_6824,N_4759,N_5388);
xnor U6825 (N_6825,N_4582,N_4693);
nand U6826 (N_6826,N_4593,N_5992);
xnor U6827 (N_6827,N_5959,N_4761);
and U6828 (N_6828,N_5447,N_5640);
nor U6829 (N_6829,N_5437,N_4721);
xnor U6830 (N_6830,N_4730,N_5413);
nand U6831 (N_6831,N_5618,N_5969);
nand U6832 (N_6832,N_5141,N_5143);
nand U6833 (N_6833,N_4532,N_4961);
nor U6834 (N_6834,N_5688,N_5195);
and U6835 (N_6835,N_5600,N_5124);
and U6836 (N_6836,N_5163,N_4530);
nor U6837 (N_6837,N_4951,N_5750);
nor U6838 (N_6838,N_4819,N_5089);
xor U6839 (N_6839,N_5978,N_5078);
nand U6840 (N_6840,N_5293,N_4983);
or U6841 (N_6841,N_4945,N_5275);
and U6842 (N_6842,N_5053,N_5896);
or U6843 (N_6843,N_5765,N_5913);
or U6844 (N_6844,N_5605,N_5564);
and U6845 (N_6845,N_4503,N_5068);
nand U6846 (N_6846,N_4823,N_5211);
or U6847 (N_6847,N_5007,N_4560);
or U6848 (N_6848,N_5288,N_4947);
nor U6849 (N_6849,N_5203,N_5470);
or U6850 (N_6850,N_5971,N_5833);
nor U6851 (N_6851,N_5600,N_5559);
xor U6852 (N_6852,N_5171,N_4571);
or U6853 (N_6853,N_5675,N_5434);
nor U6854 (N_6854,N_5086,N_5949);
nand U6855 (N_6855,N_5695,N_4607);
or U6856 (N_6856,N_5738,N_5480);
or U6857 (N_6857,N_4732,N_5429);
or U6858 (N_6858,N_5967,N_4925);
xnor U6859 (N_6859,N_5362,N_4641);
or U6860 (N_6860,N_4612,N_4697);
and U6861 (N_6861,N_5513,N_5301);
or U6862 (N_6862,N_5819,N_4743);
and U6863 (N_6863,N_4804,N_5761);
and U6864 (N_6864,N_5374,N_4913);
xnor U6865 (N_6865,N_4600,N_4915);
nand U6866 (N_6866,N_5727,N_4599);
nand U6867 (N_6867,N_5450,N_5804);
or U6868 (N_6868,N_4628,N_5812);
nand U6869 (N_6869,N_5163,N_5071);
and U6870 (N_6870,N_4543,N_5181);
nor U6871 (N_6871,N_4868,N_4723);
and U6872 (N_6872,N_4857,N_5345);
xor U6873 (N_6873,N_5619,N_4731);
nor U6874 (N_6874,N_4648,N_5367);
nand U6875 (N_6875,N_5411,N_4532);
nor U6876 (N_6876,N_5299,N_5017);
or U6877 (N_6877,N_4984,N_5285);
or U6878 (N_6878,N_5390,N_5514);
and U6879 (N_6879,N_5629,N_5328);
nor U6880 (N_6880,N_5588,N_5339);
xor U6881 (N_6881,N_4985,N_5565);
xor U6882 (N_6882,N_5180,N_4929);
nand U6883 (N_6883,N_5110,N_4842);
nor U6884 (N_6884,N_5778,N_5145);
nand U6885 (N_6885,N_4666,N_5971);
nand U6886 (N_6886,N_4878,N_4557);
xnor U6887 (N_6887,N_5460,N_5455);
or U6888 (N_6888,N_5844,N_4656);
xor U6889 (N_6889,N_5622,N_5729);
xor U6890 (N_6890,N_5357,N_5087);
nor U6891 (N_6891,N_5512,N_5469);
nor U6892 (N_6892,N_5784,N_5347);
or U6893 (N_6893,N_4886,N_5852);
nor U6894 (N_6894,N_4832,N_4793);
nand U6895 (N_6895,N_5619,N_4658);
nand U6896 (N_6896,N_5584,N_4792);
nand U6897 (N_6897,N_5067,N_5435);
or U6898 (N_6898,N_5470,N_4817);
nor U6899 (N_6899,N_5182,N_5990);
nor U6900 (N_6900,N_5633,N_5766);
and U6901 (N_6901,N_4816,N_4895);
nand U6902 (N_6902,N_5733,N_4537);
nor U6903 (N_6903,N_5793,N_5881);
or U6904 (N_6904,N_4545,N_5456);
nor U6905 (N_6905,N_4972,N_4789);
xnor U6906 (N_6906,N_5119,N_5648);
and U6907 (N_6907,N_5721,N_5388);
and U6908 (N_6908,N_5332,N_5692);
and U6909 (N_6909,N_5190,N_5964);
nand U6910 (N_6910,N_5160,N_5387);
and U6911 (N_6911,N_5396,N_5826);
or U6912 (N_6912,N_4608,N_5710);
xnor U6913 (N_6913,N_5585,N_4565);
and U6914 (N_6914,N_5392,N_5732);
nor U6915 (N_6915,N_4999,N_5110);
or U6916 (N_6916,N_5865,N_4573);
nor U6917 (N_6917,N_5977,N_4871);
and U6918 (N_6918,N_5802,N_5242);
xnor U6919 (N_6919,N_5179,N_4709);
nand U6920 (N_6920,N_5243,N_5166);
or U6921 (N_6921,N_5083,N_4558);
nor U6922 (N_6922,N_5583,N_5628);
nand U6923 (N_6923,N_5568,N_5858);
and U6924 (N_6924,N_4710,N_5582);
and U6925 (N_6925,N_4565,N_5480);
and U6926 (N_6926,N_5696,N_4576);
or U6927 (N_6927,N_5067,N_5716);
and U6928 (N_6928,N_4962,N_4569);
nor U6929 (N_6929,N_4610,N_4741);
nand U6930 (N_6930,N_4796,N_5125);
nand U6931 (N_6931,N_4944,N_4862);
nand U6932 (N_6932,N_5762,N_5751);
nand U6933 (N_6933,N_5371,N_5434);
nor U6934 (N_6934,N_5315,N_5184);
or U6935 (N_6935,N_5980,N_5881);
nand U6936 (N_6936,N_5690,N_4745);
xor U6937 (N_6937,N_4868,N_5374);
nand U6938 (N_6938,N_5039,N_5198);
nand U6939 (N_6939,N_4914,N_5963);
nor U6940 (N_6940,N_4914,N_5262);
nor U6941 (N_6941,N_4922,N_5322);
and U6942 (N_6942,N_5289,N_5212);
xnor U6943 (N_6943,N_5183,N_4689);
nor U6944 (N_6944,N_5896,N_5742);
xnor U6945 (N_6945,N_4703,N_5014);
nor U6946 (N_6946,N_5479,N_4736);
or U6947 (N_6947,N_4745,N_4660);
or U6948 (N_6948,N_4917,N_4552);
and U6949 (N_6949,N_5292,N_5387);
and U6950 (N_6950,N_5386,N_5918);
or U6951 (N_6951,N_5619,N_5655);
nor U6952 (N_6952,N_4768,N_5109);
or U6953 (N_6953,N_4915,N_4564);
nor U6954 (N_6954,N_5559,N_5972);
xnor U6955 (N_6955,N_4806,N_5880);
nand U6956 (N_6956,N_5106,N_5663);
nor U6957 (N_6957,N_5019,N_5922);
nor U6958 (N_6958,N_5099,N_5308);
nand U6959 (N_6959,N_5145,N_5487);
xnor U6960 (N_6960,N_5284,N_4755);
or U6961 (N_6961,N_5509,N_5281);
or U6962 (N_6962,N_5414,N_5218);
and U6963 (N_6963,N_5415,N_5840);
and U6964 (N_6964,N_5124,N_5037);
nor U6965 (N_6965,N_5607,N_5339);
nor U6966 (N_6966,N_5636,N_5338);
nor U6967 (N_6967,N_5416,N_5449);
xnor U6968 (N_6968,N_5590,N_5934);
nor U6969 (N_6969,N_4979,N_4580);
and U6970 (N_6970,N_5813,N_4726);
or U6971 (N_6971,N_5614,N_4906);
nor U6972 (N_6972,N_4845,N_4748);
or U6973 (N_6973,N_4998,N_5430);
xor U6974 (N_6974,N_4581,N_5445);
nand U6975 (N_6975,N_5271,N_5215);
nor U6976 (N_6976,N_5454,N_5834);
or U6977 (N_6977,N_5639,N_4757);
and U6978 (N_6978,N_4765,N_5431);
nand U6979 (N_6979,N_5712,N_5561);
or U6980 (N_6980,N_5620,N_5290);
and U6981 (N_6981,N_5834,N_4806);
and U6982 (N_6982,N_4748,N_5002);
nor U6983 (N_6983,N_5576,N_5823);
nand U6984 (N_6984,N_4795,N_5999);
or U6985 (N_6985,N_5943,N_5735);
or U6986 (N_6986,N_5558,N_5965);
xnor U6987 (N_6987,N_4557,N_4915);
or U6988 (N_6988,N_5578,N_4537);
nand U6989 (N_6989,N_5328,N_5454);
and U6990 (N_6990,N_5666,N_4933);
and U6991 (N_6991,N_5967,N_4873);
nand U6992 (N_6992,N_4850,N_5459);
and U6993 (N_6993,N_5050,N_4572);
and U6994 (N_6994,N_5962,N_5684);
nor U6995 (N_6995,N_5959,N_5216);
nand U6996 (N_6996,N_4950,N_5586);
nand U6997 (N_6997,N_5162,N_5697);
or U6998 (N_6998,N_5203,N_5512);
or U6999 (N_6999,N_5253,N_5044);
or U7000 (N_7000,N_5786,N_4577);
nor U7001 (N_7001,N_5151,N_5455);
nor U7002 (N_7002,N_4522,N_5901);
nor U7003 (N_7003,N_5196,N_4966);
or U7004 (N_7004,N_5411,N_5696);
nand U7005 (N_7005,N_5742,N_5163);
or U7006 (N_7006,N_5499,N_5925);
or U7007 (N_7007,N_5516,N_5124);
xnor U7008 (N_7008,N_5152,N_5689);
nand U7009 (N_7009,N_5515,N_5581);
xnor U7010 (N_7010,N_4761,N_5525);
nand U7011 (N_7011,N_5797,N_4909);
nand U7012 (N_7012,N_5065,N_4687);
and U7013 (N_7013,N_4621,N_5503);
and U7014 (N_7014,N_5752,N_4945);
xnor U7015 (N_7015,N_4795,N_5147);
and U7016 (N_7016,N_5991,N_5286);
xnor U7017 (N_7017,N_4554,N_4520);
xnor U7018 (N_7018,N_5396,N_5268);
or U7019 (N_7019,N_5089,N_5004);
or U7020 (N_7020,N_5792,N_4841);
nand U7021 (N_7021,N_5750,N_5859);
nor U7022 (N_7022,N_4613,N_5941);
or U7023 (N_7023,N_5489,N_4640);
or U7024 (N_7024,N_4527,N_5678);
nor U7025 (N_7025,N_4609,N_5053);
or U7026 (N_7026,N_5734,N_4635);
nand U7027 (N_7027,N_4729,N_5974);
or U7028 (N_7028,N_4530,N_5371);
and U7029 (N_7029,N_4564,N_5226);
xor U7030 (N_7030,N_5709,N_5612);
nor U7031 (N_7031,N_4602,N_5630);
and U7032 (N_7032,N_4795,N_4613);
and U7033 (N_7033,N_4752,N_5300);
or U7034 (N_7034,N_4693,N_5786);
or U7035 (N_7035,N_4727,N_5667);
and U7036 (N_7036,N_4561,N_4923);
nor U7037 (N_7037,N_5717,N_5962);
or U7038 (N_7038,N_5206,N_5440);
and U7039 (N_7039,N_4847,N_4661);
nand U7040 (N_7040,N_5143,N_4669);
xnor U7041 (N_7041,N_5906,N_5367);
or U7042 (N_7042,N_5281,N_5399);
nand U7043 (N_7043,N_5261,N_5845);
nor U7044 (N_7044,N_5189,N_5728);
nand U7045 (N_7045,N_5677,N_5276);
nand U7046 (N_7046,N_5037,N_5705);
and U7047 (N_7047,N_5721,N_4956);
and U7048 (N_7048,N_4695,N_5126);
nor U7049 (N_7049,N_4799,N_5757);
nor U7050 (N_7050,N_5653,N_4762);
and U7051 (N_7051,N_4934,N_5010);
or U7052 (N_7052,N_5567,N_5254);
nor U7053 (N_7053,N_5566,N_4764);
or U7054 (N_7054,N_5702,N_5274);
and U7055 (N_7055,N_4873,N_5174);
or U7056 (N_7056,N_5547,N_4528);
nor U7057 (N_7057,N_4821,N_5707);
or U7058 (N_7058,N_4864,N_5578);
or U7059 (N_7059,N_4757,N_5898);
nor U7060 (N_7060,N_4921,N_5366);
xnor U7061 (N_7061,N_5833,N_5362);
nand U7062 (N_7062,N_5412,N_5812);
xor U7063 (N_7063,N_5493,N_5609);
or U7064 (N_7064,N_4517,N_5378);
xnor U7065 (N_7065,N_4580,N_5247);
xor U7066 (N_7066,N_5242,N_5331);
nand U7067 (N_7067,N_5551,N_5076);
or U7068 (N_7068,N_4984,N_5897);
nor U7069 (N_7069,N_5447,N_5851);
nand U7070 (N_7070,N_5365,N_5334);
or U7071 (N_7071,N_5920,N_5115);
and U7072 (N_7072,N_4716,N_4818);
xnor U7073 (N_7073,N_5329,N_5850);
xor U7074 (N_7074,N_5651,N_5307);
nor U7075 (N_7075,N_4837,N_5537);
or U7076 (N_7076,N_5672,N_5139);
nand U7077 (N_7077,N_5875,N_4857);
nand U7078 (N_7078,N_5561,N_5113);
or U7079 (N_7079,N_5261,N_5876);
and U7080 (N_7080,N_4872,N_5720);
xor U7081 (N_7081,N_5637,N_4929);
or U7082 (N_7082,N_5946,N_5997);
and U7083 (N_7083,N_5494,N_5862);
and U7084 (N_7084,N_5908,N_5406);
and U7085 (N_7085,N_5474,N_4625);
nand U7086 (N_7086,N_4843,N_4609);
nand U7087 (N_7087,N_4983,N_5627);
nand U7088 (N_7088,N_4974,N_4849);
xor U7089 (N_7089,N_5784,N_4849);
nand U7090 (N_7090,N_5892,N_5506);
or U7091 (N_7091,N_5361,N_4624);
xnor U7092 (N_7092,N_4812,N_4964);
nor U7093 (N_7093,N_5077,N_5356);
or U7094 (N_7094,N_5583,N_5514);
and U7095 (N_7095,N_5405,N_5585);
xor U7096 (N_7096,N_4549,N_5252);
nor U7097 (N_7097,N_5672,N_4949);
or U7098 (N_7098,N_4771,N_4937);
nand U7099 (N_7099,N_4837,N_5213);
or U7100 (N_7100,N_5020,N_4608);
and U7101 (N_7101,N_4698,N_5532);
nand U7102 (N_7102,N_5909,N_5833);
xnor U7103 (N_7103,N_5131,N_4755);
nor U7104 (N_7104,N_4741,N_5433);
nor U7105 (N_7105,N_4960,N_4809);
nor U7106 (N_7106,N_5976,N_4922);
or U7107 (N_7107,N_4969,N_5156);
or U7108 (N_7108,N_5080,N_5711);
nand U7109 (N_7109,N_4507,N_5774);
or U7110 (N_7110,N_5425,N_5555);
or U7111 (N_7111,N_4825,N_5280);
or U7112 (N_7112,N_5935,N_5807);
and U7113 (N_7113,N_4945,N_5348);
and U7114 (N_7114,N_5986,N_5384);
or U7115 (N_7115,N_5419,N_5407);
nand U7116 (N_7116,N_5741,N_5568);
and U7117 (N_7117,N_5552,N_5241);
or U7118 (N_7118,N_5642,N_4565);
or U7119 (N_7119,N_5012,N_5152);
nand U7120 (N_7120,N_4582,N_5739);
and U7121 (N_7121,N_5051,N_4810);
and U7122 (N_7122,N_5791,N_4982);
nand U7123 (N_7123,N_5323,N_5945);
nand U7124 (N_7124,N_5672,N_4831);
nor U7125 (N_7125,N_5807,N_4720);
or U7126 (N_7126,N_4771,N_4708);
and U7127 (N_7127,N_5751,N_5358);
xnor U7128 (N_7128,N_4679,N_4611);
or U7129 (N_7129,N_4896,N_5323);
nor U7130 (N_7130,N_4713,N_5525);
nand U7131 (N_7131,N_5513,N_4603);
and U7132 (N_7132,N_5291,N_5942);
or U7133 (N_7133,N_5992,N_5639);
and U7134 (N_7134,N_5493,N_5091);
and U7135 (N_7135,N_5826,N_5741);
nor U7136 (N_7136,N_5850,N_5941);
or U7137 (N_7137,N_4591,N_5321);
and U7138 (N_7138,N_4630,N_5085);
nand U7139 (N_7139,N_5437,N_5480);
nor U7140 (N_7140,N_5497,N_4993);
nand U7141 (N_7141,N_4529,N_4921);
xor U7142 (N_7142,N_4500,N_5637);
nand U7143 (N_7143,N_5342,N_5538);
xnor U7144 (N_7144,N_5323,N_5000);
or U7145 (N_7145,N_4887,N_4731);
nand U7146 (N_7146,N_5407,N_5297);
nor U7147 (N_7147,N_4947,N_5584);
xnor U7148 (N_7148,N_5202,N_5568);
or U7149 (N_7149,N_4851,N_5886);
xnor U7150 (N_7150,N_5787,N_5457);
nor U7151 (N_7151,N_5198,N_4830);
xor U7152 (N_7152,N_5794,N_5021);
and U7153 (N_7153,N_5621,N_4594);
nand U7154 (N_7154,N_5958,N_5931);
xnor U7155 (N_7155,N_5689,N_5993);
nand U7156 (N_7156,N_5809,N_4726);
xnor U7157 (N_7157,N_5047,N_5839);
and U7158 (N_7158,N_5598,N_5832);
xnor U7159 (N_7159,N_5967,N_5770);
nand U7160 (N_7160,N_5193,N_4682);
nor U7161 (N_7161,N_5452,N_5712);
and U7162 (N_7162,N_5348,N_4989);
nand U7163 (N_7163,N_4790,N_5676);
nor U7164 (N_7164,N_5486,N_5663);
or U7165 (N_7165,N_5930,N_5961);
nand U7166 (N_7166,N_5409,N_5497);
nand U7167 (N_7167,N_4564,N_5332);
xnor U7168 (N_7168,N_5048,N_5535);
nor U7169 (N_7169,N_5956,N_4577);
xnor U7170 (N_7170,N_4536,N_5172);
xnor U7171 (N_7171,N_4519,N_5320);
nand U7172 (N_7172,N_4645,N_5757);
nand U7173 (N_7173,N_4940,N_5710);
xor U7174 (N_7174,N_4676,N_5062);
nor U7175 (N_7175,N_5988,N_5837);
and U7176 (N_7176,N_5398,N_5750);
and U7177 (N_7177,N_5845,N_4738);
xnor U7178 (N_7178,N_5206,N_4688);
or U7179 (N_7179,N_5711,N_5138);
and U7180 (N_7180,N_5592,N_4539);
nand U7181 (N_7181,N_4980,N_4602);
nand U7182 (N_7182,N_5863,N_5712);
nor U7183 (N_7183,N_4540,N_5860);
nand U7184 (N_7184,N_4805,N_5561);
xnor U7185 (N_7185,N_4724,N_4696);
nor U7186 (N_7186,N_4602,N_5680);
or U7187 (N_7187,N_5455,N_4593);
or U7188 (N_7188,N_5132,N_5531);
nand U7189 (N_7189,N_4913,N_5497);
or U7190 (N_7190,N_5603,N_5644);
nand U7191 (N_7191,N_5055,N_5869);
xor U7192 (N_7192,N_5925,N_5049);
xor U7193 (N_7193,N_5684,N_5700);
xnor U7194 (N_7194,N_5106,N_5570);
and U7195 (N_7195,N_5258,N_4716);
xor U7196 (N_7196,N_5678,N_5675);
xor U7197 (N_7197,N_5738,N_4559);
xnor U7198 (N_7198,N_5824,N_5116);
or U7199 (N_7199,N_5292,N_5247);
xor U7200 (N_7200,N_5232,N_5423);
or U7201 (N_7201,N_5937,N_4931);
or U7202 (N_7202,N_5257,N_5335);
xnor U7203 (N_7203,N_5180,N_5694);
nand U7204 (N_7204,N_4549,N_5367);
nand U7205 (N_7205,N_5622,N_5258);
or U7206 (N_7206,N_5899,N_5045);
and U7207 (N_7207,N_5770,N_5075);
or U7208 (N_7208,N_5581,N_5896);
nor U7209 (N_7209,N_5462,N_5510);
xnor U7210 (N_7210,N_5325,N_5263);
xnor U7211 (N_7211,N_5466,N_4922);
or U7212 (N_7212,N_5939,N_5096);
nand U7213 (N_7213,N_5367,N_5345);
or U7214 (N_7214,N_4589,N_5342);
nor U7215 (N_7215,N_5972,N_4983);
or U7216 (N_7216,N_5482,N_5250);
xor U7217 (N_7217,N_5269,N_5372);
or U7218 (N_7218,N_5733,N_4865);
and U7219 (N_7219,N_5586,N_4710);
or U7220 (N_7220,N_5446,N_5366);
or U7221 (N_7221,N_5351,N_4726);
nor U7222 (N_7222,N_5198,N_5230);
and U7223 (N_7223,N_4592,N_5271);
nand U7224 (N_7224,N_4510,N_5055);
xor U7225 (N_7225,N_4848,N_5645);
or U7226 (N_7226,N_5047,N_5423);
nor U7227 (N_7227,N_5267,N_4986);
or U7228 (N_7228,N_5925,N_5560);
nand U7229 (N_7229,N_5224,N_5222);
nor U7230 (N_7230,N_4991,N_4762);
or U7231 (N_7231,N_5446,N_5593);
nand U7232 (N_7232,N_5336,N_5558);
or U7233 (N_7233,N_5652,N_5067);
or U7234 (N_7234,N_4686,N_5416);
nor U7235 (N_7235,N_5607,N_5835);
nand U7236 (N_7236,N_5286,N_5317);
nand U7237 (N_7237,N_5957,N_5837);
nand U7238 (N_7238,N_5679,N_4798);
nor U7239 (N_7239,N_5529,N_5165);
nor U7240 (N_7240,N_5675,N_5350);
nor U7241 (N_7241,N_4998,N_5939);
and U7242 (N_7242,N_5101,N_5745);
or U7243 (N_7243,N_5410,N_4782);
and U7244 (N_7244,N_5883,N_4821);
and U7245 (N_7245,N_5400,N_4685);
nand U7246 (N_7246,N_5972,N_4549);
and U7247 (N_7247,N_5288,N_5696);
and U7248 (N_7248,N_4640,N_5042);
and U7249 (N_7249,N_4961,N_4812);
nor U7250 (N_7250,N_4721,N_4802);
nand U7251 (N_7251,N_5266,N_4589);
nand U7252 (N_7252,N_4742,N_5682);
xnor U7253 (N_7253,N_5862,N_5458);
xor U7254 (N_7254,N_4778,N_5087);
or U7255 (N_7255,N_5080,N_5092);
nand U7256 (N_7256,N_5099,N_5640);
nand U7257 (N_7257,N_4688,N_4764);
nor U7258 (N_7258,N_5960,N_4952);
and U7259 (N_7259,N_5042,N_4595);
nand U7260 (N_7260,N_5427,N_5421);
nand U7261 (N_7261,N_5668,N_4579);
nand U7262 (N_7262,N_4718,N_4750);
nor U7263 (N_7263,N_4740,N_5729);
or U7264 (N_7264,N_4570,N_5821);
nor U7265 (N_7265,N_5067,N_4928);
nor U7266 (N_7266,N_4759,N_5241);
xor U7267 (N_7267,N_4673,N_4861);
xnor U7268 (N_7268,N_5836,N_5602);
nand U7269 (N_7269,N_4750,N_5201);
or U7270 (N_7270,N_5948,N_4840);
xor U7271 (N_7271,N_5739,N_5133);
xor U7272 (N_7272,N_5814,N_5462);
xor U7273 (N_7273,N_5272,N_4818);
nor U7274 (N_7274,N_5272,N_5832);
or U7275 (N_7275,N_4785,N_5838);
nor U7276 (N_7276,N_5910,N_4700);
nor U7277 (N_7277,N_5096,N_5558);
nand U7278 (N_7278,N_5455,N_5834);
xnor U7279 (N_7279,N_4729,N_4976);
nor U7280 (N_7280,N_5230,N_5959);
xor U7281 (N_7281,N_5387,N_5715);
and U7282 (N_7282,N_5686,N_4533);
nand U7283 (N_7283,N_4604,N_5034);
or U7284 (N_7284,N_4779,N_5581);
xnor U7285 (N_7285,N_5186,N_5431);
nand U7286 (N_7286,N_4812,N_4893);
nand U7287 (N_7287,N_4973,N_4783);
and U7288 (N_7288,N_5972,N_4748);
and U7289 (N_7289,N_5088,N_4547);
xor U7290 (N_7290,N_4629,N_4748);
or U7291 (N_7291,N_5850,N_5122);
nand U7292 (N_7292,N_5635,N_4720);
nand U7293 (N_7293,N_4808,N_5363);
or U7294 (N_7294,N_5387,N_5988);
or U7295 (N_7295,N_5755,N_4961);
xor U7296 (N_7296,N_5182,N_4866);
and U7297 (N_7297,N_4698,N_5835);
or U7298 (N_7298,N_5699,N_5501);
and U7299 (N_7299,N_5613,N_5141);
and U7300 (N_7300,N_5882,N_4741);
and U7301 (N_7301,N_4830,N_5420);
xnor U7302 (N_7302,N_5276,N_4693);
xor U7303 (N_7303,N_4741,N_5315);
xor U7304 (N_7304,N_5616,N_5825);
nand U7305 (N_7305,N_5396,N_5031);
nand U7306 (N_7306,N_5992,N_5697);
or U7307 (N_7307,N_4855,N_5005);
or U7308 (N_7308,N_5622,N_4742);
or U7309 (N_7309,N_5236,N_5515);
and U7310 (N_7310,N_5649,N_4540);
and U7311 (N_7311,N_5559,N_5282);
or U7312 (N_7312,N_5274,N_5158);
xor U7313 (N_7313,N_5662,N_5660);
nor U7314 (N_7314,N_5054,N_5003);
nor U7315 (N_7315,N_5120,N_4530);
or U7316 (N_7316,N_5206,N_4795);
or U7317 (N_7317,N_5643,N_4587);
or U7318 (N_7318,N_4752,N_5942);
and U7319 (N_7319,N_5992,N_5540);
xnor U7320 (N_7320,N_5472,N_5501);
and U7321 (N_7321,N_4834,N_5331);
xnor U7322 (N_7322,N_4620,N_4734);
nand U7323 (N_7323,N_5065,N_5146);
nor U7324 (N_7324,N_5540,N_5421);
nor U7325 (N_7325,N_5797,N_5117);
or U7326 (N_7326,N_5633,N_4585);
or U7327 (N_7327,N_5607,N_5583);
and U7328 (N_7328,N_4826,N_4913);
xor U7329 (N_7329,N_5723,N_5007);
nor U7330 (N_7330,N_5056,N_5172);
or U7331 (N_7331,N_4808,N_5045);
xor U7332 (N_7332,N_5519,N_5318);
nand U7333 (N_7333,N_5032,N_5420);
or U7334 (N_7334,N_4949,N_4858);
or U7335 (N_7335,N_5323,N_5706);
xnor U7336 (N_7336,N_4537,N_5808);
nand U7337 (N_7337,N_4859,N_5947);
or U7338 (N_7338,N_5538,N_4999);
and U7339 (N_7339,N_5478,N_5612);
nand U7340 (N_7340,N_4903,N_4805);
and U7341 (N_7341,N_4659,N_5542);
xor U7342 (N_7342,N_4550,N_5334);
and U7343 (N_7343,N_4727,N_4783);
xnor U7344 (N_7344,N_4801,N_4723);
and U7345 (N_7345,N_5712,N_5358);
xnor U7346 (N_7346,N_4991,N_4960);
and U7347 (N_7347,N_4664,N_4699);
nor U7348 (N_7348,N_4612,N_5380);
nor U7349 (N_7349,N_5769,N_5074);
and U7350 (N_7350,N_5182,N_5920);
xor U7351 (N_7351,N_4983,N_4745);
and U7352 (N_7352,N_5114,N_5318);
and U7353 (N_7353,N_5082,N_5442);
xnor U7354 (N_7354,N_4709,N_5132);
nand U7355 (N_7355,N_5212,N_5613);
nand U7356 (N_7356,N_5077,N_4863);
or U7357 (N_7357,N_5077,N_5766);
nand U7358 (N_7358,N_5095,N_5330);
xor U7359 (N_7359,N_4930,N_4978);
xnor U7360 (N_7360,N_5189,N_5584);
xnor U7361 (N_7361,N_5285,N_4973);
nand U7362 (N_7362,N_4815,N_5487);
and U7363 (N_7363,N_4780,N_4747);
xnor U7364 (N_7364,N_4925,N_5797);
and U7365 (N_7365,N_4879,N_5606);
and U7366 (N_7366,N_5532,N_5933);
and U7367 (N_7367,N_5272,N_5510);
and U7368 (N_7368,N_5451,N_5954);
nor U7369 (N_7369,N_5060,N_5484);
or U7370 (N_7370,N_5073,N_5941);
or U7371 (N_7371,N_5012,N_5667);
nand U7372 (N_7372,N_4863,N_5900);
or U7373 (N_7373,N_5822,N_4819);
nor U7374 (N_7374,N_4928,N_5037);
nand U7375 (N_7375,N_5273,N_4786);
or U7376 (N_7376,N_5265,N_4558);
and U7377 (N_7377,N_5645,N_5538);
or U7378 (N_7378,N_5412,N_5690);
or U7379 (N_7379,N_5290,N_4900);
nor U7380 (N_7380,N_5932,N_4536);
or U7381 (N_7381,N_5481,N_4902);
nand U7382 (N_7382,N_5223,N_4936);
xnor U7383 (N_7383,N_4893,N_5755);
or U7384 (N_7384,N_5046,N_4983);
nor U7385 (N_7385,N_5050,N_5459);
and U7386 (N_7386,N_5454,N_4767);
nand U7387 (N_7387,N_5733,N_4634);
nand U7388 (N_7388,N_5448,N_5893);
xnor U7389 (N_7389,N_4778,N_5176);
and U7390 (N_7390,N_5291,N_5127);
and U7391 (N_7391,N_5175,N_5947);
nor U7392 (N_7392,N_5256,N_4582);
xnor U7393 (N_7393,N_5537,N_5119);
nand U7394 (N_7394,N_5950,N_5102);
nor U7395 (N_7395,N_5105,N_5450);
xnor U7396 (N_7396,N_5751,N_4693);
nand U7397 (N_7397,N_5912,N_4890);
nor U7398 (N_7398,N_4963,N_5534);
and U7399 (N_7399,N_5426,N_4840);
nor U7400 (N_7400,N_5843,N_4510);
or U7401 (N_7401,N_5553,N_4957);
nand U7402 (N_7402,N_5635,N_5776);
nand U7403 (N_7403,N_4689,N_4664);
and U7404 (N_7404,N_5517,N_5324);
nor U7405 (N_7405,N_4554,N_5693);
xor U7406 (N_7406,N_5495,N_4621);
xnor U7407 (N_7407,N_5535,N_4978);
xor U7408 (N_7408,N_5516,N_5714);
nand U7409 (N_7409,N_4874,N_4659);
xor U7410 (N_7410,N_5673,N_4826);
or U7411 (N_7411,N_5585,N_5434);
and U7412 (N_7412,N_5637,N_5058);
or U7413 (N_7413,N_5064,N_5464);
and U7414 (N_7414,N_5377,N_5237);
or U7415 (N_7415,N_5643,N_4931);
and U7416 (N_7416,N_4955,N_5997);
and U7417 (N_7417,N_5131,N_4771);
nand U7418 (N_7418,N_5724,N_5322);
nand U7419 (N_7419,N_4683,N_4581);
and U7420 (N_7420,N_5376,N_4926);
nand U7421 (N_7421,N_5443,N_5952);
nor U7422 (N_7422,N_5682,N_4943);
nor U7423 (N_7423,N_5768,N_5328);
nor U7424 (N_7424,N_5120,N_5752);
and U7425 (N_7425,N_5681,N_4954);
nor U7426 (N_7426,N_5418,N_4994);
or U7427 (N_7427,N_5044,N_5565);
and U7428 (N_7428,N_4969,N_4559);
nand U7429 (N_7429,N_5006,N_5717);
or U7430 (N_7430,N_4843,N_5277);
nand U7431 (N_7431,N_5164,N_4768);
and U7432 (N_7432,N_5024,N_5028);
xor U7433 (N_7433,N_5978,N_4507);
nor U7434 (N_7434,N_5406,N_5740);
nor U7435 (N_7435,N_4580,N_5910);
nand U7436 (N_7436,N_5631,N_4716);
nor U7437 (N_7437,N_5823,N_4836);
nand U7438 (N_7438,N_5922,N_4750);
and U7439 (N_7439,N_5638,N_5180);
xnor U7440 (N_7440,N_5537,N_5592);
or U7441 (N_7441,N_5965,N_5034);
xor U7442 (N_7442,N_4742,N_5423);
xor U7443 (N_7443,N_5962,N_5969);
nor U7444 (N_7444,N_5867,N_5746);
and U7445 (N_7445,N_5591,N_5498);
and U7446 (N_7446,N_5449,N_5516);
xnor U7447 (N_7447,N_5981,N_5636);
xor U7448 (N_7448,N_5656,N_5323);
xnor U7449 (N_7449,N_5801,N_5258);
and U7450 (N_7450,N_5318,N_5394);
nand U7451 (N_7451,N_4966,N_4553);
or U7452 (N_7452,N_5942,N_4618);
or U7453 (N_7453,N_5030,N_5603);
and U7454 (N_7454,N_4591,N_4993);
nor U7455 (N_7455,N_4870,N_4561);
nand U7456 (N_7456,N_5499,N_5394);
and U7457 (N_7457,N_5199,N_4753);
nor U7458 (N_7458,N_5555,N_5344);
nand U7459 (N_7459,N_5500,N_4535);
nor U7460 (N_7460,N_5442,N_5375);
nand U7461 (N_7461,N_5851,N_4595);
and U7462 (N_7462,N_5881,N_5828);
and U7463 (N_7463,N_5327,N_5062);
xnor U7464 (N_7464,N_5934,N_5402);
xor U7465 (N_7465,N_5650,N_5611);
xor U7466 (N_7466,N_5061,N_5116);
or U7467 (N_7467,N_5528,N_4728);
nor U7468 (N_7468,N_5149,N_5408);
and U7469 (N_7469,N_4624,N_4762);
nor U7470 (N_7470,N_5150,N_5737);
and U7471 (N_7471,N_5094,N_5522);
and U7472 (N_7472,N_5982,N_4563);
nor U7473 (N_7473,N_5204,N_4548);
and U7474 (N_7474,N_5850,N_5364);
nand U7475 (N_7475,N_4656,N_4823);
and U7476 (N_7476,N_5727,N_4710);
or U7477 (N_7477,N_5087,N_4629);
or U7478 (N_7478,N_5940,N_5512);
nor U7479 (N_7479,N_5350,N_5981);
xnor U7480 (N_7480,N_4626,N_4837);
nor U7481 (N_7481,N_5610,N_4923);
xor U7482 (N_7482,N_5847,N_5898);
nand U7483 (N_7483,N_5590,N_5449);
and U7484 (N_7484,N_5893,N_5306);
or U7485 (N_7485,N_5566,N_5700);
or U7486 (N_7486,N_4877,N_5862);
and U7487 (N_7487,N_4630,N_4856);
xor U7488 (N_7488,N_5241,N_5262);
nor U7489 (N_7489,N_4976,N_4501);
or U7490 (N_7490,N_4751,N_5830);
or U7491 (N_7491,N_5791,N_5506);
or U7492 (N_7492,N_4933,N_4970);
or U7493 (N_7493,N_5984,N_5375);
nand U7494 (N_7494,N_5823,N_5893);
nor U7495 (N_7495,N_4734,N_5225);
and U7496 (N_7496,N_4637,N_4730);
or U7497 (N_7497,N_5663,N_4834);
nor U7498 (N_7498,N_5224,N_4533);
nor U7499 (N_7499,N_5474,N_5259);
and U7500 (N_7500,N_6964,N_6310);
nand U7501 (N_7501,N_6565,N_6224);
and U7502 (N_7502,N_6408,N_7150);
nor U7503 (N_7503,N_7312,N_6568);
nor U7504 (N_7504,N_7414,N_6313);
xnor U7505 (N_7505,N_7386,N_6863);
nand U7506 (N_7506,N_6361,N_6115);
xor U7507 (N_7507,N_6033,N_6984);
and U7508 (N_7508,N_7019,N_7056);
xor U7509 (N_7509,N_6810,N_6981);
xor U7510 (N_7510,N_6303,N_7195);
or U7511 (N_7511,N_7253,N_6990);
xnor U7512 (N_7512,N_6692,N_6761);
nor U7513 (N_7513,N_6266,N_6763);
or U7514 (N_7514,N_6782,N_6021);
and U7515 (N_7515,N_7020,N_7445);
xor U7516 (N_7516,N_7130,N_6131);
and U7517 (N_7517,N_7007,N_7168);
or U7518 (N_7518,N_6913,N_6669);
nor U7519 (N_7519,N_6778,N_6958);
and U7520 (N_7520,N_6652,N_6589);
or U7521 (N_7521,N_6980,N_7144);
nand U7522 (N_7522,N_7418,N_6674);
nor U7523 (N_7523,N_7362,N_6287);
and U7524 (N_7524,N_6376,N_6952);
nand U7525 (N_7525,N_6893,N_6939);
xnor U7526 (N_7526,N_6806,N_6455);
xor U7527 (N_7527,N_6167,N_6485);
nand U7528 (N_7528,N_6610,N_6716);
xnor U7529 (N_7529,N_6114,N_7369);
or U7530 (N_7530,N_6498,N_6380);
nor U7531 (N_7531,N_6550,N_6820);
xor U7532 (N_7532,N_6542,N_7200);
nand U7533 (N_7533,N_7318,N_7354);
or U7534 (N_7534,N_7259,N_6122);
or U7535 (N_7535,N_7449,N_6070);
and U7536 (N_7536,N_7299,N_6872);
xor U7537 (N_7537,N_7399,N_6747);
or U7538 (N_7538,N_7070,N_6570);
or U7539 (N_7539,N_6165,N_6769);
nor U7540 (N_7540,N_7032,N_6600);
nand U7541 (N_7541,N_6521,N_7142);
nand U7542 (N_7542,N_6530,N_6572);
or U7543 (N_7543,N_6620,N_7274);
xor U7544 (N_7544,N_6888,N_6304);
nand U7545 (N_7545,N_6605,N_6950);
nand U7546 (N_7546,N_6489,N_6452);
or U7547 (N_7547,N_6212,N_6468);
or U7548 (N_7548,N_6546,N_6343);
nor U7549 (N_7549,N_6189,N_6428);
xor U7550 (N_7550,N_6142,N_7014);
and U7551 (N_7551,N_7066,N_6172);
nand U7552 (N_7552,N_7411,N_6848);
xnor U7553 (N_7553,N_7054,N_6002);
and U7554 (N_7554,N_7455,N_6895);
nand U7555 (N_7555,N_6393,N_7313);
nand U7556 (N_7556,N_7353,N_7151);
or U7557 (N_7557,N_6333,N_7272);
nand U7558 (N_7558,N_6196,N_6007);
nand U7559 (N_7559,N_6891,N_7423);
xnor U7560 (N_7560,N_6135,N_6098);
nand U7561 (N_7561,N_6862,N_6634);
or U7562 (N_7562,N_7232,N_6071);
nand U7563 (N_7563,N_6593,N_7461);
or U7564 (N_7564,N_6603,N_6319);
nor U7565 (N_7565,N_6868,N_7229);
nand U7566 (N_7566,N_6285,N_6749);
and U7567 (N_7567,N_7481,N_6029);
nand U7568 (N_7568,N_6999,N_6037);
xnor U7569 (N_7569,N_6798,N_6646);
or U7570 (N_7570,N_7406,N_6159);
nand U7571 (N_7571,N_6008,N_6714);
xor U7572 (N_7572,N_7492,N_6772);
nor U7573 (N_7573,N_6836,N_7286);
nor U7574 (N_7574,N_7372,N_6161);
nand U7575 (N_7575,N_6713,N_6795);
xor U7576 (N_7576,N_7012,N_6473);
nor U7577 (N_7577,N_7039,N_6458);
nor U7578 (N_7578,N_6712,N_6052);
or U7579 (N_7579,N_6857,N_6157);
nand U7580 (N_7580,N_7121,N_6997);
nor U7581 (N_7581,N_6188,N_7255);
nand U7582 (N_7582,N_7482,N_6575);
xor U7583 (N_7583,N_6225,N_6885);
nor U7584 (N_7584,N_7158,N_6378);
nor U7585 (N_7585,N_6010,N_6179);
xnor U7586 (N_7586,N_7209,N_6654);
or U7587 (N_7587,N_6364,N_7216);
nand U7588 (N_7588,N_6748,N_6075);
and U7589 (N_7589,N_7432,N_6138);
nor U7590 (N_7590,N_7293,N_7021);
and U7591 (N_7591,N_6847,N_6413);
nand U7592 (N_7592,N_6470,N_7495);
and U7593 (N_7593,N_7431,N_7361);
and U7594 (N_7594,N_6301,N_7065);
nor U7595 (N_7595,N_7278,N_7302);
and U7596 (N_7596,N_6127,N_6058);
or U7597 (N_7597,N_6426,N_7005);
nor U7598 (N_7598,N_6249,N_6438);
or U7599 (N_7599,N_7082,N_6076);
and U7600 (N_7600,N_6306,N_7045);
and U7601 (N_7601,N_7227,N_6391);
nand U7602 (N_7602,N_7008,N_7062);
xor U7603 (N_7603,N_6813,N_6594);
xnor U7604 (N_7604,N_6540,N_6811);
xor U7605 (N_7605,N_6174,N_6954);
xnor U7606 (N_7606,N_6527,N_7499);
nand U7607 (N_7607,N_6860,N_6077);
nor U7608 (N_7608,N_6396,N_7112);
and U7609 (N_7609,N_7078,N_6144);
and U7610 (N_7610,N_6124,N_7188);
and U7611 (N_7611,N_6774,N_6839);
nand U7612 (N_7612,N_7447,N_6563);
and U7613 (N_7613,N_6700,N_6584);
nor U7614 (N_7614,N_7000,N_6842);
xnor U7615 (N_7615,N_6126,N_6295);
nand U7616 (N_7616,N_6443,N_6133);
xor U7617 (N_7617,N_6015,N_7316);
and U7618 (N_7618,N_7128,N_6901);
nand U7619 (N_7619,N_6338,N_6100);
nor U7620 (N_7620,N_6957,N_6892);
or U7621 (N_7621,N_6257,N_6513);
nand U7622 (N_7622,N_6744,N_7133);
or U7623 (N_7623,N_7339,N_7389);
nor U7624 (N_7624,N_6291,N_6915);
or U7625 (N_7625,N_6934,N_6099);
nor U7626 (N_7626,N_6476,N_7109);
and U7627 (N_7627,N_7458,N_7407);
and U7628 (N_7628,N_7165,N_6185);
and U7629 (N_7629,N_6723,N_6827);
xnor U7630 (N_7630,N_7081,N_7300);
xor U7631 (N_7631,N_6996,N_6081);
and U7632 (N_7632,N_6880,N_7422);
xor U7633 (N_7633,N_6103,N_7183);
nand U7634 (N_7634,N_6539,N_6327);
or U7635 (N_7635,N_6577,N_6870);
nand U7636 (N_7636,N_7485,N_6178);
and U7637 (N_7637,N_6935,N_7113);
nand U7638 (N_7638,N_7453,N_7341);
or U7639 (N_7639,N_6499,N_7443);
or U7640 (N_7640,N_6959,N_7410);
and U7641 (N_7641,N_6379,N_7413);
and U7642 (N_7642,N_7067,N_7091);
nand U7643 (N_7643,N_6791,N_6298);
nor U7644 (N_7644,N_6139,N_7236);
nand U7645 (N_7645,N_7309,N_7192);
or U7646 (N_7646,N_7421,N_7084);
or U7647 (N_7647,N_6528,N_6556);
and U7648 (N_7648,N_6192,N_6494);
xor U7649 (N_7649,N_6263,N_6788);
nand U7650 (N_7650,N_6583,N_6785);
or U7651 (N_7651,N_6149,N_7307);
and U7652 (N_7652,N_6272,N_6125);
nand U7653 (N_7653,N_6562,N_6102);
nand U7654 (N_7654,N_6048,N_6001);
nand U7655 (N_7655,N_7285,N_6417);
xor U7656 (N_7656,N_6726,N_6328);
nand U7657 (N_7657,N_7171,N_6006);
nand U7658 (N_7658,N_6752,N_7163);
or U7659 (N_7659,N_6305,N_6201);
and U7660 (N_7660,N_6683,N_6260);
or U7661 (N_7661,N_6483,N_6615);
nor U7662 (N_7662,N_6168,N_6464);
nand U7663 (N_7663,N_7497,N_6418);
or U7664 (N_7664,N_6410,N_7017);
and U7665 (N_7665,N_6302,N_6961);
or U7666 (N_7666,N_6089,N_6436);
nand U7667 (N_7667,N_7477,N_6282);
nand U7668 (N_7668,N_6588,N_7325);
or U7669 (N_7669,N_6855,N_6832);
xnor U7670 (N_7670,N_6280,N_6977);
nand U7671 (N_7671,N_7004,N_6023);
and U7672 (N_7672,N_6423,N_7490);
nor U7673 (N_7673,N_6434,N_6936);
nand U7674 (N_7674,N_6815,N_7252);
nor U7675 (N_7675,N_7102,N_6642);
or U7676 (N_7676,N_6786,N_7427);
or U7677 (N_7677,N_7258,N_6554);
or U7678 (N_7678,N_6828,N_6720);
nor U7679 (N_7679,N_6638,N_7018);
xnor U7680 (N_7680,N_6500,N_6307);
or U7681 (N_7681,N_6350,N_6951);
or U7682 (N_7682,N_6881,N_6318);
and U7683 (N_7683,N_7024,N_7228);
nand U7684 (N_7684,N_6869,N_6826);
and U7685 (N_7685,N_6905,N_6976);
nor U7686 (N_7686,N_7474,N_7138);
and U7687 (N_7687,N_6309,N_7404);
xor U7688 (N_7688,N_7238,N_7496);
nor U7689 (N_7689,N_6523,N_6650);
nand U7690 (N_7690,N_6341,N_6852);
and U7691 (N_7691,N_6994,N_6140);
or U7692 (N_7692,N_7349,N_7304);
nand U7693 (N_7693,N_7178,N_7468);
nor U7694 (N_7694,N_7198,N_6814);
and U7695 (N_7695,N_6231,N_6060);
xor U7696 (N_7696,N_6768,N_6299);
xor U7697 (N_7697,N_7058,N_6460);
and U7698 (N_7698,N_6357,N_6315);
and U7699 (N_7699,N_7265,N_7104);
nor U7700 (N_7700,N_7378,N_6345);
xnor U7701 (N_7701,N_6118,N_6766);
nand U7702 (N_7702,N_6419,N_6359);
and U7703 (N_7703,N_6819,N_6587);
and U7704 (N_7704,N_7245,N_6439);
nor U7705 (N_7705,N_7096,N_6342);
and U7706 (N_7706,N_6035,N_6644);
or U7707 (N_7707,N_6833,N_6512);
nor U7708 (N_7708,N_6171,N_7292);
nand U7709 (N_7709,N_7011,N_7074);
nand U7710 (N_7710,N_6783,N_6399);
or U7711 (N_7711,N_6724,N_6290);
nor U7712 (N_7712,N_6850,N_6701);
and U7713 (N_7713,N_7465,N_6676);
nand U7714 (N_7714,N_7260,N_7419);
or U7715 (N_7715,N_6955,N_6496);
xor U7716 (N_7716,N_7189,N_6679);
and U7717 (N_7717,N_7220,N_6243);
or U7718 (N_7718,N_7186,N_6706);
nor U7719 (N_7719,N_6454,N_6368);
nor U7720 (N_7720,N_6900,N_6715);
and U7721 (N_7721,N_6663,N_7281);
nor U7722 (N_7722,N_6289,N_6741);
nor U7723 (N_7723,N_6339,N_6421);
nor U7724 (N_7724,N_6349,N_6404);
nand U7725 (N_7725,N_6520,N_6661);
and U7726 (N_7726,N_6169,N_6607);
xor U7727 (N_7727,N_6742,N_6845);
and U7728 (N_7728,N_6377,N_7315);
xnor U7729 (N_7729,N_6416,N_7264);
or U7730 (N_7730,N_6362,N_7098);
and U7731 (N_7731,N_6264,N_6581);
nor U7732 (N_7732,N_6698,N_6664);
and U7733 (N_7733,N_6031,N_6366);
nor U7734 (N_7734,N_7239,N_6750);
xor U7735 (N_7735,N_6406,N_7367);
or U7736 (N_7736,N_6072,N_7100);
nand U7737 (N_7737,N_6928,N_6728);
and U7738 (N_7738,N_7436,N_6865);
and U7739 (N_7739,N_6623,N_6177);
xor U7740 (N_7740,N_7089,N_7478);
or U7741 (N_7741,N_7208,N_6985);
nor U7742 (N_7742,N_6402,N_7116);
or U7743 (N_7743,N_7033,N_6804);
xor U7744 (N_7744,N_6537,N_6025);
nand U7745 (N_7745,N_6501,N_6256);
and U7746 (N_7746,N_6911,N_6942);
nand U7747 (N_7747,N_6435,N_6034);
and U7748 (N_7748,N_6737,N_7357);
xor U7749 (N_7749,N_7242,N_7322);
nor U7750 (N_7750,N_7359,N_6219);
xor U7751 (N_7751,N_6236,N_6206);
and U7752 (N_7752,N_6606,N_7051);
nand U7753 (N_7753,N_6160,N_7143);
xor U7754 (N_7754,N_6202,N_7350);
or U7755 (N_7755,N_6898,N_7043);
nor U7756 (N_7756,N_6016,N_7251);
or U7757 (N_7757,N_6867,N_7289);
or U7758 (N_7758,N_7087,N_7329);
or U7759 (N_7759,N_6383,N_7486);
and U7760 (N_7760,N_6602,N_6886);
nor U7761 (N_7761,N_7493,N_7444);
nor U7762 (N_7762,N_6381,N_7385);
nand U7763 (N_7763,N_6030,N_6471);
nand U7764 (N_7764,N_6024,N_6265);
nand U7765 (N_7765,N_6566,N_7174);
xor U7766 (N_7766,N_6722,N_7243);
and U7767 (N_7767,N_6227,N_7180);
or U7768 (N_7768,N_6158,N_6175);
or U7769 (N_7769,N_6971,N_6386);
nand U7770 (N_7770,N_6467,N_7141);
nor U7771 (N_7771,N_7092,N_6667);
nand U7772 (N_7772,N_7185,N_6397);
and U7773 (N_7773,N_7464,N_6916);
or U7774 (N_7774,N_6925,N_6281);
xnor U7775 (N_7775,N_6054,N_6555);
xnor U7776 (N_7776,N_6213,N_7129);
nor U7777 (N_7777,N_6738,N_6044);
xnor U7778 (N_7778,N_7319,N_7126);
and U7779 (N_7779,N_6877,N_7379);
and U7780 (N_7780,N_6734,N_6427);
and U7781 (N_7781,N_7470,N_6286);
nand U7782 (N_7782,N_6830,N_7226);
xor U7783 (N_7783,N_7103,N_6259);
and U7784 (N_7784,N_6505,N_6551);
nand U7785 (N_7785,N_7041,N_6414);
or U7786 (N_7786,N_7167,N_6662);
or U7787 (N_7787,N_7190,N_6472);
nor U7788 (N_7788,N_6204,N_6694);
nand U7789 (N_7789,N_7338,N_6388);
xor U7790 (N_7790,N_6109,N_7034);
xor U7791 (N_7791,N_6181,N_6049);
nand U7792 (N_7792,N_7276,N_6210);
nand U7793 (N_7793,N_7006,N_6271);
or U7794 (N_7794,N_6807,N_6776);
xor U7795 (N_7795,N_6011,N_6353);
xnor U7796 (N_7796,N_6046,N_6370);
and U7797 (N_7797,N_6982,N_7037);
or U7798 (N_7798,N_7199,N_6074);
nand U7799 (N_7799,N_6332,N_7042);
nor U7800 (N_7800,N_6340,N_7147);
or U7801 (N_7801,N_7160,N_6875);
xnor U7802 (N_7802,N_6082,N_6808);
and U7803 (N_7803,N_7262,N_6937);
nor U7804 (N_7804,N_7118,N_7273);
xnor U7805 (N_7805,N_6039,N_6214);
or U7806 (N_7806,N_7331,N_7159);
and U7807 (N_7807,N_7237,N_6549);
xor U7808 (N_7808,N_7295,N_7311);
xnor U7809 (N_7809,N_6507,N_6624);
and U7810 (N_7810,N_7127,N_7162);
and U7811 (N_7811,N_7224,N_6689);
nor U7812 (N_7812,N_7010,N_7219);
nand U7813 (N_7813,N_7451,N_7241);
xnor U7814 (N_7814,N_6365,N_6392);
and U7815 (N_7815,N_6797,N_7016);
or U7816 (N_7816,N_6938,N_7297);
xor U7817 (N_7817,N_6735,N_7348);
or U7818 (N_7818,N_7038,N_6009);
xnor U7819 (N_7819,N_6705,N_6252);
nor U7820 (N_7820,N_6107,N_6148);
or U7821 (N_7821,N_6946,N_7181);
or U7822 (N_7822,N_7221,N_6267);
xnor U7823 (N_7823,N_6538,N_7346);
nor U7824 (N_7824,N_6633,N_6800);
nand U7825 (N_7825,N_7120,N_6064);
or U7826 (N_7826,N_7393,N_6045);
nand U7827 (N_7827,N_7107,N_6322);
or U7828 (N_7828,N_7214,N_7454);
nor U7829 (N_7829,N_6482,N_7172);
and U7830 (N_7830,N_6765,N_6484);
or U7831 (N_7831,N_7029,N_6063);
xor U7832 (N_7832,N_6993,N_6730);
nand U7833 (N_7833,N_7435,N_6258);
and U7834 (N_7834,N_7110,N_7207);
and U7835 (N_7835,N_6111,N_6919);
nand U7836 (N_7836,N_7310,N_7111);
xnor U7837 (N_7837,N_6486,N_7291);
and U7838 (N_7838,N_7093,N_7155);
nor U7839 (N_7839,N_6796,N_6991);
or U7840 (N_7840,N_6004,N_6137);
or U7841 (N_7841,N_6425,N_6238);
and U7842 (N_7842,N_6759,N_7173);
or U7843 (N_7843,N_6767,N_6284);
nand U7844 (N_7844,N_6618,N_6974);
nor U7845 (N_7845,N_6805,N_6012);
xnor U7846 (N_7846,N_6586,N_6637);
and U7847 (N_7847,N_6745,N_6757);
and U7848 (N_7848,N_6608,N_6147);
nor U7849 (N_7849,N_7489,N_6824);
nand U7850 (N_7850,N_6415,N_7169);
nand U7851 (N_7851,N_6970,N_7154);
nand U7852 (N_7852,N_6817,N_6628);
and U7853 (N_7853,N_6028,N_7145);
nand U7854 (N_7854,N_6969,N_6346);
and U7855 (N_7855,N_6532,N_6330);
nand U7856 (N_7856,N_6691,N_6690);
nor U7857 (N_7857,N_6385,N_6543);
xor U7858 (N_7858,N_6226,N_6582);
and U7859 (N_7859,N_6917,N_6433);
nor U7860 (N_7860,N_6311,N_7031);
nand U7861 (N_7861,N_6323,N_7363);
and U7862 (N_7862,N_7211,N_7336);
and U7863 (N_7863,N_6896,N_7415);
nor U7864 (N_7864,N_7491,N_6274);
and U7865 (N_7865,N_6510,N_6422);
and U7866 (N_7866,N_7305,N_6444);
nor U7867 (N_7867,N_6312,N_6480);
or U7868 (N_7868,N_7213,N_6923);
nor U7869 (N_7869,N_6442,N_6649);
or U7870 (N_7870,N_6887,N_6141);
or U7871 (N_7871,N_7343,N_6609);
and U7872 (N_7872,N_7275,N_7197);
xnor U7873 (N_7873,N_7480,N_7282);
or U7874 (N_7874,N_6621,N_7382);
nand U7875 (N_7875,N_6941,N_6294);
xnor U7876 (N_7876,N_6062,N_6233);
nor U7877 (N_7877,N_7314,N_6695);
nor U7878 (N_7878,N_6851,N_6277);
nor U7879 (N_7879,N_6711,N_7135);
and U7880 (N_7880,N_6944,N_6087);
nand U7881 (N_7881,N_6186,N_6902);
nor U7882 (N_7882,N_6429,N_6405);
xnor U7883 (N_7883,N_7332,N_6506);
nand U7884 (N_7884,N_7076,N_6758);
nor U7885 (N_7885,N_6057,N_7412);
xor U7886 (N_7886,N_7269,N_6463);
xnor U7887 (N_7887,N_6446,N_6743);
and U7888 (N_7888,N_6519,N_7409);
nor U7889 (N_7889,N_7179,N_6051);
xor U7890 (N_7890,N_6710,N_7117);
xor U7891 (N_7891,N_6619,N_7069);
nand U7892 (N_7892,N_6352,N_6576);
and U7893 (N_7893,N_6574,N_6105);
or U7894 (N_7894,N_6479,N_7487);
and U7895 (N_7895,N_6678,N_6108);
or U7896 (N_7896,N_6516,N_7308);
nor U7897 (N_7897,N_7036,N_6595);
nor U7898 (N_7898,N_6943,N_7333);
nand U7899 (N_7899,N_6123,N_6130);
xnor U7900 (N_7900,N_6360,N_6921);
nor U7901 (N_7901,N_6626,N_6136);
xor U7902 (N_7902,N_7191,N_7115);
and U7903 (N_7903,N_7125,N_6073);
nor U7904 (N_7904,N_6933,N_7360);
or U7905 (N_7905,N_7201,N_6493);
and U7906 (N_7906,N_6358,N_6557);
xor U7907 (N_7907,N_6882,N_7046);
nand U7908 (N_7908,N_6134,N_6922);
and U7909 (N_7909,N_7072,N_6746);
and U7910 (N_7910,N_7187,N_6524);
and U7911 (N_7911,N_6067,N_7099);
nand U7912 (N_7912,N_7457,N_7088);
and U7913 (N_7913,N_6129,N_6545);
or U7914 (N_7914,N_6110,N_7462);
or U7915 (N_7915,N_6569,N_7114);
nor U7916 (N_7916,N_6040,N_6856);
nor U7917 (N_7917,N_6968,N_6431);
and U7918 (N_7918,N_6334,N_6490);
xor U7919 (N_7919,N_6992,N_7023);
xnor U7920 (N_7920,N_7123,N_6146);
nor U7921 (N_7921,N_7250,N_6088);
nor U7922 (N_7922,N_7047,N_6630);
nor U7923 (N_7923,N_7206,N_6270);
xnor U7924 (N_7924,N_7351,N_7079);
nor U7925 (N_7925,N_6599,N_6191);
nor U7926 (N_7926,N_6038,N_6230);
nand U7927 (N_7927,N_7044,N_7164);
or U7928 (N_7928,N_6182,N_6283);
nor U7929 (N_7929,N_6300,N_6199);
and U7930 (N_7930,N_7437,N_6056);
or U7931 (N_7931,N_7347,N_7390);
and U7932 (N_7932,N_6622,N_6837);
nand U7933 (N_7933,N_6979,N_6211);
xor U7934 (N_7934,N_6704,N_7395);
or U7935 (N_7935,N_6190,N_6255);
xnor U7936 (N_7936,N_6841,N_6878);
and U7937 (N_7937,N_6696,N_6531);
xnor U7938 (N_7938,N_6799,N_7002);
or U7939 (N_7939,N_6657,N_7015);
nand U7940 (N_7940,N_6544,N_6818);
or U7941 (N_7941,N_6998,N_7217);
xor U7942 (N_7942,N_7230,N_6879);
or U7943 (N_7943,N_6699,N_6762);
xor U7944 (N_7944,N_7321,N_7365);
nor U7945 (N_7945,N_6825,N_6205);
or U7946 (N_7946,N_6787,N_6027);
or U7947 (N_7947,N_6962,N_7405);
or U7948 (N_7948,N_6497,N_7396);
nand U7949 (N_7949,N_6792,N_6437);
nand U7950 (N_7950,N_6374,N_7153);
nor U7951 (N_7951,N_6627,N_6262);
xor U7952 (N_7952,N_6209,N_6043);
or U7953 (N_7953,N_7080,N_6170);
and U7954 (N_7954,N_6871,N_6080);
or U7955 (N_7955,N_7231,N_6207);
xnor U7956 (N_7956,N_7131,N_6119);
or U7957 (N_7957,N_7450,N_6802);
nor U7958 (N_7958,N_6020,N_6411);
or U7959 (N_7959,N_6843,N_6474);
nand U7960 (N_7960,N_6688,N_6096);
and U7961 (N_7961,N_6708,N_7335);
nor U7962 (N_7962,N_7459,N_6461);
nor U7963 (N_7963,N_6348,N_6535);
nand U7964 (N_7964,N_6789,N_7294);
xor U7965 (N_7965,N_6949,N_6612);
or U7966 (N_7966,N_6821,N_6042);
nor U7967 (N_7967,N_6235,N_6347);
nand U7968 (N_7968,N_7057,N_6719);
nor U7969 (N_7969,N_7440,N_6764);
nor U7970 (N_7970,N_6515,N_6465);
nor U7971 (N_7971,N_7149,N_7466);
or U7972 (N_7972,N_6183,N_7137);
xor U7973 (N_7973,N_7344,N_6369);
nor U7974 (N_7974,N_6061,N_7340);
xor U7975 (N_7975,N_6248,N_6509);
nor U7976 (N_7976,N_7055,N_6973);
xnor U7977 (N_7977,N_7375,N_6487);
nand U7978 (N_7978,N_6671,N_6344);
xnor U7979 (N_7979,N_6166,N_7134);
xor U7980 (N_7980,N_6790,N_7271);
xnor U7981 (N_7981,N_6153,N_6424);
nand U7982 (N_7982,N_6823,N_6351);
nor U7983 (N_7983,N_7234,N_6375);
nand U7984 (N_7984,N_6387,N_7373);
or U7985 (N_7985,N_6246,N_6803);
or U7986 (N_7986,N_6866,N_7071);
or U7987 (N_7987,N_7463,N_6194);
xnor U7988 (N_7988,N_6459,N_6400);
xor U7989 (N_7989,N_6677,N_6251);
nor U7990 (N_7990,N_7330,N_7063);
or U7991 (N_7991,N_6727,N_7064);
nand U7992 (N_7992,N_7139,N_6090);
nand U7993 (N_7993,N_7205,N_6918);
nor U7994 (N_7994,N_7196,N_6503);
or U7995 (N_7995,N_6150,N_6945);
and U7996 (N_7996,N_6559,N_6908);
nand U7997 (N_7997,N_7337,N_6232);
nor U7998 (N_7998,N_7290,N_7193);
or U7999 (N_7999,N_6656,N_6106);
and U8000 (N_8000,N_6590,N_6794);
xnor U8001 (N_8001,N_7323,N_7256);
and U8002 (N_8002,N_6631,N_6611);
or U8003 (N_8003,N_7106,N_6223);
nand U8004 (N_8004,N_6432,N_6511);
nand U8005 (N_8005,N_6093,N_6987);
and U8006 (N_8006,N_6120,N_7030);
or U8007 (N_8007,N_6036,N_6296);
or U8008 (N_8008,N_7267,N_6198);
or U8009 (N_8009,N_7059,N_6930);
nand U8010 (N_8010,N_6965,N_6187);
or U8011 (N_8011,N_6079,N_6250);
xor U8012 (N_8012,N_7218,N_7266);
nand U8013 (N_8013,N_6697,N_7049);
nand U8014 (N_8014,N_7434,N_6143);
xor U8015 (N_8015,N_6065,N_6883);
and U8016 (N_8016,N_7352,N_7381);
and U8017 (N_8017,N_6625,N_6151);
nand U8018 (N_8018,N_6491,N_7225);
nor U8019 (N_8019,N_7268,N_7342);
xnor U8020 (N_8020,N_6017,N_7428);
or U8021 (N_8021,N_6237,N_6534);
nor U8022 (N_8022,N_7140,N_7483);
xor U8023 (N_8023,N_7476,N_6317);
or U8024 (N_8024,N_7377,N_6874);
xnor U8025 (N_8025,N_6163,N_6068);
xor U8026 (N_8026,N_6740,N_6873);
xor U8027 (N_8027,N_6835,N_6326);
nor U8028 (N_8028,N_6220,N_6682);
nand U8029 (N_8029,N_6078,N_7288);
and U8030 (N_8030,N_6293,N_6536);
nor U8031 (N_8031,N_6910,N_6770);
nor U8032 (N_8032,N_6653,N_7416);
and U8033 (N_8033,N_6684,N_7441);
nor U8034 (N_8034,N_6441,N_6273);
or U8035 (N_8035,N_6447,N_6176);
xor U8036 (N_8036,N_6897,N_7371);
nor U8037 (N_8037,N_6324,N_6665);
nand U8038 (N_8038,N_7403,N_6253);
xor U8039 (N_8039,N_6755,N_6859);
nand U8040 (N_8040,N_6316,N_6989);
xnor U8041 (N_8041,N_7166,N_6389);
nand U8042 (N_8042,N_7380,N_6693);
nor U8043 (N_8043,N_7086,N_6526);
and U8044 (N_8044,N_6812,N_6420);
nor U8045 (N_8045,N_7108,N_6801);
xnor U8046 (N_8046,N_7052,N_6005);
or U8047 (N_8047,N_7182,N_6297);
or U8048 (N_8048,N_6967,N_7244);
xnor U8049 (N_8049,N_6239,N_6014);
and U8050 (N_8050,N_6707,N_6658);
nor U8051 (N_8051,N_6585,N_7027);
and U8052 (N_8052,N_6518,N_7345);
nand U8053 (N_8053,N_6552,N_7022);
or U8054 (N_8054,N_6629,N_7094);
xor U8055 (N_8055,N_6477,N_6355);
nand U8056 (N_8056,N_6929,N_6066);
and U8057 (N_8057,N_7400,N_7438);
xor U8058 (N_8058,N_7448,N_6481);
or U8059 (N_8059,N_7467,N_7025);
nand U8060 (N_8060,N_7248,N_6228);
or U8061 (N_8061,N_6966,N_6641);
or U8062 (N_8062,N_7176,N_6449);
xnor U8063 (N_8063,N_6753,N_6909);
or U8064 (N_8064,N_6846,N_6894);
or U8065 (N_8065,N_6844,N_6522);
xnor U8066 (N_8066,N_6112,N_6604);
and U8067 (N_8067,N_6907,N_6221);
nand U8068 (N_8068,N_7001,N_6469);
nor U8069 (N_8069,N_6924,N_7283);
nand U8070 (N_8070,N_6617,N_7287);
or U8071 (N_8071,N_6217,N_6195);
xnor U8072 (N_8072,N_6579,N_7254);
xnor U8073 (N_8073,N_6840,N_7040);
xor U8074 (N_8074,N_6050,N_7083);
xnor U8075 (N_8075,N_7391,N_6155);
nor U8076 (N_8076,N_7473,N_6336);
or U8077 (N_8077,N_7233,N_6725);
nor U8078 (N_8078,N_6240,N_7026);
xnor U8079 (N_8079,N_6097,N_6121);
xnor U8080 (N_8080,N_7296,N_6780);
nand U8081 (N_8081,N_7387,N_7498);
xnor U8082 (N_8082,N_6560,N_6390);
or U8083 (N_8083,N_6279,N_6222);
nand U8084 (N_8084,N_7306,N_6502);
or U8085 (N_8085,N_7355,N_6988);
xor U8086 (N_8086,N_6288,N_6104);
or U8087 (N_8087,N_6960,N_7303);
and U8088 (N_8088,N_7035,N_6229);
xnor U8089 (N_8089,N_6269,N_7152);
xor U8090 (N_8090,N_7073,N_6059);
and U8091 (N_8091,N_6983,N_6645);
or U8092 (N_8092,N_7095,N_6363);
or U8093 (N_8093,N_6261,N_6963);
xor U8094 (N_8094,N_7235,N_6533);
xnor U8095 (N_8095,N_6947,N_6972);
and U8096 (N_8096,N_7013,N_6831);
nand U8097 (N_8097,N_6448,N_6809);
and U8098 (N_8098,N_6180,N_6292);
or U8099 (N_8099,N_6597,N_6592);
nand U8100 (N_8100,N_7388,N_6128);
or U8101 (N_8101,N_7327,N_6331);
nor U8102 (N_8102,N_6659,N_6026);
nor U8103 (N_8103,N_6558,N_6314);
and U8104 (N_8104,N_6525,N_6829);
and U8105 (N_8105,N_7075,N_6244);
xor U8106 (N_8106,N_7090,N_6889);
nand U8107 (N_8107,N_6890,N_6834);
nor U8108 (N_8108,N_6648,N_7488);
xnor U8109 (N_8109,N_6703,N_6117);
and U8110 (N_8110,N_6672,N_6864);
and U8111 (N_8111,N_7446,N_7326);
nand U8112 (N_8112,N_6382,N_7301);
or U8113 (N_8113,N_6018,N_7048);
and U8114 (N_8114,N_6567,N_6218);
or U8115 (N_8115,N_6777,N_6784);
and U8116 (N_8116,N_7170,N_6573);
nor U8117 (N_8117,N_6022,N_7136);
nor U8118 (N_8118,N_6591,N_7430);
xnor U8119 (N_8119,N_6571,N_7279);
nand U8120 (N_8120,N_6660,N_7420);
xor U8121 (N_8121,N_7334,N_6488);
and U8122 (N_8122,N_7368,N_6401);
nor U8123 (N_8123,N_6553,N_7077);
nor U8124 (N_8124,N_7397,N_7061);
or U8125 (N_8125,N_6781,N_6092);
nand U8126 (N_8126,N_6216,N_6884);
nor U8127 (N_8127,N_7469,N_7222);
xor U8128 (N_8128,N_7460,N_6069);
and U8129 (N_8129,N_6561,N_6154);
nor U8130 (N_8130,N_6903,N_6614);
nand U8131 (N_8131,N_6876,N_6113);
or U8132 (N_8132,N_6858,N_7364);
or U8133 (N_8133,N_6601,N_6086);
and U8134 (N_8134,N_6906,N_6320);
nor U8135 (N_8135,N_6732,N_7161);
or U8136 (N_8136,N_6673,N_6647);
and U8137 (N_8137,N_6091,N_7328);
nand U8138 (N_8138,N_6680,N_6635);
and U8139 (N_8139,N_7215,N_7277);
nor U8140 (N_8140,N_6547,N_7204);
nor U8141 (N_8141,N_7085,N_7376);
nor U8142 (N_8142,N_6409,N_6504);
or U8143 (N_8143,N_6793,N_7394);
and U8144 (N_8144,N_6651,N_7425);
nand U8145 (N_8145,N_6203,N_7223);
xor U8146 (N_8146,N_6094,N_6047);
xor U8147 (N_8147,N_6709,N_7003);
nand U8148 (N_8148,N_6084,N_6412);
or U8149 (N_8149,N_7247,N_6729);
and U8150 (N_8150,N_6853,N_6095);
and U8151 (N_8151,N_6013,N_6854);
nand U8152 (N_8152,N_6580,N_6145);
xnor U8153 (N_8153,N_6200,N_7484);
nand U8154 (N_8154,N_6861,N_6751);
nand U8155 (N_8155,N_7249,N_6373);
xor U8156 (N_8156,N_6241,N_7175);
nor U8157 (N_8157,N_6754,N_6278);
or U8158 (N_8158,N_6495,N_6245);
nand U8159 (N_8159,N_6904,N_7132);
xnor U8160 (N_8160,N_6308,N_6517);
nand U8161 (N_8161,N_6643,N_6721);
nand U8162 (N_8162,N_7053,N_7202);
nand U8163 (N_8163,N_6456,N_6367);
nand U8164 (N_8164,N_6492,N_6242);
nand U8165 (N_8165,N_7424,N_6041);
or U8166 (N_8166,N_6986,N_6162);
nand U8167 (N_8167,N_6003,N_7494);
or U8168 (N_8168,N_6760,N_6354);
xor U8169 (N_8169,N_7298,N_7068);
and U8170 (N_8170,N_7383,N_6739);
nand U8171 (N_8171,N_6335,N_6687);
nor U8172 (N_8172,N_7417,N_7146);
xnor U8173 (N_8173,N_6975,N_6337);
nand U8174 (N_8174,N_6940,N_6899);
xor U8175 (N_8175,N_7177,N_6053);
or U8176 (N_8176,N_7122,N_6462);
or U8177 (N_8177,N_6636,N_7284);
nand U8178 (N_8178,N_6932,N_6514);
or U8179 (N_8179,N_7270,N_7401);
nor U8180 (N_8180,N_6686,N_7442);
or U8181 (N_8181,N_6453,N_6164);
nand U8182 (N_8182,N_7257,N_6101);
xor U8183 (N_8183,N_6451,N_7210);
or U8184 (N_8184,N_6640,N_6926);
nor U8185 (N_8185,N_6247,N_7324);
nand U8186 (N_8186,N_6173,N_7479);
and U8187 (N_8187,N_7194,N_6032);
or U8188 (N_8188,N_6193,N_6275);
or U8189 (N_8189,N_7261,N_7439);
nor U8190 (N_8190,N_7246,N_7280);
xnor U8191 (N_8191,N_6445,N_6655);
nand U8192 (N_8192,N_7105,N_7028);
and U8193 (N_8193,N_6234,N_7429);
and U8194 (N_8194,N_7384,N_6156);
and U8195 (N_8195,N_6718,N_6152);
xor U8196 (N_8196,N_6529,N_6849);
and U8197 (N_8197,N_6912,N_6384);
and U8198 (N_8198,N_6000,N_6995);
nand U8199 (N_8199,N_6685,N_6398);
nor U8200 (N_8200,N_6613,N_6325);
xor U8201 (N_8201,N_6356,N_6478);
nor U8202 (N_8202,N_6197,N_7317);
xor U8203 (N_8203,N_7426,N_6668);
nor U8204 (N_8204,N_7212,N_7060);
and U8205 (N_8205,N_6372,N_7374);
nor U8206 (N_8206,N_6395,N_6920);
nand U8207 (N_8207,N_7124,N_7392);
nor U8208 (N_8208,N_6816,N_6681);
and U8209 (N_8209,N_6407,N_7101);
xor U8210 (N_8210,N_7452,N_6598);
or U8211 (N_8211,N_7097,N_6717);
xor U8212 (N_8212,N_7240,N_6931);
nor U8213 (N_8213,N_7456,N_7009);
nand U8214 (N_8214,N_6756,N_6775);
and U8215 (N_8215,N_6773,N_7472);
xnor U8216 (N_8216,N_6822,N_7184);
and U8217 (N_8217,N_6508,N_6268);
or U8218 (N_8218,N_6616,N_7471);
xnor U8219 (N_8219,N_6430,N_6736);
and U8220 (N_8220,N_6394,N_6132);
nand U8221 (N_8221,N_7320,N_6675);
or U8222 (N_8222,N_7358,N_6116);
or U8223 (N_8223,N_7203,N_6019);
and U8224 (N_8224,N_6083,N_6276);
and U8225 (N_8225,N_6578,N_7433);
or U8226 (N_8226,N_6208,N_7148);
and U8227 (N_8227,N_6927,N_7408);
nand U8228 (N_8228,N_6403,N_6771);
xnor U8229 (N_8229,N_7156,N_6632);
nand U8230 (N_8230,N_7263,N_6457);
and U8231 (N_8231,N_7157,N_6948);
or U8232 (N_8232,N_6953,N_6254);
nor U8233 (N_8233,N_6838,N_6702);
xor U8234 (N_8234,N_6085,N_6733);
or U8235 (N_8235,N_6329,N_6440);
xor U8236 (N_8236,N_7366,N_6371);
and U8237 (N_8237,N_7050,N_7356);
nand U8238 (N_8238,N_6055,N_6670);
nor U8239 (N_8239,N_6914,N_7370);
and U8240 (N_8240,N_7402,N_6475);
nand U8241 (N_8241,N_6639,N_6184);
xnor U8242 (N_8242,N_6541,N_6215);
xnor U8243 (N_8243,N_7398,N_6466);
or U8244 (N_8244,N_6548,N_6596);
and U8245 (N_8245,N_7119,N_6978);
xor U8246 (N_8246,N_6956,N_6666);
or U8247 (N_8247,N_6321,N_6731);
or U8248 (N_8248,N_6779,N_7475);
or U8249 (N_8249,N_6450,N_6564);
nor U8250 (N_8250,N_7354,N_6003);
or U8251 (N_8251,N_6868,N_7362);
nand U8252 (N_8252,N_7133,N_7223);
nor U8253 (N_8253,N_6430,N_7216);
and U8254 (N_8254,N_7460,N_6870);
and U8255 (N_8255,N_6343,N_6665);
xnor U8256 (N_8256,N_6119,N_7303);
nand U8257 (N_8257,N_6173,N_7298);
nor U8258 (N_8258,N_6198,N_7208);
or U8259 (N_8259,N_6560,N_6796);
nand U8260 (N_8260,N_7362,N_6006);
nor U8261 (N_8261,N_6727,N_6898);
and U8262 (N_8262,N_6321,N_7200);
nand U8263 (N_8263,N_7381,N_7407);
and U8264 (N_8264,N_6856,N_6800);
nor U8265 (N_8265,N_6683,N_7258);
nand U8266 (N_8266,N_6665,N_6131);
xnor U8267 (N_8267,N_6939,N_6323);
and U8268 (N_8268,N_6767,N_6135);
nand U8269 (N_8269,N_6930,N_7257);
and U8270 (N_8270,N_6953,N_7202);
xor U8271 (N_8271,N_7080,N_6612);
nor U8272 (N_8272,N_7155,N_6667);
or U8273 (N_8273,N_6767,N_6777);
and U8274 (N_8274,N_7325,N_7050);
xor U8275 (N_8275,N_7104,N_7307);
or U8276 (N_8276,N_7455,N_7397);
and U8277 (N_8277,N_6006,N_6982);
or U8278 (N_8278,N_6499,N_6773);
xor U8279 (N_8279,N_7412,N_6972);
nor U8280 (N_8280,N_6887,N_6286);
and U8281 (N_8281,N_7369,N_7481);
and U8282 (N_8282,N_6989,N_7193);
and U8283 (N_8283,N_6882,N_6005);
or U8284 (N_8284,N_6679,N_6654);
and U8285 (N_8285,N_7394,N_7471);
or U8286 (N_8286,N_6404,N_7115);
nand U8287 (N_8287,N_7250,N_6854);
xor U8288 (N_8288,N_6837,N_7251);
nand U8289 (N_8289,N_7177,N_6017);
xor U8290 (N_8290,N_6563,N_6247);
xnor U8291 (N_8291,N_7303,N_6489);
xor U8292 (N_8292,N_7440,N_6142);
nor U8293 (N_8293,N_6236,N_7392);
nand U8294 (N_8294,N_7021,N_7038);
nor U8295 (N_8295,N_7384,N_7460);
xor U8296 (N_8296,N_6606,N_6307);
nor U8297 (N_8297,N_6995,N_6246);
nor U8298 (N_8298,N_7292,N_6392);
and U8299 (N_8299,N_7273,N_7153);
nor U8300 (N_8300,N_6534,N_7441);
xor U8301 (N_8301,N_6197,N_6924);
or U8302 (N_8302,N_7150,N_6496);
or U8303 (N_8303,N_6717,N_6840);
or U8304 (N_8304,N_7210,N_6935);
xnor U8305 (N_8305,N_6912,N_7119);
and U8306 (N_8306,N_6426,N_6545);
xnor U8307 (N_8307,N_6762,N_6248);
xnor U8308 (N_8308,N_7017,N_6699);
or U8309 (N_8309,N_7230,N_6463);
xnor U8310 (N_8310,N_7330,N_6677);
and U8311 (N_8311,N_7396,N_6827);
xnor U8312 (N_8312,N_7427,N_7238);
nor U8313 (N_8313,N_7144,N_7372);
and U8314 (N_8314,N_6884,N_6876);
nand U8315 (N_8315,N_7304,N_7164);
nor U8316 (N_8316,N_6176,N_7277);
or U8317 (N_8317,N_6604,N_7174);
nand U8318 (N_8318,N_7277,N_6867);
and U8319 (N_8319,N_7315,N_7350);
and U8320 (N_8320,N_6352,N_6215);
nor U8321 (N_8321,N_6778,N_6273);
nor U8322 (N_8322,N_6999,N_6879);
and U8323 (N_8323,N_6144,N_7320);
nand U8324 (N_8324,N_6202,N_6615);
and U8325 (N_8325,N_6810,N_6263);
xor U8326 (N_8326,N_7259,N_6163);
or U8327 (N_8327,N_6000,N_6760);
nor U8328 (N_8328,N_6309,N_6723);
nor U8329 (N_8329,N_6390,N_7316);
or U8330 (N_8330,N_6936,N_6448);
nand U8331 (N_8331,N_7340,N_7382);
and U8332 (N_8332,N_6630,N_6314);
xor U8333 (N_8333,N_6785,N_6348);
nor U8334 (N_8334,N_6461,N_6080);
xnor U8335 (N_8335,N_6534,N_7249);
and U8336 (N_8336,N_6182,N_7178);
or U8337 (N_8337,N_7466,N_6816);
xor U8338 (N_8338,N_6567,N_7464);
and U8339 (N_8339,N_6034,N_7188);
xor U8340 (N_8340,N_6244,N_6632);
nor U8341 (N_8341,N_7235,N_6864);
nor U8342 (N_8342,N_6806,N_6454);
nor U8343 (N_8343,N_6412,N_6900);
or U8344 (N_8344,N_6998,N_6569);
nor U8345 (N_8345,N_6247,N_6062);
and U8346 (N_8346,N_6463,N_7087);
nor U8347 (N_8347,N_7048,N_6160);
nand U8348 (N_8348,N_7263,N_6018);
and U8349 (N_8349,N_6689,N_6315);
xor U8350 (N_8350,N_6622,N_6351);
nand U8351 (N_8351,N_6261,N_7125);
nor U8352 (N_8352,N_6179,N_6015);
or U8353 (N_8353,N_7042,N_7325);
and U8354 (N_8354,N_6470,N_6233);
xor U8355 (N_8355,N_7387,N_6311);
and U8356 (N_8356,N_7392,N_6609);
and U8357 (N_8357,N_7177,N_7252);
xor U8358 (N_8358,N_6941,N_7200);
and U8359 (N_8359,N_6486,N_7207);
xnor U8360 (N_8360,N_6250,N_6106);
and U8361 (N_8361,N_7164,N_7157);
xor U8362 (N_8362,N_6001,N_7082);
nor U8363 (N_8363,N_7204,N_7493);
or U8364 (N_8364,N_7248,N_6857);
xor U8365 (N_8365,N_6466,N_6899);
and U8366 (N_8366,N_6344,N_6209);
xor U8367 (N_8367,N_6151,N_6142);
nand U8368 (N_8368,N_6847,N_6512);
or U8369 (N_8369,N_6374,N_6110);
xnor U8370 (N_8370,N_7158,N_6697);
xor U8371 (N_8371,N_6191,N_6817);
nor U8372 (N_8372,N_6509,N_7174);
or U8373 (N_8373,N_7324,N_6545);
xnor U8374 (N_8374,N_6649,N_7285);
or U8375 (N_8375,N_6588,N_6324);
nor U8376 (N_8376,N_6618,N_6713);
nand U8377 (N_8377,N_6514,N_6916);
and U8378 (N_8378,N_6381,N_7349);
and U8379 (N_8379,N_6997,N_6436);
and U8380 (N_8380,N_6144,N_7000);
nand U8381 (N_8381,N_7420,N_7345);
and U8382 (N_8382,N_6494,N_6880);
xor U8383 (N_8383,N_6187,N_6133);
nand U8384 (N_8384,N_6005,N_6645);
xor U8385 (N_8385,N_6001,N_6316);
or U8386 (N_8386,N_7122,N_6560);
or U8387 (N_8387,N_7455,N_6620);
xor U8388 (N_8388,N_6983,N_6218);
or U8389 (N_8389,N_6679,N_7442);
xor U8390 (N_8390,N_6663,N_6104);
and U8391 (N_8391,N_6483,N_6787);
nor U8392 (N_8392,N_6489,N_6673);
and U8393 (N_8393,N_6104,N_7186);
nor U8394 (N_8394,N_7188,N_6776);
xnor U8395 (N_8395,N_6409,N_6592);
and U8396 (N_8396,N_6432,N_7298);
and U8397 (N_8397,N_7042,N_6859);
nand U8398 (N_8398,N_6147,N_6328);
or U8399 (N_8399,N_6604,N_6751);
xor U8400 (N_8400,N_6857,N_6990);
and U8401 (N_8401,N_6782,N_6525);
xnor U8402 (N_8402,N_7339,N_6841);
and U8403 (N_8403,N_6486,N_7228);
or U8404 (N_8404,N_7097,N_7022);
or U8405 (N_8405,N_6755,N_6198);
xor U8406 (N_8406,N_6477,N_6016);
and U8407 (N_8407,N_7493,N_7398);
xor U8408 (N_8408,N_6445,N_6159);
nor U8409 (N_8409,N_6174,N_7135);
xnor U8410 (N_8410,N_6756,N_6154);
xor U8411 (N_8411,N_6347,N_6591);
or U8412 (N_8412,N_6859,N_7172);
and U8413 (N_8413,N_7064,N_6115);
xnor U8414 (N_8414,N_6967,N_6075);
xnor U8415 (N_8415,N_7379,N_6088);
xor U8416 (N_8416,N_6354,N_6060);
nand U8417 (N_8417,N_7384,N_6194);
xor U8418 (N_8418,N_6149,N_6094);
nand U8419 (N_8419,N_7327,N_6535);
xnor U8420 (N_8420,N_6598,N_6098);
or U8421 (N_8421,N_6073,N_7263);
nor U8422 (N_8422,N_7177,N_6830);
xor U8423 (N_8423,N_7070,N_6676);
xnor U8424 (N_8424,N_7019,N_6434);
nor U8425 (N_8425,N_6087,N_6297);
and U8426 (N_8426,N_7316,N_6076);
and U8427 (N_8427,N_6289,N_6111);
and U8428 (N_8428,N_7353,N_6490);
xor U8429 (N_8429,N_6463,N_6642);
and U8430 (N_8430,N_7097,N_6014);
xor U8431 (N_8431,N_7259,N_6453);
or U8432 (N_8432,N_6919,N_7312);
and U8433 (N_8433,N_6790,N_6571);
and U8434 (N_8434,N_6352,N_6324);
xnor U8435 (N_8435,N_6713,N_7314);
and U8436 (N_8436,N_7301,N_6490);
xnor U8437 (N_8437,N_6031,N_6050);
or U8438 (N_8438,N_6025,N_6630);
xnor U8439 (N_8439,N_6934,N_7431);
xor U8440 (N_8440,N_7462,N_6274);
nor U8441 (N_8441,N_6817,N_6205);
or U8442 (N_8442,N_6344,N_7215);
or U8443 (N_8443,N_6663,N_6053);
xnor U8444 (N_8444,N_7397,N_7255);
nand U8445 (N_8445,N_6319,N_7402);
and U8446 (N_8446,N_6784,N_7056);
nand U8447 (N_8447,N_6319,N_7403);
nand U8448 (N_8448,N_6368,N_7090);
nor U8449 (N_8449,N_6532,N_6239);
or U8450 (N_8450,N_6930,N_6110);
nand U8451 (N_8451,N_7040,N_6373);
or U8452 (N_8452,N_6618,N_7222);
or U8453 (N_8453,N_7494,N_6883);
or U8454 (N_8454,N_6431,N_6209);
nand U8455 (N_8455,N_7302,N_6529);
and U8456 (N_8456,N_6932,N_6962);
and U8457 (N_8457,N_7292,N_6274);
nand U8458 (N_8458,N_6240,N_6232);
xor U8459 (N_8459,N_6114,N_7265);
and U8460 (N_8460,N_6141,N_6784);
xor U8461 (N_8461,N_6182,N_6052);
xor U8462 (N_8462,N_6046,N_7464);
nand U8463 (N_8463,N_6025,N_6265);
and U8464 (N_8464,N_6453,N_7364);
nand U8465 (N_8465,N_7102,N_6457);
nor U8466 (N_8466,N_6928,N_6573);
or U8467 (N_8467,N_7479,N_7482);
xnor U8468 (N_8468,N_6779,N_6064);
xor U8469 (N_8469,N_6686,N_7184);
or U8470 (N_8470,N_6697,N_6451);
or U8471 (N_8471,N_7151,N_6472);
nor U8472 (N_8472,N_6307,N_6031);
and U8473 (N_8473,N_6517,N_6838);
or U8474 (N_8474,N_6403,N_6752);
and U8475 (N_8475,N_7345,N_6291);
nand U8476 (N_8476,N_7135,N_6637);
nor U8477 (N_8477,N_6802,N_6054);
and U8478 (N_8478,N_7112,N_6039);
or U8479 (N_8479,N_6669,N_6318);
or U8480 (N_8480,N_7067,N_6024);
and U8481 (N_8481,N_6917,N_6887);
and U8482 (N_8482,N_6444,N_7084);
and U8483 (N_8483,N_6049,N_6603);
xor U8484 (N_8484,N_7014,N_6226);
or U8485 (N_8485,N_6268,N_7241);
nand U8486 (N_8486,N_7104,N_7325);
or U8487 (N_8487,N_6866,N_6146);
nand U8488 (N_8488,N_7015,N_7100);
and U8489 (N_8489,N_6678,N_6062);
and U8490 (N_8490,N_7216,N_6577);
or U8491 (N_8491,N_6783,N_6536);
and U8492 (N_8492,N_6642,N_6153);
nand U8493 (N_8493,N_7026,N_7046);
nand U8494 (N_8494,N_6642,N_7432);
xor U8495 (N_8495,N_6069,N_6887);
nand U8496 (N_8496,N_6461,N_7447);
or U8497 (N_8497,N_6064,N_6462);
xnor U8498 (N_8498,N_6158,N_6068);
xnor U8499 (N_8499,N_7297,N_7222);
nand U8500 (N_8500,N_7122,N_7118);
nor U8501 (N_8501,N_6252,N_6883);
xor U8502 (N_8502,N_6839,N_6773);
nor U8503 (N_8503,N_6568,N_6685);
xnor U8504 (N_8504,N_7191,N_6660);
and U8505 (N_8505,N_6064,N_6084);
xor U8506 (N_8506,N_7209,N_6203);
nand U8507 (N_8507,N_7204,N_7378);
nand U8508 (N_8508,N_6947,N_6057);
or U8509 (N_8509,N_6820,N_6191);
nand U8510 (N_8510,N_6338,N_7349);
or U8511 (N_8511,N_6441,N_6005);
nand U8512 (N_8512,N_6549,N_6313);
or U8513 (N_8513,N_6845,N_6186);
or U8514 (N_8514,N_6094,N_6266);
xor U8515 (N_8515,N_6807,N_7016);
and U8516 (N_8516,N_6891,N_6276);
or U8517 (N_8517,N_7401,N_7156);
or U8518 (N_8518,N_6425,N_6536);
xnor U8519 (N_8519,N_6530,N_7204);
nor U8520 (N_8520,N_6881,N_7049);
or U8521 (N_8521,N_6115,N_6916);
xor U8522 (N_8522,N_6733,N_6908);
xor U8523 (N_8523,N_6561,N_6790);
nand U8524 (N_8524,N_6147,N_7381);
or U8525 (N_8525,N_7155,N_7090);
and U8526 (N_8526,N_6963,N_6094);
xor U8527 (N_8527,N_7079,N_6661);
or U8528 (N_8528,N_7440,N_6270);
nor U8529 (N_8529,N_6759,N_7248);
or U8530 (N_8530,N_7127,N_6581);
xor U8531 (N_8531,N_7213,N_6258);
xnor U8532 (N_8532,N_7390,N_6718);
and U8533 (N_8533,N_7422,N_6598);
nand U8534 (N_8534,N_6564,N_6313);
and U8535 (N_8535,N_6441,N_6740);
xnor U8536 (N_8536,N_7011,N_6308);
and U8537 (N_8537,N_6383,N_6224);
nand U8538 (N_8538,N_7269,N_7434);
nor U8539 (N_8539,N_7161,N_6452);
nand U8540 (N_8540,N_6027,N_7030);
or U8541 (N_8541,N_6572,N_6494);
nor U8542 (N_8542,N_6486,N_7038);
or U8543 (N_8543,N_6404,N_6130);
nand U8544 (N_8544,N_7247,N_7081);
xor U8545 (N_8545,N_6224,N_6876);
nor U8546 (N_8546,N_6503,N_6985);
nand U8547 (N_8547,N_6990,N_6439);
nor U8548 (N_8548,N_6795,N_6937);
or U8549 (N_8549,N_6469,N_6018);
and U8550 (N_8550,N_6553,N_6219);
and U8551 (N_8551,N_6258,N_6169);
nor U8552 (N_8552,N_6376,N_6193);
and U8553 (N_8553,N_7431,N_7176);
or U8554 (N_8554,N_6391,N_6130);
nand U8555 (N_8555,N_6067,N_6887);
or U8556 (N_8556,N_6707,N_6788);
xnor U8557 (N_8557,N_6631,N_6061);
xor U8558 (N_8558,N_6473,N_6811);
nor U8559 (N_8559,N_6064,N_6866);
xnor U8560 (N_8560,N_6319,N_6807);
or U8561 (N_8561,N_6542,N_6079);
or U8562 (N_8562,N_6829,N_6950);
nor U8563 (N_8563,N_6718,N_7440);
nor U8564 (N_8564,N_6016,N_6675);
or U8565 (N_8565,N_7304,N_7268);
nand U8566 (N_8566,N_6752,N_7129);
xor U8567 (N_8567,N_6784,N_6026);
xnor U8568 (N_8568,N_6333,N_6410);
or U8569 (N_8569,N_6199,N_6605);
nand U8570 (N_8570,N_6906,N_6433);
nor U8571 (N_8571,N_6109,N_6547);
nand U8572 (N_8572,N_7412,N_6519);
or U8573 (N_8573,N_7356,N_6895);
nand U8574 (N_8574,N_6228,N_6900);
xor U8575 (N_8575,N_6085,N_6130);
or U8576 (N_8576,N_7386,N_6919);
and U8577 (N_8577,N_7164,N_7308);
nand U8578 (N_8578,N_6176,N_6589);
nor U8579 (N_8579,N_7497,N_6755);
nor U8580 (N_8580,N_7107,N_7389);
nand U8581 (N_8581,N_7126,N_6831);
xnor U8582 (N_8582,N_6699,N_6885);
and U8583 (N_8583,N_6481,N_7053);
nor U8584 (N_8584,N_6260,N_6315);
nand U8585 (N_8585,N_6124,N_6902);
and U8586 (N_8586,N_7068,N_7324);
nand U8587 (N_8587,N_6379,N_7134);
and U8588 (N_8588,N_6819,N_7190);
or U8589 (N_8589,N_6799,N_6573);
and U8590 (N_8590,N_7067,N_6901);
nor U8591 (N_8591,N_6736,N_6954);
nor U8592 (N_8592,N_7468,N_7262);
nand U8593 (N_8593,N_6952,N_6792);
nand U8594 (N_8594,N_6478,N_6712);
nor U8595 (N_8595,N_6048,N_6019);
xnor U8596 (N_8596,N_6227,N_6521);
or U8597 (N_8597,N_6457,N_6012);
and U8598 (N_8598,N_7328,N_7237);
and U8599 (N_8599,N_6174,N_7278);
and U8600 (N_8600,N_6516,N_7300);
nand U8601 (N_8601,N_6842,N_7238);
nor U8602 (N_8602,N_6567,N_6059);
xor U8603 (N_8603,N_7291,N_6087);
nand U8604 (N_8604,N_6689,N_6324);
and U8605 (N_8605,N_6025,N_6646);
or U8606 (N_8606,N_6862,N_6131);
nand U8607 (N_8607,N_7494,N_7430);
xnor U8608 (N_8608,N_7380,N_6699);
nor U8609 (N_8609,N_7489,N_6017);
and U8610 (N_8610,N_6715,N_6234);
nor U8611 (N_8611,N_6062,N_6736);
and U8612 (N_8612,N_6409,N_6727);
nor U8613 (N_8613,N_6079,N_6047);
nand U8614 (N_8614,N_6964,N_6385);
and U8615 (N_8615,N_6581,N_7463);
nand U8616 (N_8616,N_6389,N_6553);
nor U8617 (N_8617,N_7114,N_6738);
nand U8618 (N_8618,N_7072,N_7404);
nand U8619 (N_8619,N_6743,N_6505);
or U8620 (N_8620,N_6790,N_6249);
and U8621 (N_8621,N_6921,N_7127);
xnor U8622 (N_8622,N_6227,N_7010);
nand U8623 (N_8623,N_7301,N_6225);
xnor U8624 (N_8624,N_6700,N_6392);
nor U8625 (N_8625,N_6148,N_7203);
nor U8626 (N_8626,N_6176,N_6542);
nand U8627 (N_8627,N_6346,N_7179);
xnor U8628 (N_8628,N_6810,N_6533);
nand U8629 (N_8629,N_6511,N_7147);
nor U8630 (N_8630,N_6458,N_6171);
xor U8631 (N_8631,N_6977,N_7292);
and U8632 (N_8632,N_7471,N_6707);
nor U8633 (N_8633,N_6993,N_6488);
or U8634 (N_8634,N_6179,N_6671);
or U8635 (N_8635,N_7419,N_7192);
xnor U8636 (N_8636,N_6813,N_7079);
or U8637 (N_8637,N_6540,N_6589);
xnor U8638 (N_8638,N_7359,N_7091);
and U8639 (N_8639,N_6156,N_6485);
xnor U8640 (N_8640,N_7431,N_6430);
and U8641 (N_8641,N_6671,N_6814);
or U8642 (N_8642,N_6556,N_6146);
nor U8643 (N_8643,N_7332,N_6451);
nor U8644 (N_8644,N_6490,N_7383);
or U8645 (N_8645,N_6566,N_7112);
xnor U8646 (N_8646,N_6576,N_6424);
or U8647 (N_8647,N_6639,N_6849);
xor U8648 (N_8648,N_6522,N_6956);
xor U8649 (N_8649,N_7447,N_7374);
nor U8650 (N_8650,N_6812,N_6919);
nand U8651 (N_8651,N_6336,N_6605);
xor U8652 (N_8652,N_6710,N_6182);
nor U8653 (N_8653,N_6609,N_6455);
and U8654 (N_8654,N_6356,N_6216);
nand U8655 (N_8655,N_6988,N_7103);
and U8656 (N_8656,N_6912,N_6918);
nor U8657 (N_8657,N_7483,N_6646);
nand U8658 (N_8658,N_7485,N_7420);
or U8659 (N_8659,N_7471,N_6755);
nand U8660 (N_8660,N_6885,N_7249);
nor U8661 (N_8661,N_6782,N_6156);
nor U8662 (N_8662,N_6268,N_6088);
or U8663 (N_8663,N_6165,N_6502);
or U8664 (N_8664,N_6358,N_7025);
and U8665 (N_8665,N_6798,N_6969);
or U8666 (N_8666,N_7483,N_6565);
nor U8667 (N_8667,N_6493,N_6849);
xnor U8668 (N_8668,N_6880,N_6814);
nor U8669 (N_8669,N_6239,N_6517);
xnor U8670 (N_8670,N_7011,N_6520);
xnor U8671 (N_8671,N_6191,N_7221);
or U8672 (N_8672,N_6398,N_7108);
nor U8673 (N_8673,N_7063,N_6260);
and U8674 (N_8674,N_6708,N_6031);
nor U8675 (N_8675,N_6422,N_6904);
or U8676 (N_8676,N_6221,N_6796);
or U8677 (N_8677,N_7153,N_7027);
or U8678 (N_8678,N_6535,N_7131);
or U8679 (N_8679,N_6957,N_7188);
xnor U8680 (N_8680,N_6799,N_6849);
or U8681 (N_8681,N_6172,N_6535);
and U8682 (N_8682,N_7471,N_6188);
xnor U8683 (N_8683,N_6038,N_6010);
xnor U8684 (N_8684,N_6665,N_6770);
and U8685 (N_8685,N_6698,N_6253);
xnor U8686 (N_8686,N_6244,N_7009);
and U8687 (N_8687,N_7346,N_6060);
nand U8688 (N_8688,N_7311,N_6976);
and U8689 (N_8689,N_7282,N_6605);
nand U8690 (N_8690,N_7027,N_6135);
nand U8691 (N_8691,N_6728,N_6800);
or U8692 (N_8692,N_6003,N_6870);
nor U8693 (N_8693,N_7188,N_6282);
or U8694 (N_8694,N_6311,N_6290);
or U8695 (N_8695,N_6177,N_7065);
xor U8696 (N_8696,N_7462,N_6329);
xnor U8697 (N_8697,N_6753,N_6762);
nor U8698 (N_8698,N_6056,N_6561);
or U8699 (N_8699,N_7436,N_7201);
xnor U8700 (N_8700,N_7009,N_7303);
nand U8701 (N_8701,N_6823,N_6931);
nor U8702 (N_8702,N_6867,N_7177);
nor U8703 (N_8703,N_6918,N_6972);
or U8704 (N_8704,N_7234,N_6128);
nand U8705 (N_8705,N_6009,N_6878);
nor U8706 (N_8706,N_7243,N_7333);
nor U8707 (N_8707,N_7035,N_6666);
and U8708 (N_8708,N_6568,N_6197);
nand U8709 (N_8709,N_7414,N_6740);
nor U8710 (N_8710,N_6295,N_7321);
nor U8711 (N_8711,N_6381,N_6164);
xnor U8712 (N_8712,N_6766,N_6817);
or U8713 (N_8713,N_6356,N_6652);
nor U8714 (N_8714,N_6346,N_6187);
or U8715 (N_8715,N_7190,N_6326);
nor U8716 (N_8716,N_7189,N_6554);
xor U8717 (N_8717,N_6019,N_7233);
nand U8718 (N_8718,N_6914,N_6907);
and U8719 (N_8719,N_6788,N_6162);
nand U8720 (N_8720,N_6488,N_7071);
xor U8721 (N_8721,N_6157,N_6436);
nor U8722 (N_8722,N_6349,N_6570);
xor U8723 (N_8723,N_7350,N_7462);
and U8724 (N_8724,N_7297,N_6092);
nor U8725 (N_8725,N_6725,N_6336);
or U8726 (N_8726,N_6603,N_7431);
nand U8727 (N_8727,N_6449,N_7085);
nand U8728 (N_8728,N_7144,N_6926);
and U8729 (N_8729,N_7261,N_6273);
or U8730 (N_8730,N_6452,N_6804);
xnor U8731 (N_8731,N_6536,N_7483);
or U8732 (N_8732,N_7355,N_6228);
nand U8733 (N_8733,N_7274,N_6820);
xnor U8734 (N_8734,N_7058,N_7244);
nor U8735 (N_8735,N_6511,N_6323);
and U8736 (N_8736,N_7438,N_6923);
and U8737 (N_8737,N_7299,N_6827);
and U8738 (N_8738,N_7468,N_6103);
nand U8739 (N_8739,N_6239,N_6298);
nor U8740 (N_8740,N_6534,N_6011);
nand U8741 (N_8741,N_6809,N_6691);
nand U8742 (N_8742,N_6145,N_7413);
xor U8743 (N_8743,N_7395,N_6137);
xnor U8744 (N_8744,N_7047,N_6975);
xor U8745 (N_8745,N_6800,N_6627);
xor U8746 (N_8746,N_7222,N_6987);
or U8747 (N_8747,N_6658,N_6100);
nor U8748 (N_8748,N_6369,N_6808);
nand U8749 (N_8749,N_7104,N_6337);
nand U8750 (N_8750,N_6266,N_7443);
or U8751 (N_8751,N_6935,N_6007);
and U8752 (N_8752,N_7224,N_6816);
and U8753 (N_8753,N_6926,N_7310);
and U8754 (N_8754,N_6762,N_6133);
and U8755 (N_8755,N_7200,N_6857);
nand U8756 (N_8756,N_6115,N_6687);
xor U8757 (N_8757,N_6358,N_7151);
nand U8758 (N_8758,N_6951,N_6561);
nand U8759 (N_8759,N_6192,N_6638);
nand U8760 (N_8760,N_6504,N_7088);
and U8761 (N_8761,N_6343,N_6812);
nor U8762 (N_8762,N_6506,N_7067);
nor U8763 (N_8763,N_6907,N_6085);
nor U8764 (N_8764,N_6600,N_6742);
and U8765 (N_8765,N_6109,N_6207);
nand U8766 (N_8766,N_6843,N_6750);
nand U8767 (N_8767,N_7434,N_6176);
or U8768 (N_8768,N_6650,N_6600);
and U8769 (N_8769,N_6148,N_6340);
nor U8770 (N_8770,N_7087,N_6168);
or U8771 (N_8771,N_6682,N_7385);
or U8772 (N_8772,N_6747,N_6469);
xor U8773 (N_8773,N_6624,N_6837);
xor U8774 (N_8774,N_6342,N_7302);
or U8775 (N_8775,N_6465,N_7063);
nand U8776 (N_8776,N_7485,N_6501);
or U8777 (N_8777,N_7048,N_6680);
or U8778 (N_8778,N_6010,N_6558);
xor U8779 (N_8779,N_7407,N_6875);
nor U8780 (N_8780,N_6629,N_7174);
or U8781 (N_8781,N_6321,N_7424);
or U8782 (N_8782,N_6545,N_7104);
nand U8783 (N_8783,N_7125,N_6836);
nand U8784 (N_8784,N_6491,N_6675);
or U8785 (N_8785,N_7041,N_6939);
nand U8786 (N_8786,N_6513,N_7331);
nor U8787 (N_8787,N_6829,N_7308);
and U8788 (N_8788,N_7334,N_6388);
nor U8789 (N_8789,N_7164,N_7199);
nand U8790 (N_8790,N_7174,N_6582);
xor U8791 (N_8791,N_6522,N_6231);
nand U8792 (N_8792,N_6132,N_6135);
nand U8793 (N_8793,N_6198,N_6981);
nor U8794 (N_8794,N_7011,N_6865);
nand U8795 (N_8795,N_6070,N_6212);
or U8796 (N_8796,N_6617,N_7306);
nand U8797 (N_8797,N_7119,N_6894);
and U8798 (N_8798,N_7194,N_7331);
or U8799 (N_8799,N_7235,N_7465);
nand U8800 (N_8800,N_7279,N_6287);
or U8801 (N_8801,N_6105,N_7486);
and U8802 (N_8802,N_6059,N_7101);
and U8803 (N_8803,N_6943,N_6355);
nor U8804 (N_8804,N_7234,N_7043);
and U8805 (N_8805,N_7060,N_7010);
or U8806 (N_8806,N_6885,N_6264);
xnor U8807 (N_8807,N_6902,N_7443);
nand U8808 (N_8808,N_6818,N_6951);
xnor U8809 (N_8809,N_6398,N_6360);
and U8810 (N_8810,N_7378,N_6976);
or U8811 (N_8811,N_6614,N_6654);
and U8812 (N_8812,N_7458,N_6443);
xor U8813 (N_8813,N_7462,N_6120);
xnor U8814 (N_8814,N_6386,N_7125);
nand U8815 (N_8815,N_6842,N_6368);
or U8816 (N_8816,N_7430,N_6424);
xor U8817 (N_8817,N_6637,N_6107);
or U8818 (N_8818,N_6887,N_6993);
nand U8819 (N_8819,N_6531,N_6039);
nand U8820 (N_8820,N_6136,N_7207);
xnor U8821 (N_8821,N_6197,N_7172);
and U8822 (N_8822,N_6327,N_7353);
or U8823 (N_8823,N_7274,N_7326);
or U8824 (N_8824,N_6426,N_6596);
xnor U8825 (N_8825,N_6361,N_7152);
and U8826 (N_8826,N_7134,N_6262);
or U8827 (N_8827,N_6302,N_6793);
and U8828 (N_8828,N_6674,N_6711);
nor U8829 (N_8829,N_6313,N_6997);
nand U8830 (N_8830,N_7197,N_6759);
nor U8831 (N_8831,N_6483,N_6258);
and U8832 (N_8832,N_6490,N_6707);
nor U8833 (N_8833,N_7334,N_6851);
xor U8834 (N_8834,N_6613,N_6450);
xor U8835 (N_8835,N_7442,N_6909);
nor U8836 (N_8836,N_7360,N_6229);
or U8837 (N_8837,N_6059,N_6075);
or U8838 (N_8838,N_7044,N_6026);
nor U8839 (N_8839,N_7428,N_7384);
and U8840 (N_8840,N_6332,N_7457);
nand U8841 (N_8841,N_7369,N_6684);
xnor U8842 (N_8842,N_6009,N_6418);
or U8843 (N_8843,N_6360,N_6044);
nor U8844 (N_8844,N_6373,N_6392);
or U8845 (N_8845,N_6660,N_6587);
nand U8846 (N_8846,N_6423,N_7140);
nor U8847 (N_8847,N_7182,N_6684);
nor U8848 (N_8848,N_7224,N_6159);
or U8849 (N_8849,N_7215,N_6053);
and U8850 (N_8850,N_6390,N_6872);
nor U8851 (N_8851,N_6725,N_6876);
xor U8852 (N_8852,N_6754,N_7248);
and U8853 (N_8853,N_6081,N_7351);
xnor U8854 (N_8854,N_7059,N_7235);
and U8855 (N_8855,N_7408,N_7291);
or U8856 (N_8856,N_6342,N_6640);
nor U8857 (N_8857,N_6578,N_7185);
and U8858 (N_8858,N_7262,N_6915);
xnor U8859 (N_8859,N_7222,N_7345);
and U8860 (N_8860,N_6278,N_6244);
or U8861 (N_8861,N_7356,N_7024);
or U8862 (N_8862,N_7155,N_7017);
xnor U8863 (N_8863,N_6622,N_6505);
nand U8864 (N_8864,N_6154,N_6987);
or U8865 (N_8865,N_6990,N_6490);
xor U8866 (N_8866,N_6005,N_7207);
nor U8867 (N_8867,N_6639,N_6521);
nor U8868 (N_8868,N_6631,N_6000);
and U8869 (N_8869,N_6034,N_6195);
xor U8870 (N_8870,N_6313,N_7183);
xor U8871 (N_8871,N_6376,N_7248);
or U8872 (N_8872,N_6234,N_7189);
xnor U8873 (N_8873,N_6568,N_6116);
nor U8874 (N_8874,N_7491,N_6535);
and U8875 (N_8875,N_6651,N_6751);
nor U8876 (N_8876,N_6625,N_6445);
nand U8877 (N_8877,N_6898,N_7380);
nor U8878 (N_8878,N_7292,N_6518);
nor U8879 (N_8879,N_7423,N_6746);
xnor U8880 (N_8880,N_6103,N_6327);
and U8881 (N_8881,N_7221,N_6640);
nor U8882 (N_8882,N_6836,N_6400);
nand U8883 (N_8883,N_6610,N_6034);
or U8884 (N_8884,N_6974,N_7414);
or U8885 (N_8885,N_7037,N_6372);
or U8886 (N_8886,N_6067,N_6640);
and U8887 (N_8887,N_7359,N_7410);
xor U8888 (N_8888,N_7338,N_6715);
xor U8889 (N_8889,N_6059,N_7412);
nor U8890 (N_8890,N_6883,N_6623);
xor U8891 (N_8891,N_7080,N_6324);
or U8892 (N_8892,N_7224,N_7451);
nand U8893 (N_8893,N_7464,N_6468);
nand U8894 (N_8894,N_6799,N_7247);
and U8895 (N_8895,N_6469,N_6231);
and U8896 (N_8896,N_7324,N_6236);
or U8897 (N_8897,N_7175,N_6919);
nand U8898 (N_8898,N_7299,N_7251);
and U8899 (N_8899,N_7164,N_6841);
and U8900 (N_8900,N_6894,N_6852);
xnor U8901 (N_8901,N_6017,N_7313);
xor U8902 (N_8902,N_6312,N_6627);
nor U8903 (N_8903,N_7038,N_6078);
nand U8904 (N_8904,N_6025,N_7381);
nand U8905 (N_8905,N_7187,N_6726);
and U8906 (N_8906,N_7073,N_6140);
xnor U8907 (N_8907,N_6383,N_7468);
nand U8908 (N_8908,N_6013,N_7020);
nor U8909 (N_8909,N_7425,N_6314);
and U8910 (N_8910,N_7053,N_6113);
nor U8911 (N_8911,N_6645,N_7457);
xnor U8912 (N_8912,N_6465,N_7006);
or U8913 (N_8913,N_6294,N_6397);
or U8914 (N_8914,N_6156,N_6381);
nor U8915 (N_8915,N_6319,N_6724);
nand U8916 (N_8916,N_7123,N_6065);
xor U8917 (N_8917,N_6873,N_6370);
xnor U8918 (N_8918,N_6313,N_6374);
nor U8919 (N_8919,N_6402,N_7080);
or U8920 (N_8920,N_6795,N_7152);
and U8921 (N_8921,N_6995,N_6666);
xnor U8922 (N_8922,N_6929,N_6514);
nand U8923 (N_8923,N_6112,N_6867);
and U8924 (N_8924,N_7441,N_6296);
and U8925 (N_8925,N_6666,N_7439);
xor U8926 (N_8926,N_6818,N_7448);
and U8927 (N_8927,N_6628,N_6324);
and U8928 (N_8928,N_6258,N_7409);
and U8929 (N_8929,N_7150,N_6586);
xnor U8930 (N_8930,N_7160,N_7142);
nor U8931 (N_8931,N_6869,N_6791);
nand U8932 (N_8932,N_6701,N_6142);
or U8933 (N_8933,N_7339,N_6084);
nor U8934 (N_8934,N_6235,N_7102);
nand U8935 (N_8935,N_6674,N_6860);
xor U8936 (N_8936,N_6071,N_7148);
and U8937 (N_8937,N_6162,N_6703);
and U8938 (N_8938,N_6949,N_7106);
or U8939 (N_8939,N_6289,N_6781);
or U8940 (N_8940,N_6188,N_6414);
or U8941 (N_8941,N_6855,N_7076);
xnor U8942 (N_8942,N_6475,N_7031);
xnor U8943 (N_8943,N_6563,N_6955);
or U8944 (N_8944,N_6837,N_7223);
nor U8945 (N_8945,N_6072,N_7257);
and U8946 (N_8946,N_6794,N_6459);
nand U8947 (N_8947,N_6434,N_7292);
and U8948 (N_8948,N_7449,N_7320);
and U8949 (N_8949,N_7130,N_6467);
nand U8950 (N_8950,N_6726,N_7238);
nor U8951 (N_8951,N_6839,N_6813);
xnor U8952 (N_8952,N_6062,N_6746);
nand U8953 (N_8953,N_6645,N_6467);
or U8954 (N_8954,N_6797,N_7174);
nand U8955 (N_8955,N_6175,N_6449);
nor U8956 (N_8956,N_6275,N_7395);
and U8957 (N_8957,N_6420,N_6338);
or U8958 (N_8958,N_6937,N_6074);
nand U8959 (N_8959,N_6226,N_6020);
xnor U8960 (N_8960,N_7472,N_7142);
nand U8961 (N_8961,N_6464,N_6450);
or U8962 (N_8962,N_7396,N_7478);
nor U8963 (N_8963,N_6933,N_6684);
xor U8964 (N_8964,N_6440,N_6885);
xor U8965 (N_8965,N_6426,N_6233);
nor U8966 (N_8966,N_6515,N_7021);
xnor U8967 (N_8967,N_7446,N_6984);
nand U8968 (N_8968,N_6894,N_6851);
or U8969 (N_8969,N_7322,N_6471);
and U8970 (N_8970,N_6088,N_6333);
or U8971 (N_8971,N_6887,N_6452);
nor U8972 (N_8972,N_6261,N_6896);
or U8973 (N_8973,N_6129,N_6518);
nor U8974 (N_8974,N_7127,N_6214);
nand U8975 (N_8975,N_6497,N_6184);
and U8976 (N_8976,N_7235,N_6115);
xor U8977 (N_8977,N_7242,N_6904);
xor U8978 (N_8978,N_6480,N_6140);
xnor U8979 (N_8979,N_6185,N_6873);
or U8980 (N_8980,N_6421,N_6274);
nand U8981 (N_8981,N_6085,N_6147);
nor U8982 (N_8982,N_6353,N_6833);
nand U8983 (N_8983,N_7088,N_7479);
and U8984 (N_8984,N_7158,N_6384);
nor U8985 (N_8985,N_7034,N_6030);
xnor U8986 (N_8986,N_7055,N_7224);
xnor U8987 (N_8987,N_6868,N_6802);
and U8988 (N_8988,N_6167,N_6230);
nand U8989 (N_8989,N_6585,N_6879);
nand U8990 (N_8990,N_6402,N_7118);
and U8991 (N_8991,N_6629,N_7122);
xor U8992 (N_8992,N_6725,N_7177);
nor U8993 (N_8993,N_7320,N_7390);
nor U8994 (N_8994,N_7142,N_7322);
nand U8995 (N_8995,N_6099,N_6360);
nor U8996 (N_8996,N_7469,N_7073);
xor U8997 (N_8997,N_6617,N_7293);
xor U8998 (N_8998,N_6184,N_7276);
xor U8999 (N_8999,N_7223,N_7258);
and U9000 (N_9000,N_7853,N_8270);
nand U9001 (N_9001,N_8819,N_8261);
or U9002 (N_9002,N_7822,N_8627);
xor U9003 (N_9003,N_8702,N_7752);
nand U9004 (N_9004,N_8016,N_8785);
xor U9005 (N_9005,N_8432,N_8254);
nand U9006 (N_9006,N_7651,N_8750);
and U9007 (N_9007,N_7560,N_8346);
and U9008 (N_9008,N_7602,N_7570);
nand U9009 (N_9009,N_8128,N_8781);
and U9010 (N_9010,N_8307,N_8713);
nor U9011 (N_9011,N_8291,N_8966);
nor U9012 (N_9012,N_8593,N_8917);
nand U9013 (N_9013,N_8398,N_8075);
nand U9014 (N_9014,N_7512,N_7897);
nor U9015 (N_9015,N_8096,N_7900);
or U9016 (N_9016,N_7719,N_8210);
and U9017 (N_9017,N_8960,N_8863);
xnor U9018 (N_9018,N_8453,N_8789);
nand U9019 (N_9019,N_8737,N_7640);
and U9020 (N_9020,N_8242,N_8859);
nand U9021 (N_9021,N_8824,N_8915);
nand U9022 (N_9022,N_7707,N_7524);
or U9023 (N_9023,N_8431,N_8900);
xnor U9024 (N_9024,N_7717,N_7726);
or U9025 (N_9025,N_8287,N_7561);
nor U9026 (N_9026,N_8415,N_7982);
or U9027 (N_9027,N_7873,N_7905);
or U9028 (N_9028,N_8473,N_8818);
xnor U9029 (N_9029,N_7501,N_8102);
nand U9030 (N_9030,N_8314,N_8620);
and U9031 (N_9031,N_8215,N_8400);
xnor U9032 (N_9032,N_8249,N_7795);
nand U9033 (N_9033,N_8526,N_8097);
and U9034 (N_9034,N_7755,N_8050);
xor U9035 (N_9035,N_7591,N_8366);
xnor U9036 (N_9036,N_8013,N_7589);
or U9037 (N_9037,N_8543,N_8391);
and U9038 (N_9038,N_8740,N_8823);
xor U9039 (N_9039,N_8082,N_8681);
xor U9040 (N_9040,N_8065,N_8485);
and U9041 (N_9041,N_8762,N_8411);
xnor U9042 (N_9042,N_7509,N_8561);
or U9043 (N_9043,N_8035,N_8961);
nor U9044 (N_9044,N_7709,N_7886);
nor U9045 (N_9045,N_8110,N_7653);
nor U9046 (N_9046,N_8157,N_8976);
nor U9047 (N_9047,N_8940,N_7605);
or U9048 (N_9048,N_8293,N_8661);
nor U9049 (N_9049,N_7908,N_7706);
nor U9050 (N_9050,N_8266,N_8421);
nand U9051 (N_9051,N_8038,N_7929);
xor U9052 (N_9052,N_8171,N_7997);
xor U9053 (N_9053,N_7939,N_8583);
or U9054 (N_9054,N_8904,N_8780);
nor U9055 (N_9055,N_7848,N_7926);
nor U9056 (N_9056,N_8448,N_7614);
xor U9057 (N_9057,N_8711,N_8241);
nor U9058 (N_9058,N_8497,N_8813);
nor U9059 (N_9059,N_7723,N_7683);
nor U9060 (N_9060,N_7981,N_8380);
xor U9061 (N_9061,N_7789,N_8848);
nor U9062 (N_9062,N_8343,N_8401);
xor U9063 (N_9063,N_8507,N_8897);
nand U9064 (N_9064,N_7979,N_7962);
or U9065 (N_9065,N_8833,N_8659);
xnor U9066 (N_9066,N_8150,N_7736);
or U9067 (N_9067,N_7828,N_8870);
nor U9068 (N_9068,N_8779,N_8498);
xor U9069 (N_9069,N_8902,N_8825);
xor U9070 (N_9070,N_7597,N_7663);
nand U9071 (N_9071,N_8049,N_7904);
nor U9072 (N_9072,N_8995,N_8461);
nand U9073 (N_9073,N_7955,N_7753);
nor U9074 (N_9074,N_8036,N_8696);
xor U9075 (N_9075,N_8137,N_8131);
or U9076 (N_9076,N_8104,N_8878);
xnor U9077 (N_9077,N_7840,N_8073);
nand U9078 (N_9078,N_8505,N_8258);
or U9079 (N_9079,N_8449,N_7680);
or U9080 (N_9080,N_7563,N_8211);
or U9081 (N_9081,N_8080,N_8268);
xor U9082 (N_9082,N_8633,N_7548);
nor U9083 (N_9083,N_7807,N_8120);
and U9084 (N_9084,N_8152,N_7628);
xor U9085 (N_9085,N_7880,N_7928);
nand U9086 (N_9086,N_8812,N_7881);
and U9087 (N_9087,N_8584,N_7586);
or U9088 (N_9088,N_8581,N_8807);
and U9089 (N_9089,N_8410,N_7660);
nor U9090 (N_9090,N_7610,N_8362);
nand U9091 (N_9091,N_8865,N_8041);
xnor U9092 (N_9092,N_7882,N_8020);
and U9093 (N_9093,N_8850,N_8969);
nand U9094 (N_9094,N_8439,N_8198);
and U9095 (N_9095,N_8325,N_8980);
nor U9096 (N_9096,N_8316,N_8838);
nor U9097 (N_9097,N_8193,N_8423);
nand U9098 (N_9098,N_7537,N_8712);
nor U9099 (N_9099,N_8376,N_8125);
or U9100 (N_9100,N_8588,N_8079);
and U9101 (N_9101,N_7808,N_7885);
nor U9102 (N_9102,N_7895,N_7549);
or U9103 (N_9103,N_7918,N_8668);
or U9104 (N_9104,N_8269,N_8603);
and U9105 (N_9105,N_8534,N_7684);
nand U9106 (N_9106,N_8801,N_8541);
and U9107 (N_9107,N_8882,N_8914);
and U9108 (N_9108,N_8177,N_7698);
xor U9109 (N_9109,N_8630,N_8933);
or U9110 (N_9110,N_8221,N_8414);
nor U9111 (N_9111,N_8271,N_7661);
nor U9112 (N_9112,N_7571,N_8965);
xor U9113 (N_9113,N_8085,N_7600);
and U9114 (N_9114,N_8433,N_7824);
or U9115 (N_9115,N_8815,N_8623);
xor U9116 (N_9116,N_8679,N_8790);
and U9117 (N_9117,N_7843,N_8393);
and U9118 (N_9118,N_8354,N_8090);
and U9119 (N_9119,N_8178,N_8014);
or U9120 (N_9120,N_8123,N_7662);
and U9121 (N_9121,N_7894,N_8235);
nor U9122 (N_9122,N_8800,N_8992);
xor U9123 (N_9123,N_7791,N_8109);
and U9124 (N_9124,N_7629,N_8430);
nand U9125 (N_9125,N_7656,N_8911);
nor U9126 (N_9126,N_8246,N_7826);
nand U9127 (N_9127,N_8635,N_8662);
nor U9128 (N_9128,N_8412,N_8309);
and U9129 (N_9129,N_8394,N_7715);
xor U9130 (N_9130,N_7788,N_7971);
nand U9131 (N_9131,N_8738,N_7530);
nor U9132 (N_9132,N_8765,N_7952);
xnor U9133 (N_9133,N_7510,N_8143);
xnor U9134 (N_9134,N_8548,N_8753);
xnor U9135 (N_9135,N_8010,N_8760);
nor U9136 (N_9136,N_8745,N_7506);
nor U9137 (N_9137,N_8579,N_8338);
xor U9138 (N_9138,N_8467,N_8634);
and U9139 (N_9139,N_8536,N_8606);
nor U9140 (N_9140,N_8101,N_7677);
or U9141 (N_9141,N_7500,N_8283);
or U9142 (N_9142,N_8893,N_7859);
and U9143 (N_9143,N_7792,N_8926);
xor U9144 (N_9144,N_7575,N_7743);
nor U9145 (N_9145,N_7737,N_8272);
xnor U9146 (N_9146,N_8000,N_7849);
and U9147 (N_9147,N_7529,N_8564);
or U9148 (N_9148,N_8227,N_7767);
and U9149 (N_9149,N_7672,N_7654);
nor U9150 (N_9150,N_7691,N_8983);
and U9151 (N_9151,N_8032,N_7572);
nand U9152 (N_9152,N_8234,N_8512);
and U9153 (N_9153,N_7593,N_7784);
nand U9154 (N_9154,N_8490,N_8127);
and U9155 (N_9155,N_7679,N_7686);
or U9156 (N_9156,N_8250,N_8788);
nor U9157 (N_9157,N_7712,N_8726);
and U9158 (N_9158,N_7626,N_8098);
nand U9159 (N_9159,N_8912,N_7527);
xor U9160 (N_9160,N_8087,N_8532);
or U9161 (N_9161,N_8697,N_8390);
nor U9162 (N_9162,N_7727,N_8628);
nand U9163 (N_9163,N_8600,N_8347);
nor U9164 (N_9164,N_8670,N_8148);
xnor U9165 (N_9165,N_8169,N_7724);
nor U9166 (N_9166,N_8147,N_8315);
nor U9167 (N_9167,N_7794,N_8442);
xnor U9168 (N_9168,N_8744,N_8212);
and U9169 (N_9169,N_8359,N_8903);
nor U9170 (N_9170,N_7685,N_7811);
xor U9171 (N_9171,N_7985,N_8365);
or U9172 (N_9172,N_8048,N_8948);
and U9173 (N_9173,N_7934,N_7528);
and U9174 (N_9174,N_7816,N_8378);
nor U9175 (N_9175,N_8407,N_8674);
nor U9176 (N_9176,N_8067,N_7809);
and U9177 (N_9177,N_8886,N_8806);
and U9178 (N_9178,N_7821,N_8290);
nor U9179 (N_9179,N_7925,N_7523);
nand U9180 (N_9180,N_8220,N_8786);
and U9181 (N_9181,N_8066,N_7995);
nand U9182 (N_9182,N_8846,N_8970);
nand U9183 (N_9183,N_7573,N_8962);
nor U9184 (N_9184,N_8129,N_8099);
xor U9185 (N_9185,N_8729,N_8340);
or U9186 (N_9186,N_8351,N_7567);
nand U9187 (N_9187,N_8121,N_7568);
xnor U9188 (N_9188,N_7692,N_8070);
xnor U9189 (N_9189,N_8213,N_8208);
nor U9190 (N_9190,N_8621,N_8769);
or U9191 (N_9191,N_8420,N_7675);
nor U9192 (N_9192,N_8587,N_7915);
xnor U9193 (N_9193,N_8476,N_8292);
nor U9194 (N_9194,N_8923,N_7787);
nor U9195 (N_9195,N_7750,N_8231);
xor U9196 (N_9196,N_8791,N_8763);
xnor U9197 (N_9197,N_8454,N_7766);
xor U9198 (N_9198,N_8182,N_8689);
xnor U9199 (N_9199,N_8030,N_8530);
xor U9200 (N_9200,N_7992,N_8792);
xor U9201 (N_9201,N_8667,N_7746);
or U9202 (N_9202,N_7818,N_8081);
nand U9203 (N_9203,N_7862,N_8011);
xor U9204 (N_9204,N_8286,N_7508);
or U9205 (N_9205,N_8611,N_7919);
nand U9206 (N_9206,N_7790,N_8112);
xor U9207 (N_9207,N_8440,N_7837);
and U9208 (N_9208,N_8984,N_8409);
and U9209 (N_9209,N_7596,N_7768);
nand U9210 (N_9210,N_8925,N_8331);
nand U9211 (N_9211,N_8861,N_8710);
or U9212 (N_9212,N_8179,N_8063);
xor U9213 (N_9213,N_7973,N_7783);
or U9214 (N_9214,N_7899,N_8388);
nor U9215 (N_9215,N_7940,N_8385);
and U9216 (N_9216,N_8648,N_8799);
nand U9217 (N_9217,N_8350,N_7913);
nand U9218 (N_9218,N_7810,N_8489);
and U9219 (N_9219,N_8219,N_8285);
or U9220 (N_9220,N_8739,N_8209);
xor U9221 (N_9221,N_8238,N_7613);
nand U9222 (N_9222,N_8071,N_8168);
or U9223 (N_9223,N_8342,N_8529);
and U9224 (N_9224,N_7503,N_8578);
nor U9225 (N_9225,N_8397,N_8173);
and U9226 (N_9226,N_7565,N_8721);
xnor U9227 (N_9227,N_8462,N_7583);
nor U9228 (N_9228,N_8021,N_8972);
and U9229 (N_9229,N_7553,N_8226);
nor U9230 (N_9230,N_8160,N_8869);
and U9231 (N_9231,N_7650,N_7517);
or U9232 (N_9232,N_8973,N_8503);
nand U9233 (N_9233,N_8988,N_8422);
and U9234 (N_9234,N_8263,N_7731);
nor U9235 (N_9235,N_7936,N_7927);
xor U9236 (N_9236,N_8051,N_8959);
nand U9237 (N_9237,N_8308,N_8332);
xor U9238 (N_9238,N_7638,N_8054);
nand U9239 (N_9239,N_8488,N_8426);
and U9240 (N_9240,N_8985,N_7521);
nor U9241 (N_9241,N_8282,N_8688);
xor U9242 (N_9242,N_8591,N_8652);
and U9243 (N_9243,N_8544,N_7742);
and U9244 (N_9244,N_8336,N_8055);
or U9245 (N_9245,N_8187,N_8967);
or U9246 (N_9246,N_8546,N_8370);
and U9247 (N_9247,N_8368,N_8577);
and U9248 (N_9248,N_8749,N_8909);
nand U9249 (N_9249,N_8906,N_8408);
nor U9250 (N_9250,N_8664,N_8899);
or U9251 (N_9251,N_8138,N_8733);
nand U9252 (N_9252,N_8344,N_7556);
nand U9253 (N_9253,N_7612,N_7907);
nand U9254 (N_9254,N_7889,N_7765);
and U9255 (N_9255,N_7544,N_8236);
xor U9256 (N_9256,N_8253,N_8078);
nor U9257 (N_9257,N_8974,N_8665);
and U9258 (N_9258,N_8977,N_7836);
nor U9259 (N_9259,N_8164,N_8306);
nor U9260 (N_9260,N_8758,N_8542);
xnor U9261 (N_9261,N_8317,N_8436);
nor U9262 (N_9262,N_7869,N_8624);
xor U9263 (N_9263,N_8480,N_8279);
nand U9264 (N_9264,N_8170,N_7676);
nand U9265 (N_9265,N_8596,N_7857);
or U9266 (N_9266,N_8319,N_8284);
xor U9267 (N_9267,N_8997,N_7655);
nand U9268 (N_9268,N_8517,N_8954);
nand U9269 (N_9269,N_7956,N_7999);
nor U9270 (N_9270,N_7621,N_8845);
or U9271 (N_9271,N_8894,N_8704);
or U9272 (N_9272,N_8708,N_7892);
or U9273 (N_9273,N_8192,N_8558);
or U9274 (N_9274,N_8715,N_8553);
and U9275 (N_9275,N_7964,N_8853);
and U9276 (N_9276,N_8029,N_7633);
nand U9277 (N_9277,N_7631,N_8794);
and U9278 (N_9278,N_8040,N_8849);
nand U9279 (N_9279,N_8165,N_8053);
xor U9280 (N_9280,N_8022,N_8056);
nor U9281 (N_9281,N_7734,N_8932);
nand U9282 (N_9282,N_8262,N_7515);
xnor U9283 (N_9283,N_7601,N_8993);
nand U9284 (N_9284,N_7938,N_8951);
nor U9285 (N_9285,N_8255,N_8881);
nor U9286 (N_9286,N_8264,N_7946);
nand U9287 (N_9287,N_8039,N_8660);
xor U9288 (N_9288,N_8206,N_7536);
or U9289 (N_9289,N_8994,N_8384);
and U9290 (N_9290,N_7541,N_8130);
xor U9291 (N_9291,N_8990,N_8451);
and U9292 (N_9292,N_7786,N_8278);
nor U9293 (N_9293,N_7958,N_8329);
and U9294 (N_9294,N_8636,N_7696);
nor U9295 (N_9295,N_8741,N_8327);
or U9296 (N_9296,N_7967,N_8772);
or U9297 (N_9297,N_8883,N_7785);
or U9298 (N_9298,N_8026,N_8417);
nor U9299 (N_9299,N_7671,N_8244);
nand U9300 (N_9300,N_7701,N_8999);
xor U9301 (N_9301,N_8568,N_7961);
nor U9302 (N_9302,N_7643,N_8392);
nor U9303 (N_9303,N_8537,N_8920);
xor U9304 (N_9304,N_7942,N_8381);
nand U9305 (N_9305,N_7998,N_7987);
nor U9306 (N_9306,N_7749,N_8686);
nor U9307 (N_9307,N_8831,N_8116);
or U9308 (N_9308,N_8019,N_8939);
or U9309 (N_9309,N_8607,N_8747);
or U9310 (N_9310,N_7815,N_7745);
and U9311 (N_9311,N_8770,N_8533);
or U9312 (N_9312,N_8144,N_7825);
xnor U9313 (N_9313,N_8191,N_7806);
and U9314 (N_9314,N_7834,N_8673);
and U9315 (N_9315,N_8303,N_8028);
and U9316 (N_9316,N_8119,N_7874);
and U9317 (N_9317,N_8465,N_8678);
nand U9318 (N_9318,N_8434,N_8455);
nor U9319 (N_9319,N_7920,N_8535);
and U9320 (N_9320,N_8683,N_8690);
and U9321 (N_9321,N_8377,N_8547);
nor U9322 (N_9322,N_7850,N_8851);
nand U9323 (N_9323,N_8438,N_8924);
xor U9324 (N_9324,N_7871,N_8330);
nor U9325 (N_9325,N_7805,N_8570);
and U9326 (N_9326,N_7914,N_7921);
xnor U9327 (N_9327,N_8222,N_7812);
nand U9328 (N_9328,N_8816,N_7797);
nor U9329 (N_9329,N_8281,N_7770);
nand U9330 (N_9330,N_8829,N_8200);
xnor U9331 (N_9331,N_7716,N_8566);
nand U9332 (N_9332,N_7851,N_8416);
xor U9333 (N_9333,N_8632,N_8515);
and U9334 (N_9334,N_8294,N_7539);
nor U9335 (N_9335,N_8217,N_7522);
or U9336 (N_9336,N_8625,N_8650);
nor U9337 (N_9337,N_7923,N_8093);
nand U9338 (N_9338,N_8842,N_7681);
nor U9339 (N_9339,N_8975,N_7877);
or U9340 (N_9340,N_8511,N_8864);
and U9341 (N_9341,N_7801,N_8345);
and U9342 (N_9342,N_8509,N_7514);
and U9343 (N_9343,N_8840,N_7838);
nor U9344 (N_9344,N_8405,N_8117);
nand U9345 (N_9345,N_7953,N_8274);
or U9346 (N_9346,N_8725,N_7728);
or U9347 (N_9347,N_7798,N_8761);
xor U9348 (N_9348,N_8224,N_8204);
nor U9349 (N_9349,N_8172,N_8874);
and U9350 (N_9350,N_8134,N_8707);
nor U9351 (N_9351,N_8855,N_8240);
and U9352 (N_9352,N_8484,N_8887);
or U9353 (N_9353,N_8580,N_8671);
or U9354 (N_9354,N_8867,N_8756);
nor U9355 (N_9355,N_8444,N_8888);
and U9356 (N_9356,N_8202,N_8706);
nand U9357 (N_9357,N_7930,N_7625);
or U9358 (N_9358,N_7518,N_7710);
nand U9359 (N_9359,N_8701,N_7866);
xnor U9360 (N_9360,N_8590,N_7933);
nand U9361 (N_9361,N_8176,N_7619);
nor U9362 (N_9362,N_8379,N_7963);
nor U9363 (N_9363,N_8225,N_7996);
or U9364 (N_9364,N_8002,N_7846);
nand U9365 (N_9365,N_7659,N_8692);
nand U9366 (N_9366,N_8037,N_7901);
nor U9367 (N_9367,N_8399,N_7988);
and U9368 (N_9368,N_7757,N_7665);
nand U9369 (N_9369,N_7781,N_8305);
and U9370 (N_9370,N_8796,N_7504);
xnor U9371 (N_9371,N_8699,N_8539);
nor U9372 (N_9372,N_7703,N_8716);
nand U9373 (N_9373,N_8328,N_7608);
and U9374 (N_9374,N_7616,N_8337);
or U9375 (N_9375,N_8901,N_8310);
nor U9376 (N_9376,N_8095,N_8797);
or U9377 (N_9377,N_8514,N_8520);
or U9378 (N_9378,N_7554,N_8300);
and U9379 (N_9379,N_8554,N_8989);
or U9380 (N_9380,N_8868,N_8839);
nand U9381 (N_9381,N_8425,N_8871);
or U9382 (N_9382,N_8730,N_7804);
nor U9383 (N_9383,N_8356,N_8647);
xor U9384 (N_9384,N_8614,N_7759);
or U9385 (N_9385,N_8736,N_8248);
nor U9386 (N_9386,N_7764,N_8754);
nand U9387 (N_9387,N_8827,N_7668);
xor U9388 (N_9388,N_7902,N_7772);
nor U9389 (N_9389,N_8069,N_8044);
nor U9390 (N_9390,N_8031,N_8913);
xnor U9391 (N_9391,N_8188,N_8012);
nor U9392 (N_9392,N_8348,N_7636);
or U9393 (N_9393,N_7931,N_8991);
and U9394 (N_9394,N_7690,N_8709);
nor U9395 (N_9395,N_7694,N_7688);
nor U9396 (N_9396,N_8086,N_8857);
or U9397 (N_9397,N_7558,N_7863);
xor U9398 (N_9398,N_8928,N_8675);
or U9399 (N_9399,N_8445,N_8589);
and U9400 (N_9400,N_8477,N_8252);
and U9401 (N_9401,N_8251,N_7891);
nor U9402 (N_9402,N_8927,N_8302);
nor U9403 (N_9403,N_8513,N_8201);
nand U9404 (N_9404,N_8180,N_8575);
xnor U9405 (N_9405,N_8685,N_7776);
or U9406 (N_9406,N_7546,N_8396);
xnor U9407 (N_9407,N_7584,N_8207);
nand U9408 (N_9408,N_8622,N_8427);
nand U9409 (N_9409,N_8321,N_8540);
or U9410 (N_9410,N_8907,N_8460);
nor U9411 (N_9411,N_7947,N_7858);
nor U9412 (N_9412,N_8245,N_8804);
nand U9413 (N_9413,N_7578,N_7855);
nand U9414 (N_9414,N_8656,N_8826);
nor U9415 (N_9415,N_8929,N_8091);
nor U9416 (N_9416,N_7603,N_8835);
or U9417 (N_9417,N_8156,N_8830);
and U9418 (N_9418,N_7802,N_8854);
xnor U9419 (N_9419,N_7666,N_8617);
nor U9420 (N_9420,N_8776,N_7576);
xnor U9421 (N_9421,N_8931,N_8259);
xnor U9422 (N_9422,N_8731,N_7994);
nand U9423 (N_9423,N_8778,N_8952);
nor U9424 (N_9424,N_7718,N_7909);
xor U9425 (N_9425,N_8684,N_8382);
nand U9426 (N_9426,N_8956,N_7898);
nor U9427 (N_9427,N_7965,N_7569);
nand U9428 (N_9428,N_8482,N_8717);
nor U9429 (N_9429,N_8705,N_8809);
or U9430 (N_9430,N_7714,N_7562);
and U9431 (N_9431,N_7657,N_8657);
and U9432 (N_9432,N_7552,N_7580);
xnor U9433 (N_9433,N_8103,N_8277);
nor U9434 (N_9434,N_8518,N_7951);
or U9435 (N_9435,N_8371,N_8654);
or U9436 (N_9436,N_7989,N_7689);
xor U9437 (N_9437,N_7754,N_8446);
xnor U9438 (N_9438,N_8203,N_8162);
nor U9439 (N_9439,N_7827,N_8122);
xor U9440 (N_9440,N_7673,N_8146);
nand U9441 (N_9441,N_7835,N_8885);
nor U9442 (N_9442,N_8805,N_7954);
xor U9443 (N_9443,N_8549,N_8074);
xnor U9444 (N_9444,N_8986,N_8471);
nor U9445 (N_9445,N_8437,N_8149);
and U9446 (N_9446,N_8061,N_8950);
nand U9447 (N_9447,N_7547,N_8774);
and U9448 (N_9448,N_8493,N_8185);
xor U9449 (N_9449,N_8458,N_8218);
nor U9450 (N_9450,N_8937,N_8189);
nand U9451 (N_9451,N_7648,N_7511);
or U9452 (N_9452,N_8979,N_8527);
xor U9453 (N_9453,N_8586,N_8230);
nor U9454 (N_9454,N_8059,N_8486);
and U9455 (N_9455,N_7559,N_7819);
or U9456 (N_9456,N_8111,N_8510);
and U9457 (N_9457,N_8357,N_7704);
nor U9458 (N_9458,N_8042,N_8299);
or U9459 (N_9459,N_8304,N_8602);
xnor U9460 (N_9460,N_7916,N_7888);
nor U9461 (N_9461,N_8556,N_8256);
or U9462 (N_9462,N_8229,N_8113);
xnor U9463 (N_9463,N_7760,N_8934);
or U9464 (N_9464,N_7957,N_8413);
or U9465 (N_9465,N_8115,N_8677);
nand U9466 (N_9466,N_8076,N_8808);
or U9467 (N_9467,N_7800,N_7966);
or U9468 (N_9468,N_8793,N_8158);
nand U9469 (N_9469,N_8133,N_7639);
xnor U9470 (N_9470,N_8495,N_8429);
or U9471 (N_9471,N_8349,N_8077);
and U9472 (N_9472,N_7896,N_8508);
or U9473 (N_9473,N_8597,N_8060);
or U9474 (N_9474,N_8764,N_8610);
and U9475 (N_9475,N_7868,N_7856);
nand U9476 (N_9476,N_7598,N_7682);
or U9477 (N_9477,N_7630,N_7606);
and U9478 (N_9478,N_8008,N_7977);
nor U9479 (N_9479,N_8064,N_8612);
nor U9480 (N_9480,N_8135,N_8562);
nor U9481 (N_9481,N_7984,N_7738);
and U9482 (N_9482,N_8971,N_8574);
and U9483 (N_9483,N_7566,N_8441);
nor U9484 (N_9484,N_8599,N_7658);
xor U9485 (N_9485,N_8698,N_7972);
xnor U9486 (N_9486,N_8428,N_7551);
and U9487 (N_9487,N_8944,N_7588);
or U9488 (N_9488,N_8267,N_8223);
xnor U9489 (N_9489,N_8601,N_7813);
and U9490 (N_9490,N_8964,N_8297);
nor U9491 (N_9491,N_7970,N_8009);
and U9492 (N_9492,N_8862,N_8216);
nand U9493 (N_9493,N_8810,N_8908);
nor U9494 (N_9494,N_8296,N_7974);
nor U9495 (N_9495,N_8118,N_8418);
and U9496 (N_9496,N_7702,N_8619);
and U9497 (N_9497,N_8033,N_7543);
or U9498 (N_9498,N_7617,N_8167);
nand U9499 (N_9499,N_7950,N_8629);
or U9500 (N_9500,N_8866,N_8856);
nand U9501 (N_9501,N_8598,N_7581);
xor U9502 (N_9502,N_8884,N_8817);
nand U9503 (N_9503,N_8565,N_7879);
xor U9504 (N_9504,N_8483,N_8047);
xor U9505 (N_9505,N_8363,N_8007);
or U9506 (N_9506,N_8470,N_7618);
nand U9507 (N_9507,N_7599,N_8723);
nand U9508 (N_9508,N_8140,N_8094);
nand U9509 (N_9509,N_8742,N_7878);
nand U9510 (N_9510,N_8693,N_7649);
xnor U9511 (N_9511,N_7944,N_8555);
or U9512 (N_9512,N_7968,N_8214);
or U9513 (N_9513,N_8159,N_8298);
xor U9514 (N_9514,N_8642,N_7637);
xnor U9515 (N_9515,N_8355,N_8276);
nor U9516 (N_9516,N_8106,N_8771);
xor U9517 (N_9517,N_8595,N_8154);
nor U9518 (N_9518,N_8083,N_8746);
nor U9519 (N_9519,N_8957,N_8694);
or U9520 (N_9520,N_8194,N_7642);
nand U9521 (N_9521,N_8100,N_8573);
nor U9522 (N_9522,N_7645,N_7622);
nor U9523 (N_9523,N_7611,N_8424);
xnor U9524 (N_9524,N_8501,N_8232);
and U9525 (N_9525,N_8052,N_8001);
or U9526 (N_9526,N_8015,N_8773);
nor U9527 (N_9527,N_7519,N_7609);
or U9528 (N_9528,N_7579,N_8237);
or U9529 (N_9529,N_7587,N_8034);
nand U9530 (N_9530,N_7711,N_8666);
nor U9531 (N_9531,N_7713,N_8360);
nand U9532 (N_9532,N_8492,N_8889);
nand U9533 (N_9533,N_8528,N_7820);
or U9534 (N_9534,N_8481,N_8639);
and U9535 (N_9535,N_8843,N_8643);
xnor U9536 (N_9536,N_8641,N_8858);
and U9537 (N_9537,N_8720,N_8576);
nand U9538 (N_9538,N_7604,N_8186);
xor U9539 (N_9539,N_8672,N_7670);
xnor U9540 (N_9540,N_8891,N_7779);
nand U9541 (N_9541,N_8978,N_8335);
nand U9542 (N_9542,N_8943,N_8089);
xor U9543 (N_9543,N_8025,N_7730);
nand U9544 (N_9544,N_8538,N_8727);
or U9545 (N_9545,N_8872,N_7761);
nand U9546 (N_9546,N_8027,N_7635);
nor U9547 (N_9547,N_7782,N_8567);
nor U9548 (N_9548,N_7832,N_7763);
xnor U9549 (N_9549,N_7538,N_8844);
xnor U9550 (N_9550,N_8205,N_8402);
and U9551 (N_9551,N_7887,N_7864);
nor U9552 (N_9552,N_7872,N_8457);
or U9553 (N_9553,N_8582,N_7870);
nand U9554 (N_9554,N_7502,N_7993);
xnor U9555 (N_9555,N_8464,N_7883);
xnor U9556 (N_9556,N_8155,N_7793);
nor U9557 (N_9557,N_7695,N_8605);
xor U9558 (N_9558,N_8560,N_7669);
nor U9559 (N_9559,N_8372,N_7976);
nand U9560 (N_9560,N_8735,N_8452);
xor U9561 (N_9561,N_8719,N_8751);
and U9562 (N_9562,N_8691,N_8847);
or U9563 (N_9563,N_8166,N_7535);
nor U9564 (N_9564,N_8821,N_7540);
nor U9565 (N_9565,N_8334,N_7577);
nor U9566 (N_9566,N_7740,N_8880);
nand U9567 (N_9567,N_7935,N_7741);
nor U9568 (N_9568,N_8637,N_8728);
or U9569 (N_9569,N_8820,N_8775);
and U9570 (N_9570,N_8798,N_8126);
xor U9571 (N_9571,N_8879,N_8387);
xnor U9572 (N_9572,N_7735,N_7744);
and U9573 (N_9573,N_8557,N_8324);
or U9574 (N_9574,N_8982,N_7520);
nand U9575 (N_9575,N_8947,N_8873);
nor U9576 (N_9576,N_8921,N_8613);
or U9577 (N_9577,N_8499,N_8676);
and U9578 (N_9578,N_8353,N_8289);
and U9579 (N_9579,N_8163,N_8836);
and U9580 (N_9580,N_8531,N_7620);
nand U9581 (N_9581,N_7747,N_8124);
or U9582 (N_9582,N_8942,N_7842);
nand U9583 (N_9583,N_8935,N_7852);
nand U9584 (N_9584,N_8004,N_8875);
or U9585 (N_9585,N_7943,N_7632);
and U9586 (N_9586,N_8572,N_8644);
nor U9587 (N_9587,N_8174,N_7932);
and U9588 (N_9588,N_8139,N_8784);
and U9589 (N_9589,N_8748,N_7594);
xor U9590 (N_9590,N_8955,N_8197);
xnor U9591 (N_9591,N_8996,N_8386);
xor U9592 (N_9592,N_8898,N_8594);
or U9593 (N_9593,N_8803,N_7550);
nor U9594 (N_9594,N_8105,N_8640);
nand U9595 (N_9595,N_7721,N_8787);
or U9596 (N_9596,N_8062,N_7557);
and U9597 (N_9597,N_7861,N_8472);
and U9598 (N_9598,N_7980,N_8703);
xnor U9599 (N_9599,N_8058,N_8545);
nand U9600 (N_9600,N_8777,N_7564);
nand U9601 (N_9601,N_7774,N_8890);
or U9602 (N_9602,N_7555,N_7533);
xnor U9603 (N_9603,N_8318,N_7991);
and U9604 (N_9604,N_7796,N_7830);
nand U9605 (N_9605,N_8247,N_8003);
nor U9606 (N_9606,N_7725,N_7799);
nor U9607 (N_9607,N_8722,N_8953);
nor U9608 (N_9608,N_8968,N_8743);
and U9609 (N_9609,N_8447,N_7959);
nor U9610 (N_9610,N_8896,N_8153);
nand U9611 (N_9611,N_7641,N_7705);
nand U9612 (N_9612,N_8494,N_8195);
and U9613 (N_9613,N_8496,N_8136);
or U9614 (N_9614,N_7876,N_8522);
nor U9615 (N_9615,N_8841,N_8043);
nand U9616 (N_9616,N_8005,N_7960);
xor U9617 (N_9617,N_8759,N_8288);
or U9618 (N_9618,N_8895,N_8651);
nor U9619 (N_9619,N_8519,N_8687);
and U9620 (N_9620,N_8766,N_8521);
nand U9621 (N_9621,N_8456,N_8958);
nand U9622 (N_9622,N_8616,N_8404);
nor U9623 (N_9623,N_8822,N_8700);
and U9624 (N_9624,N_7590,N_8023);
nand U9625 (N_9625,N_8184,N_8233);
or U9626 (N_9626,N_8322,N_8320);
or U9627 (N_9627,N_7922,N_8468);
nand U9628 (N_9628,N_7615,N_8892);
nand U9629 (N_9629,N_7574,N_8311);
and U9630 (N_9630,N_8228,N_8280);
xor U9631 (N_9631,N_8569,N_8275);
and U9632 (N_9632,N_7937,N_7674);
nand U9633 (N_9633,N_7829,N_7906);
and U9634 (N_9634,N_8608,N_7911);
nand U9635 (N_9635,N_7945,N_8987);
nor U9636 (N_9636,N_8295,N_8383);
nand U9637 (N_9637,N_8714,N_8592);
or U9638 (N_9638,N_8945,N_8618);
or U9639 (N_9639,N_8474,N_8876);
nand U9640 (N_9640,N_8523,N_7693);
nor U9641 (N_9641,N_8190,N_8088);
or U9642 (N_9642,N_8132,N_7531);
xnor U9643 (N_9643,N_8585,N_7507);
nor U9644 (N_9644,N_8767,N_8443);
nand U9645 (N_9645,N_8491,N_8877);
or U9646 (N_9646,N_7729,N_8814);
or U9647 (N_9647,N_7623,N_8175);
nand U9648 (N_9648,N_8732,N_8466);
and U9649 (N_9649,N_7627,N_7983);
xnor U9650 (N_9650,N_8487,N_7733);
or U9651 (N_9651,N_7924,N_8369);
or U9652 (N_9652,N_8919,N_8755);
xnor U9653 (N_9653,N_8981,N_7844);
nand U9654 (N_9654,N_8918,N_8257);
xor U9655 (N_9655,N_8916,N_8389);
nor U9656 (N_9656,N_7860,N_7775);
nand U9657 (N_9657,N_8949,N_8183);
xor U9658 (N_9658,N_8516,N_8795);
and U9659 (N_9659,N_7646,N_8141);
and U9660 (N_9660,N_7678,N_8946);
xor U9661 (N_9661,N_8963,N_7516);
nor U9662 (N_9662,N_7582,N_7751);
or U9663 (N_9663,N_8046,N_7525);
and U9664 (N_9664,N_7762,N_8524);
xnor U9665 (N_9665,N_8017,N_8361);
nor U9666 (N_9666,N_7720,N_8367);
or U9667 (N_9667,N_7773,N_7526);
or U9668 (N_9668,N_8506,N_7534);
nand U9669 (N_9669,N_8341,N_7833);
nor U9670 (N_9670,N_7893,N_7756);
nor U9671 (N_9671,N_7780,N_8695);
nand U9672 (N_9672,N_7505,N_8718);
xnor U9673 (N_9673,N_8352,N_8551);
or U9674 (N_9674,N_8752,N_8323);
xor U9675 (N_9675,N_7910,N_8301);
xnor U9676 (N_9676,N_8459,N_7697);
or U9677 (N_9677,N_7803,N_7949);
or U9678 (N_9678,N_8682,N_8783);
nand U9679 (N_9679,N_8782,N_8604);
xnor U9680 (N_9680,N_7823,N_8658);
xor U9681 (N_9681,N_7700,N_8450);
or U9682 (N_9682,N_8419,N_8563);
xor U9683 (N_9683,N_7585,N_7990);
or U9684 (N_9684,N_8151,N_8358);
nor U9685 (N_9685,N_7875,N_8680);
and U9686 (N_9686,N_7814,N_8504);
or U9687 (N_9687,N_7732,N_8832);
xnor U9688 (N_9688,N_7917,N_8313);
and U9689 (N_9689,N_7903,N_8930);
or U9690 (N_9690,N_7652,N_8478);
nand U9691 (N_9691,N_8941,N_7978);
xor U9692 (N_9692,N_8406,N_8333);
and U9693 (N_9693,N_8828,N_8312);
nor U9694 (N_9694,N_8811,N_7644);
or U9695 (N_9695,N_7841,N_7831);
or U9696 (N_9696,N_7986,N_8626);
nor U9697 (N_9697,N_8006,N_8243);
nor U9698 (N_9698,N_8196,N_7771);
or U9699 (N_9699,N_8273,N_7708);
nand U9700 (N_9700,N_8018,N_7513);
or U9701 (N_9701,N_8550,N_8998);
nor U9702 (N_9702,N_7817,N_7592);
nor U9703 (N_9703,N_8649,N_7769);
nor U9704 (N_9704,N_8609,N_7975);
or U9705 (N_9705,N_8631,N_7948);
nor U9706 (N_9706,N_8559,N_8463);
and U9707 (N_9707,N_8435,N_8479);
and U9708 (N_9708,N_7664,N_8852);
and U9709 (N_9709,N_8108,N_8469);
nor U9710 (N_9710,N_7607,N_7758);
and U9711 (N_9711,N_8375,N_8114);
xnor U9712 (N_9712,N_8265,N_8142);
and U9713 (N_9713,N_7777,N_7845);
nor U9714 (N_9714,N_8475,N_8936);
and U9715 (N_9715,N_8024,N_8145);
and U9716 (N_9716,N_7890,N_8655);
and U9717 (N_9717,N_8373,N_7699);
or U9718 (N_9718,N_7595,N_8757);
xor U9719 (N_9719,N_8638,N_8669);
nor U9720 (N_9720,N_7847,N_8938);
nor U9721 (N_9721,N_8107,N_8768);
nor U9722 (N_9722,N_8326,N_7532);
nor U9723 (N_9723,N_8045,N_7839);
and U9724 (N_9724,N_8653,N_7748);
nor U9725 (N_9725,N_8395,N_7739);
and U9726 (N_9726,N_8834,N_8860);
xnor U9727 (N_9727,N_8571,N_8734);
nand U9728 (N_9728,N_8068,N_7884);
nor U9729 (N_9729,N_7867,N_8663);
or U9730 (N_9730,N_7624,N_8615);
and U9731 (N_9731,N_8910,N_7647);
nor U9732 (N_9732,N_7687,N_7912);
and U9733 (N_9733,N_8837,N_8724);
or U9734 (N_9734,N_8922,N_8525);
and U9735 (N_9735,N_8161,N_8239);
xnor U9736 (N_9736,N_7969,N_8181);
nor U9737 (N_9737,N_8802,N_7865);
nor U9738 (N_9738,N_8084,N_8092);
or U9739 (N_9739,N_7542,N_8374);
nand U9740 (N_9740,N_7941,N_7667);
and U9741 (N_9741,N_8364,N_8905);
or U9742 (N_9742,N_8646,N_8260);
and U9743 (N_9743,N_8645,N_8072);
or U9744 (N_9744,N_7722,N_8552);
xnor U9745 (N_9745,N_7634,N_8057);
xnor U9746 (N_9746,N_8500,N_7545);
nor U9747 (N_9747,N_8339,N_7778);
xnor U9748 (N_9748,N_7854,N_8403);
nor U9749 (N_9749,N_8502,N_8199);
or U9750 (N_9750,N_7726,N_8031);
nor U9751 (N_9751,N_8700,N_8156);
xor U9752 (N_9752,N_7940,N_8418);
nor U9753 (N_9753,N_7907,N_8600);
or U9754 (N_9754,N_8737,N_8648);
xnor U9755 (N_9755,N_7786,N_7789);
xor U9756 (N_9756,N_8879,N_8975);
xor U9757 (N_9757,N_8519,N_8267);
or U9758 (N_9758,N_8784,N_8581);
or U9759 (N_9759,N_8186,N_7553);
nand U9760 (N_9760,N_8657,N_7942);
or U9761 (N_9761,N_8467,N_7786);
or U9762 (N_9762,N_8547,N_8078);
and U9763 (N_9763,N_8656,N_8050);
and U9764 (N_9764,N_8888,N_8545);
nand U9765 (N_9765,N_8257,N_8978);
nor U9766 (N_9766,N_7894,N_8640);
nor U9767 (N_9767,N_8591,N_8857);
and U9768 (N_9768,N_8580,N_8874);
xnor U9769 (N_9769,N_7794,N_8421);
nand U9770 (N_9770,N_8070,N_8431);
xnor U9771 (N_9771,N_7845,N_7647);
xor U9772 (N_9772,N_8756,N_8190);
xnor U9773 (N_9773,N_8427,N_8219);
nand U9774 (N_9774,N_7589,N_8939);
nand U9775 (N_9775,N_8552,N_7771);
and U9776 (N_9776,N_7730,N_8128);
and U9777 (N_9777,N_7653,N_7708);
xnor U9778 (N_9778,N_7977,N_8333);
and U9779 (N_9779,N_8383,N_8656);
xnor U9780 (N_9780,N_8897,N_8162);
or U9781 (N_9781,N_8845,N_7648);
xor U9782 (N_9782,N_7746,N_8906);
or U9783 (N_9783,N_8969,N_7552);
and U9784 (N_9784,N_8166,N_8525);
and U9785 (N_9785,N_7717,N_8819);
and U9786 (N_9786,N_7616,N_8170);
or U9787 (N_9787,N_8987,N_8156);
or U9788 (N_9788,N_7921,N_7729);
and U9789 (N_9789,N_7877,N_8382);
and U9790 (N_9790,N_8787,N_8363);
or U9791 (N_9791,N_7982,N_8447);
and U9792 (N_9792,N_7888,N_7815);
nor U9793 (N_9793,N_8075,N_8220);
or U9794 (N_9794,N_7674,N_8826);
and U9795 (N_9795,N_8539,N_8097);
or U9796 (N_9796,N_7534,N_8017);
xnor U9797 (N_9797,N_8995,N_8386);
nor U9798 (N_9798,N_8283,N_8373);
xnor U9799 (N_9799,N_8397,N_7597);
nor U9800 (N_9800,N_8724,N_8288);
and U9801 (N_9801,N_8598,N_8411);
nor U9802 (N_9802,N_7779,N_8124);
nand U9803 (N_9803,N_8028,N_8237);
nor U9804 (N_9804,N_8635,N_7796);
and U9805 (N_9805,N_7666,N_7727);
xor U9806 (N_9806,N_8036,N_7797);
and U9807 (N_9807,N_7586,N_8472);
or U9808 (N_9808,N_8919,N_7531);
xnor U9809 (N_9809,N_8276,N_8800);
xor U9810 (N_9810,N_8844,N_7555);
nand U9811 (N_9811,N_8371,N_7500);
nand U9812 (N_9812,N_7560,N_8604);
and U9813 (N_9813,N_8239,N_8280);
nor U9814 (N_9814,N_8526,N_7734);
nand U9815 (N_9815,N_8249,N_8839);
xor U9816 (N_9816,N_7739,N_7644);
nor U9817 (N_9817,N_8448,N_7820);
or U9818 (N_9818,N_8702,N_8909);
nand U9819 (N_9819,N_8345,N_7591);
xnor U9820 (N_9820,N_7870,N_7772);
nand U9821 (N_9821,N_7608,N_8065);
nand U9822 (N_9822,N_7832,N_7687);
xor U9823 (N_9823,N_7638,N_8225);
or U9824 (N_9824,N_8604,N_8085);
and U9825 (N_9825,N_7539,N_7921);
or U9826 (N_9826,N_8112,N_8547);
or U9827 (N_9827,N_7792,N_8878);
or U9828 (N_9828,N_8494,N_7765);
nor U9829 (N_9829,N_8567,N_7733);
nand U9830 (N_9830,N_7575,N_8644);
or U9831 (N_9831,N_8418,N_8979);
nand U9832 (N_9832,N_8653,N_7882);
nor U9833 (N_9833,N_7500,N_8534);
and U9834 (N_9834,N_8809,N_7616);
nand U9835 (N_9835,N_8330,N_8126);
nand U9836 (N_9836,N_7986,N_8092);
or U9837 (N_9837,N_8352,N_8936);
nand U9838 (N_9838,N_8281,N_8154);
and U9839 (N_9839,N_7525,N_8381);
xnor U9840 (N_9840,N_7532,N_8999);
and U9841 (N_9841,N_7622,N_8682);
nand U9842 (N_9842,N_7668,N_7607);
and U9843 (N_9843,N_7933,N_8378);
or U9844 (N_9844,N_8232,N_8823);
and U9845 (N_9845,N_8079,N_8387);
nor U9846 (N_9846,N_8333,N_8202);
xor U9847 (N_9847,N_7933,N_7728);
nor U9848 (N_9848,N_7848,N_8538);
and U9849 (N_9849,N_7568,N_8001);
or U9850 (N_9850,N_7850,N_7789);
xor U9851 (N_9851,N_8130,N_8949);
xor U9852 (N_9852,N_8718,N_8027);
xnor U9853 (N_9853,N_8033,N_7960);
xor U9854 (N_9854,N_8676,N_8821);
or U9855 (N_9855,N_8074,N_8926);
nand U9856 (N_9856,N_7921,N_7944);
and U9857 (N_9857,N_8062,N_7927);
nand U9858 (N_9858,N_8446,N_8324);
nor U9859 (N_9859,N_8190,N_7860);
nand U9860 (N_9860,N_7608,N_8494);
or U9861 (N_9861,N_7652,N_7741);
and U9862 (N_9862,N_8342,N_7765);
xnor U9863 (N_9863,N_8398,N_8686);
and U9864 (N_9864,N_8667,N_7566);
xor U9865 (N_9865,N_7635,N_8646);
xnor U9866 (N_9866,N_8136,N_8684);
and U9867 (N_9867,N_8074,N_8233);
nand U9868 (N_9868,N_7698,N_7995);
nor U9869 (N_9869,N_8993,N_7614);
nand U9870 (N_9870,N_8041,N_8411);
or U9871 (N_9871,N_7671,N_8521);
and U9872 (N_9872,N_8671,N_8894);
nand U9873 (N_9873,N_8256,N_8263);
xor U9874 (N_9874,N_8388,N_7955);
nor U9875 (N_9875,N_8559,N_8379);
nor U9876 (N_9876,N_8689,N_7993);
nand U9877 (N_9877,N_8130,N_8720);
nor U9878 (N_9878,N_8969,N_8168);
or U9879 (N_9879,N_8679,N_8407);
or U9880 (N_9880,N_8296,N_8018);
and U9881 (N_9881,N_8995,N_8037);
nor U9882 (N_9882,N_8185,N_8910);
nor U9883 (N_9883,N_8693,N_8539);
or U9884 (N_9884,N_8464,N_8241);
or U9885 (N_9885,N_8663,N_8315);
nand U9886 (N_9886,N_8605,N_8681);
or U9887 (N_9887,N_8986,N_8174);
or U9888 (N_9888,N_8719,N_7944);
nand U9889 (N_9889,N_8912,N_8907);
nor U9890 (N_9890,N_8319,N_7678);
xor U9891 (N_9891,N_7985,N_8302);
nor U9892 (N_9892,N_8605,N_7594);
or U9893 (N_9893,N_7608,N_7596);
or U9894 (N_9894,N_8701,N_7628);
nand U9895 (N_9895,N_8387,N_8094);
and U9896 (N_9896,N_7964,N_8346);
nor U9897 (N_9897,N_8697,N_7695);
nand U9898 (N_9898,N_8361,N_8176);
nor U9899 (N_9899,N_8109,N_8128);
xor U9900 (N_9900,N_7938,N_7855);
xor U9901 (N_9901,N_7788,N_7659);
xnor U9902 (N_9902,N_8082,N_8786);
nor U9903 (N_9903,N_8700,N_7548);
and U9904 (N_9904,N_8997,N_7629);
or U9905 (N_9905,N_8315,N_8458);
or U9906 (N_9906,N_7896,N_7647);
nor U9907 (N_9907,N_7843,N_8305);
nand U9908 (N_9908,N_8862,N_8812);
nand U9909 (N_9909,N_8945,N_7841);
or U9910 (N_9910,N_8955,N_7996);
or U9911 (N_9911,N_8256,N_7697);
xnor U9912 (N_9912,N_8052,N_8917);
and U9913 (N_9913,N_8642,N_8262);
nor U9914 (N_9914,N_8628,N_7516);
and U9915 (N_9915,N_8239,N_7552);
nand U9916 (N_9916,N_8986,N_7627);
xnor U9917 (N_9917,N_7606,N_8674);
nand U9918 (N_9918,N_8313,N_8604);
nor U9919 (N_9919,N_8517,N_8643);
and U9920 (N_9920,N_7966,N_8000);
or U9921 (N_9921,N_8729,N_8066);
nand U9922 (N_9922,N_8675,N_8976);
nand U9923 (N_9923,N_8542,N_8765);
and U9924 (N_9924,N_8300,N_8695);
or U9925 (N_9925,N_7766,N_8409);
nor U9926 (N_9926,N_8620,N_7972);
nor U9927 (N_9927,N_8140,N_8148);
nor U9928 (N_9928,N_7990,N_8186);
xor U9929 (N_9929,N_7583,N_8534);
nand U9930 (N_9930,N_7778,N_8467);
or U9931 (N_9931,N_7966,N_8577);
nor U9932 (N_9932,N_8802,N_8040);
nor U9933 (N_9933,N_7739,N_8680);
nand U9934 (N_9934,N_8119,N_8433);
or U9935 (N_9935,N_8696,N_8954);
or U9936 (N_9936,N_8540,N_8181);
or U9937 (N_9937,N_7709,N_7922);
or U9938 (N_9938,N_7830,N_8938);
nand U9939 (N_9939,N_8963,N_8061);
xnor U9940 (N_9940,N_7832,N_8959);
xor U9941 (N_9941,N_8800,N_8374);
nand U9942 (N_9942,N_8011,N_8280);
nand U9943 (N_9943,N_8891,N_7693);
or U9944 (N_9944,N_7595,N_8749);
nor U9945 (N_9945,N_7875,N_7577);
xnor U9946 (N_9946,N_7671,N_7708);
xor U9947 (N_9947,N_7672,N_7664);
nor U9948 (N_9948,N_7823,N_8955);
or U9949 (N_9949,N_7516,N_7783);
nor U9950 (N_9950,N_8940,N_7766);
and U9951 (N_9951,N_8727,N_8265);
or U9952 (N_9952,N_8836,N_8212);
xor U9953 (N_9953,N_8364,N_8865);
and U9954 (N_9954,N_8877,N_8265);
nand U9955 (N_9955,N_7736,N_8410);
or U9956 (N_9956,N_8142,N_8025);
and U9957 (N_9957,N_8128,N_7941);
xor U9958 (N_9958,N_7684,N_7880);
and U9959 (N_9959,N_8921,N_8022);
xnor U9960 (N_9960,N_7883,N_8280);
and U9961 (N_9961,N_8431,N_8809);
nand U9962 (N_9962,N_8667,N_8060);
nand U9963 (N_9963,N_7803,N_8339);
or U9964 (N_9964,N_8163,N_8710);
and U9965 (N_9965,N_8356,N_8800);
or U9966 (N_9966,N_8948,N_8590);
and U9967 (N_9967,N_8178,N_8466);
xor U9968 (N_9968,N_7711,N_7970);
or U9969 (N_9969,N_7601,N_7783);
nand U9970 (N_9970,N_8013,N_8011);
and U9971 (N_9971,N_8756,N_8969);
xor U9972 (N_9972,N_8538,N_7961);
or U9973 (N_9973,N_8880,N_8162);
and U9974 (N_9974,N_8925,N_8899);
nand U9975 (N_9975,N_7673,N_7882);
or U9976 (N_9976,N_7841,N_7684);
nor U9977 (N_9977,N_7865,N_7588);
and U9978 (N_9978,N_8323,N_8811);
nand U9979 (N_9979,N_7846,N_7556);
nand U9980 (N_9980,N_8792,N_8421);
nor U9981 (N_9981,N_8428,N_8871);
nand U9982 (N_9982,N_8464,N_8670);
nor U9983 (N_9983,N_7717,N_8972);
or U9984 (N_9984,N_8824,N_8528);
xor U9985 (N_9985,N_8281,N_8449);
and U9986 (N_9986,N_8464,N_7689);
or U9987 (N_9987,N_8037,N_8695);
xor U9988 (N_9988,N_7641,N_8586);
or U9989 (N_9989,N_7715,N_8339);
nor U9990 (N_9990,N_7520,N_8244);
or U9991 (N_9991,N_8231,N_8131);
xnor U9992 (N_9992,N_8482,N_8159);
and U9993 (N_9993,N_8662,N_8220);
and U9994 (N_9994,N_7718,N_8540);
and U9995 (N_9995,N_8663,N_8787);
xor U9996 (N_9996,N_8455,N_8424);
nand U9997 (N_9997,N_8729,N_8768);
nor U9998 (N_9998,N_7826,N_8068);
nand U9999 (N_9999,N_8065,N_8124);
nor U10000 (N_10000,N_8297,N_8744);
or U10001 (N_10001,N_8933,N_8180);
nand U10002 (N_10002,N_8083,N_7530);
nor U10003 (N_10003,N_8831,N_8745);
nor U10004 (N_10004,N_8106,N_7834);
nor U10005 (N_10005,N_8278,N_8645);
and U10006 (N_10006,N_8360,N_8277);
or U10007 (N_10007,N_8851,N_8428);
or U10008 (N_10008,N_8037,N_8314);
or U10009 (N_10009,N_7960,N_8634);
and U10010 (N_10010,N_8772,N_8943);
and U10011 (N_10011,N_7953,N_7752);
nor U10012 (N_10012,N_7646,N_8669);
or U10013 (N_10013,N_8431,N_8014);
and U10014 (N_10014,N_8106,N_7545);
or U10015 (N_10015,N_8465,N_8207);
nand U10016 (N_10016,N_8494,N_8217);
nor U10017 (N_10017,N_7639,N_8574);
and U10018 (N_10018,N_8245,N_8068);
nor U10019 (N_10019,N_8324,N_7684);
or U10020 (N_10020,N_8529,N_7827);
and U10021 (N_10021,N_8227,N_8650);
nand U10022 (N_10022,N_8434,N_7894);
or U10023 (N_10023,N_7717,N_8864);
nor U10024 (N_10024,N_8239,N_7557);
nand U10025 (N_10025,N_8054,N_8698);
nand U10026 (N_10026,N_7658,N_8292);
xor U10027 (N_10027,N_7994,N_8035);
or U10028 (N_10028,N_8584,N_7560);
and U10029 (N_10029,N_7714,N_8521);
nor U10030 (N_10030,N_8822,N_8515);
xnor U10031 (N_10031,N_8107,N_7993);
xnor U10032 (N_10032,N_8346,N_8734);
nor U10033 (N_10033,N_8603,N_8373);
or U10034 (N_10034,N_8307,N_8088);
xnor U10035 (N_10035,N_8611,N_7818);
nor U10036 (N_10036,N_8424,N_8315);
and U10037 (N_10037,N_8151,N_7714);
or U10038 (N_10038,N_8225,N_8662);
and U10039 (N_10039,N_8010,N_8538);
xor U10040 (N_10040,N_8321,N_8824);
and U10041 (N_10041,N_7515,N_8920);
xor U10042 (N_10042,N_8195,N_8858);
xnor U10043 (N_10043,N_8514,N_8046);
nor U10044 (N_10044,N_8908,N_8394);
xor U10045 (N_10045,N_8814,N_8028);
and U10046 (N_10046,N_8650,N_8095);
xnor U10047 (N_10047,N_8529,N_8661);
and U10048 (N_10048,N_8388,N_8596);
or U10049 (N_10049,N_8492,N_8704);
nand U10050 (N_10050,N_8352,N_8120);
or U10051 (N_10051,N_7843,N_7619);
or U10052 (N_10052,N_8128,N_8506);
nor U10053 (N_10053,N_8848,N_7897);
nand U10054 (N_10054,N_8418,N_8538);
and U10055 (N_10055,N_8294,N_8121);
and U10056 (N_10056,N_8771,N_8117);
xor U10057 (N_10057,N_8552,N_8914);
and U10058 (N_10058,N_8797,N_8569);
or U10059 (N_10059,N_8228,N_7972);
and U10060 (N_10060,N_8111,N_8921);
or U10061 (N_10061,N_7761,N_7684);
nand U10062 (N_10062,N_8997,N_8785);
nor U10063 (N_10063,N_8264,N_8845);
nor U10064 (N_10064,N_8810,N_8329);
nand U10065 (N_10065,N_8058,N_8806);
xnor U10066 (N_10066,N_8743,N_8903);
nand U10067 (N_10067,N_7812,N_8908);
or U10068 (N_10068,N_8148,N_8426);
or U10069 (N_10069,N_8763,N_8152);
and U10070 (N_10070,N_7799,N_8206);
or U10071 (N_10071,N_7521,N_7579);
or U10072 (N_10072,N_8305,N_7766);
or U10073 (N_10073,N_8727,N_8722);
nor U10074 (N_10074,N_8457,N_7683);
or U10075 (N_10075,N_8909,N_8395);
and U10076 (N_10076,N_8542,N_8792);
xor U10077 (N_10077,N_8526,N_7752);
nor U10078 (N_10078,N_7858,N_7838);
nand U10079 (N_10079,N_7527,N_8137);
nor U10080 (N_10080,N_8666,N_8763);
or U10081 (N_10081,N_8919,N_7581);
or U10082 (N_10082,N_8601,N_8697);
xnor U10083 (N_10083,N_8310,N_8738);
nor U10084 (N_10084,N_8484,N_8695);
nand U10085 (N_10085,N_8543,N_7722);
or U10086 (N_10086,N_8084,N_8851);
nor U10087 (N_10087,N_8436,N_8294);
or U10088 (N_10088,N_8280,N_7939);
or U10089 (N_10089,N_8305,N_8219);
and U10090 (N_10090,N_7767,N_7836);
or U10091 (N_10091,N_7913,N_8558);
and U10092 (N_10092,N_7689,N_8630);
nor U10093 (N_10093,N_7957,N_8690);
xor U10094 (N_10094,N_8597,N_8556);
or U10095 (N_10095,N_8932,N_8352);
and U10096 (N_10096,N_8196,N_8607);
or U10097 (N_10097,N_8610,N_8902);
or U10098 (N_10098,N_8437,N_8406);
nor U10099 (N_10099,N_8696,N_8334);
nand U10100 (N_10100,N_8656,N_7749);
or U10101 (N_10101,N_8899,N_7728);
nor U10102 (N_10102,N_8117,N_8467);
or U10103 (N_10103,N_7801,N_7694);
or U10104 (N_10104,N_8440,N_7590);
nand U10105 (N_10105,N_8386,N_8223);
xnor U10106 (N_10106,N_8466,N_8298);
xor U10107 (N_10107,N_7860,N_8571);
and U10108 (N_10108,N_7881,N_8728);
nand U10109 (N_10109,N_7750,N_8233);
nor U10110 (N_10110,N_8161,N_8792);
or U10111 (N_10111,N_8084,N_7925);
or U10112 (N_10112,N_8922,N_7722);
or U10113 (N_10113,N_8042,N_8117);
and U10114 (N_10114,N_7665,N_7703);
xor U10115 (N_10115,N_7513,N_8822);
xor U10116 (N_10116,N_8644,N_7522);
or U10117 (N_10117,N_8871,N_7733);
nand U10118 (N_10118,N_7667,N_8151);
xor U10119 (N_10119,N_8310,N_8984);
and U10120 (N_10120,N_7784,N_7974);
and U10121 (N_10121,N_7734,N_8485);
and U10122 (N_10122,N_8771,N_8883);
or U10123 (N_10123,N_8971,N_8520);
or U10124 (N_10124,N_8804,N_8039);
or U10125 (N_10125,N_7652,N_8755);
nand U10126 (N_10126,N_8507,N_7945);
nor U10127 (N_10127,N_8665,N_8873);
nand U10128 (N_10128,N_8679,N_8020);
nand U10129 (N_10129,N_8400,N_7734);
nand U10130 (N_10130,N_8538,N_8303);
nand U10131 (N_10131,N_8068,N_8162);
xnor U10132 (N_10132,N_8555,N_8757);
nor U10133 (N_10133,N_8801,N_8438);
or U10134 (N_10134,N_8889,N_8328);
and U10135 (N_10135,N_8114,N_7937);
and U10136 (N_10136,N_8803,N_8919);
xor U10137 (N_10137,N_8710,N_8770);
xnor U10138 (N_10138,N_8206,N_8169);
nor U10139 (N_10139,N_8809,N_8153);
nand U10140 (N_10140,N_8922,N_8995);
nand U10141 (N_10141,N_7702,N_7859);
nor U10142 (N_10142,N_7975,N_7572);
and U10143 (N_10143,N_7646,N_8133);
xnor U10144 (N_10144,N_8023,N_8936);
or U10145 (N_10145,N_8002,N_8120);
xnor U10146 (N_10146,N_7604,N_8556);
and U10147 (N_10147,N_8641,N_8755);
nor U10148 (N_10148,N_7508,N_7953);
xnor U10149 (N_10149,N_8291,N_8086);
xor U10150 (N_10150,N_8876,N_7547);
nand U10151 (N_10151,N_7569,N_8963);
or U10152 (N_10152,N_8894,N_8389);
and U10153 (N_10153,N_7918,N_8903);
and U10154 (N_10154,N_8410,N_8002);
and U10155 (N_10155,N_7572,N_8840);
nand U10156 (N_10156,N_8121,N_8462);
or U10157 (N_10157,N_8938,N_8530);
and U10158 (N_10158,N_8268,N_8587);
nand U10159 (N_10159,N_7906,N_8147);
nand U10160 (N_10160,N_7909,N_8592);
and U10161 (N_10161,N_8539,N_8978);
nor U10162 (N_10162,N_8034,N_7605);
xor U10163 (N_10163,N_8152,N_8644);
or U10164 (N_10164,N_8632,N_8629);
nand U10165 (N_10165,N_8645,N_7533);
or U10166 (N_10166,N_7947,N_8793);
and U10167 (N_10167,N_8861,N_8170);
or U10168 (N_10168,N_8607,N_8292);
nand U10169 (N_10169,N_8119,N_7724);
and U10170 (N_10170,N_7701,N_8258);
xor U10171 (N_10171,N_8280,N_7526);
nor U10172 (N_10172,N_8286,N_8956);
xor U10173 (N_10173,N_8813,N_8207);
nor U10174 (N_10174,N_8868,N_8450);
and U10175 (N_10175,N_8337,N_8327);
and U10176 (N_10176,N_8934,N_8664);
or U10177 (N_10177,N_8381,N_8190);
nor U10178 (N_10178,N_8126,N_8674);
or U10179 (N_10179,N_8052,N_8806);
nor U10180 (N_10180,N_8793,N_8468);
nor U10181 (N_10181,N_8647,N_8736);
or U10182 (N_10182,N_8664,N_8016);
nand U10183 (N_10183,N_7570,N_8001);
or U10184 (N_10184,N_7584,N_8692);
nand U10185 (N_10185,N_8007,N_7980);
nand U10186 (N_10186,N_8039,N_8857);
nand U10187 (N_10187,N_7681,N_7850);
or U10188 (N_10188,N_8555,N_7789);
nor U10189 (N_10189,N_7991,N_8569);
xnor U10190 (N_10190,N_8238,N_8293);
or U10191 (N_10191,N_7997,N_7561);
xor U10192 (N_10192,N_7836,N_8362);
or U10193 (N_10193,N_8172,N_7854);
and U10194 (N_10194,N_8639,N_8716);
nand U10195 (N_10195,N_8289,N_8526);
nand U10196 (N_10196,N_7891,N_7969);
xor U10197 (N_10197,N_8715,N_7874);
nor U10198 (N_10198,N_8339,N_8529);
nand U10199 (N_10199,N_8554,N_8527);
xnor U10200 (N_10200,N_8927,N_8646);
xnor U10201 (N_10201,N_7693,N_8342);
and U10202 (N_10202,N_8036,N_8204);
and U10203 (N_10203,N_7914,N_8512);
and U10204 (N_10204,N_7739,N_8804);
and U10205 (N_10205,N_8753,N_8398);
nor U10206 (N_10206,N_8427,N_8073);
or U10207 (N_10207,N_8455,N_7814);
nor U10208 (N_10208,N_8233,N_8661);
nor U10209 (N_10209,N_7992,N_8467);
and U10210 (N_10210,N_7905,N_7533);
nor U10211 (N_10211,N_8602,N_7546);
nor U10212 (N_10212,N_8216,N_7796);
nor U10213 (N_10213,N_7809,N_8732);
or U10214 (N_10214,N_8916,N_7734);
xnor U10215 (N_10215,N_7951,N_7818);
or U10216 (N_10216,N_8407,N_8813);
nand U10217 (N_10217,N_8575,N_8470);
xor U10218 (N_10218,N_8058,N_8142);
nor U10219 (N_10219,N_8254,N_8408);
or U10220 (N_10220,N_7669,N_7887);
and U10221 (N_10221,N_8008,N_7548);
nand U10222 (N_10222,N_8274,N_7712);
xor U10223 (N_10223,N_7623,N_8231);
nand U10224 (N_10224,N_8712,N_7847);
nand U10225 (N_10225,N_8460,N_7588);
xor U10226 (N_10226,N_8818,N_8697);
nand U10227 (N_10227,N_7697,N_7698);
nor U10228 (N_10228,N_7835,N_8537);
nand U10229 (N_10229,N_8727,N_8928);
nor U10230 (N_10230,N_8637,N_8936);
xnor U10231 (N_10231,N_7766,N_7991);
nor U10232 (N_10232,N_7652,N_7906);
or U10233 (N_10233,N_8440,N_8633);
nand U10234 (N_10234,N_8322,N_8673);
xor U10235 (N_10235,N_8946,N_7569);
nand U10236 (N_10236,N_8159,N_8071);
nand U10237 (N_10237,N_7937,N_8502);
nand U10238 (N_10238,N_8360,N_7720);
or U10239 (N_10239,N_8320,N_8598);
nor U10240 (N_10240,N_8500,N_8977);
xor U10241 (N_10241,N_7851,N_8122);
and U10242 (N_10242,N_8894,N_8060);
nor U10243 (N_10243,N_8666,N_7656);
and U10244 (N_10244,N_7898,N_7738);
or U10245 (N_10245,N_8564,N_8880);
nor U10246 (N_10246,N_8352,N_8559);
and U10247 (N_10247,N_8712,N_8311);
or U10248 (N_10248,N_8768,N_7881);
xor U10249 (N_10249,N_8102,N_8103);
and U10250 (N_10250,N_8260,N_8184);
and U10251 (N_10251,N_8377,N_8983);
or U10252 (N_10252,N_7700,N_8635);
and U10253 (N_10253,N_7634,N_8328);
nand U10254 (N_10254,N_7760,N_7530);
and U10255 (N_10255,N_8483,N_8587);
xnor U10256 (N_10256,N_8377,N_7675);
nand U10257 (N_10257,N_8832,N_8011);
and U10258 (N_10258,N_8072,N_8025);
nor U10259 (N_10259,N_8452,N_8701);
and U10260 (N_10260,N_8731,N_8630);
xor U10261 (N_10261,N_7928,N_7788);
nor U10262 (N_10262,N_7540,N_8869);
or U10263 (N_10263,N_7647,N_8191);
xnor U10264 (N_10264,N_8654,N_7558);
and U10265 (N_10265,N_8381,N_8348);
nand U10266 (N_10266,N_8072,N_8716);
or U10267 (N_10267,N_7744,N_8712);
nand U10268 (N_10268,N_7931,N_8817);
or U10269 (N_10269,N_7646,N_8423);
nand U10270 (N_10270,N_8522,N_7677);
and U10271 (N_10271,N_8157,N_8453);
or U10272 (N_10272,N_8946,N_7830);
nand U10273 (N_10273,N_8681,N_8330);
xnor U10274 (N_10274,N_8341,N_7717);
nand U10275 (N_10275,N_7695,N_8014);
nand U10276 (N_10276,N_8318,N_8134);
nor U10277 (N_10277,N_8819,N_8942);
and U10278 (N_10278,N_7663,N_8206);
or U10279 (N_10279,N_8086,N_8743);
nand U10280 (N_10280,N_7701,N_8534);
nand U10281 (N_10281,N_7525,N_8686);
or U10282 (N_10282,N_8015,N_8591);
and U10283 (N_10283,N_7623,N_8931);
or U10284 (N_10284,N_8714,N_7716);
xor U10285 (N_10285,N_8891,N_8184);
nand U10286 (N_10286,N_8364,N_8040);
nand U10287 (N_10287,N_8039,N_7628);
nor U10288 (N_10288,N_8685,N_8929);
or U10289 (N_10289,N_8727,N_7864);
xor U10290 (N_10290,N_8025,N_7935);
nand U10291 (N_10291,N_7525,N_7884);
or U10292 (N_10292,N_8412,N_7894);
or U10293 (N_10293,N_8449,N_8912);
nand U10294 (N_10294,N_8143,N_8461);
nor U10295 (N_10295,N_8940,N_8991);
nand U10296 (N_10296,N_8707,N_8603);
nand U10297 (N_10297,N_8046,N_7945);
xnor U10298 (N_10298,N_7675,N_8614);
xor U10299 (N_10299,N_8936,N_8953);
or U10300 (N_10300,N_7878,N_8221);
or U10301 (N_10301,N_7814,N_8044);
xor U10302 (N_10302,N_8292,N_8324);
xor U10303 (N_10303,N_8544,N_7945);
and U10304 (N_10304,N_7780,N_8679);
and U10305 (N_10305,N_8654,N_8730);
xnor U10306 (N_10306,N_8291,N_7551);
xor U10307 (N_10307,N_7714,N_8306);
xor U10308 (N_10308,N_8463,N_7573);
or U10309 (N_10309,N_7587,N_7997);
or U10310 (N_10310,N_7708,N_8456);
and U10311 (N_10311,N_8241,N_8872);
and U10312 (N_10312,N_7760,N_7667);
or U10313 (N_10313,N_8751,N_8122);
xor U10314 (N_10314,N_8526,N_8211);
nor U10315 (N_10315,N_8293,N_8674);
nor U10316 (N_10316,N_8342,N_8935);
nand U10317 (N_10317,N_7618,N_8447);
or U10318 (N_10318,N_7708,N_8088);
and U10319 (N_10319,N_8797,N_8687);
nand U10320 (N_10320,N_8696,N_8628);
or U10321 (N_10321,N_8822,N_8406);
nor U10322 (N_10322,N_7619,N_8160);
nor U10323 (N_10323,N_8767,N_8054);
nand U10324 (N_10324,N_8951,N_8590);
nand U10325 (N_10325,N_8728,N_7579);
nand U10326 (N_10326,N_7984,N_8770);
nand U10327 (N_10327,N_8642,N_8749);
and U10328 (N_10328,N_7864,N_8246);
nand U10329 (N_10329,N_8595,N_8409);
nand U10330 (N_10330,N_8867,N_8116);
nor U10331 (N_10331,N_8373,N_7590);
and U10332 (N_10332,N_8785,N_8767);
and U10333 (N_10333,N_7989,N_8190);
and U10334 (N_10334,N_8283,N_8020);
xor U10335 (N_10335,N_7717,N_8806);
or U10336 (N_10336,N_8397,N_8761);
nand U10337 (N_10337,N_7860,N_8323);
nor U10338 (N_10338,N_8097,N_7560);
nor U10339 (N_10339,N_8661,N_8544);
xor U10340 (N_10340,N_7537,N_8866);
or U10341 (N_10341,N_8835,N_8236);
or U10342 (N_10342,N_7876,N_8258);
or U10343 (N_10343,N_7537,N_8431);
or U10344 (N_10344,N_8657,N_7815);
and U10345 (N_10345,N_8822,N_8607);
or U10346 (N_10346,N_8817,N_7917);
nor U10347 (N_10347,N_8892,N_7826);
nor U10348 (N_10348,N_8829,N_7564);
nor U10349 (N_10349,N_8906,N_8959);
xnor U10350 (N_10350,N_8768,N_8966);
nand U10351 (N_10351,N_8467,N_8187);
nand U10352 (N_10352,N_8325,N_8413);
nand U10353 (N_10353,N_7695,N_7892);
and U10354 (N_10354,N_8498,N_8827);
xor U10355 (N_10355,N_7756,N_7878);
nand U10356 (N_10356,N_8403,N_8469);
nand U10357 (N_10357,N_8402,N_8619);
xor U10358 (N_10358,N_7754,N_8928);
nor U10359 (N_10359,N_8293,N_8405);
nand U10360 (N_10360,N_8496,N_8386);
or U10361 (N_10361,N_7670,N_7972);
nor U10362 (N_10362,N_8686,N_7978);
nand U10363 (N_10363,N_8362,N_8555);
or U10364 (N_10364,N_8700,N_8474);
or U10365 (N_10365,N_8108,N_8258);
or U10366 (N_10366,N_8701,N_7769);
xor U10367 (N_10367,N_8791,N_7694);
nand U10368 (N_10368,N_7976,N_8510);
xor U10369 (N_10369,N_7822,N_8316);
nand U10370 (N_10370,N_7667,N_7951);
or U10371 (N_10371,N_7662,N_7726);
or U10372 (N_10372,N_7623,N_8958);
or U10373 (N_10373,N_8039,N_7977);
nand U10374 (N_10374,N_8323,N_7630);
or U10375 (N_10375,N_8946,N_7786);
xor U10376 (N_10376,N_7694,N_8667);
xor U10377 (N_10377,N_7536,N_8169);
xor U10378 (N_10378,N_7858,N_8126);
or U10379 (N_10379,N_8637,N_8530);
and U10380 (N_10380,N_8634,N_8688);
or U10381 (N_10381,N_7747,N_8883);
or U10382 (N_10382,N_8119,N_7590);
nand U10383 (N_10383,N_8225,N_7852);
xnor U10384 (N_10384,N_8042,N_8503);
or U10385 (N_10385,N_7629,N_7604);
nor U10386 (N_10386,N_8253,N_7926);
nor U10387 (N_10387,N_8509,N_8971);
nand U10388 (N_10388,N_7969,N_8095);
and U10389 (N_10389,N_8804,N_7689);
and U10390 (N_10390,N_8101,N_8683);
nor U10391 (N_10391,N_8110,N_8900);
nand U10392 (N_10392,N_8962,N_8454);
or U10393 (N_10393,N_7633,N_8395);
and U10394 (N_10394,N_7556,N_8203);
nor U10395 (N_10395,N_8831,N_8615);
xnor U10396 (N_10396,N_7526,N_8751);
nand U10397 (N_10397,N_8081,N_7957);
nor U10398 (N_10398,N_8140,N_7587);
and U10399 (N_10399,N_7800,N_8580);
nor U10400 (N_10400,N_7784,N_7801);
nor U10401 (N_10401,N_8466,N_7529);
xnor U10402 (N_10402,N_8827,N_8822);
xor U10403 (N_10403,N_8998,N_8609);
nand U10404 (N_10404,N_8271,N_7945);
nor U10405 (N_10405,N_8254,N_8193);
nand U10406 (N_10406,N_7577,N_8676);
or U10407 (N_10407,N_8519,N_8611);
and U10408 (N_10408,N_8720,N_8348);
nor U10409 (N_10409,N_8011,N_8988);
nand U10410 (N_10410,N_7614,N_7720);
xor U10411 (N_10411,N_8001,N_8473);
xnor U10412 (N_10412,N_7789,N_7798);
or U10413 (N_10413,N_8020,N_8758);
nor U10414 (N_10414,N_7657,N_8972);
or U10415 (N_10415,N_7720,N_7830);
and U10416 (N_10416,N_7663,N_8556);
or U10417 (N_10417,N_8170,N_8352);
xor U10418 (N_10418,N_8308,N_8134);
nor U10419 (N_10419,N_7775,N_8580);
nor U10420 (N_10420,N_8917,N_8837);
nand U10421 (N_10421,N_8742,N_7841);
xnor U10422 (N_10422,N_8821,N_7949);
nor U10423 (N_10423,N_8563,N_7792);
nand U10424 (N_10424,N_8622,N_8857);
nor U10425 (N_10425,N_8823,N_7615);
xor U10426 (N_10426,N_8521,N_7781);
nor U10427 (N_10427,N_8821,N_8308);
or U10428 (N_10428,N_8901,N_8628);
nand U10429 (N_10429,N_8458,N_8038);
xor U10430 (N_10430,N_8199,N_8447);
nand U10431 (N_10431,N_7673,N_8141);
xor U10432 (N_10432,N_7985,N_8286);
xor U10433 (N_10433,N_7982,N_8862);
nor U10434 (N_10434,N_7972,N_7820);
xnor U10435 (N_10435,N_8584,N_7793);
and U10436 (N_10436,N_8779,N_7672);
and U10437 (N_10437,N_8374,N_8002);
or U10438 (N_10438,N_7818,N_8105);
nand U10439 (N_10439,N_8750,N_7925);
or U10440 (N_10440,N_8277,N_8045);
and U10441 (N_10441,N_7542,N_7671);
xor U10442 (N_10442,N_8932,N_8172);
nor U10443 (N_10443,N_8960,N_8553);
or U10444 (N_10444,N_8850,N_8263);
xnor U10445 (N_10445,N_8723,N_8014);
nor U10446 (N_10446,N_8098,N_7963);
nand U10447 (N_10447,N_8216,N_7723);
and U10448 (N_10448,N_7899,N_8383);
nor U10449 (N_10449,N_8284,N_8056);
or U10450 (N_10450,N_8214,N_8022);
or U10451 (N_10451,N_8298,N_7668);
or U10452 (N_10452,N_8224,N_7913);
xor U10453 (N_10453,N_8750,N_7590);
nor U10454 (N_10454,N_7500,N_8219);
and U10455 (N_10455,N_8448,N_7985);
or U10456 (N_10456,N_8298,N_7777);
xnor U10457 (N_10457,N_8200,N_7847);
nand U10458 (N_10458,N_8493,N_7500);
or U10459 (N_10459,N_8906,N_8558);
nand U10460 (N_10460,N_8173,N_7991);
nand U10461 (N_10461,N_8427,N_8148);
xor U10462 (N_10462,N_8527,N_8730);
or U10463 (N_10463,N_8904,N_7590);
nand U10464 (N_10464,N_8452,N_8037);
and U10465 (N_10465,N_8393,N_7869);
or U10466 (N_10466,N_8857,N_7596);
nand U10467 (N_10467,N_8971,N_8569);
or U10468 (N_10468,N_7801,N_8820);
nand U10469 (N_10469,N_7789,N_8903);
xor U10470 (N_10470,N_8342,N_8911);
nor U10471 (N_10471,N_7699,N_7868);
xnor U10472 (N_10472,N_8876,N_7638);
nor U10473 (N_10473,N_8073,N_7745);
or U10474 (N_10474,N_7909,N_8915);
nand U10475 (N_10475,N_8768,N_8170);
and U10476 (N_10476,N_8094,N_8014);
xnor U10477 (N_10477,N_8502,N_7679);
and U10478 (N_10478,N_7833,N_8795);
xnor U10479 (N_10479,N_8126,N_7990);
nor U10480 (N_10480,N_8042,N_8254);
xnor U10481 (N_10481,N_8018,N_8274);
xor U10482 (N_10482,N_8673,N_8257);
nor U10483 (N_10483,N_8118,N_8583);
xor U10484 (N_10484,N_8154,N_8229);
or U10485 (N_10485,N_8357,N_8424);
and U10486 (N_10486,N_8586,N_7725);
nand U10487 (N_10487,N_7716,N_8561);
nor U10488 (N_10488,N_8423,N_8733);
xnor U10489 (N_10489,N_7870,N_7800);
xor U10490 (N_10490,N_8100,N_7920);
or U10491 (N_10491,N_8802,N_7838);
or U10492 (N_10492,N_8357,N_8852);
xnor U10493 (N_10493,N_8826,N_8160);
xor U10494 (N_10494,N_8226,N_8081);
and U10495 (N_10495,N_8834,N_8240);
nor U10496 (N_10496,N_7808,N_8428);
or U10497 (N_10497,N_8089,N_8163);
xnor U10498 (N_10498,N_8674,N_8204);
and U10499 (N_10499,N_8139,N_7951);
nor U10500 (N_10500,N_9019,N_9784);
xor U10501 (N_10501,N_10091,N_10420);
and U10502 (N_10502,N_9177,N_10114);
or U10503 (N_10503,N_9059,N_9945);
and U10504 (N_10504,N_10185,N_10059);
nor U10505 (N_10505,N_10055,N_10498);
nor U10506 (N_10506,N_9874,N_9325);
nand U10507 (N_10507,N_9733,N_9852);
nor U10508 (N_10508,N_10208,N_10268);
nor U10509 (N_10509,N_10011,N_10123);
nor U10510 (N_10510,N_10269,N_9749);
and U10511 (N_10511,N_9965,N_9846);
or U10512 (N_10512,N_10166,N_9682);
nand U10513 (N_10513,N_10009,N_9831);
nand U10514 (N_10514,N_9201,N_10158);
xor U10515 (N_10515,N_10494,N_10015);
nor U10516 (N_10516,N_9514,N_10386);
or U10517 (N_10517,N_9274,N_10225);
or U10518 (N_10518,N_9227,N_9293);
or U10519 (N_10519,N_10312,N_9995);
nand U10520 (N_10520,N_10242,N_9543);
or U10521 (N_10521,N_9459,N_9480);
nor U10522 (N_10522,N_10265,N_10130);
xnor U10523 (N_10523,N_9661,N_9979);
and U10524 (N_10524,N_10263,N_9968);
xnor U10525 (N_10525,N_10186,N_9786);
nand U10526 (N_10526,N_10108,N_9599);
nor U10527 (N_10527,N_9820,N_9387);
nand U10528 (N_10528,N_9550,N_9930);
xnor U10529 (N_10529,N_9612,N_10047);
xor U10530 (N_10530,N_9693,N_9239);
and U10531 (N_10531,N_9537,N_9624);
xnor U10532 (N_10532,N_10464,N_10314);
xor U10533 (N_10533,N_10082,N_9590);
xnor U10534 (N_10534,N_9611,N_10140);
nor U10535 (N_10535,N_9845,N_9213);
nor U10536 (N_10536,N_9620,N_10323);
nand U10537 (N_10537,N_9904,N_9070);
nor U10538 (N_10538,N_10425,N_9674);
xnor U10539 (N_10539,N_9091,N_9894);
and U10540 (N_10540,N_10241,N_9681);
nor U10541 (N_10541,N_9403,N_9074);
and U10542 (N_10542,N_10345,N_10488);
nand U10543 (N_10543,N_9423,N_10448);
xor U10544 (N_10544,N_9440,N_9349);
and U10545 (N_10545,N_9408,N_9896);
or U10546 (N_10546,N_9604,N_10137);
or U10547 (N_10547,N_9708,N_10276);
nor U10548 (N_10548,N_9415,N_9526);
or U10549 (N_10549,N_10061,N_9544);
or U10550 (N_10550,N_9337,N_9909);
or U10551 (N_10551,N_9960,N_9678);
and U10552 (N_10552,N_9967,N_9504);
and U10553 (N_10553,N_10104,N_9993);
nand U10554 (N_10554,N_9384,N_10077);
xnor U10555 (N_10555,N_9574,N_9161);
and U10556 (N_10556,N_9591,N_9052);
xnor U10557 (N_10557,N_10384,N_9441);
and U10558 (N_10558,N_9969,N_9527);
nor U10559 (N_10559,N_9030,N_9252);
and U10560 (N_10560,N_10178,N_10196);
nand U10561 (N_10561,N_10167,N_10480);
nand U10562 (N_10562,N_10266,N_9169);
nor U10563 (N_10563,N_10238,N_10328);
nor U10564 (N_10564,N_10232,N_9147);
xor U10565 (N_10565,N_9367,N_10457);
or U10566 (N_10566,N_9464,N_10107);
or U10567 (N_10567,N_10446,N_9485);
xor U10568 (N_10568,N_10035,N_9889);
xor U10569 (N_10569,N_9218,N_9012);
or U10570 (N_10570,N_10002,N_9760);
nand U10571 (N_10571,N_10151,N_10418);
nand U10572 (N_10572,N_10252,N_10294);
and U10573 (N_10573,N_9154,N_10304);
nand U10574 (N_10574,N_10003,N_9949);
or U10575 (N_10575,N_10333,N_9915);
and U10576 (N_10576,N_10400,N_9621);
or U10577 (N_10577,N_9469,N_10454);
nand U10578 (N_10578,N_9069,N_9868);
and U10579 (N_10579,N_9054,N_9882);
nand U10580 (N_10580,N_9466,N_10295);
xnor U10581 (N_10581,N_9586,N_9938);
nand U10582 (N_10582,N_9181,N_9734);
nor U10583 (N_10583,N_9880,N_9843);
xnor U10584 (N_10584,N_10024,N_10182);
or U10585 (N_10585,N_10377,N_10244);
nand U10586 (N_10586,N_10354,N_9566);
xor U10587 (N_10587,N_9520,N_10168);
nand U10588 (N_10588,N_9873,N_10470);
and U10589 (N_10589,N_10391,N_9297);
or U10590 (N_10590,N_10375,N_9515);
xnor U10591 (N_10591,N_10068,N_9008);
and U10592 (N_10592,N_10073,N_9329);
nand U10593 (N_10593,N_9572,N_9496);
or U10594 (N_10594,N_10303,N_9926);
or U10595 (N_10595,N_9862,N_9275);
or U10596 (N_10596,N_10098,N_9263);
and U10597 (N_10597,N_9972,N_10109);
xor U10598 (N_10598,N_9997,N_9007);
and U10599 (N_10599,N_10030,N_9507);
or U10600 (N_10600,N_9004,N_9602);
xnor U10601 (N_10601,N_9090,N_9769);
and U10602 (N_10602,N_9068,N_10398);
or U10603 (N_10603,N_9476,N_9001);
and U10604 (N_10604,N_10117,N_9456);
and U10605 (N_10605,N_9088,N_9197);
nand U10606 (N_10606,N_10297,N_9306);
or U10607 (N_10607,N_9848,N_9009);
nor U10608 (N_10608,N_10366,N_9037);
nand U10609 (N_10609,N_9955,N_9105);
xnor U10610 (N_10610,N_9954,N_10436);
xor U10611 (N_10611,N_10496,N_9535);
or U10612 (N_10612,N_9302,N_10143);
or U10613 (N_10613,N_9372,N_10311);
or U10614 (N_10614,N_9966,N_9639);
nand U10615 (N_10615,N_9659,N_10359);
xor U10616 (N_10616,N_9066,N_9588);
and U10617 (N_10617,N_10272,N_10084);
and U10618 (N_10618,N_9511,N_9338);
nand U10619 (N_10619,N_10210,N_9438);
nor U10620 (N_10620,N_9094,N_10234);
xnor U10621 (N_10621,N_9232,N_9803);
nand U10622 (N_10622,N_9101,N_9719);
or U10623 (N_10623,N_9203,N_10288);
nand U10624 (N_10624,N_10142,N_9351);
xnor U10625 (N_10625,N_9023,N_9489);
xor U10626 (N_10626,N_9772,N_9770);
nor U10627 (N_10627,N_9623,N_10067);
and U10628 (N_10628,N_9474,N_9392);
nand U10629 (N_10629,N_9864,N_10426);
and U10630 (N_10630,N_9892,N_10257);
or U10631 (N_10631,N_9911,N_9596);
and U10632 (N_10632,N_9086,N_9819);
nand U10633 (N_10633,N_9175,N_9190);
or U10634 (N_10634,N_9119,N_10414);
nor U10635 (N_10635,N_9890,N_9805);
nor U10636 (N_10636,N_10408,N_9432);
nor U10637 (N_10637,N_9249,N_9342);
xor U10638 (N_10638,N_10489,N_10412);
nor U10639 (N_10639,N_10023,N_9935);
and U10640 (N_10640,N_9560,N_10334);
nor U10641 (N_10641,N_9288,N_9794);
nand U10642 (N_10642,N_9584,N_9136);
nand U10643 (N_10643,N_9562,N_10293);
or U10644 (N_10644,N_9646,N_9667);
or U10645 (N_10645,N_9187,N_10235);
xnor U10646 (N_10646,N_10487,N_9886);
nor U10647 (N_10647,N_10099,N_9398);
xnor U10648 (N_10648,N_9461,N_9724);
xor U10649 (N_10649,N_9752,N_9345);
nand U10650 (N_10650,N_9220,N_10455);
nand U10651 (N_10651,N_9563,N_9626);
nand U10652 (N_10652,N_9625,N_9617);
or U10653 (N_10653,N_9264,N_9893);
and U10654 (N_10654,N_10152,N_9282);
and U10655 (N_10655,N_9080,N_9923);
xnor U10656 (N_10656,N_9242,N_9251);
xor U10657 (N_10657,N_9981,N_9947);
xor U10658 (N_10658,N_10236,N_9561);
xor U10659 (N_10659,N_10437,N_9108);
and U10660 (N_10660,N_9594,N_9773);
nor U10661 (N_10661,N_9900,N_9692);
or U10662 (N_10662,N_10092,N_10421);
and U10663 (N_10663,N_9310,N_9391);
nor U10664 (N_10664,N_10356,N_9268);
nand U10665 (N_10665,N_10041,N_9067);
and U10666 (N_10666,N_9823,N_9258);
or U10667 (N_10667,N_9771,N_9484);
nor U10668 (N_10668,N_9236,N_10462);
nand U10669 (N_10669,N_9179,N_9013);
or U10670 (N_10670,N_9056,N_9425);
or U10671 (N_10671,N_9097,N_10013);
and U10672 (N_10672,N_10136,N_10253);
nor U10673 (N_10673,N_10461,N_9669);
and U10674 (N_10674,N_9528,N_9478);
and U10675 (N_10675,N_9658,N_9221);
or U10676 (N_10676,N_9782,N_9357);
xor U10677 (N_10677,N_9301,N_10180);
and U10678 (N_10678,N_9278,N_9853);
or U10679 (N_10679,N_9324,N_10118);
xor U10680 (N_10680,N_10486,N_10262);
or U10681 (N_10681,N_9370,N_9641);
or U10682 (N_10682,N_10057,N_9280);
nor U10683 (N_10683,N_10207,N_10326);
or U10684 (N_10684,N_9645,N_10170);
nand U10685 (N_10685,N_9698,N_9867);
nor U10686 (N_10686,N_9437,N_9043);
and U10687 (N_10687,N_9344,N_9756);
nor U10688 (N_10688,N_9018,N_9011);
or U10689 (N_10689,N_9695,N_10231);
xnor U10690 (N_10690,N_9891,N_10138);
nor U10691 (N_10691,N_9615,N_9273);
or U10692 (N_10692,N_10267,N_9810);
and U10693 (N_10693,N_9943,N_10049);
xor U10694 (N_10694,N_9608,N_10336);
and U10695 (N_10695,N_9081,N_10441);
nand U10696 (N_10696,N_10471,N_9589);
nand U10697 (N_10697,N_10169,N_9905);
and U10698 (N_10698,N_9942,N_10435);
and U10699 (N_10699,N_10342,N_9445);
xor U10700 (N_10700,N_9106,N_10075);
nand U10701 (N_10701,N_9558,N_9534);
or U10702 (N_10702,N_9956,N_9854);
and U10703 (N_10703,N_9287,N_10282);
or U10704 (N_10704,N_10439,N_10365);
and U10705 (N_10705,N_9871,N_10032);
nor U10706 (N_10706,N_10237,N_10321);
or U10707 (N_10707,N_9200,N_10349);
and U10708 (N_10708,N_9058,N_9725);
or U10709 (N_10709,N_9498,N_10353);
and U10710 (N_10710,N_9033,N_10249);
nand U10711 (N_10711,N_10329,N_9276);
xor U10712 (N_10712,N_10051,N_9736);
and U10713 (N_10713,N_10407,N_10179);
nor U10714 (N_10714,N_9555,N_9934);
nand U10715 (N_10715,N_9903,N_9414);
xnor U10716 (N_10716,N_9679,N_9075);
or U10717 (N_10717,N_9259,N_9546);
nor U10718 (N_10718,N_9042,N_9637);
nand U10719 (N_10719,N_9257,N_9533);
and U10720 (N_10720,N_9811,N_9665);
nor U10721 (N_10721,N_9508,N_10383);
nor U10722 (N_10722,N_9493,N_9718);
and U10723 (N_10723,N_9532,N_9517);
nor U10724 (N_10724,N_10279,N_9652);
and U10725 (N_10725,N_9120,N_9036);
and U10726 (N_10726,N_10256,N_10116);
and U10727 (N_10727,N_9858,N_9285);
and U10728 (N_10728,N_10373,N_9813);
or U10729 (N_10729,N_9899,N_9283);
nand U10730 (N_10730,N_10226,N_9807);
or U10731 (N_10731,N_10331,N_10291);
or U10732 (N_10732,N_9330,N_9230);
nor U10733 (N_10733,N_9305,N_9204);
xnor U10734 (N_10734,N_10004,N_9098);
or U10735 (N_10735,N_9921,N_10451);
nand U10736 (N_10736,N_10144,N_9666);
or U10737 (N_10737,N_9341,N_10478);
and U10738 (N_10738,N_10278,N_9248);
nor U10739 (N_10739,N_9444,N_9318);
or U10740 (N_10740,N_9368,N_9542);
xor U10741 (N_10741,N_10173,N_9799);
and U10742 (N_10742,N_10103,N_9241);
and U10743 (N_10743,N_10358,N_9159);
nor U10744 (N_10744,N_9454,N_9936);
or U10745 (N_10745,N_9486,N_9928);
nand U10746 (N_10746,N_10401,N_9518);
xor U10747 (N_10747,N_10381,N_9991);
nand U10748 (N_10748,N_9835,N_10125);
and U10749 (N_10749,N_9135,N_9279);
nand U10750 (N_10750,N_10095,N_10162);
nor U10751 (N_10751,N_9226,N_9920);
xnor U10752 (N_10752,N_9578,N_9595);
xor U10753 (N_10753,N_10021,N_9790);
xnor U10754 (N_10754,N_10369,N_10285);
nor U10755 (N_10755,N_10012,N_9924);
xnor U10756 (N_10756,N_10434,N_9064);
nor U10757 (N_10757,N_10034,N_9163);
or U10758 (N_10758,N_9855,N_9312);
xor U10759 (N_10759,N_10330,N_9340);
and U10760 (N_10760,N_9460,N_10080);
and U10761 (N_10761,N_9628,N_10120);
or U10762 (N_10762,N_9818,N_9744);
nand U10763 (N_10763,N_10155,N_9700);
nand U10764 (N_10764,N_9394,N_9217);
and U10765 (N_10765,N_9609,N_9815);
and U10766 (N_10766,N_10370,N_10473);
and U10767 (N_10767,N_9360,N_9152);
xnor U10768 (N_10768,N_9869,N_9379);
nor U10769 (N_10769,N_9322,N_9291);
nor U10770 (N_10770,N_9296,N_9545);
and U10771 (N_10771,N_9806,N_9730);
and U10772 (N_10772,N_10133,N_10467);
xnor U10773 (N_10773,N_9980,N_9026);
or U10774 (N_10774,N_9465,N_10281);
xor U10775 (N_10775,N_9919,N_9839);
nor U10776 (N_10776,N_9950,N_9601);
xor U10777 (N_10777,N_10110,N_9999);
or U10778 (N_10778,N_10205,N_10469);
xor U10779 (N_10779,N_10154,N_9684);
or U10780 (N_10780,N_10485,N_10203);
nand U10781 (N_10781,N_9475,N_9082);
xor U10782 (N_10782,N_9856,N_10124);
nand U10783 (N_10783,N_9549,N_9798);
and U10784 (N_10784,N_9737,N_9613);
or U10785 (N_10785,N_9706,N_10450);
xnor U10786 (N_10786,N_9976,N_9582);
nor U10787 (N_10787,N_9103,N_10147);
nor U10788 (N_10788,N_9047,N_9577);
xnor U10789 (N_10789,N_9717,N_10122);
or U10790 (N_10790,N_9401,N_9153);
nor U10791 (N_10791,N_9024,N_10191);
or U10792 (N_10792,N_10399,N_10044);
nor U10793 (N_10793,N_9606,N_9580);
or U10794 (N_10794,N_9100,N_10490);
or U10795 (N_10795,N_10102,N_9359);
or U10796 (N_10796,N_9450,N_9878);
or U10797 (N_10797,N_9307,N_9078);
xor U10798 (N_10798,N_10352,N_9974);
nand U10799 (N_10799,N_9126,N_10033);
nor U10800 (N_10800,N_9184,N_9172);
or U10801 (N_10801,N_9162,N_9751);
nand U10802 (N_10802,N_9512,N_9160);
xnor U10803 (N_10803,N_10146,N_9038);
xnor U10804 (N_10804,N_9850,N_9132);
or U10805 (N_10805,N_9110,N_10322);
nor U10806 (N_10806,N_9509,N_9714);
nand U10807 (N_10807,N_9761,N_10442);
and U10808 (N_10808,N_9783,N_9716);
and U10809 (N_10809,N_9238,N_9683);
nand U10810 (N_10810,N_9523,N_10097);
or U10811 (N_10811,N_9188,N_9376);
and U10812 (N_10812,N_9115,N_10230);
and U10813 (N_10813,N_9944,N_9795);
nand U10814 (N_10814,N_9836,N_9709);
or U10815 (N_10815,N_9468,N_10199);
xnor U10816 (N_10816,N_9849,N_10335);
nand U10817 (N_10817,N_9910,N_10223);
and U10818 (N_10818,N_10422,N_9726);
or U10819 (N_10819,N_10112,N_9364);
xor U10820 (N_10820,N_9842,N_9421);
nand U10821 (N_10821,N_9431,N_9198);
nor U10822 (N_10822,N_10211,N_10376);
and U10823 (N_10823,N_10126,N_9859);
nand U10824 (N_10824,N_9299,N_9035);
nand U10825 (N_10825,N_9743,N_9722);
or U10826 (N_10826,N_10209,N_9568);
and U10827 (N_10827,N_9888,N_9530);
nor U10828 (N_10828,N_9347,N_10299);
or U10829 (N_10829,N_10395,N_10064);
nand U10830 (N_10830,N_10096,N_9045);
nand U10831 (N_10831,N_10479,N_10460);
or U10832 (N_10832,N_10119,N_10465);
nand U10833 (N_10833,N_10001,N_10348);
and U10834 (N_10834,N_9791,N_10387);
and U10835 (N_10835,N_9671,N_9490);
xor U10836 (N_10836,N_9458,N_9155);
nor U10837 (N_10837,N_9605,N_10048);
or U10838 (N_10838,N_9128,N_10309);
nor U10839 (N_10839,N_10008,N_10433);
and U10840 (N_10840,N_10074,N_10066);
and U10841 (N_10841,N_10200,N_10043);
xor U10842 (N_10842,N_10415,N_9146);
nor U10843 (N_10843,N_9107,N_9304);
nand U10844 (N_10844,N_9348,N_9978);
nand U10845 (N_10845,N_9907,N_10127);
and U10846 (N_10846,N_9118,N_10357);
xnor U10847 (N_10847,N_9261,N_9863);
nor U10848 (N_10848,N_9233,N_9000);
nand U10849 (N_10849,N_10307,N_9313);
nand U10850 (N_10850,N_9173,N_10087);
nor U10851 (N_10851,N_10393,N_9696);
and U10852 (N_10852,N_9483,N_10315);
nor U10853 (N_10853,N_10324,N_10429);
xor U10854 (N_10854,N_9961,N_9127);
nand U10855 (N_10855,N_9303,N_9990);
or U10856 (N_10856,N_9383,N_9689);
nor U10857 (N_10857,N_9122,N_10083);
and U10858 (N_10858,N_9102,N_9959);
nor U10859 (N_10859,N_10411,N_9397);
or U10860 (N_10860,N_9284,N_9985);
nand U10861 (N_10861,N_9071,N_10484);
nor U10862 (N_10862,N_9247,N_9872);
xor U10863 (N_10863,N_10258,N_9206);
and U10864 (N_10864,N_10456,N_9228);
xnor U10865 (N_10865,N_10385,N_9657);
or U10866 (N_10866,N_10388,N_10089);
nand U10867 (N_10867,N_10476,N_9185);
or U10868 (N_10868,N_9446,N_9319);
xnor U10869 (N_10869,N_10273,N_10183);
and U10870 (N_10870,N_9673,N_9662);
and U10871 (N_10871,N_9723,N_9089);
nor U10872 (N_10872,N_10344,N_9130);
xnor U10873 (N_10873,N_9426,N_9627);
and U10874 (N_10874,N_9254,N_10174);
and U10875 (N_10875,N_9352,N_9632);
nor U10876 (N_10876,N_9448,N_10343);
and U10877 (N_10877,N_9525,N_9655);
or U10878 (N_10878,N_10093,N_9884);
or U10879 (N_10879,N_9712,N_9720);
nor U10880 (N_10880,N_9491,N_9237);
xnor U10881 (N_10881,N_10022,N_9986);
nand U10882 (N_10882,N_9758,N_9837);
xnor U10883 (N_10883,N_9964,N_9208);
and U10884 (N_10884,N_9742,N_9062);
and U10885 (N_10885,N_9998,N_9390);
and U10886 (N_10886,N_9416,N_9272);
nor U10887 (N_10887,N_10197,N_10371);
nand U10888 (N_10888,N_10475,N_10313);
nand U10889 (N_10889,N_9610,N_9766);
nor U10890 (N_10890,N_9113,N_9320);
or U10891 (N_10891,N_10016,N_9912);
xnor U10892 (N_10892,N_9021,N_9400);
nand U10893 (N_10893,N_10007,N_9687);
and U10894 (N_10894,N_10260,N_9876);
nor U10895 (N_10895,N_10251,N_9439);
and U10896 (N_10896,N_9638,N_9195);
or U10897 (N_10897,N_9371,N_9245);
nand U10898 (N_10898,N_9650,N_9660);
nor U10899 (N_10899,N_10363,N_9653);
and U10900 (N_10900,N_10431,N_10430);
and U10901 (N_10901,N_9634,N_9452);
nand U10902 (N_10902,N_9143,N_9328);
xor U10903 (N_10903,N_9207,N_9151);
nand U10904 (N_10904,N_10010,N_10403);
nand U10905 (N_10905,N_10037,N_9281);
xor U10906 (N_10906,N_10443,N_9095);
nor U10907 (N_10907,N_9025,N_10337);
and U10908 (N_10908,N_9901,N_9327);
and U10909 (N_10909,N_9366,N_10079);
nand U10910 (N_10910,N_9883,N_10214);
xnor U10911 (N_10911,N_9738,N_9885);
nor U10912 (N_10912,N_9768,N_9686);
and U10913 (N_10913,N_9183,N_9240);
xor U10914 (N_10914,N_10458,N_9642);
nor U10915 (N_10915,N_9804,N_10243);
nor U10916 (N_10916,N_9670,N_9614);
nor U10917 (N_10917,N_10396,N_9917);
xnor U10918 (N_10918,N_9564,N_9962);
nand U10919 (N_10919,N_9753,N_9699);
xor U10920 (N_10920,N_9702,N_9003);
xnor U10921 (N_10921,N_9028,N_9405);
nand U10922 (N_10922,N_9732,N_10440);
nor U10923 (N_10923,N_9457,N_10132);
nor U10924 (N_10924,N_10220,N_9192);
xnor U10925 (N_10925,N_10270,N_10452);
nor U10926 (N_10926,N_9838,N_9253);
nand U10927 (N_10927,N_9711,N_10317);
or U10928 (N_10928,N_10000,N_9918);
nor U10929 (N_10929,N_10229,N_9418);
nand U10930 (N_10930,N_9168,N_9697);
nor U10931 (N_10931,N_9745,N_9797);
xor U10932 (N_10932,N_9256,N_10134);
xor U10933 (N_10933,N_9556,N_10424);
nor U10934 (N_10934,N_9027,N_9044);
nand U10935 (N_10935,N_9809,N_9728);
xnor U10936 (N_10936,N_10040,N_10367);
nand U10937 (N_10937,N_9521,N_10397);
nor U10938 (N_10938,N_10392,N_9104);
nand U10939 (N_10939,N_9501,N_9112);
nand U10940 (N_10940,N_9587,N_9355);
nand U10941 (N_10941,N_9266,N_9295);
and U10942 (N_10942,N_10275,N_10069);
and U10943 (N_10943,N_9411,N_9703);
nand U10944 (N_10944,N_9430,N_9442);
or U10945 (N_10945,N_9635,N_9656);
or U10946 (N_10946,N_9781,N_9987);
xor U10947 (N_10947,N_9933,N_10159);
nand U10948 (N_10948,N_10379,N_9093);
nor U10949 (N_10949,N_9579,N_10198);
and U10950 (N_10950,N_9034,N_9234);
nor U10951 (N_10951,N_10261,N_9243);
xor U10952 (N_10952,N_10088,N_9205);
or U10953 (N_10953,N_9260,N_10351);
and U10954 (N_10954,N_10121,N_9774);
and U10955 (N_10955,N_9727,N_9522);
or U10956 (N_10956,N_9860,N_9988);
or U10957 (N_10957,N_10217,N_10062);
or U10958 (N_10958,N_10239,N_9166);
and U10959 (N_10959,N_9470,N_9603);
xnor U10960 (N_10960,N_9449,N_10050);
and U10961 (N_10961,N_9321,N_10042);
nand U10962 (N_10962,N_9757,N_9111);
or U10963 (N_10963,N_9040,N_9246);
or U10964 (N_10964,N_10347,N_9404);
or U10965 (N_10965,N_9643,N_10320);
xor U10966 (N_10966,N_10360,N_9816);
or U10967 (N_10967,N_9897,N_10482);
or U10968 (N_10968,N_9829,N_9503);
and U10969 (N_10969,N_9925,N_9554);
or U10970 (N_10970,N_9970,N_10005);
xor U10971 (N_10971,N_10145,N_10039);
xnor U10972 (N_10972,N_10025,N_9750);
nand U10973 (N_10973,N_9017,N_9710);
and U10974 (N_10974,N_9677,N_9651);
nand U10975 (N_10975,N_9079,N_9808);
or U10976 (N_10976,N_9540,N_9597);
xnor U10977 (N_10977,N_10063,N_10072);
and U10978 (N_10978,N_10060,N_9553);
nor U10979 (N_10979,N_10156,N_9547);
nand U10980 (N_10980,N_9354,N_9747);
nor U10981 (N_10981,N_9735,N_10157);
and U10982 (N_10982,N_9524,N_10240);
nand U10983 (N_10983,N_9570,N_10427);
nand U10984 (N_10984,N_9531,N_10254);
xnor U10985 (N_10985,N_10105,N_10459);
xor U10986 (N_10986,N_9482,N_9870);
nor U10987 (N_10987,N_9085,N_10417);
and U10988 (N_10988,N_9114,N_9701);
or U10989 (N_10989,N_9765,N_9565);
xor U10990 (N_10990,N_9740,N_9339);
or U10991 (N_10991,N_10382,N_9332);
nand U10992 (N_10992,N_10245,N_10447);
xor U10993 (N_10993,N_9209,N_9462);
xor U10994 (N_10994,N_10419,N_9477);
or U10995 (N_10995,N_10378,N_9092);
xor U10996 (N_10996,N_9487,N_9427);
xor U10997 (N_10997,N_9049,N_10100);
nor U10998 (N_10998,N_9381,N_9764);
and U10999 (N_10999,N_9824,N_10189);
or U11000 (N_11000,N_9908,N_9668);
nand U11001 (N_11001,N_10036,N_10227);
or U11002 (N_11002,N_9137,N_9419);
xnor U11003 (N_11003,N_10491,N_10497);
nor U11004 (N_11004,N_10316,N_9971);
nand U11005 (N_11005,N_9219,N_9417);
nand U11006 (N_11006,N_10289,N_9982);
xor U11007 (N_11007,N_9255,N_9361);
nor U11008 (N_11008,N_9409,N_10492);
nor U11009 (N_11009,N_10340,N_9927);
nand U11010 (N_11010,N_9014,N_9144);
xor U11011 (N_11011,N_10194,N_9800);
or U11012 (N_11012,N_10216,N_9061);
nor U11013 (N_11013,N_10318,N_9046);
nor U11014 (N_11014,N_9946,N_9472);
xnor U11015 (N_11015,N_10054,N_9244);
nor U11016 (N_11016,N_9399,N_9833);
and U11017 (N_11017,N_9776,N_9453);
nor U11018 (N_11018,N_9913,N_9225);
or U11019 (N_11019,N_10339,N_9539);
xor U11020 (N_11020,N_9270,N_9694);
xnor U11021 (N_11021,N_9202,N_9680);
nand U11022 (N_11022,N_9224,N_9331);
xor U11023 (N_11023,N_9378,N_9451);
xor U11024 (N_11024,N_10319,N_9099);
nor U11025 (N_11025,N_10029,N_10374);
or U11026 (N_11026,N_9828,N_9977);
xnor U11027 (N_11027,N_9552,N_10246);
and U11028 (N_11028,N_9350,N_10212);
nand U11029 (N_11029,N_9267,N_9413);
nor U11030 (N_11030,N_9395,N_9428);
nand U11031 (N_11031,N_9881,N_10175);
or U11032 (N_11032,N_10201,N_9455);
nand U11033 (N_11033,N_10327,N_9992);
and U11034 (N_11034,N_9315,N_10463);
and U11035 (N_11035,N_9433,N_10019);
nor U11036 (N_11036,N_9607,N_9193);
xor U11037 (N_11037,N_10149,N_9210);
nor U11038 (N_11038,N_10362,N_9336);
and U11039 (N_11039,N_10006,N_9356);
xor U11040 (N_11040,N_10111,N_9975);
xnor U11041 (N_11041,N_10466,N_9386);
and U11042 (N_11042,N_10028,N_10065);
nor U11043 (N_11043,N_10221,N_9581);
and U11044 (N_11044,N_10171,N_9005);
xnor U11045 (N_11045,N_9494,N_9393);
or U11046 (N_11046,N_9473,N_9631);
nor U11047 (N_11047,N_10389,N_9865);
xnor U11048 (N_11048,N_10052,N_9649);
nor U11049 (N_11049,N_9138,N_9053);
and U11050 (N_11050,N_9269,N_10284);
xor U11051 (N_11051,N_9953,N_9164);
and U11052 (N_11052,N_9022,N_9567);
xnor U11053 (N_11053,N_9644,N_9664);
nor U11054 (N_11054,N_9375,N_9952);
and U11055 (N_11055,N_10499,N_10153);
or U11056 (N_11056,N_10453,N_9145);
nand U11057 (N_11057,N_10405,N_9940);
nor U11058 (N_11058,N_9057,N_10404);
xor U11059 (N_11059,N_9600,N_9569);
nor U11060 (N_11060,N_9174,N_9077);
and U11061 (N_11061,N_9083,N_9754);
nor U11062 (N_11062,N_10292,N_9292);
nor U11063 (N_11063,N_10493,N_9124);
and U11064 (N_11064,N_10432,N_10090);
nor U11065 (N_11065,N_9002,N_9141);
or U11066 (N_11066,N_9029,N_9290);
or U11067 (N_11067,N_9958,N_9840);
nand U11068 (N_11068,N_9429,N_10271);
or U11069 (N_11069,N_9402,N_10495);
nor U11070 (N_11070,N_9479,N_10181);
nand U11071 (N_11071,N_9422,N_9117);
or U11072 (N_11072,N_9731,N_10364);
or U11073 (N_11073,N_9759,N_9707);
nor U11074 (N_11074,N_10026,N_9389);
and U11075 (N_11075,N_10195,N_10139);
or U11076 (N_11076,N_10045,N_10361);
and U11077 (N_11077,N_9063,N_9619);
nor U11078 (N_11078,N_9616,N_9385);
xnor U11079 (N_11079,N_9801,N_9369);
and U11080 (N_11080,N_9443,N_10172);
and U11081 (N_11081,N_10101,N_9396);
nor U11082 (N_11082,N_9311,N_10286);
xor U11083 (N_11083,N_9447,N_9688);
nor U11084 (N_11084,N_9294,N_10163);
or U11085 (N_11085,N_9506,N_10224);
nand U11086 (N_11086,N_9289,N_9412);
nand U11087 (N_11087,N_9559,N_9640);
nor U11088 (N_11088,N_10071,N_10394);
xnor U11089 (N_11089,N_10416,N_9538);
or U11090 (N_11090,N_9779,N_9231);
nor U11091 (N_11091,N_10094,N_9065);
and U11092 (N_11092,N_9133,N_10076);
nand U11093 (N_11093,N_9778,N_9629);
nand U11094 (N_11094,N_9353,N_9170);
and U11095 (N_11095,N_9994,N_10020);
or U11096 (N_11096,N_10280,N_9500);
xor U11097 (N_11097,N_9076,N_9648);
and U11098 (N_11098,N_9434,N_9931);
and U11099 (N_11099,N_10014,N_9675);
xnor U11100 (N_11100,N_9300,N_9158);
nor U11101 (N_11101,N_9866,N_9377);
nand U11102 (N_11102,N_9150,N_10115);
xnor U11103 (N_11103,N_9826,N_9041);
nand U11104 (N_11104,N_10402,N_10259);
nor U11105 (N_11105,N_9314,N_9180);
and U11106 (N_11106,N_9156,N_9898);
nand U11107 (N_11107,N_9598,N_9087);
nor U11108 (N_11108,N_10298,N_9084);
and U11109 (N_11109,N_9196,N_9729);
nor U11110 (N_11110,N_9495,N_9211);
or U11111 (N_11111,N_9182,N_9499);
xor U11112 (N_11112,N_9186,N_9121);
nand U11113 (N_11113,N_10255,N_10070);
and U11114 (N_11114,N_9505,N_9051);
nand U11115 (N_11115,N_9055,N_10031);
nor U11116 (N_11116,N_9157,N_9123);
or U11117 (N_11117,N_9792,N_9763);
nor U11118 (N_11118,N_10131,N_9690);
nand U11119 (N_11119,N_9420,N_10113);
xnor U11120 (N_11120,N_9887,N_9436);
and U11121 (N_11121,N_9777,N_10380);
or U11122 (N_11122,N_9497,N_10160);
nand U11123 (N_11123,N_9767,N_9215);
nand U11124 (N_11124,N_9902,N_10164);
or U11125 (N_11125,N_9541,N_9463);
nand U11126 (N_11126,N_9851,N_9793);
and U11127 (N_11127,N_9636,N_10222);
and U11128 (N_11128,N_9171,N_9149);
nor U11129 (N_11129,N_9705,N_10078);
nor U11130 (N_11130,N_9571,N_10150);
or U11131 (N_11131,N_9374,N_10438);
nand U11132 (N_11132,N_9576,N_10018);
nor U11133 (N_11133,N_9814,N_9335);
and U11134 (N_11134,N_9812,N_9212);
nor U11135 (N_11135,N_9821,N_9822);
nand U11136 (N_11136,N_9510,N_10206);
nand U11137 (N_11137,N_10081,N_9176);
or U11138 (N_11138,N_9031,N_9229);
nor U11139 (N_11139,N_9875,N_9148);
xor U11140 (N_11140,N_10287,N_10129);
xor U11141 (N_11141,N_9139,N_9308);
xnor U11142 (N_11142,N_10449,N_9265);
and U11143 (N_11143,N_10228,N_9125);
nand U11144 (N_11144,N_9746,N_9373);
and U11145 (N_11145,N_10277,N_9672);
nand U11146 (N_11146,N_10250,N_9326);
and U11147 (N_11147,N_9762,N_10332);
and U11148 (N_11148,N_9323,N_10283);
xor U11149 (N_11149,N_9963,N_10264);
and U11150 (N_11150,N_10409,N_9895);
xor U11151 (N_11151,N_9557,N_9948);
nor U11152 (N_11152,N_9973,N_10053);
nor U11153 (N_11153,N_9789,N_9519);
or U11154 (N_11154,N_9406,N_10310);
or U11155 (N_11155,N_10274,N_9073);
xnor U11156 (N_11156,N_9109,N_9787);
nand U11157 (N_11157,N_10204,N_9830);
xnor U11158 (N_11158,N_9471,N_9932);
and U11159 (N_11159,N_10027,N_9333);
xnor U11160 (N_11160,N_9715,N_10483);
nand U11161 (N_11161,N_9222,N_10128);
or U11162 (N_11162,N_9010,N_10017);
or U11163 (N_11163,N_9116,N_9647);
nor U11164 (N_11164,N_9841,N_9879);
nor U11165 (N_11165,N_9223,N_9131);
nor U11166 (N_11166,N_9548,N_10165);
and U11167 (N_11167,N_9189,N_9334);
nand U11168 (N_11168,N_9575,N_9827);
nand U11169 (N_11169,N_9861,N_9298);
or U11170 (N_11170,N_10477,N_10141);
or U11171 (N_11171,N_10305,N_9583);
xnor U11172 (N_11172,N_9286,N_9020);
or U11173 (N_11173,N_9488,N_9817);
or U11174 (N_11174,N_10445,N_9739);
xnor U11175 (N_11175,N_10390,N_9362);
xor U11176 (N_11176,N_9343,N_9957);
or U11177 (N_11177,N_9060,N_9380);
or U11178 (N_11178,N_9914,N_9407);
and U11179 (N_11179,N_9502,N_9015);
or U11180 (N_11180,N_9676,N_9622);
nand U11181 (N_11181,N_9006,N_10472);
or U11182 (N_11182,N_9941,N_9424);
xnor U11183 (N_11183,N_10190,N_9235);
and U11184 (N_11184,N_9214,N_9796);
nor U11185 (N_11185,N_9032,N_9016);
or U11186 (N_11186,N_9250,N_9536);
or U11187 (N_11187,N_9050,N_9513);
nand U11188 (N_11188,N_9039,N_10296);
nand U11189 (N_11189,N_10444,N_9346);
and U11190 (N_11190,N_9785,N_10413);
nor U11191 (N_11191,N_10350,N_9663);
nand U11192 (N_11192,N_9435,N_10474);
or U11193 (N_11193,N_9516,N_9630);
nor U11194 (N_11194,N_9388,N_10176);
nor U11195 (N_11195,N_9142,N_10248);
xnor U11196 (N_11196,N_9691,N_10302);
xor U11197 (N_11197,N_9316,N_9984);
or U11198 (N_11198,N_9048,N_9685);
xnor U11199 (N_11199,N_9467,N_9618);
and U11200 (N_11200,N_10058,N_9802);
nand U11201 (N_11201,N_9365,N_9877);
nand U11202 (N_11202,N_10038,N_9922);
nor U11203 (N_11203,N_9194,N_9788);
and U11204 (N_11204,N_10193,N_9633);
and U11205 (N_11205,N_9167,N_9199);
and U11206 (N_11206,N_9382,N_10233);
or U11207 (N_11207,N_10423,N_9072);
nor U11208 (N_11208,N_10202,N_9216);
xor U11209 (N_11209,N_10300,N_10056);
or U11210 (N_11210,N_10410,N_9939);
xor U11211 (N_11211,N_10148,N_9271);
xor U11212 (N_11212,N_9165,N_10468);
nor U11213 (N_11213,N_10187,N_10372);
and U11214 (N_11214,N_9847,N_9704);
or U11215 (N_11215,N_9593,N_9916);
and U11216 (N_11216,N_9825,N_9721);
nand U11217 (N_11217,N_9996,N_9191);
and U11218 (N_11218,N_9780,N_9573);
xor U11219 (N_11219,N_10085,N_9713);
and U11220 (N_11220,N_10192,N_9983);
nor U11221 (N_11221,N_9989,N_10086);
nor U11222 (N_11222,N_9834,N_10338);
or U11223 (N_11223,N_9551,N_10046);
nand U11224 (N_11224,N_9481,N_9937);
or U11225 (N_11225,N_9492,N_10184);
and U11226 (N_11226,N_10481,N_10341);
or U11227 (N_11227,N_9178,N_9755);
or U11228 (N_11228,N_9363,N_10215);
nor U11229 (N_11229,N_10161,N_9929);
nor U11230 (N_11230,N_10290,N_9592);
and U11231 (N_11231,N_9857,N_9134);
and U11232 (N_11232,N_10219,N_10218);
xor U11233 (N_11233,N_10106,N_9832);
xor U11234 (N_11234,N_10177,N_10406);
nor U11235 (N_11235,N_10213,N_9410);
xnor U11236 (N_11236,N_10355,N_9140);
nand U11237 (N_11237,N_9748,N_10188);
nor U11238 (N_11238,N_9654,N_10247);
xnor U11239 (N_11239,N_9309,N_9358);
or U11240 (N_11240,N_10306,N_10301);
and U11241 (N_11241,N_10346,N_9741);
nor U11242 (N_11242,N_9585,N_10325);
xnor U11243 (N_11243,N_9129,N_10428);
nand U11244 (N_11244,N_9277,N_10368);
nor U11245 (N_11245,N_10135,N_9951);
nand U11246 (N_11246,N_9317,N_9262);
xor U11247 (N_11247,N_9775,N_9096);
or U11248 (N_11248,N_10308,N_9906);
nor U11249 (N_11249,N_9529,N_9844);
xnor U11250 (N_11250,N_9215,N_9921);
or U11251 (N_11251,N_9908,N_9072);
or U11252 (N_11252,N_9975,N_10134);
and U11253 (N_11253,N_10454,N_9577);
or U11254 (N_11254,N_9481,N_10144);
xnor U11255 (N_11255,N_9249,N_9163);
xnor U11256 (N_11256,N_9964,N_9804);
nor U11257 (N_11257,N_9464,N_9211);
nand U11258 (N_11258,N_9746,N_9483);
xor U11259 (N_11259,N_10070,N_9050);
and U11260 (N_11260,N_10494,N_9081);
nor U11261 (N_11261,N_9472,N_10176);
or U11262 (N_11262,N_10432,N_9863);
xnor U11263 (N_11263,N_9061,N_9696);
and U11264 (N_11264,N_9169,N_9897);
nand U11265 (N_11265,N_9656,N_9936);
xor U11266 (N_11266,N_10217,N_10116);
and U11267 (N_11267,N_9680,N_9110);
xnor U11268 (N_11268,N_10195,N_10260);
xnor U11269 (N_11269,N_10128,N_9796);
nand U11270 (N_11270,N_9332,N_9275);
xnor U11271 (N_11271,N_10271,N_9161);
and U11272 (N_11272,N_10239,N_10344);
xor U11273 (N_11273,N_10220,N_9983);
xnor U11274 (N_11274,N_9441,N_10428);
and U11275 (N_11275,N_10492,N_9657);
or U11276 (N_11276,N_9414,N_9743);
and U11277 (N_11277,N_10243,N_9049);
and U11278 (N_11278,N_9825,N_9680);
and U11279 (N_11279,N_10023,N_9767);
or U11280 (N_11280,N_10123,N_9182);
and U11281 (N_11281,N_10496,N_9710);
nand U11282 (N_11282,N_9808,N_9498);
xnor U11283 (N_11283,N_9865,N_9328);
or U11284 (N_11284,N_10273,N_9416);
nor U11285 (N_11285,N_10480,N_9139);
nor U11286 (N_11286,N_9210,N_9171);
and U11287 (N_11287,N_9231,N_9963);
nand U11288 (N_11288,N_9930,N_9219);
nor U11289 (N_11289,N_10094,N_9127);
or U11290 (N_11290,N_9502,N_10132);
and U11291 (N_11291,N_9926,N_10139);
and U11292 (N_11292,N_9729,N_9104);
nand U11293 (N_11293,N_9870,N_9844);
and U11294 (N_11294,N_9008,N_10106);
xnor U11295 (N_11295,N_9558,N_9857);
xor U11296 (N_11296,N_9346,N_9758);
nand U11297 (N_11297,N_9237,N_9064);
nor U11298 (N_11298,N_10300,N_9711);
and U11299 (N_11299,N_10034,N_10321);
nor U11300 (N_11300,N_9725,N_9880);
xor U11301 (N_11301,N_9601,N_9213);
or U11302 (N_11302,N_9348,N_9314);
nand U11303 (N_11303,N_9445,N_10322);
and U11304 (N_11304,N_9171,N_10211);
nor U11305 (N_11305,N_9898,N_10384);
and U11306 (N_11306,N_10101,N_9835);
nor U11307 (N_11307,N_10425,N_9753);
nand U11308 (N_11308,N_9132,N_9292);
xnor U11309 (N_11309,N_9448,N_9251);
nor U11310 (N_11310,N_9604,N_9894);
xor U11311 (N_11311,N_9424,N_9367);
or U11312 (N_11312,N_9071,N_10102);
nor U11313 (N_11313,N_9851,N_10132);
and U11314 (N_11314,N_10058,N_9189);
and U11315 (N_11315,N_10269,N_10275);
nand U11316 (N_11316,N_9971,N_10198);
xor U11317 (N_11317,N_9486,N_9412);
nand U11318 (N_11318,N_9471,N_9465);
and U11319 (N_11319,N_10138,N_10309);
and U11320 (N_11320,N_9264,N_10346);
nand U11321 (N_11321,N_9393,N_9985);
nor U11322 (N_11322,N_9437,N_9714);
or U11323 (N_11323,N_9283,N_10057);
xor U11324 (N_11324,N_9379,N_9071);
nor U11325 (N_11325,N_9746,N_10196);
nand U11326 (N_11326,N_9943,N_9276);
or U11327 (N_11327,N_9793,N_10224);
and U11328 (N_11328,N_9515,N_9434);
xnor U11329 (N_11329,N_9574,N_10321);
nand U11330 (N_11330,N_10313,N_9898);
nand U11331 (N_11331,N_9926,N_9512);
or U11332 (N_11332,N_9153,N_9786);
nand U11333 (N_11333,N_10470,N_10201);
xnor U11334 (N_11334,N_9133,N_10411);
nand U11335 (N_11335,N_9406,N_9407);
or U11336 (N_11336,N_10098,N_9283);
and U11337 (N_11337,N_10305,N_9989);
nor U11338 (N_11338,N_9074,N_9180);
nand U11339 (N_11339,N_10108,N_9751);
or U11340 (N_11340,N_9324,N_9919);
or U11341 (N_11341,N_9074,N_10025);
or U11342 (N_11342,N_9241,N_9638);
or U11343 (N_11343,N_9354,N_9893);
and U11344 (N_11344,N_10029,N_9891);
and U11345 (N_11345,N_10251,N_10245);
nor U11346 (N_11346,N_9605,N_9251);
nor U11347 (N_11347,N_10344,N_9575);
xor U11348 (N_11348,N_9054,N_9091);
nand U11349 (N_11349,N_10378,N_9951);
or U11350 (N_11350,N_10306,N_10436);
and U11351 (N_11351,N_9010,N_9546);
xor U11352 (N_11352,N_10320,N_9849);
nor U11353 (N_11353,N_9185,N_10405);
nand U11354 (N_11354,N_10165,N_9151);
nor U11355 (N_11355,N_10297,N_9841);
or U11356 (N_11356,N_10129,N_9089);
or U11357 (N_11357,N_9457,N_9076);
or U11358 (N_11358,N_10216,N_9223);
nand U11359 (N_11359,N_9590,N_9710);
nand U11360 (N_11360,N_9372,N_9828);
or U11361 (N_11361,N_10239,N_9811);
nand U11362 (N_11362,N_10239,N_10018);
nor U11363 (N_11363,N_9967,N_9352);
xor U11364 (N_11364,N_9533,N_9589);
nand U11365 (N_11365,N_9009,N_9903);
and U11366 (N_11366,N_9525,N_9069);
or U11367 (N_11367,N_9266,N_10411);
or U11368 (N_11368,N_10023,N_9853);
and U11369 (N_11369,N_9272,N_9586);
xor U11370 (N_11370,N_9477,N_9493);
nor U11371 (N_11371,N_10134,N_9390);
nand U11372 (N_11372,N_9502,N_10332);
nand U11373 (N_11373,N_9038,N_9296);
nor U11374 (N_11374,N_9433,N_10454);
nand U11375 (N_11375,N_10009,N_10186);
nor U11376 (N_11376,N_9065,N_10225);
xnor U11377 (N_11377,N_10305,N_9940);
or U11378 (N_11378,N_10030,N_9271);
or U11379 (N_11379,N_10398,N_9021);
nor U11380 (N_11380,N_9407,N_10085);
and U11381 (N_11381,N_9823,N_9781);
and U11382 (N_11382,N_10149,N_9480);
and U11383 (N_11383,N_9345,N_9519);
or U11384 (N_11384,N_9370,N_9330);
and U11385 (N_11385,N_10071,N_9275);
and U11386 (N_11386,N_9593,N_9208);
xnor U11387 (N_11387,N_9019,N_9608);
xor U11388 (N_11388,N_10093,N_10075);
or U11389 (N_11389,N_10079,N_10195);
xnor U11390 (N_11390,N_9083,N_10074);
nand U11391 (N_11391,N_9254,N_10472);
or U11392 (N_11392,N_9888,N_9980);
xor U11393 (N_11393,N_9734,N_10376);
and U11394 (N_11394,N_10223,N_10422);
nand U11395 (N_11395,N_9823,N_9378);
nor U11396 (N_11396,N_9475,N_9627);
or U11397 (N_11397,N_9707,N_9686);
and U11398 (N_11398,N_9977,N_9701);
and U11399 (N_11399,N_9880,N_9696);
or U11400 (N_11400,N_9047,N_9289);
nand U11401 (N_11401,N_9089,N_9762);
xor U11402 (N_11402,N_10210,N_9299);
nor U11403 (N_11403,N_10458,N_10485);
xnor U11404 (N_11404,N_10075,N_10321);
and U11405 (N_11405,N_10033,N_10476);
and U11406 (N_11406,N_9397,N_9614);
nand U11407 (N_11407,N_9896,N_10452);
or U11408 (N_11408,N_9127,N_10225);
and U11409 (N_11409,N_9535,N_9121);
xnor U11410 (N_11410,N_10164,N_9986);
or U11411 (N_11411,N_10253,N_9315);
and U11412 (N_11412,N_10328,N_10284);
xnor U11413 (N_11413,N_9609,N_9749);
and U11414 (N_11414,N_9928,N_10230);
and U11415 (N_11415,N_9493,N_10170);
nand U11416 (N_11416,N_9739,N_10197);
nor U11417 (N_11417,N_9677,N_10152);
xnor U11418 (N_11418,N_9419,N_9268);
xor U11419 (N_11419,N_10268,N_9771);
nor U11420 (N_11420,N_10397,N_9449);
xor U11421 (N_11421,N_9390,N_9304);
nand U11422 (N_11422,N_9391,N_9872);
nand U11423 (N_11423,N_9908,N_10176);
and U11424 (N_11424,N_9134,N_9886);
and U11425 (N_11425,N_9102,N_10250);
xnor U11426 (N_11426,N_9446,N_10001);
nor U11427 (N_11427,N_9919,N_9345);
nand U11428 (N_11428,N_9972,N_10265);
xor U11429 (N_11429,N_9673,N_9505);
nor U11430 (N_11430,N_9656,N_9693);
xor U11431 (N_11431,N_10409,N_10371);
nand U11432 (N_11432,N_9068,N_9183);
or U11433 (N_11433,N_9392,N_10200);
and U11434 (N_11434,N_9321,N_9918);
and U11435 (N_11435,N_10420,N_9121);
nor U11436 (N_11436,N_9811,N_9697);
or U11437 (N_11437,N_9978,N_9136);
or U11438 (N_11438,N_9234,N_9327);
nor U11439 (N_11439,N_10225,N_9412);
nor U11440 (N_11440,N_9677,N_9702);
nand U11441 (N_11441,N_9494,N_9668);
or U11442 (N_11442,N_9858,N_9115);
nor U11443 (N_11443,N_10022,N_9723);
nand U11444 (N_11444,N_9641,N_9663);
and U11445 (N_11445,N_10127,N_9182);
xnor U11446 (N_11446,N_9660,N_9223);
or U11447 (N_11447,N_9252,N_9451);
nor U11448 (N_11448,N_10215,N_9773);
nor U11449 (N_11449,N_9691,N_9960);
and U11450 (N_11450,N_10103,N_10083);
nand U11451 (N_11451,N_10386,N_10403);
xnor U11452 (N_11452,N_10348,N_10362);
xor U11453 (N_11453,N_9522,N_10412);
and U11454 (N_11454,N_9459,N_9293);
nand U11455 (N_11455,N_10070,N_10193);
nor U11456 (N_11456,N_9447,N_10336);
and U11457 (N_11457,N_10130,N_9730);
nand U11458 (N_11458,N_9345,N_10015);
xor U11459 (N_11459,N_9928,N_9984);
nor U11460 (N_11460,N_10483,N_9094);
or U11461 (N_11461,N_9534,N_9224);
nand U11462 (N_11462,N_9886,N_9114);
and U11463 (N_11463,N_9400,N_9541);
xnor U11464 (N_11464,N_9628,N_10012);
or U11465 (N_11465,N_9386,N_10417);
or U11466 (N_11466,N_9526,N_9802);
xor U11467 (N_11467,N_9104,N_9543);
or U11468 (N_11468,N_9665,N_10019);
nor U11469 (N_11469,N_9589,N_9731);
nor U11470 (N_11470,N_9617,N_10338);
and U11471 (N_11471,N_10287,N_9535);
nor U11472 (N_11472,N_9471,N_9390);
nor U11473 (N_11473,N_10207,N_9425);
nand U11474 (N_11474,N_10369,N_9872);
xnor U11475 (N_11475,N_10353,N_9091);
or U11476 (N_11476,N_10424,N_9776);
xnor U11477 (N_11477,N_9731,N_9454);
or U11478 (N_11478,N_10291,N_9317);
xnor U11479 (N_11479,N_9368,N_10487);
and U11480 (N_11480,N_9099,N_10394);
and U11481 (N_11481,N_10159,N_9610);
nand U11482 (N_11482,N_10287,N_9359);
nand U11483 (N_11483,N_9497,N_9384);
nor U11484 (N_11484,N_9103,N_9219);
or U11485 (N_11485,N_9344,N_9885);
nor U11486 (N_11486,N_10238,N_9546);
nand U11487 (N_11487,N_9665,N_9049);
and U11488 (N_11488,N_9586,N_9483);
nand U11489 (N_11489,N_10132,N_10139);
nor U11490 (N_11490,N_10381,N_9978);
and U11491 (N_11491,N_9967,N_10349);
nor U11492 (N_11492,N_9470,N_10262);
nand U11493 (N_11493,N_9745,N_9598);
nand U11494 (N_11494,N_10053,N_9735);
xor U11495 (N_11495,N_9414,N_9283);
and U11496 (N_11496,N_9287,N_9722);
nor U11497 (N_11497,N_9769,N_9747);
and U11498 (N_11498,N_9255,N_10204);
and U11499 (N_11499,N_9597,N_9623);
nor U11500 (N_11500,N_9624,N_10336);
xnor U11501 (N_11501,N_9719,N_9959);
nand U11502 (N_11502,N_9843,N_10475);
nand U11503 (N_11503,N_9511,N_10052);
nor U11504 (N_11504,N_9259,N_9896);
nor U11505 (N_11505,N_9672,N_9663);
and U11506 (N_11506,N_9145,N_9853);
and U11507 (N_11507,N_9413,N_9233);
nand U11508 (N_11508,N_9535,N_9858);
or U11509 (N_11509,N_9717,N_9587);
nand U11510 (N_11510,N_10413,N_9085);
and U11511 (N_11511,N_9276,N_10221);
or U11512 (N_11512,N_9007,N_9271);
nand U11513 (N_11513,N_9005,N_10406);
or U11514 (N_11514,N_10150,N_10422);
nand U11515 (N_11515,N_9591,N_10363);
xnor U11516 (N_11516,N_9422,N_9458);
or U11517 (N_11517,N_9653,N_9337);
nor U11518 (N_11518,N_10123,N_9430);
xor U11519 (N_11519,N_9216,N_9864);
nand U11520 (N_11520,N_10286,N_10004);
xor U11521 (N_11521,N_10255,N_10106);
or U11522 (N_11522,N_9027,N_9244);
nand U11523 (N_11523,N_9065,N_10010);
nand U11524 (N_11524,N_9200,N_10061);
nor U11525 (N_11525,N_10042,N_9864);
xnor U11526 (N_11526,N_9382,N_10279);
and U11527 (N_11527,N_9806,N_9162);
and U11528 (N_11528,N_9987,N_9184);
or U11529 (N_11529,N_9344,N_10383);
nor U11530 (N_11530,N_9923,N_10024);
nor U11531 (N_11531,N_9597,N_9554);
and U11532 (N_11532,N_9899,N_9326);
nor U11533 (N_11533,N_10387,N_10363);
and U11534 (N_11534,N_10291,N_10265);
xor U11535 (N_11535,N_10476,N_9463);
nand U11536 (N_11536,N_10011,N_9625);
and U11537 (N_11537,N_9739,N_10361);
nor U11538 (N_11538,N_9278,N_9935);
nand U11539 (N_11539,N_10117,N_9462);
nor U11540 (N_11540,N_10073,N_10040);
or U11541 (N_11541,N_9156,N_9610);
or U11542 (N_11542,N_9835,N_9090);
and U11543 (N_11543,N_9310,N_9109);
xnor U11544 (N_11544,N_9215,N_9793);
and U11545 (N_11545,N_10199,N_9670);
and U11546 (N_11546,N_9624,N_9397);
and U11547 (N_11547,N_10499,N_10474);
xor U11548 (N_11548,N_9552,N_10018);
xnor U11549 (N_11549,N_10177,N_9738);
nand U11550 (N_11550,N_9205,N_9822);
nand U11551 (N_11551,N_10427,N_9470);
or U11552 (N_11552,N_9586,N_10166);
nor U11553 (N_11553,N_10431,N_10022);
or U11554 (N_11554,N_9544,N_9484);
nand U11555 (N_11555,N_9186,N_9983);
or U11556 (N_11556,N_9467,N_9787);
xor U11557 (N_11557,N_9328,N_9988);
nand U11558 (N_11558,N_10237,N_10346);
and U11559 (N_11559,N_9754,N_10291);
or U11560 (N_11560,N_10359,N_10064);
or U11561 (N_11561,N_9279,N_9802);
and U11562 (N_11562,N_9653,N_9392);
and U11563 (N_11563,N_9177,N_9278);
and U11564 (N_11564,N_9846,N_9657);
or U11565 (N_11565,N_10021,N_9604);
and U11566 (N_11566,N_9393,N_9090);
and U11567 (N_11567,N_9520,N_10288);
nor U11568 (N_11568,N_9533,N_9234);
nand U11569 (N_11569,N_9703,N_9341);
or U11570 (N_11570,N_9509,N_9949);
xnor U11571 (N_11571,N_9541,N_9698);
or U11572 (N_11572,N_9668,N_9931);
nand U11573 (N_11573,N_9947,N_9692);
or U11574 (N_11574,N_9641,N_9591);
xor U11575 (N_11575,N_9294,N_9128);
nand U11576 (N_11576,N_10483,N_9653);
nand U11577 (N_11577,N_10034,N_9788);
xnor U11578 (N_11578,N_10313,N_9892);
or U11579 (N_11579,N_9713,N_9324);
nand U11580 (N_11580,N_10185,N_9345);
xor U11581 (N_11581,N_10278,N_10118);
xor U11582 (N_11582,N_10470,N_10185);
nor U11583 (N_11583,N_9627,N_9755);
nand U11584 (N_11584,N_10454,N_9708);
or U11585 (N_11585,N_9835,N_10186);
and U11586 (N_11586,N_9988,N_9999);
nand U11587 (N_11587,N_10177,N_9146);
and U11588 (N_11588,N_10400,N_10290);
nor U11589 (N_11589,N_9570,N_9741);
or U11590 (N_11590,N_9348,N_10263);
nand U11591 (N_11591,N_9363,N_9109);
or U11592 (N_11592,N_10039,N_9591);
xnor U11593 (N_11593,N_9826,N_9606);
or U11594 (N_11594,N_9012,N_9799);
or U11595 (N_11595,N_10091,N_9822);
and U11596 (N_11596,N_9145,N_10353);
nand U11597 (N_11597,N_9060,N_9955);
nor U11598 (N_11598,N_9210,N_9512);
xnor U11599 (N_11599,N_10250,N_9540);
xnor U11600 (N_11600,N_10496,N_9227);
xor U11601 (N_11601,N_9125,N_9538);
or U11602 (N_11602,N_9162,N_10497);
or U11603 (N_11603,N_9583,N_9095);
or U11604 (N_11604,N_9349,N_10497);
xor U11605 (N_11605,N_9495,N_9679);
and U11606 (N_11606,N_10265,N_9545);
nor U11607 (N_11607,N_10098,N_10336);
and U11608 (N_11608,N_9156,N_10157);
or U11609 (N_11609,N_10181,N_9741);
xnor U11610 (N_11610,N_10403,N_10354);
nor U11611 (N_11611,N_9944,N_9015);
nor U11612 (N_11612,N_9559,N_10335);
nor U11613 (N_11613,N_9310,N_9870);
or U11614 (N_11614,N_10281,N_10133);
nor U11615 (N_11615,N_9466,N_9344);
xor U11616 (N_11616,N_9190,N_9344);
nand U11617 (N_11617,N_9316,N_9732);
nor U11618 (N_11618,N_9729,N_10385);
nor U11619 (N_11619,N_10463,N_10215);
nor U11620 (N_11620,N_10430,N_10035);
nand U11621 (N_11621,N_9026,N_9030);
nand U11622 (N_11622,N_9368,N_9247);
nor U11623 (N_11623,N_9253,N_10387);
nor U11624 (N_11624,N_9078,N_10340);
and U11625 (N_11625,N_9947,N_9963);
or U11626 (N_11626,N_9973,N_10116);
nor U11627 (N_11627,N_10388,N_9890);
nor U11628 (N_11628,N_9795,N_9697);
nor U11629 (N_11629,N_9712,N_10011);
or U11630 (N_11630,N_9182,N_9262);
nor U11631 (N_11631,N_9096,N_9232);
nor U11632 (N_11632,N_10359,N_10155);
nor U11633 (N_11633,N_9116,N_10050);
nor U11634 (N_11634,N_10222,N_9889);
xnor U11635 (N_11635,N_9210,N_9750);
or U11636 (N_11636,N_10017,N_9661);
xor U11637 (N_11637,N_10276,N_9057);
xnor U11638 (N_11638,N_9369,N_9851);
and U11639 (N_11639,N_9910,N_9390);
nand U11640 (N_11640,N_9287,N_9707);
and U11641 (N_11641,N_9634,N_9302);
nand U11642 (N_11642,N_9243,N_9820);
nor U11643 (N_11643,N_9666,N_10140);
nand U11644 (N_11644,N_9672,N_10265);
or U11645 (N_11645,N_9583,N_10246);
xor U11646 (N_11646,N_9850,N_10139);
nand U11647 (N_11647,N_10286,N_9937);
and U11648 (N_11648,N_9046,N_10430);
xnor U11649 (N_11649,N_9304,N_9110);
or U11650 (N_11650,N_9945,N_9581);
xnor U11651 (N_11651,N_10484,N_10048);
or U11652 (N_11652,N_9729,N_10441);
xor U11653 (N_11653,N_9545,N_10489);
or U11654 (N_11654,N_9484,N_10110);
xor U11655 (N_11655,N_9429,N_9153);
xor U11656 (N_11656,N_10024,N_9676);
nand U11657 (N_11657,N_9126,N_9371);
xnor U11658 (N_11658,N_9708,N_10080);
nand U11659 (N_11659,N_9568,N_10447);
or U11660 (N_11660,N_10044,N_9067);
or U11661 (N_11661,N_10112,N_9441);
xnor U11662 (N_11662,N_9655,N_10157);
nand U11663 (N_11663,N_9627,N_9354);
or U11664 (N_11664,N_9156,N_9996);
and U11665 (N_11665,N_9279,N_9349);
nor U11666 (N_11666,N_9005,N_10064);
or U11667 (N_11667,N_9756,N_9706);
nand U11668 (N_11668,N_10053,N_10157);
nor U11669 (N_11669,N_9712,N_9424);
xor U11670 (N_11670,N_9436,N_9135);
or U11671 (N_11671,N_9962,N_9593);
xnor U11672 (N_11672,N_10115,N_9063);
nor U11673 (N_11673,N_9604,N_9571);
and U11674 (N_11674,N_9967,N_10026);
xnor U11675 (N_11675,N_9157,N_10098);
nor U11676 (N_11676,N_10272,N_9230);
nand U11677 (N_11677,N_9146,N_9706);
and U11678 (N_11678,N_10315,N_10091);
nand U11679 (N_11679,N_9364,N_9816);
nor U11680 (N_11680,N_10310,N_10410);
nand U11681 (N_11681,N_9034,N_9660);
nor U11682 (N_11682,N_9988,N_9787);
nor U11683 (N_11683,N_9776,N_9102);
nor U11684 (N_11684,N_10111,N_9411);
nor U11685 (N_11685,N_10070,N_9168);
or U11686 (N_11686,N_10405,N_9608);
and U11687 (N_11687,N_10119,N_9906);
xor U11688 (N_11688,N_9031,N_10111);
or U11689 (N_11689,N_9512,N_10166);
xor U11690 (N_11690,N_9746,N_9015);
xor U11691 (N_11691,N_9013,N_10323);
or U11692 (N_11692,N_9959,N_9629);
and U11693 (N_11693,N_9250,N_9538);
xnor U11694 (N_11694,N_10047,N_10149);
or U11695 (N_11695,N_10371,N_9465);
nor U11696 (N_11696,N_9835,N_9055);
nand U11697 (N_11697,N_10013,N_10418);
or U11698 (N_11698,N_9676,N_9727);
xnor U11699 (N_11699,N_10113,N_10202);
nor U11700 (N_11700,N_9776,N_9588);
nand U11701 (N_11701,N_10190,N_9692);
and U11702 (N_11702,N_9971,N_10435);
nand U11703 (N_11703,N_9587,N_10002);
nand U11704 (N_11704,N_9692,N_9789);
nor U11705 (N_11705,N_10365,N_9339);
nor U11706 (N_11706,N_9347,N_10203);
nand U11707 (N_11707,N_9802,N_10023);
nor U11708 (N_11708,N_10321,N_10289);
and U11709 (N_11709,N_9410,N_10238);
nand U11710 (N_11710,N_10150,N_9094);
and U11711 (N_11711,N_9561,N_10444);
or U11712 (N_11712,N_10120,N_9029);
xnor U11713 (N_11713,N_10270,N_9906);
and U11714 (N_11714,N_9544,N_10247);
or U11715 (N_11715,N_9637,N_9138);
and U11716 (N_11716,N_10208,N_9403);
nor U11717 (N_11717,N_10465,N_9342);
nor U11718 (N_11718,N_9433,N_10106);
nand U11719 (N_11719,N_10149,N_10174);
nand U11720 (N_11720,N_10052,N_10115);
xnor U11721 (N_11721,N_9652,N_10473);
or U11722 (N_11722,N_10250,N_10221);
xor U11723 (N_11723,N_9445,N_9871);
xor U11724 (N_11724,N_9198,N_10146);
xnor U11725 (N_11725,N_9622,N_9972);
or U11726 (N_11726,N_9629,N_9563);
nand U11727 (N_11727,N_10267,N_9791);
and U11728 (N_11728,N_9775,N_9263);
nor U11729 (N_11729,N_10125,N_9007);
or U11730 (N_11730,N_9775,N_9434);
nand U11731 (N_11731,N_9705,N_9954);
nand U11732 (N_11732,N_9234,N_9526);
or U11733 (N_11733,N_10491,N_9801);
or U11734 (N_11734,N_9487,N_9573);
xnor U11735 (N_11735,N_9564,N_10016);
or U11736 (N_11736,N_9922,N_9561);
or U11737 (N_11737,N_9049,N_10326);
nand U11738 (N_11738,N_9844,N_10429);
and U11739 (N_11739,N_9420,N_9472);
xor U11740 (N_11740,N_9847,N_10349);
xnor U11741 (N_11741,N_9019,N_10029);
or U11742 (N_11742,N_9224,N_10384);
or U11743 (N_11743,N_9003,N_9457);
xnor U11744 (N_11744,N_10050,N_9077);
nor U11745 (N_11745,N_9247,N_9519);
nand U11746 (N_11746,N_9453,N_10265);
and U11747 (N_11747,N_10100,N_10144);
xor U11748 (N_11748,N_9733,N_10455);
nor U11749 (N_11749,N_10358,N_9680);
or U11750 (N_11750,N_10250,N_10495);
or U11751 (N_11751,N_9148,N_10490);
or U11752 (N_11752,N_9095,N_9322);
or U11753 (N_11753,N_10212,N_10451);
or U11754 (N_11754,N_9101,N_9854);
nand U11755 (N_11755,N_9460,N_9233);
nor U11756 (N_11756,N_9798,N_9673);
or U11757 (N_11757,N_10355,N_9015);
xnor U11758 (N_11758,N_9902,N_9195);
or U11759 (N_11759,N_10069,N_9692);
xnor U11760 (N_11760,N_10118,N_9061);
or U11761 (N_11761,N_10219,N_9795);
and U11762 (N_11762,N_10064,N_10483);
nor U11763 (N_11763,N_10497,N_9638);
or U11764 (N_11764,N_9020,N_9863);
nand U11765 (N_11765,N_9432,N_9299);
nor U11766 (N_11766,N_9110,N_10169);
nor U11767 (N_11767,N_9668,N_9963);
or U11768 (N_11768,N_10453,N_9922);
xnor U11769 (N_11769,N_10400,N_9469);
nand U11770 (N_11770,N_10430,N_9008);
xor U11771 (N_11771,N_10096,N_10205);
or U11772 (N_11772,N_9975,N_10215);
or U11773 (N_11773,N_9652,N_10084);
nor U11774 (N_11774,N_9429,N_10031);
or U11775 (N_11775,N_9289,N_9253);
xor U11776 (N_11776,N_9072,N_9842);
or U11777 (N_11777,N_9962,N_10008);
xnor U11778 (N_11778,N_10181,N_9243);
and U11779 (N_11779,N_10048,N_10021);
xnor U11780 (N_11780,N_9511,N_9544);
nand U11781 (N_11781,N_9954,N_10393);
nand U11782 (N_11782,N_9560,N_9200);
xnor U11783 (N_11783,N_9932,N_9231);
or U11784 (N_11784,N_10137,N_9002);
nor U11785 (N_11785,N_10282,N_9318);
xnor U11786 (N_11786,N_9680,N_10472);
nand U11787 (N_11787,N_9405,N_9044);
nand U11788 (N_11788,N_9257,N_10094);
and U11789 (N_11789,N_9498,N_9755);
nor U11790 (N_11790,N_10260,N_9582);
xor U11791 (N_11791,N_10260,N_10095);
nand U11792 (N_11792,N_10258,N_9651);
nand U11793 (N_11793,N_10410,N_10003);
nor U11794 (N_11794,N_10126,N_10142);
or U11795 (N_11795,N_10222,N_9139);
and U11796 (N_11796,N_9866,N_10353);
nand U11797 (N_11797,N_9565,N_9369);
or U11798 (N_11798,N_9807,N_9022);
xnor U11799 (N_11799,N_9892,N_9999);
xnor U11800 (N_11800,N_9270,N_9232);
xnor U11801 (N_11801,N_9233,N_10107);
and U11802 (N_11802,N_9594,N_10144);
or U11803 (N_11803,N_10083,N_9971);
or U11804 (N_11804,N_10387,N_9535);
and U11805 (N_11805,N_9486,N_9091);
xor U11806 (N_11806,N_10203,N_9989);
xor U11807 (N_11807,N_9305,N_9493);
nand U11808 (N_11808,N_10282,N_10461);
xnor U11809 (N_11809,N_10118,N_9688);
nand U11810 (N_11810,N_9136,N_10344);
or U11811 (N_11811,N_9699,N_9581);
or U11812 (N_11812,N_9596,N_10491);
and U11813 (N_11813,N_10345,N_9610);
nand U11814 (N_11814,N_9933,N_9175);
nand U11815 (N_11815,N_9755,N_9757);
or U11816 (N_11816,N_9426,N_9691);
nand U11817 (N_11817,N_9291,N_9243);
nand U11818 (N_11818,N_10031,N_10488);
and U11819 (N_11819,N_9712,N_10018);
nand U11820 (N_11820,N_10357,N_10411);
and U11821 (N_11821,N_9869,N_9501);
nor U11822 (N_11822,N_10239,N_10140);
xnor U11823 (N_11823,N_9516,N_9568);
xor U11824 (N_11824,N_9000,N_9017);
nor U11825 (N_11825,N_9958,N_9279);
xor U11826 (N_11826,N_9007,N_9586);
nand U11827 (N_11827,N_10251,N_9075);
xnor U11828 (N_11828,N_9885,N_9240);
xor U11829 (N_11829,N_10308,N_10085);
nand U11830 (N_11830,N_9285,N_9206);
nand U11831 (N_11831,N_10493,N_9955);
nor U11832 (N_11832,N_9673,N_9877);
or U11833 (N_11833,N_9324,N_9939);
and U11834 (N_11834,N_10018,N_9486);
or U11835 (N_11835,N_10330,N_9956);
and U11836 (N_11836,N_10028,N_10364);
nand U11837 (N_11837,N_10475,N_10082);
xor U11838 (N_11838,N_9845,N_9661);
nor U11839 (N_11839,N_10294,N_9142);
nor U11840 (N_11840,N_9158,N_9137);
nor U11841 (N_11841,N_9835,N_10399);
xnor U11842 (N_11842,N_9390,N_9500);
nor U11843 (N_11843,N_9783,N_10291);
and U11844 (N_11844,N_10395,N_9855);
nand U11845 (N_11845,N_9852,N_9939);
or U11846 (N_11846,N_9810,N_10075);
xor U11847 (N_11847,N_9243,N_9157);
nand U11848 (N_11848,N_9368,N_10020);
or U11849 (N_11849,N_9166,N_9870);
xnor U11850 (N_11850,N_9231,N_9948);
xor U11851 (N_11851,N_9022,N_9638);
nand U11852 (N_11852,N_10307,N_10073);
nor U11853 (N_11853,N_9778,N_10221);
nor U11854 (N_11854,N_9218,N_9665);
and U11855 (N_11855,N_9981,N_10337);
and U11856 (N_11856,N_9593,N_9414);
nor U11857 (N_11857,N_9085,N_10496);
nand U11858 (N_11858,N_9582,N_9387);
or U11859 (N_11859,N_9583,N_9305);
nand U11860 (N_11860,N_9766,N_9324);
xor U11861 (N_11861,N_9033,N_9791);
or U11862 (N_11862,N_9982,N_10263);
nand U11863 (N_11863,N_10065,N_9311);
nand U11864 (N_11864,N_9890,N_9929);
nor U11865 (N_11865,N_9924,N_10028);
and U11866 (N_11866,N_9967,N_10051);
or U11867 (N_11867,N_9911,N_10247);
or U11868 (N_11868,N_9252,N_9756);
and U11869 (N_11869,N_10227,N_10381);
or U11870 (N_11870,N_9685,N_9873);
xnor U11871 (N_11871,N_9372,N_9470);
nand U11872 (N_11872,N_10271,N_10138);
nand U11873 (N_11873,N_9187,N_9480);
xnor U11874 (N_11874,N_9680,N_10363);
nor U11875 (N_11875,N_9388,N_10299);
or U11876 (N_11876,N_9476,N_9366);
and U11877 (N_11877,N_9833,N_10044);
xor U11878 (N_11878,N_9927,N_9425);
and U11879 (N_11879,N_10168,N_9512);
or U11880 (N_11880,N_9745,N_9408);
and U11881 (N_11881,N_9674,N_10101);
and U11882 (N_11882,N_9963,N_9245);
nand U11883 (N_11883,N_9906,N_10076);
nor U11884 (N_11884,N_9635,N_10221);
or U11885 (N_11885,N_10355,N_10127);
or U11886 (N_11886,N_9098,N_10154);
and U11887 (N_11887,N_10066,N_10342);
and U11888 (N_11888,N_9991,N_9000);
nand U11889 (N_11889,N_10066,N_9716);
and U11890 (N_11890,N_9269,N_9978);
nand U11891 (N_11891,N_10135,N_9325);
and U11892 (N_11892,N_10240,N_9356);
nand U11893 (N_11893,N_9900,N_10401);
and U11894 (N_11894,N_9618,N_9516);
nor U11895 (N_11895,N_9830,N_9504);
xor U11896 (N_11896,N_10371,N_10479);
and U11897 (N_11897,N_10169,N_9863);
and U11898 (N_11898,N_10129,N_10254);
nor U11899 (N_11899,N_9562,N_9947);
nand U11900 (N_11900,N_10252,N_9444);
xor U11901 (N_11901,N_9980,N_9001);
nor U11902 (N_11902,N_10203,N_9495);
and U11903 (N_11903,N_10143,N_10204);
nand U11904 (N_11904,N_10177,N_9951);
xor U11905 (N_11905,N_9018,N_9912);
xor U11906 (N_11906,N_9542,N_10391);
xor U11907 (N_11907,N_10416,N_10022);
or U11908 (N_11908,N_9485,N_10027);
or U11909 (N_11909,N_10163,N_9314);
nand U11910 (N_11910,N_9992,N_9443);
and U11911 (N_11911,N_9863,N_10404);
or U11912 (N_11912,N_10353,N_10318);
xnor U11913 (N_11913,N_9170,N_10074);
nor U11914 (N_11914,N_9973,N_9240);
and U11915 (N_11915,N_9141,N_9224);
nor U11916 (N_11916,N_9484,N_10323);
nor U11917 (N_11917,N_9056,N_10393);
nor U11918 (N_11918,N_9738,N_9189);
nand U11919 (N_11919,N_10170,N_9406);
or U11920 (N_11920,N_9225,N_10448);
and U11921 (N_11921,N_10410,N_10291);
and U11922 (N_11922,N_9193,N_10051);
and U11923 (N_11923,N_9687,N_10317);
nor U11924 (N_11924,N_9528,N_9500);
nor U11925 (N_11925,N_9959,N_10140);
nand U11926 (N_11926,N_9276,N_10267);
nor U11927 (N_11927,N_9541,N_9830);
nand U11928 (N_11928,N_9008,N_9311);
nor U11929 (N_11929,N_9909,N_10082);
nand U11930 (N_11930,N_9210,N_9784);
or U11931 (N_11931,N_9378,N_9598);
nor U11932 (N_11932,N_9048,N_9615);
xor U11933 (N_11933,N_9112,N_9128);
nand U11934 (N_11934,N_9866,N_9341);
nand U11935 (N_11935,N_9754,N_10228);
nand U11936 (N_11936,N_9563,N_9293);
nor U11937 (N_11937,N_9058,N_9338);
nor U11938 (N_11938,N_9650,N_9017);
and U11939 (N_11939,N_10245,N_9211);
nand U11940 (N_11940,N_10326,N_9912);
or U11941 (N_11941,N_9789,N_9790);
nor U11942 (N_11942,N_10379,N_9953);
and U11943 (N_11943,N_10193,N_9779);
and U11944 (N_11944,N_9891,N_9811);
nor U11945 (N_11945,N_9554,N_9600);
xnor U11946 (N_11946,N_9894,N_10296);
nor U11947 (N_11947,N_9753,N_9743);
nand U11948 (N_11948,N_9816,N_10310);
or U11949 (N_11949,N_9732,N_9145);
xnor U11950 (N_11950,N_9237,N_10417);
nor U11951 (N_11951,N_9914,N_9950);
nor U11952 (N_11952,N_9215,N_9126);
nand U11953 (N_11953,N_9433,N_9041);
xor U11954 (N_11954,N_9104,N_9513);
and U11955 (N_11955,N_9319,N_9795);
or U11956 (N_11956,N_9141,N_9470);
nand U11957 (N_11957,N_9146,N_10336);
and U11958 (N_11958,N_9693,N_9306);
xor U11959 (N_11959,N_10109,N_9630);
nand U11960 (N_11960,N_9866,N_9376);
nand U11961 (N_11961,N_9036,N_9786);
nor U11962 (N_11962,N_9283,N_10014);
nand U11963 (N_11963,N_9758,N_9067);
or U11964 (N_11964,N_10477,N_10302);
and U11965 (N_11965,N_9284,N_10136);
or U11966 (N_11966,N_9495,N_10223);
and U11967 (N_11967,N_10473,N_10060);
or U11968 (N_11968,N_9195,N_9456);
and U11969 (N_11969,N_9082,N_9747);
nand U11970 (N_11970,N_10347,N_10446);
or U11971 (N_11971,N_10114,N_9911);
nor U11972 (N_11972,N_10348,N_9055);
nor U11973 (N_11973,N_10342,N_10329);
or U11974 (N_11974,N_9503,N_9092);
nor U11975 (N_11975,N_9090,N_9830);
nor U11976 (N_11976,N_9950,N_10312);
or U11977 (N_11977,N_9327,N_9737);
nand U11978 (N_11978,N_9988,N_9089);
xor U11979 (N_11979,N_9659,N_10200);
or U11980 (N_11980,N_9798,N_9318);
or U11981 (N_11981,N_9882,N_9447);
or U11982 (N_11982,N_9950,N_10325);
and U11983 (N_11983,N_9856,N_9976);
nand U11984 (N_11984,N_10218,N_10084);
or U11985 (N_11985,N_9711,N_10292);
xor U11986 (N_11986,N_9535,N_9328);
and U11987 (N_11987,N_9176,N_10117);
and U11988 (N_11988,N_9426,N_9047);
xnor U11989 (N_11989,N_9641,N_9475);
nor U11990 (N_11990,N_10183,N_10097);
and U11991 (N_11991,N_9069,N_9545);
or U11992 (N_11992,N_10151,N_9431);
xor U11993 (N_11993,N_9848,N_9880);
nor U11994 (N_11994,N_9527,N_9998);
nand U11995 (N_11995,N_9997,N_9454);
and U11996 (N_11996,N_10309,N_9134);
xnor U11997 (N_11997,N_9437,N_9995);
nor U11998 (N_11998,N_9645,N_9878);
nand U11999 (N_11999,N_9073,N_10389);
or U12000 (N_12000,N_11231,N_10872);
nor U12001 (N_12001,N_11431,N_11025);
and U12002 (N_12002,N_11796,N_11126);
nand U12003 (N_12003,N_10887,N_11228);
or U12004 (N_12004,N_10953,N_10636);
and U12005 (N_12005,N_11168,N_11605);
nor U12006 (N_12006,N_11562,N_11744);
and U12007 (N_12007,N_10974,N_11230);
xnor U12008 (N_12008,N_11476,N_11805);
nand U12009 (N_12009,N_11650,N_11935);
nor U12010 (N_12010,N_11814,N_11586);
and U12011 (N_12011,N_11189,N_11350);
xnor U12012 (N_12012,N_10770,N_11873);
and U12013 (N_12013,N_11296,N_11089);
xnor U12014 (N_12014,N_11149,N_11694);
nor U12015 (N_12015,N_11234,N_11898);
and U12016 (N_12016,N_11250,N_11018);
xor U12017 (N_12017,N_11278,N_11647);
nor U12018 (N_12018,N_11836,N_11968);
xnor U12019 (N_12019,N_11897,N_10731);
nand U12020 (N_12020,N_10534,N_11566);
or U12021 (N_12021,N_11884,N_11090);
nand U12022 (N_12022,N_11901,N_11116);
nor U12023 (N_12023,N_11499,N_11298);
xnor U12024 (N_12024,N_10748,N_11014);
xor U12025 (N_12025,N_10524,N_10620);
and U12026 (N_12026,N_10564,N_11715);
nand U12027 (N_12027,N_11921,N_11141);
nand U12028 (N_12028,N_10734,N_11057);
or U12029 (N_12029,N_11672,N_10909);
nor U12030 (N_12030,N_11508,N_10836);
nor U12031 (N_12031,N_11438,N_11464);
and U12032 (N_12032,N_11105,N_11345);
or U12033 (N_12033,N_11415,N_11594);
xor U12034 (N_12034,N_11505,N_11076);
or U12035 (N_12035,N_11319,N_10581);
and U12036 (N_12036,N_10789,N_10772);
or U12037 (N_12037,N_10787,N_11035);
and U12038 (N_12038,N_11943,N_11385);
nor U12039 (N_12039,N_11946,N_10604);
nor U12040 (N_12040,N_11860,N_11172);
nand U12041 (N_12041,N_10759,N_11227);
and U12042 (N_12042,N_11434,N_10739);
nor U12043 (N_12043,N_11933,N_11569);
or U12044 (N_12044,N_11810,N_11367);
nor U12045 (N_12045,N_10784,N_11161);
or U12046 (N_12046,N_11100,N_11206);
xor U12047 (N_12047,N_11140,N_11045);
or U12048 (N_12048,N_11176,N_10624);
nor U12049 (N_12049,N_10967,N_11005);
or U12050 (N_12050,N_11478,N_11584);
nand U12051 (N_12051,N_11770,N_10705);
nand U12052 (N_12052,N_10573,N_10845);
or U12053 (N_12053,N_10990,N_11288);
nand U12054 (N_12054,N_11396,N_10584);
xor U12055 (N_12055,N_11155,N_10950);
and U12056 (N_12056,N_11371,N_11775);
xor U12057 (N_12057,N_11183,N_10798);
nor U12058 (N_12058,N_10861,N_11754);
and U12059 (N_12059,N_10969,N_10778);
and U12060 (N_12060,N_10569,N_10609);
nor U12061 (N_12061,N_11244,N_10767);
and U12062 (N_12062,N_11877,N_11497);
nand U12063 (N_12063,N_11443,N_11670);
nand U12064 (N_12064,N_10886,N_11555);
xnor U12065 (N_12065,N_10833,N_11620);
and U12066 (N_12066,N_11633,N_10648);
nand U12067 (N_12067,N_11286,N_10780);
or U12068 (N_12068,N_11147,N_11993);
and U12069 (N_12069,N_10629,N_11614);
or U12070 (N_12070,N_10781,N_11047);
nand U12071 (N_12071,N_11980,N_10782);
or U12072 (N_12072,N_11468,N_10677);
nand U12073 (N_12073,N_10854,N_10832);
xnor U12074 (N_12074,N_11655,N_11695);
and U12075 (N_12075,N_11195,N_11406);
nor U12076 (N_12076,N_11626,N_11440);
and U12077 (N_12077,N_11861,N_11124);
xnor U12078 (N_12078,N_11779,N_11202);
nand U12079 (N_12079,N_10575,N_11737);
nand U12080 (N_12080,N_11846,N_10560);
and U12081 (N_12081,N_10699,N_11556);
nor U12082 (N_12082,N_11920,N_11848);
or U12083 (N_12083,N_11346,N_11245);
nand U12084 (N_12084,N_11200,N_11144);
and U12085 (N_12085,N_11341,N_11524);
and U12086 (N_12086,N_10906,N_11673);
nand U12087 (N_12087,N_11482,N_10571);
nor U12088 (N_12088,N_11241,N_11099);
or U12089 (N_12089,N_11996,N_11173);
nand U12090 (N_12090,N_11948,N_10709);
xnor U12091 (N_12091,N_10725,N_10991);
xnor U12092 (N_12092,N_10915,N_11021);
xnor U12093 (N_12093,N_10639,N_10989);
nand U12094 (N_12094,N_10727,N_10779);
nand U12095 (N_12095,N_11030,N_11764);
nand U12096 (N_12096,N_11666,N_10650);
or U12097 (N_12097,N_11563,N_11617);
nand U12098 (N_12098,N_11882,N_11447);
and U12099 (N_12099,N_11128,N_10985);
and U12100 (N_12100,N_11553,N_11326);
xor U12101 (N_12101,N_11711,N_10970);
xnor U12102 (N_12102,N_10956,N_11171);
nand U12103 (N_12103,N_11889,N_10519);
xnor U12104 (N_12104,N_10557,N_10755);
nor U12105 (N_12105,N_11780,N_11928);
nand U12106 (N_12106,N_11034,N_10653);
xnor U12107 (N_12107,N_11874,N_11693);
and U12108 (N_12108,N_10714,N_11940);
and U12109 (N_12109,N_11668,N_11747);
and U12110 (N_12110,N_11749,N_10976);
and U12111 (N_12111,N_10592,N_11890);
nand U12112 (N_12112,N_11932,N_11104);
nor U12113 (N_12113,N_10535,N_11062);
or U12114 (N_12114,N_10599,N_11334);
or U12115 (N_12115,N_11040,N_11262);
and U12116 (N_12116,N_10687,N_10975);
and U12117 (N_12117,N_10747,N_11287);
xnor U12118 (N_12118,N_11274,N_10914);
nand U12119 (N_12119,N_11409,N_11221);
nor U12120 (N_12120,N_11959,N_11750);
and U12121 (N_12121,N_11652,N_10590);
or U12122 (N_12122,N_11109,N_11813);
xor U12123 (N_12123,N_11857,N_10785);
or U12124 (N_12124,N_11769,N_10550);
nand U12125 (N_12125,N_10753,N_11284);
xor U12126 (N_12126,N_11953,N_11645);
nor U12127 (N_12127,N_11981,N_11625);
xor U12128 (N_12128,N_10695,N_11131);
nor U12129 (N_12129,N_11280,N_11448);
xor U12130 (N_12130,N_11748,N_11259);
or U12131 (N_12131,N_10948,N_10683);
and U12132 (N_12132,N_11717,N_10822);
nor U12133 (N_12133,N_11338,N_10882);
nor U12134 (N_12134,N_10973,N_10533);
and U12135 (N_12135,N_11362,N_11190);
nor U12136 (N_12136,N_11597,N_11085);
or U12137 (N_12137,N_11060,N_11847);
nor U12138 (N_12138,N_10506,N_10566);
or U12139 (N_12139,N_10972,N_11979);
and U12140 (N_12140,N_11480,N_11222);
nor U12141 (N_12141,N_11707,N_11546);
xor U12142 (N_12142,N_11927,N_11947);
and U12143 (N_12143,N_11148,N_11308);
xor U12144 (N_12144,N_11488,N_11723);
nor U12145 (N_12145,N_11379,N_10978);
xor U12146 (N_12146,N_10844,N_11667);
or U12147 (N_12147,N_11533,N_11500);
nand U12148 (N_12148,N_11636,N_11321);
nand U12149 (N_12149,N_10689,N_11971);
nand U12150 (N_12150,N_11268,N_11427);
and U12151 (N_12151,N_11213,N_10589);
xnor U12152 (N_12152,N_11355,N_11054);
xnor U12153 (N_12153,N_10513,N_10823);
nand U12154 (N_12154,N_10966,N_11318);
nand U12155 (N_12155,N_10563,N_10987);
xor U12156 (N_12156,N_11013,N_11094);
xor U12157 (N_12157,N_11194,N_10863);
xnor U12158 (N_12158,N_11329,N_10723);
or U12159 (N_12159,N_11201,N_10955);
nand U12160 (N_12160,N_11960,N_11470);
nand U12161 (N_12161,N_11519,N_10512);
and U12162 (N_12162,N_10543,N_10527);
nor U12163 (N_12163,N_11984,N_11938);
or U12164 (N_12164,N_11604,N_11905);
xor U12165 (N_12165,N_11640,N_11511);
nand U12166 (N_12166,N_11618,N_11530);
nor U12167 (N_12167,N_10879,N_11998);
xor U12168 (N_12168,N_11179,N_11619);
nor U12169 (N_12169,N_10889,N_10595);
and U12170 (N_12170,N_11883,N_11070);
or U12171 (N_12171,N_11079,N_10913);
nand U12172 (N_12172,N_10858,N_11380);
or U12173 (N_12173,N_10711,N_11224);
or U12174 (N_12174,N_10774,N_10801);
nor U12175 (N_12175,N_11044,N_11106);
nor U12176 (N_12176,N_10792,N_11364);
nand U12177 (N_12177,N_11212,N_11314);
nor U12178 (N_12178,N_11657,N_11292);
nor U12179 (N_12179,N_11487,N_11247);
nand U12180 (N_12180,N_10530,N_10936);
nor U12181 (N_12181,N_11559,N_11554);
xnor U12182 (N_12182,N_11075,N_10610);
or U12183 (N_12183,N_10971,N_11065);
nand U12184 (N_12184,N_10529,N_11637);
and U12185 (N_12185,N_11606,N_11359);
and U12186 (N_12186,N_11610,N_10795);
and U12187 (N_12187,N_11229,N_11537);
and U12188 (N_12188,N_10540,N_11127);
or U12189 (N_12189,N_11714,N_10875);
nand U12190 (N_12190,N_10605,N_10596);
nand U12191 (N_12191,N_10908,N_11818);
and U12192 (N_12192,N_10791,N_10911);
nor U12193 (N_12193,N_11356,N_10883);
and U12194 (N_12194,N_11773,N_11370);
nand U12195 (N_12195,N_11452,N_11630);
or U12196 (N_12196,N_10958,N_10903);
and U12197 (N_12197,N_11022,N_10657);
nor U12198 (N_12198,N_10598,N_11365);
nand U12199 (N_12199,N_11387,N_10600);
xnor U12200 (N_12200,N_11215,N_11774);
nand U12201 (N_12201,N_10752,N_11139);
and U12202 (N_12202,N_10613,N_10904);
nor U12203 (N_12203,N_10665,N_11941);
xor U12204 (N_12204,N_11975,N_10902);
nand U12205 (N_12205,N_10864,N_11395);
or U12206 (N_12206,N_11899,N_11491);
nand U12207 (N_12207,N_11567,N_11097);
nand U12208 (N_12208,N_11677,N_11002);
nand U12209 (N_12209,N_11969,N_11801);
nand U12210 (N_12210,N_11523,N_10988);
and U12211 (N_12211,N_11320,N_10635);
xnor U12212 (N_12212,N_11248,N_11307);
or U12213 (N_12213,N_11674,N_11735);
nand U12214 (N_12214,N_11990,N_11242);
nor U12215 (N_12215,N_10541,N_10628);
and U12216 (N_12216,N_11428,N_11407);
or U12217 (N_12217,N_11669,N_11392);
xnor U12218 (N_12218,N_10706,N_11738);
and U12219 (N_12219,N_11421,N_10814);
and U12220 (N_12220,N_11337,N_11028);
xor U12221 (N_12221,N_11671,N_11059);
and U12222 (N_12222,N_11624,N_11797);
xnor U12223 (N_12223,N_11056,N_11023);
nand U12224 (N_12224,N_11285,N_10831);
and U12225 (N_12225,N_11820,N_10995);
nor U12226 (N_12226,N_11143,N_11454);
and U12227 (N_12227,N_11725,N_11513);
xnor U12228 (N_12228,N_11203,N_11474);
xor U12229 (N_12229,N_10926,N_11378);
nor U12230 (N_12230,N_11120,N_10675);
and U12231 (N_12231,N_11015,N_10796);
nand U12232 (N_12232,N_11880,N_11217);
nor U12233 (N_12233,N_11053,N_11261);
or U12234 (N_12234,N_10996,N_11084);
xor U12235 (N_12235,N_11269,N_10673);
xor U12236 (N_12236,N_10521,N_10894);
or U12237 (N_12237,N_11507,N_11289);
nor U12238 (N_12238,N_11302,N_10511);
xor U12239 (N_12239,N_10503,N_10878);
and U12240 (N_12240,N_11441,N_11628);
nand U12241 (N_12241,N_10749,N_11974);
xnor U12242 (N_12242,N_11728,N_11449);
nor U12243 (N_12243,N_10952,N_10729);
or U12244 (N_12244,N_11697,N_11265);
nand U12245 (N_12245,N_11542,N_11658);
or U12246 (N_12246,N_11483,N_11389);
xor U12247 (N_12247,N_10551,N_11003);
nand U12248 (N_12248,N_11082,N_10686);
or U12249 (N_12249,N_10777,N_10855);
xnor U12250 (N_12250,N_10680,N_11829);
or U12251 (N_12251,N_11032,N_10884);
nand U12252 (N_12252,N_11133,N_11756);
and U12253 (N_12253,N_10984,N_11914);
nand U12254 (N_12254,N_11540,N_10502);
and U12255 (N_12255,N_10807,N_10678);
xor U12256 (N_12256,N_11486,N_10559);
and U12257 (N_12257,N_11757,N_10642);
xor U12258 (N_12258,N_11646,N_11574);
and U12259 (N_12259,N_11220,N_10745);
nand U12260 (N_12260,N_11664,N_11623);
and U12261 (N_12261,N_11451,N_11130);
and U12262 (N_12262,N_10769,N_10916);
nand U12263 (N_12263,N_11967,N_11167);
or U12264 (N_12264,N_11521,N_10580);
nand U12265 (N_12265,N_11453,N_10800);
nand U12266 (N_12266,N_11855,N_11595);
and U12267 (N_12267,N_11180,N_11550);
and U12268 (N_12268,N_11408,N_10700);
nand U12269 (N_12269,N_11039,N_11216);
or U12270 (N_12270,N_11635,N_11575);
nor U12271 (N_12271,N_11322,N_11985);
and U12272 (N_12272,N_11659,N_11276);
nor U12273 (N_12273,N_10603,N_10582);
nand U12274 (N_12274,N_10640,N_11510);
nor U12275 (N_12275,N_11751,N_10799);
and U12276 (N_12276,N_11119,N_10641);
nand U12277 (N_12277,N_11209,N_11459);
and U12278 (N_12278,N_11484,N_10572);
or U12279 (N_12279,N_10773,N_10834);
nor U12280 (N_12280,N_11323,N_10929);
and U12281 (N_12281,N_11924,N_10962);
and U12282 (N_12282,N_11436,N_11893);
xnor U12283 (N_12283,N_11724,N_11509);
and U12284 (N_12284,N_11410,N_10842);
xor U12285 (N_12285,N_11405,N_10998);
xor U12286 (N_12286,N_11174,N_11376);
and U12287 (N_12287,N_10556,N_11954);
and U12288 (N_12288,N_11918,N_11534);
nor U12289 (N_12289,N_11598,N_11976);
xnor U12290 (N_12290,N_11786,N_11989);
nand U12291 (N_12291,N_11926,N_10744);
nand U12292 (N_12292,N_11351,N_10611);
and U12293 (N_12293,N_11742,N_10786);
xor U12294 (N_12294,N_10539,N_10910);
or U12295 (N_12295,N_11834,N_11781);
nor U12296 (N_12296,N_11856,N_10715);
and U12297 (N_12297,N_10549,N_11049);
nor U12298 (N_12298,N_11762,N_10632);
nor U12299 (N_12299,N_10526,N_11547);
or U12300 (N_12300,N_10586,N_11184);
and U12301 (N_12301,N_11822,N_11461);
nand U12302 (N_12302,N_11311,N_11923);
nor U12303 (N_12303,N_11493,N_11435);
or U12304 (N_12304,N_10552,N_11166);
or U12305 (N_12305,N_11029,N_11279);
or U12306 (N_12306,N_10713,N_11214);
xor U12307 (N_12307,N_11886,N_10824);
nand U12308 (N_12308,N_11473,N_11732);
nor U12309 (N_12309,N_11275,N_11688);
and U12310 (N_12310,N_11768,N_11821);
and U12311 (N_12311,N_11479,N_10664);
nand U12312 (N_12312,N_11577,N_11456);
or U12313 (N_12313,N_11251,N_11024);
xor U12314 (N_12314,N_10757,N_11186);
and U12315 (N_12315,N_10803,N_11064);
xor U12316 (N_12316,N_11541,N_11680);
xor U12317 (N_12317,N_10579,N_10758);
or U12318 (N_12318,N_11336,N_11026);
xor U12319 (N_12319,N_11072,N_11807);
nor U12320 (N_12320,N_10827,N_10923);
and U12321 (N_12321,N_11613,N_10718);
xor U12322 (N_12322,N_11368,N_11369);
and U12323 (N_12323,N_11420,N_11360);
xor U12324 (N_12324,N_11503,N_10776);
or U12325 (N_12325,N_11593,N_11504);
nor U12326 (N_12326,N_11066,N_11578);
xnor U12327 (N_12327,N_11506,N_10558);
xor U12328 (N_12328,N_11687,N_11226);
and U12329 (N_12329,N_11357,N_10587);
nand U12330 (N_12330,N_11611,N_10965);
xnor U12331 (N_12331,N_11588,N_11086);
nand U12332 (N_12332,N_10652,N_11766);
and U12333 (N_12333,N_11839,N_11293);
and U12334 (N_12334,N_10726,N_11239);
and U12335 (N_12335,N_11381,N_10930);
nor U12336 (N_12336,N_11718,N_11632);
nor U12337 (N_12337,N_11243,N_10655);
and U12338 (N_12338,N_10743,N_10514);
nor U12339 (N_12339,N_10765,N_11403);
or U12340 (N_12340,N_10545,N_10574);
nor U12341 (N_12341,N_10746,N_10577);
nor U12342 (N_12342,N_11397,N_10934);
nand U12343 (N_12343,N_10829,N_11008);
xor U12344 (N_12344,N_10896,N_11570);
and U12345 (N_12345,N_11587,N_10666);
or U12346 (N_12346,N_11910,N_10616);
xor U12347 (N_12347,N_10736,N_11412);
nor U12348 (N_12348,N_11661,N_11612);
or U12349 (N_12349,N_10907,N_10835);
or U12350 (N_12350,N_11437,N_10501);
xor U12351 (N_12351,N_11763,N_11518);
nand U12352 (N_12352,N_11722,N_11363);
or U12353 (N_12353,N_10555,N_10703);
xnor U12354 (N_12354,N_11837,N_11665);
nor U12355 (N_12355,N_10704,N_11160);
or U12356 (N_12356,N_11529,N_11375);
nand U12357 (N_12357,N_10670,N_11970);
and U12358 (N_12358,N_10638,N_11930);
or U12359 (N_12359,N_11912,N_11581);
nor U12360 (N_12360,N_11414,N_11755);
nand U12361 (N_12361,N_11061,N_10523);
nor U12362 (N_12362,N_11372,N_11142);
nor U12363 (N_12363,N_11073,N_11411);
nor U12364 (N_12364,N_11966,N_11867);
nor U12365 (N_12365,N_11048,N_11467);
nor U12366 (N_12366,N_11153,N_11398);
nand U12367 (N_12367,N_11445,N_10818);
xnor U12368 (N_12368,N_10721,N_11418);
nand U12369 (N_12369,N_11643,N_10669);
xnor U12370 (N_12370,N_11599,N_10672);
and U12371 (N_12371,N_10717,N_11739);
nor U12372 (N_12372,N_11016,N_10849);
or U12373 (N_12373,N_10510,N_11549);
or U12374 (N_12374,N_11299,N_10805);
nand U12375 (N_12375,N_10869,N_11696);
xnor U12376 (N_12376,N_11425,N_11639);
xor U12377 (N_12377,N_10701,N_10623);
or U12378 (N_12378,N_11169,N_10821);
or U12379 (N_12379,N_10698,N_11263);
xnor U12380 (N_12380,N_11908,N_10917);
or U12381 (N_12381,N_11423,N_11961);
or U12382 (N_12382,N_11791,N_11713);
nand U12383 (N_12383,N_11006,N_11151);
or U12384 (N_12384,N_10728,N_11907);
and U12385 (N_12385,N_11330,N_11041);
nand U12386 (N_12386,N_11621,N_11616);
nand U12387 (N_12387,N_10959,N_11733);
nand U12388 (N_12388,N_11760,N_11827);
nand U12389 (N_12389,N_10820,N_10994);
and U12390 (N_12390,N_11600,N_10977);
xnor U12391 (N_12391,N_11734,N_11038);
xor U12392 (N_12392,N_11706,N_11838);
and U12393 (N_12393,N_11548,N_11798);
xor U12394 (N_12394,N_10614,N_11007);
or U12395 (N_12395,N_11701,N_10839);
nor U12396 (N_12396,N_11878,N_10515);
and U12397 (N_12397,N_10576,N_10671);
nand U12398 (N_12398,N_10895,N_11352);
and U12399 (N_12399,N_10602,N_11753);
nand U12400 (N_12400,N_10750,N_10964);
xor U12401 (N_12401,N_11196,N_11283);
or U12402 (N_12402,N_11936,N_11746);
or U12403 (N_12403,N_11137,N_11324);
and U12404 (N_12404,N_11477,N_11156);
nor U12405 (N_12405,N_11875,N_11651);
nor U12406 (N_12406,N_11433,N_10509);
and U12407 (N_12407,N_11122,N_11349);
xor U12408 (N_12408,N_11102,N_11784);
nand U12409 (N_12409,N_11913,N_10618);
xnor U12410 (N_12410,N_11152,N_11977);
and U12411 (N_12411,N_11642,N_10740);
or U12412 (N_12412,N_10825,N_11270);
nor U12413 (N_12413,N_11121,N_11896);
nand U12414 (N_12414,N_10817,N_10627);
and U12415 (N_12415,N_11656,N_11281);
and U12416 (N_12416,N_10681,N_11863);
nor U12417 (N_12417,N_11291,N_10856);
nor U12418 (N_12418,N_10591,N_11799);
and U12419 (N_12419,N_11009,N_10848);
nand U12420 (N_12420,N_11193,N_10897);
xor U12421 (N_12421,N_11917,N_10500);
nor U12422 (N_12422,N_11675,N_11726);
or U12423 (N_12423,N_10522,N_10583);
and U12424 (N_12424,N_10871,N_11973);
or U12425 (N_12425,N_10568,N_11700);
or U12426 (N_12426,N_11450,N_11851);
nor U12427 (N_12427,N_11986,N_11388);
xor U12428 (N_12428,N_11809,N_11267);
nand U12429 (N_12429,N_11660,N_10763);
or U12430 (N_12430,N_11096,N_10925);
nand U12431 (N_12431,N_11017,N_11699);
and U12432 (N_12432,N_10517,N_11223);
and U12433 (N_12433,N_11854,N_11939);
nand U12434 (N_12434,N_10532,N_11178);
nor U12435 (N_12435,N_11934,N_11498);
or U12436 (N_12436,N_11042,N_11512);
nand U12437 (N_12437,N_11295,N_11835);
nor U12438 (N_12438,N_10935,N_11561);
nand U12439 (N_12439,N_11629,N_11489);
and U12440 (N_12440,N_11788,N_10608);
xor U12441 (N_12441,N_11424,N_11374);
nand U12442 (N_12442,N_11911,N_10567);
nor U12443 (N_12443,N_11138,N_10853);
or U12444 (N_12444,N_11958,N_11782);
nand U12445 (N_12445,N_11937,N_10830);
and U12446 (N_12446,N_10860,N_10708);
xnor U12447 (N_12447,N_11390,N_11125);
nand U12448 (N_12448,N_10943,N_11771);
xor U12449 (N_12449,N_11163,N_10813);
nor U12450 (N_12450,N_10697,N_10667);
nand U12451 (N_12451,N_11870,N_11343);
nor U12452 (N_12452,N_10730,N_11956);
nand U12453 (N_12453,N_11852,N_11087);
nor U12454 (N_12454,N_11585,N_10643);
and U12455 (N_12455,N_11806,N_10901);
xor U12456 (N_12456,N_10561,N_11310);
nand U12457 (N_12457,N_10866,N_11686);
or U12458 (N_12458,N_11532,N_11078);
and U12459 (N_12459,N_11384,N_10660);
nor U12460 (N_12460,N_10986,N_11853);
and U12461 (N_12461,N_11526,N_11945);
and U12462 (N_12462,N_10644,N_11134);
nor U12463 (N_12463,N_11145,N_10797);
and U12464 (N_12464,N_11068,N_10979);
or U12465 (N_12465,N_11010,N_11466);
or U12466 (N_12466,N_10742,N_11313);
nand U12467 (N_12467,N_11260,N_11536);
and U12468 (N_12468,N_11012,N_10649);
nor U12469 (N_12469,N_11793,N_11649);
nor U12470 (N_12470,N_10954,N_11634);
and U12471 (N_12471,N_11601,N_10615);
xor U12472 (N_12472,N_10659,N_10508);
nor U12473 (N_12473,N_10651,N_11290);
and U12474 (N_12474,N_11312,N_11638);
xor U12475 (N_12475,N_11074,N_10597);
or U12476 (N_12476,N_10656,N_11077);
and U12477 (N_12477,N_10867,N_11164);
nand U12478 (N_12478,N_11582,N_11849);
and U12479 (N_12479,N_11790,N_11787);
nand U12480 (N_12480,N_11386,N_10585);
or U12481 (N_12481,N_11492,N_11783);
and U12482 (N_12482,N_11465,N_11462);
nor U12483 (N_12483,N_11182,N_11277);
nand U12484 (N_12484,N_11864,N_11271);
nor U12485 (N_12485,N_10946,N_11903);
and U12486 (N_12486,N_11309,N_11811);
or U12487 (N_12487,N_10525,N_11915);
or U12488 (N_12488,N_11922,N_11394);
or U12489 (N_12489,N_11112,N_10963);
nor U12490 (N_12490,N_11894,N_11900);
xor U12491 (N_12491,N_11995,N_11758);
nor U12492 (N_12492,N_10981,N_10809);
nand U12493 (N_12493,N_11545,N_11929);
nand U12494 (N_12494,N_11335,N_11705);
or U12495 (N_12495,N_11716,N_11020);
xnor U12496 (N_12496,N_11063,N_11676);
and U12497 (N_12497,N_11111,N_10768);
nor U12498 (N_12498,N_11218,N_10528);
nor U12499 (N_12499,N_11342,N_11273);
or U12500 (N_12500,N_10548,N_10949);
or U12501 (N_12501,N_11490,N_11955);
nor U12502 (N_12502,N_10815,N_11794);
nor U12503 (N_12503,N_11093,N_11430);
nand U12504 (N_12504,N_11358,N_10588);
xor U12505 (N_12505,N_11515,N_11475);
nand U12506 (N_12506,N_11992,N_11957);
or U12507 (N_12507,N_10601,N_11303);
or U12508 (N_12508,N_11058,N_11816);
nand U12509 (N_12509,N_11383,N_10980);
xor U12510 (N_12510,N_10951,N_11727);
xor U12511 (N_12511,N_11108,N_11501);
and U12512 (N_12512,N_11238,N_10928);
or U12513 (N_12513,N_11817,N_11983);
and U12514 (N_12514,N_10852,N_11256);
and U12515 (N_12515,N_11327,N_10612);
nor U12516 (N_12516,N_11869,N_11107);
xor U12517 (N_12517,N_10788,N_11804);
nand U12518 (N_12518,N_11177,N_11257);
and U12519 (N_12519,N_10668,N_11404);
nor U12520 (N_12520,N_11573,N_10968);
or U12521 (N_12521,N_10812,N_11564);
or U12522 (N_12522,N_11157,N_11181);
nand U12523 (N_12523,N_10536,N_11580);
nor U12524 (N_12524,N_11426,N_10937);
nor U12525 (N_12525,N_10982,N_10637);
nand U12526 (N_12526,N_10507,N_11951);
or U12527 (N_12527,N_11833,N_10870);
nand U12528 (N_12528,N_11495,N_11046);
or U12529 (N_12529,N_10735,N_11158);
nand U12530 (N_12530,N_10881,N_11252);
or U12531 (N_12531,N_11906,N_10868);
or U12532 (N_12532,N_10537,N_11683);
and U12533 (N_12533,N_11027,N_11712);
nand U12534 (N_12534,N_10793,N_11325);
nor U12535 (N_12535,N_10716,N_11653);
xor U12536 (N_12536,N_11494,N_10760);
nor U12537 (N_12537,N_10762,N_11258);
and U12538 (N_12538,N_10947,N_11964);
nand U12539 (N_12539,N_11830,N_11233);
nand U12540 (N_12540,N_10684,N_10546);
nor U12541 (N_12541,N_10538,N_11463);
xor U12542 (N_12542,N_11778,N_11691);
nand U12543 (N_12543,N_10857,N_10693);
and U12544 (N_12544,N_10626,N_11795);
xnor U12545 (N_12545,N_10737,N_11871);
and U12546 (N_12546,N_11887,N_11709);
xor U12547 (N_12547,N_11997,N_11785);
xnor U12548 (N_12548,N_11069,N_10761);
nand U12549 (N_12549,N_11682,N_10764);
and U12550 (N_12550,N_10837,N_10544);
nand U12551 (N_12551,N_11333,N_10617);
nand U12552 (N_12552,N_11885,N_11496);
or U12553 (N_12553,N_11963,N_10846);
and U12554 (N_12554,N_10859,N_11347);
xnor U12555 (N_12555,N_10553,N_10920);
xnor U12556 (N_12556,N_10804,N_11842);
or U12557 (N_12557,N_11083,N_11031);
xnor U12558 (N_12558,N_11949,N_10808);
nand U12559 (N_12559,N_10927,N_11710);
nor U12560 (N_12560,N_10658,N_10775);
nand U12561 (N_12561,N_11592,N_10874);
and U12562 (N_12562,N_11191,N_11551);
nand U12563 (N_12563,N_11607,N_10766);
nor U12564 (N_12564,N_11353,N_11609);
and U12565 (N_12565,N_10806,N_11249);
nand U12566 (N_12566,N_10662,N_11051);
nor U12567 (N_12567,N_11824,N_11457);
and U12568 (N_12568,N_10520,N_11819);
nor U12569 (N_12569,N_11999,N_11132);
nand U12570 (N_12570,N_10933,N_10674);
or U12571 (N_12571,N_10783,N_11080);
xnor U12572 (N_12572,N_11001,N_10654);
or U12573 (N_12573,N_10819,N_10945);
nor U12574 (N_12574,N_10504,N_10547);
nor U12575 (N_12575,N_11568,N_11197);
nor U12576 (N_12576,N_11517,N_11469);
and U12577 (N_12577,N_11516,N_10692);
xor U12578 (N_12578,N_11088,N_11402);
nand U12579 (N_12579,N_11590,N_11055);
xor U12580 (N_12580,N_11123,N_11685);
xor U12581 (N_12581,N_11692,N_11232);
nand U12582 (N_12582,N_10924,N_11876);
or U12583 (N_12583,N_11684,N_10944);
nand U12584 (N_12584,N_10843,N_10724);
xor U12585 (N_12585,N_11815,N_11615);
and U12586 (N_12586,N_11340,N_11401);
or U12587 (N_12587,N_10905,N_10690);
xor U12588 (N_12588,N_10921,N_11208);
or U12589 (N_12589,N_11165,N_11067);
or U12590 (N_12590,N_11205,N_10594);
nor U12591 (N_12591,N_11422,N_11831);
xor U12592 (N_12592,N_11004,N_10802);
nand U12593 (N_12593,N_11731,N_11916);
and U12594 (N_12594,N_11520,N_10961);
and U12595 (N_12595,N_10992,N_11522);
nand U12596 (N_12596,N_11828,N_11098);
nand U12597 (N_12597,N_11419,N_11919);
and U12598 (N_12598,N_11019,N_10531);
or U12599 (N_12599,N_10661,N_11301);
nor U12600 (N_12600,N_11091,N_11662);
nand U12601 (N_12601,N_11572,N_10794);
nor U12602 (N_12602,N_11240,N_11527);
nand U12603 (N_12603,N_11825,N_11832);
nand U12604 (N_12604,N_10877,N_10719);
or U12605 (N_12605,N_10828,N_10873);
nand U12606 (N_12606,N_11845,N_10696);
nand U12607 (N_12607,N_10771,N_11136);
and U12608 (N_12608,N_10607,N_10516);
nor U12609 (N_12609,N_10505,N_11777);
or U12610 (N_12610,N_11235,N_10754);
nand U12611 (N_12611,N_11192,N_10518);
xor U12612 (N_12612,N_11879,N_11859);
nor U12613 (N_12613,N_11101,N_11344);
xor U12614 (N_12614,N_11339,N_11211);
nor U12615 (N_12615,N_11052,N_11439);
or U12616 (N_12616,N_11316,N_11865);
or U12617 (N_12617,N_11648,N_11972);
nand U12618 (N_12618,N_11502,N_11185);
and U12619 (N_12619,N_11095,N_10663);
and U12620 (N_12620,N_10741,N_11690);
and U12621 (N_12621,N_11952,N_11154);
xor U12622 (N_12622,N_10542,N_11987);
nor U12623 (N_12623,N_11862,N_11560);
nand U12624 (N_12624,N_11579,N_11317);
nand U12625 (N_12625,N_10679,N_10841);
or U12626 (N_12626,N_11354,N_11902);
xor U12627 (N_12627,N_11752,N_10810);
and U12628 (N_12628,N_11789,N_10562);
xnor U12629 (N_12629,N_11531,N_11366);
nor U12630 (N_12630,N_11033,N_10918);
or U12631 (N_12631,N_11219,N_11772);
and U12632 (N_12632,N_11942,N_11826);
nand U12633 (N_12633,N_10676,N_11071);
nand U12634 (N_12634,N_11382,N_11802);
or U12635 (N_12635,N_11565,N_11377);
or U12636 (N_12636,N_10622,N_11118);
xnor U12637 (N_12637,N_10922,N_11603);
nor U12638 (N_12638,N_10633,N_10941);
nor U12639 (N_12639,N_11442,N_10756);
nand U12640 (N_12640,N_11803,N_10912);
nand U12641 (N_12641,N_10646,N_10876);
or U12642 (N_12642,N_11622,N_11679);
or U12643 (N_12643,N_11162,N_11730);
nand U12644 (N_12644,N_11925,N_11300);
xor U12645 (N_12645,N_10862,N_11472);
or U12646 (N_12646,N_11708,N_11187);
nand U12647 (N_12647,N_11535,N_11294);
xor U12648 (N_12648,N_10625,N_11641);
nor U12649 (N_12649,N_10826,N_11866);
xor U12650 (N_12650,N_10865,N_11850);
or U12651 (N_12651,N_11543,N_10880);
and U12652 (N_12652,N_11800,N_10630);
nor U12653 (N_12653,N_11808,N_10751);
and U12654 (N_12654,N_11204,N_10645);
and U12655 (N_12655,N_11841,N_11332);
nor U12656 (N_12656,N_11305,N_11150);
nor U12657 (N_12657,N_11272,N_10631);
and U12658 (N_12658,N_11631,N_11868);
or U12659 (N_12659,N_11888,N_10957);
or U12660 (N_12660,N_11416,N_11114);
and U12661 (N_12661,N_10606,N_10983);
nor U12662 (N_12662,N_11931,N_11481);
xnor U12663 (N_12663,N_10940,N_11198);
and U12664 (N_12664,N_10720,N_11736);
nor U12665 (N_12665,N_10885,N_10847);
nand U12666 (N_12666,N_11978,N_10816);
xor U12667 (N_12667,N_11988,N_10712);
nor U12668 (N_12668,N_10634,N_11444);
xnor U12669 (N_12669,N_11282,N_11237);
nor U12670 (N_12670,N_11188,N_11199);
or U12671 (N_12671,N_11895,N_11602);
and U12672 (N_12672,N_11103,N_11589);
nand U12673 (N_12673,N_10932,N_11525);
and U12674 (N_12674,N_11721,N_10554);
or U12675 (N_12675,N_11654,N_11417);
or U12676 (N_12676,N_11429,N_10722);
nor U12677 (N_12677,N_11904,N_11225);
or U12678 (N_12678,N_10738,N_11663);
nand U12679 (N_12679,N_11236,N_11720);
or U12680 (N_12680,N_11740,N_11315);
nand U12681 (N_12681,N_11644,N_11891);
and U12682 (N_12682,N_10942,N_10931);
or U12683 (N_12683,N_11812,N_10891);
or U12684 (N_12684,N_11844,N_11348);
nor U12685 (N_12685,N_10997,N_11982);
and U12686 (N_12686,N_11254,N_11702);
or U12687 (N_12687,N_10899,N_10685);
nand U12688 (N_12688,N_11050,N_10898);
and U12689 (N_12689,N_11858,N_11117);
and U12690 (N_12690,N_11092,N_10688);
nor U12691 (N_12691,N_11965,N_11991);
nand U12692 (N_12692,N_11110,N_10593);
xor U12693 (N_12693,N_11792,N_11892);
xor U12694 (N_12694,N_11328,N_11264);
or U12695 (N_12695,N_11704,N_11460);
xnor U12696 (N_12696,N_11538,N_11011);
xnor U12697 (N_12697,N_11596,N_11331);
xor U12698 (N_12698,N_10850,N_10811);
nor U12699 (N_12699,N_11207,N_10694);
or U12700 (N_12700,N_11306,N_11297);
xor U12701 (N_12701,N_11761,N_11557);
nand U12702 (N_12702,N_11591,N_10893);
or U12703 (N_12703,N_10892,N_11391);
or U12704 (N_12704,N_11255,N_10732);
xor U12705 (N_12705,N_11266,N_11681);
nor U12706 (N_12706,N_10960,N_10919);
nand U12707 (N_12707,N_11246,N_11253);
or U12708 (N_12708,N_11729,N_11765);
xnor U12709 (N_12709,N_11571,N_11393);
nand U12710 (N_12710,N_11159,N_10570);
and U12711 (N_12711,N_11994,N_10707);
xor U12712 (N_12712,N_11944,N_11471);
and U12713 (N_12713,N_11608,N_11000);
nand U12714 (N_12714,N_11719,N_11135);
nor U12715 (N_12715,N_10938,N_11399);
nand U12716 (N_12716,N_11759,N_11146);
nand U12717 (N_12717,N_10702,N_11552);
or U12718 (N_12718,N_11843,N_11576);
xnor U12719 (N_12719,N_10838,N_10851);
nor U12720 (N_12720,N_11113,N_10790);
and U12721 (N_12721,N_11115,N_11458);
xor U12722 (N_12722,N_11745,N_10619);
and U12723 (N_12723,N_11909,N_10999);
nand U12724 (N_12724,N_11840,N_10647);
and U12725 (N_12725,N_11872,N_11304);
and U12726 (N_12726,N_10890,N_11036);
xnor U12727 (N_12727,N_10565,N_11776);
xor U12728 (N_12728,N_11703,N_10578);
or U12729 (N_12729,N_10733,N_10682);
nand U12730 (N_12730,N_11698,N_11823);
or U12731 (N_12731,N_10939,N_11361);
xor U12732 (N_12732,N_11170,N_11950);
nand U12733 (N_12733,N_11583,N_11558);
or U12734 (N_12734,N_11881,N_11175);
nand U12735 (N_12735,N_11485,N_11043);
and U12736 (N_12736,N_10710,N_10840);
and U12737 (N_12737,N_11743,N_11528);
xor U12738 (N_12738,N_11446,N_11962);
and U12739 (N_12739,N_11210,N_10888);
nand U12740 (N_12740,N_11037,N_10621);
or U12741 (N_12741,N_11081,N_11129);
nand U12742 (N_12742,N_11373,N_11539);
nor U12743 (N_12743,N_11400,N_11544);
xor U12744 (N_12744,N_10993,N_11741);
xnor U12745 (N_12745,N_11514,N_11767);
or U12746 (N_12746,N_11455,N_11413);
nand U12747 (N_12747,N_11689,N_11432);
xor U12748 (N_12748,N_10900,N_10691);
nand U12749 (N_12749,N_11627,N_11678);
nor U12750 (N_12750,N_10665,N_11842);
nand U12751 (N_12751,N_11162,N_11478);
xnor U12752 (N_12752,N_11822,N_11686);
and U12753 (N_12753,N_11547,N_11255);
or U12754 (N_12754,N_11956,N_11411);
xnor U12755 (N_12755,N_10860,N_11071);
and U12756 (N_12756,N_11093,N_10576);
and U12757 (N_12757,N_10684,N_10605);
and U12758 (N_12758,N_10635,N_11516);
or U12759 (N_12759,N_11165,N_10896);
and U12760 (N_12760,N_11553,N_10790);
xor U12761 (N_12761,N_11141,N_11155);
and U12762 (N_12762,N_11627,N_10686);
or U12763 (N_12763,N_11247,N_11097);
xnor U12764 (N_12764,N_11078,N_10742);
nand U12765 (N_12765,N_11546,N_10829);
or U12766 (N_12766,N_11125,N_10567);
or U12767 (N_12767,N_11302,N_11703);
nor U12768 (N_12768,N_10742,N_11211);
and U12769 (N_12769,N_11064,N_11686);
xnor U12770 (N_12770,N_10596,N_11891);
xor U12771 (N_12771,N_11243,N_11797);
and U12772 (N_12772,N_10589,N_11370);
xnor U12773 (N_12773,N_11364,N_10732);
nor U12774 (N_12774,N_10793,N_11928);
nand U12775 (N_12775,N_11612,N_10891);
and U12776 (N_12776,N_11381,N_11667);
xnor U12777 (N_12777,N_10760,N_11599);
nand U12778 (N_12778,N_11799,N_11666);
and U12779 (N_12779,N_11984,N_11913);
and U12780 (N_12780,N_10533,N_11729);
nand U12781 (N_12781,N_11725,N_11838);
xor U12782 (N_12782,N_11818,N_11166);
xnor U12783 (N_12783,N_11600,N_10577);
nor U12784 (N_12784,N_10883,N_10581);
nor U12785 (N_12785,N_11080,N_11773);
or U12786 (N_12786,N_10865,N_11344);
and U12787 (N_12787,N_11549,N_11332);
nand U12788 (N_12788,N_11333,N_11076);
or U12789 (N_12789,N_11611,N_11946);
nor U12790 (N_12790,N_10817,N_11941);
nor U12791 (N_12791,N_11688,N_10936);
nor U12792 (N_12792,N_11444,N_11068);
xnor U12793 (N_12793,N_10654,N_10945);
xnor U12794 (N_12794,N_10983,N_11804);
xor U12795 (N_12795,N_11596,N_10511);
or U12796 (N_12796,N_11843,N_10823);
or U12797 (N_12797,N_10508,N_11621);
xor U12798 (N_12798,N_11546,N_11272);
nand U12799 (N_12799,N_11577,N_11301);
nand U12800 (N_12800,N_11815,N_11991);
xnor U12801 (N_12801,N_11510,N_11161);
xor U12802 (N_12802,N_11484,N_11731);
nor U12803 (N_12803,N_11572,N_11986);
nor U12804 (N_12804,N_11412,N_11369);
nor U12805 (N_12805,N_11115,N_10526);
and U12806 (N_12806,N_11791,N_11583);
or U12807 (N_12807,N_11018,N_10681);
or U12808 (N_12808,N_10548,N_11909);
and U12809 (N_12809,N_11465,N_11764);
or U12810 (N_12810,N_11847,N_10785);
or U12811 (N_12811,N_11208,N_11501);
or U12812 (N_12812,N_11271,N_11244);
nand U12813 (N_12813,N_11989,N_11961);
nand U12814 (N_12814,N_11749,N_10677);
and U12815 (N_12815,N_11805,N_10807);
nand U12816 (N_12816,N_10805,N_10538);
nand U12817 (N_12817,N_11926,N_10751);
nand U12818 (N_12818,N_10684,N_10601);
nand U12819 (N_12819,N_10638,N_11266);
xor U12820 (N_12820,N_11319,N_11930);
or U12821 (N_12821,N_10947,N_11071);
nand U12822 (N_12822,N_11569,N_11703);
nor U12823 (N_12823,N_10731,N_10695);
and U12824 (N_12824,N_10669,N_11917);
or U12825 (N_12825,N_10859,N_11560);
nand U12826 (N_12826,N_11831,N_11869);
and U12827 (N_12827,N_10605,N_11916);
and U12828 (N_12828,N_11295,N_11865);
nor U12829 (N_12829,N_10811,N_11071);
and U12830 (N_12830,N_11480,N_10783);
and U12831 (N_12831,N_10560,N_11849);
xor U12832 (N_12832,N_11245,N_11475);
nor U12833 (N_12833,N_11497,N_11070);
and U12834 (N_12834,N_11887,N_10623);
and U12835 (N_12835,N_10621,N_10763);
nand U12836 (N_12836,N_11828,N_10938);
and U12837 (N_12837,N_10964,N_10968);
xnor U12838 (N_12838,N_11528,N_11888);
and U12839 (N_12839,N_10969,N_11556);
or U12840 (N_12840,N_11679,N_11652);
and U12841 (N_12841,N_11281,N_11151);
or U12842 (N_12842,N_11716,N_11293);
nor U12843 (N_12843,N_11866,N_11643);
or U12844 (N_12844,N_10640,N_10703);
and U12845 (N_12845,N_11562,N_11636);
nand U12846 (N_12846,N_10688,N_11894);
xor U12847 (N_12847,N_11645,N_11379);
or U12848 (N_12848,N_10543,N_11177);
nor U12849 (N_12849,N_11666,N_11989);
and U12850 (N_12850,N_10929,N_10593);
nor U12851 (N_12851,N_11800,N_11454);
or U12852 (N_12852,N_11333,N_11865);
nor U12853 (N_12853,N_11575,N_11269);
and U12854 (N_12854,N_11147,N_11004);
nand U12855 (N_12855,N_11870,N_10946);
and U12856 (N_12856,N_10881,N_10893);
nand U12857 (N_12857,N_11740,N_10855);
xnor U12858 (N_12858,N_11300,N_11561);
xnor U12859 (N_12859,N_11628,N_11800);
nand U12860 (N_12860,N_10769,N_11320);
or U12861 (N_12861,N_11157,N_11479);
nor U12862 (N_12862,N_11871,N_10577);
nor U12863 (N_12863,N_11181,N_10990);
xor U12864 (N_12864,N_10546,N_11616);
and U12865 (N_12865,N_11949,N_11571);
or U12866 (N_12866,N_11660,N_10895);
nor U12867 (N_12867,N_11657,N_11202);
nor U12868 (N_12868,N_11430,N_11284);
or U12869 (N_12869,N_11300,N_11135);
or U12870 (N_12870,N_11113,N_11074);
nor U12871 (N_12871,N_11599,N_10539);
nand U12872 (N_12872,N_11152,N_11485);
nand U12873 (N_12873,N_11486,N_10658);
nor U12874 (N_12874,N_11162,N_11743);
or U12875 (N_12875,N_11909,N_11846);
nand U12876 (N_12876,N_10941,N_11974);
xor U12877 (N_12877,N_11923,N_10777);
or U12878 (N_12878,N_10762,N_10712);
xnor U12879 (N_12879,N_10840,N_11048);
and U12880 (N_12880,N_11435,N_11617);
or U12881 (N_12881,N_11448,N_11799);
xnor U12882 (N_12882,N_11270,N_11681);
xor U12883 (N_12883,N_11336,N_10596);
and U12884 (N_12884,N_11819,N_10585);
nor U12885 (N_12885,N_10679,N_10769);
xor U12886 (N_12886,N_11009,N_10918);
nand U12887 (N_12887,N_11050,N_10978);
xnor U12888 (N_12888,N_10953,N_10693);
and U12889 (N_12889,N_11770,N_11086);
and U12890 (N_12890,N_11180,N_11472);
and U12891 (N_12891,N_11275,N_11093);
nand U12892 (N_12892,N_11700,N_11189);
xor U12893 (N_12893,N_10605,N_11662);
or U12894 (N_12894,N_10514,N_11390);
nand U12895 (N_12895,N_11407,N_11565);
or U12896 (N_12896,N_11462,N_11519);
or U12897 (N_12897,N_11951,N_11075);
xnor U12898 (N_12898,N_11596,N_11626);
nor U12899 (N_12899,N_11250,N_10914);
nand U12900 (N_12900,N_11408,N_11068);
or U12901 (N_12901,N_11364,N_11675);
nor U12902 (N_12902,N_11114,N_11909);
and U12903 (N_12903,N_11807,N_11163);
or U12904 (N_12904,N_11039,N_11893);
nand U12905 (N_12905,N_11550,N_10695);
and U12906 (N_12906,N_10801,N_10503);
nor U12907 (N_12907,N_11977,N_10683);
nand U12908 (N_12908,N_10560,N_11688);
and U12909 (N_12909,N_10837,N_10655);
nand U12910 (N_12910,N_11307,N_11460);
nand U12911 (N_12911,N_11299,N_11701);
xor U12912 (N_12912,N_10740,N_11869);
nor U12913 (N_12913,N_10767,N_11545);
or U12914 (N_12914,N_10585,N_11740);
or U12915 (N_12915,N_10974,N_10932);
xor U12916 (N_12916,N_11841,N_10619);
and U12917 (N_12917,N_10866,N_11009);
nand U12918 (N_12918,N_11936,N_11390);
nand U12919 (N_12919,N_11740,N_11348);
and U12920 (N_12920,N_11744,N_11108);
or U12921 (N_12921,N_11774,N_11169);
nor U12922 (N_12922,N_11112,N_11128);
nand U12923 (N_12923,N_11125,N_11265);
xnor U12924 (N_12924,N_10622,N_11284);
and U12925 (N_12925,N_11534,N_11925);
or U12926 (N_12926,N_10735,N_11094);
and U12927 (N_12927,N_11858,N_11086);
and U12928 (N_12928,N_11949,N_11516);
and U12929 (N_12929,N_11055,N_11659);
nand U12930 (N_12930,N_11651,N_11548);
or U12931 (N_12931,N_11620,N_11968);
or U12932 (N_12932,N_11256,N_10729);
or U12933 (N_12933,N_11032,N_11237);
or U12934 (N_12934,N_11773,N_11310);
nand U12935 (N_12935,N_11612,N_11965);
nand U12936 (N_12936,N_10720,N_10850);
and U12937 (N_12937,N_11822,N_11200);
xnor U12938 (N_12938,N_11155,N_11961);
or U12939 (N_12939,N_11673,N_11610);
or U12940 (N_12940,N_11472,N_11804);
and U12941 (N_12941,N_11519,N_10516);
or U12942 (N_12942,N_11166,N_11595);
nor U12943 (N_12943,N_11740,N_10951);
or U12944 (N_12944,N_11290,N_11646);
nand U12945 (N_12945,N_11643,N_11923);
nor U12946 (N_12946,N_11353,N_11938);
and U12947 (N_12947,N_10824,N_10587);
or U12948 (N_12948,N_10987,N_11900);
nor U12949 (N_12949,N_11665,N_11797);
nand U12950 (N_12950,N_11491,N_10782);
or U12951 (N_12951,N_11867,N_11918);
nor U12952 (N_12952,N_11151,N_11109);
or U12953 (N_12953,N_11034,N_10679);
or U12954 (N_12954,N_11247,N_11161);
nand U12955 (N_12955,N_11571,N_11756);
nand U12956 (N_12956,N_11613,N_10889);
xnor U12957 (N_12957,N_11063,N_11309);
and U12958 (N_12958,N_11916,N_11841);
nand U12959 (N_12959,N_10773,N_11669);
and U12960 (N_12960,N_11295,N_11029);
or U12961 (N_12961,N_11100,N_11156);
nor U12962 (N_12962,N_10790,N_11833);
or U12963 (N_12963,N_11334,N_11776);
nor U12964 (N_12964,N_11814,N_11095);
nand U12965 (N_12965,N_11445,N_11514);
and U12966 (N_12966,N_11675,N_11272);
xor U12967 (N_12967,N_10547,N_11276);
and U12968 (N_12968,N_10982,N_10685);
xor U12969 (N_12969,N_11681,N_10858);
nor U12970 (N_12970,N_10544,N_10640);
xnor U12971 (N_12971,N_11302,N_10788);
or U12972 (N_12972,N_10566,N_10527);
and U12973 (N_12973,N_10674,N_10979);
nor U12974 (N_12974,N_11553,N_11643);
nor U12975 (N_12975,N_11099,N_11881);
xor U12976 (N_12976,N_11179,N_11071);
nand U12977 (N_12977,N_11729,N_11080);
nor U12978 (N_12978,N_10944,N_11131);
nand U12979 (N_12979,N_11659,N_11506);
and U12980 (N_12980,N_11099,N_11375);
nand U12981 (N_12981,N_11677,N_11558);
xor U12982 (N_12982,N_11197,N_10941);
or U12983 (N_12983,N_11742,N_11776);
and U12984 (N_12984,N_11548,N_11807);
or U12985 (N_12985,N_10549,N_11712);
or U12986 (N_12986,N_10909,N_10649);
xnor U12987 (N_12987,N_11255,N_10665);
nand U12988 (N_12988,N_11470,N_11234);
and U12989 (N_12989,N_10742,N_10890);
or U12990 (N_12990,N_11295,N_11012);
xnor U12991 (N_12991,N_11465,N_11142);
or U12992 (N_12992,N_11647,N_11828);
nand U12993 (N_12993,N_10853,N_11429);
and U12994 (N_12994,N_11501,N_11832);
and U12995 (N_12995,N_11460,N_11084);
nand U12996 (N_12996,N_11618,N_11443);
xnor U12997 (N_12997,N_11264,N_10670);
nor U12998 (N_12998,N_10524,N_11862);
nor U12999 (N_12999,N_10717,N_11955);
nor U13000 (N_13000,N_11974,N_11595);
and U13001 (N_13001,N_10707,N_11753);
xor U13002 (N_13002,N_11013,N_11276);
nor U13003 (N_13003,N_11419,N_11709);
nor U13004 (N_13004,N_10885,N_11271);
nand U13005 (N_13005,N_10968,N_11311);
xor U13006 (N_13006,N_11640,N_10722);
and U13007 (N_13007,N_11932,N_11108);
nor U13008 (N_13008,N_10796,N_11988);
xor U13009 (N_13009,N_10671,N_11930);
and U13010 (N_13010,N_10608,N_11341);
nand U13011 (N_13011,N_10553,N_10867);
or U13012 (N_13012,N_11416,N_11061);
and U13013 (N_13013,N_11755,N_10797);
nand U13014 (N_13014,N_11053,N_10947);
nand U13015 (N_13015,N_11551,N_11118);
and U13016 (N_13016,N_11489,N_11375);
and U13017 (N_13017,N_11612,N_11946);
xor U13018 (N_13018,N_10663,N_11126);
and U13019 (N_13019,N_11607,N_10709);
nor U13020 (N_13020,N_11500,N_10513);
nand U13021 (N_13021,N_11933,N_11786);
or U13022 (N_13022,N_11694,N_10648);
xnor U13023 (N_13023,N_11070,N_11840);
or U13024 (N_13024,N_11537,N_11464);
and U13025 (N_13025,N_11079,N_11084);
or U13026 (N_13026,N_11214,N_11720);
nor U13027 (N_13027,N_11643,N_10971);
nand U13028 (N_13028,N_11220,N_11522);
and U13029 (N_13029,N_11504,N_10503);
or U13030 (N_13030,N_10956,N_11640);
or U13031 (N_13031,N_10563,N_11162);
xor U13032 (N_13032,N_11488,N_10894);
nor U13033 (N_13033,N_10811,N_10539);
nand U13034 (N_13034,N_11615,N_10973);
and U13035 (N_13035,N_11869,N_11875);
nor U13036 (N_13036,N_10740,N_10667);
or U13037 (N_13037,N_10946,N_11381);
nand U13038 (N_13038,N_11419,N_11828);
nand U13039 (N_13039,N_10557,N_11942);
and U13040 (N_13040,N_11033,N_10774);
and U13041 (N_13041,N_11624,N_11719);
nand U13042 (N_13042,N_10510,N_10943);
nor U13043 (N_13043,N_11075,N_10935);
nor U13044 (N_13044,N_11468,N_11907);
nor U13045 (N_13045,N_11745,N_11000);
and U13046 (N_13046,N_11525,N_10521);
xnor U13047 (N_13047,N_11096,N_11971);
and U13048 (N_13048,N_10982,N_11797);
xnor U13049 (N_13049,N_10892,N_11738);
xor U13050 (N_13050,N_11847,N_10940);
and U13051 (N_13051,N_11056,N_11723);
nand U13052 (N_13052,N_11682,N_11809);
and U13053 (N_13053,N_11538,N_11764);
and U13054 (N_13054,N_11489,N_10788);
nor U13055 (N_13055,N_10604,N_10778);
nor U13056 (N_13056,N_11829,N_10586);
nand U13057 (N_13057,N_11646,N_11893);
xnor U13058 (N_13058,N_10786,N_10591);
nor U13059 (N_13059,N_11801,N_11398);
nor U13060 (N_13060,N_11129,N_11043);
nand U13061 (N_13061,N_11017,N_11936);
nor U13062 (N_13062,N_10583,N_10852);
and U13063 (N_13063,N_11866,N_10647);
nor U13064 (N_13064,N_11081,N_11964);
nand U13065 (N_13065,N_10600,N_11330);
or U13066 (N_13066,N_10767,N_10717);
and U13067 (N_13067,N_11185,N_11739);
or U13068 (N_13068,N_10750,N_11770);
xnor U13069 (N_13069,N_11662,N_11062);
nor U13070 (N_13070,N_11564,N_11729);
nor U13071 (N_13071,N_11095,N_11107);
nor U13072 (N_13072,N_11712,N_11398);
nor U13073 (N_13073,N_10689,N_11943);
or U13074 (N_13074,N_10553,N_11468);
nand U13075 (N_13075,N_11728,N_11077);
or U13076 (N_13076,N_10864,N_11029);
nand U13077 (N_13077,N_10821,N_11715);
xnor U13078 (N_13078,N_11507,N_11462);
nor U13079 (N_13079,N_10792,N_10653);
nand U13080 (N_13080,N_10901,N_11391);
or U13081 (N_13081,N_11783,N_11597);
or U13082 (N_13082,N_11953,N_11005);
and U13083 (N_13083,N_11386,N_11054);
nor U13084 (N_13084,N_10563,N_10973);
nor U13085 (N_13085,N_11711,N_11979);
or U13086 (N_13086,N_11653,N_11710);
xor U13087 (N_13087,N_11834,N_10899);
nand U13088 (N_13088,N_11966,N_10706);
nor U13089 (N_13089,N_11890,N_11141);
or U13090 (N_13090,N_11287,N_11962);
or U13091 (N_13091,N_10841,N_10980);
and U13092 (N_13092,N_10680,N_11967);
or U13093 (N_13093,N_10661,N_11468);
xor U13094 (N_13094,N_11786,N_11171);
nor U13095 (N_13095,N_10768,N_10678);
and U13096 (N_13096,N_11991,N_11878);
nand U13097 (N_13097,N_11891,N_11862);
and U13098 (N_13098,N_10971,N_11969);
and U13099 (N_13099,N_11941,N_10765);
nor U13100 (N_13100,N_11732,N_11448);
xnor U13101 (N_13101,N_11009,N_11803);
nor U13102 (N_13102,N_11444,N_11223);
nand U13103 (N_13103,N_11014,N_10952);
nand U13104 (N_13104,N_11174,N_11583);
xnor U13105 (N_13105,N_11958,N_10774);
xnor U13106 (N_13106,N_11582,N_10528);
xor U13107 (N_13107,N_10778,N_11364);
or U13108 (N_13108,N_10974,N_11669);
and U13109 (N_13109,N_11679,N_11597);
xnor U13110 (N_13110,N_10723,N_11338);
nand U13111 (N_13111,N_11771,N_11880);
nor U13112 (N_13112,N_11219,N_11949);
or U13113 (N_13113,N_11222,N_10608);
nand U13114 (N_13114,N_11140,N_11878);
nor U13115 (N_13115,N_10689,N_11966);
or U13116 (N_13116,N_10854,N_11829);
or U13117 (N_13117,N_11882,N_11981);
and U13118 (N_13118,N_10573,N_10899);
nor U13119 (N_13119,N_11805,N_11729);
xnor U13120 (N_13120,N_10622,N_11369);
nor U13121 (N_13121,N_11399,N_11789);
nor U13122 (N_13122,N_10840,N_11160);
or U13123 (N_13123,N_10702,N_10603);
nor U13124 (N_13124,N_10699,N_11079);
or U13125 (N_13125,N_10818,N_11514);
nand U13126 (N_13126,N_11774,N_11402);
nand U13127 (N_13127,N_11671,N_11655);
nand U13128 (N_13128,N_11997,N_11543);
xor U13129 (N_13129,N_11255,N_10850);
nand U13130 (N_13130,N_11937,N_11134);
and U13131 (N_13131,N_10519,N_10722);
nand U13132 (N_13132,N_10889,N_11819);
nand U13133 (N_13133,N_11634,N_11334);
xnor U13134 (N_13134,N_11462,N_11756);
xnor U13135 (N_13135,N_11870,N_11866);
nor U13136 (N_13136,N_11637,N_10600);
xor U13137 (N_13137,N_11729,N_11288);
nand U13138 (N_13138,N_10915,N_11208);
nor U13139 (N_13139,N_11764,N_11855);
nand U13140 (N_13140,N_11262,N_11715);
xor U13141 (N_13141,N_11225,N_10905);
xor U13142 (N_13142,N_10861,N_11712);
or U13143 (N_13143,N_11058,N_11228);
or U13144 (N_13144,N_10651,N_11732);
xnor U13145 (N_13145,N_11266,N_11453);
nor U13146 (N_13146,N_11960,N_11623);
nand U13147 (N_13147,N_10948,N_11177);
xnor U13148 (N_13148,N_11635,N_11302);
xor U13149 (N_13149,N_11575,N_11213);
nor U13150 (N_13150,N_11853,N_10553);
and U13151 (N_13151,N_10945,N_10781);
or U13152 (N_13152,N_10667,N_11833);
xnor U13153 (N_13153,N_10972,N_11310);
or U13154 (N_13154,N_10758,N_11181);
nor U13155 (N_13155,N_11314,N_11877);
and U13156 (N_13156,N_10922,N_11732);
xnor U13157 (N_13157,N_10946,N_10860);
nand U13158 (N_13158,N_11645,N_11007);
nand U13159 (N_13159,N_10508,N_10740);
or U13160 (N_13160,N_11902,N_11667);
nor U13161 (N_13161,N_11721,N_10714);
nand U13162 (N_13162,N_11269,N_11670);
xnor U13163 (N_13163,N_10560,N_11564);
and U13164 (N_13164,N_11820,N_10632);
xor U13165 (N_13165,N_11874,N_10799);
and U13166 (N_13166,N_11529,N_11789);
xnor U13167 (N_13167,N_11156,N_11072);
nor U13168 (N_13168,N_11015,N_11889);
and U13169 (N_13169,N_10534,N_11181);
and U13170 (N_13170,N_11598,N_11202);
and U13171 (N_13171,N_11022,N_11343);
and U13172 (N_13172,N_11272,N_11318);
and U13173 (N_13173,N_11494,N_10800);
xor U13174 (N_13174,N_11485,N_10715);
and U13175 (N_13175,N_10980,N_11280);
nor U13176 (N_13176,N_11392,N_11212);
xor U13177 (N_13177,N_11072,N_10817);
xnor U13178 (N_13178,N_10936,N_11092);
nand U13179 (N_13179,N_10897,N_11498);
xor U13180 (N_13180,N_11028,N_11095);
nor U13181 (N_13181,N_11478,N_10917);
nand U13182 (N_13182,N_11704,N_10752);
or U13183 (N_13183,N_11274,N_10627);
nor U13184 (N_13184,N_11664,N_11564);
nor U13185 (N_13185,N_11023,N_11364);
and U13186 (N_13186,N_10807,N_10806);
nor U13187 (N_13187,N_10771,N_10920);
and U13188 (N_13188,N_11118,N_10813);
and U13189 (N_13189,N_10719,N_10669);
nor U13190 (N_13190,N_11277,N_10682);
nand U13191 (N_13191,N_11293,N_11648);
nor U13192 (N_13192,N_11518,N_10929);
and U13193 (N_13193,N_10609,N_11289);
nand U13194 (N_13194,N_11149,N_11557);
and U13195 (N_13195,N_10623,N_11249);
nor U13196 (N_13196,N_10673,N_11085);
nand U13197 (N_13197,N_10593,N_10858);
nor U13198 (N_13198,N_11607,N_11928);
nor U13199 (N_13199,N_11406,N_10644);
or U13200 (N_13200,N_11751,N_10842);
nand U13201 (N_13201,N_11462,N_11682);
nor U13202 (N_13202,N_11833,N_11665);
nor U13203 (N_13203,N_10851,N_11913);
nor U13204 (N_13204,N_11853,N_11489);
nand U13205 (N_13205,N_11059,N_11083);
nand U13206 (N_13206,N_11542,N_11000);
and U13207 (N_13207,N_10521,N_11553);
nor U13208 (N_13208,N_11421,N_10989);
nor U13209 (N_13209,N_10610,N_10665);
or U13210 (N_13210,N_11867,N_11409);
or U13211 (N_13211,N_10995,N_11259);
xor U13212 (N_13212,N_11995,N_10597);
xor U13213 (N_13213,N_11734,N_11917);
xnor U13214 (N_13214,N_10674,N_11927);
nor U13215 (N_13215,N_11111,N_11655);
and U13216 (N_13216,N_11323,N_11028);
xor U13217 (N_13217,N_11667,N_11479);
or U13218 (N_13218,N_10504,N_10793);
and U13219 (N_13219,N_11987,N_10992);
xor U13220 (N_13220,N_10570,N_11184);
nor U13221 (N_13221,N_10741,N_11128);
or U13222 (N_13222,N_10637,N_11202);
nor U13223 (N_13223,N_11298,N_10996);
or U13224 (N_13224,N_11838,N_10560);
nand U13225 (N_13225,N_10596,N_10712);
and U13226 (N_13226,N_11800,N_11691);
xor U13227 (N_13227,N_10997,N_10522);
or U13228 (N_13228,N_11267,N_11333);
nor U13229 (N_13229,N_11296,N_11029);
and U13230 (N_13230,N_11321,N_10907);
and U13231 (N_13231,N_11671,N_11658);
or U13232 (N_13232,N_11485,N_11146);
nor U13233 (N_13233,N_10933,N_11942);
and U13234 (N_13234,N_10763,N_11587);
and U13235 (N_13235,N_11902,N_10565);
and U13236 (N_13236,N_11874,N_10837);
nor U13237 (N_13237,N_11686,N_11153);
or U13238 (N_13238,N_10917,N_10715);
nor U13239 (N_13239,N_11621,N_10964);
nor U13240 (N_13240,N_10921,N_10883);
or U13241 (N_13241,N_10627,N_11521);
and U13242 (N_13242,N_10705,N_11879);
xnor U13243 (N_13243,N_11199,N_11355);
or U13244 (N_13244,N_10649,N_10840);
or U13245 (N_13245,N_11130,N_10713);
or U13246 (N_13246,N_11901,N_11885);
nor U13247 (N_13247,N_10502,N_11057);
nor U13248 (N_13248,N_11787,N_11847);
and U13249 (N_13249,N_10805,N_10947);
nand U13250 (N_13250,N_11949,N_10911);
nand U13251 (N_13251,N_11764,N_11895);
or U13252 (N_13252,N_10696,N_11828);
nor U13253 (N_13253,N_11348,N_11709);
nor U13254 (N_13254,N_10772,N_10868);
nor U13255 (N_13255,N_11586,N_11244);
or U13256 (N_13256,N_10576,N_11372);
or U13257 (N_13257,N_11266,N_10847);
and U13258 (N_13258,N_10801,N_10895);
nor U13259 (N_13259,N_10841,N_10772);
or U13260 (N_13260,N_11165,N_11927);
and U13261 (N_13261,N_11932,N_11203);
nor U13262 (N_13262,N_11533,N_11371);
nor U13263 (N_13263,N_10890,N_11446);
or U13264 (N_13264,N_10926,N_11056);
and U13265 (N_13265,N_11325,N_11752);
nor U13266 (N_13266,N_11541,N_10655);
xor U13267 (N_13267,N_11401,N_11642);
and U13268 (N_13268,N_11761,N_11902);
nand U13269 (N_13269,N_10643,N_10891);
or U13270 (N_13270,N_10621,N_10599);
xor U13271 (N_13271,N_10899,N_11713);
xor U13272 (N_13272,N_10992,N_10578);
nor U13273 (N_13273,N_10668,N_10888);
and U13274 (N_13274,N_11847,N_10742);
and U13275 (N_13275,N_10652,N_11455);
or U13276 (N_13276,N_11416,N_11266);
xnor U13277 (N_13277,N_11025,N_11880);
and U13278 (N_13278,N_11537,N_10870);
and U13279 (N_13279,N_11333,N_11973);
and U13280 (N_13280,N_10797,N_11973);
or U13281 (N_13281,N_10784,N_11173);
and U13282 (N_13282,N_10756,N_11303);
nor U13283 (N_13283,N_10529,N_11950);
and U13284 (N_13284,N_11941,N_11132);
nand U13285 (N_13285,N_11154,N_11591);
xor U13286 (N_13286,N_11979,N_11972);
nor U13287 (N_13287,N_11910,N_10950);
xnor U13288 (N_13288,N_11343,N_10989);
and U13289 (N_13289,N_11391,N_10591);
nor U13290 (N_13290,N_10996,N_10754);
xnor U13291 (N_13291,N_10935,N_11199);
or U13292 (N_13292,N_10598,N_10914);
nor U13293 (N_13293,N_11615,N_10722);
nor U13294 (N_13294,N_11400,N_11965);
xor U13295 (N_13295,N_10918,N_10554);
or U13296 (N_13296,N_11630,N_11668);
or U13297 (N_13297,N_11608,N_10750);
nand U13298 (N_13298,N_11163,N_10960);
or U13299 (N_13299,N_10578,N_10887);
nor U13300 (N_13300,N_11730,N_11101);
or U13301 (N_13301,N_11603,N_10924);
or U13302 (N_13302,N_11213,N_11792);
nor U13303 (N_13303,N_10665,N_11567);
or U13304 (N_13304,N_11782,N_11377);
nor U13305 (N_13305,N_11563,N_11858);
and U13306 (N_13306,N_10698,N_10776);
xor U13307 (N_13307,N_11445,N_10940);
nor U13308 (N_13308,N_11354,N_11833);
or U13309 (N_13309,N_10945,N_11567);
nor U13310 (N_13310,N_11482,N_10854);
nand U13311 (N_13311,N_11729,N_11270);
nand U13312 (N_13312,N_11754,N_11401);
or U13313 (N_13313,N_11676,N_11463);
or U13314 (N_13314,N_11581,N_11864);
nand U13315 (N_13315,N_11006,N_11381);
nor U13316 (N_13316,N_10798,N_11215);
nand U13317 (N_13317,N_11663,N_11145);
nand U13318 (N_13318,N_11286,N_11414);
and U13319 (N_13319,N_11275,N_11032);
or U13320 (N_13320,N_11172,N_11652);
xnor U13321 (N_13321,N_11745,N_10825);
xor U13322 (N_13322,N_11190,N_11120);
nor U13323 (N_13323,N_10604,N_10795);
xnor U13324 (N_13324,N_10578,N_11453);
and U13325 (N_13325,N_10675,N_11261);
or U13326 (N_13326,N_10831,N_11925);
xor U13327 (N_13327,N_10997,N_11847);
xnor U13328 (N_13328,N_11331,N_11334);
and U13329 (N_13329,N_11990,N_10710);
nor U13330 (N_13330,N_10804,N_11164);
nor U13331 (N_13331,N_11832,N_11029);
nand U13332 (N_13332,N_10537,N_11721);
and U13333 (N_13333,N_11244,N_10815);
xor U13334 (N_13334,N_11371,N_11401);
xnor U13335 (N_13335,N_10990,N_11780);
nand U13336 (N_13336,N_11796,N_11220);
xnor U13337 (N_13337,N_11028,N_11308);
and U13338 (N_13338,N_11878,N_11349);
and U13339 (N_13339,N_11423,N_11752);
or U13340 (N_13340,N_11541,N_11100);
nor U13341 (N_13341,N_11467,N_11221);
nand U13342 (N_13342,N_10685,N_11037);
xor U13343 (N_13343,N_11911,N_10713);
nand U13344 (N_13344,N_11751,N_11804);
and U13345 (N_13345,N_11613,N_11499);
nand U13346 (N_13346,N_11053,N_11752);
nand U13347 (N_13347,N_11332,N_10944);
and U13348 (N_13348,N_10864,N_10904);
and U13349 (N_13349,N_10781,N_11686);
or U13350 (N_13350,N_10792,N_11562);
or U13351 (N_13351,N_11843,N_10835);
nand U13352 (N_13352,N_11214,N_11513);
nor U13353 (N_13353,N_11370,N_10960);
nor U13354 (N_13354,N_11368,N_10688);
nand U13355 (N_13355,N_10743,N_10719);
and U13356 (N_13356,N_10862,N_10780);
nand U13357 (N_13357,N_11384,N_11402);
nand U13358 (N_13358,N_11047,N_10679);
and U13359 (N_13359,N_10638,N_11367);
nand U13360 (N_13360,N_10984,N_11657);
and U13361 (N_13361,N_11573,N_10885);
nor U13362 (N_13362,N_10945,N_11933);
nand U13363 (N_13363,N_11048,N_11577);
nor U13364 (N_13364,N_11887,N_10612);
nor U13365 (N_13365,N_11477,N_11305);
nor U13366 (N_13366,N_11185,N_11195);
xor U13367 (N_13367,N_11834,N_10983);
nand U13368 (N_13368,N_11506,N_10931);
or U13369 (N_13369,N_11535,N_11613);
and U13370 (N_13370,N_11707,N_11999);
or U13371 (N_13371,N_10645,N_10737);
nand U13372 (N_13372,N_11312,N_11770);
or U13373 (N_13373,N_10829,N_10935);
nand U13374 (N_13374,N_11403,N_10956);
xnor U13375 (N_13375,N_11953,N_11908);
nand U13376 (N_13376,N_10553,N_11987);
and U13377 (N_13377,N_10946,N_11504);
nand U13378 (N_13378,N_10757,N_11131);
or U13379 (N_13379,N_10525,N_10651);
and U13380 (N_13380,N_11788,N_11589);
xnor U13381 (N_13381,N_11436,N_11043);
xor U13382 (N_13382,N_11762,N_10674);
xnor U13383 (N_13383,N_10795,N_11391);
nand U13384 (N_13384,N_11869,N_10520);
and U13385 (N_13385,N_10902,N_11823);
and U13386 (N_13386,N_11861,N_11750);
xor U13387 (N_13387,N_10845,N_11424);
nor U13388 (N_13388,N_10809,N_11756);
nand U13389 (N_13389,N_10799,N_11601);
xor U13390 (N_13390,N_10740,N_10761);
or U13391 (N_13391,N_10896,N_10549);
xnor U13392 (N_13392,N_11242,N_10879);
or U13393 (N_13393,N_11705,N_10660);
or U13394 (N_13394,N_10716,N_11199);
and U13395 (N_13395,N_11823,N_10818);
or U13396 (N_13396,N_10670,N_11782);
xnor U13397 (N_13397,N_11715,N_10820);
nand U13398 (N_13398,N_10983,N_11779);
and U13399 (N_13399,N_11189,N_10700);
and U13400 (N_13400,N_11074,N_11847);
nor U13401 (N_13401,N_11978,N_10714);
and U13402 (N_13402,N_11712,N_11219);
xor U13403 (N_13403,N_11333,N_11086);
nor U13404 (N_13404,N_10909,N_10919);
nor U13405 (N_13405,N_11236,N_11269);
or U13406 (N_13406,N_11621,N_11673);
or U13407 (N_13407,N_11753,N_11372);
or U13408 (N_13408,N_11445,N_10744);
xor U13409 (N_13409,N_11093,N_11225);
or U13410 (N_13410,N_10591,N_11113);
nand U13411 (N_13411,N_11758,N_10667);
or U13412 (N_13412,N_11647,N_11220);
nor U13413 (N_13413,N_11276,N_11987);
or U13414 (N_13414,N_11516,N_11985);
nand U13415 (N_13415,N_11431,N_11551);
nor U13416 (N_13416,N_10706,N_11056);
nor U13417 (N_13417,N_10604,N_11576);
nand U13418 (N_13418,N_10845,N_11092);
nand U13419 (N_13419,N_11924,N_11040);
nor U13420 (N_13420,N_11507,N_11776);
and U13421 (N_13421,N_11287,N_10898);
and U13422 (N_13422,N_10724,N_11451);
nand U13423 (N_13423,N_10657,N_11582);
nand U13424 (N_13424,N_11492,N_10820);
nand U13425 (N_13425,N_11286,N_10850);
nand U13426 (N_13426,N_11215,N_11688);
xnor U13427 (N_13427,N_10580,N_11760);
xor U13428 (N_13428,N_11527,N_10579);
xnor U13429 (N_13429,N_11469,N_10721);
nor U13430 (N_13430,N_11505,N_11491);
or U13431 (N_13431,N_10557,N_11628);
and U13432 (N_13432,N_10548,N_10538);
nor U13433 (N_13433,N_10725,N_11829);
nand U13434 (N_13434,N_11900,N_11385);
xor U13435 (N_13435,N_11212,N_10814);
nor U13436 (N_13436,N_11298,N_11981);
nand U13437 (N_13437,N_11903,N_10626);
or U13438 (N_13438,N_11811,N_11494);
xor U13439 (N_13439,N_11721,N_11220);
nor U13440 (N_13440,N_10884,N_11753);
xor U13441 (N_13441,N_11662,N_10596);
nand U13442 (N_13442,N_11192,N_11944);
xnor U13443 (N_13443,N_11697,N_11149);
xor U13444 (N_13444,N_11694,N_11044);
nor U13445 (N_13445,N_10543,N_11404);
nor U13446 (N_13446,N_11900,N_11940);
xnor U13447 (N_13447,N_11672,N_11815);
xnor U13448 (N_13448,N_11873,N_10922);
and U13449 (N_13449,N_11290,N_11062);
and U13450 (N_13450,N_11298,N_11456);
nor U13451 (N_13451,N_10502,N_11459);
nand U13452 (N_13452,N_11678,N_11964);
nor U13453 (N_13453,N_11062,N_11483);
nor U13454 (N_13454,N_11523,N_11342);
nor U13455 (N_13455,N_10819,N_11722);
and U13456 (N_13456,N_11457,N_11082);
or U13457 (N_13457,N_11579,N_11568);
or U13458 (N_13458,N_11569,N_10680);
xnor U13459 (N_13459,N_10950,N_11058);
nor U13460 (N_13460,N_11732,N_11539);
nand U13461 (N_13461,N_11912,N_11745);
or U13462 (N_13462,N_10915,N_10609);
xor U13463 (N_13463,N_11748,N_11520);
or U13464 (N_13464,N_11106,N_11899);
and U13465 (N_13465,N_11866,N_11020);
nor U13466 (N_13466,N_11560,N_11160);
or U13467 (N_13467,N_11275,N_11492);
nand U13468 (N_13468,N_11484,N_10965);
xnor U13469 (N_13469,N_11842,N_11579);
nor U13470 (N_13470,N_10936,N_10856);
or U13471 (N_13471,N_11471,N_11959);
xnor U13472 (N_13472,N_11913,N_11960);
or U13473 (N_13473,N_11017,N_11305);
and U13474 (N_13474,N_11301,N_11670);
or U13475 (N_13475,N_11630,N_11653);
nand U13476 (N_13476,N_11793,N_10964);
xor U13477 (N_13477,N_10657,N_11962);
or U13478 (N_13478,N_10514,N_11047);
nor U13479 (N_13479,N_11434,N_10594);
and U13480 (N_13480,N_11022,N_10746);
xor U13481 (N_13481,N_11408,N_11122);
nor U13482 (N_13482,N_11570,N_11523);
or U13483 (N_13483,N_11262,N_11798);
or U13484 (N_13484,N_11271,N_11358);
xnor U13485 (N_13485,N_11539,N_11825);
xor U13486 (N_13486,N_11569,N_11772);
nor U13487 (N_13487,N_11741,N_11000);
nor U13488 (N_13488,N_10550,N_11317);
or U13489 (N_13489,N_11614,N_11522);
nor U13490 (N_13490,N_11055,N_10571);
xor U13491 (N_13491,N_11864,N_11038);
xnor U13492 (N_13492,N_11237,N_10520);
xnor U13493 (N_13493,N_11179,N_10783);
or U13494 (N_13494,N_11169,N_11410);
nand U13495 (N_13495,N_11572,N_11703);
xor U13496 (N_13496,N_11524,N_11375);
nor U13497 (N_13497,N_11804,N_11758);
or U13498 (N_13498,N_11939,N_10870);
xnor U13499 (N_13499,N_11362,N_11148);
nor U13500 (N_13500,N_12396,N_12416);
and U13501 (N_13501,N_12253,N_12483);
xor U13502 (N_13502,N_13105,N_12673);
nor U13503 (N_13503,N_13146,N_12127);
or U13504 (N_13504,N_12714,N_12315);
nand U13505 (N_13505,N_12776,N_12816);
and U13506 (N_13506,N_13142,N_12247);
and U13507 (N_13507,N_13394,N_12112);
nor U13508 (N_13508,N_12033,N_13433);
xnor U13509 (N_13509,N_12849,N_12382);
xor U13510 (N_13510,N_12448,N_12554);
xor U13511 (N_13511,N_12392,N_12370);
nand U13512 (N_13512,N_12348,N_13084);
and U13513 (N_13513,N_12410,N_12181);
or U13514 (N_13514,N_13415,N_13033);
xnor U13515 (N_13515,N_13274,N_13235);
and U13516 (N_13516,N_12552,N_12055);
nor U13517 (N_13517,N_13068,N_12868);
xor U13518 (N_13518,N_12739,N_13216);
nand U13519 (N_13519,N_12399,N_12526);
and U13520 (N_13520,N_12901,N_13438);
and U13521 (N_13521,N_12944,N_13054);
nand U13522 (N_13522,N_12060,N_13237);
and U13523 (N_13523,N_12621,N_13183);
nand U13524 (N_13524,N_13390,N_12708);
nor U13525 (N_13525,N_12069,N_12845);
or U13526 (N_13526,N_13449,N_12299);
nand U13527 (N_13527,N_12777,N_12211);
xnor U13528 (N_13528,N_12210,N_12185);
or U13529 (N_13529,N_13171,N_12962);
or U13530 (N_13530,N_12974,N_12682);
xnor U13531 (N_13531,N_12472,N_12403);
and U13532 (N_13532,N_12276,N_13089);
nor U13533 (N_13533,N_12627,N_12930);
xnor U13534 (N_13534,N_12763,N_13116);
nand U13535 (N_13535,N_12109,N_12238);
nand U13536 (N_13536,N_12351,N_12030);
and U13537 (N_13537,N_12164,N_12497);
xor U13538 (N_13538,N_12218,N_12435);
xor U13539 (N_13539,N_12307,N_12766);
xor U13540 (N_13540,N_12861,N_13258);
nor U13541 (N_13541,N_12327,N_12848);
nand U13542 (N_13542,N_13189,N_12574);
xor U13543 (N_13543,N_13331,N_13031);
xnor U13544 (N_13544,N_12313,N_12473);
and U13545 (N_13545,N_12778,N_13200);
nor U13546 (N_13546,N_13012,N_12465);
or U13547 (N_13547,N_12791,N_12545);
nor U13548 (N_13548,N_12258,N_12373);
nand U13549 (N_13549,N_13174,N_12636);
or U13550 (N_13550,N_13225,N_13292);
nor U13551 (N_13551,N_12368,N_13080);
xor U13552 (N_13552,N_12369,N_12136);
nand U13553 (N_13553,N_12927,N_12444);
and U13554 (N_13554,N_12407,N_12801);
and U13555 (N_13555,N_12101,N_13231);
xor U13556 (N_13556,N_12830,N_13276);
nor U13557 (N_13557,N_13322,N_13404);
or U13558 (N_13558,N_12987,N_13414);
and U13559 (N_13559,N_13297,N_12853);
nand U13560 (N_13560,N_13056,N_13419);
and U13561 (N_13561,N_12051,N_13338);
nand U13562 (N_13562,N_12786,N_12843);
xnor U13563 (N_13563,N_12793,N_12455);
nand U13564 (N_13564,N_13355,N_12479);
nand U13565 (N_13565,N_12590,N_13232);
and U13566 (N_13566,N_13079,N_12144);
or U13567 (N_13567,N_13468,N_12108);
nor U13568 (N_13568,N_12720,N_12192);
nand U13569 (N_13569,N_12635,N_13147);
nor U13570 (N_13570,N_12934,N_12639);
nor U13571 (N_13571,N_13017,N_12198);
nor U13572 (N_13572,N_12730,N_12963);
nand U13573 (N_13573,N_12893,N_13153);
nand U13574 (N_13574,N_13076,N_12279);
nor U13575 (N_13575,N_12610,N_12584);
and U13576 (N_13576,N_12311,N_13161);
nand U13577 (N_13577,N_12452,N_12489);
or U13578 (N_13578,N_12814,N_12922);
nor U13579 (N_13579,N_13362,N_13024);
xor U13580 (N_13580,N_12980,N_12289);
or U13581 (N_13581,N_13233,N_13382);
nor U13582 (N_13582,N_12072,N_12291);
and U13583 (N_13583,N_12550,N_12029);
and U13584 (N_13584,N_12260,N_12268);
or U13585 (N_13585,N_12269,N_13179);
xor U13586 (N_13586,N_12297,N_13278);
or U13587 (N_13587,N_13374,N_12756);
or U13588 (N_13588,N_13169,N_12388);
xnor U13589 (N_13589,N_12773,N_12468);
and U13590 (N_13590,N_12383,N_12310);
nand U13591 (N_13591,N_12850,N_12954);
xnor U13592 (N_13592,N_12424,N_13097);
nor U13593 (N_13593,N_13234,N_12910);
nor U13594 (N_13594,N_12747,N_13317);
nor U13595 (N_13595,N_13475,N_12607);
nor U13596 (N_13596,N_12240,N_12804);
nand U13597 (N_13597,N_13125,N_12488);
nand U13598 (N_13598,N_12623,N_13485);
nor U13599 (N_13599,N_12300,N_12949);
or U13600 (N_13600,N_12705,N_12825);
and U13601 (N_13601,N_13295,N_12264);
or U13602 (N_13602,N_13436,N_13144);
xnor U13603 (N_13603,N_12414,N_12047);
xor U13604 (N_13604,N_12429,N_13482);
or U13605 (N_13605,N_13474,N_13110);
nand U13606 (N_13606,N_12738,N_12490);
nor U13607 (N_13607,N_12042,N_13040);
nand U13608 (N_13608,N_13069,N_13151);
or U13609 (N_13609,N_12575,N_13220);
nor U13610 (N_13610,N_12255,N_12604);
and U13611 (N_13611,N_13026,N_12691);
and U13612 (N_13612,N_12937,N_12785);
and U13613 (N_13613,N_13440,N_12257);
nand U13614 (N_13614,N_12733,N_12151);
and U13615 (N_13615,N_12376,N_12725);
nand U13616 (N_13616,N_13127,N_12066);
and U13617 (N_13617,N_12206,N_12446);
xor U13618 (N_13618,N_12209,N_13120);
xnor U13619 (N_13619,N_12881,N_13444);
and U13620 (N_13620,N_12728,N_13280);
xor U13621 (N_13621,N_12835,N_13326);
and U13622 (N_13622,N_13473,N_12262);
xnor U13623 (N_13623,N_13000,N_12261);
nor U13624 (N_13624,N_12915,N_12891);
and U13625 (N_13625,N_12753,N_13316);
or U13626 (N_13626,N_12317,N_12229);
nor U13627 (N_13627,N_12035,N_13310);
nor U13628 (N_13628,N_12221,N_13128);
and U13629 (N_13629,N_12692,N_13308);
xnor U13630 (N_13630,N_13238,N_12961);
nor U13631 (N_13631,N_13427,N_12250);
nor U13632 (N_13632,N_12338,N_12665);
nor U13633 (N_13633,N_13006,N_12063);
xnor U13634 (N_13634,N_12886,N_13187);
nor U13635 (N_13635,N_12009,N_13300);
nor U13636 (N_13636,N_12088,N_13284);
nor U13637 (N_13637,N_13249,N_12393);
nor U13638 (N_13638,N_13018,N_12999);
or U13639 (N_13639,N_13401,N_13157);
xnor U13640 (N_13640,N_12654,N_12609);
or U13641 (N_13641,N_12456,N_12983);
and U13642 (N_13642,N_12558,N_12427);
and U13643 (N_13643,N_13202,N_13311);
and U13644 (N_13644,N_12844,N_13286);
or U13645 (N_13645,N_12031,N_13405);
nor U13646 (N_13646,N_13424,N_12406);
xnor U13647 (N_13647,N_12367,N_13288);
xor U13648 (N_13648,N_13357,N_12592);
nor U13649 (N_13649,N_13451,N_12286);
nor U13650 (N_13650,N_12715,N_12381);
and U13651 (N_13651,N_12235,N_12595);
or U13652 (N_13652,N_12606,N_13333);
nand U13653 (N_13653,N_12411,N_13453);
nand U13654 (N_13654,N_12233,N_12345);
and U13655 (N_13655,N_12401,N_13484);
nor U13656 (N_13656,N_12453,N_13004);
and U13657 (N_13657,N_12277,N_12026);
nor U13658 (N_13658,N_12308,N_13376);
or U13659 (N_13659,N_13201,N_12205);
nor U13660 (N_13660,N_12293,N_12531);
or U13661 (N_13661,N_12764,N_12973);
and U13662 (N_13662,N_12875,N_13291);
or U13663 (N_13663,N_13098,N_12573);
nor U13664 (N_13664,N_12833,N_12813);
or U13665 (N_13665,N_12677,N_12660);
nor U13666 (N_13666,N_13339,N_12160);
or U13667 (N_13667,N_13063,N_12391);
xnor U13668 (N_13668,N_12278,N_13042);
xor U13669 (N_13669,N_12306,N_13090);
nand U13670 (N_13670,N_13259,N_13458);
nor U13671 (N_13671,N_13119,N_13193);
xnor U13672 (N_13672,N_12827,N_13389);
nor U13673 (N_13673,N_12467,N_12896);
and U13674 (N_13674,N_13494,N_12956);
or U13675 (N_13675,N_12865,N_13448);
xor U13676 (N_13676,N_12423,N_12321);
or U13677 (N_13677,N_13269,N_12135);
nor U13678 (N_13678,N_13315,N_12740);
nor U13679 (N_13679,N_13454,N_12460);
xnor U13680 (N_13680,N_13122,N_12203);
nor U13681 (N_13681,N_13388,N_12994);
xnor U13682 (N_13682,N_13099,N_12661);
and U13683 (N_13683,N_12624,N_12049);
or U13684 (N_13684,N_12405,N_12282);
nor U13685 (N_13685,N_12281,N_12167);
nor U13686 (N_13686,N_12758,N_12626);
and U13687 (N_13687,N_12890,N_12729);
nor U13688 (N_13688,N_12642,N_12462);
nand U13689 (N_13689,N_12271,N_12569);
and U13690 (N_13690,N_13011,N_12750);
nor U13691 (N_13691,N_12143,N_12716);
and U13692 (N_13692,N_12062,N_13210);
xnor U13693 (N_13693,N_12248,N_12923);
and U13694 (N_13694,N_13456,N_13219);
and U13695 (N_13695,N_12292,N_13176);
nand U13696 (N_13696,N_12826,N_13057);
xnor U13697 (N_13697,N_12323,N_12092);
xnor U13698 (N_13698,N_12008,N_13184);
and U13699 (N_13699,N_12808,N_13420);
xor U13700 (N_13700,N_12476,N_12091);
and U13701 (N_13701,N_12908,N_12698);
or U13702 (N_13702,N_12765,N_13132);
xor U13703 (N_13703,N_12613,N_12749);
or U13704 (N_13704,N_13464,N_12084);
xnor U13705 (N_13705,N_12017,N_12073);
or U13706 (N_13706,N_12180,N_12529);
and U13707 (N_13707,N_13010,N_13375);
nand U13708 (N_13708,N_12123,N_13005);
xnor U13709 (N_13709,N_13402,N_12877);
xor U13710 (N_13710,N_12751,N_12491);
nand U13711 (N_13711,N_12475,N_13182);
or U13712 (N_13712,N_12717,N_12968);
or U13713 (N_13713,N_13460,N_12111);
xnor U13714 (N_13714,N_12537,N_12141);
or U13715 (N_13715,N_12847,N_12099);
and U13716 (N_13716,N_12770,N_12230);
nand U13717 (N_13717,N_12204,N_12806);
or U13718 (N_13718,N_12217,N_12413);
xnor U13719 (N_13719,N_12982,N_12957);
nor U13720 (N_13720,N_12839,N_13411);
or U13721 (N_13721,N_12556,N_12544);
nor U13722 (N_13722,N_12440,N_13499);
and U13723 (N_13723,N_12430,N_13324);
nand U13724 (N_13724,N_12421,N_12878);
nor U13725 (N_13725,N_13072,N_13013);
xor U13726 (N_13726,N_13203,N_12741);
xnor U13727 (N_13727,N_13467,N_12970);
and U13728 (N_13728,N_12418,N_12993);
nand U13729 (N_13729,N_12128,N_13378);
or U13730 (N_13730,N_12285,N_12582);
and U13731 (N_13731,N_13022,N_13156);
xor U13732 (N_13732,N_12676,N_12898);
or U13733 (N_13733,N_12105,N_13163);
nand U13734 (N_13734,N_12187,N_12649);
and U13735 (N_13735,N_12653,N_12477);
and U13736 (N_13736,N_12674,N_13043);
xnor U13737 (N_13737,N_13229,N_12384);
xnor U13738 (N_13738,N_12213,N_12334);
and U13739 (N_13739,N_13067,N_12340);
or U13740 (N_13740,N_12940,N_12829);
or U13741 (N_13741,N_12882,N_13205);
nand U13742 (N_13742,N_12666,N_13254);
nor U13743 (N_13743,N_13177,N_12718);
and U13744 (N_13744,N_13020,N_13188);
nor U13745 (N_13745,N_13262,N_12638);
nor U13746 (N_13746,N_12459,N_13393);
nor U13747 (N_13747,N_13275,N_13164);
xor U13748 (N_13748,N_13277,N_12798);
and U13749 (N_13749,N_12598,N_12528);
and U13750 (N_13750,N_12670,N_12214);
xor U13751 (N_13751,N_12939,N_12001);
xnor U13752 (N_13752,N_13091,N_13062);
nand U13753 (N_13753,N_13296,N_13348);
or U13754 (N_13754,N_12050,N_12918);
xnor U13755 (N_13755,N_12006,N_13065);
and U13756 (N_13756,N_12270,N_12436);
nand U13757 (N_13757,N_12612,N_12960);
xor U13758 (N_13758,N_12183,N_13071);
and U13759 (N_13759,N_13384,N_13445);
xor U13760 (N_13760,N_13369,N_13423);
nand U13761 (N_13761,N_13126,N_12736);
nor U13762 (N_13762,N_13046,N_12619);
nand U13763 (N_13763,N_12320,N_12837);
and U13764 (N_13764,N_12536,N_12864);
nor U13765 (N_13765,N_12565,N_13094);
xnor U13766 (N_13766,N_12580,N_12888);
nor U13767 (N_13767,N_13273,N_12754);
or U13768 (N_13768,N_13434,N_13197);
and U13769 (N_13769,N_12792,N_12104);
xor U13770 (N_13770,N_13349,N_12737);
or U13771 (N_13771,N_13323,N_12095);
xor U13772 (N_13772,N_13034,N_12471);
or U13773 (N_13773,N_12011,N_12114);
nand U13774 (N_13774,N_12120,N_13299);
and U13775 (N_13775,N_12336,N_13383);
or U13776 (N_13776,N_13078,N_13016);
nand U13777 (N_13777,N_12745,N_13015);
nor U13778 (N_13778,N_12669,N_13287);
nor U13779 (N_13779,N_12083,N_13143);
or U13780 (N_13780,N_12899,N_12046);
nor U13781 (N_13781,N_13104,N_12971);
xnor U13782 (N_13782,N_12805,N_12815);
nand U13783 (N_13783,N_12681,N_13239);
or U13784 (N_13784,N_13074,N_12428);
xnor U13785 (N_13785,N_12059,N_13082);
or U13786 (N_13786,N_13400,N_12486);
nor U13787 (N_13787,N_13486,N_12876);
and U13788 (N_13788,N_12130,N_13431);
nor U13789 (N_13789,N_12995,N_12779);
nor U13790 (N_13790,N_13093,N_12759);
nor U13791 (N_13791,N_12194,N_12439);
and U13792 (N_13792,N_13328,N_12316);
nor U13793 (N_13793,N_12675,N_12178);
and U13794 (N_13794,N_12838,N_12690);
and U13795 (N_13795,N_12375,N_13439);
nor U13796 (N_13796,N_12602,N_12236);
nor U13797 (N_13797,N_13107,N_13466);
nor U13798 (N_13798,N_13002,N_13447);
nand U13799 (N_13799,N_13092,N_12216);
xor U13800 (N_13800,N_12228,N_12967);
nand U13801 (N_13801,N_13135,N_12678);
xnor U13802 (N_13802,N_12579,N_13498);
and U13803 (N_13803,N_13003,N_12858);
and U13804 (N_13804,N_12614,N_12894);
nand U13805 (N_13805,N_13246,N_12871);
nor U13806 (N_13806,N_12911,N_13133);
or U13807 (N_13807,N_13257,N_13211);
and U13808 (N_13808,N_12931,N_12324);
nor U13809 (N_13809,N_13019,N_13070);
nand U13810 (N_13810,N_12506,N_12823);
xor U13811 (N_13811,N_12726,N_12684);
nor U13812 (N_13812,N_12094,N_12567);
nand U13813 (N_13813,N_12789,N_12975);
nor U13814 (N_13814,N_12080,N_12470);
nor U13815 (N_13815,N_12984,N_12451);
or U13816 (N_13816,N_13181,N_12727);
xnor U13817 (N_13817,N_12224,N_13425);
or U13818 (N_13818,N_12431,N_13285);
nor U13819 (N_13819,N_13283,N_13463);
nand U13820 (N_13820,N_12075,N_13047);
xnor U13821 (N_13821,N_13111,N_12457);
xor U13822 (N_13822,N_12622,N_12836);
or U13823 (N_13823,N_12625,N_12869);
nor U13824 (N_13824,N_13334,N_13198);
or U13825 (N_13825,N_12152,N_13204);
nor U13826 (N_13826,N_12339,N_13061);
nand U13827 (N_13827,N_13083,N_12965);
nor U13828 (N_13828,N_13367,N_12570);
and U13829 (N_13829,N_12053,N_12781);
nor U13830 (N_13830,N_12860,N_13170);
nand U13831 (N_13831,N_12484,N_12137);
and U13832 (N_13832,N_12672,N_12329);
and U13833 (N_13833,N_12952,N_13282);
nand U13834 (N_13834,N_12562,N_12985);
nand U13835 (N_13835,N_13136,N_12232);
or U13836 (N_13836,N_12755,N_12515);
nor U13837 (N_13837,N_12731,N_12146);
and U13838 (N_13838,N_12663,N_12846);
xnor U13839 (N_13839,N_12319,N_12933);
xnor U13840 (N_13840,N_12979,N_13325);
nor U13841 (N_13841,N_12265,N_12702);
xnor U13842 (N_13842,N_12605,N_12118);
or U13843 (N_13843,N_13085,N_12748);
and U13844 (N_13844,N_12352,N_13049);
and U13845 (N_13845,N_13207,N_13408);
and U13846 (N_13846,N_12618,N_12350);
nor U13847 (N_13847,N_13281,N_12189);
or U13848 (N_13848,N_12153,N_12074);
nor U13849 (N_13849,N_13217,N_12054);
xor U13850 (N_13850,N_12664,N_13138);
xor U13851 (N_13851,N_12337,N_13346);
nor U13852 (N_13852,N_12929,N_12913);
xor U13853 (N_13853,N_12113,N_12986);
nand U13854 (N_13854,N_13462,N_12176);
nand U13855 (N_13855,N_12832,N_12723);
and U13856 (N_13856,N_12689,N_12936);
nor U13857 (N_13857,N_12364,N_13461);
nand U13858 (N_13858,N_12463,N_12070);
nor U13859 (N_13859,N_13437,N_13196);
nand U13860 (N_13860,N_12948,N_12196);
nor U13861 (N_13861,N_13483,N_12977);
or U13862 (N_13862,N_12495,N_12841);
or U13863 (N_13863,N_12964,N_13245);
nand U13864 (N_13864,N_12711,N_12207);
and U13865 (N_13865,N_12566,N_12301);
xor U13866 (N_13866,N_13155,N_12513);
nor U13867 (N_13867,N_12419,N_12555);
or U13868 (N_13868,N_13452,N_12857);
nor U13869 (N_13869,N_12599,N_13368);
or U13870 (N_13870,N_12916,N_13185);
nor U13871 (N_13871,N_13387,N_12142);
nand U13872 (N_13872,N_12818,N_12821);
nor U13873 (N_13873,N_12107,N_12110);
nor U13874 (N_13874,N_12007,N_12628);
and U13875 (N_13875,N_12199,N_12155);
nor U13876 (N_13876,N_12346,N_13457);
nor U13877 (N_13877,N_13493,N_12374);
nand U13878 (N_13878,N_12527,N_12700);
and U13879 (N_13879,N_13150,N_13397);
nor U13880 (N_13880,N_13309,N_12634);
xor U13881 (N_13881,N_12305,N_12389);
xnor U13882 (N_13882,N_12824,N_12325);
nor U13883 (N_13883,N_12201,N_12647);
nor U13884 (N_13884,N_12950,N_12769);
nor U13885 (N_13885,N_12503,N_12466);
or U13886 (N_13886,N_13496,N_13476);
and U13887 (N_13887,N_13021,N_12662);
nand U13888 (N_13888,N_13344,N_13027);
nand U13889 (N_13889,N_12856,N_13410);
or U13890 (N_13890,N_12991,N_12150);
nand U13891 (N_13891,N_12795,N_12656);
and U13892 (N_13892,N_12903,N_12713);
nand U13893 (N_13893,N_13271,N_13113);
or U13894 (N_13894,N_13430,N_12941);
and U13895 (N_13895,N_12231,N_12693);
or U13896 (N_13896,N_13130,N_13103);
nand U13897 (N_13897,N_12790,N_13053);
xnor U13898 (N_13898,N_12699,N_12811);
and U13899 (N_13899,N_12784,N_13264);
or U13900 (N_13900,N_12227,N_12521);
nand U13901 (N_13901,N_12275,N_12378);
or U13902 (N_13902,N_12617,N_12025);
and U13903 (N_13903,N_13115,N_13363);
nand U13904 (N_13904,N_13096,N_12461);
xnor U13905 (N_13905,N_12512,N_12244);
nor U13906 (N_13906,N_13168,N_13228);
or U13907 (N_13907,N_13441,N_13131);
or U13908 (N_13908,N_13180,N_12796);
nand U13909 (N_13909,N_12441,N_12658);
and U13910 (N_13910,N_12184,N_12024);
nand U13911 (N_13911,N_12583,N_13301);
and U13912 (N_13912,N_12173,N_12762);
nand U13913 (N_13913,N_13480,N_12190);
xor U13914 (N_13914,N_12443,N_12045);
nand U13915 (N_13915,N_13361,N_12831);
or U13916 (N_13916,N_12655,N_12997);
xor U13917 (N_13917,N_12398,N_13266);
nand U13918 (N_13918,N_12274,N_12298);
or U13919 (N_13919,N_12302,N_12400);
xnor U13920 (N_13920,N_12098,N_12377);
xor U13921 (N_13921,N_12012,N_12166);
or U13922 (N_13922,N_12992,N_13172);
or U13923 (N_13923,N_12147,N_12318);
nand U13924 (N_13924,N_13337,N_13370);
and U13925 (N_13925,N_12018,N_12129);
or U13926 (N_13926,N_12121,N_12354);
nand U13927 (N_13927,N_12267,N_12505);
or U13928 (N_13928,N_13114,N_12577);
nor U13929 (N_13929,N_13121,N_12097);
or U13930 (N_13930,N_13175,N_13109);
and U13931 (N_13931,N_13426,N_12182);
or U13932 (N_13932,N_12314,N_12543);
or U13933 (N_13933,N_12998,N_12897);
xnor U13934 (N_13934,N_12458,N_12568);
and U13935 (N_13935,N_12912,N_13208);
and U13936 (N_13936,N_12593,N_12819);
xnor U13937 (N_13937,N_12056,N_12280);
and U13938 (N_13938,N_13029,N_12892);
xor U13939 (N_13939,N_13218,N_12454);
or U13940 (N_13940,N_12140,N_12581);
and U13941 (N_13941,N_12016,N_12695);
or U13942 (N_13942,N_12179,N_12591);
nand U13943 (N_13943,N_12362,N_12328);
or U13944 (N_13944,N_12358,N_13224);
and U13945 (N_13945,N_13251,N_12402);
xnor U13946 (N_13946,N_13432,N_12014);
and U13947 (N_13947,N_12330,N_12879);
xor U13948 (N_13948,N_12988,N_13372);
nand U13949 (N_13949,N_13395,N_12701);
xor U13950 (N_13950,N_13058,N_12810);
xor U13951 (N_13951,N_12644,N_13243);
or U13952 (N_13952,N_13478,N_12082);
or U13953 (N_13953,N_13154,N_12522);
nand U13954 (N_13954,N_12616,N_12077);
nand U13955 (N_13955,N_12165,N_12906);
nor U13956 (N_13956,N_12041,N_12646);
nor U13957 (N_13957,N_13192,N_12175);
nand U13958 (N_13958,N_13087,N_13459);
and U13959 (N_13959,N_12290,N_12532);
xor U13960 (N_13960,N_12343,N_12990);
and U13961 (N_13961,N_12548,N_12215);
xor U13962 (N_13962,N_12498,N_12052);
nand U13963 (N_13963,N_13226,N_12048);
nor U13964 (N_13964,N_12546,N_12078);
and U13965 (N_13965,N_12951,N_12076);
nand U13966 (N_13966,N_12516,N_12571);
and U13967 (N_13967,N_12520,N_12239);
xnor U13968 (N_13968,N_12197,N_12594);
nor U13969 (N_13969,N_12820,N_12283);
and U13970 (N_13970,N_12028,N_12686);
nand U13971 (N_13971,N_12349,N_12685);
nand U13972 (N_13972,N_12071,N_12442);
nor U13973 (N_13973,N_12259,N_13081);
xor U13974 (N_13974,N_13320,N_12633);
or U13975 (N_13975,N_12415,N_12643);
nor U13976 (N_13976,N_12501,N_12530);
or U13977 (N_13977,N_13117,N_13435);
nand U13978 (N_13978,N_12417,N_13028);
nand U13979 (N_13979,N_12601,N_13159);
nand U13980 (N_13980,N_13413,N_12559);
xor U13981 (N_13981,N_12955,N_13086);
xor U13982 (N_13982,N_12862,N_12220);
and U13983 (N_13983,N_13148,N_13446);
and U13984 (N_13984,N_12359,N_12222);
or U13985 (N_13985,N_12828,N_12953);
nor U13986 (N_13986,N_12139,N_13140);
or U13987 (N_13987,N_12734,N_13442);
nor U13988 (N_13988,N_13318,N_13256);
xnor U13989 (N_13989,N_12037,N_12551);
and U13990 (N_13990,N_13222,N_13353);
xnor U13991 (N_13991,N_12921,N_12671);
and U13992 (N_13992,N_12807,N_12464);
nor U13993 (N_13993,N_13227,N_13488);
xor U13994 (N_13994,N_12600,N_12822);
and U13995 (N_13995,N_13479,N_13359);
and U13996 (N_13996,N_12068,N_12437);
nor U13997 (N_13997,N_12395,N_13298);
xor U13998 (N_13998,N_13455,N_12379);
and U13999 (N_13999,N_12086,N_12386);
xnor U14000 (N_14000,N_12926,N_12500);
xnor U14001 (N_14001,N_12043,N_12163);
nand U14002 (N_14002,N_12885,N_12966);
and U14003 (N_14003,N_12782,N_12036);
or U14004 (N_14004,N_12586,N_13036);
or U14005 (N_14005,N_12799,N_12519);
or U14006 (N_14006,N_13321,N_12093);
nor U14007 (N_14007,N_13341,N_13244);
and U14008 (N_14008,N_12226,N_12866);
nor U14009 (N_14009,N_12287,N_12003);
and U14010 (N_14010,N_12703,N_12969);
xor U14011 (N_14011,N_13343,N_12161);
xnor U14012 (N_14012,N_12688,N_12783);
nor U14013 (N_14013,N_13307,N_12668);
nand U14014 (N_14014,N_12208,N_12039);
nor U14015 (N_14015,N_12707,N_13495);
nor U14016 (N_14016,N_12597,N_12852);
nand U14017 (N_14017,N_12648,N_12637);
nor U14018 (N_14018,N_13186,N_13167);
or U14019 (N_14019,N_13134,N_13267);
nor U14020 (N_14020,N_12251,N_12564);
xor U14021 (N_14021,N_12044,N_12202);
nand U14022 (N_14022,N_12978,N_13306);
and U14023 (N_14023,N_12508,N_12761);
nand U14024 (N_14024,N_12744,N_13014);
or U14025 (N_14025,N_12245,N_12057);
xnor U14026 (N_14026,N_13421,N_12387);
nor U14027 (N_14027,N_13329,N_12064);
and U14028 (N_14028,N_13360,N_12719);
or U14029 (N_14029,N_12780,N_12394);
xnor U14030 (N_14030,N_12303,N_12022);
nor U14031 (N_14031,N_12630,N_13303);
and U14032 (N_14032,N_13236,N_13260);
or U14033 (N_14033,N_12000,N_12704);
nor U14034 (N_14034,N_12576,N_12735);
or U14035 (N_14035,N_12241,N_13380);
and U14036 (N_14036,N_13240,N_12124);
and U14037 (N_14037,N_13327,N_12225);
and U14038 (N_14038,N_12263,N_12117);
and U14039 (N_14039,N_13492,N_13491);
or U14040 (N_14040,N_12549,N_12304);
nor U14041 (N_14041,N_13409,N_12863);
or U14042 (N_14042,N_12502,N_13373);
and U14043 (N_14043,N_12895,N_13302);
xor U14044 (N_14044,N_12942,N_12335);
xnor U14045 (N_14045,N_12432,N_12840);
and U14046 (N_14046,N_13051,N_13088);
or U14047 (N_14047,N_12907,N_12694);
xnor U14048 (N_14048,N_12480,N_13305);
xor U14049 (N_14049,N_12524,N_13009);
nor U14050 (N_14050,N_12237,N_13165);
nor U14051 (N_14051,N_12585,N_12040);
xor U14052 (N_14052,N_12487,N_12132);
nor U14053 (N_14053,N_13252,N_12972);
nand U14054 (N_14054,N_12511,N_12365);
xor U14055 (N_14055,N_12611,N_12924);
and U14056 (N_14056,N_12021,N_12482);
nor U14057 (N_14057,N_12015,N_12794);
nand U14058 (N_14058,N_12768,N_12817);
and U14059 (N_14059,N_12938,N_12884);
nor U14060 (N_14060,N_12195,N_12177);
or U14061 (N_14061,N_12873,N_12115);
nand U14062 (N_14062,N_12900,N_13398);
or U14063 (N_14063,N_12507,N_13312);
or U14064 (N_14064,N_13342,N_13223);
or U14065 (N_14065,N_12445,N_12019);
xor U14066 (N_14066,N_12872,N_12020);
nor U14067 (N_14067,N_12273,N_12859);
and U14068 (N_14068,N_12469,N_12883);
and U14069 (N_14069,N_12588,N_13095);
nand U14070 (N_14070,N_13064,N_12067);
or U14071 (N_14071,N_12547,N_12657);
nor U14072 (N_14072,N_12904,N_13160);
nand U14073 (N_14073,N_13045,N_12802);
nor U14074 (N_14074,N_12385,N_13330);
xor U14075 (N_14075,N_12361,N_12408);
and U14076 (N_14076,N_13450,N_12752);
and U14077 (N_14077,N_12412,N_12032);
or U14078 (N_14078,N_12058,N_12631);
xor U14079 (N_14079,N_12169,N_12525);
or U14080 (N_14080,N_12803,N_12680);
xnor U14081 (N_14081,N_13422,N_12493);
xor U14082 (N_14082,N_13101,N_12603);
nand U14083 (N_14083,N_12170,N_12296);
nor U14084 (N_14084,N_13336,N_12065);
xnor U14085 (N_14085,N_12162,N_12148);
xor U14086 (N_14086,N_12038,N_12563);
xor U14087 (N_14087,N_12331,N_13470);
and U14088 (N_14088,N_13152,N_13412);
or U14089 (N_14089,N_13190,N_13158);
or U14090 (N_14090,N_13313,N_12834);
or U14091 (N_14091,N_13212,N_12560);
or U14092 (N_14092,N_13497,N_12145);
xor U14093 (N_14093,N_13407,N_13129);
xnor U14094 (N_14094,N_12809,N_13112);
xor U14095 (N_14095,N_12332,N_12775);
or U14096 (N_14096,N_13418,N_12131);
and U14097 (N_14097,N_13429,N_13396);
xnor U14098 (N_14098,N_12420,N_12333);
xor U14099 (N_14099,N_12535,N_12958);
nor U14100 (N_14100,N_12326,N_12854);
nor U14101 (N_14101,N_12356,N_12919);
or U14102 (N_14102,N_12589,N_12851);
and U14103 (N_14103,N_13052,N_12126);
xor U14104 (N_14104,N_12288,N_13489);
or U14105 (N_14105,N_13041,N_12422);
nand U14106 (N_14106,N_12932,N_12855);
nor U14107 (N_14107,N_13199,N_13354);
nor U14108 (N_14108,N_12742,N_12004);
and U14109 (N_14109,N_12640,N_13351);
nand U14110 (N_14110,N_12002,N_13141);
nand U14111 (N_14111,N_13221,N_13030);
nor U14112 (N_14112,N_12171,N_12492);
or U14113 (N_14113,N_12920,N_12724);
and U14114 (N_14114,N_12561,N_12578);
xnor U14115 (N_14115,N_12710,N_12344);
nor U14116 (N_14116,N_12596,N_13032);
and U14117 (N_14117,N_13060,N_12608);
xor U14118 (N_14118,N_12867,N_12149);
and U14119 (N_14119,N_13366,N_12917);
and U14120 (N_14120,N_12504,N_13173);
nand U14121 (N_14121,N_12397,N_13139);
xor U14122 (N_14122,N_13392,N_12959);
and U14123 (N_14123,N_12553,N_12434);
and U14124 (N_14124,N_12322,N_12005);
xor U14125 (N_14125,N_13118,N_13073);
or U14126 (N_14126,N_13314,N_13039);
nand U14127 (N_14127,N_13206,N_12168);
nand U14128 (N_14128,N_12341,N_12797);
or U14129 (N_14129,N_13371,N_13215);
or U14130 (N_14130,N_12587,N_12134);
xor U14131 (N_14131,N_13035,N_12887);
xnor U14132 (N_14132,N_12174,N_13075);
nand U14133 (N_14133,N_13106,N_12172);
nand U14134 (N_14134,N_13023,N_12757);
xor U14135 (N_14135,N_12243,N_12061);
nand U14136 (N_14136,N_12478,N_13417);
xnor U14137 (N_14137,N_12156,N_13241);
nor U14138 (N_14138,N_13386,N_12212);
and U14139 (N_14139,N_13356,N_13025);
nand U14140 (N_14140,N_12721,N_12481);
and U14141 (N_14141,N_13472,N_13213);
and U14142 (N_14142,N_13209,N_12106);
nand U14143 (N_14143,N_12295,N_12100);
and U14144 (N_14144,N_13038,N_13465);
and U14145 (N_14145,N_12771,N_13481);
xnor U14146 (N_14146,N_12138,N_12133);
nand U14147 (N_14147,N_12371,N_12363);
nand U14148 (N_14148,N_12294,N_12023);
xnor U14149 (N_14149,N_12523,N_12309);
xor U14150 (N_14150,N_13340,N_13195);
nor U14151 (N_14151,N_12494,N_13268);
nand U14152 (N_14152,N_12659,N_13166);
and U14153 (N_14153,N_12902,N_12372);
or U14154 (N_14154,N_12709,N_13044);
nand U14155 (N_14155,N_12404,N_13428);
or U14156 (N_14156,N_13399,N_13248);
nand U14157 (N_14157,N_12102,N_12650);
xor U14158 (N_14158,N_13123,N_12485);
or U14159 (N_14159,N_12687,N_13250);
nand U14160 (N_14160,N_13191,N_13270);
or U14161 (N_14161,N_12760,N_12870);
nor U14162 (N_14162,N_12200,N_12812);
nand U14163 (N_14163,N_12242,N_12188);
or U14164 (N_14164,N_12557,N_13477);
nor U14165 (N_14165,N_12474,N_12645);
or U14166 (N_14166,N_12787,N_12509);
and U14167 (N_14167,N_13365,N_12909);
or U14168 (N_14168,N_12905,N_13487);
and U14169 (N_14169,N_12947,N_12125);
or U14170 (N_14170,N_12256,N_12889);
or U14171 (N_14171,N_12652,N_12945);
xnor U14172 (N_14172,N_13364,N_13050);
xor U14173 (N_14173,N_12928,N_12103);
xor U14174 (N_14174,N_12946,N_13385);
and U14175 (N_14175,N_13048,N_12629);
nand U14176 (N_14176,N_12925,N_12935);
nand U14177 (N_14177,N_12390,N_13279);
xnor U14178 (N_14178,N_12347,N_12158);
nand U14179 (N_14179,N_12842,N_13381);
nand U14180 (N_14180,N_12712,N_13059);
and U14181 (N_14181,N_12116,N_12542);
or U14182 (N_14182,N_12010,N_12767);
and U14183 (N_14183,N_13350,N_12157);
nand U14184 (N_14184,N_12119,N_12743);
xor U14185 (N_14185,N_13077,N_13406);
or U14186 (N_14186,N_12540,N_12272);
nor U14187 (N_14187,N_13272,N_12013);
nand U14188 (N_14188,N_13335,N_13352);
and U14189 (N_14189,N_13345,N_12772);
or U14190 (N_14190,N_12651,N_12357);
nand U14191 (N_14191,N_13255,N_12499);
nand U14192 (N_14192,N_12683,N_12366);
or U14193 (N_14193,N_12433,N_12380);
nor U14194 (N_14194,N_12087,N_13247);
or U14195 (N_14195,N_12219,N_12081);
nor U14196 (N_14196,N_13294,N_13001);
and U14197 (N_14197,N_12027,N_13102);
or U14198 (N_14198,N_13008,N_12533);
nand U14199 (N_14199,N_13214,N_12122);
or U14200 (N_14200,N_13145,N_12615);
and U14201 (N_14201,N_13289,N_12874);
or U14202 (N_14202,N_13055,N_12266);
nor U14203 (N_14203,N_12976,N_12154);
and U14204 (N_14204,N_13469,N_13253);
and U14205 (N_14205,N_13358,N_12667);
nand U14206 (N_14206,N_12981,N_12538);
or U14207 (N_14207,N_12632,N_12746);
and U14208 (N_14208,N_12254,N_13100);
nor U14209 (N_14209,N_12706,N_13242);
and U14210 (N_14210,N_12193,N_12249);
nor U14211 (N_14211,N_12539,N_12186);
nor U14212 (N_14212,N_12722,N_13319);
nor U14213 (N_14213,N_12943,N_12517);
nor U14214 (N_14214,N_12089,N_13471);
nand U14215 (N_14215,N_13490,N_13066);
nand U14216 (N_14216,N_12079,N_12880);
and U14217 (N_14217,N_12355,N_13416);
nand U14218 (N_14218,N_12996,N_13304);
nand U14219 (N_14219,N_12800,N_12496);
or U14220 (N_14220,N_12312,N_12426);
or U14221 (N_14221,N_12246,N_12449);
and U14222 (N_14222,N_12159,N_12914);
nand U14223 (N_14223,N_12447,N_12284);
and U14224 (N_14224,N_12510,N_13332);
nand U14225 (N_14225,N_12620,N_13108);
nand U14226 (N_14226,N_12518,N_12409);
nand U14227 (N_14227,N_12360,N_13137);
nand U14228 (N_14228,N_13443,N_13230);
nor U14229 (N_14229,N_13290,N_12191);
and U14230 (N_14230,N_12252,N_13037);
xor U14231 (N_14231,N_12697,N_13391);
nand U14232 (N_14232,N_12514,N_12534);
xnor U14233 (N_14233,N_13194,N_13178);
and U14234 (N_14234,N_12085,N_12425);
nand U14235 (N_14235,N_12989,N_13377);
or U14236 (N_14236,N_13162,N_13261);
or U14237 (N_14237,N_12788,N_13124);
and U14238 (N_14238,N_12541,N_12090);
or U14239 (N_14239,N_12438,N_12732);
or U14240 (N_14240,N_12679,N_13007);
nor U14241 (N_14241,N_13149,N_12696);
xor U14242 (N_14242,N_12774,N_13263);
xnor U14243 (N_14243,N_13403,N_12641);
xnor U14244 (N_14244,N_12034,N_13265);
or U14245 (N_14245,N_12450,N_13379);
xor U14246 (N_14246,N_12572,N_12234);
nor U14247 (N_14247,N_12342,N_12223);
nor U14248 (N_14248,N_12353,N_13347);
nor U14249 (N_14249,N_12096,N_13293);
and U14250 (N_14250,N_12410,N_12072);
nor U14251 (N_14251,N_12322,N_12983);
nor U14252 (N_14252,N_12334,N_13307);
nand U14253 (N_14253,N_12815,N_12016);
or U14254 (N_14254,N_12171,N_12693);
or U14255 (N_14255,N_13186,N_12360);
or U14256 (N_14256,N_12146,N_13341);
or U14257 (N_14257,N_12054,N_13082);
or U14258 (N_14258,N_12364,N_13419);
xnor U14259 (N_14259,N_12733,N_12880);
or U14260 (N_14260,N_13220,N_12639);
and U14261 (N_14261,N_13336,N_12475);
nor U14262 (N_14262,N_12999,N_13473);
xor U14263 (N_14263,N_12656,N_12898);
nor U14264 (N_14264,N_13186,N_12073);
xnor U14265 (N_14265,N_13409,N_12345);
and U14266 (N_14266,N_13277,N_12239);
nor U14267 (N_14267,N_12652,N_12273);
xnor U14268 (N_14268,N_12901,N_13104);
xor U14269 (N_14269,N_12697,N_12897);
and U14270 (N_14270,N_13058,N_12186);
or U14271 (N_14271,N_13485,N_12494);
nand U14272 (N_14272,N_12040,N_13404);
nor U14273 (N_14273,N_12260,N_13438);
nor U14274 (N_14274,N_12722,N_12440);
xnor U14275 (N_14275,N_12503,N_13062);
or U14276 (N_14276,N_13383,N_12309);
or U14277 (N_14277,N_13473,N_13495);
nor U14278 (N_14278,N_12863,N_13047);
or U14279 (N_14279,N_12817,N_12513);
nor U14280 (N_14280,N_12699,N_12798);
or U14281 (N_14281,N_12422,N_12364);
and U14282 (N_14282,N_12229,N_13272);
nand U14283 (N_14283,N_13131,N_12534);
xnor U14284 (N_14284,N_12704,N_12605);
xnor U14285 (N_14285,N_13237,N_13400);
nand U14286 (N_14286,N_13289,N_12421);
nand U14287 (N_14287,N_12023,N_13163);
nor U14288 (N_14288,N_13328,N_12738);
nand U14289 (N_14289,N_13093,N_12739);
nor U14290 (N_14290,N_12092,N_13002);
xnor U14291 (N_14291,N_12569,N_12733);
and U14292 (N_14292,N_12578,N_13238);
and U14293 (N_14293,N_13048,N_12743);
nor U14294 (N_14294,N_12423,N_12429);
nor U14295 (N_14295,N_12963,N_12251);
xor U14296 (N_14296,N_13394,N_12937);
or U14297 (N_14297,N_12209,N_13314);
nand U14298 (N_14298,N_12579,N_12611);
xor U14299 (N_14299,N_12188,N_12472);
or U14300 (N_14300,N_12945,N_13433);
xnor U14301 (N_14301,N_13210,N_12814);
or U14302 (N_14302,N_13163,N_12636);
or U14303 (N_14303,N_12832,N_12642);
or U14304 (N_14304,N_13468,N_12192);
nand U14305 (N_14305,N_12843,N_13192);
and U14306 (N_14306,N_13221,N_12046);
nor U14307 (N_14307,N_12188,N_12204);
xor U14308 (N_14308,N_12487,N_12936);
nor U14309 (N_14309,N_12068,N_12444);
or U14310 (N_14310,N_13030,N_12940);
nor U14311 (N_14311,N_12025,N_12702);
and U14312 (N_14312,N_13199,N_13074);
nor U14313 (N_14313,N_13301,N_13033);
and U14314 (N_14314,N_12435,N_12227);
or U14315 (N_14315,N_13462,N_12046);
nand U14316 (N_14316,N_12297,N_12453);
and U14317 (N_14317,N_12699,N_12823);
nor U14318 (N_14318,N_13177,N_12356);
nand U14319 (N_14319,N_13128,N_12986);
and U14320 (N_14320,N_12729,N_12891);
nand U14321 (N_14321,N_12134,N_12390);
nand U14322 (N_14322,N_13404,N_12956);
xor U14323 (N_14323,N_12104,N_12174);
or U14324 (N_14324,N_13150,N_13137);
or U14325 (N_14325,N_13091,N_12875);
or U14326 (N_14326,N_13307,N_12173);
nor U14327 (N_14327,N_13347,N_12766);
nor U14328 (N_14328,N_13390,N_12375);
and U14329 (N_14329,N_13361,N_13086);
or U14330 (N_14330,N_12465,N_12001);
or U14331 (N_14331,N_12650,N_12861);
xnor U14332 (N_14332,N_13276,N_12889);
nand U14333 (N_14333,N_13065,N_13380);
nand U14334 (N_14334,N_12241,N_12311);
xor U14335 (N_14335,N_12724,N_12878);
or U14336 (N_14336,N_12570,N_12266);
xnor U14337 (N_14337,N_12330,N_12987);
xnor U14338 (N_14338,N_12778,N_12722);
nor U14339 (N_14339,N_12178,N_12009);
or U14340 (N_14340,N_13475,N_13425);
nor U14341 (N_14341,N_13124,N_12834);
nor U14342 (N_14342,N_12889,N_12915);
nor U14343 (N_14343,N_12518,N_13119);
and U14344 (N_14344,N_12450,N_12645);
nand U14345 (N_14345,N_12931,N_12264);
xor U14346 (N_14346,N_13121,N_12516);
and U14347 (N_14347,N_12792,N_13130);
and U14348 (N_14348,N_13026,N_12503);
nand U14349 (N_14349,N_12736,N_13022);
or U14350 (N_14350,N_13259,N_12887);
and U14351 (N_14351,N_12976,N_12727);
nor U14352 (N_14352,N_12004,N_13046);
or U14353 (N_14353,N_12445,N_12902);
and U14354 (N_14354,N_12027,N_13473);
and U14355 (N_14355,N_12264,N_12664);
xor U14356 (N_14356,N_12042,N_13005);
and U14357 (N_14357,N_12424,N_12054);
nand U14358 (N_14358,N_12804,N_12539);
nor U14359 (N_14359,N_13495,N_13307);
nor U14360 (N_14360,N_13276,N_12764);
nor U14361 (N_14361,N_13170,N_13423);
nor U14362 (N_14362,N_12549,N_12144);
and U14363 (N_14363,N_12470,N_12375);
or U14364 (N_14364,N_13211,N_13438);
or U14365 (N_14365,N_13068,N_12834);
and U14366 (N_14366,N_12518,N_12694);
nor U14367 (N_14367,N_12001,N_13273);
nor U14368 (N_14368,N_12500,N_12999);
nor U14369 (N_14369,N_13080,N_13425);
or U14370 (N_14370,N_12922,N_12650);
or U14371 (N_14371,N_12827,N_13440);
xnor U14372 (N_14372,N_12983,N_13498);
and U14373 (N_14373,N_12115,N_13001);
xor U14374 (N_14374,N_12503,N_13107);
or U14375 (N_14375,N_12544,N_13166);
nor U14376 (N_14376,N_12068,N_12806);
nor U14377 (N_14377,N_13298,N_13056);
nor U14378 (N_14378,N_12412,N_13462);
or U14379 (N_14379,N_13294,N_12559);
or U14380 (N_14380,N_12201,N_13180);
nand U14381 (N_14381,N_12396,N_12414);
xnor U14382 (N_14382,N_12356,N_12804);
or U14383 (N_14383,N_12602,N_13434);
or U14384 (N_14384,N_12489,N_13211);
or U14385 (N_14385,N_12324,N_12676);
xor U14386 (N_14386,N_12718,N_12713);
nand U14387 (N_14387,N_13028,N_12354);
nor U14388 (N_14388,N_13453,N_12930);
nor U14389 (N_14389,N_12883,N_13002);
nor U14390 (N_14390,N_12649,N_12844);
nand U14391 (N_14391,N_12400,N_13350);
and U14392 (N_14392,N_12585,N_12746);
xnor U14393 (N_14393,N_12209,N_12617);
or U14394 (N_14394,N_12224,N_13168);
nor U14395 (N_14395,N_13159,N_13104);
and U14396 (N_14396,N_12046,N_12979);
and U14397 (N_14397,N_13488,N_12529);
or U14398 (N_14398,N_13216,N_13498);
and U14399 (N_14399,N_12107,N_12892);
xnor U14400 (N_14400,N_12166,N_12682);
and U14401 (N_14401,N_12022,N_12860);
and U14402 (N_14402,N_12237,N_13009);
and U14403 (N_14403,N_12672,N_13474);
or U14404 (N_14404,N_12357,N_12746);
xor U14405 (N_14405,N_12358,N_12264);
or U14406 (N_14406,N_12427,N_12817);
or U14407 (N_14407,N_13232,N_12741);
nand U14408 (N_14408,N_12358,N_12459);
nand U14409 (N_14409,N_13167,N_12347);
nor U14410 (N_14410,N_12119,N_12496);
nor U14411 (N_14411,N_12163,N_12265);
xor U14412 (N_14412,N_13188,N_12695);
nand U14413 (N_14413,N_12108,N_12808);
or U14414 (N_14414,N_12336,N_12509);
and U14415 (N_14415,N_13064,N_12528);
nand U14416 (N_14416,N_13015,N_12995);
and U14417 (N_14417,N_13442,N_12302);
xor U14418 (N_14418,N_12026,N_12823);
and U14419 (N_14419,N_12246,N_12035);
and U14420 (N_14420,N_12897,N_12955);
nor U14421 (N_14421,N_12176,N_13329);
or U14422 (N_14422,N_13067,N_12380);
nor U14423 (N_14423,N_13384,N_12258);
nand U14424 (N_14424,N_12184,N_12215);
nor U14425 (N_14425,N_12584,N_12161);
nor U14426 (N_14426,N_12037,N_13044);
nor U14427 (N_14427,N_13216,N_13277);
or U14428 (N_14428,N_12953,N_13442);
xnor U14429 (N_14429,N_13358,N_12947);
nand U14430 (N_14430,N_13365,N_12160);
nand U14431 (N_14431,N_12186,N_12354);
nor U14432 (N_14432,N_12973,N_12043);
and U14433 (N_14433,N_12130,N_12786);
nand U14434 (N_14434,N_12444,N_12988);
nor U14435 (N_14435,N_13111,N_13388);
nor U14436 (N_14436,N_13250,N_13465);
or U14437 (N_14437,N_12844,N_12535);
or U14438 (N_14438,N_12860,N_12701);
nand U14439 (N_14439,N_13431,N_12017);
xnor U14440 (N_14440,N_12837,N_13398);
nor U14441 (N_14441,N_12364,N_12476);
nand U14442 (N_14442,N_12622,N_12758);
nor U14443 (N_14443,N_13188,N_13416);
and U14444 (N_14444,N_12111,N_12750);
and U14445 (N_14445,N_12564,N_13031);
or U14446 (N_14446,N_12413,N_13055);
and U14447 (N_14447,N_13224,N_12758);
or U14448 (N_14448,N_13178,N_12749);
nor U14449 (N_14449,N_12541,N_12152);
or U14450 (N_14450,N_12830,N_12837);
or U14451 (N_14451,N_12655,N_12391);
xor U14452 (N_14452,N_13236,N_12163);
or U14453 (N_14453,N_12918,N_13138);
and U14454 (N_14454,N_12644,N_12584);
xor U14455 (N_14455,N_12130,N_12302);
and U14456 (N_14456,N_12850,N_13489);
nand U14457 (N_14457,N_12863,N_12178);
or U14458 (N_14458,N_12878,N_12310);
nor U14459 (N_14459,N_12710,N_13405);
nand U14460 (N_14460,N_12429,N_13172);
or U14461 (N_14461,N_12920,N_12830);
and U14462 (N_14462,N_12883,N_12117);
and U14463 (N_14463,N_12563,N_12153);
xor U14464 (N_14464,N_12959,N_13328);
and U14465 (N_14465,N_12340,N_12111);
or U14466 (N_14466,N_12729,N_13479);
or U14467 (N_14467,N_12091,N_12644);
and U14468 (N_14468,N_12857,N_13440);
xor U14469 (N_14469,N_13065,N_12133);
or U14470 (N_14470,N_13122,N_12226);
nand U14471 (N_14471,N_12151,N_12487);
xor U14472 (N_14472,N_12803,N_12439);
or U14473 (N_14473,N_13131,N_12448);
nand U14474 (N_14474,N_12250,N_12738);
xor U14475 (N_14475,N_12873,N_12378);
or U14476 (N_14476,N_13201,N_13267);
xnor U14477 (N_14477,N_13081,N_12726);
nand U14478 (N_14478,N_12195,N_12738);
xnor U14479 (N_14479,N_12319,N_13320);
xor U14480 (N_14480,N_13190,N_12509);
or U14481 (N_14481,N_12734,N_13020);
or U14482 (N_14482,N_12813,N_13236);
xor U14483 (N_14483,N_13280,N_12524);
nor U14484 (N_14484,N_13474,N_13118);
nor U14485 (N_14485,N_12786,N_13306);
nor U14486 (N_14486,N_13195,N_12736);
nand U14487 (N_14487,N_12362,N_12341);
nor U14488 (N_14488,N_12568,N_12794);
or U14489 (N_14489,N_12948,N_13154);
nand U14490 (N_14490,N_12565,N_13078);
or U14491 (N_14491,N_12581,N_13393);
or U14492 (N_14492,N_12558,N_12451);
nand U14493 (N_14493,N_12634,N_12636);
nand U14494 (N_14494,N_12559,N_12726);
or U14495 (N_14495,N_13318,N_12520);
or U14496 (N_14496,N_12963,N_12231);
or U14497 (N_14497,N_12436,N_12001);
xnor U14498 (N_14498,N_13341,N_12586);
or U14499 (N_14499,N_12089,N_12240);
or U14500 (N_14500,N_12176,N_12829);
nor U14501 (N_14501,N_12459,N_12889);
xor U14502 (N_14502,N_12424,N_12458);
nand U14503 (N_14503,N_12707,N_12723);
or U14504 (N_14504,N_13356,N_13158);
nand U14505 (N_14505,N_13187,N_13320);
nor U14506 (N_14506,N_12699,N_12753);
nand U14507 (N_14507,N_12782,N_12291);
nand U14508 (N_14508,N_12028,N_12431);
and U14509 (N_14509,N_13439,N_12285);
nand U14510 (N_14510,N_12563,N_12258);
and U14511 (N_14511,N_12086,N_13296);
nor U14512 (N_14512,N_12084,N_13232);
and U14513 (N_14513,N_12332,N_12982);
and U14514 (N_14514,N_13308,N_12286);
or U14515 (N_14515,N_12361,N_13088);
nor U14516 (N_14516,N_12578,N_12845);
or U14517 (N_14517,N_12719,N_13056);
nor U14518 (N_14518,N_12168,N_12018);
nand U14519 (N_14519,N_12085,N_13209);
xor U14520 (N_14520,N_12700,N_13005);
or U14521 (N_14521,N_12648,N_12182);
and U14522 (N_14522,N_12421,N_12252);
and U14523 (N_14523,N_12131,N_12941);
nand U14524 (N_14524,N_13436,N_12555);
xor U14525 (N_14525,N_12499,N_13156);
nand U14526 (N_14526,N_13176,N_12221);
xor U14527 (N_14527,N_13486,N_12072);
xor U14528 (N_14528,N_12133,N_12584);
or U14529 (N_14529,N_12683,N_12739);
or U14530 (N_14530,N_12735,N_13072);
or U14531 (N_14531,N_12111,N_12807);
nand U14532 (N_14532,N_12187,N_13461);
nor U14533 (N_14533,N_12140,N_13144);
and U14534 (N_14534,N_13142,N_12665);
and U14535 (N_14535,N_13112,N_12123);
nand U14536 (N_14536,N_13160,N_12515);
nand U14537 (N_14537,N_12484,N_13318);
or U14538 (N_14538,N_12543,N_12489);
and U14539 (N_14539,N_12521,N_12729);
xnor U14540 (N_14540,N_12129,N_12636);
or U14541 (N_14541,N_12296,N_13089);
nor U14542 (N_14542,N_13096,N_13137);
and U14543 (N_14543,N_12733,N_13414);
and U14544 (N_14544,N_12977,N_12337);
and U14545 (N_14545,N_12135,N_12188);
xor U14546 (N_14546,N_13467,N_13095);
xnor U14547 (N_14547,N_12318,N_13015);
and U14548 (N_14548,N_13331,N_13329);
nand U14549 (N_14549,N_13304,N_12561);
nand U14550 (N_14550,N_12992,N_12120);
nor U14551 (N_14551,N_12973,N_12726);
or U14552 (N_14552,N_13225,N_13446);
nand U14553 (N_14553,N_12451,N_12333);
nor U14554 (N_14554,N_12049,N_12679);
or U14555 (N_14555,N_12553,N_12023);
and U14556 (N_14556,N_12977,N_12433);
xnor U14557 (N_14557,N_13432,N_13196);
nand U14558 (N_14558,N_13319,N_12309);
or U14559 (N_14559,N_12772,N_13232);
and U14560 (N_14560,N_12145,N_12105);
and U14561 (N_14561,N_13210,N_12411);
or U14562 (N_14562,N_13253,N_13337);
xnor U14563 (N_14563,N_13479,N_13024);
or U14564 (N_14564,N_12048,N_12193);
nor U14565 (N_14565,N_12867,N_13487);
xor U14566 (N_14566,N_12613,N_12018);
nand U14567 (N_14567,N_12953,N_13324);
or U14568 (N_14568,N_12859,N_12586);
or U14569 (N_14569,N_13090,N_13203);
or U14570 (N_14570,N_12872,N_12922);
and U14571 (N_14571,N_12424,N_13170);
xnor U14572 (N_14572,N_12764,N_12027);
and U14573 (N_14573,N_12123,N_13276);
nand U14574 (N_14574,N_12746,N_12183);
nand U14575 (N_14575,N_13459,N_12646);
xnor U14576 (N_14576,N_12734,N_12190);
nor U14577 (N_14577,N_12563,N_12113);
or U14578 (N_14578,N_13191,N_12126);
nand U14579 (N_14579,N_12348,N_12539);
nor U14580 (N_14580,N_13160,N_13299);
nor U14581 (N_14581,N_13142,N_13238);
nor U14582 (N_14582,N_13021,N_12427);
or U14583 (N_14583,N_12927,N_12110);
xnor U14584 (N_14584,N_12070,N_12217);
nor U14585 (N_14585,N_12050,N_13124);
xnor U14586 (N_14586,N_13078,N_12545);
or U14587 (N_14587,N_12424,N_12556);
xor U14588 (N_14588,N_12199,N_13425);
and U14589 (N_14589,N_13411,N_12930);
nor U14590 (N_14590,N_12682,N_12081);
and U14591 (N_14591,N_13131,N_12041);
or U14592 (N_14592,N_13378,N_12721);
or U14593 (N_14593,N_12955,N_12337);
xor U14594 (N_14594,N_12526,N_12617);
or U14595 (N_14595,N_12799,N_12286);
nor U14596 (N_14596,N_13235,N_13200);
and U14597 (N_14597,N_12472,N_12989);
nand U14598 (N_14598,N_12879,N_13294);
xor U14599 (N_14599,N_13229,N_12027);
nor U14600 (N_14600,N_12619,N_12669);
xnor U14601 (N_14601,N_12062,N_12345);
and U14602 (N_14602,N_12094,N_12486);
and U14603 (N_14603,N_13435,N_12790);
nand U14604 (N_14604,N_12399,N_13020);
and U14605 (N_14605,N_13289,N_12711);
and U14606 (N_14606,N_13473,N_12121);
nand U14607 (N_14607,N_12701,N_12641);
nand U14608 (N_14608,N_13462,N_13430);
xnor U14609 (N_14609,N_12840,N_12754);
or U14610 (N_14610,N_13125,N_12268);
nor U14611 (N_14611,N_12992,N_12196);
nor U14612 (N_14612,N_12954,N_12928);
nand U14613 (N_14613,N_12408,N_12120);
or U14614 (N_14614,N_13143,N_12421);
and U14615 (N_14615,N_12829,N_12413);
nand U14616 (N_14616,N_12053,N_12838);
nor U14617 (N_14617,N_12992,N_13129);
nor U14618 (N_14618,N_12457,N_12467);
nand U14619 (N_14619,N_12123,N_13272);
nand U14620 (N_14620,N_12911,N_12219);
nor U14621 (N_14621,N_12902,N_12591);
nand U14622 (N_14622,N_12601,N_12931);
nor U14623 (N_14623,N_13036,N_12817);
nor U14624 (N_14624,N_13278,N_13346);
nand U14625 (N_14625,N_13230,N_12273);
nor U14626 (N_14626,N_13211,N_13320);
xnor U14627 (N_14627,N_12587,N_12941);
nand U14628 (N_14628,N_13053,N_12850);
nor U14629 (N_14629,N_12008,N_13296);
and U14630 (N_14630,N_12030,N_12196);
or U14631 (N_14631,N_12766,N_12774);
nor U14632 (N_14632,N_13149,N_13374);
xor U14633 (N_14633,N_12846,N_12135);
nor U14634 (N_14634,N_12819,N_12634);
nand U14635 (N_14635,N_12929,N_12820);
nand U14636 (N_14636,N_13389,N_12293);
and U14637 (N_14637,N_12043,N_12590);
nor U14638 (N_14638,N_12116,N_12894);
nand U14639 (N_14639,N_13419,N_13312);
and U14640 (N_14640,N_12624,N_12610);
nor U14641 (N_14641,N_12865,N_12522);
or U14642 (N_14642,N_12132,N_12147);
and U14643 (N_14643,N_12582,N_12201);
xnor U14644 (N_14644,N_12739,N_12219);
nor U14645 (N_14645,N_12318,N_13162);
nand U14646 (N_14646,N_12486,N_12491);
xnor U14647 (N_14647,N_12187,N_12258);
nand U14648 (N_14648,N_13277,N_13248);
xor U14649 (N_14649,N_13222,N_12438);
xnor U14650 (N_14650,N_12341,N_12359);
nand U14651 (N_14651,N_12098,N_13288);
nor U14652 (N_14652,N_13293,N_12568);
or U14653 (N_14653,N_12022,N_12863);
xor U14654 (N_14654,N_13147,N_13085);
nand U14655 (N_14655,N_13436,N_12987);
and U14656 (N_14656,N_12656,N_12126);
xnor U14657 (N_14657,N_12900,N_12093);
nor U14658 (N_14658,N_12269,N_12933);
xnor U14659 (N_14659,N_12499,N_13146);
and U14660 (N_14660,N_12351,N_12710);
and U14661 (N_14661,N_12625,N_12770);
and U14662 (N_14662,N_12993,N_12845);
and U14663 (N_14663,N_13445,N_13472);
nor U14664 (N_14664,N_12224,N_12264);
nand U14665 (N_14665,N_12950,N_12540);
and U14666 (N_14666,N_13218,N_12341);
or U14667 (N_14667,N_13129,N_12282);
nand U14668 (N_14668,N_12132,N_12198);
and U14669 (N_14669,N_12024,N_12033);
or U14670 (N_14670,N_12395,N_12775);
and U14671 (N_14671,N_13288,N_12996);
nor U14672 (N_14672,N_13243,N_12149);
or U14673 (N_14673,N_13326,N_13309);
and U14674 (N_14674,N_13402,N_12375);
xor U14675 (N_14675,N_12576,N_12388);
or U14676 (N_14676,N_13361,N_12491);
or U14677 (N_14677,N_12458,N_12617);
xnor U14678 (N_14678,N_13127,N_13285);
xor U14679 (N_14679,N_12642,N_12317);
and U14680 (N_14680,N_13383,N_12982);
or U14681 (N_14681,N_13358,N_12920);
or U14682 (N_14682,N_12211,N_12652);
or U14683 (N_14683,N_13202,N_12462);
nand U14684 (N_14684,N_13450,N_12975);
nand U14685 (N_14685,N_13394,N_12702);
or U14686 (N_14686,N_13042,N_13458);
or U14687 (N_14687,N_13026,N_12448);
xnor U14688 (N_14688,N_13038,N_12127);
xor U14689 (N_14689,N_12562,N_12442);
nor U14690 (N_14690,N_13369,N_13135);
nand U14691 (N_14691,N_13446,N_12818);
xor U14692 (N_14692,N_13187,N_12785);
nand U14693 (N_14693,N_12633,N_12764);
nand U14694 (N_14694,N_12403,N_12375);
and U14695 (N_14695,N_12627,N_12952);
nand U14696 (N_14696,N_12636,N_12561);
xnor U14697 (N_14697,N_13252,N_12525);
and U14698 (N_14698,N_13230,N_12094);
or U14699 (N_14699,N_13239,N_12346);
nor U14700 (N_14700,N_12101,N_12349);
or U14701 (N_14701,N_12269,N_12083);
nor U14702 (N_14702,N_12454,N_13055);
xnor U14703 (N_14703,N_12210,N_12199);
or U14704 (N_14704,N_12102,N_13321);
xnor U14705 (N_14705,N_12671,N_12350);
nor U14706 (N_14706,N_12819,N_12832);
nor U14707 (N_14707,N_12372,N_12976);
or U14708 (N_14708,N_13474,N_12697);
nand U14709 (N_14709,N_13314,N_12781);
and U14710 (N_14710,N_12869,N_12170);
nor U14711 (N_14711,N_13196,N_12695);
or U14712 (N_14712,N_13075,N_12971);
nor U14713 (N_14713,N_12608,N_12257);
and U14714 (N_14714,N_13179,N_12076);
xnor U14715 (N_14715,N_12493,N_12137);
nor U14716 (N_14716,N_13158,N_12446);
nor U14717 (N_14717,N_13457,N_13066);
nor U14718 (N_14718,N_13363,N_12997);
and U14719 (N_14719,N_12056,N_12916);
xnor U14720 (N_14720,N_13294,N_12336);
xor U14721 (N_14721,N_12158,N_12567);
and U14722 (N_14722,N_13298,N_12134);
or U14723 (N_14723,N_13426,N_12001);
nor U14724 (N_14724,N_12682,N_12610);
and U14725 (N_14725,N_12827,N_12369);
and U14726 (N_14726,N_12798,N_12631);
and U14727 (N_14727,N_12308,N_12874);
nor U14728 (N_14728,N_12739,N_12835);
nor U14729 (N_14729,N_12204,N_12995);
nor U14730 (N_14730,N_12894,N_12541);
nand U14731 (N_14731,N_13481,N_12411);
xnor U14732 (N_14732,N_12781,N_13155);
nand U14733 (N_14733,N_13076,N_13209);
nor U14734 (N_14734,N_12211,N_12900);
xnor U14735 (N_14735,N_12394,N_13087);
and U14736 (N_14736,N_13120,N_12486);
nor U14737 (N_14737,N_12839,N_12177);
nand U14738 (N_14738,N_12142,N_12554);
or U14739 (N_14739,N_13497,N_12907);
or U14740 (N_14740,N_13089,N_12956);
and U14741 (N_14741,N_12158,N_13168);
or U14742 (N_14742,N_12986,N_13378);
and U14743 (N_14743,N_12987,N_12820);
or U14744 (N_14744,N_13243,N_13050);
xnor U14745 (N_14745,N_13463,N_13488);
nand U14746 (N_14746,N_13319,N_12257);
nand U14747 (N_14747,N_12987,N_12467);
and U14748 (N_14748,N_12962,N_12677);
nor U14749 (N_14749,N_12184,N_12765);
and U14750 (N_14750,N_12113,N_12446);
and U14751 (N_14751,N_13097,N_13137);
xor U14752 (N_14752,N_13201,N_12061);
or U14753 (N_14753,N_12513,N_12944);
xnor U14754 (N_14754,N_13309,N_12662);
or U14755 (N_14755,N_12450,N_13033);
nor U14756 (N_14756,N_13351,N_12479);
nand U14757 (N_14757,N_12310,N_12157);
or U14758 (N_14758,N_12455,N_13214);
xnor U14759 (N_14759,N_12971,N_12720);
xor U14760 (N_14760,N_12004,N_13136);
nor U14761 (N_14761,N_12652,N_12360);
or U14762 (N_14762,N_12603,N_12772);
or U14763 (N_14763,N_13104,N_13079);
or U14764 (N_14764,N_13487,N_12541);
nand U14765 (N_14765,N_12837,N_13079);
nand U14766 (N_14766,N_13470,N_12961);
or U14767 (N_14767,N_13096,N_13076);
and U14768 (N_14768,N_12987,N_12727);
nor U14769 (N_14769,N_12315,N_12338);
nand U14770 (N_14770,N_13441,N_12106);
nand U14771 (N_14771,N_12523,N_13027);
xor U14772 (N_14772,N_12358,N_12311);
and U14773 (N_14773,N_12049,N_13045);
xor U14774 (N_14774,N_12828,N_12473);
nand U14775 (N_14775,N_13420,N_12728);
xor U14776 (N_14776,N_12820,N_13179);
nor U14777 (N_14777,N_12875,N_12220);
nor U14778 (N_14778,N_12025,N_12679);
and U14779 (N_14779,N_12221,N_12049);
nor U14780 (N_14780,N_12015,N_12678);
nand U14781 (N_14781,N_13179,N_12711);
nor U14782 (N_14782,N_12350,N_12082);
nand U14783 (N_14783,N_13257,N_12398);
nand U14784 (N_14784,N_13210,N_13416);
and U14785 (N_14785,N_12926,N_12594);
nor U14786 (N_14786,N_12935,N_12803);
xnor U14787 (N_14787,N_13095,N_12193);
nor U14788 (N_14788,N_12190,N_12207);
and U14789 (N_14789,N_12582,N_12287);
and U14790 (N_14790,N_12273,N_12457);
nand U14791 (N_14791,N_13339,N_12430);
nor U14792 (N_14792,N_13172,N_12692);
or U14793 (N_14793,N_13072,N_12997);
nand U14794 (N_14794,N_13430,N_12730);
xnor U14795 (N_14795,N_12407,N_12665);
and U14796 (N_14796,N_12806,N_13117);
and U14797 (N_14797,N_12706,N_12761);
and U14798 (N_14798,N_12418,N_13467);
nand U14799 (N_14799,N_12229,N_12488);
nand U14800 (N_14800,N_12806,N_12454);
and U14801 (N_14801,N_13269,N_13330);
nor U14802 (N_14802,N_12475,N_13473);
nand U14803 (N_14803,N_13192,N_13246);
and U14804 (N_14804,N_13382,N_13304);
nand U14805 (N_14805,N_13119,N_13411);
or U14806 (N_14806,N_13126,N_12018);
nor U14807 (N_14807,N_12667,N_13445);
and U14808 (N_14808,N_12272,N_12561);
and U14809 (N_14809,N_12655,N_12328);
xnor U14810 (N_14810,N_13343,N_12411);
nand U14811 (N_14811,N_12197,N_13431);
xnor U14812 (N_14812,N_12866,N_12714);
nand U14813 (N_14813,N_13094,N_13323);
or U14814 (N_14814,N_12827,N_12325);
nand U14815 (N_14815,N_12002,N_13306);
and U14816 (N_14816,N_13155,N_12822);
nand U14817 (N_14817,N_13072,N_12307);
or U14818 (N_14818,N_12934,N_13411);
xor U14819 (N_14819,N_12638,N_12568);
nor U14820 (N_14820,N_13288,N_12088);
nor U14821 (N_14821,N_12072,N_13077);
and U14822 (N_14822,N_13432,N_12950);
xor U14823 (N_14823,N_13019,N_12943);
and U14824 (N_14824,N_12089,N_13016);
and U14825 (N_14825,N_13488,N_12517);
nor U14826 (N_14826,N_12262,N_12837);
xnor U14827 (N_14827,N_13116,N_12709);
nor U14828 (N_14828,N_12760,N_13041);
nand U14829 (N_14829,N_12616,N_12497);
nand U14830 (N_14830,N_12915,N_13016);
and U14831 (N_14831,N_12166,N_12292);
and U14832 (N_14832,N_12510,N_13108);
nor U14833 (N_14833,N_12823,N_13316);
xor U14834 (N_14834,N_12230,N_13429);
nand U14835 (N_14835,N_13297,N_12565);
nand U14836 (N_14836,N_12522,N_13395);
nand U14837 (N_14837,N_13158,N_13399);
and U14838 (N_14838,N_12449,N_12584);
or U14839 (N_14839,N_13329,N_13101);
or U14840 (N_14840,N_13027,N_12453);
nand U14841 (N_14841,N_13171,N_12218);
or U14842 (N_14842,N_13027,N_12881);
nand U14843 (N_14843,N_12178,N_12096);
nor U14844 (N_14844,N_13257,N_12204);
or U14845 (N_14845,N_12156,N_12603);
and U14846 (N_14846,N_12268,N_12563);
and U14847 (N_14847,N_13416,N_13071);
and U14848 (N_14848,N_12737,N_13468);
nor U14849 (N_14849,N_12038,N_12566);
nand U14850 (N_14850,N_13442,N_12211);
xnor U14851 (N_14851,N_12473,N_12987);
and U14852 (N_14852,N_12212,N_13468);
and U14853 (N_14853,N_13452,N_13286);
nor U14854 (N_14854,N_13364,N_12085);
nand U14855 (N_14855,N_13385,N_13069);
or U14856 (N_14856,N_12209,N_13009);
nand U14857 (N_14857,N_12590,N_13059);
and U14858 (N_14858,N_12355,N_13167);
xor U14859 (N_14859,N_12151,N_12236);
nand U14860 (N_14860,N_12691,N_12954);
and U14861 (N_14861,N_12239,N_13469);
nand U14862 (N_14862,N_13373,N_12857);
xor U14863 (N_14863,N_12301,N_13481);
nand U14864 (N_14864,N_12872,N_13217);
or U14865 (N_14865,N_13348,N_12286);
or U14866 (N_14866,N_13496,N_12783);
or U14867 (N_14867,N_12920,N_12513);
nand U14868 (N_14868,N_13327,N_13176);
or U14869 (N_14869,N_12857,N_12119);
and U14870 (N_14870,N_12859,N_13069);
or U14871 (N_14871,N_12335,N_12792);
xnor U14872 (N_14872,N_12486,N_12476);
nor U14873 (N_14873,N_12365,N_12209);
nor U14874 (N_14874,N_12579,N_12146);
or U14875 (N_14875,N_13131,N_12856);
nand U14876 (N_14876,N_12902,N_12906);
nand U14877 (N_14877,N_13224,N_12900);
and U14878 (N_14878,N_12790,N_12474);
or U14879 (N_14879,N_12893,N_12845);
and U14880 (N_14880,N_13058,N_12360);
xnor U14881 (N_14881,N_12803,N_12048);
or U14882 (N_14882,N_12069,N_12019);
or U14883 (N_14883,N_12024,N_12550);
nand U14884 (N_14884,N_13277,N_12965);
xor U14885 (N_14885,N_13007,N_12294);
or U14886 (N_14886,N_13479,N_12439);
and U14887 (N_14887,N_13150,N_12656);
or U14888 (N_14888,N_12686,N_12143);
or U14889 (N_14889,N_12224,N_12517);
nor U14890 (N_14890,N_12314,N_13004);
or U14891 (N_14891,N_13145,N_12316);
xor U14892 (N_14892,N_12346,N_12390);
nor U14893 (N_14893,N_13427,N_12775);
xnor U14894 (N_14894,N_13190,N_13064);
nand U14895 (N_14895,N_13326,N_13499);
and U14896 (N_14896,N_12622,N_12515);
nand U14897 (N_14897,N_13345,N_13102);
nor U14898 (N_14898,N_13154,N_12764);
xnor U14899 (N_14899,N_12565,N_12002);
xor U14900 (N_14900,N_13476,N_12185);
nor U14901 (N_14901,N_12124,N_12364);
or U14902 (N_14902,N_12745,N_12649);
nor U14903 (N_14903,N_12498,N_13181);
nor U14904 (N_14904,N_12957,N_13085);
nor U14905 (N_14905,N_12127,N_12198);
and U14906 (N_14906,N_12062,N_12954);
and U14907 (N_14907,N_12547,N_13336);
and U14908 (N_14908,N_13399,N_12777);
or U14909 (N_14909,N_13347,N_12828);
nand U14910 (N_14910,N_12863,N_13020);
nand U14911 (N_14911,N_12815,N_12082);
xor U14912 (N_14912,N_13033,N_12022);
xnor U14913 (N_14913,N_13485,N_12998);
nor U14914 (N_14914,N_12660,N_12234);
xnor U14915 (N_14915,N_12491,N_12648);
and U14916 (N_14916,N_12542,N_12449);
or U14917 (N_14917,N_13070,N_12229);
and U14918 (N_14918,N_12915,N_13310);
or U14919 (N_14919,N_13430,N_12547);
and U14920 (N_14920,N_13148,N_12865);
or U14921 (N_14921,N_12446,N_12866);
nand U14922 (N_14922,N_13421,N_12801);
xor U14923 (N_14923,N_12099,N_12051);
and U14924 (N_14924,N_13177,N_12064);
xnor U14925 (N_14925,N_12271,N_12416);
nor U14926 (N_14926,N_12135,N_13348);
or U14927 (N_14927,N_12619,N_12009);
nor U14928 (N_14928,N_12586,N_12448);
xnor U14929 (N_14929,N_12093,N_12357);
xnor U14930 (N_14930,N_12878,N_12222);
nor U14931 (N_14931,N_13021,N_13034);
or U14932 (N_14932,N_12748,N_12066);
and U14933 (N_14933,N_12414,N_12678);
or U14934 (N_14934,N_12609,N_13366);
and U14935 (N_14935,N_12373,N_12116);
and U14936 (N_14936,N_13267,N_12849);
nor U14937 (N_14937,N_12740,N_13119);
nor U14938 (N_14938,N_12128,N_12367);
and U14939 (N_14939,N_12562,N_12694);
and U14940 (N_14940,N_12636,N_12695);
and U14941 (N_14941,N_12791,N_12675);
or U14942 (N_14942,N_13277,N_13213);
nor U14943 (N_14943,N_13032,N_12145);
nand U14944 (N_14944,N_13015,N_12291);
and U14945 (N_14945,N_13388,N_12541);
nor U14946 (N_14946,N_12924,N_12535);
xor U14947 (N_14947,N_13121,N_12542);
or U14948 (N_14948,N_12096,N_13080);
nor U14949 (N_14949,N_12015,N_13198);
nand U14950 (N_14950,N_12777,N_12984);
nand U14951 (N_14951,N_12831,N_12710);
nand U14952 (N_14952,N_13065,N_12295);
nand U14953 (N_14953,N_12589,N_13160);
xor U14954 (N_14954,N_12460,N_12528);
xnor U14955 (N_14955,N_12203,N_12293);
nor U14956 (N_14956,N_12177,N_12014);
or U14957 (N_14957,N_12261,N_12929);
nor U14958 (N_14958,N_12125,N_13361);
nor U14959 (N_14959,N_12413,N_13091);
and U14960 (N_14960,N_12336,N_12162);
nor U14961 (N_14961,N_13397,N_13465);
and U14962 (N_14962,N_12219,N_12131);
nand U14963 (N_14963,N_13293,N_13047);
nand U14964 (N_14964,N_13183,N_13264);
xnor U14965 (N_14965,N_12310,N_12350);
and U14966 (N_14966,N_12804,N_13479);
nand U14967 (N_14967,N_13326,N_12772);
and U14968 (N_14968,N_12074,N_12809);
xor U14969 (N_14969,N_12287,N_12172);
nor U14970 (N_14970,N_13185,N_12815);
nor U14971 (N_14971,N_12601,N_12160);
and U14972 (N_14972,N_12846,N_12305);
nor U14973 (N_14973,N_13132,N_13298);
xnor U14974 (N_14974,N_13119,N_12166);
and U14975 (N_14975,N_12822,N_13396);
xor U14976 (N_14976,N_12116,N_13354);
or U14977 (N_14977,N_12854,N_12275);
xnor U14978 (N_14978,N_13260,N_12374);
xnor U14979 (N_14979,N_12950,N_12543);
and U14980 (N_14980,N_13294,N_13444);
nor U14981 (N_14981,N_12070,N_12907);
nand U14982 (N_14982,N_12040,N_13056);
xnor U14983 (N_14983,N_12055,N_12412);
xnor U14984 (N_14984,N_12975,N_13271);
nor U14985 (N_14985,N_12779,N_12693);
or U14986 (N_14986,N_12479,N_12660);
and U14987 (N_14987,N_12909,N_13175);
nor U14988 (N_14988,N_12157,N_12390);
or U14989 (N_14989,N_12543,N_12185);
nor U14990 (N_14990,N_12617,N_12461);
nor U14991 (N_14991,N_12226,N_13410);
or U14992 (N_14992,N_12097,N_12362);
and U14993 (N_14993,N_12178,N_12348);
nand U14994 (N_14994,N_13135,N_12735);
xor U14995 (N_14995,N_13221,N_12676);
xnor U14996 (N_14996,N_12294,N_12389);
and U14997 (N_14997,N_13362,N_12085);
xor U14998 (N_14998,N_12242,N_13352);
nor U14999 (N_14999,N_12782,N_12484);
or UO_0 (O_0,N_14354,N_14522);
nor UO_1 (O_1,N_13573,N_14271);
nor UO_2 (O_2,N_14793,N_14349);
nor UO_3 (O_3,N_13776,N_14829);
and UO_4 (O_4,N_14119,N_13762);
nor UO_5 (O_5,N_13992,N_13564);
and UO_6 (O_6,N_14079,N_14238);
nand UO_7 (O_7,N_14042,N_13753);
nor UO_8 (O_8,N_14671,N_14039);
nor UO_9 (O_9,N_13632,N_13526);
or UO_10 (O_10,N_14732,N_14748);
xor UO_11 (O_11,N_14987,N_14853);
and UO_12 (O_12,N_14951,N_14610);
xor UO_13 (O_13,N_13706,N_14935);
nor UO_14 (O_14,N_13689,N_14067);
and UO_15 (O_15,N_14063,N_14364);
xor UO_16 (O_16,N_13915,N_13543);
nor UO_17 (O_17,N_13590,N_14996);
or UO_18 (O_18,N_14177,N_13935);
and UO_19 (O_19,N_14579,N_13880);
or UO_20 (O_20,N_14554,N_14778);
nor UO_21 (O_21,N_13549,N_14415);
xnor UO_22 (O_22,N_14991,N_13922);
nand UO_23 (O_23,N_14603,N_14241);
nand UO_24 (O_24,N_14166,N_14841);
nand UO_25 (O_25,N_14871,N_14561);
or UO_26 (O_26,N_14879,N_14002);
or UO_27 (O_27,N_14792,N_13875);
or UO_28 (O_28,N_14993,N_14453);
nand UO_29 (O_29,N_14282,N_14151);
and UO_30 (O_30,N_14441,N_13657);
or UO_31 (O_31,N_14660,N_14198);
and UO_32 (O_32,N_14806,N_14190);
xnor UO_33 (O_33,N_14494,N_13997);
nand UO_34 (O_34,N_14967,N_13783);
xor UO_35 (O_35,N_14051,N_14308);
xnor UO_36 (O_36,N_13606,N_13866);
xor UO_37 (O_37,N_14008,N_13594);
or UO_38 (O_38,N_14287,N_14585);
and UO_39 (O_39,N_14304,N_13629);
xnor UO_40 (O_40,N_13546,N_13605);
or UO_41 (O_41,N_14673,N_14280);
or UO_42 (O_42,N_14722,N_14962);
nand UO_43 (O_43,N_13509,N_13604);
and UO_44 (O_44,N_13624,N_14680);
xor UO_45 (O_45,N_14390,N_14456);
and UO_46 (O_46,N_13799,N_14694);
nand UO_47 (O_47,N_14399,N_14046);
and UO_48 (O_48,N_13775,N_13717);
xor UO_49 (O_49,N_13570,N_13773);
nand UO_50 (O_50,N_13533,N_13741);
or UO_51 (O_51,N_14716,N_14633);
nor UO_52 (O_52,N_14977,N_13530);
and UO_53 (O_53,N_14614,N_14837);
and UO_54 (O_54,N_13868,N_14139);
nand UO_55 (O_55,N_13884,N_14122);
nor UO_56 (O_56,N_13987,N_13595);
and UO_57 (O_57,N_14362,N_14876);
xnor UO_58 (O_58,N_14222,N_14847);
nand UO_59 (O_59,N_14896,N_14616);
xor UO_60 (O_60,N_14725,N_14321);
and UO_61 (O_61,N_14875,N_14358);
xor UO_62 (O_62,N_14500,N_13758);
and UO_63 (O_63,N_13575,N_14677);
xor UO_64 (O_64,N_13644,N_13923);
and UO_65 (O_65,N_13821,N_13557);
nor UO_66 (O_66,N_14934,N_14767);
nor UO_67 (O_67,N_14164,N_14484);
or UO_68 (O_68,N_14517,N_13619);
nor UO_69 (O_69,N_14467,N_13610);
nor UO_70 (O_70,N_14104,N_14918);
nand UO_71 (O_71,N_13983,N_14638);
and UO_72 (O_72,N_14314,N_14857);
and UO_73 (O_73,N_14683,N_14531);
nor UO_74 (O_74,N_14734,N_14943);
or UO_75 (O_75,N_13695,N_14931);
or UO_76 (O_76,N_13791,N_14325);
and UO_77 (O_77,N_14376,N_14626);
nand UO_78 (O_78,N_14125,N_13804);
nor UO_79 (O_79,N_14604,N_13505);
xor UO_80 (O_80,N_14503,N_13842);
or UO_81 (O_81,N_14232,N_13643);
and UO_82 (O_82,N_13609,N_14634);
nand UO_83 (O_83,N_14632,N_14985);
or UO_84 (O_84,N_14518,N_14773);
xor UO_85 (O_85,N_13906,N_13954);
nor UO_86 (O_86,N_14450,N_14592);
nor UO_87 (O_87,N_14299,N_13955);
nor UO_88 (O_88,N_13951,N_13944);
or UO_89 (O_89,N_14091,N_14652);
xnor UO_90 (O_90,N_13535,N_14499);
or UO_91 (O_91,N_14455,N_14403);
nor UO_92 (O_92,N_13539,N_13646);
and UO_93 (O_93,N_14726,N_14012);
nor UO_94 (O_94,N_14435,N_13919);
xor UO_95 (O_95,N_13810,N_14609);
nor UO_96 (O_96,N_14893,N_13611);
xnor UO_97 (O_97,N_13928,N_14075);
nor UO_98 (O_98,N_14662,N_13642);
xor UO_99 (O_99,N_14537,N_13903);
xnor UO_100 (O_100,N_14410,N_14463);
nand UO_101 (O_101,N_14261,N_14318);
nand UO_102 (O_102,N_13649,N_14252);
nand UO_103 (O_103,N_14307,N_14586);
xnor UO_104 (O_104,N_14718,N_14440);
and UO_105 (O_105,N_14698,N_14229);
nand UO_106 (O_106,N_14926,N_14345);
xnor UO_107 (O_107,N_14197,N_13542);
nand UO_108 (O_108,N_14711,N_14708);
nand UO_109 (O_109,N_13692,N_13978);
xor UO_110 (O_110,N_14451,N_13559);
nor UO_111 (O_111,N_14393,N_14955);
nand UO_112 (O_112,N_13713,N_13973);
nand UO_113 (O_113,N_13628,N_14940);
or UO_114 (O_114,N_14407,N_14596);
nor UO_115 (O_115,N_14277,N_14024);
or UO_116 (O_116,N_13874,N_13664);
and UO_117 (O_117,N_13946,N_14069);
nor UO_118 (O_118,N_14647,N_14589);
xor UO_119 (O_119,N_14515,N_14344);
and UO_120 (O_120,N_14357,N_13872);
nand UO_121 (O_121,N_13888,N_14846);
nand UO_122 (O_122,N_13848,N_14565);
or UO_123 (O_123,N_13967,N_14527);
nand UO_124 (O_124,N_14446,N_14873);
nand UO_125 (O_125,N_13516,N_14825);
nor UO_126 (O_126,N_13852,N_13726);
nor UO_127 (O_127,N_14427,N_14553);
and UO_128 (O_128,N_14386,N_14965);
nor UO_129 (O_129,N_13749,N_13898);
or UO_130 (O_130,N_13699,N_14103);
or UO_131 (O_131,N_13743,N_14902);
or UO_132 (O_132,N_14986,N_13620);
and UO_133 (O_133,N_14741,N_14646);
nand UO_134 (O_134,N_14739,N_13788);
and UO_135 (O_135,N_13508,N_14640);
or UO_136 (O_136,N_14860,N_14712);
nor UO_137 (O_137,N_13540,N_13932);
or UO_138 (O_138,N_13588,N_14900);
xor UO_139 (O_139,N_14236,N_14476);
nor UO_140 (O_140,N_13538,N_13563);
nand UO_141 (O_141,N_13529,N_14776);
xnor UO_142 (O_142,N_14950,N_13995);
or UO_143 (O_143,N_14359,N_14421);
xor UO_144 (O_144,N_14021,N_13789);
and UO_145 (O_145,N_13910,N_14856);
xnor UO_146 (O_146,N_14599,N_14402);
or UO_147 (O_147,N_14279,N_14310);
or UO_148 (O_148,N_14738,N_14283);
nor UO_149 (O_149,N_13793,N_14108);
nand UO_150 (O_150,N_14128,N_14056);
xnor UO_151 (O_151,N_13969,N_14289);
xor UO_152 (O_152,N_14823,N_13761);
nor UO_153 (O_153,N_14350,N_14227);
or UO_154 (O_154,N_14705,N_14802);
or UO_155 (O_155,N_13800,N_13635);
nand UO_156 (O_156,N_14704,N_14872);
and UO_157 (O_157,N_13895,N_14272);
or UO_158 (O_158,N_14858,N_14765);
or UO_159 (O_159,N_14813,N_13621);
or UO_160 (O_160,N_14367,N_14989);
nand UO_161 (O_161,N_14188,N_14798);
nand UO_162 (O_162,N_14093,N_13865);
nor UO_163 (O_163,N_14100,N_14506);
nor UO_164 (O_164,N_14173,N_14581);
xor UO_165 (O_165,N_14066,N_13669);
nand UO_166 (O_166,N_14249,N_13837);
nand UO_167 (O_167,N_14883,N_13845);
nand UO_168 (O_168,N_13721,N_14297);
and UO_169 (O_169,N_14462,N_14752);
nor UO_170 (O_170,N_13577,N_13510);
xor UO_171 (O_171,N_14408,N_14011);
xor UO_172 (O_172,N_14709,N_14162);
nand UO_173 (O_173,N_14974,N_14013);
and UO_174 (O_174,N_14891,N_13633);
xor UO_175 (O_175,N_14356,N_13527);
nand UO_176 (O_176,N_13679,N_13990);
nand UO_177 (O_177,N_14405,N_13740);
nor UO_178 (O_178,N_14217,N_14388);
nand UO_179 (O_179,N_13686,N_14723);
nand UO_180 (O_180,N_14040,N_13772);
nor UO_181 (O_181,N_14292,N_14085);
xor UO_182 (O_182,N_14719,N_14485);
nand UO_183 (O_183,N_14265,N_13964);
nand UO_184 (O_184,N_13545,N_13603);
and UO_185 (O_185,N_13598,N_14504);
nand UO_186 (O_186,N_14658,N_13576);
and UO_187 (O_187,N_14790,N_14821);
and UO_188 (O_188,N_13602,N_13752);
nand UO_189 (O_189,N_14092,N_14366);
nor UO_190 (O_190,N_14687,N_14973);
and UO_191 (O_191,N_14000,N_14735);
nor UO_192 (O_192,N_14195,N_14601);
nor UO_193 (O_193,N_14584,N_14539);
xnor UO_194 (O_194,N_13707,N_14497);
nor UO_195 (O_195,N_14513,N_14266);
and UO_196 (O_196,N_13911,N_14165);
and UO_197 (O_197,N_13913,N_14302);
nor UO_198 (O_198,N_14483,N_14233);
and UO_199 (O_199,N_14720,N_14322);
or UO_200 (O_200,N_13774,N_14324);
xnor UO_201 (O_201,N_14111,N_14913);
nor UO_202 (O_202,N_14548,N_13870);
or UO_203 (O_203,N_13806,N_14618);
and UO_204 (O_204,N_14216,N_13511);
and UO_205 (O_205,N_14114,N_13853);
and UO_206 (O_206,N_13803,N_13962);
and UO_207 (O_207,N_13663,N_14438);
nand UO_208 (O_208,N_13712,N_13579);
xor UO_209 (O_209,N_14521,N_13892);
nor UO_210 (O_210,N_13826,N_14892);
or UO_211 (O_211,N_13766,N_13668);
or UO_212 (O_212,N_14413,N_14378);
nor UO_213 (O_213,N_14098,N_13625);
xnor UO_214 (O_214,N_14509,N_14210);
and UO_215 (O_215,N_14577,N_13769);
or UO_216 (O_216,N_14360,N_14980);
nor UO_217 (O_217,N_13930,N_14078);
or UO_218 (O_218,N_14171,N_14831);
and UO_219 (O_219,N_14574,N_14583);
or UO_220 (O_220,N_14706,N_14512);
nor UO_221 (O_221,N_13856,N_13981);
nor UO_222 (O_222,N_14482,N_14001);
nand UO_223 (O_223,N_14670,N_14562);
nand UO_224 (O_224,N_14084,N_14186);
nor UO_225 (O_225,N_13864,N_14248);
xor UO_226 (O_226,N_14436,N_14460);
xor UO_227 (O_227,N_14775,N_13936);
xnor UO_228 (O_228,N_14144,N_14043);
nand UO_229 (O_229,N_13512,N_14118);
or UO_230 (O_230,N_14044,N_14404);
xor UO_231 (O_231,N_14432,N_14120);
and UO_232 (O_232,N_14061,N_14760);
and UO_233 (O_233,N_14999,N_14839);
or UO_234 (O_234,N_14071,N_14192);
or UO_235 (O_235,N_14886,N_14443);
xnor UO_236 (O_236,N_13777,N_13506);
or UO_237 (O_237,N_14113,N_14555);
and UO_238 (O_238,N_14153,N_14073);
nand UO_239 (O_239,N_14717,N_13671);
xor UO_240 (O_240,N_14771,N_14495);
nand UO_241 (O_241,N_14933,N_14552);
nor UO_242 (O_242,N_13939,N_14897);
and UO_243 (O_243,N_13807,N_14083);
xnor UO_244 (O_244,N_14035,N_13797);
nor UO_245 (O_245,N_14150,N_14631);
and UO_246 (O_246,N_14678,N_14142);
and UO_247 (O_247,N_13569,N_13927);
and UO_248 (O_248,N_14156,N_13654);
nand UO_249 (O_249,N_14146,N_14780);
nor UO_250 (O_250,N_13659,N_14988);
nand UO_251 (O_251,N_13578,N_14323);
or UO_252 (O_252,N_13836,N_13976);
nand UO_253 (O_253,N_13980,N_13878);
nor UO_254 (O_254,N_14025,N_14105);
and UO_255 (O_255,N_13961,N_13725);
and UO_256 (O_256,N_13891,N_13942);
nand UO_257 (O_257,N_13732,N_14370);
xor UO_258 (O_258,N_13798,N_14077);
or UO_259 (O_259,N_14203,N_13727);
and UO_260 (O_260,N_13907,N_13677);
nand UO_261 (O_261,N_14528,N_14546);
nor UO_262 (O_262,N_14914,N_14258);
nand UO_263 (O_263,N_13617,N_13688);
or UO_264 (O_264,N_14907,N_13716);
xor UO_265 (O_265,N_14511,N_14840);
xnor UO_266 (O_266,N_14617,N_14742);
and UO_267 (O_267,N_13770,N_13839);
nand UO_268 (O_268,N_13887,N_14273);
or UO_269 (O_269,N_14941,N_14567);
nor UO_270 (O_270,N_13994,N_14690);
and UO_271 (O_271,N_14576,N_14910);
or UO_272 (O_272,N_14795,N_13912);
xnor UO_273 (O_273,N_14536,N_14923);
nor UO_274 (O_274,N_14041,N_13672);
xnor UO_275 (O_275,N_13702,N_14863);
and UO_276 (O_276,N_14101,N_14976);
and UO_277 (O_277,N_14491,N_14486);
or UO_278 (O_278,N_14140,N_14389);
xnor UO_279 (O_279,N_13885,N_14267);
xor UO_280 (O_280,N_14956,N_14983);
or UO_281 (O_281,N_13568,N_14757);
nand UO_282 (O_282,N_13627,N_14761);
and UO_283 (O_283,N_14473,N_14667);
or UO_284 (O_284,N_13520,N_14196);
nor UO_285 (O_285,N_13794,N_14607);
and UO_286 (O_286,N_14303,N_14559);
or UO_287 (O_287,N_13673,N_14906);
or UO_288 (O_288,N_13670,N_14317);
xor UO_289 (O_289,N_14990,N_13722);
or UO_290 (O_290,N_14619,N_14147);
or UO_291 (O_291,N_14434,N_14335);
and UO_292 (O_292,N_14047,N_13824);
or UO_293 (O_293,N_13862,N_14855);
or UO_294 (O_294,N_14492,N_14580);
and UO_295 (O_295,N_13830,N_14107);
xor UO_296 (O_296,N_14901,N_14866);
xor UO_297 (O_297,N_14268,N_14057);
nor UO_298 (O_298,N_13996,N_14545);
nand UO_299 (O_299,N_14411,N_13984);
and UO_300 (O_300,N_13703,N_14137);
nor UO_301 (O_301,N_13801,N_14049);
or UO_302 (O_302,N_13534,N_13586);
xor UO_303 (O_303,N_14759,N_13678);
and UO_304 (O_304,N_14072,N_14478);
or UO_305 (O_305,N_14808,N_13823);
nor UO_306 (O_306,N_14600,N_14627);
or UO_307 (O_307,N_14365,N_14744);
nand UO_308 (O_308,N_14055,N_14372);
and UO_309 (O_309,N_14966,N_14593);
xnor UO_310 (O_310,N_14178,N_14161);
and UO_311 (O_311,N_14288,N_14703);
or UO_312 (O_312,N_13600,N_14648);
or UO_313 (O_313,N_14656,N_13813);
nor UO_314 (O_314,N_13735,N_14895);
or UO_315 (O_315,N_14613,N_14070);
and UO_316 (O_316,N_14911,N_14929);
or UO_317 (O_317,N_14348,N_14332);
and UO_318 (O_318,N_13708,N_14721);
xnor UO_319 (O_319,N_13675,N_14384);
xnor UO_320 (O_320,N_14624,N_13661);
nor UO_321 (O_321,N_13645,N_13763);
xnor UO_322 (O_322,N_14927,N_13811);
and UO_323 (O_323,N_14729,N_13841);
xor UO_324 (O_324,N_14014,N_14031);
and UO_325 (O_325,N_14163,N_14250);
and UO_326 (O_326,N_14822,N_13715);
nand UO_327 (O_327,N_14020,N_14397);
xnor UO_328 (O_328,N_14076,N_14889);
xor UO_329 (O_329,N_13503,N_14769);
or UO_330 (O_330,N_14159,N_14804);
nand UO_331 (O_331,N_14787,N_14968);
nor UO_332 (O_332,N_14916,N_14637);
nand UO_333 (O_333,N_13759,N_13623);
or UO_334 (O_334,N_13779,N_14884);
nor UO_335 (O_335,N_13851,N_14796);
or UO_336 (O_336,N_14836,N_14810);
nand UO_337 (O_337,N_14121,N_14228);
xnor UO_338 (O_338,N_13737,N_14595);
nand UO_339 (O_339,N_14507,N_13867);
or UO_340 (O_340,N_13631,N_14645);
xnor UO_341 (O_341,N_14374,N_14168);
xnor UO_342 (O_342,N_14587,N_13982);
and UO_343 (O_343,N_14204,N_14665);
nand UO_344 (O_344,N_13745,N_14758);
nor UO_345 (O_345,N_13795,N_13714);
or UO_346 (O_346,N_13653,N_14942);
nor UO_347 (O_347,N_13551,N_14737);
and UO_348 (O_348,N_14036,N_14343);
nor UO_349 (O_349,N_13731,N_13698);
nor UO_350 (O_350,N_14949,N_14109);
or UO_351 (O_351,N_14112,N_14447);
xnor UO_352 (O_352,N_14394,N_14791);
nand UO_353 (O_353,N_14848,N_14026);
and UO_354 (O_354,N_13765,N_13989);
or UO_355 (O_355,N_14959,N_14992);
nor UO_356 (O_356,N_13691,N_13815);
or UO_357 (O_357,N_14116,N_13683);
nor UO_358 (O_358,N_14028,N_13889);
nand UO_359 (O_359,N_13816,N_14242);
xnor UO_360 (O_360,N_13616,N_14239);
xnor UO_361 (O_361,N_14751,N_13728);
or UO_362 (O_362,N_14193,N_13700);
nor UO_363 (O_363,N_14978,N_14245);
and UO_364 (O_364,N_14423,N_13941);
nor UO_365 (O_365,N_14557,N_14060);
and UO_366 (O_366,N_14685,N_13519);
xnor UO_367 (O_367,N_14532,N_14642);
or UO_368 (O_368,N_14675,N_14925);
and UO_369 (O_369,N_14176,N_14650);
and UO_370 (O_370,N_13730,N_14459);
xor UO_371 (O_371,N_13724,N_14206);
and UO_372 (O_372,N_14213,N_14936);
or UO_373 (O_373,N_13787,N_14448);
and UO_374 (O_374,N_14611,N_13778);
nand UO_375 (O_375,N_14952,N_13681);
and UO_376 (O_376,N_14033,N_14605);
nor UO_377 (O_377,N_14960,N_14298);
and UO_378 (O_378,N_14696,N_13914);
xnor UO_379 (O_379,N_13719,N_14255);
nand UO_380 (O_380,N_14591,N_13917);
nand UO_381 (O_381,N_14797,N_14805);
nor UO_382 (O_382,N_14286,N_14305);
xor UO_383 (O_383,N_13697,N_13952);
nor UO_384 (O_384,N_14032,N_13883);
and UO_385 (O_385,N_13701,N_13612);
nand UO_386 (O_386,N_13524,N_13918);
xnor UO_387 (O_387,N_14371,N_13750);
xor UO_388 (O_388,N_14948,N_14425);
or UO_389 (O_389,N_13979,N_13585);
xor UO_390 (O_390,N_14309,N_13709);
or UO_391 (O_391,N_14353,N_13608);
nand UO_392 (O_392,N_14320,N_14668);
nor UO_393 (O_393,N_14127,N_14004);
and UO_394 (O_394,N_14003,N_14082);
and UO_395 (O_395,N_14200,N_14030);
xnor UO_396 (O_396,N_14006,N_14488);
and UO_397 (O_397,N_13515,N_14569);
nand UO_398 (O_398,N_13667,N_13718);
xnor UO_399 (O_399,N_14746,N_14050);
nor UO_400 (O_400,N_14590,N_13756);
and UO_401 (O_401,N_14938,N_14158);
nor UO_402 (O_402,N_14749,N_14623);
xnor UO_403 (O_403,N_13869,N_13630);
and UO_404 (O_404,N_14606,N_14682);
nand UO_405 (O_405,N_13921,N_14149);
or UO_406 (O_406,N_13764,N_14409);
xor UO_407 (O_407,N_14334,N_14867);
nor UO_408 (O_408,N_13550,N_13786);
or UO_409 (O_409,N_14625,N_13838);
nand UO_410 (O_410,N_14890,N_14674);
nand UO_411 (O_411,N_14449,N_14899);
nand UO_412 (O_412,N_14887,N_14905);
and UO_413 (O_413,N_14219,N_13890);
nor UO_414 (O_414,N_13920,N_14480);
xnor UO_415 (O_415,N_14772,N_14519);
nand UO_416 (O_416,N_13968,N_13855);
and UO_417 (O_417,N_14274,N_14909);
or UO_418 (O_418,N_13849,N_14920);
and UO_419 (O_419,N_14947,N_14754);
xor UO_420 (O_420,N_14541,N_13662);
or UO_421 (O_421,N_14336,N_13581);
and UO_422 (O_422,N_13583,N_14412);
and UO_423 (O_423,N_14740,N_14733);
nor UO_424 (O_424,N_14745,N_14556);
or UO_425 (O_425,N_14629,N_13881);
xnor UO_426 (O_426,N_13782,N_13947);
or UO_427 (O_427,N_14770,N_14669);
or UO_428 (O_428,N_14870,N_14898);
nor UO_429 (O_429,N_14995,N_14016);
nor UO_430 (O_430,N_13641,N_13760);
xnor UO_431 (O_431,N_13513,N_13957);
nand UO_432 (O_432,N_13544,N_14816);
nor UO_433 (O_433,N_14766,N_14445);
nand UO_434 (O_434,N_14523,N_13685);
or UO_435 (O_435,N_13666,N_14183);
and UO_436 (O_436,N_13501,N_13558);
nand UO_437 (O_437,N_14202,N_14089);
or UO_438 (O_438,N_14293,N_13742);
or UO_439 (O_439,N_14275,N_14630);
nor UO_440 (O_440,N_14908,N_13850);
and UO_441 (O_441,N_13565,N_14534);
nand UO_442 (O_442,N_14930,N_14628);
nand UO_443 (O_443,N_14005,N_14661);
nand UO_444 (O_444,N_13747,N_14243);
xor UO_445 (O_445,N_14380,N_14037);
xnor UO_446 (O_446,N_14131,N_14540);
and UO_447 (O_447,N_13814,N_14845);
nor UO_448 (O_448,N_14134,N_14352);
nand UO_449 (O_449,N_14928,N_14466);
nand UO_450 (O_450,N_13829,N_13999);
and UO_451 (O_451,N_14379,N_14807);
nor UO_452 (O_452,N_14396,N_14110);
xnor UO_453 (O_453,N_14919,N_13933);
nand UO_454 (O_454,N_14833,N_13860);
or UO_455 (O_455,N_13656,N_13648);
nor UO_456 (O_456,N_14383,N_14487);
nand UO_457 (O_457,N_14672,N_14710);
and UO_458 (O_458,N_14319,N_14525);
xnor UO_459 (O_459,N_14981,N_14641);
or UO_460 (O_460,N_14558,N_14885);
nand UO_461 (O_461,N_14375,N_14785);
xor UO_462 (O_462,N_14199,N_14263);
and UO_463 (O_463,N_13553,N_14655);
nand UO_464 (O_464,N_14997,N_14803);
nand UO_465 (O_465,N_14074,N_14835);
and UO_466 (O_466,N_13704,N_14094);
nand UO_467 (O_467,N_14713,N_13537);
nor UO_468 (O_468,N_13827,N_14223);
nor UO_469 (O_469,N_14081,N_14854);
nand UO_470 (O_470,N_14417,N_14442);
xor UO_471 (O_471,N_14699,N_14994);
and UO_472 (O_472,N_14437,N_14180);
or UO_473 (O_473,N_14062,N_13991);
xnor UO_474 (O_474,N_14849,N_13820);
and UO_475 (O_475,N_14240,N_14817);
nor UO_476 (O_476,N_13723,N_13953);
nand UO_477 (O_477,N_13945,N_13833);
or UO_478 (O_478,N_13899,N_14464);
nor UO_479 (O_479,N_14964,N_13871);
nor UO_480 (O_480,N_14922,N_13596);
and UO_481 (O_481,N_13861,N_13736);
nand UO_482 (O_482,N_13940,N_14174);
and UO_483 (O_483,N_14657,N_14194);
xnor UO_484 (O_484,N_13532,N_13835);
and UO_485 (O_485,N_14979,N_14054);
nor UO_486 (O_486,N_14602,N_13916);
and UO_487 (O_487,N_14294,N_14145);
xnor UO_488 (O_488,N_14201,N_13567);
and UO_489 (O_489,N_13638,N_13859);
or UO_490 (O_490,N_14419,N_14788);
nor UO_491 (O_491,N_14123,N_14903);
and UO_492 (O_492,N_13528,N_13802);
nand UO_493 (O_493,N_13658,N_13636);
xor UO_494 (O_494,N_14007,N_13705);
nand UO_495 (O_495,N_14862,N_14824);
nor UO_496 (O_496,N_13963,N_14363);
or UO_497 (O_497,N_14526,N_14315);
nand UO_498 (O_498,N_14578,N_14970);
or UO_499 (O_499,N_14251,N_14226);
and UO_500 (O_500,N_14038,N_13680);
or UO_501 (O_501,N_14235,N_13909);
or UO_502 (O_502,N_14571,N_14794);
nand UO_503 (O_503,N_14560,N_14747);
and UO_504 (O_504,N_14842,N_14819);
or UO_505 (O_505,N_14017,N_14736);
and UO_506 (O_506,N_14764,N_14398);
xnor UO_507 (O_507,N_14470,N_14337);
or UO_508 (O_508,N_14015,N_14088);
nand UO_509 (O_509,N_14373,N_14779);
and UO_510 (O_510,N_13767,N_14326);
and UO_511 (O_511,N_13817,N_13796);
nor UO_512 (O_512,N_13893,N_14452);
and UO_513 (O_513,N_13846,N_13647);
nand UO_514 (O_514,N_14888,N_14355);
or UO_515 (O_515,N_13985,N_14946);
nor UO_516 (O_516,N_13655,N_14939);
and UO_517 (O_517,N_13554,N_14185);
xnor UO_518 (O_518,N_13938,N_14237);
nor UO_519 (O_519,N_14136,N_13809);
nand UO_520 (O_520,N_14530,N_14333);
and UO_521 (O_521,N_13572,N_14877);
or UO_522 (O_522,N_13857,N_14649);
or UO_523 (O_523,N_14851,N_14784);
and UO_524 (O_524,N_13552,N_13956);
xnor UO_525 (O_525,N_13751,N_14461);
xnor UO_526 (O_526,N_14207,N_14368);
or UO_527 (O_527,N_14212,N_13729);
nor UO_528 (O_528,N_14568,N_14086);
nor UO_529 (O_529,N_13626,N_14209);
xnor UO_530 (O_530,N_14850,N_14457);
xnor UO_531 (O_531,N_13819,N_14573);
and UO_532 (O_532,N_14904,N_14542);
nor UO_533 (O_533,N_14291,N_13970);
or UO_534 (O_534,N_14285,N_14786);
or UO_535 (O_535,N_13618,N_14278);
or UO_536 (O_536,N_13858,N_13593);
xnor UO_537 (O_537,N_14852,N_13843);
nand UO_538 (O_538,N_13755,N_14707);
nand UO_539 (O_539,N_14489,N_14401);
and UO_540 (O_540,N_14815,N_14944);
or UO_541 (O_541,N_14130,N_14533);
and UO_542 (O_542,N_13547,N_13971);
and UO_543 (O_543,N_13790,N_14099);
nand UO_544 (O_544,N_14516,N_14097);
xnor UO_545 (O_545,N_14594,N_14869);
or UO_546 (O_546,N_13525,N_14975);
nor UO_547 (O_547,N_13882,N_14126);
or UO_548 (O_548,N_13556,N_14215);
xor UO_549 (O_549,N_13925,N_14340);
nand UO_550 (O_550,N_14688,N_13665);
xnor UO_551 (O_551,N_14882,N_13902);
or UO_552 (O_552,N_14187,N_13582);
nor UO_553 (O_553,N_14915,N_13504);
nand UO_554 (O_554,N_14912,N_14958);
and UO_555 (O_555,N_14762,N_13682);
or UO_556 (O_556,N_14431,N_14316);
nor UO_557 (O_557,N_14957,N_14827);
and UO_558 (O_558,N_14689,N_14598);
and UO_559 (O_559,N_13639,N_14505);
nor UO_560 (O_560,N_14874,N_13847);
and UO_561 (O_561,N_14564,N_14880);
xor UO_562 (O_562,N_14653,N_14208);
nand UO_563 (O_563,N_13960,N_13660);
and UO_564 (O_564,N_14018,N_14878);
xor UO_565 (O_565,N_14406,N_14471);
nor UO_566 (O_566,N_14259,N_13739);
nor UO_567 (O_567,N_14755,N_14189);
nand UO_568 (O_568,N_13517,N_14838);
xnor UO_569 (O_569,N_13744,N_14644);
or UO_570 (O_570,N_14472,N_14416);
nor UO_571 (O_571,N_14244,N_14768);
nand UO_572 (O_572,N_14290,N_14894);
or UO_573 (O_573,N_14231,N_14179);
or UO_574 (O_574,N_14998,N_14799);
and UO_575 (O_575,N_14148,N_14566);
and UO_576 (O_576,N_14022,N_13863);
nand UO_577 (O_577,N_14064,N_14172);
nand UO_578 (O_578,N_14830,N_14544);
nand UO_579 (O_579,N_14296,N_13748);
xor UO_580 (O_580,N_14052,N_14924);
xor UO_581 (O_581,N_14058,N_13834);
xor UO_582 (O_582,N_14684,N_14023);
and UO_583 (O_583,N_13904,N_14392);
and UO_584 (O_584,N_14861,N_14330);
and UO_585 (O_585,N_14221,N_14588);
nor UO_586 (O_586,N_14338,N_13840);
or UO_587 (O_587,N_14498,N_14454);
and UO_588 (O_588,N_14117,N_14679);
and UO_589 (O_589,N_14800,N_14395);
nor UO_590 (O_590,N_14954,N_14253);
nor UO_591 (O_591,N_14385,N_14256);
xnor UO_592 (O_592,N_13825,N_14102);
nand UO_593 (O_593,N_13768,N_13958);
nand UO_594 (O_594,N_14643,N_13988);
nor UO_595 (O_595,N_14774,N_13690);
nand UO_596 (O_596,N_14563,N_13822);
nor UO_597 (O_597,N_14422,N_13757);
and UO_598 (O_598,N_14247,N_14262);
nand UO_599 (O_599,N_14400,N_14420);
or UO_600 (O_600,N_13738,N_14458);
nand UO_601 (O_601,N_13746,N_14477);
or UO_602 (O_602,N_13650,N_14479);
xnor UO_603 (O_603,N_14175,N_13589);
nand UO_604 (O_604,N_14937,N_13901);
xor UO_605 (O_605,N_14812,N_13937);
nand UO_606 (O_606,N_14218,N_13502);
nor UO_607 (O_607,N_14681,N_14575);
or UO_608 (O_608,N_13676,N_13754);
and UO_609 (O_609,N_14859,N_14191);
xor UO_610 (O_610,N_13949,N_14972);
nand UO_611 (O_611,N_14155,N_13687);
xnor UO_612 (O_612,N_14481,N_14834);
nor UO_613 (O_613,N_14465,N_13587);
xnor UO_614 (O_614,N_13818,N_14468);
or UO_615 (O_615,N_13832,N_14182);
xnor UO_616 (O_616,N_14341,N_14439);
nand UO_617 (O_617,N_14695,N_13693);
and UO_618 (O_618,N_13924,N_14493);
nand UO_619 (O_619,N_14135,N_14701);
or UO_620 (O_620,N_14832,N_14496);
xor UO_621 (O_621,N_14789,N_13652);
xor UO_622 (O_622,N_14971,N_13879);
and UO_623 (O_623,N_14750,N_13908);
nor UO_624 (O_624,N_13784,N_13771);
nand UO_625 (O_625,N_14214,N_14387);
and UO_626 (O_626,N_14529,N_14129);
xor UO_627 (O_627,N_14666,N_13710);
xnor UO_628 (O_628,N_14635,N_14692);
nand UO_629 (O_629,N_13523,N_13972);
or UO_630 (O_630,N_14714,N_14693);
nand UO_631 (O_631,N_14433,N_14059);
or UO_632 (O_632,N_14230,N_14826);
nor UO_633 (O_633,N_13514,N_13905);
nor UO_634 (O_634,N_14429,N_13897);
nor UO_635 (O_635,N_14510,N_13828);
xnor UO_636 (O_636,N_14132,N_14300);
nor UO_637 (O_637,N_14697,N_13854);
nand UO_638 (O_638,N_14312,N_14414);
xor UO_639 (O_639,N_14782,N_14205);
nor UO_640 (O_640,N_13584,N_13696);
and UO_641 (O_641,N_14953,N_14170);
nand UO_642 (O_642,N_13929,N_14087);
nor UO_643 (O_643,N_14246,N_14328);
and UO_644 (O_644,N_14106,N_14543);
xor UO_645 (O_645,N_14284,N_13876);
nand UO_646 (O_646,N_13844,N_13634);
nand UO_647 (O_647,N_14730,N_13622);
or UO_648 (O_648,N_13792,N_14276);
or UO_649 (O_649,N_13948,N_14608);
nor UO_650 (O_650,N_14524,N_14783);
xor UO_651 (O_651,N_13812,N_14048);
and UO_652 (O_652,N_14444,N_14295);
nand UO_653 (O_653,N_14382,N_14391);
or UO_654 (O_654,N_14426,N_13521);
nor UO_655 (O_655,N_13574,N_13711);
and UO_656 (O_656,N_13561,N_14181);
and UO_657 (O_657,N_14639,N_14430);
xnor UO_658 (O_658,N_14844,N_14377);
nor UO_659 (O_659,N_13560,N_14550);
nand UO_660 (O_660,N_14095,N_14663);
or UO_661 (O_661,N_14702,N_14763);
and UO_662 (O_662,N_14868,N_14490);
or UO_663 (O_663,N_13518,N_14029);
and UO_664 (O_664,N_13805,N_14691);
nand UO_665 (O_665,N_13873,N_13966);
or UO_666 (O_666,N_14224,N_14753);
or UO_667 (O_667,N_13566,N_13615);
xor UO_668 (O_668,N_14820,N_14811);
nor UO_669 (O_669,N_14381,N_14651);
xnor UO_670 (O_670,N_13720,N_14361);
and UO_671 (O_671,N_14184,N_13733);
xor UO_672 (O_672,N_14961,N_13684);
xor UO_673 (O_673,N_14814,N_14865);
nor UO_674 (O_674,N_13975,N_14264);
nand UO_675 (O_675,N_14010,N_13500);
nor UO_676 (O_676,N_14301,N_13886);
nand UO_677 (O_677,N_14167,N_14982);
and UO_678 (O_678,N_14547,N_14715);
xnor UO_679 (O_679,N_13877,N_14514);
xor UO_680 (O_680,N_14963,N_14143);
and UO_681 (O_681,N_14351,N_13592);
and UO_682 (O_682,N_13896,N_14306);
or UO_683 (O_683,N_14572,N_14369);
nand UO_684 (O_684,N_14743,N_14281);
or UO_685 (O_685,N_14154,N_13541);
nor UO_686 (O_686,N_14428,N_13651);
nor UO_687 (O_687,N_13926,N_13931);
and UO_688 (O_688,N_14053,N_14664);
nor UO_689 (O_689,N_13780,N_14597);
nand UO_690 (O_690,N_13580,N_13571);
and UO_691 (O_691,N_14932,N_14475);
and UO_692 (O_692,N_14921,N_14700);
or UO_693 (O_693,N_13781,N_14809);
nor UO_694 (O_694,N_14731,N_14969);
nor UO_695 (O_695,N_13894,N_14234);
nor UO_696 (O_696,N_13808,N_14881);
nor UO_697 (O_697,N_14068,N_14945);
or UO_698 (O_698,N_14339,N_13900);
nand UO_699 (O_699,N_14917,N_14169);
or UO_700 (O_700,N_14311,N_14612);
and UO_701 (O_701,N_13993,N_14027);
nor UO_702 (O_702,N_14327,N_13950);
and UO_703 (O_703,N_13640,N_14615);
nand UO_704 (O_704,N_14801,N_13562);
and UO_705 (O_705,N_14828,N_14133);
nand UO_706 (O_706,N_14342,N_13998);
or UO_707 (O_707,N_14270,N_13597);
xnor UO_708 (O_708,N_14329,N_13607);
nand UO_709 (O_709,N_13548,N_14080);
or UO_710 (O_710,N_13831,N_14843);
or UO_711 (O_711,N_13785,N_13531);
nand UO_712 (O_712,N_14501,N_14220);
nor UO_713 (O_713,N_14724,N_13555);
nand UO_714 (O_714,N_14090,N_13974);
xor UO_715 (O_715,N_14502,N_14034);
xnor UO_716 (O_716,N_13965,N_14260);
nand UO_717 (O_717,N_14621,N_13986);
nand UO_718 (O_718,N_14636,N_14818);
or UO_719 (O_719,N_13977,N_13591);
xnor UO_720 (O_720,N_14727,N_14347);
or UO_721 (O_721,N_14570,N_14864);
or UO_722 (O_722,N_14549,N_14654);
or UO_723 (O_723,N_14418,N_13674);
or UO_724 (O_724,N_14538,N_14728);
xor UO_725 (O_725,N_14676,N_14009);
xor UO_726 (O_726,N_13943,N_14469);
and UO_727 (O_727,N_14551,N_14781);
nor UO_728 (O_728,N_14124,N_13601);
nand UO_729 (O_729,N_14152,N_14225);
xor UO_730 (O_730,N_14424,N_14045);
nand UO_731 (O_731,N_14269,N_13507);
nand UO_732 (O_732,N_14620,N_13536);
or UO_733 (O_733,N_14254,N_14346);
nand UO_734 (O_734,N_14474,N_14257);
nor UO_735 (O_735,N_14096,N_14582);
or UO_736 (O_736,N_13599,N_14138);
nor UO_737 (O_737,N_14756,N_14535);
nand UO_738 (O_738,N_13637,N_14160);
and UO_739 (O_739,N_14313,N_13934);
nor UO_740 (O_740,N_14777,N_14508);
or UO_741 (O_741,N_14019,N_14211);
nor UO_742 (O_742,N_14984,N_14065);
xnor UO_743 (O_743,N_13959,N_13694);
xor UO_744 (O_744,N_14157,N_13614);
nand UO_745 (O_745,N_14520,N_14331);
nand UO_746 (O_746,N_14141,N_14622);
and UO_747 (O_747,N_14659,N_14115);
or UO_748 (O_748,N_13613,N_13734);
and UO_749 (O_749,N_14686,N_13522);
or UO_750 (O_750,N_13997,N_14818);
nor UO_751 (O_751,N_14480,N_14160);
xnor UO_752 (O_752,N_14454,N_14319);
or UO_753 (O_753,N_14990,N_14657);
xor UO_754 (O_754,N_14123,N_13746);
nor UO_755 (O_755,N_14115,N_14441);
nor UO_756 (O_756,N_14027,N_13947);
nand UO_757 (O_757,N_13616,N_14491);
nor UO_758 (O_758,N_14929,N_14172);
and UO_759 (O_759,N_14999,N_14368);
xor UO_760 (O_760,N_13870,N_14150);
nand UO_761 (O_761,N_13773,N_14751);
xor UO_762 (O_762,N_14406,N_14540);
xor UO_763 (O_763,N_14521,N_13869);
nor UO_764 (O_764,N_14784,N_14882);
nand UO_765 (O_765,N_14337,N_14019);
and UO_766 (O_766,N_14996,N_14294);
or UO_767 (O_767,N_13549,N_14280);
or UO_768 (O_768,N_14534,N_14377);
nand UO_769 (O_769,N_13999,N_14677);
and UO_770 (O_770,N_13923,N_14310);
nand UO_771 (O_771,N_14146,N_14510);
nor UO_772 (O_772,N_13674,N_14839);
nor UO_773 (O_773,N_14156,N_13689);
or UO_774 (O_774,N_13643,N_14526);
xnor UO_775 (O_775,N_13531,N_14384);
or UO_776 (O_776,N_14950,N_14872);
nor UO_777 (O_777,N_13855,N_14596);
nand UO_778 (O_778,N_13835,N_14849);
nor UO_779 (O_779,N_13598,N_13912);
nor UO_780 (O_780,N_14116,N_13657);
nand UO_781 (O_781,N_13552,N_13809);
xnor UO_782 (O_782,N_14960,N_14745);
nor UO_783 (O_783,N_14930,N_13819);
nand UO_784 (O_784,N_13650,N_14906);
or UO_785 (O_785,N_13767,N_13601);
nor UO_786 (O_786,N_14608,N_14008);
and UO_787 (O_787,N_14666,N_14824);
or UO_788 (O_788,N_13974,N_14145);
xor UO_789 (O_789,N_13954,N_13918);
nand UO_790 (O_790,N_13551,N_14788);
nor UO_791 (O_791,N_14273,N_14955);
xor UO_792 (O_792,N_13950,N_14415);
and UO_793 (O_793,N_14615,N_14684);
nor UO_794 (O_794,N_14557,N_13973);
xor UO_795 (O_795,N_14423,N_13921);
nor UO_796 (O_796,N_14134,N_13741);
xor UO_797 (O_797,N_14283,N_14232);
nor UO_798 (O_798,N_13757,N_14241);
nand UO_799 (O_799,N_13679,N_13883);
or UO_800 (O_800,N_13623,N_13986);
and UO_801 (O_801,N_14562,N_14317);
nand UO_802 (O_802,N_13745,N_13871);
xor UO_803 (O_803,N_13628,N_13963);
nor UO_804 (O_804,N_14534,N_13777);
nand UO_805 (O_805,N_13916,N_13671);
and UO_806 (O_806,N_14726,N_14350);
xnor UO_807 (O_807,N_13781,N_13527);
or UO_808 (O_808,N_14037,N_13760);
and UO_809 (O_809,N_14396,N_14378);
or UO_810 (O_810,N_14730,N_14784);
and UO_811 (O_811,N_14098,N_13812);
xnor UO_812 (O_812,N_14489,N_14956);
or UO_813 (O_813,N_14014,N_14371);
nand UO_814 (O_814,N_14153,N_13669);
and UO_815 (O_815,N_14683,N_14118);
or UO_816 (O_816,N_13857,N_14798);
or UO_817 (O_817,N_13975,N_13671);
xor UO_818 (O_818,N_14205,N_14653);
or UO_819 (O_819,N_14534,N_14337);
nand UO_820 (O_820,N_14236,N_13572);
nand UO_821 (O_821,N_13672,N_14146);
xnor UO_822 (O_822,N_14875,N_14716);
nor UO_823 (O_823,N_14324,N_13823);
nor UO_824 (O_824,N_14875,N_14735);
nor UO_825 (O_825,N_13916,N_13748);
nor UO_826 (O_826,N_14388,N_13671);
xor UO_827 (O_827,N_14156,N_14346);
nand UO_828 (O_828,N_13605,N_14728);
or UO_829 (O_829,N_13964,N_14187);
nor UO_830 (O_830,N_13693,N_13681);
nor UO_831 (O_831,N_14286,N_13635);
nand UO_832 (O_832,N_14353,N_14974);
nor UO_833 (O_833,N_14239,N_14774);
nor UO_834 (O_834,N_13733,N_14169);
xor UO_835 (O_835,N_14783,N_14032);
and UO_836 (O_836,N_14085,N_14673);
nor UO_837 (O_837,N_14310,N_14262);
nor UO_838 (O_838,N_13796,N_14807);
xor UO_839 (O_839,N_13918,N_14666);
and UO_840 (O_840,N_13724,N_14164);
xnor UO_841 (O_841,N_14049,N_13874);
nand UO_842 (O_842,N_14382,N_14562);
and UO_843 (O_843,N_13710,N_13688);
nor UO_844 (O_844,N_14852,N_14579);
or UO_845 (O_845,N_14072,N_14712);
xnor UO_846 (O_846,N_14501,N_14795);
or UO_847 (O_847,N_14643,N_14071);
nand UO_848 (O_848,N_13648,N_14776);
and UO_849 (O_849,N_14526,N_13894);
or UO_850 (O_850,N_14819,N_13512);
or UO_851 (O_851,N_13856,N_14720);
nand UO_852 (O_852,N_14397,N_13558);
nand UO_853 (O_853,N_14250,N_13766);
or UO_854 (O_854,N_14607,N_13565);
xnor UO_855 (O_855,N_14739,N_14787);
or UO_856 (O_856,N_14934,N_14107);
or UO_857 (O_857,N_14149,N_13754);
nand UO_858 (O_858,N_13898,N_14352);
or UO_859 (O_859,N_14029,N_14086);
or UO_860 (O_860,N_14028,N_14317);
nand UO_861 (O_861,N_13530,N_13982);
or UO_862 (O_862,N_14851,N_14925);
nand UO_863 (O_863,N_14129,N_13761);
and UO_864 (O_864,N_13754,N_13823);
and UO_865 (O_865,N_14522,N_14909);
and UO_866 (O_866,N_14668,N_13749);
nor UO_867 (O_867,N_14776,N_14454);
and UO_868 (O_868,N_14936,N_13821);
or UO_869 (O_869,N_14149,N_14289);
xnor UO_870 (O_870,N_13849,N_14528);
and UO_871 (O_871,N_14510,N_14093);
xnor UO_872 (O_872,N_13543,N_14753);
or UO_873 (O_873,N_14894,N_14985);
and UO_874 (O_874,N_14111,N_13835);
xor UO_875 (O_875,N_14025,N_14600);
nand UO_876 (O_876,N_14375,N_14967);
nor UO_877 (O_877,N_13992,N_13713);
nor UO_878 (O_878,N_13897,N_14742);
nand UO_879 (O_879,N_14249,N_13811);
nor UO_880 (O_880,N_14304,N_13610);
nand UO_881 (O_881,N_14308,N_13991);
or UO_882 (O_882,N_14088,N_13836);
or UO_883 (O_883,N_13563,N_14113);
nand UO_884 (O_884,N_13904,N_14808);
nor UO_885 (O_885,N_14752,N_14932);
and UO_886 (O_886,N_13732,N_14389);
nand UO_887 (O_887,N_14077,N_13612);
xor UO_888 (O_888,N_14354,N_14430);
or UO_889 (O_889,N_14103,N_14113);
nor UO_890 (O_890,N_13646,N_14838);
or UO_891 (O_891,N_14670,N_14633);
xnor UO_892 (O_892,N_14287,N_14956);
nand UO_893 (O_893,N_14704,N_13615);
and UO_894 (O_894,N_14963,N_14531);
and UO_895 (O_895,N_13928,N_13827);
nand UO_896 (O_896,N_14142,N_14730);
or UO_897 (O_897,N_13928,N_14529);
and UO_898 (O_898,N_13898,N_14760);
nand UO_899 (O_899,N_14939,N_14469);
or UO_900 (O_900,N_13555,N_14347);
xor UO_901 (O_901,N_13603,N_14526);
nor UO_902 (O_902,N_14882,N_13531);
xnor UO_903 (O_903,N_14758,N_14445);
xor UO_904 (O_904,N_14588,N_14240);
nand UO_905 (O_905,N_14887,N_13854);
nand UO_906 (O_906,N_14043,N_14129);
nor UO_907 (O_907,N_13734,N_13601);
nand UO_908 (O_908,N_14303,N_13894);
xnor UO_909 (O_909,N_13672,N_14069);
nand UO_910 (O_910,N_13674,N_14097);
nand UO_911 (O_911,N_14662,N_14468);
and UO_912 (O_912,N_13639,N_14278);
nand UO_913 (O_913,N_13766,N_13814);
nor UO_914 (O_914,N_13836,N_13591);
and UO_915 (O_915,N_14678,N_13530);
nor UO_916 (O_916,N_14675,N_14181);
xor UO_917 (O_917,N_14360,N_14391);
or UO_918 (O_918,N_14783,N_14618);
nor UO_919 (O_919,N_14660,N_13895);
or UO_920 (O_920,N_13919,N_13699);
or UO_921 (O_921,N_13814,N_13992);
xnor UO_922 (O_922,N_14535,N_14095);
nand UO_923 (O_923,N_14301,N_13803);
or UO_924 (O_924,N_13753,N_13880);
xnor UO_925 (O_925,N_14928,N_13803);
or UO_926 (O_926,N_13873,N_14470);
xor UO_927 (O_927,N_14304,N_13866);
or UO_928 (O_928,N_13580,N_13863);
or UO_929 (O_929,N_14621,N_14187);
and UO_930 (O_930,N_13655,N_14492);
xor UO_931 (O_931,N_14299,N_13981);
and UO_932 (O_932,N_14108,N_14952);
nand UO_933 (O_933,N_14400,N_13773);
xor UO_934 (O_934,N_14370,N_13807);
nor UO_935 (O_935,N_13617,N_14573);
and UO_936 (O_936,N_13660,N_14102);
xnor UO_937 (O_937,N_13703,N_13665);
and UO_938 (O_938,N_14956,N_14628);
nor UO_939 (O_939,N_14076,N_14758);
and UO_940 (O_940,N_14408,N_14001);
and UO_941 (O_941,N_14527,N_14764);
xnor UO_942 (O_942,N_14248,N_14464);
xnor UO_943 (O_943,N_14598,N_14766);
nand UO_944 (O_944,N_13680,N_14757);
xnor UO_945 (O_945,N_13575,N_13878);
nand UO_946 (O_946,N_13664,N_13881);
xnor UO_947 (O_947,N_14827,N_14738);
and UO_948 (O_948,N_14042,N_13911);
nor UO_949 (O_949,N_14152,N_14086);
and UO_950 (O_950,N_14224,N_14263);
xor UO_951 (O_951,N_14689,N_14063);
nor UO_952 (O_952,N_14919,N_14967);
nor UO_953 (O_953,N_14502,N_13870);
and UO_954 (O_954,N_13577,N_14625);
xor UO_955 (O_955,N_14094,N_14121);
nor UO_956 (O_956,N_14949,N_14955);
and UO_957 (O_957,N_14712,N_13521);
nor UO_958 (O_958,N_14973,N_14191);
nand UO_959 (O_959,N_14166,N_14176);
or UO_960 (O_960,N_13720,N_14324);
nor UO_961 (O_961,N_14081,N_14272);
and UO_962 (O_962,N_14473,N_14406);
nand UO_963 (O_963,N_14058,N_14812);
xor UO_964 (O_964,N_13541,N_14122);
and UO_965 (O_965,N_14592,N_14113);
nand UO_966 (O_966,N_13509,N_14046);
and UO_967 (O_967,N_14229,N_13785);
or UO_968 (O_968,N_13678,N_14442);
nor UO_969 (O_969,N_13994,N_14886);
and UO_970 (O_970,N_13675,N_13538);
or UO_971 (O_971,N_14163,N_13919);
nor UO_972 (O_972,N_14333,N_13900);
and UO_973 (O_973,N_14639,N_14774);
and UO_974 (O_974,N_13627,N_14283);
and UO_975 (O_975,N_14952,N_14799);
or UO_976 (O_976,N_13596,N_13909);
nor UO_977 (O_977,N_14869,N_14994);
nand UO_978 (O_978,N_14372,N_13689);
and UO_979 (O_979,N_14765,N_14178);
or UO_980 (O_980,N_13924,N_14754);
and UO_981 (O_981,N_14059,N_13590);
xor UO_982 (O_982,N_13701,N_14383);
nand UO_983 (O_983,N_14438,N_14319);
or UO_984 (O_984,N_14123,N_14800);
or UO_985 (O_985,N_13668,N_14575);
nand UO_986 (O_986,N_13765,N_14010);
nor UO_987 (O_987,N_14730,N_14965);
nand UO_988 (O_988,N_14113,N_13600);
and UO_989 (O_989,N_14079,N_14264);
xnor UO_990 (O_990,N_13625,N_14767);
or UO_991 (O_991,N_13985,N_13576);
nand UO_992 (O_992,N_14627,N_13659);
and UO_993 (O_993,N_14074,N_14987);
and UO_994 (O_994,N_14214,N_14198);
nor UO_995 (O_995,N_14538,N_14611);
and UO_996 (O_996,N_14510,N_14032);
or UO_997 (O_997,N_14746,N_14382);
xnor UO_998 (O_998,N_14320,N_13899);
and UO_999 (O_999,N_13667,N_14671);
or UO_1000 (O_1000,N_14415,N_14452);
nor UO_1001 (O_1001,N_14348,N_13755);
nor UO_1002 (O_1002,N_14300,N_14887);
or UO_1003 (O_1003,N_13956,N_13547);
nor UO_1004 (O_1004,N_14404,N_13504);
nor UO_1005 (O_1005,N_14350,N_13800);
xnor UO_1006 (O_1006,N_14753,N_13500);
xor UO_1007 (O_1007,N_14076,N_13532);
or UO_1008 (O_1008,N_14390,N_14698);
and UO_1009 (O_1009,N_14857,N_14093);
or UO_1010 (O_1010,N_14016,N_13717);
xnor UO_1011 (O_1011,N_14563,N_13870);
xor UO_1012 (O_1012,N_14498,N_14509);
xor UO_1013 (O_1013,N_14193,N_14535);
and UO_1014 (O_1014,N_14566,N_13578);
and UO_1015 (O_1015,N_14007,N_14890);
and UO_1016 (O_1016,N_14929,N_14765);
xor UO_1017 (O_1017,N_13789,N_14605);
and UO_1018 (O_1018,N_13627,N_14223);
nand UO_1019 (O_1019,N_14343,N_13966);
nor UO_1020 (O_1020,N_14290,N_14888);
and UO_1021 (O_1021,N_14847,N_14525);
or UO_1022 (O_1022,N_14817,N_13541);
nand UO_1023 (O_1023,N_13593,N_14245);
nand UO_1024 (O_1024,N_14421,N_13779);
and UO_1025 (O_1025,N_13779,N_13605);
xnor UO_1026 (O_1026,N_13931,N_13716);
nand UO_1027 (O_1027,N_13960,N_13610);
nand UO_1028 (O_1028,N_14001,N_14888);
nand UO_1029 (O_1029,N_14337,N_14221);
nand UO_1030 (O_1030,N_13652,N_14911);
xnor UO_1031 (O_1031,N_14032,N_14416);
and UO_1032 (O_1032,N_14886,N_14249);
and UO_1033 (O_1033,N_14464,N_13716);
nand UO_1034 (O_1034,N_14432,N_13948);
xnor UO_1035 (O_1035,N_13677,N_14109);
or UO_1036 (O_1036,N_14903,N_14482);
and UO_1037 (O_1037,N_14586,N_14427);
and UO_1038 (O_1038,N_13578,N_13736);
and UO_1039 (O_1039,N_14022,N_13831);
and UO_1040 (O_1040,N_14648,N_13560);
or UO_1041 (O_1041,N_14375,N_14051);
nor UO_1042 (O_1042,N_14414,N_13540);
nor UO_1043 (O_1043,N_14445,N_13545);
and UO_1044 (O_1044,N_14389,N_14546);
xor UO_1045 (O_1045,N_13842,N_14115);
and UO_1046 (O_1046,N_14629,N_14867);
xor UO_1047 (O_1047,N_14608,N_14276);
nor UO_1048 (O_1048,N_14299,N_14987);
xnor UO_1049 (O_1049,N_14933,N_14733);
or UO_1050 (O_1050,N_13988,N_13570);
and UO_1051 (O_1051,N_14708,N_14138);
nor UO_1052 (O_1052,N_14463,N_14842);
nor UO_1053 (O_1053,N_13738,N_14944);
and UO_1054 (O_1054,N_13777,N_14803);
nor UO_1055 (O_1055,N_13995,N_14029);
nand UO_1056 (O_1056,N_13913,N_14473);
nand UO_1057 (O_1057,N_14411,N_14815);
xnor UO_1058 (O_1058,N_14274,N_13762);
or UO_1059 (O_1059,N_13987,N_14892);
or UO_1060 (O_1060,N_14654,N_14691);
xor UO_1061 (O_1061,N_14360,N_14529);
xnor UO_1062 (O_1062,N_14118,N_14545);
or UO_1063 (O_1063,N_14900,N_14106);
xor UO_1064 (O_1064,N_14876,N_14971);
and UO_1065 (O_1065,N_13720,N_13704);
nor UO_1066 (O_1066,N_14115,N_13995);
nand UO_1067 (O_1067,N_14794,N_14376);
nor UO_1068 (O_1068,N_14892,N_13844);
nor UO_1069 (O_1069,N_14577,N_14475);
nor UO_1070 (O_1070,N_13781,N_13552);
or UO_1071 (O_1071,N_14540,N_14134);
and UO_1072 (O_1072,N_13942,N_14551);
xor UO_1073 (O_1073,N_14613,N_14063);
xor UO_1074 (O_1074,N_14998,N_14748);
and UO_1075 (O_1075,N_14509,N_14000);
or UO_1076 (O_1076,N_14912,N_13766);
nand UO_1077 (O_1077,N_13745,N_14290);
nand UO_1078 (O_1078,N_13727,N_13571);
or UO_1079 (O_1079,N_13693,N_14117);
and UO_1080 (O_1080,N_13979,N_14487);
nand UO_1081 (O_1081,N_14433,N_14888);
xor UO_1082 (O_1082,N_14365,N_13930);
nand UO_1083 (O_1083,N_14469,N_14607);
nand UO_1084 (O_1084,N_14454,N_13533);
xnor UO_1085 (O_1085,N_14235,N_14258);
or UO_1086 (O_1086,N_13990,N_14645);
xor UO_1087 (O_1087,N_14677,N_13687);
nand UO_1088 (O_1088,N_14577,N_14816);
nand UO_1089 (O_1089,N_14473,N_14721);
nand UO_1090 (O_1090,N_13934,N_14109);
nor UO_1091 (O_1091,N_14570,N_14533);
and UO_1092 (O_1092,N_13503,N_13578);
and UO_1093 (O_1093,N_13693,N_14408);
and UO_1094 (O_1094,N_14700,N_14901);
and UO_1095 (O_1095,N_13685,N_14835);
or UO_1096 (O_1096,N_14232,N_14836);
nand UO_1097 (O_1097,N_13988,N_14558);
nand UO_1098 (O_1098,N_13838,N_14858);
nand UO_1099 (O_1099,N_14930,N_13795);
or UO_1100 (O_1100,N_13546,N_13954);
nor UO_1101 (O_1101,N_14046,N_14053);
nor UO_1102 (O_1102,N_13729,N_13937);
nand UO_1103 (O_1103,N_14842,N_13545);
nand UO_1104 (O_1104,N_14401,N_13776);
and UO_1105 (O_1105,N_14373,N_14818);
nor UO_1106 (O_1106,N_14669,N_13982);
or UO_1107 (O_1107,N_14876,N_14020);
and UO_1108 (O_1108,N_13787,N_14962);
nand UO_1109 (O_1109,N_13631,N_14298);
and UO_1110 (O_1110,N_14405,N_14678);
or UO_1111 (O_1111,N_14120,N_14720);
and UO_1112 (O_1112,N_14579,N_14974);
xnor UO_1113 (O_1113,N_14816,N_14290);
xnor UO_1114 (O_1114,N_13841,N_13647);
xor UO_1115 (O_1115,N_13894,N_14864);
or UO_1116 (O_1116,N_14040,N_13763);
and UO_1117 (O_1117,N_13768,N_13674);
and UO_1118 (O_1118,N_14568,N_13604);
nor UO_1119 (O_1119,N_14217,N_14863);
xnor UO_1120 (O_1120,N_13756,N_14339);
and UO_1121 (O_1121,N_13890,N_14356);
nor UO_1122 (O_1122,N_14967,N_14442);
nor UO_1123 (O_1123,N_14760,N_14793);
xor UO_1124 (O_1124,N_14742,N_14305);
nor UO_1125 (O_1125,N_14305,N_14748);
and UO_1126 (O_1126,N_13600,N_14704);
nor UO_1127 (O_1127,N_14891,N_14039);
nor UO_1128 (O_1128,N_13629,N_14602);
and UO_1129 (O_1129,N_14244,N_14372);
xor UO_1130 (O_1130,N_14728,N_14547);
and UO_1131 (O_1131,N_13520,N_14133);
nand UO_1132 (O_1132,N_14967,N_14342);
xor UO_1133 (O_1133,N_14115,N_14752);
nand UO_1134 (O_1134,N_14629,N_14191);
xor UO_1135 (O_1135,N_14738,N_14580);
nand UO_1136 (O_1136,N_14889,N_14920);
nand UO_1137 (O_1137,N_13828,N_14772);
xor UO_1138 (O_1138,N_14946,N_13676);
and UO_1139 (O_1139,N_14864,N_13899);
nor UO_1140 (O_1140,N_13636,N_13661);
or UO_1141 (O_1141,N_13544,N_13690);
nor UO_1142 (O_1142,N_13828,N_14936);
nand UO_1143 (O_1143,N_14620,N_14666);
or UO_1144 (O_1144,N_13855,N_14952);
xnor UO_1145 (O_1145,N_13991,N_14874);
and UO_1146 (O_1146,N_13922,N_14407);
xnor UO_1147 (O_1147,N_13684,N_13857);
or UO_1148 (O_1148,N_14155,N_13858);
or UO_1149 (O_1149,N_14664,N_14131);
xor UO_1150 (O_1150,N_13745,N_14057);
xor UO_1151 (O_1151,N_14581,N_14876);
xor UO_1152 (O_1152,N_14210,N_14444);
and UO_1153 (O_1153,N_14828,N_13754);
nand UO_1154 (O_1154,N_13633,N_14766);
xnor UO_1155 (O_1155,N_14144,N_13500);
xnor UO_1156 (O_1156,N_13640,N_13776);
xor UO_1157 (O_1157,N_14706,N_14777);
and UO_1158 (O_1158,N_13577,N_13615);
or UO_1159 (O_1159,N_14292,N_13513);
nor UO_1160 (O_1160,N_14457,N_14648);
nand UO_1161 (O_1161,N_14614,N_13757);
xnor UO_1162 (O_1162,N_14593,N_13839);
and UO_1163 (O_1163,N_14831,N_14271);
nand UO_1164 (O_1164,N_14417,N_14238);
or UO_1165 (O_1165,N_14765,N_14574);
nor UO_1166 (O_1166,N_13544,N_13953);
or UO_1167 (O_1167,N_13966,N_14520);
nor UO_1168 (O_1168,N_13560,N_14176);
and UO_1169 (O_1169,N_13779,N_14065);
and UO_1170 (O_1170,N_13888,N_13851);
and UO_1171 (O_1171,N_13936,N_14911);
xnor UO_1172 (O_1172,N_14418,N_14670);
nor UO_1173 (O_1173,N_14316,N_14440);
nand UO_1174 (O_1174,N_13650,N_14252);
xor UO_1175 (O_1175,N_14718,N_13757);
xor UO_1176 (O_1176,N_14162,N_14422);
nand UO_1177 (O_1177,N_13886,N_14514);
nor UO_1178 (O_1178,N_13857,N_14027);
xor UO_1179 (O_1179,N_13910,N_14228);
nand UO_1180 (O_1180,N_14055,N_14346);
and UO_1181 (O_1181,N_14923,N_14660);
and UO_1182 (O_1182,N_13938,N_13631);
nor UO_1183 (O_1183,N_13633,N_13996);
or UO_1184 (O_1184,N_14628,N_14072);
or UO_1185 (O_1185,N_14845,N_14640);
nor UO_1186 (O_1186,N_13900,N_14031);
nor UO_1187 (O_1187,N_14523,N_14531);
xnor UO_1188 (O_1188,N_13788,N_13930);
nor UO_1189 (O_1189,N_13729,N_14017);
nor UO_1190 (O_1190,N_13962,N_14277);
and UO_1191 (O_1191,N_13804,N_14110);
or UO_1192 (O_1192,N_14124,N_13947);
xor UO_1193 (O_1193,N_14064,N_13633);
xor UO_1194 (O_1194,N_14520,N_13883);
or UO_1195 (O_1195,N_13968,N_14293);
and UO_1196 (O_1196,N_14598,N_13695);
nor UO_1197 (O_1197,N_14980,N_14361);
xor UO_1198 (O_1198,N_14299,N_13861);
xnor UO_1199 (O_1199,N_13975,N_13940);
xnor UO_1200 (O_1200,N_14794,N_14487);
xor UO_1201 (O_1201,N_14886,N_13712);
or UO_1202 (O_1202,N_13521,N_14099);
xor UO_1203 (O_1203,N_14629,N_14458);
xor UO_1204 (O_1204,N_13909,N_13779);
xnor UO_1205 (O_1205,N_14246,N_14753);
nand UO_1206 (O_1206,N_14782,N_14379);
nor UO_1207 (O_1207,N_13746,N_14054);
xnor UO_1208 (O_1208,N_14035,N_14586);
nor UO_1209 (O_1209,N_13829,N_14082);
nor UO_1210 (O_1210,N_14500,N_13621);
and UO_1211 (O_1211,N_13792,N_14967);
nand UO_1212 (O_1212,N_14642,N_13782);
nand UO_1213 (O_1213,N_14767,N_13628);
nand UO_1214 (O_1214,N_13820,N_14825);
or UO_1215 (O_1215,N_13750,N_14738);
xnor UO_1216 (O_1216,N_14451,N_14094);
or UO_1217 (O_1217,N_14345,N_14491);
xor UO_1218 (O_1218,N_14527,N_13884);
or UO_1219 (O_1219,N_14363,N_14584);
or UO_1220 (O_1220,N_14087,N_13651);
or UO_1221 (O_1221,N_14623,N_14479);
xor UO_1222 (O_1222,N_14422,N_14684);
nand UO_1223 (O_1223,N_13872,N_13577);
nor UO_1224 (O_1224,N_14678,N_13577);
and UO_1225 (O_1225,N_14106,N_14484);
xnor UO_1226 (O_1226,N_14337,N_14409);
nor UO_1227 (O_1227,N_14774,N_14174);
and UO_1228 (O_1228,N_14623,N_14143);
nor UO_1229 (O_1229,N_14383,N_14871);
and UO_1230 (O_1230,N_14810,N_14556);
and UO_1231 (O_1231,N_13749,N_14222);
nand UO_1232 (O_1232,N_14547,N_13934);
and UO_1233 (O_1233,N_13624,N_13795);
and UO_1234 (O_1234,N_14680,N_13913);
nand UO_1235 (O_1235,N_14943,N_13592);
nor UO_1236 (O_1236,N_14766,N_14060);
nand UO_1237 (O_1237,N_14937,N_14558);
nor UO_1238 (O_1238,N_14833,N_13568);
and UO_1239 (O_1239,N_14302,N_13818);
nor UO_1240 (O_1240,N_14349,N_14241);
nor UO_1241 (O_1241,N_14029,N_14403);
or UO_1242 (O_1242,N_14147,N_14280);
nand UO_1243 (O_1243,N_14608,N_14984);
and UO_1244 (O_1244,N_13978,N_13984);
nand UO_1245 (O_1245,N_13905,N_14377);
nand UO_1246 (O_1246,N_13814,N_13850);
or UO_1247 (O_1247,N_14474,N_13918);
xor UO_1248 (O_1248,N_14826,N_14981);
or UO_1249 (O_1249,N_13805,N_14074);
nand UO_1250 (O_1250,N_13981,N_14439);
nand UO_1251 (O_1251,N_13786,N_14639);
nand UO_1252 (O_1252,N_14295,N_14268);
or UO_1253 (O_1253,N_13737,N_14614);
nor UO_1254 (O_1254,N_13792,N_13868);
nor UO_1255 (O_1255,N_13931,N_14890);
nor UO_1256 (O_1256,N_13687,N_14867);
nand UO_1257 (O_1257,N_14076,N_14631);
or UO_1258 (O_1258,N_13956,N_14604);
xnor UO_1259 (O_1259,N_13542,N_14799);
or UO_1260 (O_1260,N_13996,N_14924);
and UO_1261 (O_1261,N_14434,N_14823);
nand UO_1262 (O_1262,N_13602,N_14623);
or UO_1263 (O_1263,N_14712,N_13713);
xor UO_1264 (O_1264,N_14550,N_14725);
xor UO_1265 (O_1265,N_13607,N_14395);
nand UO_1266 (O_1266,N_14733,N_13594);
or UO_1267 (O_1267,N_14381,N_13839);
and UO_1268 (O_1268,N_14871,N_14458);
xnor UO_1269 (O_1269,N_14241,N_14104);
nor UO_1270 (O_1270,N_14512,N_13818);
nor UO_1271 (O_1271,N_14277,N_14761);
xor UO_1272 (O_1272,N_14249,N_14302);
nor UO_1273 (O_1273,N_14141,N_14716);
nand UO_1274 (O_1274,N_13887,N_14198);
xor UO_1275 (O_1275,N_14971,N_13903);
nand UO_1276 (O_1276,N_14621,N_13723);
and UO_1277 (O_1277,N_14011,N_14818);
xor UO_1278 (O_1278,N_14418,N_14542);
and UO_1279 (O_1279,N_14079,N_14650);
xor UO_1280 (O_1280,N_14213,N_13526);
nand UO_1281 (O_1281,N_13944,N_14722);
and UO_1282 (O_1282,N_14640,N_13883);
nand UO_1283 (O_1283,N_13725,N_14868);
xnor UO_1284 (O_1284,N_14687,N_13972);
xnor UO_1285 (O_1285,N_14174,N_14312);
xor UO_1286 (O_1286,N_14506,N_14466);
xor UO_1287 (O_1287,N_14653,N_14678);
or UO_1288 (O_1288,N_14333,N_13609);
or UO_1289 (O_1289,N_14749,N_13616);
nand UO_1290 (O_1290,N_14320,N_14667);
nor UO_1291 (O_1291,N_13511,N_13544);
or UO_1292 (O_1292,N_13834,N_14051);
or UO_1293 (O_1293,N_14189,N_14352);
and UO_1294 (O_1294,N_13585,N_14002);
or UO_1295 (O_1295,N_13587,N_14603);
xor UO_1296 (O_1296,N_14782,N_13521);
nand UO_1297 (O_1297,N_13858,N_13937);
nor UO_1298 (O_1298,N_14156,N_13933);
nand UO_1299 (O_1299,N_13729,N_14071);
xor UO_1300 (O_1300,N_14456,N_14168);
nand UO_1301 (O_1301,N_14279,N_14864);
or UO_1302 (O_1302,N_14375,N_14539);
xor UO_1303 (O_1303,N_14451,N_14668);
nand UO_1304 (O_1304,N_14390,N_13799);
nand UO_1305 (O_1305,N_14174,N_14262);
and UO_1306 (O_1306,N_13609,N_14514);
or UO_1307 (O_1307,N_14685,N_14947);
nor UO_1308 (O_1308,N_14767,N_13863);
or UO_1309 (O_1309,N_14448,N_13945);
nor UO_1310 (O_1310,N_14983,N_13942);
nor UO_1311 (O_1311,N_13655,N_13573);
or UO_1312 (O_1312,N_14658,N_14843);
and UO_1313 (O_1313,N_14240,N_13921);
and UO_1314 (O_1314,N_14764,N_14891);
xor UO_1315 (O_1315,N_14277,N_13830);
nor UO_1316 (O_1316,N_13522,N_14771);
nand UO_1317 (O_1317,N_13898,N_13992);
or UO_1318 (O_1318,N_14114,N_14478);
and UO_1319 (O_1319,N_14609,N_13781);
xor UO_1320 (O_1320,N_14789,N_13666);
or UO_1321 (O_1321,N_14692,N_14643);
or UO_1322 (O_1322,N_14392,N_14211);
or UO_1323 (O_1323,N_14501,N_14109);
nand UO_1324 (O_1324,N_14938,N_13824);
and UO_1325 (O_1325,N_14461,N_14816);
nor UO_1326 (O_1326,N_13811,N_14758);
or UO_1327 (O_1327,N_14982,N_14484);
and UO_1328 (O_1328,N_13509,N_14716);
xnor UO_1329 (O_1329,N_13930,N_13736);
nand UO_1330 (O_1330,N_14202,N_13619);
nor UO_1331 (O_1331,N_13619,N_13656);
or UO_1332 (O_1332,N_14907,N_14958);
or UO_1333 (O_1333,N_13978,N_14815);
xnor UO_1334 (O_1334,N_13927,N_13634);
and UO_1335 (O_1335,N_14144,N_14278);
xor UO_1336 (O_1336,N_14277,N_14376);
and UO_1337 (O_1337,N_14555,N_13859);
nand UO_1338 (O_1338,N_14399,N_13815);
or UO_1339 (O_1339,N_14252,N_13792);
xor UO_1340 (O_1340,N_14645,N_14799);
or UO_1341 (O_1341,N_14337,N_13875);
nor UO_1342 (O_1342,N_13878,N_14690);
and UO_1343 (O_1343,N_14793,N_14479);
nor UO_1344 (O_1344,N_14658,N_13754);
nand UO_1345 (O_1345,N_14946,N_14108);
nand UO_1346 (O_1346,N_14529,N_13559);
nand UO_1347 (O_1347,N_14170,N_14783);
nor UO_1348 (O_1348,N_13559,N_13831);
and UO_1349 (O_1349,N_14247,N_14057);
nand UO_1350 (O_1350,N_14969,N_14641);
or UO_1351 (O_1351,N_13547,N_14877);
or UO_1352 (O_1352,N_14646,N_14843);
xnor UO_1353 (O_1353,N_13521,N_13672);
nor UO_1354 (O_1354,N_13958,N_14162);
nor UO_1355 (O_1355,N_13740,N_14553);
nand UO_1356 (O_1356,N_14638,N_14281);
xnor UO_1357 (O_1357,N_13784,N_13778);
and UO_1358 (O_1358,N_13508,N_14651);
or UO_1359 (O_1359,N_14845,N_14104);
xnor UO_1360 (O_1360,N_14921,N_14141);
and UO_1361 (O_1361,N_14956,N_14259);
and UO_1362 (O_1362,N_13765,N_14678);
nor UO_1363 (O_1363,N_14350,N_13905);
nor UO_1364 (O_1364,N_14136,N_13640);
nand UO_1365 (O_1365,N_13571,N_13839);
or UO_1366 (O_1366,N_14082,N_13526);
and UO_1367 (O_1367,N_14286,N_14338);
xnor UO_1368 (O_1368,N_14516,N_13724);
nor UO_1369 (O_1369,N_14997,N_14870);
xor UO_1370 (O_1370,N_14430,N_14658);
nor UO_1371 (O_1371,N_14357,N_14541);
or UO_1372 (O_1372,N_13941,N_14902);
xor UO_1373 (O_1373,N_14340,N_13890);
or UO_1374 (O_1374,N_13503,N_14831);
or UO_1375 (O_1375,N_14490,N_14996);
xnor UO_1376 (O_1376,N_14975,N_14221);
nor UO_1377 (O_1377,N_14055,N_14151);
nand UO_1378 (O_1378,N_14830,N_14332);
xor UO_1379 (O_1379,N_14611,N_13558);
and UO_1380 (O_1380,N_14206,N_14659);
nand UO_1381 (O_1381,N_14447,N_14224);
nor UO_1382 (O_1382,N_14291,N_13671);
nand UO_1383 (O_1383,N_13908,N_14259);
xnor UO_1384 (O_1384,N_14849,N_13873);
and UO_1385 (O_1385,N_14089,N_13758);
or UO_1386 (O_1386,N_14971,N_13667);
xor UO_1387 (O_1387,N_14545,N_14960);
or UO_1388 (O_1388,N_14240,N_14575);
nor UO_1389 (O_1389,N_14078,N_13862);
or UO_1390 (O_1390,N_13632,N_14748);
or UO_1391 (O_1391,N_13930,N_14637);
nor UO_1392 (O_1392,N_14276,N_13696);
xor UO_1393 (O_1393,N_14988,N_13929);
xnor UO_1394 (O_1394,N_13640,N_14434);
nor UO_1395 (O_1395,N_14966,N_14115);
and UO_1396 (O_1396,N_14693,N_14375);
or UO_1397 (O_1397,N_13782,N_14076);
nand UO_1398 (O_1398,N_14173,N_13723);
xor UO_1399 (O_1399,N_14214,N_14225);
xnor UO_1400 (O_1400,N_13752,N_13744);
nor UO_1401 (O_1401,N_14264,N_13595);
nand UO_1402 (O_1402,N_13671,N_14504);
nand UO_1403 (O_1403,N_13548,N_14075);
nor UO_1404 (O_1404,N_13675,N_14830);
nor UO_1405 (O_1405,N_13863,N_14061);
or UO_1406 (O_1406,N_14431,N_14662);
nor UO_1407 (O_1407,N_13799,N_14815);
nand UO_1408 (O_1408,N_13818,N_13597);
nor UO_1409 (O_1409,N_13534,N_13617);
and UO_1410 (O_1410,N_14870,N_14069);
nor UO_1411 (O_1411,N_13748,N_14197);
and UO_1412 (O_1412,N_14646,N_14523);
xnor UO_1413 (O_1413,N_14235,N_14377);
and UO_1414 (O_1414,N_14080,N_13675);
nor UO_1415 (O_1415,N_13642,N_14507);
and UO_1416 (O_1416,N_13666,N_14710);
and UO_1417 (O_1417,N_14810,N_13803);
and UO_1418 (O_1418,N_14462,N_13753);
xnor UO_1419 (O_1419,N_13966,N_14240);
or UO_1420 (O_1420,N_13534,N_13771);
and UO_1421 (O_1421,N_13757,N_14925);
nor UO_1422 (O_1422,N_14160,N_14604);
xor UO_1423 (O_1423,N_14657,N_13830);
xor UO_1424 (O_1424,N_14974,N_13824);
nand UO_1425 (O_1425,N_14516,N_13523);
nor UO_1426 (O_1426,N_14067,N_13570);
nand UO_1427 (O_1427,N_14517,N_14439);
or UO_1428 (O_1428,N_14748,N_14766);
or UO_1429 (O_1429,N_13643,N_13765);
nor UO_1430 (O_1430,N_14452,N_14535);
or UO_1431 (O_1431,N_13717,N_14898);
xnor UO_1432 (O_1432,N_13656,N_13770);
and UO_1433 (O_1433,N_14312,N_14209);
xnor UO_1434 (O_1434,N_14682,N_13638);
nor UO_1435 (O_1435,N_14171,N_13704);
xor UO_1436 (O_1436,N_13617,N_14004);
and UO_1437 (O_1437,N_13898,N_14874);
nand UO_1438 (O_1438,N_14520,N_13869);
nand UO_1439 (O_1439,N_13628,N_14268);
xnor UO_1440 (O_1440,N_14593,N_14197);
nor UO_1441 (O_1441,N_14651,N_14538);
nor UO_1442 (O_1442,N_14721,N_13765);
or UO_1443 (O_1443,N_13555,N_14282);
or UO_1444 (O_1444,N_14308,N_14671);
nor UO_1445 (O_1445,N_14110,N_14195);
nand UO_1446 (O_1446,N_13803,N_13513);
or UO_1447 (O_1447,N_14439,N_14771);
nand UO_1448 (O_1448,N_14066,N_14007);
nor UO_1449 (O_1449,N_14482,N_13951);
xor UO_1450 (O_1450,N_13845,N_13602);
and UO_1451 (O_1451,N_14385,N_14305);
or UO_1452 (O_1452,N_13964,N_13599);
xnor UO_1453 (O_1453,N_13936,N_14983);
xor UO_1454 (O_1454,N_14555,N_14343);
or UO_1455 (O_1455,N_14487,N_14174);
nand UO_1456 (O_1456,N_14086,N_13530);
or UO_1457 (O_1457,N_13731,N_13682);
xor UO_1458 (O_1458,N_13850,N_13594);
nor UO_1459 (O_1459,N_14938,N_14821);
nor UO_1460 (O_1460,N_14146,N_13918);
nand UO_1461 (O_1461,N_14409,N_14525);
or UO_1462 (O_1462,N_13772,N_14383);
or UO_1463 (O_1463,N_14468,N_13596);
xnor UO_1464 (O_1464,N_13550,N_13644);
nor UO_1465 (O_1465,N_14218,N_14460);
xnor UO_1466 (O_1466,N_13980,N_14836);
and UO_1467 (O_1467,N_14125,N_14789);
nand UO_1468 (O_1468,N_14834,N_14873);
nor UO_1469 (O_1469,N_13508,N_14462);
and UO_1470 (O_1470,N_14391,N_14563);
nand UO_1471 (O_1471,N_14395,N_14140);
xor UO_1472 (O_1472,N_13701,N_13509);
nand UO_1473 (O_1473,N_14513,N_14135);
nand UO_1474 (O_1474,N_14370,N_13687);
nor UO_1475 (O_1475,N_14331,N_14553);
and UO_1476 (O_1476,N_14877,N_14543);
nand UO_1477 (O_1477,N_14916,N_13599);
nor UO_1478 (O_1478,N_13829,N_14456);
xnor UO_1479 (O_1479,N_13558,N_13784);
and UO_1480 (O_1480,N_13718,N_13778);
nor UO_1481 (O_1481,N_13544,N_14906);
xnor UO_1482 (O_1482,N_14535,N_14692);
xnor UO_1483 (O_1483,N_14335,N_13569);
nor UO_1484 (O_1484,N_13558,N_14092);
xor UO_1485 (O_1485,N_14781,N_14265);
nand UO_1486 (O_1486,N_14875,N_14459);
nor UO_1487 (O_1487,N_13956,N_13775);
and UO_1488 (O_1488,N_14060,N_14583);
nor UO_1489 (O_1489,N_14060,N_14467);
and UO_1490 (O_1490,N_14279,N_13737);
nor UO_1491 (O_1491,N_14570,N_14966);
and UO_1492 (O_1492,N_13565,N_14097);
nor UO_1493 (O_1493,N_13708,N_14057);
nor UO_1494 (O_1494,N_14066,N_13912);
and UO_1495 (O_1495,N_14951,N_13970);
nor UO_1496 (O_1496,N_14222,N_13870);
xnor UO_1497 (O_1497,N_14752,N_14758);
and UO_1498 (O_1498,N_13743,N_14314);
xor UO_1499 (O_1499,N_13707,N_14832);
or UO_1500 (O_1500,N_14208,N_14081);
xor UO_1501 (O_1501,N_13879,N_14943);
nor UO_1502 (O_1502,N_14774,N_14671);
nor UO_1503 (O_1503,N_14359,N_13752);
nor UO_1504 (O_1504,N_14971,N_13650);
xor UO_1505 (O_1505,N_14293,N_14452);
nand UO_1506 (O_1506,N_14861,N_13531);
or UO_1507 (O_1507,N_14246,N_14423);
or UO_1508 (O_1508,N_14663,N_14584);
nor UO_1509 (O_1509,N_14357,N_13507);
nand UO_1510 (O_1510,N_14085,N_14656);
and UO_1511 (O_1511,N_13665,N_14384);
xor UO_1512 (O_1512,N_13730,N_14965);
or UO_1513 (O_1513,N_14370,N_13658);
or UO_1514 (O_1514,N_14117,N_14151);
or UO_1515 (O_1515,N_14894,N_14240);
and UO_1516 (O_1516,N_14287,N_13970);
xor UO_1517 (O_1517,N_13594,N_13555);
xnor UO_1518 (O_1518,N_14065,N_14459);
and UO_1519 (O_1519,N_13758,N_13935);
and UO_1520 (O_1520,N_13761,N_13795);
and UO_1521 (O_1521,N_14207,N_14288);
or UO_1522 (O_1522,N_13790,N_13814);
and UO_1523 (O_1523,N_13584,N_14329);
xnor UO_1524 (O_1524,N_13534,N_13774);
or UO_1525 (O_1525,N_14479,N_13804);
xor UO_1526 (O_1526,N_13915,N_13654);
nor UO_1527 (O_1527,N_14583,N_14687);
or UO_1528 (O_1528,N_14201,N_14417);
or UO_1529 (O_1529,N_13961,N_14656);
xnor UO_1530 (O_1530,N_14518,N_13894);
and UO_1531 (O_1531,N_14069,N_13785);
and UO_1532 (O_1532,N_14971,N_13772);
and UO_1533 (O_1533,N_13899,N_13500);
nand UO_1534 (O_1534,N_14670,N_14258);
xnor UO_1535 (O_1535,N_14821,N_14029);
or UO_1536 (O_1536,N_14225,N_14047);
and UO_1537 (O_1537,N_14362,N_14137);
or UO_1538 (O_1538,N_13627,N_13863);
xor UO_1539 (O_1539,N_13709,N_14678);
and UO_1540 (O_1540,N_14144,N_14742);
or UO_1541 (O_1541,N_13795,N_14080);
xnor UO_1542 (O_1542,N_14063,N_13796);
nand UO_1543 (O_1543,N_14794,N_14630);
or UO_1544 (O_1544,N_13829,N_14331);
or UO_1545 (O_1545,N_14648,N_14316);
and UO_1546 (O_1546,N_13917,N_14603);
nor UO_1547 (O_1547,N_14828,N_14434);
and UO_1548 (O_1548,N_14245,N_13833);
xnor UO_1549 (O_1549,N_14894,N_13695);
and UO_1550 (O_1550,N_14271,N_13867);
or UO_1551 (O_1551,N_13554,N_13894);
nor UO_1552 (O_1552,N_13601,N_14724);
nand UO_1553 (O_1553,N_14048,N_14146);
and UO_1554 (O_1554,N_14006,N_14017);
nor UO_1555 (O_1555,N_14504,N_14735);
nand UO_1556 (O_1556,N_14549,N_14126);
xnor UO_1557 (O_1557,N_14995,N_13900);
nor UO_1558 (O_1558,N_14522,N_14852);
nor UO_1559 (O_1559,N_13746,N_13822);
or UO_1560 (O_1560,N_14675,N_14535);
and UO_1561 (O_1561,N_14413,N_13902);
and UO_1562 (O_1562,N_13895,N_14798);
nor UO_1563 (O_1563,N_14034,N_14328);
nor UO_1564 (O_1564,N_14739,N_13526);
and UO_1565 (O_1565,N_14931,N_14710);
nor UO_1566 (O_1566,N_14467,N_14515);
nand UO_1567 (O_1567,N_14751,N_14989);
nor UO_1568 (O_1568,N_14161,N_14313);
nand UO_1569 (O_1569,N_14575,N_14287);
nor UO_1570 (O_1570,N_13787,N_13661);
xnor UO_1571 (O_1571,N_13680,N_14028);
nor UO_1572 (O_1572,N_14442,N_14882);
xor UO_1573 (O_1573,N_13634,N_13971);
xor UO_1574 (O_1574,N_13629,N_13648);
nand UO_1575 (O_1575,N_13604,N_14369);
and UO_1576 (O_1576,N_14814,N_13747);
nor UO_1577 (O_1577,N_13836,N_14004);
nor UO_1578 (O_1578,N_13715,N_14755);
nand UO_1579 (O_1579,N_14757,N_14795);
nand UO_1580 (O_1580,N_14458,N_14417);
nor UO_1581 (O_1581,N_13847,N_13792);
or UO_1582 (O_1582,N_13576,N_14783);
xor UO_1583 (O_1583,N_14991,N_14778);
xor UO_1584 (O_1584,N_14380,N_14370);
nor UO_1585 (O_1585,N_14014,N_14894);
nand UO_1586 (O_1586,N_14759,N_13957);
xnor UO_1587 (O_1587,N_13953,N_13938);
xnor UO_1588 (O_1588,N_14440,N_14471);
nor UO_1589 (O_1589,N_14389,N_14661);
xnor UO_1590 (O_1590,N_14848,N_13561);
nor UO_1591 (O_1591,N_14397,N_14956);
or UO_1592 (O_1592,N_13985,N_13801);
or UO_1593 (O_1593,N_14329,N_13643);
and UO_1594 (O_1594,N_13701,N_13622);
nand UO_1595 (O_1595,N_13997,N_14604);
or UO_1596 (O_1596,N_13885,N_14580);
nor UO_1597 (O_1597,N_13940,N_14750);
and UO_1598 (O_1598,N_14256,N_13918);
and UO_1599 (O_1599,N_14659,N_14984);
nor UO_1600 (O_1600,N_14045,N_14676);
xnor UO_1601 (O_1601,N_14925,N_13788);
xnor UO_1602 (O_1602,N_14052,N_14928);
xnor UO_1603 (O_1603,N_13784,N_13848);
or UO_1604 (O_1604,N_13508,N_14328);
and UO_1605 (O_1605,N_14302,N_14639);
nand UO_1606 (O_1606,N_13632,N_14984);
nor UO_1607 (O_1607,N_14483,N_13558);
nand UO_1608 (O_1608,N_14772,N_14913);
nor UO_1609 (O_1609,N_14268,N_14867);
nand UO_1610 (O_1610,N_13959,N_14617);
nor UO_1611 (O_1611,N_14000,N_14233);
nor UO_1612 (O_1612,N_14386,N_14784);
nand UO_1613 (O_1613,N_14942,N_13795);
xnor UO_1614 (O_1614,N_13558,N_13914);
xor UO_1615 (O_1615,N_14517,N_13622);
nor UO_1616 (O_1616,N_14511,N_14104);
nand UO_1617 (O_1617,N_14554,N_13751);
nand UO_1618 (O_1618,N_14671,N_14736);
or UO_1619 (O_1619,N_14762,N_14160);
xor UO_1620 (O_1620,N_14894,N_13985);
nor UO_1621 (O_1621,N_13711,N_14949);
nand UO_1622 (O_1622,N_14665,N_13987);
nor UO_1623 (O_1623,N_13658,N_14862);
xor UO_1624 (O_1624,N_13532,N_13993);
or UO_1625 (O_1625,N_14364,N_14437);
nor UO_1626 (O_1626,N_14995,N_14626);
and UO_1627 (O_1627,N_13610,N_13630);
nor UO_1628 (O_1628,N_14071,N_14032);
nand UO_1629 (O_1629,N_14644,N_13938);
nor UO_1630 (O_1630,N_14801,N_14379);
and UO_1631 (O_1631,N_14448,N_14810);
nor UO_1632 (O_1632,N_13951,N_14082);
xor UO_1633 (O_1633,N_14294,N_14689);
xor UO_1634 (O_1634,N_14517,N_13874);
xor UO_1635 (O_1635,N_14403,N_14729);
nand UO_1636 (O_1636,N_13932,N_13692);
and UO_1637 (O_1637,N_13981,N_13766);
xnor UO_1638 (O_1638,N_14109,N_14996);
nor UO_1639 (O_1639,N_14530,N_13766);
xnor UO_1640 (O_1640,N_14385,N_13781);
and UO_1641 (O_1641,N_14772,N_14215);
nor UO_1642 (O_1642,N_13962,N_14349);
or UO_1643 (O_1643,N_13951,N_13620);
nand UO_1644 (O_1644,N_13624,N_13844);
or UO_1645 (O_1645,N_14697,N_13663);
xor UO_1646 (O_1646,N_14985,N_14612);
nor UO_1647 (O_1647,N_14658,N_13868);
nor UO_1648 (O_1648,N_14984,N_13781);
xor UO_1649 (O_1649,N_14703,N_14677);
and UO_1650 (O_1650,N_14508,N_14750);
and UO_1651 (O_1651,N_14390,N_14821);
or UO_1652 (O_1652,N_14092,N_13569);
xnor UO_1653 (O_1653,N_13719,N_13515);
nor UO_1654 (O_1654,N_14239,N_13892);
or UO_1655 (O_1655,N_14380,N_14715);
nor UO_1656 (O_1656,N_14927,N_14736);
nor UO_1657 (O_1657,N_14341,N_14850);
nor UO_1658 (O_1658,N_14740,N_13618);
nor UO_1659 (O_1659,N_14447,N_14091);
nor UO_1660 (O_1660,N_14031,N_13717);
or UO_1661 (O_1661,N_14815,N_14892);
xor UO_1662 (O_1662,N_14008,N_13766);
and UO_1663 (O_1663,N_13779,N_14559);
or UO_1664 (O_1664,N_14597,N_14222);
or UO_1665 (O_1665,N_14970,N_14712);
and UO_1666 (O_1666,N_13677,N_14716);
nand UO_1667 (O_1667,N_14590,N_14550);
xnor UO_1668 (O_1668,N_14710,N_14197);
or UO_1669 (O_1669,N_14962,N_13935);
xnor UO_1670 (O_1670,N_14605,N_14716);
nor UO_1671 (O_1671,N_14950,N_14072);
or UO_1672 (O_1672,N_13889,N_13928);
nand UO_1673 (O_1673,N_14903,N_14479);
or UO_1674 (O_1674,N_14497,N_14767);
or UO_1675 (O_1675,N_14722,N_14406);
xor UO_1676 (O_1676,N_13881,N_14409);
nor UO_1677 (O_1677,N_13940,N_13695);
nor UO_1678 (O_1678,N_13550,N_14461);
and UO_1679 (O_1679,N_14389,N_14201);
and UO_1680 (O_1680,N_13812,N_13884);
xnor UO_1681 (O_1681,N_13866,N_13509);
nor UO_1682 (O_1682,N_14124,N_14894);
and UO_1683 (O_1683,N_14264,N_14692);
nor UO_1684 (O_1684,N_14083,N_14751);
or UO_1685 (O_1685,N_14665,N_14366);
xor UO_1686 (O_1686,N_13644,N_13693);
nand UO_1687 (O_1687,N_13968,N_14906);
xnor UO_1688 (O_1688,N_14237,N_13600);
xor UO_1689 (O_1689,N_14166,N_14760);
nand UO_1690 (O_1690,N_13779,N_14903);
nor UO_1691 (O_1691,N_14661,N_14739);
nor UO_1692 (O_1692,N_13958,N_14614);
and UO_1693 (O_1693,N_13999,N_13675);
nand UO_1694 (O_1694,N_14400,N_14460);
and UO_1695 (O_1695,N_14073,N_13697);
nor UO_1696 (O_1696,N_14420,N_14207);
or UO_1697 (O_1697,N_13713,N_14918);
and UO_1698 (O_1698,N_14288,N_14830);
nor UO_1699 (O_1699,N_13578,N_13663);
and UO_1700 (O_1700,N_14843,N_14838);
and UO_1701 (O_1701,N_13601,N_14079);
xnor UO_1702 (O_1702,N_13678,N_14075);
xor UO_1703 (O_1703,N_14671,N_14778);
or UO_1704 (O_1704,N_14348,N_14309);
xor UO_1705 (O_1705,N_14155,N_13925);
and UO_1706 (O_1706,N_13523,N_14671);
or UO_1707 (O_1707,N_13696,N_14057);
xor UO_1708 (O_1708,N_13589,N_14694);
and UO_1709 (O_1709,N_14246,N_13844);
or UO_1710 (O_1710,N_14449,N_13579);
nand UO_1711 (O_1711,N_14793,N_13594);
or UO_1712 (O_1712,N_13574,N_13958);
nor UO_1713 (O_1713,N_14606,N_14220);
or UO_1714 (O_1714,N_14789,N_14136);
nand UO_1715 (O_1715,N_14319,N_13618);
nand UO_1716 (O_1716,N_14412,N_14139);
nor UO_1717 (O_1717,N_14626,N_13811);
nand UO_1718 (O_1718,N_14396,N_13946);
xnor UO_1719 (O_1719,N_13578,N_13937);
nor UO_1720 (O_1720,N_14176,N_14861);
nor UO_1721 (O_1721,N_14398,N_14446);
nand UO_1722 (O_1722,N_14678,N_14079);
nor UO_1723 (O_1723,N_14094,N_13863);
and UO_1724 (O_1724,N_14246,N_14876);
nand UO_1725 (O_1725,N_14025,N_14854);
xnor UO_1726 (O_1726,N_14909,N_14329);
nand UO_1727 (O_1727,N_13650,N_14841);
xnor UO_1728 (O_1728,N_14182,N_14081);
nand UO_1729 (O_1729,N_14417,N_14425);
or UO_1730 (O_1730,N_14379,N_14684);
or UO_1731 (O_1731,N_13600,N_13942);
and UO_1732 (O_1732,N_14202,N_13734);
or UO_1733 (O_1733,N_14605,N_13967);
xnor UO_1734 (O_1734,N_14593,N_14262);
nand UO_1735 (O_1735,N_13594,N_13889);
nor UO_1736 (O_1736,N_14604,N_13951);
xor UO_1737 (O_1737,N_14135,N_14982);
xnor UO_1738 (O_1738,N_14690,N_13563);
and UO_1739 (O_1739,N_13771,N_14542);
nor UO_1740 (O_1740,N_14976,N_13674);
and UO_1741 (O_1741,N_13868,N_14567);
nand UO_1742 (O_1742,N_13728,N_13986);
xnor UO_1743 (O_1743,N_13507,N_13617);
or UO_1744 (O_1744,N_13595,N_14697);
xor UO_1745 (O_1745,N_14569,N_14125);
xor UO_1746 (O_1746,N_13824,N_14512);
or UO_1747 (O_1747,N_14963,N_14053);
xor UO_1748 (O_1748,N_13689,N_13787);
nor UO_1749 (O_1749,N_14436,N_14280);
or UO_1750 (O_1750,N_13570,N_13894);
and UO_1751 (O_1751,N_14269,N_14773);
and UO_1752 (O_1752,N_14488,N_14408);
and UO_1753 (O_1753,N_13998,N_14625);
xor UO_1754 (O_1754,N_14292,N_14391);
nor UO_1755 (O_1755,N_13644,N_13626);
xor UO_1756 (O_1756,N_14898,N_13678);
nand UO_1757 (O_1757,N_13532,N_14202);
xor UO_1758 (O_1758,N_13541,N_14335);
nand UO_1759 (O_1759,N_14129,N_13714);
xnor UO_1760 (O_1760,N_14630,N_13534);
nand UO_1761 (O_1761,N_13550,N_14296);
xnor UO_1762 (O_1762,N_14434,N_13637);
xnor UO_1763 (O_1763,N_14132,N_13707);
nand UO_1764 (O_1764,N_14414,N_13509);
xor UO_1765 (O_1765,N_13932,N_14569);
xnor UO_1766 (O_1766,N_14548,N_13772);
xor UO_1767 (O_1767,N_13747,N_13907);
or UO_1768 (O_1768,N_14325,N_14115);
xor UO_1769 (O_1769,N_14936,N_14551);
or UO_1770 (O_1770,N_14977,N_13780);
and UO_1771 (O_1771,N_13584,N_14914);
or UO_1772 (O_1772,N_13759,N_14883);
xnor UO_1773 (O_1773,N_14172,N_13748);
and UO_1774 (O_1774,N_14987,N_14193);
nand UO_1775 (O_1775,N_14576,N_14481);
nand UO_1776 (O_1776,N_14553,N_14269);
nand UO_1777 (O_1777,N_13713,N_14573);
nand UO_1778 (O_1778,N_14439,N_14748);
xnor UO_1779 (O_1779,N_14026,N_14370);
nor UO_1780 (O_1780,N_14885,N_13996);
and UO_1781 (O_1781,N_14720,N_13531);
nand UO_1782 (O_1782,N_13659,N_14735);
nand UO_1783 (O_1783,N_14168,N_14230);
nor UO_1784 (O_1784,N_14782,N_13626);
and UO_1785 (O_1785,N_14397,N_13757);
or UO_1786 (O_1786,N_14804,N_14698);
or UO_1787 (O_1787,N_13969,N_14839);
nand UO_1788 (O_1788,N_13526,N_14804);
xnor UO_1789 (O_1789,N_14326,N_13950);
xnor UO_1790 (O_1790,N_14474,N_14989);
nor UO_1791 (O_1791,N_14491,N_14207);
xor UO_1792 (O_1792,N_14147,N_14089);
xnor UO_1793 (O_1793,N_14848,N_14005);
nor UO_1794 (O_1794,N_14841,N_14197);
and UO_1795 (O_1795,N_13899,N_13934);
nand UO_1796 (O_1796,N_14475,N_13952);
nand UO_1797 (O_1797,N_14715,N_14420);
nor UO_1798 (O_1798,N_14393,N_14458);
or UO_1799 (O_1799,N_13549,N_14420);
and UO_1800 (O_1800,N_14445,N_13892);
nand UO_1801 (O_1801,N_14049,N_13530);
nor UO_1802 (O_1802,N_13683,N_13695);
or UO_1803 (O_1803,N_14534,N_13892);
and UO_1804 (O_1804,N_13952,N_14174);
and UO_1805 (O_1805,N_14322,N_13891);
xor UO_1806 (O_1806,N_13833,N_14425);
nand UO_1807 (O_1807,N_14947,N_14652);
or UO_1808 (O_1808,N_13893,N_13933);
or UO_1809 (O_1809,N_14064,N_14896);
xor UO_1810 (O_1810,N_13721,N_14240);
or UO_1811 (O_1811,N_13911,N_14438);
nand UO_1812 (O_1812,N_14568,N_14805);
nor UO_1813 (O_1813,N_14156,N_13630);
and UO_1814 (O_1814,N_14137,N_13774);
nand UO_1815 (O_1815,N_14270,N_14218);
or UO_1816 (O_1816,N_14380,N_14084);
and UO_1817 (O_1817,N_13719,N_13962);
or UO_1818 (O_1818,N_13566,N_14759);
nand UO_1819 (O_1819,N_14334,N_13745);
nand UO_1820 (O_1820,N_14839,N_14522);
and UO_1821 (O_1821,N_14587,N_14349);
nor UO_1822 (O_1822,N_14855,N_14610);
nand UO_1823 (O_1823,N_14377,N_13732);
and UO_1824 (O_1824,N_14253,N_14673);
nor UO_1825 (O_1825,N_14248,N_13732);
nand UO_1826 (O_1826,N_14599,N_13570);
nand UO_1827 (O_1827,N_13746,N_13858);
nand UO_1828 (O_1828,N_14053,N_13774);
nor UO_1829 (O_1829,N_13543,N_14044);
and UO_1830 (O_1830,N_13764,N_14454);
nor UO_1831 (O_1831,N_13666,N_13839);
nor UO_1832 (O_1832,N_14220,N_14660);
nand UO_1833 (O_1833,N_14298,N_14160);
xor UO_1834 (O_1834,N_13969,N_14061);
and UO_1835 (O_1835,N_14452,N_13552);
xor UO_1836 (O_1836,N_14543,N_13871);
xnor UO_1837 (O_1837,N_13926,N_14954);
nand UO_1838 (O_1838,N_14801,N_14783);
nand UO_1839 (O_1839,N_14285,N_13871);
nor UO_1840 (O_1840,N_14059,N_13624);
xor UO_1841 (O_1841,N_13626,N_13684);
or UO_1842 (O_1842,N_14483,N_14153);
and UO_1843 (O_1843,N_14715,N_14668);
xnor UO_1844 (O_1844,N_13943,N_14680);
and UO_1845 (O_1845,N_13831,N_14942);
nor UO_1846 (O_1846,N_14382,N_14683);
and UO_1847 (O_1847,N_14339,N_14531);
nor UO_1848 (O_1848,N_13845,N_14983);
and UO_1849 (O_1849,N_14210,N_14807);
or UO_1850 (O_1850,N_13542,N_14289);
and UO_1851 (O_1851,N_14341,N_14927);
nand UO_1852 (O_1852,N_14255,N_13534);
xor UO_1853 (O_1853,N_14634,N_13738);
and UO_1854 (O_1854,N_13932,N_13690);
or UO_1855 (O_1855,N_13640,N_14417);
or UO_1856 (O_1856,N_13524,N_14649);
and UO_1857 (O_1857,N_14253,N_13560);
nand UO_1858 (O_1858,N_14449,N_13687);
xor UO_1859 (O_1859,N_14424,N_14811);
nand UO_1860 (O_1860,N_14080,N_14881);
or UO_1861 (O_1861,N_14425,N_13650);
or UO_1862 (O_1862,N_13707,N_13897);
and UO_1863 (O_1863,N_14037,N_13547);
xor UO_1864 (O_1864,N_14429,N_13611);
nor UO_1865 (O_1865,N_14599,N_14497);
nor UO_1866 (O_1866,N_13891,N_13539);
nand UO_1867 (O_1867,N_14592,N_14829);
or UO_1868 (O_1868,N_14109,N_14551);
nand UO_1869 (O_1869,N_13727,N_14683);
and UO_1870 (O_1870,N_14515,N_14301);
nor UO_1871 (O_1871,N_13954,N_14648);
or UO_1872 (O_1872,N_14425,N_14261);
nor UO_1873 (O_1873,N_14873,N_14093);
nand UO_1874 (O_1874,N_13799,N_13776);
xnor UO_1875 (O_1875,N_14345,N_14298);
xnor UO_1876 (O_1876,N_14913,N_14475);
nor UO_1877 (O_1877,N_13652,N_14104);
or UO_1878 (O_1878,N_14870,N_14167);
nor UO_1879 (O_1879,N_14305,N_13985);
and UO_1880 (O_1880,N_14081,N_13645);
and UO_1881 (O_1881,N_14697,N_14702);
and UO_1882 (O_1882,N_14711,N_13626);
nand UO_1883 (O_1883,N_14199,N_14907);
xor UO_1884 (O_1884,N_14915,N_13928);
or UO_1885 (O_1885,N_13807,N_14317);
xnor UO_1886 (O_1886,N_14687,N_13716);
or UO_1887 (O_1887,N_13642,N_13934);
or UO_1888 (O_1888,N_14776,N_14479);
nand UO_1889 (O_1889,N_14747,N_13929);
xnor UO_1890 (O_1890,N_13674,N_14413);
or UO_1891 (O_1891,N_14024,N_14027);
nand UO_1892 (O_1892,N_14949,N_13719);
and UO_1893 (O_1893,N_14647,N_13576);
nor UO_1894 (O_1894,N_13815,N_13606);
and UO_1895 (O_1895,N_14527,N_13510);
and UO_1896 (O_1896,N_14266,N_13804);
nand UO_1897 (O_1897,N_14731,N_13876);
or UO_1898 (O_1898,N_13744,N_14427);
xnor UO_1899 (O_1899,N_14318,N_14794);
nand UO_1900 (O_1900,N_14405,N_13824);
or UO_1901 (O_1901,N_14225,N_13986);
or UO_1902 (O_1902,N_14416,N_13952);
or UO_1903 (O_1903,N_13990,N_13615);
and UO_1904 (O_1904,N_14489,N_14928);
nand UO_1905 (O_1905,N_13694,N_14679);
or UO_1906 (O_1906,N_14982,N_13954);
nor UO_1907 (O_1907,N_14156,N_13661);
or UO_1908 (O_1908,N_13834,N_14539);
xnor UO_1909 (O_1909,N_14477,N_14052);
nand UO_1910 (O_1910,N_14463,N_14769);
or UO_1911 (O_1911,N_14453,N_14474);
nand UO_1912 (O_1912,N_14225,N_14166);
and UO_1913 (O_1913,N_14190,N_13707);
or UO_1914 (O_1914,N_13615,N_14762);
or UO_1915 (O_1915,N_13543,N_14973);
xor UO_1916 (O_1916,N_13980,N_13770);
nor UO_1917 (O_1917,N_14004,N_13565);
nor UO_1918 (O_1918,N_14129,N_13852);
or UO_1919 (O_1919,N_14395,N_13577);
nor UO_1920 (O_1920,N_14246,N_14633);
and UO_1921 (O_1921,N_14432,N_14073);
nand UO_1922 (O_1922,N_14652,N_14372);
and UO_1923 (O_1923,N_14552,N_14965);
nand UO_1924 (O_1924,N_14474,N_14729);
xor UO_1925 (O_1925,N_14639,N_14725);
or UO_1926 (O_1926,N_14693,N_14730);
or UO_1927 (O_1927,N_13943,N_14335);
or UO_1928 (O_1928,N_14869,N_13567);
nand UO_1929 (O_1929,N_14563,N_14465);
nand UO_1930 (O_1930,N_14759,N_14277);
nand UO_1931 (O_1931,N_13699,N_14633);
nor UO_1932 (O_1932,N_13648,N_14828);
or UO_1933 (O_1933,N_14050,N_13916);
nand UO_1934 (O_1934,N_14687,N_13813);
and UO_1935 (O_1935,N_13744,N_14240);
nand UO_1936 (O_1936,N_14110,N_13546);
nand UO_1937 (O_1937,N_14949,N_14002);
or UO_1938 (O_1938,N_14612,N_13584);
and UO_1939 (O_1939,N_14566,N_14250);
nor UO_1940 (O_1940,N_14714,N_13873);
nand UO_1941 (O_1941,N_14707,N_13956);
nor UO_1942 (O_1942,N_14901,N_13547);
and UO_1943 (O_1943,N_13646,N_14674);
and UO_1944 (O_1944,N_14855,N_13709);
or UO_1945 (O_1945,N_14860,N_14793);
nor UO_1946 (O_1946,N_14206,N_14126);
nand UO_1947 (O_1947,N_14697,N_14704);
nand UO_1948 (O_1948,N_14787,N_14431);
or UO_1949 (O_1949,N_14361,N_13769);
or UO_1950 (O_1950,N_14824,N_13694);
or UO_1951 (O_1951,N_14965,N_14510);
nor UO_1952 (O_1952,N_13964,N_14831);
nand UO_1953 (O_1953,N_13582,N_14356);
nor UO_1954 (O_1954,N_14860,N_14992);
xnor UO_1955 (O_1955,N_14743,N_13969);
nor UO_1956 (O_1956,N_13766,N_14600);
and UO_1957 (O_1957,N_14594,N_13937);
xor UO_1958 (O_1958,N_14515,N_14761);
nand UO_1959 (O_1959,N_14108,N_13757);
or UO_1960 (O_1960,N_14282,N_14296);
or UO_1961 (O_1961,N_14236,N_14837);
nor UO_1962 (O_1962,N_13815,N_14197);
and UO_1963 (O_1963,N_14965,N_14639);
and UO_1964 (O_1964,N_14984,N_14128);
and UO_1965 (O_1965,N_13845,N_14197);
nand UO_1966 (O_1966,N_13973,N_14301);
or UO_1967 (O_1967,N_14442,N_14103);
or UO_1968 (O_1968,N_14617,N_13872);
or UO_1969 (O_1969,N_14280,N_14539);
and UO_1970 (O_1970,N_14272,N_14344);
nor UO_1971 (O_1971,N_13521,N_14658);
nand UO_1972 (O_1972,N_14387,N_14805);
xor UO_1973 (O_1973,N_14876,N_13986);
xnor UO_1974 (O_1974,N_14634,N_13931);
and UO_1975 (O_1975,N_14691,N_14878);
or UO_1976 (O_1976,N_14825,N_13709);
or UO_1977 (O_1977,N_13963,N_14120);
nand UO_1978 (O_1978,N_14790,N_13577);
and UO_1979 (O_1979,N_13682,N_14189);
nor UO_1980 (O_1980,N_14769,N_13939);
or UO_1981 (O_1981,N_14852,N_14497);
and UO_1982 (O_1982,N_14483,N_14332);
nand UO_1983 (O_1983,N_14884,N_14448);
or UO_1984 (O_1984,N_14096,N_13596);
or UO_1985 (O_1985,N_14080,N_14336);
nor UO_1986 (O_1986,N_14396,N_14291);
nand UO_1987 (O_1987,N_13772,N_14296);
and UO_1988 (O_1988,N_14610,N_13948);
and UO_1989 (O_1989,N_14706,N_14434);
xor UO_1990 (O_1990,N_13910,N_14947);
nor UO_1991 (O_1991,N_14428,N_13608);
nor UO_1992 (O_1992,N_13669,N_13661);
nand UO_1993 (O_1993,N_13569,N_13590);
xnor UO_1994 (O_1994,N_14245,N_13909);
nor UO_1995 (O_1995,N_14580,N_13934);
and UO_1996 (O_1996,N_14114,N_14292);
nand UO_1997 (O_1997,N_14295,N_14042);
or UO_1998 (O_1998,N_14749,N_14525);
xor UO_1999 (O_1999,N_14490,N_14202);
endmodule