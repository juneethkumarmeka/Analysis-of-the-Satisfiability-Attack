module basic_750_5000_1000_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_446,In_76);
nor U1 (N_1,In_80,In_612);
or U2 (N_2,In_509,In_244);
xnor U3 (N_3,In_510,In_77);
and U4 (N_4,In_280,In_196);
and U5 (N_5,In_368,In_684);
or U6 (N_6,In_719,In_473);
or U7 (N_7,In_407,In_350);
nand U8 (N_8,In_456,In_31);
and U9 (N_9,In_655,In_262);
nand U10 (N_10,In_391,In_599);
nand U11 (N_11,In_142,In_463);
nor U12 (N_12,In_543,In_455);
or U13 (N_13,In_98,In_563);
and U14 (N_14,In_21,In_157);
nor U15 (N_15,In_439,In_480);
or U16 (N_16,In_13,In_339);
nand U17 (N_17,In_689,In_188);
or U18 (N_18,In_397,In_377);
nand U19 (N_19,In_56,In_499);
nand U20 (N_20,In_422,In_99);
or U21 (N_21,In_131,In_29);
and U22 (N_22,In_41,In_506);
and U23 (N_23,In_575,In_421);
nand U24 (N_24,In_315,In_481);
nand U25 (N_25,In_235,In_383);
or U26 (N_26,In_395,In_225);
and U27 (N_27,In_534,In_667);
nor U28 (N_28,In_597,In_695);
xnor U29 (N_29,In_322,In_501);
nor U30 (N_30,In_606,In_125);
nand U31 (N_31,In_173,In_554);
nor U32 (N_32,In_55,In_431);
or U33 (N_33,In_347,In_51);
or U34 (N_34,In_603,In_618);
and U35 (N_35,In_406,In_177);
or U36 (N_36,In_284,In_57);
xor U37 (N_37,In_527,In_307);
nor U38 (N_38,In_592,In_148);
nand U39 (N_39,In_78,In_326);
or U40 (N_40,In_290,In_283);
nand U41 (N_41,In_355,In_140);
xnor U42 (N_42,In_102,In_171);
nand U43 (N_43,In_662,In_46);
nor U44 (N_44,In_11,In_664);
nor U45 (N_45,In_726,In_692);
or U46 (N_46,In_268,In_614);
nand U47 (N_47,In_237,In_564);
and U48 (N_48,In_649,In_738);
or U49 (N_49,In_622,In_277);
or U50 (N_50,In_601,In_310);
nand U51 (N_51,In_404,In_303);
or U52 (N_52,In_35,In_149);
nor U53 (N_53,In_258,In_490);
xnor U54 (N_54,In_578,In_112);
and U55 (N_55,In_716,In_454);
nor U56 (N_56,In_351,In_519);
nand U57 (N_57,In_241,In_432);
or U58 (N_58,In_119,In_441);
or U59 (N_59,In_591,In_278);
or U60 (N_60,In_718,In_660);
or U61 (N_61,In_194,In_184);
and U62 (N_62,In_38,In_747);
and U63 (N_63,In_589,In_590);
and U64 (N_64,In_359,In_211);
nand U65 (N_65,In_634,In_478);
and U66 (N_66,In_423,In_84);
and U67 (N_67,In_338,In_321);
xnor U68 (N_68,In_525,In_593);
nor U69 (N_69,In_353,In_114);
nor U70 (N_70,In_661,In_741);
and U71 (N_71,In_174,In_104);
nor U72 (N_72,In_728,In_433);
and U73 (N_73,In_528,In_693);
and U74 (N_74,In_229,In_491);
or U75 (N_75,In_16,In_744);
or U76 (N_76,In_633,In_610);
or U77 (N_77,In_238,In_524);
or U78 (N_78,In_115,In_37);
nand U79 (N_79,In_79,In_546);
xnor U80 (N_80,In_308,In_387);
nor U81 (N_81,In_32,In_122);
nand U82 (N_82,In_95,In_65);
or U83 (N_83,In_420,In_152);
and U84 (N_84,In_495,In_86);
or U85 (N_85,In_652,In_153);
nand U86 (N_86,In_130,In_675);
nor U87 (N_87,In_573,In_743);
or U88 (N_88,In_145,In_568);
xnor U89 (N_89,In_212,In_105);
and U90 (N_90,In_584,In_256);
and U91 (N_91,In_511,In_700);
nor U92 (N_92,In_451,In_430);
and U93 (N_93,In_208,In_87);
nand U94 (N_94,In_317,In_413);
xor U95 (N_95,In_643,In_545);
xnor U96 (N_96,In_602,In_236);
nor U97 (N_97,In_414,In_139);
or U98 (N_98,In_740,In_199);
xor U99 (N_99,In_657,In_269);
nand U100 (N_100,In_20,In_556);
nor U101 (N_101,In_734,In_103);
and U102 (N_102,In_467,In_62);
and U103 (N_103,In_222,In_34);
and U104 (N_104,In_348,In_642);
xnor U105 (N_105,In_267,In_720);
or U106 (N_106,In_617,In_565);
or U107 (N_107,In_129,In_245);
or U108 (N_108,In_386,In_405);
nor U109 (N_109,In_567,In_61);
or U110 (N_110,In_475,In_620);
nand U111 (N_111,In_521,In_52);
and U112 (N_112,In_189,In_448);
or U113 (N_113,In_155,In_717);
and U114 (N_114,In_44,In_66);
and U115 (N_115,In_676,In_198);
nor U116 (N_116,In_619,In_374);
or U117 (N_117,In_558,In_42);
nand U118 (N_118,In_291,In_381);
nor U119 (N_119,In_186,In_214);
and U120 (N_120,In_444,In_605);
nor U121 (N_121,In_6,In_319);
or U122 (N_122,In_513,In_12);
and U123 (N_123,In_557,In_588);
nor U124 (N_124,In_396,In_698);
or U125 (N_125,In_88,In_312);
xor U126 (N_126,In_496,In_365);
and U127 (N_127,In_113,In_489);
nand U128 (N_128,In_637,In_181);
nand U129 (N_129,In_232,In_197);
nor U130 (N_130,In_272,In_116);
nor U131 (N_131,In_394,In_179);
nand U132 (N_132,In_43,In_626);
nand U133 (N_133,In_725,In_533);
or U134 (N_134,In_638,In_261);
and U135 (N_135,In_274,In_449);
nor U136 (N_136,In_111,In_409);
or U137 (N_137,In_343,In_378);
nor U138 (N_138,In_349,In_702);
xor U139 (N_139,In_639,In_295);
or U140 (N_140,In_629,In_540);
or U141 (N_141,In_252,In_459);
or U142 (N_142,In_26,In_17);
nand U143 (N_143,In_608,In_399);
and U144 (N_144,In_561,In_324);
and U145 (N_145,In_10,In_100);
nor U146 (N_146,In_276,In_221);
and U147 (N_147,In_625,In_271);
xor U148 (N_148,In_93,In_254);
or U149 (N_149,In_537,In_223);
nand U150 (N_150,In_745,In_306);
xor U151 (N_151,In_215,In_328);
nor U152 (N_152,In_685,In_60);
nor U153 (N_153,In_83,In_724);
xor U154 (N_154,In_668,In_220);
or U155 (N_155,In_192,In_504);
or U156 (N_156,In_33,In_231);
and U157 (N_157,In_243,In_183);
and U158 (N_158,In_392,In_275);
nor U159 (N_159,In_364,In_666);
nor U160 (N_160,In_40,In_7);
nor U161 (N_161,In_550,In_90);
xnor U162 (N_162,In_436,In_299);
nand U163 (N_163,In_671,In_327);
or U164 (N_164,In_48,In_216);
nor U165 (N_165,In_24,In_503);
nand U166 (N_166,In_346,In_279);
nor U167 (N_167,In_107,In_358);
xor U168 (N_168,In_170,In_27);
nand U169 (N_169,In_703,In_551);
and U170 (N_170,In_670,In_710);
and U171 (N_171,In_401,In_89);
or U172 (N_172,In_623,In_193);
nor U173 (N_173,In_128,In_403);
or U174 (N_174,In_426,In_70);
or U175 (N_175,In_304,In_721);
and U176 (N_176,In_389,In_722);
xor U177 (N_177,In_538,In_30);
nand U178 (N_178,In_361,In_577);
or U179 (N_179,In_182,In_539);
and U180 (N_180,In_371,In_445);
nor U181 (N_181,In_167,In_560);
nand U182 (N_182,In_472,In_418);
nor U183 (N_183,In_143,In_410);
nor U184 (N_184,In_690,In_663);
nor U185 (N_185,In_302,In_206);
or U186 (N_186,In_484,In_479);
nor U187 (N_187,In_621,In_323);
nor U188 (N_188,In_305,In_627);
and U189 (N_189,In_201,In_651);
nor U190 (N_190,In_428,In_169);
xnor U191 (N_191,In_466,In_69);
xnor U192 (N_192,In_226,In_332);
and U193 (N_193,In_178,In_101);
nand U194 (N_194,In_248,In_260);
and U195 (N_195,In_645,In_136);
or U196 (N_196,In_94,In_207);
nor U197 (N_197,In_462,In_458);
nor U198 (N_198,In_541,In_314);
nor U199 (N_199,In_1,In_320);
xnor U200 (N_200,In_486,In_334);
and U201 (N_201,In_450,In_265);
nand U202 (N_202,In_150,In_544);
nor U203 (N_203,In_356,In_416);
nor U204 (N_204,In_75,In_542);
or U205 (N_205,In_301,In_58);
or U206 (N_206,In_483,In_240);
and U207 (N_207,In_616,In_408);
or U208 (N_208,In_553,In_108);
nand U209 (N_209,In_357,In_659);
or U210 (N_210,In_636,In_270);
and U211 (N_211,In_714,In_293);
nor U212 (N_212,In_576,In_735);
or U213 (N_213,In_678,In_653);
nor U214 (N_214,In_109,In_205);
nand U215 (N_215,In_646,In_8);
or U216 (N_216,In_388,In_202);
nand U217 (N_217,In_172,In_613);
or U218 (N_218,In_574,In_712);
or U219 (N_219,In_286,In_36);
nor U220 (N_220,In_727,In_134);
nand U221 (N_221,In_273,In_673);
and U222 (N_222,In_373,In_683);
nand U223 (N_223,In_195,In_729);
xnor U224 (N_224,In_746,In_672);
and U225 (N_225,In_434,In_22);
nand U226 (N_226,In_300,In_96);
nor U227 (N_227,In_631,In_23);
nand U228 (N_228,In_352,In_2);
and U229 (N_229,In_390,In_159);
xnor U230 (N_230,In_289,In_429);
nor U231 (N_231,In_19,In_340);
nand U232 (N_232,In_674,In_309);
nor U233 (N_233,In_0,In_367);
nand U234 (N_234,In_505,In_705);
nand U235 (N_235,In_635,In_609);
nor U236 (N_236,In_200,In_247);
nand U237 (N_237,In_447,In_120);
and U238 (N_238,In_526,In_18);
or U239 (N_239,In_28,In_748);
or U240 (N_240,In_679,In_572);
nand U241 (N_241,In_411,In_742);
and U242 (N_242,In_213,In_438);
nor U243 (N_243,In_331,In_158);
and U244 (N_244,In_342,In_681);
nor U245 (N_245,In_474,In_9);
nor U246 (N_246,In_123,In_264);
nor U247 (N_247,In_682,In_72);
nor U248 (N_248,In_644,In_117);
nand U249 (N_249,In_250,In_4);
and U250 (N_250,In_384,In_126);
or U251 (N_251,In_691,In_464);
and U252 (N_252,In_677,In_628);
or U253 (N_253,In_485,In_156);
nor U254 (N_254,In_147,In_380);
and U255 (N_255,In_562,In_417);
nor U256 (N_256,In_571,In_106);
and U257 (N_257,In_427,In_335);
nor U258 (N_258,In_594,In_209);
and U259 (N_259,In_369,In_731);
xor U260 (N_260,In_512,In_285);
nand U261 (N_261,In_641,In_366);
nand U262 (N_262,In_482,In_569);
nand U263 (N_263,In_730,In_507);
and U264 (N_264,In_375,In_15);
nand U265 (N_265,In_598,In_529);
nand U266 (N_266,In_687,In_354);
nand U267 (N_267,In_230,In_749);
or U268 (N_268,In_453,In_522);
xor U269 (N_269,In_282,In_360);
or U270 (N_270,In_471,In_686);
nand U271 (N_271,In_63,In_469);
nor U272 (N_272,In_607,In_688);
nand U273 (N_273,In_732,In_502);
or U274 (N_274,In_135,In_137);
and U275 (N_275,In_736,In_337);
nor U276 (N_276,In_118,In_465);
and U277 (N_277,In_74,In_85);
nand U278 (N_278,In_615,In_457);
and U279 (N_279,In_523,In_699);
or U280 (N_280,In_313,In_316);
nor U281 (N_281,In_548,In_73);
or U282 (N_282,In_493,In_253);
nand U283 (N_283,In_624,In_582);
nand U284 (N_284,In_739,In_233);
or U285 (N_285,In_92,In_723);
nor U286 (N_286,In_587,In_376);
nor U287 (N_287,In_25,In_440);
nor U288 (N_288,In_133,In_711);
or U289 (N_289,In_210,In_494);
and U290 (N_290,In_124,In_266);
nor U291 (N_291,In_217,In_552);
or U292 (N_292,In_547,In_345);
and U293 (N_293,In_706,In_497);
nand U294 (N_294,In_249,In_654);
or U295 (N_295,In_701,In_650);
nor U296 (N_296,In_658,In_400);
nor U297 (N_297,In_532,In_680);
nor U298 (N_298,In_175,In_185);
or U299 (N_299,In_168,In_97);
nor U300 (N_300,In_53,In_425);
or U301 (N_301,In_251,In_508);
nand U302 (N_302,In_536,In_604);
nand U303 (N_303,In_515,In_39);
nor U304 (N_304,In_516,In_498);
nand U305 (N_305,In_336,In_398);
nor U306 (N_306,In_733,In_443);
nor U307 (N_307,In_127,In_500);
xor U308 (N_308,In_632,In_470);
nand U309 (N_309,In_227,In_435);
and U310 (N_310,In_535,In_224);
and U311 (N_311,In_370,In_234);
nand U312 (N_312,In_330,In_585);
or U313 (N_313,In_419,In_296);
or U314 (N_314,In_242,In_715);
xor U315 (N_315,In_294,In_492);
nand U316 (N_316,In_518,In_611);
xor U317 (N_317,In_586,In_549);
or U318 (N_318,In_514,In_218);
or U319 (N_319,In_737,In_144);
xnor U320 (N_320,In_697,In_530);
nand U321 (N_321,In_154,In_596);
nand U322 (N_322,In_110,In_67);
nor U323 (N_323,In_559,In_442);
and U324 (N_324,In_713,In_176);
or U325 (N_325,In_50,In_257);
and U326 (N_326,In_708,In_341);
and U327 (N_327,In_583,In_520);
or U328 (N_328,In_59,In_311);
nand U329 (N_329,In_477,In_160);
and U330 (N_330,In_630,In_318);
xor U331 (N_331,In_298,In_647);
nor U332 (N_332,In_68,In_146);
or U333 (N_333,In_49,In_191);
xor U334 (N_334,In_372,In_344);
and U335 (N_335,In_91,In_468);
nand U336 (N_336,In_228,In_437);
xor U337 (N_337,In_424,In_166);
nor U338 (N_338,In_694,In_488);
nor U339 (N_339,In_190,In_476);
and U340 (N_340,In_709,In_385);
or U341 (N_341,In_333,In_600);
nor U342 (N_342,In_180,In_5);
or U343 (N_343,In_580,In_460);
nand U344 (N_344,In_555,In_292);
nor U345 (N_345,In_203,In_161);
xor U346 (N_346,In_415,In_204);
xor U347 (N_347,In_696,In_121);
and U348 (N_348,In_665,In_581);
or U349 (N_349,In_393,In_141);
and U350 (N_350,In_412,In_640);
nor U351 (N_351,In_82,In_255);
nor U352 (N_352,In_566,In_362);
nor U353 (N_353,In_281,In_138);
and U354 (N_354,In_297,In_595);
or U355 (N_355,In_263,In_163);
and U356 (N_356,In_151,In_579);
nand U357 (N_357,In_487,In_402);
nand U358 (N_358,In_239,In_81);
and U359 (N_359,In_162,In_246);
or U360 (N_360,In_219,In_45);
and U361 (N_361,In_187,In_707);
and U362 (N_362,In_164,In_656);
nor U363 (N_363,In_288,In_54);
nand U364 (N_364,In_3,In_132);
nand U365 (N_365,In_64,In_329);
nor U366 (N_366,In_363,In_382);
nand U367 (N_367,In_517,In_165);
and U368 (N_368,In_669,In_704);
nor U369 (N_369,In_570,In_531);
nor U370 (N_370,In_47,In_379);
and U371 (N_371,In_452,In_648);
nand U372 (N_372,In_14,In_461);
and U373 (N_373,In_71,In_325);
nand U374 (N_374,In_259,In_287);
and U375 (N_375,In_357,In_419);
and U376 (N_376,In_482,In_395);
and U377 (N_377,In_632,In_180);
and U378 (N_378,In_515,In_354);
nor U379 (N_379,In_567,In_204);
xor U380 (N_380,In_586,In_494);
nor U381 (N_381,In_25,In_281);
or U382 (N_382,In_37,In_363);
or U383 (N_383,In_17,In_285);
and U384 (N_384,In_729,In_715);
and U385 (N_385,In_501,In_675);
and U386 (N_386,In_599,In_2);
nand U387 (N_387,In_249,In_286);
nand U388 (N_388,In_186,In_85);
xnor U389 (N_389,In_53,In_738);
nor U390 (N_390,In_739,In_497);
xor U391 (N_391,In_513,In_191);
and U392 (N_392,In_744,In_562);
and U393 (N_393,In_10,In_225);
or U394 (N_394,In_505,In_598);
nor U395 (N_395,In_302,In_151);
and U396 (N_396,In_281,In_374);
xor U397 (N_397,In_328,In_618);
and U398 (N_398,In_605,In_45);
nor U399 (N_399,In_9,In_180);
or U400 (N_400,In_191,In_729);
or U401 (N_401,In_411,In_403);
nand U402 (N_402,In_108,In_90);
nor U403 (N_403,In_235,In_641);
nor U404 (N_404,In_337,In_399);
or U405 (N_405,In_138,In_696);
nor U406 (N_406,In_664,In_259);
or U407 (N_407,In_338,In_152);
xnor U408 (N_408,In_634,In_34);
nor U409 (N_409,In_622,In_134);
nand U410 (N_410,In_512,In_17);
or U411 (N_411,In_661,In_433);
or U412 (N_412,In_652,In_741);
nor U413 (N_413,In_654,In_691);
nor U414 (N_414,In_154,In_466);
or U415 (N_415,In_620,In_698);
nand U416 (N_416,In_255,In_4);
nand U417 (N_417,In_302,In_286);
xor U418 (N_418,In_416,In_365);
nand U419 (N_419,In_450,In_494);
and U420 (N_420,In_369,In_255);
nand U421 (N_421,In_505,In_434);
nor U422 (N_422,In_614,In_470);
or U423 (N_423,In_22,In_593);
or U424 (N_424,In_603,In_328);
xor U425 (N_425,In_658,In_403);
nand U426 (N_426,In_490,In_499);
nand U427 (N_427,In_320,In_293);
and U428 (N_428,In_112,In_388);
nor U429 (N_429,In_643,In_629);
nand U430 (N_430,In_620,In_520);
nand U431 (N_431,In_74,In_24);
nor U432 (N_432,In_110,In_631);
nor U433 (N_433,In_26,In_330);
or U434 (N_434,In_82,In_622);
nand U435 (N_435,In_729,In_182);
nor U436 (N_436,In_344,In_233);
or U437 (N_437,In_164,In_612);
nor U438 (N_438,In_181,In_258);
xor U439 (N_439,In_133,In_681);
and U440 (N_440,In_209,In_723);
or U441 (N_441,In_221,In_161);
or U442 (N_442,In_566,In_28);
nand U443 (N_443,In_123,In_544);
nand U444 (N_444,In_246,In_31);
nor U445 (N_445,In_517,In_140);
or U446 (N_446,In_273,In_113);
or U447 (N_447,In_323,In_382);
xor U448 (N_448,In_292,In_631);
nor U449 (N_449,In_596,In_607);
nand U450 (N_450,In_708,In_643);
or U451 (N_451,In_220,In_257);
nor U452 (N_452,In_146,In_634);
nor U453 (N_453,In_588,In_630);
or U454 (N_454,In_190,In_523);
or U455 (N_455,In_398,In_558);
xor U456 (N_456,In_259,In_728);
nand U457 (N_457,In_559,In_353);
and U458 (N_458,In_737,In_91);
nor U459 (N_459,In_4,In_67);
nand U460 (N_460,In_312,In_637);
and U461 (N_461,In_526,In_626);
or U462 (N_462,In_704,In_515);
nand U463 (N_463,In_664,In_573);
nor U464 (N_464,In_109,In_670);
nand U465 (N_465,In_733,In_442);
nand U466 (N_466,In_19,In_465);
and U467 (N_467,In_742,In_437);
nor U468 (N_468,In_549,In_651);
or U469 (N_469,In_376,In_433);
nand U470 (N_470,In_431,In_179);
and U471 (N_471,In_331,In_672);
nand U472 (N_472,In_466,In_736);
nor U473 (N_473,In_466,In_512);
or U474 (N_474,In_42,In_463);
nor U475 (N_475,In_231,In_482);
or U476 (N_476,In_138,In_279);
nor U477 (N_477,In_376,In_21);
nor U478 (N_478,In_653,In_8);
nand U479 (N_479,In_683,In_161);
or U480 (N_480,In_110,In_138);
nor U481 (N_481,In_698,In_741);
nand U482 (N_482,In_114,In_611);
nand U483 (N_483,In_466,In_302);
or U484 (N_484,In_85,In_306);
nand U485 (N_485,In_173,In_194);
xor U486 (N_486,In_57,In_11);
xnor U487 (N_487,In_652,In_228);
and U488 (N_488,In_648,In_626);
and U489 (N_489,In_661,In_303);
or U490 (N_490,In_649,In_87);
or U491 (N_491,In_327,In_102);
nor U492 (N_492,In_429,In_362);
or U493 (N_493,In_188,In_60);
xor U494 (N_494,In_466,In_172);
nor U495 (N_495,In_708,In_244);
xor U496 (N_496,In_85,In_420);
and U497 (N_497,In_633,In_552);
nor U498 (N_498,In_693,In_74);
nand U499 (N_499,In_431,In_502);
or U500 (N_500,In_207,In_4);
xor U501 (N_501,In_491,In_353);
or U502 (N_502,In_465,In_59);
nor U503 (N_503,In_713,In_282);
and U504 (N_504,In_99,In_500);
or U505 (N_505,In_472,In_387);
and U506 (N_506,In_237,In_480);
or U507 (N_507,In_647,In_498);
and U508 (N_508,In_721,In_226);
and U509 (N_509,In_655,In_511);
nand U510 (N_510,In_141,In_544);
and U511 (N_511,In_303,In_451);
or U512 (N_512,In_354,In_210);
nand U513 (N_513,In_286,In_301);
or U514 (N_514,In_626,In_308);
and U515 (N_515,In_468,In_194);
or U516 (N_516,In_329,In_362);
nand U517 (N_517,In_0,In_607);
xnor U518 (N_518,In_426,In_644);
and U519 (N_519,In_151,In_504);
nand U520 (N_520,In_406,In_196);
and U521 (N_521,In_569,In_285);
xnor U522 (N_522,In_682,In_235);
or U523 (N_523,In_709,In_212);
xnor U524 (N_524,In_717,In_606);
or U525 (N_525,In_710,In_142);
or U526 (N_526,In_19,In_717);
nor U527 (N_527,In_726,In_1);
nor U528 (N_528,In_584,In_599);
or U529 (N_529,In_530,In_38);
xnor U530 (N_530,In_248,In_689);
nand U531 (N_531,In_519,In_672);
nand U532 (N_532,In_568,In_99);
and U533 (N_533,In_604,In_164);
nor U534 (N_534,In_612,In_236);
nor U535 (N_535,In_484,In_148);
nand U536 (N_536,In_392,In_183);
or U537 (N_537,In_136,In_102);
nand U538 (N_538,In_619,In_643);
nand U539 (N_539,In_423,In_42);
or U540 (N_540,In_618,In_191);
nor U541 (N_541,In_137,In_46);
and U542 (N_542,In_415,In_583);
nand U543 (N_543,In_426,In_442);
xor U544 (N_544,In_51,In_138);
and U545 (N_545,In_470,In_729);
or U546 (N_546,In_374,In_420);
or U547 (N_547,In_318,In_138);
nand U548 (N_548,In_16,In_634);
and U549 (N_549,In_623,In_584);
or U550 (N_550,In_178,In_471);
nand U551 (N_551,In_254,In_147);
nor U552 (N_552,In_316,In_651);
and U553 (N_553,In_694,In_593);
or U554 (N_554,In_353,In_99);
and U555 (N_555,In_7,In_556);
nor U556 (N_556,In_701,In_735);
nand U557 (N_557,In_72,In_591);
nand U558 (N_558,In_31,In_744);
nor U559 (N_559,In_705,In_151);
nor U560 (N_560,In_138,In_167);
nor U561 (N_561,In_132,In_138);
nor U562 (N_562,In_544,In_639);
or U563 (N_563,In_84,In_596);
or U564 (N_564,In_199,In_235);
and U565 (N_565,In_620,In_444);
and U566 (N_566,In_660,In_203);
xnor U567 (N_567,In_50,In_488);
nand U568 (N_568,In_65,In_477);
nand U569 (N_569,In_266,In_262);
or U570 (N_570,In_618,In_737);
and U571 (N_571,In_72,In_242);
or U572 (N_572,In_98,In_194);
and U573 (N_573,In_168,In_3);
nand U574 (N_574,In_570,In_431);
and U575 (N_575,In_659,In_77);
nor U576 (N_576,In_697,In_484);
nand U577 (N_577,In_478,In_620);
nand U578 (N_578,In_436,In_729);
or U579 (N_579,In_742,In_699);
and U580 (N_580,In_742,In_102);
nand U581 (N_581,In_611,In_63);
nor U582 (N_582,In_192,In_275);
xnor U583 (N_583,In_103,In_0);
and U584 (N_584,In_382,In_259);
nor U585 (N_585,In_714,In_145);
or U586 (N_586,In_31,In_352);
or U587 (N_587,In_608,In_406);
nand U588 (N_588,In_55,In_619);
and U589 (N_589,In_742,In_199);
or U590 (N_590,In_589,In_554);
nand U591 (N_591,In_575,In_734);
xor U592 (N_592,In_103,In_49);
nand U593 (N_593,In_353,In_378);
nand U594 (N_594,In_514,In_528);
xnor U595 (N_595,In_719,In_397);
or U596 (N_596,In_216,In_480);
nor U597 (N_597,In_684,In_294);
nand U598 (N_598,In_269,In_501);
nor U599 (N_599,In_356,In_681);
nor U600 (N_600,In_585,In_716);
nand U601 (N_601,In_322,In_621);
nand U602 (N_602,In_405,In_57);
nor U603 (N_603,In_164,In_667);
and U604 (N_604,In_485,In_95);
and U605 (N_605,In_689,In_622);
and U606 (N_606,In_149,In_38);
and U607 (N_607,In_369,In_22);
or U608 (N_608,In_364,In_343);
nand U609 (N_609,In_729,In_280);
nand U610 (N_610,In_132,In_306);
or U611 (N_611,In_455,In_432);
and U612 (N_612,In_532,In_629);
nand U613 (N_613,In_256,In_253);
nor U614 (N_614,In_456,In_718);
nand U615 (N_615,In_648,In_481);
nand U616 (N_616,In_268,In_49);
xor U617 (N_617,In_93,In_200);
xor U618 (N_618,In_613,In_65);
or U619 (N_619,In_471,In_509);
or U620 (N_620,In_82,In_661);
nand U621 (N_621,In_5,In_62);
nand U622 (N_622,In_146,In_749);
nand U623 (N_623,In_523,In_522);
nor U624 (N_624,In_504,In_325);
nor U625 (N_625,In_696,In_332);
or U626 (N_626,In_708,In_375);
or U627 (N_627,In_672,In_201);
and U628 (N_628,In_79,In_19);
nor U629 (N_629,In_567,In_333);
nor U630 (N_630,In_631,In_597);
and U631 (N_631,In_542,In_561);
and U632 (N_632,In_617,In_430);
nor U633 (N_633,In_221,In_325);
nor U634 (N_634,In_507,In_617);
or U635 (N_635,In_164,In_615);
or U636 (N_636,In_380,In_737);
and U637 (N_637,In_119,In_158);
nor U638 (N_638,In_628,In_16);
nand U639 (N_639,In_281,In_346);
and U640 (N_640,In_252,In_369);
xor U641 (N_641,In_335,In_212);
nand U642 (N_642,In_308,In_613);
nand U643 (N_643,In_53,In_445);
nor U644 (N_644,In_385,In_346);
and U645 (N_645,In_39,In_706);
nand U646 (N_646,In_688,In_53);
or U647 (N_647,In_706,In_682);
or U648 (N_648,In_463,In_597);
xor U649 (N_649,In_582,In_441);
or U650 (N_650,In_365,In_574);
nor U651 (N_651,In_729,In_555);
and U652 (N_652,In_46,In_428);
nand U653 (N_653,In_738,In_692);
or U654 (N_654,In_649,In_52);
nor U655 (N_655,In_123,In_607);
and U656 (N_656,In_424,In_227);
xor U657 (N_657,In_367,In_118);
and U658 (N_658,In_106,In_369);
nand U659 (N_659,In_211,In_113);
xnor U660 (N_660,In_138,In_418);
nand U661 (N_661,In_748,In_691);
nor U662 (N_662,In_160,In_115);
or U663 (N_663,In_168,In_69);
nand U664 (N_664,In_293,In_524);
xor U665 (N_665,In_285,In_428);
nor U666 (N_666,In_312,In_17);
nand U667 (N_667,In_80,In_357);
or U668 (N_668,In_494,In_143);
and U669 (N_669,In_370,In_406);
nand U670 (N_670,In_79,In_330);
nor U671 (N_671,In_434,In_77);
and U672 (N_672,In_113,In_213);
nand U673 (N_673,In_199,In_317);
xor U674 (N_674,In_157,In_332);
nand U675 (N_675,In_361,In_94);
or U676 (N_676,In_194,In_604);
or U677 (N_677,In_719,In_582);
nand U678 (N_678,In_13,In_725);
and U679 (N_679,In_278,In_615);
nand U680 (N_680,In_692,In_274);
and U681 (N_681,In_395,In_559);
and U682 (N_682,In_718,In_484);
nand U683 (N_683,In_568,In_57);
nand U684 (N_684,In_134,In_490);
and U685 (N_685,In_73,In_174);
and U686 (N_686,In_498,In_511);
and U687 (N_687,In_167,In_706);
nand U688 (N_688,In_391,In_473);
nand U689 (N_689,In_404,In_233);
and U690 (N_690,In_300,In_158);
or U691 (N_691,In_316,In_274);
nand U692 (N_692,In_174,In_128);
and U693 (N_693,In_558,In_397);
nor U694 (N_694,In_732,In_578);
xor U695 (N_695,In_522,In_337);
and U696 (N_696,In_640,In_405);
nand U697 (N_697,In_28,In_493);
nor U698 (N_698,In_343,In_353);
nor U699 (N_699,In_444,In_295);
xor U700 (N_700,In_662,In_282);
nand U701 (N_701,In_666,In_674);
or U702 (N_702,In_155,In_213);
nand U703 (N_703,In_312,In_675);
and U704 (N_704,In_605,In_160);
nand U705 (N_705,In_574,In_727);
or U706 (N_706,In_261,In_78);
nand U707 (N_707,In_447,In_607);
nand U708 (N_708,In_640,In_316);
nand U709 (N_709,In_279,In_2);
nand U710 (N_710,In_503,In_593);
xnor U711 (N_711,In_11,In_175);
xnor U712 (N_712,In_207,In_428);
nor U713 (N_713,In_366,In_355);
or U714 (N_714,In_192,In_263);
and U715 (N_715,In_176,In_546);
or U716 (N_716,In_55,In_555);
xor U717 (N_717,In_277,In_109);
and U718 (N_718,In_637,In_378);
and U719 (N_719,In_256,In_721);
and U720 (N_720,In_11,In_319);
and U721 (N_721,In_76,In_572);
or U722 (N_722,In_298,In_27);
nor U723 (N_723,In_245,In_337);
xor U724 (N_724,In_724,In_492);
or U725 (N_725,In_635,In_179);
nand U726 (N_726,In_175,In_349);
nor U727 (N_727,In_354,In_455);
or U728 (N_728,In_642,In_609);
nand U729 (N_729,In_733,In_521);
or U730 (N_730,In_127,In_268);
xor U731 (N_731,In_245,In_554);
nor U732 (N_732,In_446,In_110);
nand U733 (N_733,In_426,In_668);
and U734 (N_734,In_5,In_232);
xnor U735 (N_735,In_455,In_318);
nor U736 (N_736,In_586,In_246);
nand U737 (N_737,In_89,In_462);
or U738 (N_738,In_237,In_464);
xnor U739 (N_739,In_280,In_592);
nor U740 (N_740,In_321,In_97);
or U741 (N_741,In_259,In_634);
and U742 (N_742,In_59,In_234);
nand U743 (N_743,In_0,In_88);
nor U744 (N_744,In_362,In_116);
and U745 (N_745,In_747,In_579);
or U746 (N_746,In_683,In_206);
nor U747 (N_747,In_496,In_313);
and U748 (N_748,In_68,In_731);
or U749 (N_749,In_713,In_493);
and U750 (N_750,In_685,In_707);
nor U751 (N_751,In_577,In_206);
or U752 (N_752,In_659,In_514);
nand U753 (N_753,In_662,In_146);
nor U754 (N_754,In_303,In_706);
nand U755 (N_755,In_94,In_623);
and U756 (N_756,In_357,In_638);
nor U757 (N_757,In_115,In_208);
nand U758 (N_758,In_157,In_435);
xnor U759 (N_759,In_640,In_686);
or U760 (N_760,In_551,In_699);
nand U761 (N_761,In_414,In_440);
and U762 (N_762,In_318,In_215);
nor U763 (N_763,In_548,In_495);
nor U764 (N_764,In_209,In_155);
and U765 (N_765,In_272,In_423);
nor U766 (N_766,In_736,In_138);
and U767 (N_767,In_745,In_402);
and U768 (N_768,In_547,In_62);
and U769 (N_769,In_654,In_392);
nor U770 (N_770,In_552,In_410);
and U771 (N_771,In_150,In_129);
or U772 (N_772,In_714,In_579);
nor U773 (N_773,In_156,In_716);
and U774 (N_774,In_509,In_548);
nand U775 (N_775,In_249,In_495);
or U776 (N_776,In_194,In_615);
or U777 (N_777,In_435,In_444);
nand U778 (N_778,In_696,In_711);
and U779 (N_779,In_532,In_481);
nor U780 (N_780,In_652,In_698);
and U781 (N_781,In_556,In_386);
or U782 (N_782,In_284,In_268);
or U783 (N_783,In_510,In_560);
or U784 (N_784,In_320,In_362);
nand U785 (N_785,In_654,In_69);
nor U786 (N_786,In_715,In_480);
and U787 (N_787,In_569,In_462);
or U788 (N_788,In_28,In_258);
nand U789 (N_789,In_684,In_273);
or U790 (N_790,In_511,In_237);
nand U791 (N_791,In_181,In_427);
nor U792 (N_792,In_243,In_169);
or U793 (N_793,In_637,In_537);
nand U794 (N_794,In_184,In_607);
and U795 (N_795,In_692,In_691);
nor U796 (N_796,In_28,In_55);
and U797 (N_797,In_112,In_285);
nor U798 (N_798,In_454,In_695);
nand U799 (N_799,In_197,In_352);
nor U800 (N_800,In_435,In_272);
nor U801 (N_801,In_632,In_641);
nand U802 (N_802,In_289,In_242);
xor U803 (N_803,In_367,In_263);
xor U804 (N_804,In_466,In_147);
nor U805 (N_805,In_727,In_639);
or U806 (N_806,In_168,In_717);
nand U807 (N_807,In_615,In_508);
xnor U808 (N_808,In_649,In_748);
or U809 (N_809,In_682,In_189);
and U810 (N_810,In_493,In_298);
xnor U811 (N_811,In_170,In_597);
and U812 (N_812,In_12,In_537);
nor U813 (N_813,In_541,In_646);
and U814 (N_814,In_674,In_420);
nor U815 (N_815,In_700,In_283);
and U816 (N_816,In_321,In_719);
and U817 (N_817,In_552,In_86);
or U818 (N_818,In_15,In_32);
or U819 (N_819,In_57,In_490);
or U820 (N_820,In_523,In_222);
and U821 (N_821,In_574,In_190);
and U822 (N_822,In_604,In_378);
and U823 (N_823,In_517,In_412);
nand U824 (N_824,In_250,In_489);
nor U825 (N_825,In_477,In_558);
and U826 (N_826,In_353,In_500);
and U827 (N_827,In_329,In_270);
nor U828 (N_828,In_671,In_18);
or U829 (N_829,In_167,In_134);
xor U830 (N_830,In_581,In_745);
nor U831 (N_831,In_677,In_247);
nor U832 (N_832,In_361,In_529);
nand U833 (N_833,In_531,In_642);
and U834 (N_834,In_541,In_56);
nor U835 (N_835,In_238,In_102);
or U836 (N_836,In_272,In_649);
nor U837 (N_837,In_142,In_459);
or U838 (N_838,In_688,In_576);
and U839 (N_839,In_726,In_351);
and U840 (N_840,In_149,In_295);
nand U841 (N_841,In_118,In_46);
nor U842 (N_842,In_509,In_39);
xnor U843 (N_843,In_648,In_374);
and U844 (N_844,In_299,In_438);
or U845 (N_845,In_708,In_77);
nor U846 (N_846,In_144,In_178);
nand U847 (N_847,In_204,In_321);
or U848 (N_848,In_310,In_670);
nand U849 (N_849,In_502,In_398);
nand U850 (N_850,In_340,In_667);
or U851 (N_851,In_458,In_343);
or U852 (N_852,In_112,In_49);
or U853 (N_853,In_255,In_113);
nor U854 (N_854,In_721,In_224);
nand U855 (N_855,In_52,In_730);
nand U856 (N_856,In_409,In_119);
nand U857 (N_857,In_692,In_514);
and U858 (N_858,In_651,In_605);
nor U859 (N_859,In_503,In_92);
or U860 (N_860,In_749,In_2);
or U861 (N_861,In_331,In_646);
xor U862 (N_862,In_271,In_370);
nor U863 (N_863,In_682,In_707);
or U864 (N_864,In_682,In_83);
and U865 (N_865,In_248,In_658);
and U866 (N_866,In_352,In_457);
and U867 (N_867,In_140,In_555);
nor U868 (N_868,In_530,In_445);
xnor U869 (N_869,In_651,In_664);
nand U870 (N_870,In_373,In_137);
or U871 (N_871,In_41,In_1);
and U872 (N_872,In_576,In_640);
nor U873 (N_873,In_291,In_571);
nor U874 (N_874,In_71,In_464);
or U875 (N_875,In_683,In_185);
xnor U876 (N_876,In_292,In_710);
or U877 (N_877,In_298,In_484);
or U878 (N_878,In_228,In_425);
nor U879 (N_879,In_209,In_409);
and U880 (N_880,In_632,In_573);
nand U881 (N_881,In_718,In_317);
nand U882 (N_882,In_677,In_687);
xor U883 (N_883,In_482,In_366);
nor U884 (N_884,In_555,In_547);
and U885 (N_885,In_567,In_622);
nor U886 (N_886,In_265,In_602);
or U887 (N_887,In_314,In_476);
and U888 (N_888,In_624,In_238);
and U889 (N_889,In_330,In_356);
nor U890 (N_890,In_401,In_369);
or U891 (N_891,In_194,In_346);
xor U892 (N_892,In_408,In_600);
nor U893 (N_893,In_57,In_91);
nor U894 (N_894,In_589,In_259);
or U895 (N_895,In_65,In_716);
nand U896 (N_896,In_379,In_281);
and U897 (N_897,In_410,In_492);
or U898 (N_898,In_652,In_3);
or U899 (N_899,In_717,In_306);
nand U900 (N_900,In_194,In_160);
or U901 (N_901,In_87,In_150);
and U902 (N_902,In_154,In_481);
nor U903 (N_903,In_267,In_548);
or U904 (N_904,In_528,In_122);
nor U905 (N_905,In_349,In_345);
or U906 (N_906,In_598,In_560);
nand U907 (N_907,In_499,In_467);
nor U908 (N_908,In_89,In_147);
or U909 (N_909,In_369,In_344);
or U910 (N_910,In_637,In_141);
nand U911 (N_911,In_639,In_623);
and U912 (N_912,In_150,In_185);
or U913 (N_913,In_294,In_562);
or U914 (N_914,In_398,In_266);
and U915 (N_915,In_293,In_384);
nand U916 (N_916,In_72,In_523);
or U917 (N_917,In_231,In_81);
nand U918 (N_918,In_23,In_285);
and U919 (N_919,In_96,In_731);
or U920 (N_920,In_370,In_229);
and U921 (N_921,In_428,In_59);
or U922 (N_922,In_143,In_681);
xor U923 (N_923,In_515,In_386);
or U924 (N_924,In_653,In_394);
and U925 (N_925,In_376,In_693);
nand U926 (N_926,In_180,In_449);
and U927 (N_927,In_268,In_575);
nand U928 (N_928,In_371,In_238);
nor U929 (N_929,In_479,In_745);
or U930 (N_930,In_41,In_644);
and U931 (N_931,In_179,In_138);
nand U932 (N_932,In_439,In_190);
nor U933 (N_933,In_681,In_195);
and U934 (N_934,In_259,In_192);
nand U935 (N_935,In_604,In_558);
nor U936 (N_936,In_590,In_523);
and U937 (N_937,In_384,In_52);
or U938 (N_938,In_517,In_102);
and U939 (N_939,In_102,In_521);
and U940 (N_940,In_582,In_383);
and U941 (N_941,In_231,In_712);
nor U942 (N_942,In_51,In_317);
and U943 (N_943,In_406,In_538);
and U944 (N_944,In_117,In_680);
nand U945 (N_945,In_54,In_100);
or U946 (N_946,In_417,In_223);
nand U947 (N_947,In_418,In_272);
and U948 (N_948,In_516,In_75);
or U949 (N_949,In_500,In_616);
nand U950 (N_950,In_103,In_464);
or U951 (N_951,In_29,In_478);
nor U952 (N_952,In_692,In_312);
and U953 (N_953,In_4,In_267);
or U954 (N_954,In_329,In_632);
and U955 (N_955,In_652,In_165);
nor U956 (N_956,In_511,In_524);
or U957 (N_957,In_732,In_344);
and U958 (N_958,In_514,In_145);
nand U959 (N_959,In_643,In_315);
and U960 (N_960,In_647,In_48);
nor U961 (N_961,In_463,In_456);
or U962 (N_962,In_236,In_301);
xor U963 (N_963,In_372,In_378);
or U964 (N_964,In_458,In_246);
nand U965 (N_965,In_735,In_209);
xnor U966 (N_966,In_467,In_547);
xor U967 (N_967,In_218,In_208);
nor U968 (N_968,In_327,In_119);
and U969 (N_969,In_172,In_483);
or U970 (N_970,In_658,In_573);
or U971 (N_971,In_179,In_110);
and U972 (N_972,In_567,In_210);
xnor U973 (N_973,In_422,In_136);
and U974 (N_974,In_146,In_442);
and U975 (N_975,In_268,In_737);
xor U976 (N_976,In_652,In_511);
or U977 (N_977,In_373,In_528);
nor U978 (N_978,In_484,In_96);
nor U979 (N_979,In_561,In_644);
nand U980 (N_980,In_529,In_179);
nor U981 (N_981,In_428,In_271);
or U982 (N_982,In_717,In_536);
nand U983 (N_983,In_280,In_508);
nand U984 (N_984,In_254,In_349);
nand U985 (N_985,In_27,In_747);
nor U986 (N_986,In_43,In_602);
or U987 (N_987,In_724,In_408);
and U988 (N_988,In_633,In_307);
and U989 (N_989,In_374,In_204);
and U990 (N_990,In_509,In_532);
and U991 (N_991,In_116,In_308);
or U992 (N_992,In_217,In_143);
nand U993 (N_993,In_234,In_258);
or U994 (N_994,In_652,In_609);
nand U995 (N_995,In_18,In_329);
nor U996 (N_996,In_680,In_651);
nor U997 (N_997,In_518,In_167);
or U998 (N_998,In_523,In_271);
nor U999 (N_999,In_564,In_193);
and U1000 (N_1000,N_560,N_545);
nand U1001 (N_1001,N_904,N_426);
or U1002 (N_1002,N_215,N_171);
nand U1003 (N_1003,N_11,N_351);
and U1004 (N_1004,N_411,N_816);
nand U1005 (N_1005,N_820,N_988);
nand U1006 (N_1006,N_562,N_228);
nand U1007 (N_1007,N_658,N_864);
nand U1008 (N_1008,N_291,N_367);
nand U1009 (N_1009,N_42,N_389);
and U1010 (N_1010,N_143,N_59);
nor U1011 (N_1011,N_309,N_927);
xor U1012 (N_1012,N_428,N_718);
or U1013 (N_1013,N_721,N_583);
or U1014 (N_1014,N_916,N_992);
nor U1015 (N_1015,N_870,N_568);
or U1016 (N_1016,N_628,N_674);
nor U1017 (N_1017,N_585,N_517);
or U1018 (N_1018,N_182,N_914);
nor U1019 (N_1019,N_778,N_746);
xor U1020 (N_1020,N_414,N_344);
nand U1021 (N_1021,N_555,N_989);
nor U1022 (N_1022,N_233,N_556);
xor U1023 (N_1023,N_515,N_226);
nor U1024 (N_1024,N_489,N_177);
nand U1025 (N_1025,N_943,N_464);
and U1026 (N_1026,N_485,N_73);
nor U1027 (N_1027,N_796,N_969);
and U1028 (N_1028,N_981,N_536);
or U1029 (N_1029,N_187,N_5);
and U1030 (N_1030,N_317,N_93);
and U1031 (N_1031,N_833,N_297);
or U1032 (N_1032,N_249,N_624);
or U1033 (N_1033,N_172,N_645);
and U1034 (N_1034,N_807,N_72);
or U1035 (N_1035,N_479,N_600);
nor U1036 (N_1036,N_200,N_936);
or U1037 (N_1037,N_96,N_92);
and U1038 (N_1038,N_885,N_263);
or U1039 (N_1039,N_27,N_311);
and U1040 (N_1040,N_61,N_293);
nand U1041 (N_1041,N_980,N_691);
xor U1042 (N_1042,N_451,N_483);
and U1043 (N_1043,N_576,N_437);
xnor U1044 (N_1044,N_315,N_621);
nor U1045 (N_1045,N_396,N_97);
nor U1046 (N_1046,N_74,N_518);
or U1047 (N_1047,N_281,N_731);
nor U1048 (N_1048,N_789,N_363);
nand U1049 (N_1049,N_754,N_636);
nor U1050 (N_1050,N_951,N_30);
and U1051 (N_1051,N_136,N_52);
and U1052 (N_1052,N_629,N_592);
or U1053 (N_1053,N_186,N_204);
or U1054 (N_1054,N_429,N_610);
nor U1055 (N_1055,N_111,N_823);
nand U1056 (N_1056,N_727,N_28);
nand U1057 (N_1057,N_745,N_524);
nand U1058 (N_1058,N_597,N_366);
nor U1059 (N_1059,N_374,N_880);
xnor U1060 (N_1060,N_874,N_328);
and U1061 (N_1061,N_193,N_741);
xor U1062 (N_1062,N_318,N_744);
or U1063 (N_1063,N_57,N_888);
and U1064 (N_1064,N_595,N_675);
or U1065 (N_1065,N_492,N_825);
nor U1066 (N_1066,N_540,N_609);
or U1067 (N_1067,N_493,N_156);
nand U1068 (N_1068,N_323,N_973);
nand U1069 (N_1069,N_514,N_769);
nor U1070 (N_1070,N_46,N_991);
or U1071 (N_1071,N_574,N_605);
nand U1072 (N_1072,N_158,N_997);
or U1073 (N_1073,N_704,N_761);
or U1074 (N_1074,N_245,N_216);
nor U1075 (N_1075,N_314,N_112);
or U1076 (N_1076,N_584,N_655);
or U1077 (N_1077,N_896,N_640);
and U1078 (N_1078,N_693,N_300);
or U1079 (N_1079,N_47,N_902);
or U1080 (N_1080,N_108,N_661);
and U1081 (N_1081,N_89,N_627);
or U1082 (N_1082,N_252,N_801);
and U1083 (N_1083,N_931,N_787);
nor U1084 (N_1084,N_855,N_151);
and U1085 (N_1085,N_792,N_550);
nand U1086 (N_1086,N_841,N_569);
or U1087 (N_1087,N_41,N_697);
nor U1088 (N_1088,N_406,N_333);
and U1089 (N_1089,N_180,N_626);
nand U1090 (N_1090,N_734,N_821);
or U1091 (N_1091,N_917,N_152);
nor U1092 (N_1092,N_482,N_69);
xnor U1093 (N_1093,N_901,N_157);
or U1094 (N_1094,N_958,N_781);
and U1095 (N_1095,N_543,N_455);
nor U1096 (N_1096,N_993,N_702);
or U1097 (N_1097,N_649,N_207);
and U1098 (N_1098,N_651,N_33);
and U1099 (N_1099,N_898,N_647);
nor U1100 (N_1100,N_998,N_891);
nand U1101 (N_1101,N_736,N_673);
and U1102 (N_1102,N_394,N_461);
and U1103 (N_1103,N_18,N_928);
nor U1104 (N_1104,N_847,N_672);
nand U1105 (N_1105,N_742,N_375);
nor U1106 (N_1106,N_994,N_387);
nand U1107 (N_1107,N_504,N_979);
or U1108 (N_1108,N_716,N_341);
nand U1109 (N_1109,N_282,N_267);
and U1110 (N_1110,N_759,N_836);
or U1111 (N_1111,N_619,N_680);
and U1112 (N_1112,N_557,N_856);
and U1113 (N_1113,N_722,N_308);
and U1114 (N_1114,N_195,N_580);
or U1115 (N_1115,N_260,N_830);
nand U1116 (N_1116,N_723,N_444);
and U1117 (N_1117,N_85,N_918);
nand U1118 (N_1118,N_203,N_764);
nor U1119 (N_1119,N_51,N_295);
and U1120 (N_1120,N_503,N_133);
and U1121 (N_1121,N_468,N_635);
or U1122 (N_1122,N_714,N_607);
nor U1123 (N_1123,N_662,N_831);
nor U1124 (N_1124,N_280,N_412);
and U1125 (N_1125,N_911,N_832);
and U1126 (N_1126,N_961,N_601);
nor U1127 (N_1127,N_95,N_471);
nand U1128 (N_1128,N_330,N_554);
and U1129 (N_1129,N_337,N_110);
and U1130 (N_1130,N_866,N_138);
and U1131 (N_1131,N_279,N_301);
and U1132 (N_1132,N_433,N_729);
nand U1133 (N_1133,N_168,N_408);
nand U1134 (N_1134,N_712,N_613);
xnor U1135 (N_1135,N_771,N_534);
xnor U1136 (N_1136,N_586,N_677);
nor U1137 (N_1137,N_477,N_620);
or U1138 (N_1138,N_499,N_878);
nand U1139 (N_1139,N_999,N_386);
nor U1140 (N_1140,N_713,N_840);
or U1141 (N_1141,N_893,N_941);
and U1142 (N_1142,N_511,N_952);
nand U1143 (N_1143,N_405,N_895);
nor U1144 (N_1144,N_505,N_530);
nand U1145 (N_1145,N_425,N_197);
or U1146 (N_1146,N_362,N_750);
nor U1147 (N_1147,N_379,N_715);
nor U1148 (N_1148,N_273,N_546);
xor U1149 (N_1149,N_810,N_685);
and U1150 (N_1150,N_756,N_101);
nand U1151 (N_1151,N_278,N_173);
and U1152 (N_1152,N_860,N_488);
nor U1153 (N_1153,N_711,N_378);
nor U1154 (N_1154,N_522,N_799);
nor U1155 (N_1155,N_826,N_208);
xor U1156 (N_1156,N_82,N_637);
or U1157 (N_1157,N_946,N_127);
or U1158 (N_1158,N_292,N_25);
nand U1159 (N_1159,N_932,N_806);
or U1160 (N_1160,N_798,N_912);
and U1161 (N_1161,N_835,N_247);
and U1162 (N_1162,N_364,N_758);
nor U1163 (N_1163,N_706,N_719);
nor U1164 (N_1164,N_76,N_191);
nor U1165 (N_1165,N_659,N_199);
nor U1166 (N_1166,N_447,N_298);
nor U1167 (N_1167,N_147,N_126);
and U1168 (N_1168,N_224,N_415);
and U1169 (N_1169,N_780,N_777);
or U1170 (N_1170,N_162,N_211);
nand U1171 (N_1171,N_985,N_897);
or U1172 (N_1172,N_10,N_288);
xnor U1173 (N_1173,N_296,N_819);
or U1174 (N_1174,N_873,N_683);
xor U1175 (N_1175,N_2,N_434);
xor U1176 (N_1176,N_340,N_575);
and U1177 (N_1177,N_814,N_150);
nand U1178 (N_1178,N_775,N_632);
and U1179 (N_1179,N_502,N_265);
and U1180 (N_1180,N_383,N_606);
and U1181 (N_1181,N_472,N_903);
and U1182 (N_1182,N_995,N_497);
and U1183 (N_1183,N_776,N_269);
nor U1184 (N_1184,N_53,N_329);
nand U1185 (N_1185,N_264,N_109);
nand U1186 (N_1186,N_13,N_421);
or U1187 (N_1187,N_102,N_871);
or U1188 (N_1188,N_214,N_360);
nor U1189 (N_1189,N_839,N_889);
or U1190 (N_1190,N_377,N_356);
nand U1191 (N_1191,N_846,N_921);
and U1192 (N_1192,N_339,N_937);
nand U1193 (N_1193,N_805,N_652);
or U1194 (N_1194,N_163,N_972);
nor U1195 (N_1195,N_748,N_62);
nor U1196 (N_1196,N_132,N_355);
xnor U1197 (N_1197,N_441,N_35);
and U1198 (N_1198,N_246,N_751);
or U1199 (N_1199,N_749,N_578);
nand U1200 (N_1200,N_306,N_582);
nand U1201 (N_1201,N_347,N_469);
nand U1202 (N_1202,N_188,N_241);
or U1203 (N_1203,N_519,N_869);
xor U1204 (N_1204,N_420,N_178);
nand U1205 (N_1205,N_240,N_788);
nor U1206 (N_1206,N_385,N_770);
or U1207 (N_1207,N_445,N_802);
nor U1208 (N_1208,N_474,N_181);
or U1209 (N_1209,N_567,N_164);
xnor U1210 (N_1210,N_60,N_894);
nor U1211 (N_1211,N_539,N_122);
and U1212 (N_1212,N_665,N_448);
and U1213 (N_1213,N_38,N_75);
nor U1214 (N_1214,N_320,N_700);
nor U1215 (N_1215,N_531,N_4);
nand U1216 (N_1216,N_201,N_392);
nand U1217 (N_1217,N_752,N_290);
xnor U1218 (N_1218,N_521,N_454);
xnor U1219 (N_1219,N_361,N_648);
nand U1220 (N_1220,N_862,N_274);
and U1221 (N_1221,N_91,N_354);
or U1222 (N_1222,N_822,N_236);
or U1223 (N_1223,N_848,N_343);
or U1224 (N_1224,N_81,N_452);
nor U1225 (N_1225,N_432,N_671);
or U1226 (N_1226,N_579,N_622);
or U1227 (N_1227,N_460,N_844);
nor U1228 (N_1228,N_940,N_430);
nand U1229 (N_1229,N_922,N_99);
nand U1230 (N_1230,N_310,N_17);
nor U1231 (N_1231,N_496,N_221);
nor U1232 (N_1232,N_528,N_66);
nand U1233 (N_1233,N_321,N_403);
nand U1234 (N_1234,N_743,N_467);
and U1235 (N_1235,N_0,N_950);
nand U1236 (N_1236,N_65,N_970);
nor U1237 (N_1237,N_209,N_986);
xnor U1238 (N_1238,N_537,N_368);
nand U1239 (N_1239,N_148,N_319);
or U1240 (N_1240,N_602,N_312);
xor U1241 (N_1241,N_436,N_890);
nand U1242 (N_1242,N_774,N_174);
or U1243 (N_1243,N_755,N_68);
nor U1244 (N_1244,N_786,N_538);
nor U1245 (N_1245,N_114,N_220);
and U1246 (N_1246,N_234,N_948);
or U1247 (N_1247,N_254,N_695);
or U1248 (N_1248,N_768,N_210);
or U1249 (N_1249,N_262,N_813);
nand U1250 (N_1250,N_56,N_868);
or U1251 (N_1251,N_160,N_924);
nor U1252 (N_1252,N_527,N_990);
and U1253 (N_1253,N_116,N_123);
nand U1254 (N_1254,N_884,N_244);
nor U1255 (N_1255,N_54,N_762);
or U1256 (N_1256,N_849,N_974);
nand U1257 (N_1257,N_283,N_303);
nor U1258 (N_1258,N_790,N_535);
and U1259 (N_1259,N_212,N_670);
or U1260 (N_1260,N_570,N_760);
nand U1261 (N_1261,N_190,N_881);
nor U1262 (N_1262,N_299,N_703);
and U1263 (N_1263,N_735,N_106);
nor U1264 (N_1264,N_803,N_266);
nand U1265 (N_1265,N_612,N_842);
nand U1266 (N_1266,N_161,N_663);
nor U1267 (N_1267,N_45,N_407);
or U1268 (N_1268,N_782,N_446);
nor U1269 (N_1269,N_380,N_603);
nand U1270 (N_1270,N_804,N_596);
and U1271 (N_1271,N_653,N_906);
nor U1272 (N_1272,N_410,N_625);
nor U1273 (N_1273,N_36,N_508);
or U1274 (N_1274,N_591,N_564);
or U1275 (N_1275,N_643,N_84);
nand U1276 (N_1276,N_581,N_747);
and U1277 (N_1277,N_128,N_382);
or U1278 (N_1278,N_144,N_589);
or U1279 (N_1279,N_783,N_867);
and U1280 (N_1280,N_975,N_23);
and U1281 (N_1281,N_397,N_934);
nand U1282 (N_1282,N_276,N_231);
or U1283 (N_1283,N_863,N_573);
and U1284 (N_1284,N_795,N_342);
or U1285 (N_1285,N_325,N_409);
or U1286 (N_1286,N_944,N_359);
xor U1287 (N_1287,N_498,N_724);
nand U1288 (N_1288,N_525,N_271);
nor U1289 (N_1289,N_456,N_400);
or U1290 (N_1290,N_646,N_939);
nor U1291 (N_1291,N_717,N_352);
xor U1292 (N_1292,N_614,N_561);
and U1293 (N_1293,N_563,N_834);
nor U1294 (N_1294,N_350,N_476);
nor U1295 (N_1295,N_542,N_141);
nand U1296 (N_1296,N_376,N_399);
and U1297 (N_1297,N_851,N_86);
or U1298 (N_1298,N_277,N_590);
nor U1299 (N_1299,N_935,N_63);
or U1300 (N_1300,N_919,N_817);
nand U1301 (N_1301,N_113,N_19);
or U1302 (N_1302,N_370,N_316);
nand U1303 (N_1303,N_184,N_552);
nand U1304 (N_1304,N_500,N_529);
xor U1305 (N_1305,N_966,N_78);
or U1306 (N_1306,N_64,N_737);
nor U1307 (N_1307,N_879,N_920);
or U1308 (N_1308,N_598,N_438);
and U1309 (N_1309,N_43,N_235);
xor U1310 (N_1310,N_681,N_690);
xnor U1311 (N_1311,N_326,N_779);
xor U1312 (N_1312,N_139,N_965);
and U1313 (N_1313,N_617,N_730);
or U1314 (N_1314,N_194,N_733);
nor U1315 (N_1315,N_431,N_166);
nand U1316 (N_1316,N_983,N_140);
nand U1317 (N_1317,N_219,N_812);
xnor U1318 (N_1318,N_899,N_103);
nor U1319 (N_1319,N_587,N_107);
and U1320 (N_1320,N_694,N_21);
nand U1321 (N_1321,N_401,N_687);
or U1322 (N_1322,N_322,N_845);
or U1323 (N_1323,N_887,N_79);
nand U1324 (N_1324,N_442,N_134);
or U1325 (N_1325,N_766,N_506);
and U1326 (N_1326,N_424,N_439);
and U1327 (N_1327,N_689,N_270);
nand U1328 (N_1328,N_559,N_686);
nand U1329 (N_1329,N_630,N_149);
and U1330 (N_1330,N_900,N_459);
xor U1331 (N_1331,N_213,N_544);
nand U1332 (N_1332,N_242,N_512);
nand U1333 (N_1333,N_551,N_237);
and U1334 (N_1334,N_227,N_656);
nor U1335 (N_1335,N_167,N_302);
or U1336 (N_1336,N_800,N_416);
xnor U1337 (N_1337,N_883,N_185);
nor U1338 (N_1338,N_668,N_791);
nand U1339 (N_1339,N_594,N_55);
xnor U1340 (N_1340,N_962,N_83);
xor U1341 (N_1341,N_772,N_960);
or U1342 (N_1342,N_501,N_6);
nand U1343 (N_1343,N_473,N_809);
and U1344 (N_1344,N_169,N_858);
and U1345 (N_1345,N_165,N_117);
or U1346 (N_1346,N_324,N_877);
and U1347 (N_1347,N_558,N_34);
nand U1348 (N_1348,N_657,N_593);
nor U1349 (N_1349,N_478,N_987);
nor U1350 (N_1350,N_876,N_153);
or U1351 (N_1351,N_955,N_608);
or U1352 (N_1352,N_577,N_358);
nor U1353 (N_1353,N_49,N_572);
or U1354 (N_1354,N_440,N_910);
nor U1355 (N_1355,N_963,N_953);
nor U1356 (N_1356,N_29,N_229);
nand U1357 (N_1357,N_225,N_119);
xnor U1358 (N_1358,N_696,N_838);
xnor U1359 (N_1359,N_740,N_450);
and U1360 (N_1360,N_170,N_913);
nand U1361 (N_1361,N_548,N_159);
and U1362 (N_1362,N_331,N_682);
and U1363 (N_1363,N_604,N_865);
and U1364 (N_1364,N_907,N_205);
or U1365 (N_1365,N_80,N_7);
or U1366 (N_1366,N_175,N_176);
or U1367 (N_1367,N_285,N_705);
or U1368 (N_1368,N_239,N_115);
and U1369 (N_1369,N_349,N_335);
and U1370 (N_1370,N_815,N_892);
and U1371 (N_1371,N_490,N_419);
nor U1372 (N_1372,N_667,N_230);
and U1373 (N_1373,N_692,N_268);
and U1374 (N_1374,N_125,N_391);
nor U1375 (N_1375,N_94,N_785);
nor U1376 (N_1376,N_3,N_763);
or U1377 (N_1377,N_929,N_384);
xnor U1378 (N_1378,N_256,N_725);
or U1379 (N_1379,N_824,N_925);
nor U1380 (N_1380,N_676,N_124);
and U1381 (N_1381,N_954,N_611);
nand U1382 (N_1382,N_688,N_765);
and U1383 (N_1383,N_753,N_644);
nand U1384 (N_1384,N_257,N_549);
nor U1385 (N_1385,N_872,N_395);
nand U1386 (N_1386,N_250,N_357);
or U1387 (N_1387,N_369,N_470);
and U1388 (N_1388,N_571,N_307);
or U1389 (N_1389,N_660,N_336);
nor U1390 (N_1390,N_684,N_238);
and U1391 (N_1391,N_413,N_243);
nor U1392 (N_1392,N_664,N_218);
nand U1393 (N_1393,N_404,N_793);
and U1394 (N_1394,N_466,N_398);
and U1395 (N_1395,N_313,N_50);
or U1396 (N_1396,N_457,N_289);
nor U1397 (N_1397,N_393,N_372);
nand U1398 (N_1398,N_631,N_137);
nor U1399 (N_1399,N_509,N_638);
nor U1400 (N_1400,N_70,N_859);
or U1401 (N_1401,N_48,N_487);
xnor U1402 (N_1402,N_959,N_390);
or U1403 (N_1403,N_131,N_930);
nand U1404 (N_1404,N_971,N_305);
and U1405 (N_1405,N_808,N_978);
and U1406 (N_1406,N_633,N_259);
nand U1407 (N_1407,N_905,N_192);
nand U1408 (N_1408,N_67,N_945);
and U1409 (N_1409,N_738,N_728);
nor U1410 (N_1410,N_679,N_222);
nor U1411 (N_1411,N_850,N_258);
xor U1412 (N_1412,N_526,N_449);
nand U1413 (N_1413,N_135,N_964);
nand U1414 (N_1414,N_44,N_784);
xor U1415 (N_1415,N_698,N_565);
or U1416 (N_1416,N_32,N_829);
xor U1417 (N_1417,N_853,N_287);
nor U1418 (N_1418,N_938,N_516);
nor U1419 (N_1419,N_20,N_486);
nand U1420 (N_1420,N_31,N_491);
nor U1421 (N_1421,N_926,N_286);
nand U1422 (N_1422,N_272,N_707);
nand U1423 (N_1423,N_566,N_861);
and U1424 (N_1424,N_666,N_304);
nor U1425 (N_1425,N_957,N_701);
and U1426 (N_1426,N_121,N_22);
nand U1427 (N_1427,N_251,N_402);
and U1428 (N_1428,N_739,N_26);
xor U1429 (N_1429,N_933,N_422);
nand U1430 (N_1430,N_183,N_154);
and U1431 (N_1431,N_353,N_206);
nor U1432 (N_1432,N_923,N_494);
and U1433 (N_1433,N_767,N_942);
or U1434 (N_1434,N_248,N_130);
and U1435 (N_1435,N_513,N_435);
or U1436 (N_1436,N_484,N_720);
xor U1437 (N_1437,N_843,N_507);
and U1438 (N_1438,N_155,N_345);
nor U1439 (N_1439,N_547,N_196);
nand U1440 (N_1440,N_373,N_875);
nand U1441 (N_1441,N_996,N_275);
and U1442 (N_1442,N_857,N_223);
and U1443 (N_1443,N_24,N_37);
and U1444 (N_1444,N_261,N_423);
or U1445 (N_1445,N_886,N_16);
or U1446 (N_1446,N_198,N_797);
and U1447 (N_1447,N_618,N_202);
xor U1448 (N_1448,N_388,N_982);
xor U1449 (N_1449,N_338,N_427);
or U1450 (N_1450,N_98,N_811);
nand U1451 (N_1451,N_87,N_40);
nand U1452 (N_1452,N_709,N_827);
or U1453 (N_1453,N_699,N_616);
and U1454 (N_1454,N_118,N_773);
nor U1455 (N_1455,N_977,N_332);
nand U1456 (N_1456,N_854,N_669);
nor U1457 (N_1457,N_453,N_348);
nor U1458 (N_1458,N_599,N_284);
nand U1459 (N_1459,N_634,N_179);
nand U1460 (N_1460,N_142,N_371);
and U1461 (N_1461,N_481,N_523);
nor U1462 (N_1462,N_949,N_255);
or U1463 (N_1463,N_678,N_463);
xnor U1464 (N_1464,N_732,N_458);
nand U1465 (N_1465,N_346,N_253);
or U1466 (N_1466,N_757,N_976);
and U1467 (N_1467,N_837,N_294);
nor U1468 (N_1468,N_710,N_708);
or U1469 (N_1469,N_532,N_908);
or U1470 (N_1470,N_105,N_984);
nand U1471 (N_1471,N_641,N_381);
nor U1472 (N_1472,N_553,N_129);
nor U1473 (N_1473,N_623,N_9);
and U1474 (N_1474,N_462,N_510);
or U1475 (N_1475,N_520,N_654);
or U1476 (N_1476,N_642,N_967);
nor U1477 (N_1477,N_968,N_475);
nand U1478 (N_1478,N_947,N_852);
nand U1479 (N_1479,N_465,N_639);
nand U1480 (N_1480,N_480,N_327);
and U1481 (N_1481,N_915,N_818);
and U1482 (N_1482,N_71,N_145);
nor U1483 (N_1483,N_726,N_232);
xor U1484 (N_1484,N_533,N_146);
nand U1485 (N_1485,N_58,N_541);
nand U1486 (N_1486,N_650,N_1);
or U1487 (N_1487,N_365,N_334);
or U1488 (N_1488,N_588,N_909);
or U1489 (N_1489,N_15,N_120);
or U1490 (N_1490,N_100,N_39);
or U1491 (N_1491,N_828,N_615);
xor U1492 (N_1492,N_104,N_88);
and U1493 (N_1493,N_14,N_443);
or U1494 (N_1494,N_417,N_495);
nor U1495 (N_1495,N_90,N_794);
xnor U1496 (N_1496,N_189,N_418);
or U1497 (N_1497,N_882,N_956);
nand U1498 (N_1498,N_8,N_217);
xor U1499 (N_1499,N_77,N_12);
or U1500 (N_1500,N_451,N_530);
or U1501 (N_1501,N_285,N_895);
nor U1502 (N_1502,N_583,N_584);
nand U1503 (N_1503,N_327,N_674);
or U1504 (N_1504,N_965,N_76);
or U1505 (N_1505,N_889,N_55);
nand U1506 (N_1506,N_156,N_714);
and U1507 (N_1507,N_520,N_9);
nand U1508 (N_1508,N_383,N_838);
or U1509 (N_1509,N_813,N_56);
or U1510 (N_1510,N_946,N_704);
xor U1511 (N_1511,N_933,N_887);
nor U1512 (N_1512,N_131,N_139);
or U1513 (N_1513,N_643,N_442);
nor U1514 (N_1514,N_16,N_990);
nor U1515 (N_1515,N_950,N_377);
nor U1516 (N_1516,N_653,N_384);
nor U1517 (N_1517,N_334,N_854);
nor U1518 (N_1518,N_336,N_481);
xnor U1519 (N_1519,N_957,N_200);
nor U1520 (N_1520,N_963,N_26);
nand U1521 (N_1521,N_268,N_816);
or U1522 (N_1522,N_243,N_961);
or U1523 (N_1523,N_118,N_777);
nand U1524 (N_1524,N_505,N_838);
and U1525 (N_1525,N_798,N_485);
or U1526 (N_1526,N_880,N_810);
and U1527 (N_1527,N_706,N_380);
and U1528 (N_1528,N_36,N_808);
and U1529 (N_1529,N_459,N_845);
or U1530 (N_1530,N_638,N_394);
and U1531 (N_1531,N_768,N_494);
nand U1532 (N_1532,N_278,N_540);
nand U1533 (N_1533,N_898,N_225);
or U1534 (N_1534,N_301,N_706);
nor U1535 (N_1535,N_742,N_618);
and U1536 (N_1536,N_718,N_852);
and U1537 (N_1537,N_541,N_605);
nand U1538 (N_1538,N_956,N_818);
and U1539 (N_1539,N_546,N_973);
nand U1540 (N_1540,N_336,N_499);
nor U1541 (N_1541,N_278,N_771);
and U1542 (N_1542,N_854,N_802);
and U1543 (N_1543,N_255,N_155);
and U1544 (N_1544,N_909,N_729);
or U1545 (N_1545,N_21,N_921);
nand U1546 (N_1546,N_535,N_240);
nor U1547 (N_1547,N_586,N_714);
and U1548 (N_1548,N_732,N_289);
nor U1549 (N_1549,N_482,N_862);
nand U1550 (N_1550,N_991,N_948);
or U1551 (N_1551,N_621,N_421);
nor U1552 (N_1552,N_192,N_975);
nor U1553 (N_1553,N_604,N_386);
nor U1554 (N_1554,N_692,N_166);
xnor U1555 (N_1555,N_204,N_966);
and U1556 (N_1556,N_621,N_583);
nor U1557 (N_1557,N_491,N_821);
nand U1558 (N_1558,N_159,N_248);
and U1559 (N_1559,N_12,N_290);
or U1560 (N_1560,N_96,N_940);
nand U1561 (N_1561,N_846,N_419);
nor U1562 (N_1562,N_354,N_85);
or U1563 (N_1563,N_509,N_376);
or U1564 (N_1564,N_564,N_671);
or U1565 (N_1565,N_859,N_968);
nand U1566 (N_1566,N_68,N_439);
and U1567 (N_1567,N_724,N_855);
and U1568 (N_1568,N_643,N_803);
xor U1569 (N_1569,N_490,N_165);
or U1570 (N_1570,N_654,N_345);
nor U1571 (N_1571,N_848,N_483);
nor U1572 (N_1572,N_889,N_823);
nand U1573 (N_1573,N_659,N_114);
xnor U1574 (N_1574,N_213,N_755);
and U1575 (N_1575,N_851,N_659);
and U1576 (N_1576,N_691,N_160);
nor U1577 (N_1577,N_2,N_27);
xnor U1578 (N_1578,N_488,N_569);
nor U1579 (N_1579,N_400,N_883);
nor U1580 (N_1580,N_312,N_234);
nand U1581 (N_1581,N_844,N_208);
nor U1582 (N_1582,N_859,N_112);
xor U1583 (N_1583,N_415,N_691);
nand U1584 (N_1584,N_954,N_604);
and U1585 (N_1585,N_929,N_332);
xor U1586 (N_1586,N_927,N_725);
nor U1587 (N_1587,N_788,N_349);
nand U1588 (N_1588,N_252,N_362);
and U1589 (N_1589,N_926,N_339);
and U1590 (N_1590,N_320,N_119);
nand U1591 (N_1591,N_393,N_241);
and U1592 (N_1592,N_445,N_134);
xnor U1593 (N_1593,N_237,N_127);
or U1594 (N_1594,N_310,N_701);
or U1595 (N_1595,N_303,N_157);
or U1596 (N_1596,N_86,N_467);
nor U1597 (N_1597,N_944,N_984);
and U1598 (N_1598,N_405,N_102);
nand U1599 (N_1599,N_328,N_154);
nand U1600 (N_1600,N_114,N_412);
and U1601 (N_1601,N_101,N_457);
or U1602 (N_1602,N_732,N_524);
nor U1603 (N_1603,N_841,N_301);
nand U1604 (N_1604,N_316,N_343);
or U1605 (N_1605,N_458,N_476);
xnor U1606 (N_1606,N_195,N_124);
nor U1607 (N_1607,N_94,N_403);
and U1608 (N_1608,N_473,N_248);
nor U1609 (N_1609,N_609,N_857);
and U1610 (N_1610,N_819,N_226);
or U1611 (N_1611,N_99,N_459);
or U1612 (N_1612,N_272,N_904);
nand U1613 (N_1613,N_518,N_311);
nor U1614 (N_1614,N_251,N_307);
nand U1615 (N_1615,N_234,N_211);
nor U1616 (N_1616,N_999,N_715);
or U1617 (N_1617,N_100,N_362);
xor U1618 (N_1618,N_657,N_157);
or U1619 (N_1619,N_138,N_163);
xnor U1620 (N_1620,N_738,N_694);
or U1621 (N_1621,N_634,N_118);
and U1622 (N_1622,N_131,N_410);
nand U1623 (N_1623,N_970,N_443);
nor U1624 (N_1624,N_727,N_4);
or U1625 (N_1625,N_134,N_731);
xor U1626 (N_1626,N_251,N_41);
xor U1627 (N_1627,N_804,N_911);
and U1628 (N_1628,N_527,N_273);
nor U1629 (N_1629,N_492,N_953);
and U1630 (N_1630,N_115,N_273);
xor U1631 (N_1631,N_131,N_285);
nor U1632 (N_1632,N_462,N_458);
nand U1633 (N_1633,N_129,N_62);
and U1634 (N_1634,N_156,N_148);
or U1635 (N_1635,N_342,N_208);
nand U1636 (N_1636,N_879,N_562);
nor U1637 (N_1637,N_164,N_328);
nor U1638 (N_1638,N_76,N_124);
nor U1639 (N_1639,N_664,N_962);
and U1640 (N_1640,N_667,N_50);
and U1641 (N_1641,N_866,N_195);
nand U1642 (N_1642,N_555,N_967);
or U1643 (N_1643,N_886,N_438);
or U1644 (N_1644,N_992,N_118);
or U1645 (N_1645,N_156,N_26);
or U1646 (N_1646,N_84,N_203);
and U1647 (N_1647,N_967,N_696);
or U1648 (N_1648,N_90,N_311);
nor U1649 (N_1649,N_108,N_401);
or U1650 (N_1650,N_382,N_129);
nor U1651 (N_1651,N_892,N_918);
nand U1652 (N_1652,N_384,N_494);
and U1653 (N_1653,N_991,N_157);
nor U1654 (N_1654,N_737,N_754);
xnor U1655 (N_1655,N_307,N_451);
nor U1656 (N_1656,N_364,N_876);
and U1657 (N_1657,N_833,N_240);
xor U1658 (N_1658,N_405,N_119);
or U1659 (N_1659,N_153,N_410);
or U1660 (N_1660,N_592,N_138);
and U1661 (N_1661,N_660,N_233);
xnor U1662 (N_1662,N_174,N_909);
nand U1663 (N_1663,N_351,N_94);
and U1664 (N_1664,N_638,N_170);
and U1665 (N_1665,N_145,N_55);
nand U1666 (N_1666,N_755,N_903);
nand U1667 (N_1667,N_308,N_821);
and U1668 (N_1668,N_589,N_875);
nand U1669 (N_1669,N_853,N_122);
nor U1670 (N_1670,N_763,N_647);
and U1671 (N_1671,N_682,N_832);
and U1672 (N_1672,N_267,N_249);
xnor U1673 (N_1673,N_186,N_830);
nand U1674 (N_1674,N_664,N_547);
or U1675 (N_1675,N_598,N_918);
or U1676 (N_1676,N_903,N_435);
nand U1677 (N_1677,N_649,N_254);
or U1678 (N_1678,N_502,N_838);
nor U1679 (N_1679,N_135,N_656);
nand U1680 (N_1680,N_306,N_564);
nor U1681 (N_1681,N_289,N_719);
xnor U1682 (N_1682,N_677,N_647);
nand U1683 (N_1683,N_976,N_25);
or U1684 (N_1684,N_185,N_930);
nand U1685 (N_1685,N_465,N_58);
nand U1686 (N_1686,N_506,N_649);
nor U1687 (N_1687,N_155,N_899);
nand U1688 (N_1688,N_393,N_72);
nor U1689 (N_1689,N_718,N_800);
or U1690 (N_1690,N_656,N_276);
or U1691 (N_1691,N_908,N_348);
and U1692 (N_1692,N_916,N_474);
nor U1693 (N_1693,N_379,N_417);
nand U1694 (N_1694,N_303,N_94);
and U1695 (N_1695,N_85,N_79);
and U1696 (N_1696,N_973,N_476);
or U1697 (N_1697,N_113,N_314);
nor U1698 (N_1698,N_551,N_168);
or U1699 (N_1699,N_393,N_982);
nor U1700 (N_1700,N_371,N_434);
nand U1701 (N_1701,N_603,N_976);
and U1702 (N_1702,N_385,N_145);
xor U1703 (N_1703,N_986,N_570);
or U1704 (N_1704,N_973,N_667);
or U1705 (N_1705,N_733,N_255);
or U1706 (N_1706,N_386,N_606);
or U1707 (N_1707,N_137,N_655);
nor U1708 (N_1708,N_191,N_359);
or U1709 (N_1709,N_98,N_303);
and U1710 (N_1710,N_155,N_473);
nor U1711 (N_1711,N_136,N_0);
xor U1712 (N_1712,N_885,N_915);
or U1713 (N_1713,N_750,N_145);
nand U1714 (N_1714,N_857,N_178);
and U1715 (N_1715,N_721,N_586);
xor U1716 (N_1716,N_863,N_307);
and U1717 (N_1717,N_162,N_919);
and U1718 (N_1718,N_981,N_602);
or U1719 (N_1719,N_984,N_611);
nand U1720 (N_1720,N_703,N_394);
and U1721 (N_1721,N_641,N_499);
or U1722 (N_1722,N_529,N_816);
nor U1723 (N_1723,N_803,N_814);
and U1724 (N_1724,N_474,N_709);
xor U1725 (N_1725,N_364,N_206);
or U1726 (N_1726,N_495,N_82);
or U1727 (N_1727,N_865,N_99);
or U1728 (N_1728,N_861,N_675);
or U1729 (N_1729,N_287,N_569);
and U1730 (N_1730,N_483,N_529);
nor U1731 (N_1731,N_277,N_694);
or U1732 (N_1732,N_315,N_437);
and U1733 (N_1733,N_181,N_486);
and U1734 (N_1734,N_330,N_263);
and U1735 (N_1735,N_249,N_781);
xor U1736 (N_1736,N_455,N_310);
or U1737 (N_1737,N_705,N_4);
nand U1738 (N_1738,N_244,N_229);
and U1739 (N_1739,N_515,N_862);
nor U1740 (N_1740,N_413,N_649);
nand U1741 (N_1741,N_591,N_709);
and U1742 (N_1742,N_710,N_961);
or U1743 (N_1743,N_4,N_332);
or U1744 (N_1744,N_95,N_920);
nor U1745 (N_1745,N_670,N_519);
and U1746 (N_1746,N_79,N_631);
and U1747 (N_1747,N_978,N_517);
nor U1748 (N_1748,N_851,N_388);
or U1749 (N_1749,N_825,N_166);
or U1750 (N_1750,N_380,N_445);
and U1751 (N_1751,N_865,N_538);
and U1752 (N_1752,N_908,N_517);
and U1753 (N_1753,N_364,N_851);
nor U1754 (N_1754,N_718,N_480);
nor U1755 (N_1755,N_895,N_447);
nor U1756 (N_1756,N_299,N_576);
or U1757 (N_1757,N_812,N_787);
nor U1758 (N_1758,N_904,N_883);
or U1759 (N_1759,N_759,N_286);
or U1760 (N_1760,N_999,N_159);
and U1761 (N_1761,N_430,N_269);
xor U1762 (N_1762,N_472,N_833);
and U1763 (N_1763,N_820,N_314);
or U1764 (N_1764,N_517,N_584);
and U1765 (N_1765,N_927,N_827);
nor U1766 (N_1766,N_51,N_164);
and U1767 (N_1767,N_15,N_193);
xor U1768 (N_1768,N_184,N_861);
or U1769 (N_1769,N_509,N_445);
or U1770 (N_1770,N_211,N_285);
or U1771 (N_1771,N_143,N_930);
xor U1772 (N_1772,N_730,N_767);
nand U1773 (N_1773,N_533,N_802);
and U1774 (N_1774,N_781,N_537);
nand U1775 (N_1775,N_467,N_403);
and U1776 (N_1776,N_17,N_545);
xnor U1777 (N_1777,N_387,N_689);
nand U1778 (N_1778,N_406,N_409);
and U1779 (N_1779,N_34,N_116);
nand U1780 (N_1780,N_376,N_613);
nor U1781 (N_1781,N_675,N_833);
and U1782 (N_1782,N_929,N_889);
xnor U1783 (N_1783,N_814,N_724);
and U1784 (N_1784,N_18,N_189);
nor U1785 (N_1785,N_699,N_623);
or U1786 (N_1786,N_996,N_18);
xor U1787 (N_1787,N_211,N_664);
xor U1788 (N_1788,N_624,N_362);
nor U1789 (N_1789,N_707,N_871);
nor U1790 (N_1790,N_39,N_443);
xor U1791 (N_1791,N_198,N_600);
xor U1792 (N_1792,N_644,N_425);
and U1793 (N_1793,N_481,N_995);
or U1794 (N_1794,N_646,N_776);
or U1795 (N_1795,N_633,N_769);
and U1796 (N_1796,N_951,N_579);
nor U1797 (N_1797,N_493,N_192);
nor U1798 (N_1798,N_105,N_898);
nor U1799 (N_1799,N_504,N_181);
and U1800 (N_1800,N_184,N_67);
nor U1801 (N_1801,N_494,N_871);
and U1802 (N_1802,N_373,N_643);
or U1803 (N_1803,N_536,N_521);
xor U1804 (N_1804,N_887,N_753);
nand U1805 (N_1805,N_688,N_626);
nor U1806 (N_1806,N_957,N_949);
nor U1807 (N_1807,N_242,N_892);
nand U1808 (N_1808,N_584,N_989);
xor U1809 (N_1809,N_687,N_864);
and U1810 (N_1810,N_51,N_410);
nand U1811 (N_1811,N_675,N_320);
nor U1812 (N_1812,N_880,N_586);
or U1813 (N_1813,N_274,N_454);
and U1814 (N_1814,N_862,N_891);
xor U1815 (N_1815,N_428,N_936);
and U1816 (N_1816,N_368,N_349);
nor U1817 (N_1817,N_605,N_416);
xnor U1818 (N_1818,N_851,N_650);
nor U1819 (N_1819,N_238,N_364);
xor U1820 (N_1820,N_68,N_747);
and U1821 (N_1821,N_505,N_276);
nand U1822 (N_1822,N_131,N_235);
nand U1823 (N_1823,N_698,N_952);
nand U1824 (N_1824,N_720,N_749);
and U1825 (N_1825,N_218,N_868);
and U1826 (N_1826,N_973,N_806);
and U1827 (N_1827,N_801,N_967);
and U1828 (N_1828,N_509,N_20);
nand U1829 (N_1829,N_928,N_807);
or U1830 (N_1830,N_84,N_420);
xor U1831 (N_1831,N_280,N_396);
and U1832 (N_1832,N_499,N_438);
nand U1833 (N_1833,N_942,N_795);
nand U1834 (N_1834,N_884,N_700);
xor U1835 (N_1835,N_518,N_121);
or U1836 (N_1836,N_351,N_118);
and U1837 (N_1837,N_701,N_467);
nor U1838 (N_1838,N_845,N_591);
and U1839 (N_1839,N_348,N_668);
nor U1840 (N_1840,N_323,N_820);
and U1841 (N_1841,N_88,N_161);
and U1842 (N_1842,N_302,N_371);
nand U1843 (N_1843,N_938,N_734);
and U1844 (N_1844,N_908,N_192);
nor U1845 (N_1845,N_461,N_799);
nor U1846 (N_1846,N_297,N_974);
nand U1847 (N_1847,N_110,N_715);
nand U1848 (N_1848,N_173,N_562);
xor U1849 (N_1849,N_1,N_322);
or U1850 (N_1850,N_477,N_112);
and U1851 (N_1851,N_442,N_612);
nand U1852 (N_1852,N_461,N_656);
nand U1853 (N_1853,N_855,N_758);
nand U1854 (N_1854,N_937,N_207);
and U1855 (N_1855,N_26,N_947);
and U1856 (N_1856,N_361,N_666);
or U1857 (N_1857,N_628,N_641);
and U1858 (N_1858,N_556,N_810);
and U1859 (N_1859,N_671,N_676);
or U1860 (N_1860,N_450,N_674);
or U1861 (N_1861,N_574,N_582);
and U1862 (N_1862,N_404,N_684);
nand U1863 (N_1863,N_19,N_909);
nor U1864 (N_1864,N_225,N_905);
or U1865 (N_1865,N_691,N_127);
nand U1866 (N_1866,N_379,N_146);
nand U1867 (N_1867,N_570,N_151);
or U1868 (N_1868,N_795,N_366);
and U1869 (N_1869,N_784,N_903);
nor U1870 (N_1870,N_746,N_231);
nand U1871 (N_1871,N_704,N_939);
nand U1872 (N_1872,N_498,N_352);
nand U1873 (N_1873,N_890,N_648);
and U1874 (N_1874,N_214,N_356);
nor U1875 (N_1875,N_363,N_239);
nand U1876 (N_1876,N_663,N_812);
nand U1877 (N_1877,N_338,N_747);
nor U1878 (N_1878,N_573,N_972);
nor U1879 (N_1879,N_433,N_23);
nor U1880 (N_1880,N_234,N_172);
and U1881 (N_1881,N_890,N_38);
nand U1882 (N_1882,N_753,N_207);
nand U1883 (N_1883,N_647,N_338);
nor U1884 (N_1884,N_455,N_814);
and U1885 (N_1885,N_398,N_633);
or U1886 (N_1886,N_833,N_174);
nand U1887 (N_1887,N_87,N_283);
and U1888 (N_1888,N_812,N_677);
nand U1889 (N_1889,N_413,N_175);
nor U1890 (N_1890,N_343,N_112);
or U1891 (N_1891,N_838,N_744);
nor U1892 (N_1892,N_679,N_395);
nand U1893 (N_1893,N_275,N_304);
nand U1894 (N_1894,N_904,N_351);
nand U1895 (N_1895,N_635,N_574);
or U1896 (N_1896,N_495,N_544);
xnor U1897 (N_1897,N_705,N_991);
and U1898 (N_1898,N_102,N_982);
and U1899 (N_1899,N_588,N_764);
nor U1900 (N_1900,N_291,N_630);
and U1901 (N_1901,N_644,N_508);
or U1902 (N_1902,N_919,N_962);
nor U1903 (N_1903,N_91,N_15);
nor U1904 (N_1904,N_80,N_9);
nand U1905 (N_1905,N_649,N_392);
nand U1906 (N_1906,N_997,N_927);
nand U1907 (N_1907,N_187,N_885);
nand U1908 (N_1908,N_187,N_92);
nand U1909 (N_1909,N_836,N_941);
or U1910 (N_1910,N_283,N_304);
nor U1911 (N_1911,N_900,N_96);
and U1912 (N_1912,N_860,N_799);
or U1913 (N_1913,N_533,N_8);
nor U1914 (N_1914,N_581,N_758);
nor U1915 (N_1915,N_820,N_690);
nand U1916 (N_1916,N_354,N_545);
xor U1917 (N_1917,N_274,N_636);
and U1918 (N_1918,N_289,N_214);
nor U1919 (N_1919,N_49,N_80);
nand U1920 (N_1920,N_527,N_327);
nand U1921 (N_1921,N_820,N_449);
and U1922 (N_1922,N_769,N_128);
or U1923 (N_1923,N_79,N_894);
nand U1924 (N_1924,N_773,N_906);
or U1925 (N_1925,N_332,N_612);
nand U1926 (N_1926,N_682,N_45);
xnor U1927 (N_1927,N_777,N_414);
or U1928 (N_1928,N_476,N_155);
and U1929 (N_1929,N_299,N_574);
nand U1930 (N_1930,N_990,N_40);
and U1931 (N_1931,N_31,N_233);
xnor U1932 (N_1932,N_189,N_406);
and U1933 (N_1933,N_376,N_190);
nor U1934 (N_1934,N_404,N_406);
and U1935 (N_1935,N_982,N_22);
or U1936 (N_1936,N_8,N_339);
and U1937 (N_1937,N_3,N_490);
xor U1938 (N_1938,N_272,N_42);
or U1939 (N_1939,N_467,N_203);
and U1940 (N_1940,N_226,N_250);
xor U1941 (N_1941,N_897,N_625);
or U1942 (N_1942,N_530,N_741);
nand U1943 (N_1943,N_574,N_157);
nand U1944 (N_1944,N_607,N_177);
nand U1945 (N_1945,N_975,N_933);
nand U1946 (N_1946,N_292,N_447);
xnor U1947 (N_1947,N_763,N_208);
or U1948 (N_1948,N_405,N_438);
nand U1949 (N_1949,N_788,N_808);
or U1950 (N_1950,N_773,N_411);
or U1951 (N_1951,N_401,N_272);
nand U1952 (N_1952,N_619,N_974);
or U1953 (N_1953,N_721,N_657);
or U1954 (N_1954,N_194,N_528);
nor U1955 (N_1955,N_307,N_839);
and U1956 (N_1956,N_800,N_898);
nor U1957 (N_1957,N_541,N_150);
and U1958 (N_1958,N_346,N_177);
and U1959 (N_1959,N_838,N_144);
or U1960 (N_1960,N_159,N_574);
and U1961 (N_1961,N_133,N_57);
xnor U1962 (N_1962,N_720,N_910);
or U1963 (N_1963,N_837,N_279);
nand U1964 (N_1964,N_220,N_806);
or U1965 (N_1965,N_364,N_475);
and U1966 (N_1966,N_81,N_251);
nor U1967 (N_1967,N_938,N_814);
xnor U1968 (N_1968,N_942,N_239);
or U1969 (N_1969,N_755,N_367);
nor U1970 (N_1970,N_497,N_748);
nand U1971 (N_1971,N_863,N_741);
and U1972 (N_1972,N_928,N_614);
nor U1973 (N_1973,N_69,N_219);
and U1974 (N_1974,N_746,N_319);
and U1975 (N_1975,N_873,N_227);
nor U1976 (N_1976,N_790,N_54);
nor U1977 (N_1977,N_19,N_109);
or U1978 (N_1978,N_916,N_897);
and U1979 (N_1979,N_439,N_368);
xor U1980 (N_1980,N_545,N_865);
or U1981 (N_1981,N_782,N_394);
xor U1982 (N_1982,N_852,N_733);
or U1983 (N_1983,N_407,N_258);
or U1984 (N_1984,N_476,N_901);
nor U1985 (N_1985,N_62,N_715);
or U1986 (N_1986,N_556,N_917);
and U1987 (N_1987,N_858,N_941);
nor U1988 (N_1988,N_577,N_810);
and U1989 (N_1989,N_863,N_216);
or U1990 (N_1990,N_908,N_320);
or U1991 (N_1991,N_233,N_720);
nor U1992 (N_1992,N_666,N_629);
and U1993 (N_1993,N_122,N_753);
and U1994 (N_1994,N_173,N_421);
xor U1995 (N_1995,N_91,N_228);
nand U1996 (N_1996,N_805,N_852);
xor U1997 (N_1997,N_182,N_17);
nand U1998 (N_1998,N_801,N_699);
nand U1999 (N_1999,N_556,N_847);
nand U2000 (N_2000,N_1264,N_1136);
nand U2001 (N_2001,N_1344,N_1154);
or U2002 (N_2002,N_1823,N_1884);
nand U2003 (N_2003,N_1695,N_1503);
and U2004 (N_2004,N_1747,N_1453);
or U2005 (N_2005,N_1149,N_1245);
nand U2006 (N_2006,N_1458,N_1696);
or U2007 (N_2007,N_1253,N_1235);
nor U2008 (N_2008,N_1677,N_1815);
nor U2009 (N_2009,N_1929,N_1732);
and U2010 (N_2010,N_1090,N_1414);
and U2011 (N_2011,N_1988,N_1128);
nand U2012 (N_2012,N_1763,N_1442);
nor U2013 (N_2013,N_1200,N_1863);
nor U2014 (N_2014,N_1222,N_1326);
nand U2015 (N_2015,N_1980,N_1350);
nor U2016 (N_2016,N_1471,N_1457);
nand U2017 (N_2017,N_1361,N_1383);
or U2018 (N_2018,N_1179,N_1315);
or U2019 (N_2019,N_1436,N_1932);
xor U2020 (N_2020,N_1666,N_1964);
nor U2021 (N_2021,N_1752,N_1722);
nand U2022 (N_2022,N_1920,N_1827);
nand U2023 (N_2023,N_1196,N_1723);
nor U2024 (N_2024,N_1584,N_1277);
or U2025 (N_2025,N_1516,N_1117);
nand U2026 (N_2026,N_1492,N_1995);
nand U2027 (N_2027,N_1340,N_1889);
and U2028 (N_2028,N_1711,N_1989);
and U2029 (N_2029,N_1215,N_1699);
and U2030 (N_2030,N_1655,N_1586);
nand U2031 (N_2031,N_1690,N_1820);
or U2032 (N_2032,N_1505,N_1243);
nand U2033 (N_2033,N_1106,N_1712);
nor U2034 (N_2034,N_1892,N_1422);
nor U2035 (N_2035,N_1802,N_1318);
nand U2036 (N_2036,N_1204,N_1259);
nor U2037 (N_2037,N_1992,N_1119);
and U2038 (N_2038,N_1688,N_1596);
nor U2039 (N_2039,N_1103,N_1578);
nor U2040 (N_2040,N_1237,N_1770);
nor U2041 (N_2041,N_1267,N_1464);
and U2042 (N_2042,N_1911,N_1506);
and U2043 (N_2043,N_1956,N_1399);
xor U2044 (N_2044,N_1675,N_1330);
nand U2045 (N_2045,N_1319,N_1170);
and U2046 (N_2046,N_1285,N_1969);
nand U2047 (N_2047,N_1362,N_1073);
or U2048 (N_2048,N_1122,N_1841);
and U2049 (N_2049,N_1120,N_1633);
xnor U2050 (N_2050,N_1166,N_1062);
nor U2051 (N_2051,N_1926,N_1611);
nor U2052 (N_2052,N_1602,N_1782);
or U2053 (N_2053,N_1329,N_1490);
and U2054 (N_2054,N_1387,N_1757);
nor U2055 (N_2055,N_1412,N_1910);
nor U2056 (N_2056,N_1191,N_1931);
nor U2057 (N_2057,N_1298,N_1445);
xor U2058 (N_2058,N_1135,N_1908);
nand U2059 (N_2059,N_1208,N_1303);
nor U2060 (N_2060,N_1576,N_1023);
or U2061 (N_2061,N_1811,N_1451);
nor U2062 (N_2062,N_1067,N_1369);
and U2063 (N_2063,N_1323,N_1226);
and U2064 (N_2064,N_1255,N_1982);
nand U2065 (N_2065,N_1297,N_1801);
nor U2066 (N_2066,N_1526,N_1483);
nand U2067 (N_2067,N_1129,N_1877);
nand U2068 (N_2068,N_1685,N_1545);
or U2069 (N_2069,N_1052,N_1003);
nand U2070 (N_2070,N_1523,N_1580);
nor U2071 (N_2071,N_1496,N_1241);
nor U2072 (N_2072,N_1733,N_1554);
or U2073 (N_2073,N_1021,N_1086);
nor U2074 (N_2074,N_1089,N_1131);
and U2075 (N_2075,N_1017,N_1402);
nor U2076 (N_2076,N_1567,N_1831);
nand U2077 (N_2077,N_1941,N_1721);
nor U2078 (N_2078,N_1574,N_1477);
nor U2079 (N_2079,N_1797,N_1371);
nand U2080 (N_2080,N_1434,N_1391);
and U2081 (N_2081,N_1682,N_1439);
xnor U2082 (N_2082,N_1651,N_1702);
or U2083 (N_2083,N_1906,N_1985);
or U2084 (N_2084,N_1459,N_1251);
nand U2085 (N_2085,N_1172,N_1587);
and U2086 (N_2086,N_1001,N_1118);
or U2087 (N_2087,N_1869,N_1847);
nor U2088 (N_2088,N_1175,N_1948);
xor U2089 (N_2089,N_1799,N_1474);
xnor U2090 (N_2090,N_1798,N_1718);
nor U2091 (N_2091,N_1609,N_1991);
nand U2092 (N_2092,N_1978,N_1758);
nand U2093 (N_2093,N_1355,N_1654);
nand U2094 (N_2094,N_1463,N_1857);
or U2095 (N_2095,N_1337,N_1058);
nor U2096 (N_2096,N_1328,N_1614);
and U2097 (N_2097,N_1002,N_1977);
and U2098 (N_2098,N_1697,N_1376);
nand U2099 (N_2099,N_1787,N_1748);
nor U2100 (N_2100,N_1745,N_1449);
nor U2101 (N_2101,N_1683,N_1829);
and U2102 (N_2102,N_1937,N_1499);
or U2103 (N_2103,N_1384,N_1060);
nor U2104 (N_2104,N_1153,N_1138);
or U2105 (N_2105,N_1512,N_1261);
and U2106 (N_2106,N_1999,N_1854);
nor U2107 (N_2107,N_1377,N_1844);
nor U2108 (N_2108,N_1921,N_1312);
nor U2109 (N_2109,N_1148,N_1256);
or U2110 (N_2110,N_1856,N_1278);
nand U2111 (N_2111,N_1491,N_1364);
or U2112 (N_2112,N_1788,N_1342);
xor U2113 (N_2113,N_1380,N_1585);
xnor U2114 (N_2114,N_1821,N_1145);
nor U2115 (N_2115,N_1132,N_1552);
or U2116 (N_2116,N_1481,N_1600);
and U2117 (N_2117,N_1398,N_1053);
nor U2118 (N_2118,N_1033,N_1955);
or U2119 (N_2119,N_1944,N_1984);
nand U2120 (N_2120,N_1194,N_1431);
nand U2121 (N_2121,N_1368,N_1625);
nor U2122 (N_2122,N_1075,N_1227);
nand U2123 (N_2123,N_1216,N_1834);
nand U2124 (N_2124,N_1260,N_1054);
or U2125 (N_2125,N_1346,N_1959);
nor U2126 (N_2126,N_1700,N_1643);
or U2127 (N_2127,N_1411,N_1949);
nand U2128 (N_2128,N_1324,N_1167);
xor U2129 (N_2129,N_1236,N_1012);
xor U2130 (N_2130,N_1427,N_1000);
nor U2131 (N_2131,N_1206,N_1659);
nor U2132 (N_2132,N_1026,N_1538);
xnor U2133 (N_2133,N_1963,N_1645);
and U2134 (N_2134,N_1217,N_1565);
and U2135 (N_2135,N_1934,N_1307);
nor U2136 (N_2136,N_1727,N_1389);
nand U2137 (N_2137,N_1694,N_1852);
xor U2138 (N_2138,N_1497,N_1930);
nand U2139 (N_2139,N_1112,N_1905);
nor U2140 (N_2140,N_1108,N_1055);
or U2141 (N_2141,N_1846,N_1916);
and U2142 (N_2142,N_1967,N_1657);
nand U2143 (N_2143,N_1005,N_1562);
or U2144 (N_2144,N_1940,N_1192);
nor U2145 (N_2145,N_1169,N_1945);
and U2146 (N_2146,N_1410,N_1593);
or U2147 (N_2147,N_1348,N_1031);
xor U2148 (N_2148,N_1317,N_1936);
and U2149 (N_2149,N_1238,N_1818);
and U2150 (N_2150,N_1165,N_1246);
nor U2151 (N_2151,N_1443,N_1724);
nand U2152 (N_2152,N_1358,N_1363);
nand U2153 (N_2153,N_1189,N_1147);
nand U2154 (N_2154,N_1366,N_1603);
or U2155 (N_2155,N_1302,N_1095);
or U2156 (N_2156,N_1468,N_1656);
nor U2157 (N_2157,N_1019,N_1294);
or U2158 (N_2158,N_1572,N_1740);
xnor U2159 (N_2159,N_1601,N_1873);
nor U2160 (N_2160,N_1311,N_1527);
nor U2161 (N_2161,N_1343,N_1452);
or U2162 (N_2162,N_1310,N_1824);
or U2163 (N_2163,N_1197,N_1791);
or U2164 (N_2164,N_1960,N_1163);
xnor U2165 (N_2165,N_1401,N_1855);
xnor U2166 (N_2166,N_1731,N_1726);
nor U2167 (N_2167,N_1088,N_1141);
and U2168 (N_2168,N_1705,N_1515);
nor U2169 (N_2169,N_1007,N_1093);
and U2170 (N_2170,N_1622,N_1071);
nand U2171 (N_2171,N_1152,N_1157);
xnor U2172 (N_2172,N_1182,N_1299);
and U2173 (N_2173,N_1777,N_1283);
or U2174 (N_2174,N_1478,N_1063);
and U2175 (N_2175,N_1164,N_1664);
and U2176 (N_2176,N_1385,N_1448);
nand U2177 (N_2177,N_1848,N_1306);
nor U2178 (N_2178,N_1804,N_1687);
nor U2179 (N_2179,N_1495,N_1134);
xor U2180 (N_2180,N_1010,N_1072);
and U2181 (N_2181,N_1529,N_1270);
or U2182 (N_2182,N_1094,N_1456);
nor U2183 (N_2183,N_1274,N_1279);
or U2184 (N_2184,N_1974,N_1943);
and U2185 (N_2185,N_1714,N_1321);
nand U2186 (N_2186,N_1590,N_1566);
nor U2187 (N_2187,N_1997,N_1866);
or U2188 (N_2188,N_1907,N_1043);
or U2189 (N_2189,N_1900,N_1785);
nor U2190 (N_2190,N_1742,N_1830);
xor U2191 (N_2191,N_1653,N_1105);
and U2192 (N_2192,N_1588,N_1313);
or U2193 (N_2193,N_1500,N_1524);
or U2194 (N_2194,N_1560,N_1379);
nand U2195 (N_2195,N_1883,N_1314);
nor U2196 (N_2196,N_1465,N_1864);
nand U2197 (N_2197,N_1660,N_1082);
and U2198 (N_2198,N_1915,N_1594);
nand U2199 (N_2199,N_1455,N_1564);
or U2200 (N_2200,N_1473,N_1553);
xnor U2201 (N_2201,N_1887,N_1417);
and U2202 (N_2202,N_1498,N_1607);
nand U2203 (N_2203,N_1973,N_1339);
or U2204 (N_2204,N_1004,N_1466);
or U2205 (N_2205,N_1382,N_1766);
and U2206 (N_2206,N_1015,N_1142);
nor U2207 (N_2207,N_1640,N_1998);
and U2208 (N_2208,N_1140,N_1174);
or U2209 (N_2209,N_1316,N_1901);
or U2210 (N_2210,N_1924,N_1835);
nor U2211 (N_2211,N_1220,N_1667);
or U2212 (N_2212,N_1867,N_1796);
or U2213 (N_2213,N_1396,N_1130);
or U2214 (N_2214,N_1234,N_1333);
nor U2215 (N_2215,N_1751,N_1244);
and U2216 (N_2216,N_1897,N_1469);
and U2217 (N_2217,N_1680,N_1247);
or U2218 (N_2218,N_1292,N_1239);
and U2219 (N_2219,N_1504,N_1305);
or U2220 (N_2220,N_1909,N_1703);
nor U2221 (N_2221,N_1104,N_1780);
or U2222 (N_2222,N_1853,N_1263);
and U2223 (N_2223,N_1630,N_1738);
nor U2224 (N_2224,N_1741,N_1430);
nor U2225 (N_2225,N_1707,N_1405);
nand U2226 (N_2226,N_1617,N_1919);
or U2227 (N_2227,N_1177,N_1535);
nand U2228 (N_2228,N_1444,N_1893);
xor U2229 (N_2229,N_1137,N_1254);
and U2230 (N_2230,N_1860,N_1493);
xor U2231 (N_2231,N_1485,N_1626);
or U2232 (N_2232,N_1352,N_1281);
xnor U2233 (N_2233,N_1461,N_1024);
xor U2234 (N_2234,N_1390,N_1440);
nor U2235 (N_2235,N_1735,N_1301);
and U2236 (N_2236,N_1533,N_1115);
nand U2237 (N_2237,N_1610,N_1953);
or U2238 (N_2238,N_1833,N_1794);
and U2239 (N_2239,N_1813,N_1544);
or U2240 (N_2240,N_1879,N_1331);
nor U2241 (N_2241,N_1290,N_1096);
and U2242 (N_2242,N_1968,N_1193);
and U2243 (N_2243,N_1224,N_1064);
nor U2244 (N_2244,N_1265,N_1536);
nor U2245 (N_2245,N_1761,N_1036);
and U2246 (N_2246,N_1708,N_1039);
and U2247 (N_2247,N_1756,N_1408);
or U2248 (N_2248,N_1904,N_1876);
or U2249 (N_2249,N_1028,N_1151);
and U2250 (N_2250,N_1304,N_1139);
or U2251 (N_2251,N_1836,N_1472);
nor U2252 (N_2252,N_1765,N_1037);
and U2253 (N_2253,N_1228,N_1575);
or U2254 (N_2254,N_1240,N_1400);
nand U2255 (N_2255,N_1684,N_1979);
nand U2256 (N_2256,N_1420,N_1962);
nor U2257 (N_2257,N_1933,N_1816);
nand U2258 (N_2258,N_1706,N_1532);
nand U2259 (N_2259,N_1693,N_1808);
or U2260 (N_2260,N_1098,N_1334);
or U2261 (N_2261,N_1276,N_1789);
or U2262 (N_2262,N_1038,N_1636);
nand U2263 (N_2263,N_1649,N_1746);
or U2264 (N_2264,N_1365,N_1522);
nand U2265 (N_2265,N_1143,N_1713);
nand U2266 (N_2266,N_1599,N_1604);
nor U2267 (N_2267,N_1009,N_1729);
or U2268 (N_2268,N_1672,N_1212);
nand U2269 (N_2269,N_1262,N_1386);
nand U2270 (N_2270,N_1013,N_1958);
nor U2271 (N_2271,N_1309,N_1403);
xor U2272 (N_2272,N_1100,N_1205);
nor U2273 (N_2273,N_1187,N_1547);
nand U2274 (N_2274,N_1034,N_1381);
nor U2275 (N_2275,N_1620,N_1102);
or U2276 (N_2276,N_1885,N_1595);
and U2277 (N_2277,N_1671,N_1429);
and U2278 (N_2278,N_1537,N_1233);
or U2279 (N_2279,N_1838,N_1198);
nand U2280 (N_2280,N_1819,N_1083);
nor U2281 (N_2281,N_1810,N_1156);
xor U2282 (N_2282,N_1983,N_1437);
and U2283 (N_2283,N_1210,N_1395);
xor U2284 (N_2284,N_1209,N_1759);
and U2285 (N_2285,N_1016,N_1881);
and U2286 (N_2286,N_1786,N_1938);
nand U2287 (N_2287,N_1616,N_1511);
nand U2288 (N_2288,N_1242,N_1519);
and U2289 (N_2289,N_1621,N_1608);
xnor U2290 (N_2290,N_1639,N_1704);
xnor U2291 (N_2291,N_1635,N_1744);
or U2292 (N_2292,N_1993,N_1928);
nand U2293 (N_2293,N_1011,N_1902);
or U2294 (N_2294,N_1423,N_1618);
nand U2295 (N_2295,N_1406,N_1202);
nor U2296 (N_2296,N_1338,N_1716);
and U2297 (N_2297,N_1539,N_1289);
or U2298 (N_2298,N_1415,N_1336);
nor U2299 (N_2299,N_1698,N_1895);
and U2300 (N_2300,N_1849,N_1479);
nand U2301 (N_2301,N_1950,N_1046);
nor U2302 (N_2302,N_1870,N_1433);
and U2303 (N_2303,N_1571,N_1606);
nor U2304 (N_2304,N_1397,N_1300);
and U2305 (N_2305,N_1475,N_1840);
nor U2306 (N_2306,N_1040,N_1917);
nand U2307 (N_2307,N_1032,N_1619);
and U2308 (N_2308,N_1581,N_1470);
nor U2309 (N_2309,N_1087,N_1689);
xnor U2310 (N_2310,N_1809,N_1951);
nor U2311 (N_2311,N_1665,N_1085);
and U2312 (N_2312,N_1668,N_1612);
nand U2313 (N_2313,N_1644,N_1772);
nor U2314 (N_2314,N_1996,N_1513);
and U2315 (N_2315,N_1543,N_1125);
and U2316 (N_2316,N_1378,N_1990);
or U2317 (N_2317,N_1678,N_1308);
nand U2318 (N_2318,N_1550,N_1124);
and U2319 (N_2319,N_1425,N_1832);
and U2320 (N_2320,N_1070,N_1435);
nor U2321 (N_2321,N_1520,N_1441);
or U2322 (N_2322,N_1710,N_1632);
or U2323 (N_2323,N_1720,N_1476);
or U2324 (N_2324,N_1923,N_1896);
or U2325 (N_2325,N_1027,N_1322);
and U2326 (N_2326,N_1570,N_1269);
or U2327 (N_2327,N_1822,N_1669);
xnor U2328 (N_2328,N_1284,N_1935);
or U2329 (N_2329,N_1426,N_1627);
and U2330 (N_2330,N_1252,N_1681);
nor U2331 (N_2331,N_1502,N_1341);
nand U2332 (N_2332,N_1190,N_1375);
nor U2333 (N_2333,N_1486,N_1514);
nor U2334 (N_2334,N_1195,N_1661);
nand U2335 (N_2335,N_1020,N_1691);
nand U2336 (N_2336,N_1061,N_1859);
nand U2337 (N_2337,N_1845,N_1354);
and U2338 (N_2338,N_1737,N_1219);
or U2339 (N_2339,N_1784,N_1501);
and U2340 (N_2340,N_1159,N_1325);
and U2341 (N_2341,N_1035,N_1771);
xor U2342 (N_2342,N_1109,N_1409);
or U2343 (N_2343,N_1050,N_1029);
or U2344 (N_2344,N_1629,N_1760);
and U2345 (N_2345,N_1257,N_1987);
nor U2346 (N_2346,N_1871,N_1663);
or U2347 (N_2347,N_1957,N_1767);
or U2348 (N_2348,N_1510,N_1872);
and U2349 (N_2349,N_1356,N_1248);
nand U2350 (N_2350,N_1986,N_1807);
nor U2351 (N_2351,N_1332,N_1946);
nand U2352 (N_2352,N_1286,N_1814);
xnor U2353 (N_2353,N_1432,N_1994);
and U2354 (N_2354,N_1018,N_1843);
or U2355 (N_2355,N_1373,N_1184);
nand U2356 (N_2356,N_1223,N_1008);
and U2357 (N_2357,N_1803,N_1898);
nor U2358 (N_2358,N_1764,N_1558);
nand U2359 (N_2359,N_1970,N_1976);
or U2360 (N_2360,N_1826,N_1878);
and U2361 (N_2361,N_1351,N_1280);
and U2362 (N_2362,N_1173,N_1388);
xnor U2363 (N_2363,N_1428,N_1250);
nor U2364 (N_2364,N_1066,N_1800);
nor U2365 (N_2365,N_1111,N_1779);
and U2366 (N_2366,N_1273,N_1939);
nand U2367 (N_2367,N_1418,N_1899);
nand U2368 (N_2368,N_1882,N_1068);
and U2369 (N_2369,N_1851,N_1296);
or U2370 (N_2370,N_1171,N_1769);
nand U2371 (N_2371,N_1113,N_1709);
or U2372 (N_2372,N_1230,N_1912);
and U2373 (N_2373,N_1631,N_1180);
and U2374 (N_2374,N_1730,N_1942);
and U2375 (N_2375,N_1890,N_1214);
and U2376 (N_2376,N_1692,N_1293);
xnor U2377 (N_2377,N_1488,N_1719);
nor U2378 (N_2378,N_1271,N_1868);
and U2379 (N_2379,N_1282,N_1370);
nor U2380 (N_2380,N_1345,N_1874);
nand U2381 (N_2381,N_1728,N_1218);
or U2382 (N_2382,N_1817,N_1144);
xnor U2383 (N_2383,N_1837,N_1161);
nand U2384 (N_2384,N_1679,N_1446);
or U2385 (N_2385,N_1101,N_1521);
nand U2386 (N_2386,N_1894,N_1743);
or U2387 (N_2387,N_1842,N_1628);
or U2388 (N_2388,N_1487,N_1918);
or U2389 (N_2389,N_1121,N_1839);
xor U2390 (N_2390,N_1828,N_1762);
nand U2391 (N_2391,N_1518,N_1126);
nand U2392 (N_2392,N_1715,N_1123);
or U2393 (N_2393,N_1127,N_1971);
and U2394 (N_2394,N_1773,N_1107);
or U2395 (N_2395,N_1952,N_1181);
nand U2396 (N_2396,N_1078,N_1221);
and U2397 (N_2397,N_1641,N_1875);
or U2398 (N_2398,N_1042,N_1006);
nand U2399 (N_2399,N_1790,N_1701);
xor U2400 (N_2400,N_1579,N_1110);
or U2401 (N_2401,N_1349,N_1965);
and U2402 (N_2402,N_1288,N_1025);
or U2403 (N_2403,N_1676,N_1438);
xor U2404 (N_2404,N_1793,N_1229);
nor U2405 (N_2405,N_1534,N_1557);
xnor U2406 (N_2406,N_1494,N_1768);
nor U2407 (N_2407,N_1650,N_1638);
or U2408 (N_2408,N_1615,N_1850);
nand U2409 (N_2409,N_1199,N_1091);
nand U2410 (N_2410,N_1981,N_1749);
nor U2411 (N_2411,N_1597,N_1392);
nor U2412 (N_2412,N_1739,N_1542);
or U2413 (N_2413,N_1858,N_1213);
or U2414 (N_2414,N_1972,N_1582);
nand U2415 (N_2415,N_1407,N_1736);
and U2416 (N_2416,N_1734,N_1569);
and U2417 (N_2417,N_1421,N_1048);
and U2418 (N_2418,N_1022,N_1394);
nor U2419 (N_2419,N_1658,N_1642);
nor U2420 (N_2420,N_1605,N_1416);
xnor U2421 (N_2421,N_1045,N_1168);
nand U2422 (N_2422,N_1903,N_1158);
or U2423 (N_2423,N_1914,N_1862);
or U2424 (N_2424,N_1374,N_1489);
or U2425 (N_2425,N_1335,N_1162);
nor U2426 (N_2426,N_1133,N_1778);
nand U2427 (N_2427,N_1556,N_1275);
nor U2428 (N_2428,N_1755,N_1674);
nand U2429 (N_2429,N_1065,N_1372);
nor U2430 (N_2430,N_1367,N_1116);
nor U2431 (N_2431,N_1913,N_1551);
nand U2432 (N_2432,N_1272,N_1795);
nor U2433 (N_2433,N_1546,N_1750);
xor U2434 (N_2434,N_1084,N_1188);
or U2435 (N_2435,N_1865,N_1531);
or U2436 (N_2436,N_1077,N_1686);
xor U2437 (N_2437,N_1076,N_1753);
or U2438 (N_2438,N_1563,N_1225);
or U2439 (N_2439,N_1646,N_1652);
and U2440 (N_2440,N_1207,N_1092);
xor U2441 (N_2441,N_1266,N_1647);
xnor U2442 (N_2442,N_1327,N_1781);
nand U2443 (N_2443,N_1249,N_1583);
and U2444 (N_2444,N_1482,N_1540);
nor U2445 (N_2445,N_1555,N_1662);
nand U2446 (N_2446,N_1961,N_1648);
xnor U2447 (N_2447,N_1484,N_1975);
or U2448 (N_2448,N_1454,N_1549);
and U2449 (N_2449,N_1447,N_1231);
nor U2450 (N_2450,N_1462,N_1393);
nand U2451 (N_2451,N_1203,N_1783);
nor U2452 (N_2452,N_1509,N_1360);
nor U2453 (N_2453,N_1568,N_1186);
nand U2454 (N_2454,N_1725,N_1947);
nor U2455 (N_2455,N_1888,N_1861);
xor U2456 (N_2456,N_1480,N_1424);
and U2457 (N_2457,N_1891,N_1577);
nor U2458 (N_2458,N_1069,N_1954);
nor U2459 (N_2459,N_1922,N_1927);
nand U2460 (N_2460,N_1886,N_1591);
nand U2461 (N_2461,N_1232,N_1211);
nor U2462 (N_2462,N_1258,N_1041);
nand U2463 (N_2463,N_1925,N_1057);
or U2464 (N_2464,N_1178,N_1030);
nand U2465 (N_2465,N_1051,N_1776);
or U2466 (N_2466,N_1623,N_1775);
or U2467 (N_2467,N_1047,N_1097);
nor U2468 (N_2468,N_1201,N_1613);
or U2469 (N_2469,N_1637,N_1080);
nor U2470 (N_2470,N_1825,N_1268);
nor U2471 (N_2471,N_1359,N_1413);
nand U2472 (N_2472,N_1357,N_1673);
nand U2473 (N_2473,N_1320,N_1508);
nor U2474 (N_2474,N_1966,N_1291);
nor U2475 (N_2475,N_1081,N_1805);
or U2476 (N_2476,N_1049,N_1056);
nor U2477 (N_2477,N_1598,N_1561);
nand U2478 (N_2478,N_1347,N_1517);
or U2479 (N_2479,N_1146,N_1287);
xor U2480 (N_2480,N_1754,N_1634);
or U2481 (N_2481,N_1589,N_1507);
nand U2482 (N_2482,N_1548,N_1044);
or U2483 (N_2483,N_1670,N_1155);
nand U2484 (N_2484,N_1160,N_1559);
nor U2485 (N_2485,N_1150,N_1450);
nand U2486 (N_2486,N_1530,N_1717);
and U2487 (N_2487,N_1099,N_1880);
and U2488 (N_2488,N_1812,N_1528);
nor U2489 (N_2489,N_1541,N_1059);
nor U2490 (N_2490,N_1525,N_1419);
and U2491 (N_2491,N_1806,N_1074);
or U2492 (N_2492,N_1460,N_1792);
and U2493 (N_2493,N_1467,N_1573);
or U2494 (N_2494,N_1185,N_1176);
and U2495 (N_2495,N_1404,N_1295);
nor U2496 (N_2496,N_1014,N_1079);
xnor U2497 (N_2497,N_1624,N_1114);
or U2498 (N_2498,N_1183,N_1774);
or U2499 (N_2499,N_1592,N_1353);
nor U2500 (N_2500,N_1200,N_1492);
nand U2501 (N_2501,N_1678,N_1878);
and U2502 (N_2502,N_1394,N_1726);
or U2503 (N_2503,N_1232,N_1508);
nor U2504 (N_2504,N_1471,N_1319);
and U2505 (N_2505,N_1845,N_1657);
or U2506 (N_2506,N_1368,N_1061);
and U2507 (N_2507,N_1984,N_1052);
nand U2508 (N_2508,N_1022,N_1091);
and U2509 (N_2509,N_1657,N_1461);
nand U2510 (N_2510,N_1187,N_1317);
or U2511 (N_2511,N_1455,N_1556);
xnor U2512 (N_2512,N_1286,N_1850);
and U2513 (N_2513,N_1334,N_1308);
nand U2514 (N_2514,N_1984,N_1011);
and U2515 (N_2515,N_1089,N_1121);
nand U2516 (N_2516,N_1256,N_1362);
nand U2517 (N_2517,N_1563,N_1603);
and U2518 (N_2518,N_1345,N_1859);
and U2519 (N_2519,N_1764,N_1740);
or U2520 (N_2520,N_1761,N_1729);
and U2521 (N_2521,N_1925,N_1832);
and U2522 (N_2522,N_1255,N_1487);
nand U2523 (N_2523,N_1570,N_1373);
and U2524 (N_2524,N_1926,N_1620);
nor U2525 (N_2525,N_1789,N_1734);
or U2526 (N_2526,N_1948,N_1646);
and U2527 (N_2527,N_1575,N_1257);
nand U2528 (N_2528,N_1224,N_1589);
or U2529 (N_2529,N_1356,N_1000);
nand U2530 (N_2530,N_1925,N_1302);
and U2531 (N_2531,N_1944,N_1974);
or U2532 (N_2532,N_1883,N_1255);
nor U2533 (N_2533,N_1151,N_1944);
nor U2534 (N_2534,N_1783,N_1579);
or U2535 (N_2535,N_1227,N_1320);
and U2536 (N_2536,N_1965,N_1647);
and U2537 (N_2537,N_1036,N_1529);
and U2538 (N_2538,N_1697,N_1492);
xnor U2539 (N_2539,N_1222,N_1640);
or U2540 (N_2540,N_1888,N_1356);
or U2541 (N_2541,N_1989,N_1791);
or U2542 (N_2542,N_1153,N_1320);
or U2543 (N_2543,N_1328,N_1581);
nand U2544 (N_2544,N_1113,N_1753);
nor U2545 (N_2545,N_1441,N_1118);
xnor U2546 (N_2546,N_1733,N_1878);
xnor U2547 (N_2547,N_1702,N_1340);
and U2548 (N_2548,N_1831,N_1461);
and U2549 (N_2549,N_1876,N_1337);
nor U2550 (N_2550,N_1733,N_1421);
or U2551 (N_2551,N_1267,N_1618);
and U2552 (N_2552,N_1447,N_1263);
nor U2553 (N_2553,N_1342,N_1127);
or U2554 (N_2554,N_1956,N_1525);
nor U2555 (N_2555,N_1740,N_1817);
nor U2556 (N_2556,N_1916,N_1142);
and U2557 (N_2557,N_1710,N_1559);
nor U2558 (N_2558,N_1562,N_1102);
or U2559 (N_2559,N_1664,N_1077);
nor U2560 (N_2560,N_1435,N_1587);
xnor U2561 (N_2561,N_1736,N_1638);
and U2562 (N_2562,N_1876,N_1774);
xor U2563 (N_2563,N_1080,N_1680);
or U2564 (N_2564,N_1498,N_1297);
xnor U2565 (N_2565,N_1677,N_1316);
and U2566 (N_2566,N_1844,N_1531);
nand U2567 (N_2567,N_1075,N_1014);
or U2568 (N_2568,N_1465,N_1694);
nand U2569 (N_2569,N_1207,N_1123);
nand U2570 (N_2570,N_1927,N_1025);
or U2571 (N_2571,N_1536,N_1160);
xnor U2572 (N_2572,N_1022,N_1743);
nand U2573 (N_2573,N_1636,N_1383);
nor U2574 (N_2574,N_1612,N_1170);
nor U2575 (N_2575,N_1113,N_1935);
nor U2576 (N_2576,N_1615,N_1221);
or U2577 (N_2577,N_1321,N_1820);
nor U2578 (N_2578,N_1970,N_1084);
nand U2579 (N_2579,N_1795,N_1769);
nand U2580 (N_2580,N_1983,N_1328);
or U2581 (N_2581,N_1182,N_1854);
and U2582 (N_2582,N_1494,N_1543);
and U2583 (N_2583,N_1046,N_1188);
nand U2584 (N_2584,N_1336,N_1699);
nand U2585 (N_2585,N_1834,N_1142);
xnor U2586 (N_2586,N_1181,N_1475);
nor U2587 (N_2587,N_1922,N_1437);
xor U2588 (N_2588,N_1420,N_1562);
or U2589 (N_2589,N_1780,N_1971);
nor U2590 (N_2590,N_1553,N_1076);
nand U2591 (N_2591,N_1686,N_1290);
nand U2592 (N_2592,N_1845,N_1745);
nand U2593 (N_2593,N_1574,N_1231);
nor U2594 (N_2594,N_1344,N_1198);
or U2595 (N_2595,N_1418,N_1074);
or U2596 (N_2596,N_1859,N_1011);
xor U2597 (N_2597,N_1534,N_1870);
nor U2598 (N_2598,N_1876,N_1098);
and U2599 (N_2599,N_1603,N_1802);
and U2600 (N_2600,N_1188,N_1956);
nor U2601 (N_2601,N_1521,N_1391);
or U2602 (N_2602,N_1761,N_1969);
nor U2603 (N_2603,N_1581,N_1491);
nor U2604 (N_2604,N_1314,N_1610);
nor U2605 (N_2605,N_1587,N_1084);
nand U2606 (N_2606,N_1990,N_1711);
nand U2607 (N_2607,N_1950,N_1819);
or U2608 (N_2608,N_1988,N_1445);
or U2609 (N_2609,N_1588,N_1556);
or U2610 (N_2610,N_1680,N_1419);
nor U2611 (N_2611,N_1179,N_1752);
nand U2612 (N_2612,N_1873,N_1501);
or U2613 (N_2613,N_1425,N_1223);
xor U2614 (N_2614,N_1046,N_1330);
nand U2615 (N_2615,N_1997,N_1889);
or U2616 (N_2616,N_1448,N_1157);
and U2617 (N_2617,N_1103,N_1569);
or U2618 (N_2618,N_1528,N_1852);
or U2619 (N_2619,N_1090,N_1272);
and U2620 (N_2620,N_1004,N_1107);
and U2621 (N_2621,N_1864,N_1106);
and U2622 (N_2622,N_1215,N_1194);
nor U2623 (N_2623,N_1952,N_1426);
xor U2624 (N_2624,N_1426,N_1835);
nor U2625 (N_2625,N_1038,N_1191);
nor U2626 (N_2626,N_1266,N_1830);
and U2627 (N_2627,N_1282,N_1854);
and U2628 (N_2628,N_1096,N_1671);
or U2629 (N_2629,N_1687,N_1214);
or U2630 (N_2630,N_1917,N_1424);
or U2631 (N_2631,N_1829,N_1909);
or U2632 (N_2632,N_1500,N_1309);
nor U2633 (N_2633,N_1744,N_1408);
nor U2634 (N_2634,N_1635,N_1946);
nor U2635 (N_2635,N_1376,N_1622);
nor U2636 (N_2636,N_1074,N_1025);
nor U2637 (N_2637,N_1064,N_1519);
xor U2638 (N_2638,N_1868,N_1334);
nand U2639 (N_2639,N_1796,N_1573);
and U2640 (N_2640,N_1628,N_1849);
or U2641 (N_2641,N_1240,N_1663);
or U2642 (N_2642,N_1758,N_1699);
nor U2643 (N_2643,N_1831,N_1015);
nor U2644 (N_2644,N_1929,N_1299);
nor U2645 (N_2645,N_1532,N_1277);
nand U2646 (N_2646,N_1610,N_1697);
or U2647 (N_2647,N_1317,N_1824);
nand U2648 (N_2648,N_1597,N_1593);
or U2649 (N_2649,N_1566,N_1261);
nand U2650 (N_2650,N_1389,N_1173);
or U2651 (N_2651,N_1055,N_1900);
nor U2652 (N_2652,N_1023,N_1474);
or U2653 (N_2653,N_1853,N_1073);
or U2654 (N_2654,N_1974,N_1568);
and U2655 (N_2655,N_1385,N_1806);
and U2656 (N_2656,N_1481,N_1332);
nand U2657 (N_2657,N_1377,N_1533);
or U2658 (N_2658,N_1480,N_1086);
xor U2659 (N_2659,N_1545,N_1503);
nor U2660 (N_2660,N_1046,N_1345);
or U2661 (N_2661,N_1872,N_1344);
or U2662 (N_2662,N_1293,N_1899);
xnor U2663 (N_2663,N_1156,N_1740);
and U2664 (N_2664,N_1459,N_1472);
and U2665 (N_2665,N_1480,N_1033);
and U2666 (N_2666,N_1394,N_1473);
nand U2667 (N_2667,N_1174,N_1888);
and U2668 (N_2668,N_1563,N_1730);
and U2669 (N_2669,N_1003,N_1074);
and U2670 (N_2670,N_1852,N_1518);
and U2671 (N_2671,N_1519,N_1409);
xor U2672 (N_2672,N_1045,N_1101);
nor U2673 (N_2673,N_1792,N_1321);
xnor U2674 (N_2674,N_1997,N_1419);
nand U2675 (N_2675,N_1760,N_1428);
nor U2676 (N_2676,N_1828,N_1419);
nand U2677 (N_2677,N_1130,N_1577);
nor U2678 (N_2678,N_1872,N_1259);
nor U2679 (N_2679,N_1593,N_1937);
nor U2680 (N_2680,N_1321,N_1188);
or U2681 (N_2681,N_1732,N_1738);
nand U2682 (N_2682,N_1245,N_1659);
and U2683 (N_2683,N_1618,N_1234);
nand U2684 (N_2684,N_1259,N_1923);
and U2685 (N_2685,N_1368,N_1127);
or U2686 (N_2686,N_1074,N_1239);
and U2687 (N_2687,N_1823,N_1662);
xnor U2688 (N_2688,N_1988,N_1793);
and U2689 (N_2689,N_1902,N_1101);
nand U2690 (N_2690,N_1469,N_1899);
nor U2691 (N_2691,N_1463,N_1275);
nor U2692 (N_2692,N_1172,N_1614);
nor U2693 (N_2693,N_1323,N_1767);
xor U2694 (N_2694,N_1899,N_1902);
nor U2695 (N_2695,N_1974,N_1475);
nand U2696 (N_2696,N_1169,N_1918);
and U2697 (N_2697,N_1218,N_1088);
and U2698 (N_2698,N_1662,N_1034);
xnor U2699 (N_2699,N_1679,N_1201);
and U2700 (N_2700,N_1589,N_1761);
nor U2701 (N_2701,N_1344,N_1327);
nor U2702 (N_2702,N_1853,N_1181);
or U2703 (N_2703,N_1327,N_1322);
xnor U2704 (N_2704,N_1623,N_1265);
nor U2705 (N_2705,N_1058,N_1624);
or U2706 (N_2706,N_1789,N_1094);
or U2707 (N_2707,N_1941,N_1041);
and U2708 (N_2708,N_1556,N_1682);
nor U2709 (N_2709,N_1452,N_1832);
or U2710 (N_2710,N_1557,N_1400);
xnor U2711 (N_2711,N_1062,N_1413);
and U2712 (N_2712,N_1024,N_1143);
or U2713 (N_2713,N_1718,N_1772);
or U2714 (N_2714,N_1724,N_1058);
and U2715 (N_2715,N_1850,N_1341);
or U2716 (N_2716,N_1604,N_1497);
nor U2717 (N_2717,N_1507,N_1085);
nand U2718 (N_2718,N_1803,N_1255);
nand U2719 (N_2719,N_1463,N_1297);
nand U2720 (N_2720,N_1212,N_1705);
xor U2721 (N_2721,N_1024,N_1781);
or U2722 (N_2722,N_1432,N_1259);
xnor U2723 (N_2723,N_1812,N_1468);
nor U2724 (N_2724,N_1682,N_1836);
nand U2725 (N_2725,N_1976,N_1499);
or U2726 (N_2726,N_1123,N_1080);
or U2727 (N_2727,N_1123,N_1766);
xor U2728 (N_2728,N_1089,N_1884);
and U2729 (N_2729,N_1388,N_1573);
and U2730 (N_2730,N_1315,N_1430);
and U2731 (N_2731,N_1489,N_1781);
and U2732 (N_2732,N_1860,N_1852);
xnor U2733 (N_2733,N_1471,N_1222);
xor U2734 (N_2734,N_1779,N_1051);
and U2735 (N_2735,N_1811,N_1244);
nand U2736 (N_2736,N_1241,N_1300);
xor U2737 (N_2737,N_1494,N_1941);
or U2738 (N_2738,N_1982,N_1399);
nor U2739 (N_2739,N_1839,N_1772);
nand U2740 (N_2740,N_1195,N_1135);
xnor U2741 (N_2741,N_1199,N_1842);
nand U2742 (N_2742,N_1731,N_1985);
or U2743 (N_2743,N_1852,N_1373);
and U2744 (N_2744,N_1571,N_1032);
nor U2745 (N_2745,N_1415,N_1222);
xor U2746 (N_2746,N_1338,N_1859);
and U2747 (N_2747,N_1020,N_1897);
nor U2748 (N_2748,N_1995,N_1897);
xor U2749 (N_2749,N_1920,N_1117);
nand U2750 (N_2750,N_1240,N_1221);
nand U2751 (N_2751,N_1762,N_1920);
or U2752 (N_2752,N_1240,N_1557);
and U2753 (N_2753,N_1502,N_1102);
nor U2754 (N_2754,N_1008,N_1279);
nand U2755 (N_2755,N_1291,N_1078);
and U2756 (N_2756,N_1288,N_1066);
or U2757 (N_2757,N_1461,N_1136);
nand U2758 (N_2758,N_1080,N_1056);
nand U2759 (N_2759,N_1849,N_1092);
xor U2760 (N_2760,N_1010,N_1577);
and U2761 (N_2761,N_1522,N_1768);
xnor U2762 (N_2762,N_1362,N_1979);
or U2763 (N_2763,N_1940,N_1663);
or U2764 (N_2764,N_1197,N_1980);
nor U2765 (N_2765,N_1143,N_1828);
and U2766 (N_2766,N_1686,N_1895);
and U2767 (N_2767,N_1591,N_1191);
nor U2768 (N_2768,N_1649,N_1308);
nand U2769 (N_2769,N_1683,N_1455);
and U2770 (N_2770,N_1860,N_1835);
or U2771 (N_2771,N_1511,N_1332);
and U2772 (N_2772,N_1090,N_1888);
or U2773 (N_2773,N_1205,N_1936);
nor U2774 (N_2774,N_1160,N_1817);
nor U2775 (N_2775,N_1248,N_1847);
xor U2776 (N_2776,N_1874,N_1736);
nand U2777 (N_2777,N_1170,N_1905);
or U2778 (N_2778,N_1022,N_1641);
and U2779 (N_2779,N_1406,N_1362);
and U2780 (N_2780,N_1856,N_1653);
nand U2781 (N_2781,N_1219,N_1686);
nor U2782 (N_2782,N_1851,N_1361);
and U2783 (N_2783,N_1501,N_1175);
and U2784 (N_2784,N_1256,N_1666);
nand U2785 (N_2785,N_1649,N_1984);
nor U2786 (N_2786,N_1979,N_1284);
or U2787 (N_2787,N_1711,N_1487);
nand U2788 (N_2788,N_1761,N_1804);
nand U2789 (N_2789,N_1409,N_1886);
and U2790 (N_2790,N_1248,N_1601);
or U2791 (N_2791,N_1215,N_1318);
and U2792 (N_2792,N_1984,N_1267);
or U2793 (N_2793,N_1436,N_1476);
and U2794 (N_2794,N_1302,N_1727);
xor U2795 (N_2795,N_1998,N_1499);
nand U2796 (N_2796,N_1002,N_1786);
xor U2797 (N_2797,N_1429,N_1229);
or U2798 (N_2798,N_1582,N_1861);
nand U2799 (N_2799,N_1055,N_1715);
nand U2800 (N_2800,N_1346,N_1785);
nor U2801 (N_2801,N_1419,N_1881);
xnor U2802 (N_2802,N_1402,N_1656);
or U2803 (N_2803,N_1302,N_1900);
or U2804 (N_2804,N_1693,N_1676);
nand U2805 (N_2805,N_1824,N_1657);
or U2806 (N_2806,N_1832,N_1196);
xnor U2807 (N_2807,N_1564,N_1304);
nand U2808 (N_2808,N_1921,N_1994);
and U2809 (N_2809,N_1549,N_1933);
or U2810 (N_2810,N_1197,N_1637);
xor U2811 (N_2811,N_1579,N_1106);
xor U2812 (N_2812,N_1486,N_1005);
nor U2813 (N_2813,N_1818,N_1206);
and U2814 (N_2814,N_1508,N_1854);
and U2815 (N_2815,N_1114,N_1294);
nor U2816 (N_2816,N_1377,N_1564);
nor U2817 (N_2817,N_1282,N_1425);
nand U2818 (N_2818,N_1798,N_1636);
nor U2819 (N_2819,N_1510,N_1633);
or U2820 (N_2820,N_1732,N_1062);
nor U2821 (N_2821,N_1462,N_1797);
or U2822 (N_2822,N_1647,N_1352);
nand U2823 (N_2823,N_1474,N_1677);
nor U2824 (N_2824,N_1000,N_1087);
nand U2825 (N_2825,N_1238,N_1329);
nor U2826 (N_2826,N_1494,N_1604);
nand U2827 (N_2827,N_1890,N_1828);
nor U2828 (N_2828,N_1464,N_1329);
nor U2829 (N_2829,N_1091,N_1344);
or U2830 (N_2830,N_1964,N_1672);
or U2831 (N_2831,N_1424,N_1296);
nor U2832 (N_2832,N_1124,N_1975);
and U2833 (N_2833,N_1232,N_1693);
or U2834 (N_2834,N_1709,N_1532);
xnor U2835 (N_2835,N_1085,N_1133);
nand U2836 (N_2836,N_1528,N_1296);
nand U2837 (N_2837,N_1149,N_1651);
nand U2838 (N_2838,N_1441,N_1461);
nand U2839 (N_2839,N_1310,N_1512);
or U2840 (N_2840,N_1206,N_1565);
and U2841 (N_2841,N_1566,N_1926);
xnor U2842 (N_2842,N_1843,N_1767);
nor U2843 (N_2843,N_1373,N_1021);
nand U2844 (N_2844,N_1540,N_1862);
nor U2845 (N_2845,N_1146,N_1364);
nand U2846 (N_2846,N_1122,N_1284);
nand U2847 (N_2847,N_1578,N_1935);
and U2848 (N_2848,N_1406,N_1002);
and U2849 (N_2849,N_1705,N_1370);
and U2850 (N_2850,N_1525,N_1986);
xnor U2851 (N_2851,N_1914,N_1100);
or U2852 (N_2852,N_1427,N_1143);
or U2853 (N_2853,N_1202,N_1985);
or U2854 (N_2854,N_1299,N_1271);
and U2855 (N_2855,N_1517,N_1729);
nor U2856 (N_2856,N_1692,N_1697);
nor U2857 (N_2857,N_1844,N_1489);
or U2858 (N_2858,N_1458,N_1608);
nor U2859 (N_2859,N_1166,N_1673);
or U2860 (N_2860,N_1345,N_1032);
or U2861 (N_2861,N_1439,N_1413);
nor U2862 (N_2862,N_1445,N_1818);
or U2863 (N_2863,N_1300,N_1279);
nand U2864 (N_2864,N_1890,N_1193);
xor U2865 (N_2865,N_1537,N_1201);
and U2866 (N_2866,N_1226,N_1306);
nor U2867 (N_2867,N_1056,N_1605);
nand U2868 (N_2868,N_1134,N_1119);
or U2869 (N_2869,N_1930,N_1906);
nand U2870 (N_2870,N_1380,N_1632);
nand U2871 (N_2871,N_1082,N_1910);
and U2872 (N_2872,N_1052,N_1833);
nand U2873 (N_2873,N_1107,N_1480);
nand U2874 (N_2874,N_1042,N_1854);
and U2875 (N_2875,N_1450,N_1863);
nor U2876 (N_2876,N_1890,N_1085);
or U2877 (N_2877,N_1577,N_1719);
or U2878 (N_2878,N_1920,N_1327);
or U2879 (N_2879,N_1014,N_1144);
and U2880 (N_2880,N_1826,N_1386);
nand U2881 (N_2881,N_1373,N_1154);
or U2882 (N_2882,N_1060,N_1126);
nor U2883 (N_2883,N_1363,N_1669);
or U2884 (N_2884,N_1729,N_1201);
nand U2885 (N_2885,N_1238,N_1009);
nor U2886 (N_2886,N_1897,N_1514);
nand U2887 (N_2887,N_1741,N_1302);
nand U2888 (N_2888,N_1998,N_1924);
or U2889 (N_2889,N_1870,N_1948);
and U2890 (N_2890,N_1607,N_1723);
nor U2891 (N_2891,N_1612,N_1685);
nand U2892 (N_2892,N_1694,N_1405);
xor U2893 (N_2893,N_1401,N_1261);
and U2894 (N_2894,N_1580,N_1958);
or U2895 (N_2895,N_1154,N_1609);
nor U2896 (N_2896,N_1280,N_1925);
and U2897 (N_2897,N_1889,N_1678);
xnor U2898 (N_2898,N_1866,N_1794);
nand U2899 (N_2899,N_1421,N_1887);
nor U2900 (N_2900,N_1754,N_1010);
nand U2901 (N_2901,N_1097,N_1996);
and U2902 (N_2902,N_1019,N_1148);
nor U2903 (N_2903,N_1982,N_1607);
and U2904 (N_2904,N_1135,N_1040);
or U2905 (N_2905,N_1595,N_1680);
nand U2906 (N_2906,N_1748,N_1964);
nand U2907 (N_2907,N_1025,N_1811);
or U2908 (N_2908,N_1044,N_1989);
or U2909 (N_2909,N_1829,N_1646);
nand U2910 (N_2910,N_1238,N_1514);
and U2911 (N_2911,N_1292,N_1244);
nand U2912 (N_2912,N_1724,N_1412);
nand U2913 (N_2913,N_1429,N_1303);
and U2914 (N_2914,N_1565,N_1614);
nor U2915 (N_2915,N_1101,N_1851);
or U2916 (N_2916,N_1068,N_1825);
nand U2917 (N_2917,N_1449,N_1318);
and U2918 (N_2918,N_1489,N_1093);
nor U2919 (N_2919,N_1306,N_1954);
nor U2920 (N_2920,N_1879,N_1186);
or U2921 (N_2921,N_1290,N_1340);
or U2922 (N_2922,N_1164,N_1977);
and U2923 (N_2923,N_1723,N_1157);
or U2924 (N_2924,N_1446,N_1907);
nand U2925 (N_2925,N_1097,N_1489);
nor U2926 (N_2926,N_1494,N_1927);
xnor U2927 (N_2927,N_1854,N_1904);
xnor U2928 (N_2928,N_1567,N_1817);
nor U2929 (N_2929,N_1517,N_1313);
or U2930 (N_2930,N_1379,N_1316);
nor U2931 (N_2931,N_1215,N_1767);
nor U2932 (N_2932,N_1252,N_1882);
nor U2933 (N_2933,N_1114,N_1447);
xnor U2934 (N_2934,N_1422,N_1962);
nand U2935 (N_2935,N_1953,N_1185);
or U2936 (N_2936,N_1248,N_1739);
or U2937 (N_2937,N_1936,N_1374);
xor U2938 (N_2938,N_1634,N_1893);
and U2939 (N_2939,N_1984,N_1912);
or U2940 (N_2940,N_1334,N_1086);
and U2941 (N_2941,N_1697,N_1706);
and U2942 (N_2942,N_1070,N_1422);
and U2943 (N_2943,N_1526,N_1456);
nand U2944 (N_2944,N_1365,N_1466);
or U2945 (N_2945,N_1696,N_1464);
nor U2946 (N_2946,N_1436,N_1537);
or U2947 (N_2947,N_1033,N_1167);
and U2948 (N_2948,N_1372,N_1342);
or U2949 (N_2949,N_1517,N_1374);
nor U2950 (N_2950,N_1758,N_1614);
and U2951 (N_2951,N_1348,N_1211);
xor U2952 (N_2952,N_1699,N_1933);
nand U2953 (N_2953,N_1409,N_1401);
nand U2954 (N_2954,N_1119,N_1474);
and U2955 (N_2955,N_1937,N_1556);
nand U2956 (N_2956,N_1822,N_1273);
nand U2957 (N_2957,N_1094,N_1702);
or U2958 (N_2958,N_1334,N_1540);
nand U2959 (N_2959,N_1010,N_1384);
nand U2960 (N_2960,N_1359,N_1740);
or U2961 (N_2961,N_1498,N_1263);
or U2962 (N_2962,N_1265,N_1040);
nor U2963 (N_2963,N_1582,N_1594);
or U2964 (N_2964,N_1231,N_1995);
nand U2965 (N_2965,N_1380,N_1964);
nand U2966 (N_2966,N_1363,N_1837);
nor U2967 (N_2967,N_1596,N_1879);
xnor U2968 (N_2968,N_1871,N_1425);
or U2969 (N_2969,N_1995,N_1276);
nor U2970 (N_2970,N_1065,N_1006);
and U2971 (N_2971,N_1984,N_1648);
and U2972 (N_2972,N_1754,N_1922);
nor U2973 (N_2973,N_1670,N_1714);
xor U2974 (N_2974,N_1276,N_1923);
nand U2975 (N_2975,N_1246,N_1437);
or U2976 (N_2976,N_1316,N_1344);
or U2977 (N_2977,N_1026,N_1796);
nor U2978 (N_2978,N_1983,N_1638);
nor U2979 (N_2979,N_1582,N_1687);
xnor U2980 (N_2980,N_1707,N_1416);
nand U2981 (N_2981,N_1726,N_1780);
nand U2982 (N_2982,N_1539,N_1355);
nand U2983 (N_2983,N_1389,N_1264);
nand U2984 (N_2984,N_1093,N_1292);
and U2985 (N_2985,N_1129,N_1591);
or U2986 (N_2986,N_1163,N_1106);
nand U2987 (N_2987,N_1967,N_1393);
or U2988 (N_2988,N_1201,N_1629);
nor U2989 (N_2989,N_1232,N_1583);
nor U2990 (N_2990,N_1754,N_1240);
or U2991 (N_2991,N_1121,N_1789);
nand U2992 (N_2992,N_1951,N_1681);
nand U2993 (N_2993,N_1931,N_1489);
xor U2994 (N_2994,N_1735,N_1032);
and U2995 (N_2995,N_1359,N_1143);
or U2996 (N_2996,N_1009,N_1335);
or U2997 (N_2997,N_1151,N_1267);
nand U2998 (N_2998,N_1154,N_1144);
xnor U2999 (N_2999,N_1769,N_1963);
or U3000 (N_3000,N_2699,N_2775);
and U3001 (N_3001,N_2535,N_2786);
and U3002 (N_3002,N_2173,N_2718);
nand U3003 (N_3003,N_2659,N_2904);
xnor U3004 (N_3004,N_2208,N_2636);
or U3005 (N_3005,N_2561,N_2292);
or U3006 (N_3006,N_2562,N_2960);
nand U3007 (N_3007,N_2122,N_2119);
xor U3008 (N_3008,N_2335,N_2681);
and U3009 (N_3009,N_2186,N_2135);
nor U3010 (N_3010,N_2440,N_2226);
nor U3011 (N_3011,N_2949,N_2253);
nand U3012 (N_3012,N_2781,N_2650);
and U3013 (N_3013,N_2228,N_2583);
and U3014 (N_3014,N_2995,N_2644);
nand U3015 (N_3015,N_2570,N_2779);
or U3016 (N_3016,N_2913,N_2615);
nor U3017 (N_3017,N_2777,N_2682);
and U3018 (N_3018,N_2558,N_2569);
or U3019 (N_3019,N_2693,N_2818);
or U3020 (N_3020,N_2072,N_2540);
nor U3021 (N_3021,N_2755,N_2743);
nor U3022 (N_3022,N_2311,N_2518);
nand U3023 (N_3023,N_2478,N_2134);
nand U3024 (N_3024,N_2336,N_2056);
nor U3025 (N_3025,N_2938,N_2204);
and U3026 (N_3026,N_2288,N_2829);
or U3027 (N_3027,N_2555,N_2748);
nand U3028 (N_3028,N_2005,N_2930);
nand U3029 (N_3029,N_2945,N_2325);
nor U3030 (N_3030,N_2018,N_2340);
or U3031 (N_3031,N_2724,N_2716);
nand U3032 (N_3032,N_2798,N_2805);
and U3033 (N_3033,N_2066,N_2399);
and U3034 (N_3034,N_2679,N_2532);
nand U3035 (N_3035,N_2729,N_2692);
nor U3036 (N_3036,N_2663,N_2216);
and U3037 (N_3037,N_2011,N_2948);
nor U3038 (N_3038,N_2334,N_2922);
nor U3039 (N_3039,N_2266,N_2107);
nand U3040 (N_3040,N_2898,N_2835);
xnor U3041 (N_3041,N_2402,N_2167);
nor U3042 (N_3042,N_2617,N_2668);
nand U3043 (N_3043,N_2812,N_2227);
nand U3044 (N_3044,N_2243,N_2593);
nor U3045 (N_3045,N_2653,N_2610);
nor U3046 (N_3046,N_2050,N_2374);
nor U3047 (N_3047,N_2944,N_2851);
or U3048 (N_3048,N_2580,N_2064);
and U3049 (N_3049,N_2279,N_2907);
or U3050 (N_3050,N_2577,N_2892);
xor U3051 (N_3051,N_2806,N_2890);
xor U3052 (N_3052,N_2275,N_2665);
and U3053 (N_3053,N_2745,N_2795);
xor U3054 (N_3054,N_2021,N_2799);
and U3055 (N_3055,N_2385,N_2906);
and U3056 (N_3056,N_2029,N_2308);
nand U3057 (N_3057,N_2258,N_2883);
nand U3058 (N_3058,N_2100,N_2567);
nand U3059 (N_3059,N_2623,N_2363);
nor U3060 (N_3060,N_2655,N_2811);
and U3061 (N_3061,N_2975,N_2486);
nand U3062 (N_3062,N_2954,N_2044);
and U3063 (N_3063,N_2982,N_2759);
or U3064 (N_3064,N_2863,N_2574);
and U3065 (N_3065,N_2470,N_2888);
or U3066 (N_3066,N_2451,N_2804);
nor U3067 (N_3067,N_2246,N_2347);
and U3068 (N_3068,N_2549,N_2928);
nor U3069 (N_3069,N_2589,N_2876);
nand U3070 (N_3070,N_2645,N_2868);
and U3071 (N_3071,N_2409,N_2283);
xnor U3072 (N_3072,N_2101,N_2970);
nor U3073 (N_3073,N_2460,N_2850);
nand U3074 (N_3074,N_2112,N_2475);
and U3075 (N_3075,N_2788,N_2980);
or U3076 (N_3076,N_2421,N_2953);
or U3077 (N_3077,N_2096,N_2927);
or U3078 (N_3078,N_2143,N_2074);
xnor U3079 (N_3079,N_2834,N_2712);
nor U3080 (N_3080,N_2462,N_2778);
nor U3081 (N_3081,N_2495,N_2853);
and U3082 (N_3082,N_2452,N_2115);
or U3083 (N_3083,N_2849,N_2053);
nand U3084 (N_3084,N_2218,N_2746);
nor U3085 (N_3085,N_2092,N_2594);
and U3086 (N_3086,N_2735,N_2527);
nand U3087 (N_3087,N_2229,N_2703);
nand U3088 (N_3088,N_2999,N_2661);
nor U3089 (N_3089,N_2903,N_2916);
and U3090 (N_3090,N_2200,N_2408);
or U3091 (N_3091,N_2051,N_2274);
or U3092 (N_3092,N_2550,N_2464);
nand U3093 (N_3093,N_2894,N_2313);
nor U3094 (N_3094,N_2941,N_2762);
and U3095 (N_3095,N_2760,N_2177);
or U3096 (N_3096,N_2541,N_2384);
nor U3097 (N_3097,N_2392,N_2284);
nor U3098 (N_3098,N_2675,N_2842);
and U3099 (N_3099,N_2994,N_2217);
and U3100 (N_3100,N_2711,N_2105);
or U3101 (N_3101,N_2537,N_2819);
nand U3102 (N_3102,N_2526,N_2635);
and U3103 (N_3103,N_2738,N_2067);
nor U3104 (N_3104,N_2536,N_2696);
or U3105 (N_3105,N_2480,N_2298);
nor U3106 (N_3106,N_2024,N_2989);
or U3107 (N_3107,N_2036,N_2744);
and U3108 (N_3108,N_2225,N_2439);
or U3109 (N_3109,N_2168,N_2559);
or U3110 (N_3110,N_2694,N_2691);
nand U3111 (N_3111,N_2039,N_2078);
nor U3112 (N_3112,N_2161,N_2048);
and U3113 (N_3113,N_2068,N_2774);
nor U3114 (N_3114,N_2882,N_2169);
nand U3115 (N_3115,N_2430,N_2707);
and U3116 (N_3116,N_2341,N_2730);
nand U3117 (N_3117,N_2267,N_2909);
or U3118 (N_3118,N_2701,N_2764);
or U3119 (N_3119,N_2790,N_2905);
or U3120 (N_3120,N_2817,N_2479);
xnor U3121 (N_3121,N_2962,N_2736);
and U3122 (N_3122,N_2242,N_2089);
nor U3123 (N_3123,N_2222,N_2377);
nor U3124 (N_3124,N_2155,N_2111);
nor U3125 (N_3125,N_2420,N_2614);
and U3126 (N_3126,N_2387,N_2528);
nor U3127 (N_3127,N_2698,N_2504);
nor U3128 (N_3128,N_2171,N_2702);
xor U3129 (N_3129,N_2722,N_2734);
or U3130 (N_3130,N_2320,N_2502);
nor U3131 (N_3131,N_2471,N_2500);
or U3132 (N_3132,N_2912,N_2525);
or U3133 (N_3133,N_2448,N_2827);
nand U3134 (N_3134,N_2632,N_2847);
or U3135 (N_3135,N_2484,N_2885);
nor U3136 (N_3136,N_2856,N_2503);
and U3137 (N_3137,N_2104,N_2162);
nor U3138 (N_3138,N_2578,N_2040);
nand U3139 (N_3139,N_2412,N_2654);
or U3140 (N_3140,N_2880,N_2358);
nor U3141 (N_3141,N_2785,N_2723);
nor U3142 (N_3142,N_2010,N_2917);
nand U3143 (N_3143,N_2671,N_2741);
nand U3144 (N_3144,N_2873,N_2772);
nand U3145 (N_3145,N_2328,N_2896);
nand U3146 (N_3146,N_2605,N_2052);
xnor U3147 (N_3147,N_2359,N_2126);
nand U3148 (N_3148,N_2080,N_2860);
nand U3149 (N_3149,N_2418,N_2684);
nor U3150 (N_3150,N_2386,N_2014);
nor U3151 (N_3151,N_2611,N_2366);
nand U3152 (N_3152,N_2520,N_2269);
nand U3153 (N_3153,N_2224,N_2543);
and U3154 (N_3154,N_2351,N_2545);
nor U3155 (N_3155,N_2680,N_2996);
and U3156 (N_3156,N_2485,N_2022);
or U3157 (N_3157,N_2803,N_2895);
or U3158 (N_3158,N_2183,N_2172);
and U3159 (N_3159,N_2784,N_2330);
nand U3160 (N_3160,N_2268,N_2733);
nand U3161 (N_3161,N_2375,N_2936);
and U3162 (N_3162,N_2008,N_2765);
and U3163 (N_3163,N_2534,N_2662);
nor U3164 (N_3164,N_2416,N_2091);
nor U3165 (N_3165,N_2401,N_2031);
or U3166 (N_3166,N_2247,N_2531);
and U3167 (N_3167,N_2466,N_2754);
and U3168 (N_3168,N_2825,N_2688);
and U3169 (N_3169,N_2165,N_2767);
nor U3170 (N_3170,N_2166,N_2704);
and U3171 (N_3171,N_2087,N_2394);
nor U3172 (N_3172,N_2461,N_2564);
nor U3173 (N_3173,N_2926,N_2028);
and U3174 (N_3174,N_2816,N_2968);
nor U3175 (N_3175,N_2556,N_2921);
or U3176 (N_3176,N_2188,N_2182);
or U3177 (N_3177,N_2342,N_2059);
and U3178 (N_3178,N_2147,N_2150);
nand U3179 (N_3179,N_2411,N_2251);
or U3180 (N_3180,N_2465,N_2281);
nand U3181 (N_3181,N_2372,N_2317);
or U3182 (N_3182,N_2690,N_2318);
and U3183 (N_3183,N_2206,N_2006);
xnor U3184 (N_3184,N_2770,N_2581);
nor U3185 (N_3185,N_2306,N_2884);
or U3186 (N_3186,N_2163,N_2986);
xnor U3187 (N_3187,N_2131,N_2295);
xor U3188 (N_3188,N_2255,N_2355);
nor U3189 (N_3189,N_2133,N_2343);
or U3190 (N_3190,N_2138,N_2406);
nand U3191 (N_3191,N_2004,N_2219);
and U3192 (N_3192,N_2482,N_2547);
nand U3193 (N_3193,N_2307,N_2220);
nor U3194 (N_3194,N_2136,N_2413);
nand U3195 (N_3195,N_2338,N_2129);
and U3196 (N_3196,N_2705,N_2151);
nand U3197 (N_3197,N_2291,N_2606);
or U3198 (N_3198,N_2717,N_2700);
nand U3199 (N_3199,N_2758,N_2727);
nor U3200 (N_3200,N_2086,N_2791);
or U3201 (N_3201,N_2290,N_2557);
and U3202 (N_3202,N_2519,N_2839);
xnor U3203 (N_3203,N_2591,N_2587);
nand U3204 (N_3204,N_2472,N_2942);
or U3205 (N_3205,N_2807,N_2207);
nand U3206 (N_3206,N_2373,N_2918);
or U3207 (N_3207,N_2613,N_2981);
nor U3208 (N_3208,N_2796,N_2622);
and U3209 (N_3209,N_2859,N_2310);
nand U3210 (N_3210,N_2003,N_2449);
nor U3211 (N_3211,N_2602,N_2007);
nand U3212 (N_3212,N_2128,N_2214);
nor U3213 (N_3213,N_2881,N_2141);
and U3214 (N_3214,N_2045,N_2720);
and U3215 (N_3215,N_2508,N_2658);
and U3216 (N_3216,N_2278,N_2794);
and U3217 (N_3217,N_2752,N_2194);
or U3218 (N_3218,N_2174,N_2958);
or U3219 (N_3219,N_2315,N_2879);
nand U3220 (N_3220,N_2319,N_2552);
nor U3221 (N_3221,N_2271,N_2350);
or U3222 (N_3222,N_2084,N_2023);
nor U3223 (N_3223,N_2585,N_2117);
or U3224 (N_3224,N_2763,N_2749);
and U3225 (N_3225,N_2706,N_2400);
nand U3226 (N_3226,N_2998,N_2405);
nor U3227 (N_3227,N_2491,N_2193);
or U3228 (N_3228,N_2522,N_2599);
nor U3229 (N_3229,N_2142,N_2871);
nand U3230 (N_3230,N_2248,N_2333);
nand U3231 (N_3231,N_2265,N_2721);
and U3232 (N_3232,N_2769,N_2677);
nand U3233 (N_3233,N_2867,N_2624);
nand U3234 (N_3234,N_2047,N_2497);
and U3235 (N_3235,N_2455,N_2957);
or U3236 (N_3236,N_2349,N_2598);
xor U3237 (N_3237,N_2361,N_2002);
and U3238 (N_3238,N_2302,N_2713);
nor U3239 (N_3239,N_2590,N_2858);
xor U3240 (N_3240,N_2961,N_2951);
or U3241 (N_3241,N_2813,N_2352);
xnor U3242 (N_3242,N_2647,N_2846);
nand U3243 (N_3243,N_2893,N_2862);
or U3244 (N_3244,N_2309,N_2972);
and U3245 (N_3245,N_2203,N_2038);
nand U3246 (N_3246,N_2637,N_2297);
and U3247 (N_3247,N_2094,N_2609);
xor U3248 (N_3248,N_2260,N_2649);
or U3249 (N_3249,N_2304,N_2652);
nand U3250 (N_3250,N_2512,N_2544);
nor U3251 (N_3251,N_2822,N_2757);
nor U3252 (N_3252,N_2792,N_2563);
and U3253 (N_3253,N_2689,N_2009);
nor U3254 (N_3254,N_2037,N_2766);
and U3255 (N_3255,N_2090,N_2877);
nand U3256 (N_3256,N_2686,N_2546);
or U3257 (N_3257,N_2501,N_2487);
or U3258 (N_3258,N_2529,N_2164);
or U3259 (N_3259,N_2221,N_2034);
xnor U3260 (N_3260,N_2510,N_2118);
xnor U3261 (N_3261,N_2145,N_2296);
or U3262 (N_3262,N_2789,N_2576);
nand U3263 (N_3263,N_2293,N_2323);
or U3264 (N_3264,N_2345,N_2468);
or U3265 (N_3265,N_2483,N_2554);
or U3266 (N_3266,N_2241,N_2404);
and U3267 (N_3267,N_2857,N_2616);
nor U3268 (N_3268,N_2820,N_2499);
nor U3269 (N_3269,N_2509,N_2427);
nand U3270 (N_3270,N_2742,N_2120);
or U3271 (N_3271,N_2782,N_2425);
or U3272 (N_3272,N_2726,N_2176);
nand U3273 (N_3273,N_2852,N_2124);
xnor U3274 (N_3274,N_2673,N_2641);
nand U3275 (N_3275,N_2414,N_2236);
or U3276 (N_3276,N_2436,N_2709);
nand U3277 (N_3277,N_2127,N_2337);
and U3278 (N_3278,N_2097,N_2808);
or U3279 (N_3279,N_2521,N_2433);
xnor U3280 (N_3280,N_2821,N_2506);
xor U3281 (N_3281,N_2270,N_2728);
or U3282 (N_3282,N_2417,N_2210);
nand U3283 (N_3283,N_2215,N_2073);
and U3284 (N_3284,N_2113,N_2075);
nand U3285 (N_3285,N_2316,N_2354);
or U3286 (N_3286,N_2300,N_2910);
nor U3287 (N_3287,N_2952,N_2185);
nand U3288 (N_3288,N_2571,N_2191);
or U3289 (N_3289,N_2493,N_2380);
xnor U3290 (N_3290,N_2457,N_2940);
nor U3291 (N_3291,N_2667,N_2376);
xor U3292 (N_3292,N_2687,N_2159);
nor U3293 (N_3293,N_2058,N_2250);
and U3294 (N_3294,N_2190,N_2391);
and U3295 (N_3295,N_2395,N_2971);
nor U3296 (N_3296,N_2175,N_2178);
nand U3297 (N_3297,N_2923,N_2114);
and U3298 (N_3298,N_2230,N_2937);
and U3299 (N_3299,N_2146,N_2294);
and U3300 (N_3300,N_2530,N_2979);
and U3301 (N_3301,N_2619,N_2144);
and U3302 (N_3302,N_2331,N_2054);
xnor U3303 (N_3303,N_2625,N_2865);
or U3304 (N_3304,N_2393,N_2993);
nor U3305 (N_3305,N_2572,N_2978);
nand U3306 (N_3306,N_2033,N_2783);
xor U3307 (N_3307,N_2065,N_2327);
nor U3308 (N_3308,N_2832,N_2121);
nand U3309 (N_3309,N_2666,N_2715);
nand U3310 (N_3310,N_2170,N_2628);
nor U3311 (N_3311,N_2367,N_2833);
and U3312 (N_3312,N_2303,N_2160);
nor U3313 (N_3313,N_2780,N_2761);
and U3314 (N_3314,N_2601,N_2843);
and U3315 (N_3315,N_2339,N_2634);
nand U3316 (N_3316,N_2431,N_2276);
or U3317 (N_3317,N_2116,N_2234);
and U3318 (N_3318,N_2638,N_2596);
and U3319 (N_3319,N_2826,N_2648);
and U3320 (N_3320,N_2071,N_2751);
or U3321 (N_3321,N_2670,N_2459);
nor U3322 (N_3322,N_2125,N_2245);
nor U3323 (N_3323,N_2983,N_2244);
nor U3324 (N_3324,N_2438,N_2737);
and U3325 (N_3325,N_2069,N_2911);
and U3326 (N_3326,N_2035,N_2403);
xor U3327 (N_3327,N_2025,N_2473);
nor U3328 (N_3328,N_2429,N_2202);
nor U3329 (N_3329,N_2233,N_2565);
nor U3330 (N_3330,N_2586,N_2450);
or U3331 (N_3331,N_2061,N_2914);
nor U3332 (N_3332,N_2600,N_2189);
and U3333 (N_3333,N_2643,N_2836);
and U3334 (N_3334,N_2149,N_2332);
nand U3335 (N_3335,N_2368,N_2088);
nand U3336 (N_3336,N_2965,N_2844);
or U3337 (N_3337,N_2725,N_2442);
and U3338 (N_3338,N_2130,N_2657);
nor U3339 (N_3339,N_2838,N_2287);
or U3340 (N_3340,N_2205,N_2719);
nor U3341 (N_3341,N_2209,N_2046);
and U3342 (N_3342,N_2612,N_2568);
nor U3343 (N_3343,N_2597,N_2444);
and U3344 (N_3344,N_2592,N_2840);
or U3345 (N_3345,N_2201,N_2132);
nand U3346 (N_3346,N_2815,N_2371);
nand U3347 (N_3347,N_2063,N_2969);
and U3348 (N_3348,N_2845,N_2062);
or U3349 (N_3349,N_2157,N_2055);
nor U3350 (N_3350,N_2286,N_2192);
nand U3351 (N_3351,N_2032,N_2640);
or U3352 (N_3352,N_2180,N_2516);
or U3353 (N_3353,N_2831,N_2950);
or U3354 (N_3354,N_2110,N_2517);
nor U3355 (N_3355,N_2642,N_2030);
and U3356 (N_3356,N_2947,N_2855);
nand U3357 (N_3357,N_2966,N_2515);
xnor U3358 (N_3358,N_2618,N_2321);
xnor U3359 (N_3359,N_2507,N_2864);
nor U3360 (N_3360,N_2935,N_2049);
nor U3361 (N_3361,N_2261,N_2042);
and U3362 (N_3362,N_2977,N_2365);
nand U3363 (N_3363,N_2148,N_2277);
and U3364 (N_3364,N_2070,N_2181);
nor U3365 (N_3365,N_2664,N_2305);
nor U3366 (N_3366,N_2739,N_2262);
and U3367 (N_3367,N_2077,N_2474);
nand U3368 (N_3368,N_2870,N_2357);
and U3369 (N_3369,N_2802,N_2020);
or U3370 (N_3370,N_2874,N_2828);
xnor U3371 (N_3371,N_2076,N_2232);
nor U3372 (N_3372,N_2560,N_2902);
xnor U3373 (N_3373,N_2198,N_2083);
or U3374 (N_3374,N_2924,N_2223);
and U3375 (N_3375,N_2383,N_2633);
nand U3376 (N_3376,N_2955,N_2824);
nor U3377 (N_3377,N_2488,N_2991);
nand U3378 (N_3378,N_2946,N_2579);
nor U3379 (N_3379,N_2370,N_2551);
and U3380 (N_3380,N_2184,N_2106);
xnor U3381 (N_3381,N_2095,N_2872);
or U3382 (N_3382,N_2875,N_2239);
nor U3383 (N_3383,N_2933,N_2747);
nand U3384 (N_3384,N_2787,N_2697);
xnor U3385 (N_3385,N_2103,N_2428);
or U3386 (N_3386,N_2973,N_2801);
and U3387 (N_3387,N_2674,N_2900);
or U3388 (N_3388,N_2607,N_2109);
nand U3389 (N_3389,N_2324,N_2932);
nand U3390 (N_3390,N_2257,N_2447);
or U3391 (N_3391,N_2099,N_2443);
and U3392 (N_3392,N_2629,N_2492);
or U3393 (N_3393,N_2841,N_2771);
nand U3394 (N_3394,N_2630,N_2489);
nor U3395 (N_3395,N_2511,N_2369);
nor U3396 (N_3396,N_2273,N_2001);
and U3397 (N_3397,N_2997,N_2093);
nand U3398 (N_3398,N_2814,N_2445);
or U3399 (N_3399,N_2397,N_2732);
nand U3400 (N_3400,N_2626,N_2553);
and U3401 (N_3401,N_2582,N_2390);
or U3402 (N_3402,N_2013,N_2263);
nor U3403 (N_3403,N_2211,N_2364);
or U3404 (N_3404,N_2041,N_2710);
nand U3405 (N_3405,N_2139,N_2424);
nand U3406 (N_3406,N_2939,N_2481);
nor U3407 (N_3407,N_2823,N_2861);
nor U3408 (N_3408,N_2398,N_2179);
and U3409 (N_3409,N_2886,N_2153);
xnor U3410 (N_3410,N_2490,N_2187);
nor U3411 (N_3411,N_2282,N_2627);
or U3412 (N_3412,N_2280,N_2381);
or U3413 (N_3413,N_2695,N_2897);
nor U3414 (N_3414,N_2249,N_2158);
and U3415 (N_3415,N_2651,N_2848);
xor U3416 (N_3416,N_2683,N_2456);
or U3417 (N_3417,N_2523,N_2919);
xor U3418 (N_3418,N_2672,N_2542);
nor U3419 (N_3419,N_2348,N_2967);
and U3420 (N_3420,N_2731,N_2102);
nor U3421 (N_3421,N_2566,N_2256);
nor U3422 (N_3422,N_2943,N_2889);
nor U3423 (N_3423,N_2584,N_2869);
nor U3424 (N_3424,N_2753,N_2756);
nand U3425 (N_3425,N_2082,N_2017);
or U3426 (N_3426,N_2389,N_2797);
and U3427 (N_3427,N_2469,N_2974);
nor U3428 (N_3428,N_2353,N_2254);
or U3429 (N_3429,N_2043,N_2238);
nor U3430 (N_3430,N_2329,N_2415);
and U3431 (N_3431,N_2396,N_2407);
or U3432 (N_3432,N_2299,N_2621);
xnor U3433 (N_3433,N_2012,N_2085);
or U3434 (N_3434,N_2646,N_2656);
nand U3435 (N_3435,N_2432,N_2379);
xor U3436 (N_3436,N_2956,N_2477);
nor U3437 (N_3437,N_2603,N_2426);
or U3438 (N_3438,N_2987,N_2604);
nand U3439 (N_3439,N_2410,N_2830);
or U3440 (N_3440,N_2212,N_2513);
or U3441 (N_3441,N_2467,N_2196);
nor U3442 (N_3442,N_2199,N_2963);
nor U3443 (N_3443,N_2344,N_2362);
nor U3444 (N_3444,N_2108,N_2639);
and U3445 (N_3445,N_2524,N_2312);
and U3446 (N_3446,N_2213,N_2929);
nand U3447 (N_3447,N_2959,N_2915);
or U3448 (N_3448,N_2908,N_2750);
nor U3449 (N_3449,N_2608,N_2575);
nand U3450 (N_3450,N_2714,N_2514);
or U3451 (N_3451,N_2140,N_2195);
or U3452 (N_3452,N_2538,N_2422);
nor U3453 (N_3453,N_2154,N_2988);
nand U3454 (N_3454,N_2272,N_2285);
nand U3455 (N_3455,N_2322,N_2434);
nand U3456 (N_3456,N_2240,N_2708);
nand U3457 (N_3457,N_2346,N_2388);
xor U3458 (N_3458,N_2152,N_2081);
or U3459 (N_3459,N_2768,N_2252);
or U3460 (N_3460,N_2992,N_2231);
xor U3461 (N_3461,N_2837,N_2573);
nor U3462 (N_3462,N_2934,N_2595);
nand U3463 (N_3463,N_2548,N_2123);
xnor U3464 (N_3464,N_2446,N_2463);
or U3465 (N_3465,N_2984,N_2027);
nor U3466 (N_3466,N_2259,N_2454);
nand U3467 (N_3467,N_2423,N_2925);
nand U3468 (N_3468,N_2494,N_2015);
and U3469 (N_3469,N_2437,N_2678);
nand U3470 (N_3470,N_2079,N_2026);
nand U3471 (N_3471,N_2676,N_2990);
nor U3472 (N_3472,N_2453,N_2878);
xnor U3473 (N_3473,N_2669,N_2631);
and U3474 (N_3474,N_2901,N_2920);
and U3475 (N_3475,N_2057,N_2505);
nand U3476 (N_3476,N_2419,N_2356);
or U3477 (N_3477,N_2098,N_2314);
and U3478 (N_3478,N_2793,N_2458);
nor U3479 (N_3479,N_2533,N_2060);
or U3480 (N_3480,N_2476,N_2264);
nor U3481 (N_3481,N_2887,N_2985);
nand U3482 (N_3482,N_2289,N_2237);
and U3483 (N_3483,N_2382,N_2931);
xnor U3484 (N_3484,N_2891,N_2660);
nor U3485 (N_3485,N_2866,N_2539);
nand U3486 (N_3486,N_2588,N_2378);
nand U3487 (N_3487,N_2019,N_2441);
nand U3488 (N_3488,N_2326,N_2235);
and U3489 (N_3489,N_2435,N_2301);
nand U3490 (N_3490,N_2156,N_2620);
nor U3491 (N_3491,N_2854,N_2496);
nor U3492 (N_3492,N_2000,N_2498);
nor U3493 (N_3493,N_2809,N_2360);
nand U3494 (N_3494,N_2740,N_2137);
and U3495 (N_3495,N_2685,N_2810);
or U3496 (N_3496,N_2016,N_2776);
nand U3497 (N_3497,N_2976,N_2197);
or U3498 (N_3498,N_2800,N_2773);
nand U3499 (N_3499,N_2899,N_2964);
xnor U3500 (N_3500,N_2898,N_2427);
or U3501 (N_3501,N_2750,N_2419);
or U3502 (N_3502,N_2879,N_2244);
nand U3503 (N_3503,N_2119,N_2726);
and U3504 (N_3504,N_2744,N_2449);
or U3505 (N_3505,N_2018,N_2698);
or U3506 (N_3506,N_2857,N_2357);
and U3507 (N_3507,N_2858,N_2159);
or U3508 (N_3508,N_2134,N_2887);
and U3509 (N_3509,N_2868,N_2786);
or U3510 (N_3510,N_2539,N_2963);
xnor U3511 (N_3511,N_2691,N_2458);
and U3512 (N_3512,N_2862,N_2315);
and U3513 (N_3513,N_2351,N_2277);
nor U3514 (N_3514,N_2175,N_2825);
nand U3515 (N_3515,N_2925,N_2985);
nand U3516 (N_3516,N_2479,N_2409);
or U3517 (N_3517,N_2055,N_2684);
nor U3518 (N_3518,N_2285,N_2960);
or U3519 (N_3519,N_2595,N_2809);
and U3520 (N_3520,N_2881,N_2826);
or U3521 (N_3521,N_2797,N_2969);
and U3522 (N_3522,N_2981,N_2972);
nor U3523 (N_3523,N_2091,N_2801);
and U3524 (N_3524,N_2260,N_2822);
nor U3525 (N_3525,N_2881,N_2989);
nor U3526 (N_3526,N_2123,N_2648);
nand U3527 (N_3527,N_2323,N_2639);
and U3528 (N_3528,N_2883,N_2720);
nor U3529 (N_3529,N_2655,N_2226);
nor U3530 (N_3530,N_2421,N_2246);
and U3531 (N_3531,N_2782,N_2762);
or U3532 (N_3532,N_2486,N_2113);
nor U3533 (N_3533,N_2631,N_2390);
nand U3534 (N_3534,N_2738,N_2437);
nor U3535 (N_3535,N_2965,N_2611);
xor U3536 (N_3536,N_2283,N_2870);
nand U3537 (N_3537,N_2316,N_2489);
or U3538 (N_3538,N_2704,N_2109);
nor U3539 (N_3539,N_2871,N_2980);
and U3540 (N_3540,N_2141,N_2370);
or U3541 (N_3541,N_2091,N_2902);
nor U3542 (N_3542,N_2696,N_2036);
or U3543 (N_3543,N_2164,N_2595);
nand U3544 (N_3544,N_2200,N_2184);
nand U3545 (N_3545,N_2964,N_2735);
or U3546 (N_3546,N_2038,N_2792);
or U3547 (N_3547,N_2908,N_2266);
nand U3548 (N_3548,N_2271,N_2107);
nor U3549 (N_3549,N_2331,N_2283);
or U3550 (N_3550,N_2059,N_2154);
nand U3551 (N_3551,N_2386,N_2715);
nor U3552 (N_3552,N_2193,N_2220);
and U3553 (N_3553,N_2754,N_2052);
xnor U3554 (N_3554,N_2340,N_2906);
xnor U3555 (N_3555,N_2564,N_2578);
xnor U3556 (N_3556,N_2063,N_2299);
and U3557 (N_3557,N_2691,N_2248);
nand U3558 (N_3558,N_2264,N_2940);
and U3559 (N_3559,N_2734,N_2981);
or U3560 (N_3560,N_2004,N_2134);
nor U3561 (N_3561,N_2799,N_2972);
nor U3562 (N_3562,N_2691,N_2632);
nand U3563 (N_3563,N_2981,N_2286);
nand U3564 (N_3564,N_2857,N_2813);
xor U3565 (N_3565,N_2022,N_2470);
nand U3566 (N_3566,N_2758,N_2085);
nand U3567 (N_3567,N_2088,N_2736);
and U3568 (N_3568,N_2409,N_2793);
nor U3569 (N_3569,N_2446,N_2029);
or U3570 (N_3570,N_2241,N_2787);
nor U3571 (N_3571,N_2861,N_2599);
nand U3572 (N_3572,N_2930,N_2660);
or U3573 (N_3573,N_2625,N_2790);
or U3574 (N_3574,N_2817,N_2190);
nand U3575 (N_3575,N_2411,N_2198);
and U3576 (N_3576,N_2796,N_2204);
and U3577 (N_3577,N_2538,N_2237);
and U3578 (N_3578,N_2147,N_2542);
and U3579 (N_3579,N_2796,N_2991);
or U3580 (N_3580,N_2305,N_2484);
or U3581 (N_3581,N_2920,N_2436);
and U3582 (N_3582,N_2980,N_2719);
or U3583 (N_3583,N_2499,N_2364);
and U3584 (N_3584,N_2627,N_2820);
nand U3585 (N_3585,N_2942,N_2702);
or U3586 (N_3586,N_2187,N_2146);
nor U3587 (N_3587,N_2310,N_2609);
nand U3588 (N_3588,N_2346,N_2387);
xnor U3589 (N_3589,N_2079,N_2149);
nand U3590 (N_3590,N_2093,N_2818);
and U3591 (N_3591,N_2031,N_2554);
nor U3592 (N_3592,N_2332,N_2421);
and U3593 (N_3593,N_2112,N_2530);
nand U3594 (N_3594,N_2948,N_2585);
and U3595 (N_3595,N_2741,N_2579);
nand U3596 (N_3596,N_2137,N_2739);
or U3597 (N_3597,N_2006,N_2865);
or U3598 (N_3598,N_2331,N_2445);
and U3599 (N_3599,N_2487,N_2400);
nor U3600 (N_3600,N_2207,N_2435);
or U3601 (N_3601,N_2046,N_2216);
nor U3602 (N_3602,N_2447,N_2086);
nor U3603 (N_3603,N_2248,N_2499);
nor U3604 (N_3604,N_2695,N_2983);
nor U3605 (N_3605,N_2206,N_2007);
nand U3606 (N_3606,N_2034,N_2814);
and U3607 (N_3607,N_2787,N_2005);
nand U3608 (N_3608,N_2949,N_2515);
or U3609 (N_3609,N_2088,N_2688);
nand U3610 (N_3610,N_2606,N_2444);
or U3611 (N_3611,N_2661,N_2470);
and U3612 (N_3612,N_2148,N_2484);
or U3613 (N_3613,N_2707,N_2426);
and U3614 (N_3614,N_2476,N_2332);
nor U3615 (N_3615,N_2987,N_2935);
nor U3616 (N_3616,N_2155,N_2714);
nand U3617 (N_3617,N_2430,N_2844);
xor U3618 (N_3618,N_2681,N_2118);
nand U3619 (N_3619,N_2227,N_2195);
and U3620 (N_3620,N_2768,N_2478);
and U3621 (N_3621,N_2222,N_2291);
nor U3622 (N_3622,N_2167,N_2828);
nand U3623 (N_3623,N_2055,N_2957);
nand U3624 (N_3624,N_2939,N_2135);
and U3625 (N_3625,N_2806,N_2774);
nand U3626 (N_3626,N_2014,N_2259);
nand U3627 (N_3627,N_2988,N_2315);
or U3628 (N_3628,N_2584,N_2264);
nor U3629 (N_3629,N_2424,N_2600);
and U3630 (N_3630,N_2081,N_2669);
or U3631 (N_3631,N_2336,N_2685);
or U3632 (N_3632,N_2868,N_2322);
and U3633 (N_3633,N_2535,N_2927);
nor U3634 (N_3634,N_2229,N_2999);
nand U3635 (N_3635,N_2698,N_2845);
xnor U3636 (N_3636,N_2886,N_2257);
and U3637 (N_3637,N_2075,N_2873);
nand U3638 (N_3638,N_2856,N_2037);
and U3639 (N_3639,N_2100,N_2023);
and U3640 (N_3640,N_2346,N_2207);
nand U3641 (N_3641,N_2286,N_2432);
xor U3642 (N_3642,N_2989,N_2859);
or U3643 (N_3643,N_2798,N_2933);
or U3644 (N_3644,N_2696,N_2961);
nand U3645 (N_3645,N_2394,N_2456);
and U3646 (N_3646,N_2026,N_2484);
nand U3647 (N_3647,N_2027,N_2117);
or U3648 (N_3648,N_2131,N_2583);
nand U3649 (N_3649,N_2585,N_2078);
nand U3650 (N_3650,N_2962,N_2080);
nor U3651 (N_3651,N_2267,N_2759);
nor U3652 (N_3652,N_2090,N_2797);
or U3653 (N_3653,N_2583,N_2602);
or U3654 (N_3654,N_2263,N_2055);
nand U3655 (N_3655,N_2526,N_2427);
nor U3656 (N_3656,N_2755,N_2581);
nand U3657 (N_3657,N_2242,N_2932);
xnor U3658 (N_3658,N_2700,N_2623);
or U3659 (N_3659,N_2513,N_2321);
and U3660 (N_3660,N_2606,N_2973);
or U3661 (N_3661,N_2392,N_2717);
and U3662 (N_3662,N_2687,N_2866);
nand U3663 (N_3663,N_2565,N_2658);
nand U3664 (N_3664,N_2372,N_2349);
nand U3665 (N_3665,N_2491,N_2279);
or U3666 (N_3666,N_2851,N_2471);
nand U3667 (N_3667,N_2624,N_2734);
nor U3668 (N_3668,N_2693,N_2690);
nand U3669 (N_3669,N_2243,N_2887);
and U3670 (N_3670,N_2300,N_2812);
nor U3671 (N_3671,N_2155,N_2297);
nor U3672 (N_3672,N_2341,N_2651);
nor U3673 (N_3673,N_2003,N_2994);
or U3674 (N_3674,N_2407,N_2861);
nor U3675 (N_3675,N_2704,N_2545);
nand U3676 (N_3676,N_2586,N_2345);
and U3677 (N_3677,N_2512,N_2239);
nand U3678 (N_3678,N_2574,N_2805);
nor U3679 (N_3679,N_2013,N_2240);
or U3680 (N_3680,N_2555,N_2669);
nor U3681 (N_3681,N_2730,N_2260);
and U3682 (N_3682,N_2762,N_2812);
nand U3683 (N_3683,N_2452,N_2247);
and U3684 (N_3684,N_2055,N_2134);
nor U3685 (N_3685,N_2582,N_2974);
nand U3686 (N_3686,N_2331,N_2371);
and U3687 (N_3687,N_2132,N_2278);
nor U3688 (N_3688,N_2477,N_2877);
or U3689 (N_3689,N_2971,N_2340);
nand U3690 (N_3690,N_2597,N_2999);
or U3691 (N_3691,N_2283,N_2748);
nor U3692 (N_3692,N_2227,N_2194);
or U3693 (N_3693,N_2785,N_2749);
or U3694 (N_3694,N_2861,N_2435);
xor U3695 (N_3695,N_2265,N_2180);
and U3696 (N_3696,N_2182,N_2862);
nand U3697 (N_3697,N_2014,N_2625);
nand U3698 (N_3698,N_2635,N_2397);
or U3699 (N_3699,N_2554,N_2243);
nor U3700 (N_3700,N_2362,N_2607);
nor U3701 (N_3701,N_2133,N_2426);
nand U3702 (N_3702,N_2362,N_2611);
nor U3703 (N_3703,N_2176,N_2173);
and U3704 (N_3704,N_2893,N_2096);
and U3705 (N_3705,N_2411,N_2914);
and U3706 (N_3706,N_2936,N_2575);
or U3707 (N_3707,N_2366,N_2429);
and U3708 (N_3708,N_2904,N_2486);
and U3709 (N_3709,N_2582,N_2465);
and U3710 (N_3710,N_2448,N_2177);
xor U3711 (N_3711,N_2994,N_2947);
nand U3712 (N_3712,N_2909,N_2496);
or U3713 (N_3713,N_2418,N_2302);
nor U3714 (N_3714,N_2450,N_2542);
xnor U3715 (N_3715,N_2568,N_2031);
nor U3716 (N_3716,N_2336,N_2559);
or U3717 (N_3717,N_2920,N_2986);
or U3718 (N_3718,N_2335,N_2831);
nand U3719 (N_3719,N_2817,N_2423);
and U3720 (N_3720,N_2854,N_2522);
nand U3721 (N_3721,N_2194,N_2158);
and U3722 (N_3722,N_2843,N_2651);
nor U3723 (N_3723,N_2559,N_2843);
or U3724 (N_3724,N_2668,N_2332);
nor U3725 (N_3725,N_2544,N_2207);
nor U3726 (N_3726,N_2367,N_2222);
and U3727 (N_3727,N_2978,N_2491);
or U3728 (N_3728,N_2040,N_2151);
nor U3729 (N_3729,N_2597,N_2781);
nor U3730 (N_3730,N_2168,N_2758);
or U3731 (N_3731,N_2105,N_2795);
or U3732 (N_3732,N_2033,N_2511);
nor U3733 (N_3733,N_2188,N_2050);
nand U3734 (N_3734,N_2790,N_2729);
and U3735 (N_3735,N_2804,N_2117);
nand U3736 (N_3736,N_2305,N_2108);
or U3737 (N_3737,N_2018,N_2031);
nand U3738 (N_3738,N_2680,N_2493);
nand U3739 (N_3739,N_2929,N_2626);
and U3740 (N_3740,N_2285,N_2093);
nor U3741 (N_3741,N_2908,N_2070);
and U3742 (N_3742,N_2372,N_2890);
nor U3743 (N_3743,N_2234,N_2198);
or U3744 (N_3744,N_2200,N_2806);
nand U3745 (N_3745,N_2648,N_2928);
and U3746 (N_3746,N_2544,N_2078);
nand U3747 (N_3747,N_2053,N_2530);
nor U3748 (N_3748,N_2577,N_2120);
or U3749 (N_3749,N_2864,N_2186);
or U3750 (N_3750,N_2177,N_2717);
nand U3751 (N_3751,N_2900,N_2201);
or U3752 (N_3752,N_2886,N_2814);
nand U3753 (N_3753,N_2930,N_2109);
xnor U3754 (N_3754,N_2319,N_2731);
xnor U3755 (N_3755,N_2535,N_2430);
nor U3756 (N_3756,N_2957,N_2575);
or U3757 (N_3757,N_2898,N_2826);
nand U3758 (N_3758,N_2204,N_2334);
and U3759 (N_3759,N_2255,N_2417);
and U3760 (N_3760,N_2540,N_2933);
and U3761 (N_3761,N_2547,N_2642);
nor U3762 (N_3762,N_2883,N_2549);
or U3763 (N_3763,N_2956,N_2988);
or U3764 (N_3764,N_2226,N_2590);
nand U3765 (N_3765,N_2838,N_2760);
or U3766 (N_3766,N_2830,N_2247);
or U3767 (N_3767,N_2460,N_2155);
and U3768 (N_3768,N_2451,N_2805);
or U3769 (N_3769,N_2150,N_2134);
xnor U3770 (N_3770,N_2290,N_2837);
nand U3771 (N_3771,N_2773,N_2106);
xnor U3772 (N_3772,N_2677,N_2696);
and U3773 (N_3773,N_2892,N_2433);
nor U3774 (N_3774,N_2622,N_2940);
and U3775 (N_3775,N_2320,N_2098);
nand U3776 (N_3776,N_2129,N_2086);
nor U3777 (N_3777,N_2046,N_2981);
nand U3778 (N_3778,N_2559,N_2517);
nand U3779 (N_3779,N_2783,N_2352);
nand U3780 (N_3780,N_2095,N_2266);
nor U3781 (N_3781,N_2830,N_2240);
nand U3782 (N_3782,N_2274,N_2558);
nand U3783 (N_3783,N_2629,N_2298);
xor U3784 (N_3784,N_2563,N_2895);
or U3785 (N_3785,N_2628,N_2364);
or U3786 (N_3786,N_2449,N_2292);
nand U3787 (N_3787,N_2023,N_2241);
or U3788 (N_3788,N_2939,N_2561);
or U3789 (N_3789,N_2492,N_2075);
nor U3790 (N_3790,N_2124,N_2882);
and U3791 (N_3791,N_2933,N_2122);
nor U3792 (N_3792,N_2171,N_2749);
or U3793 (N_3793,N_2527,N_2477);
and U3794 (N_3794,N_2062,N_2550);
nor U3795 (N_3795,N_2728,N_2310);
and U3796 (N_3796,N_2639,N_2346);
xor U3797 (N_3797,N_2824,N_2722);
or U3798 (N_3798,N_2586,N_2305);
nor U3799 (N_3799,N_2493,N_2261);
and U3800 (N_3800,N_2792,N_2242);
or U3801 (N_3801,N_2820,N_2218);
or U3802 (N_3802,N_2864,N_2538);
nor U3803 (N_3803,N_2865,N_2647);
nand U3804 (N_3804,N_2091,N_2933);
xor U3805 (N_3805,N_2638,N_2849);
or U3806 (N_3806,N_2517,N_2016);
and U3807 (N_3807,N_2126,N_2304);
nor U3808 (N_3808,N_2253,N_2485);
and U3809 (N_3809,N_2459,N_2940);
or U3810 (N_3810,N_2541,N_2821);
nand U3811 (N_3811,N_2400,N_2042);
nor U3812 (N_3812,N_2470,N_2480);
nor U3813 (N_3813,N_2162,N_2907);
xnor U3814 (N_3814,N_2605,N_2017);
or U3815 (N_3815,N_2590,N_2689);
xor U3816 (N_3816,N_2948,N_2394);
nor U3817 (N_3817,N_2048,N_2227);
or U3818 (N_3818,N_2755,N_2676);
or U3819 (N_3819,N_2285,N_2525);
nand U3820 (N_3820,N_2489,N_2654);
nand U3821 (N_3821,N_2839,N_2546);
nor U3822 (N_3822,N_2778,N_2222);
xnor U3823 (N_3823,N_2914,N_2537);
nand U3824 (N_3824,N_2262,N_2699);
xnor U3825 (N_3825,N_2348,N_2615);
or U3826 (N_3826,N_2314,N_2058);
and U3827 (N_3827,N_2290,N_2194);
xor U3828 (N_3828,N_2797,N_2653);
or U3829 (N_3829,N_2204,N_2724);
and U3830 (N_3830,N_2835,N_2111);
xor U3831 (N_3831,N_2005,N_2276);
nand U3832 (N_3832,N_2918,N_2787);
nor U3833 (N_3833,N_2772,N_2828);
nor U3834 (N_3834,N_2137,N_2476);
nor U3835 (N_3835,N_2295,N_2673);
nand U3836 (N_3836,N_2036,N_2774);
nor U3837 (N_3837,N_2314,N_2439);
xor U3838 (N_3838,N_2063,N_2354);
and U3839 (N_3839,N_2878,N_2096);
xor U3840 (N_3840,N_2222,N_2255);
nor U3841 (N_3841,N_2694,N_2397);
or U3842 (N_3842,N_2678,N_2079);
xor U3843 (N_3843,N_2049,N_2647);
nand U3844 (N_3844,N_2123,N_2291);
and U3845 (N_3845,N_2754,N_2988);
nor U3846 (N_3846,N_2118,N_2066);
and U3847 (N_3847,N_2028,N_2628);
xor U3848 (N_3848,N_2423,N_2040);
nor U3849 (N_3849,N_2995,N_2417);
or U3850 (N_3850,N_2449,N_2372);
nor U3851 (N_3851,N_2187,N_2716);
nand U3852 (N_3852,N_2865,N_2109);
nor U3853 (N_3853,N_2105,N_2078);
nand U3854 (N_3854,N_2396,N_2050);
or U3855 (N_3855,N_2966,N_2794);
nand U3856 (N_3856,N_2804,N_2426);
and U3857 (N_3857,N_2469,N_2581);
and U3858 (N_3858,N_2126,N_2588);
and U3859 (N_3859,N_2016,N_2513);
xnor U3860 (N_3860,N_2229,N_2072);
nand U3861 (N_3861,N_2328,N_2897);
or U3862 (N_3862,N_2118,N_2181);
nand U3863 (N_3863,N_2043,N_2557);
nor U3864 (N_3864,N_2928,N_2605);
and U3865 (N_3865,N_2502,N_2018);
nand U3866 (N_3866,N_2416,N_2922);
nand U3867 (N_3867,N_2246,N_2997);
and U3868 (N_3868,N_2124,N_2070);
and U3869 (N_3869,N_2055,N_2155);
nand U3870 (N_3870,N_2219,N_2175);
nand U3871 (N_3871,N_2857,N_2823);
and U3872 (N_3872,N_2386,N_2124);
or U3873 (N_3873,N_2360,N_2953);
or U3874 (N_3874,N_2141,N_2417);
or U3875 (N_3875,N_2950,N_2331);
nand U3876 (N_3876,N_2114,N_2824);
and U3877 (N_3877,N_2029,N_2039);
or U3878 (N_3878,N_2568,N_2721);
nor U3879 (N_3879,N_2117,N_2684);
and U3880 (N_3880,N_2190,N_2351);
nor U3881 (N_3881,N_2451,N_2430);
or U3882 (N_3882,N_2319,N_2292);
nor U3883 (N_3883,N_2517,N_2368);
xor U3884 (N_3884,N_2061,N_2877);
nor U3885 (N_3885,N_2660,N_2223);
nand U3886 (N_3886,N_2829,N_2809);
nor U3887 (N_3887,N_2913,N_2608);
or U3888 (N_3888,N_2114,N_2164);
nand U3889 (N_3889,N_2778,N_2444);
nand U3890 (N_3890,N_2980,N_2411);
and U3891 (N_3891,N_2061,N_2608);
nor U3892 (N_3892,N_2815,N_2167);
or U3893 (N_3893,N_2844,N_2261);
or U3894 (N_3894,N_2003,N_2120);
nor U3895 (N_3895,N_2680,N_2658);
nand U3896 (N_3896,N_2859,N_2926);
and U3897 (N_3897,N_2351,N_2420);
xor U3898 (N_3898,N_2877,N_2609);
nor U3899 (N_3899,N_2502,N_2274);
or U3900 (N_3900,N_2424,N_2345);
xnor U3901 (N_3901,N_2568,N_2779);
or U3902 (N_3902,N_2501,N_2902);
nand U3903 (N_3903,N_2987,N_2645);
and U3904 (N_3904,N_2798,N_2433);
nor U3905 (N_3905,N_2212,N_2793);
or U3906 (N_3906,N_2433,N_2054);
and U3907 (N_3907,N_2677,N_2193);
or U3908 (N_3908,N_2336,N_2666);
and U3909 (N_3909,N_2550,N_2405);
and U3910 (N_3910,N_2803,N_2101);
or U3911 (N_3911,N_2951,N_2367);
or U3912 (N_3912,N_2180,N_2130);
nor U3913 (N_3913,N_2190,N_2006);
nor U3914 (N_3914,N_2080,N_2210);
nand U3915 (N_3915,N_2018,N_2591);
or U3916 (N_3916,N_2187,N_2375);
and U3917 (N_3917,N_2592,N_2485);
and U3918 (N_3918,N_2533,N_2275);
nor U3919 (N_3919,N_2229,N_2904);
nand U3920 (N_3920,N_2443,N_2368);
or U3921 (N_3921,N_2711,N_2365);
or U3922 (N_3922,N_2890,N_2379);
nor U3923 (N_3923,N_2351,N_2696);
xnor U3924 (N_3924,N_2023,N_2348);
xor U3925 (N_3925,N_2246,N_2907);
or U3926 (N_3926,N_2783,N_2863);
and U3927 (N_3927,N_2934,N_2417);
xor U3928 (N_3928,N_2844,N_2297);
nor U3929 (N_3929,N_2640,N_2868);
or U3930 (N_3930,N_2374,N_2138);
and U3931 (N_3931,N_2186,N_2673);
or U3932 (N_3932,N_2300,N_2412);
nand U3933 (N_3933,N_2849,N_2581);
xor U3934 (N_3934,N_2252,N_2298);
and U3935 (N_3935,N_2605,N_2221);
nand U3936 (N_3936,N_2781,N_2168);
or U3937 (N_3937,N_2380,N_2525);
or U3938 (N_3938,N_2611,N_2538);
and U3939 (N_3939,N_2572,N_2630);
and U3940 (N_3940,N_2931,N_2180);
and U3941 (N_3941,N_2130,N_2991);
and U3942 (N_3942,N_2075,N_2160);
nor U3943 (N_3943,N_2724,N_2050);
or U3944 (N_3944,N_2775,N_2992);
or U3945 (N_3945,N_2634,N_2069);
and U3946 (N_3946,N_2799,N_2826);
nand U3947 (N_3947,N_2530,N_2828);
and U3948 (N_3948,N_2108,N_2953);
nor U3949 (N_3949,N_2285,N_2650);
or U3950 (N_3950,N_2098,N_2553);
or U3951 (N_3951,N_2424,N_2353);
nand U3952 (N_3952,N_2372,N_2245);
or U3953 (N_3953,N_2137,N_2861);
or U3954 (N_3954,N_2925,N_2276);
and U3955 (N_3955,N_2001,N_2424);
or U3956 (N_3956,N_2021,N_2032);
xnor U3957 (N_3957,N_2033,N_2824);
or U3958 (N_3958,N_2050,N_2948);
xnor U3959 (N_3959,N_2780,N_2802);
nand U3960 (N_3960,N_2352,N_2274);
nor U3961 (N_3961,N_2946,N_2592);
nand U3962 (N_3962,N_2750,N_2752);
and U3963 (N_3963,N_2227,N_2276);
and U3964 (N_3964,N_2623,N_2616);
or U3965 (N_3965,N_2679,N_2573);
or U3966 (N_3966,N_2264,N_2646);
nor U3967 (N_3967,N_2602,N_2505);
and U3968 (N_3968,N_2239,N_2690);
nor U3969 (N_3969,N_2634,N_2968);
nor U3970 (N_3970,N_2518,N_2247);
nand U3971 (N_3971,N_2214,N_2978);
xnor U3972 (N_3972,N_2304,N_2231);
nand U3973 (N_3973,N_2613,N_2306);
xor U3974 (N_3974,N_2772,N_2078);
nor U3975 (N_3975,N_2313,N_2508);
nand U3976 (N_3976,N_2540,N_2481);
and U3977 (N_3977,N_2305,N_2024);
and U3978 (N_3978,N_2559,N_2070);
and U3979 (N_3979,N_2934,N_2566);
or U3980 (N_3980,N_2572,N_2954);
nand U3981 (N_3981,N_2211,N_2525);
nor U3982 (N_3982,N_2729,N_2296);
or U3983 (N_3983,N_2008,N_2053);
and U3984 (N_3984,N_2359,N_2477);
nor U3985 (N_3985,N_2166,N_2004);
and U3986 (N_3986,N_2751,N_2512);
or U3987 (N_3987,N_2636,N_2359);
and U3988 (N_3988,N_2487,N_2107);
nand U3989 (N_3989,N_2865,N_2080);
nor U3990 (N_3990,N_2521,N_2651);
or U3991 (N_3991,N_2794,N_2500);
nor U3992 (N_3992,N_2309,N_2135);
nand U3993 (N_3993,N_2687,N_2995);
and U3994 (N_3994,N_2458,N_2389);
nand U3995 (N_3995,N_2262,N_2422);
nand U3996 (N_3996,N_2047,N_2705);
nor U3997 (N_3997,N_2221,N_2285);
nand U3998 (N_3998,N_2246,N_2070);
nand U3999 (N_3999,N_2501,N_2384);
xnor U4000 (N_4000,N_3855,N_3265);
and U4001 (N_4001,N_3842,N_3527);
nand U4002 (N_4002,N_3726,N_3309);
or U4003 (N_4003,N_3511,N_3390);
nor U4004 (N_4004,N_3935,N_3270);
nor U4005 (N_4005,N_3933,N_3257);
or U4006 (N_4006,N_3525,N_3275);
or U4007 (N_4007,N_3762,N_3023);
or U4008 (N_4008,N_3343,N_3621);
and U4009 (N_4009,N_3807,N_3733);
nand U4010 (N_4010,N_3712,N_3802);
or U4011 (N_4011,N_3383,N_3963);
and U4012 (N_4012,N_3812,N_3339);
nor U4013 (N_4013,N_3239,N_3510);
or U4014 (N_4014,N_3185,N_3434);
or U4015 (N_4015,N_3086,N_3586);
nand U4016 (N_4016,N_3548,N_3054);
nand U4017 (N_4017,N_3610,N_3024);
and U4018 (N_4018,N_3014,N_3638);
xnor U4019 (N_4019,N_3979,N_3497);
or U4020 (N_4020,N_3908,N_3388);
nand U4021 (N_4021,N_3405,N_3191);
nor U4022 (N_4022,N_3096,N_3036);
and U4023 (N_4023,N_3231,N_3269);
and U4024 (N_4024,N_3001,N_3091);
or U4025 (N_4025,N_3941,N_3382);
xnor U4026 (N_4026,N_3290,N_3385);
nor U4027 (N_4027,N_3272,N_3079);
nor U4028 (N_4028,N_3753,N_3125);
nor U4029 (N_4029,N_3703,N_3460);
or U4030 (N_4030,N_3420,N_3003);
nor U4031 (N_4031,N_3861,N_3324);
nand U4032 (N_4032,N_3528,N_3260);
or U4033 (N_4033,N_3496,N_3954);
and U4034 (N_4034,N_3653,N_3461);
nor U4035 (N_4035,N_3619,N_3321);
and U4036 (N_4036,N_3505,N_3648);
nor U4037 (N_4037,N_3336,N_3256);
nor U4038 (N_4038,N_3323,N_3531);
nor U4039 (N_4039,N_3667,N_3217);
and U4040 (N_4040,N_3845,N_3064);
or U4041 (N_4041,N_3650,N_3234);
nand U4042 (N_4042,N_3333,N_3316);
or U4043 (N_4043,N_3216,N_3924);
xor U4044 (N_4044,N_3996,N_3228);
nor U4045 (N_4045,N_3784,N_3325);
or U4046 (N_4046,N_3870,N_3571);
nand U4047 (N_4047,N_3771,N_3347);
nor U4048 (N_4048,N_3411,N_3917);
nor U4049 (N_4049,N_3182,N_3053);
xor U4050 (N_4050,N_3635,N_3459);
xor U4051 (N_4051,N_3971,N_3015);
or U4052 (N_4052,N_3865,N_3618);
or U4053 (N_4053,N_3439,N_3089);
and U4054 (N_4054,N_3783,N_3132);
and U4055 (N_4055,N_3800,N_3428);
nand U4056 (N_4056,N_3193,N_3945);
or U4057 (N_4057,N_3106,N_3168);
or U4058 (N_4058,N_3984,N_3544);
and U4059 (N_4059,N_3210,N_3970);
nor U4060 (N_4060,N_3208,N_3821);
and U4061 (N_4061,N_3986,N_3551);
nand U4062 (N_4062,N_3837,N_3765);
or U4063 (N_4063,N_3547,N_3848);
nor U4064 (N_4064,N_3533,N_3287);
nand U4065 (N_4065,N_3903,N_3878);
nand U4066 (N_4066,N_3706,N_3133);
and U4067 (N_4067,N_3699,N_3378);
and U4068 (N_4068,N_3264,N_3647);
or U4069 (N_4069,N_3490,N_3172);
or U4070 (N_4070,N_3016,N_3143);
or U4071 (N_4071,N_3696,N_3523);
xnor U4072 (N_4072,N_3501,N_3568);
nor U4073 (N_4073,N_3404,N_3302);
or U4074 (N_4074,N_3175,N_3748);
or U4075 (N_4075,N_3009,N_3072);
or U4076 (N_4076,N_3352,N_3118);
nor U4077 (N_4077,N_3432,N_3487);
nor U4078 (N_4078,N_3906,N_3285);
nand U4079 (N_4079,N_3534,N_3214);
or U4080 (N_4080,N_3441,N_3854);
nand U4081 (N_4081,N_3494,N_3763);
and U4082 (N_4082,N_3661,N_3622);
xnor U4083 (N_4083,N_3081,N_3196);
and U4084 (N_4084,N_3169,N_3976);
and U4085 (N_4085,N_3259,N_3319);
nand U4086 (N_4086,N_3847,N_3101);
nor U4087 (N_4087,N_3593,N_3374);
nor U4088 (N_4088,N_3164,N_3499);
and U4089 (N_4089,N_3330,N_3857);
or U4090 (N_4090,N_3680,N_3102);
or U4091 (N_4091,N_3209,N_3981);
nand U4092 (N_4092,N_3485,N_3359);
nor U4093 (N_4093,N_3768,N_3243);
and U4094 (N_4094,N_3148,N_3590);
or U4095 (N_4095,N_3504,N_3577);
or U4096 (N_4096,N_3949,N_3598);
nor U4097 (N_4097,N_3017,N_3021);
nand U4098 (N_4098,N_3368,N_3881);
and U4099 (N_4099,N_3395,N_3815);
or U4100 (N_4100,N_3393,N_3891);
nor U4101 (N_4101,N_3786,N_3515);
or U4102 (N_4102,N_3227,N_3357);
xor U4103 (N_4103,N_3421,N_3772);
or U4104 (N_4104,N_3745,N_3008);
and U4105 (N_4105,N_3474,N_3962);
and U4106 (N_4106,N_3298,N_3137);
xnor U4107 (N_4107,N_3273,N_3427);
and U4108 (N_4108,N_3866,N_3927);
or U4109 (N_4109,N_3263,N_3649);
and U4110 (N_4110,N_3223,N_3714);
and U4111 (N_4111,N_3034,N_3115);
xnor U4112 (N_4112,N_3922,N_3005);
or U4113 (N_4113,N_3197,N_3671);
or U4114 (N_4114,N_3462,N_3369);
and U4115 (N_4115,N_3360,N_3039);
xnor U4116 (N_4116,N_3757,N_3261);
and U4117 (N_4117,N_3391,N_3977);
or U4118 (N_4118,N_3473,N_3356);
nand U4119 (N_4119,N_3686,N_3503);
nor U4120 (N_4120,N_3061,N_3678);
or U4121 (N_4121,N_3312,N_3565);
or U4122 (N_4122,N_3964,N_3447);
and U4123 (N_4123,N_3892,N_3297);
nor U4124 (N_4124,N_3122,N_3303);
or U4125 (N_4125,N_3063,N_3723);
or U4126 (N_4126,N_3521,N_3351);
or U4127 (N_4127,N_3479,N_3355);
nor U4128 (N_4128,N_3932,N_3628);
nor U4129 (N_4129,N_3431,N_3232);
nand U4130 (N_4130,N_3846,N_3512);
nor U4131 (N_4131,N_3481,N_3161);
nand U4132 (N_4132,N_3721,N_3119);
and U4133 (N_4133,N_3370,N_3526);
and U4134 (N_4134,N_3684,N_3727);
xnor U4135 (N_4135,N_3300,N_3978);
nor U4136 (N_4136,N_3044,N_3394);
and U4137 (N_4137,N_3792,N_3074);
and U4138 (N_4138,N_3464,N_3448);
and U4139 (N_4139,N_3488,N_3093);
and U4140 (N_4140,N_3245,N_3609);
or U4141 (N_4141,N_3444,N_3280);
and U4142 (N_4142,N_3952,N_3247);
xnor U4143 (N_4143,N_3560,N_3830);
and U4144 (N_4144,N_3697,N_3237);
nand U4145 (N_4145,N_3135,N_3946);
xor U4146 (N_4146,N_3435,N_3047);
xor U4147 (N_4147,N_3959,N_3045);
and U4148 (N_4148,N_3968,N_3563);
and U4149 (N_4149,N_3810,N_3822);
xor U4150 (N_4150,N_3990,N_3651);
nor U4151 (N_4151,N_3178,N_3665);
and U4152 (N_4152,N_3304,N_3371);
and U4153 (N_4153,N_3203,N_3708);
nor U4154 (N_4154,N_3951,N_3163);
and U4155 (N_4155,N_3989,N_3729);
or U4156 (N_4156,N_3450,N_3871);
nand U4157 (N_4157,N_3443,N_3070);
or U4158 (N_4158,N_3215,N_3670);
xnor U4159 (N_4159,N_3353,N_3627);
or U4160 (N_4160,N_3088,N_3082);
nor U4161 (N_4161,N_3475,N_3852);
nor U4162 (N_4162,N_3630,N_3159);
and U4163 (N_4163,N_3415,N_3255);
or U4164 (N_4164,N_3910,N_3246);
and U4165 (N_4165,N_3999,N_3307);
and U4166 (N_4166,N_3226,N_3294);
nor U4167 (N_4167,N_3655,N_3798);
nor U4168 (N_4168,N_3809,N_3406);
nand U4169 (N_4169,N_3037,N_3124);
and U4170 (N_4170,N_3436,N_3035);
nor U4171 (N_4171,N_3704,N_3419);
and U4172 (N_4172,N_3885,N_3663);
nand U4173 (N_4173,N_3399,N_3535);
nand U4174 (N_4174,N_3736,N_3085);
nor U4175 (N_4175,N_3506,N_3555);
xnor U4176 (N_4176,N_3914,N_3972);
nor U4177 (N_4177,N_3123,N_3605);
nor U4178 (N_4178,N_3840,N_3335);
nand U4179 (N_4179,N_3283,N_3816);
nand U4180 (N_4180,N_3337,N_3179);
nor U4181 (N_4181,N_3195,N_3907);
nand U4182 (N_4182,N_3755,N_3423);
nor U4183 (N_4183,N_3207,N_3000);
nand U4184 (N_4184,N_3416,N_3817);
nor U4185 (N_4185,N_3502,N_3863);
or U4186 (N_4186,N_3716,N_3626);
and U4187 (N_4187,N_3579,N_3874);
or U4188 (N_4188,N_3679,N_3578);
or U4189 (N_4189,N_3931,N_3732);
nand U4190 (N_4190,N_3090,N_3094);
and U4191 (N_4191,N_3925,N_3737);
xor U4192 (N_4192,N_3147,N_3904);
nor U4193 (N_4193,N_3136,N_3584);
and U4194 (N_4194,N_3340,N_3022);
or U4195 (N_4195,N_3095,N_3026);
nor U4196 (N_4196,N_3785,N_3741);
nor U4197 (N_4197,N_3433,N_3929);
xnor U4198 (N_4198,N_3545,N_3345);
and U4199 (N_4199,N_3664,N_3672);
nor U4200 (N_4200,N_3953,N_3915);
or U4201 (N_4201,N_3957,N_3117);
nand U4202 (N_4202,N_3358,N_3100);
nor U4203 (N_4203,N_3167,N_3770);
nor U4204 (N_4204,N_3581,N_3660);
or U4205 (N_4205,N_3128,N_3240);
xnor U4206 (N_4206,N_3398,N_3559);
xnor U4207 (N_4207,N_3078,N_3400);
nor U4208 (N_4208,N_3077,N_3675);
or U4209 (N_4209,N_3731,N_3975);
and U4210 (N_4210,N_3087,N_3342);
nor U4211 (N_4211,N_3508,N_3218);
nand U4212 (N_4212,N_3625,N_3006);
or U4213 (N_4213,N_3445,N_3900);
nor U4214 (N_4214,N_3381,N_3206);
nor U4215 (N_4215,N_3872,N_3198);
xnor U4216 (N_4216,N_3537,N_3774);
or U4217 (N_4217,N_3793,N_3028);
or U4218 (N_4218,N_3614,N_3029);
and U4219 (N_4219,N_3166,N_3564);
nand U4220 (N_4220,N_3483,N_3902);
nand U4221 (N_4221,N_3707,N_3219);
and U4222 (N_4222,N_3677,N_3636);
and U4223 (N_4223,N_3794,N_3552);
nor U4224 (N_4224,N_3562,N_3594);
nand U4225 (N_4225,N_3509,N_3826);
xor U4226 (N_4226,N_3131,N_3105);
or U4227 (N_4227,N_3367,N_3595);
nand U4228 (N_4228,N_3739,N_3827);
or U4229 (N_4229,N_3138,N_3403);
or U4230 (N_4230,N_3414,N_3764);
nor U4231 (N_4231,N_3801,N_3489);
xnor U4232 (N_4232,N_3442,N_3993);
nor U4233 (N_4233,N_3181,N_3624);
nor U4234 (N_4234,N_3918,N_3629);
and U4235 (N_4235,N_3928,N_3380);
or U4236 (N_4236,N_3306,N_3437);
nand U4237 (N_4237,N_3230,N_3923);
nor U4238 (N_4238,N_3010,N_3580);
or U4239 (N_4239,N_3289,N_3311);
and U4240 (N_4240,N_3788,N_3387);
and U4241 (N_4241,N_3710,N_3720);
and U4242 (N_4242,N_3153,N_3899);
and U4243 (N_4243,N_3170,N_3401);
and U4244 (N_4244,N_3517,N_3887);
xnor U4245 (N_4245,N_3637,N_3640);
nor U4246 (N_4246,N_3540,N_3092);
xor U4247 (N_4247,N_3268,N_3066);
or U4248 (N_4248,N_3282,N_3700);
or U4249 (N_4249,N_3144,N_3204);
or U4250 (N_4250,N_3747,N_3835);
or U4251 (N_4251,N_3645,N_3913);
and U4252 (N_4252,N_3575,N_3032);
nor U4253 (N_4253,N_3769,N_3690);
nand U4254 (N_4254,N_3813,N_3858);
xor U4255 (N_4255,N_3281,N_3484);
nor U4256 (N_4256,N_3749,N_3286);
or U4257 (N_4257,N_3472,N_3519);
or U4258 (N_4258,N_3375,N_3836);
or U4259 (N_4259,N_3338,N_3354);
and U4260 (N_4260,N_3500,N_3724);
xnor U4261 (N_4261,N_3599,N_3520);
and U4262 (N_4262,N_3705,N_3961);
nor U4263 (N_4263,N_3186,N_3002);
nand U4264 (N_4264,N_3825,N_3960);
nor U4265 (N_4265,N_3065,N_3759);
nor U4266 (N_4266,N_3112,N_3740);
or U4267 (N_4267,N_3220,N_3572);
xnor U4268 (N_4268,N_3947,N_3142);
nand U4269 (N_4269,N_3040,N_3602);
or U4270 (N_4270,N_3585,N_3253);
and U4271 (N_4271,N_3277,N_3372);
xor U4272 (N_4272,N_3799,N_3591);
nand U4273 (N_4273,N_3617,N_3573);
nand U4274 (N_4274,N_3266,N_3554);
xnor U4275 (N_4275,N_3344,N_3069);
nand U4276 (N_4276,N_3911,N_3407);
and U4277 (N_4277,N_3430,N_3735);
or U4278 (N_4278,N_3939,N_3200);
nand U4279 (N_4279,N_3362,N_3693);
nor U4280 (N_4280,N_3222,N_3980);
and U4281 (N_4281,N_3983,N_3652);
and U4282 (N_4282,N_3291,N_3099);
nand U4283 (N_4283,N_3901,N_3944);
nor U4284 (N_4284,N_3058,N_3296);
nor U4285 (N_4285,N_3814,N_3542);
nand U4286 (N_4286,N_3558,N_3828);
nand U4287 (N_4287,N_3030,N_3734);
and U4288 (N_4288,N_3666,N_3498);
nor U4289 (N_4289,N_3982,N_3738);
or U4290 (N_4290,N_3715,N_3429);
and U4291 (N_4291,N_3880,N_3600);
or U4292 (N_4292,N_3596,N_3157);
nand U4293 (N_4293,N_3644,N_3350);
nor U4294 (N_4294,N_3379,N_3491);
nor U4295 (N_4295,N_3725,N_3940);
and U4296 (N_4296,N_3673,N_3546);
or U4297 (N_4297,N_3152,N_3315);
nor U4298 (N_4298,N_3188,N_3458);
nor U4299 (N_4299,N_3176,N_3987);
nand U4300 (N_4300,N_3466,N_3576);
nand U4301 (N_4301,N_3041,N_3589);
and U4302 (N_4302,N_3937,N_3249);
nor U4303 (N_4303,N_3597,N_3930);
or U4304 (N_4304,N_3080,N_3662);
nor U4305 (N_4305,N_3995,N_3373);
and U4306 (N_4306,N_3305,N_3781);
or U4307 (N_4307,N_3121,N_3129);
nor U4308 (N_4308,N_3657,N_3888);
nand U4309 (N_4309,N_3921,N_3860);
nand U4310 (N_4310,N_3756,N_3364);
or U4311 (N_4311,N_3334,N_3284);
and U4312 (N_4312,N_3695,N_3412);
and U4313 (N_4313,N_3884,N_3746);
and U4314 (N_4314,N_3805,N_3457);
nand U4315 (N_4315,N_3912,N_3248);
xnor U4316 (N_4316,N_3139,N_3165);
nor U4317 (N_4317,N_3482,N_3654);
nor U4318 (N_4318,N_3177,N_3849);
or U4319 (N_4319,N_3114,N_3408);
or U4320 (N_4320,N_3212,N_3539);
and U4321 (N_4321,N_3251,N_3583);
nor U4322 (N_4322,N_3057,N_3109);
nor U4323 (N_4323,N_3623,N_3318);
nand U4324 (N_4324,N_3702,N_3905);
nor U4325 (N_4325,N_3894,N_3766);
xnor U4326 (N_4326,N_3767,N_3711);
nand U4327 (N_4327,N_3942,N_3567);
nand U4328 (N_4328,N_3607,N_3116);
nor U4329 (N_4329,N_3145,N_3553);
nor U4330 (N_4330,N_3004,N_3850);
nand U4331 (N_4331,N_3668,N_3998);
nor U4332 (N_4332,N_3997,N_3377);
nand U4333 (N_4333,N_3919,N_3031);
nand U4334 (N_4334,N_3829,N_3646);
or U4335 (N_4335,N_3779,N_3516);
nand U4336 (N_4336,N_3127,N_3752);
or U4337 (N_4337,N_3742,N_3582);
or U4338 (N_4338,N_3634,N_3110);
nand U4339 (N_4339,N_3659,N_3244);
or U4340 (N_4340,N_3824,N_3950);
and U4341 (N_4341,N_3465,N_3279);
or U4342 (N_4342,N_3478,N_3224);
and U4343 (N_4343,N_3851,N_3760);
nand U4344 (N_4344,N_3310,N_3238);
and U4345 (N_4345,N_3787,N_3068);
or U4346 (N_4346,N_3313,N_3233);
and U4347 (N_4347,N_3758,N_3754);
xor U4348 (N_4348,N_3038,N_3876);
nand U4349 (N_4349,N_3055,N_3862);
or U4350 (N_4350,N_3292,N_3570);
nor U4351 (N_4351,N_3477,N_3189);
nor U4352 (N_4352,N_3916,N_3751);
and U4353 (N_4353,N_3056,N_3409);
or U4354 (N_4354,N_3073,N_3422);
nand U4355 (N_4355,N_3790,N_3683);
nor U4356 (N_4356,N_3909,N_3797);
nand U4357 (N_4357,N_3839,N_3926);
and U4358 (N_4358,N_3384,N_3789);
nand U4359 (N_4359,N_3322,N_3823);
nand U4360 (N_4360,N_3027,N_3761);
nor U4361 (N_4361,N_3833,N_3867);
and U4362 (N_4362,N_3469,N_3187);
and U4363 (N_4363,N_3103,N_3782);
nor U4364 (N_4364,N_3843,N_3184);
xor U4365 (N_4365,N_3113,N_3241);
and U4366 (N_4366,N_3020,N_3150);
or U4367 (N_4367,N_3205,N_3966);
nor U4368 (N_4368,N_3897,N_3084);
and U4369 (N_4369,N_3221,N_3898);
nor U4370 (N_4370,N_3943,N_3561);
nand U4371 (N_4371,N_3549,N_3608);
or U4372 (N_4372,N_3493,N_3804);
or U4373 (N_4373,N_3363,N_3744);
and U4374 (N_4374,N_3495,N_3013);
nor U4375 (N_4375,N_3603,N_3098);
or U4376 (N_4376,N_3691,N_3936);
nor U4377 (N_4377,N_3076,N_3397);
and U4378 (N_4378,N_3180,N_3777);
or U4379 (N_4379,N_3620,N_3417);
and U4380 (N_4380,N_3719,N_3956);
nor U4381 (N_4381,N_3656,N_3274);
and U4382 (N_4382,N_3601,N_3538);
or U4383 (N_4383,N_3969,N_3455);
or U4384 (N_4384,N_3875,N_3468);
or U4385 (N_4385,N_3938,N_3856);
nor U4386 (N_4386,N_3514,N_3868);
nor U4387 (N_4387,N_3588,N_3155);
and U4388 (N_4388,N_3183,N_3262);
nor U4389 (N_4389,N_3994,N_3955);
nand U4390 (N_4390,N_3832,N_3235);
nand U4391 (N_4391,N_3470,N_3242);
or U4392 (N_4392,N_3791,N_3413);
nand U4393 (N_4393,N_3418,N_3574);
nor U4394 (N_4394,N_3225,N_3778);
nand U4395 (N_4395,N_3471,N_3518);
or U4396 (N_4396,N_3844,N_3171);
or U4397 (N_4397,N_3033,N_3154);
xor U4398 (N_4398,N_3326,N_3258);
and U4399 (N_4399,N_3965,N_3201);
and U4400 (N_4400,N_3838,N_3107);
nand U4401 (N_4401,N_3252,N_3365);
nor U4402 (N_4402,N_3202,N_3859);
nand U4403 (N_4403,N_3713,N_3557);
nand U4404 (N_4404,N_3346,N_3879);
nor U4405 (N_4405,N_3633,N_3543);
nor U4406 (N_4406,N_3893,N_3920);
nor U4407 (N_4407,N_3775,N_3271);
nand U4408 (N_4408,N_3709,N_3730);
or U4409 (N_4409,N_3612,N_3604);
nor U4410 (N_4410,N_3873,N_3454);
xor U4411 (N_4411,N_3146,N_3062);
or U4412 (N_4412,N_3361,N_3831);
nand U4413 (N_4413,N_3687,N_3948);
and U4414 (N_4414,N_3019,N_3111);
xnor U4415 (N_4415,N_3192,N_3295);
nand U4416 (N_4416,N_3140,N_3524);
nor U4417 (N_4417,N_3569,N_3018);
xnor U4418 (N_4418,N_3991,N_3190);
nor U4419 (N_4419,N_3476,N_3060);
nand U4420 (N_4420,N_3213,N_3550);
and U4421 (N_4421,N_3934,N_3425);
nand U4422 (N_4422,N_3049,N_3529);
nand U4423 (N_4423,N_3314,N_3194);
or U4424 (N_4424,N_3173,N_3007);
nor U4425 (N_4425,N_3278,N_3050);
and U4426 (N_4426,N_3149,N_3896);
xor U4427 (N_4427,N_3507,N_3808);
xor U4428 (N_4428,N_3676,N_3532);
nor U4429 (N_4429,N_3592,N_3890);
nand U4430 (N_4430,N_3452,N_3895);
nor U4431 (N_4431,N_3818,N_3349);
and U4432 (N_4432,N_3288,N_3083);
and U4433 (N_4433,N_3811,N_3126);
nor U4434 (N_4434,N_3396,N_3317);
or U4435 (N_4435,N_3834,N_3631);
nand U4436 (N_4436,N_3682,N_3642);
nor U4437 (N_4437,N_3780,N_3587);
and U4438 (N_4438,N_3632,N_3392);
and U4439 (N_4439,N_3877,N_3276);
xnor U4440 (N_4440,N_3566,N_3320);
and U4441 (N_4441,N_3685,N_3329);
or U4442 (N_4442,N_3681,N_3134);
nor U4443 (N_4443,N_3486,N_3615);
xnor U4444 (N_4444,N_3743,N_3042);
or U4445 (N_4445,N_3541,N_3536);
xnor U4446 (N_4446,N_3386,N_3236);
xnor U4447 (N_4447,N_3530,N_3698);
xor U4448 (N_4448,N_3160,N_3841);
and U4449 (N_4449,N_3067,N_3267);
nand U4450 (N_4450,N_3988,N_3426);
nand U4451 (N_4451,N_3331,N_3492);
nand U4452 (N_4452,N_3974,N_3104);
and U4453 (N_4453,N_3059,N_3299);
nand U4454 (N_4454,N_3046,N_3229);
nand U4455 (N_4455,N_3795,N_3641);
nor U4456 (N_4456,N_3701,N_3853);
or U4457 (N_4457,N_3440,N_3389);
nor U4458 (N_4458,N_3328,N_3438);
and U4459 (N_4459,N_3025,N_3011);
nand U4460 (N_4460,N_3130,N_3694);
nor U4461 (N_4461,N_3886,N_3410);
nand U4462 (N_4462,N_3453,N_3658);
or U4463 (N_4463,N_3556,N_3156);
and U4464 (N_4464,N_3480,N_3728);
or U4465 (N_4465,N_3254,N_3669);
nor U4466 (N_4466,N_3424,N_3674);
nand U4467 (N_4467,N_3446,N_3250);
nand U4468 (N_4468,N_3348,N_3864);
and U4469 (N_4469,N_3141,N_3819);
nand U4470 (N_4470,N_3613,N_3097);
nand U4471 (N_4471,N_3162,N_3075);
nand U4472 (N_4472,N_3451,N_3366);
nor U4473 (N_4473,N_3071,N_3985);
and U4474 (N_4474,N_3689,N_3750);
nor U4475 (N_4475,N_3151,N_3158);
nor U4476 (N_4476,N_3341,N_3958);
and U4477 (N_4477,N_3643,N_3611);
and U4478 (N_4478,N_3463,N_3051);
nand U4479 (N_4479,N_3717,N_3449);
nor U4480 (N_4480,N_3402,N_3327);
and U4481 (N_4481,N_3606,N_3803);
xnor U4482 (N_4482,N_3820,N_3688);
nand U4483 (N_4483,N_3522,N_3467);
nor U4484 (N_4484,N_3796,N_3174);
nand U4485 (N_4485,N_3211,N_3718);
nor U4486 (N_4486,N_3012,N_3332);
or U4487 (N_4487,N_3639,N_3967);
nor U4488 (N_4488,N_3048,N_3806);
nand U4489 (N_4489,N_3692,N_3973);
xor U4490 (N_4490,N_3722,N_3043);
nor U4491 (N_4491,N_3052,N_3513);
and U4492 (N_4492,N_3883,N_3199);
xor U4493 (N_4493,N_3776,N_3301);
and U4494 (N_4494,N_3376,N_3773);
nand U4495 (N_4495,N_3308,N_3992);
nand U4496 (N_4496,N_3120,N_3108);
nand U4497 (N_4497,N_3293,N_3889);
nor U4498 (N_4498,N_3869,N_3616);
nand U4499 (N_4499,N_3882,N_3456);
and U4500 (N_4500,N_3525,N_3174);
or U4501 (N_4501,N_3497,N_3809);
and U4502 (N_4502,N_3018,N_3072);
and U4503 (N_4503,N_3334,N_3838);
and U4504 (N_4504,N_3939,N_3639);
nor U4505 (N_4505,N_3630,N_3731);
xor U4506 (N_4506,N_3691,N_3529);
nor U4507 (N_4507,N_3421,N_3955);
or U4508 (N_4508,N_3726,N_3626);
and U4509 (N_4509,N_3211,N_3938);
nand U4510 (N_4510,N_3568,N_3491);
or U4511 (N_4511,N_3434,N_3946);
nand U4512 (N_4512,N_3880,N_3965);
and U4513 (N_4513,N_3994,N_3801);
nor U4514 (N_4514,N_3804,N_3613);
or U4515 (N_4515,N_3576,N_3951);
nor U4516 (N_4516,N_3848,N_3730);
nand U4517 (N_4517,N_3479,N_3697);
nor U4518 (N_4518,N_3897,N_3870);
nand U4519 (N_4519,N_3929,N_3710);
and U4520 (N_4520,N_3305,N_3317);
or U4521 (N_4521,N_3709,N_3796);
or U4522 (N_4522,N_3564,N_3041);
xor U4523 (N_4523,N_3926,N_3158);
and U4524 (N_4524,N_3574,N_3948);
nand U4525 (N_4525,N_3056,N_3996);
or U4526 (N_4526,N_3960,N_3680);
xnor U4527 (N_4527,N_3407,N_3486);
and U4528 (N_4528,N_3049,N_3408);
nor U4529 (N_4529,N_3817,N_3240);
nor U4530 (N_4530,N_3762,N_3615);
nor U4531 (N_4531,N_3727,N_3491);
nor U4532 (N_4532,N_3427,N_3008);
nor U4533 (N_4533,N_3386,N_3652);
xnor U4534 (N_4534,N_3576,N_3998);
and U4535 (N_4535,N_3775,N_3931);
or U4536 (N_4536,N_3490,N_3918);
xnor U4537 (N_4537,N_3913,N_3096);
and U4538 (N_4538,N_3194,N_3287);
nand U4539 (N_4539,N_3757,N_3483);
nand U4540 (N_4540,N_3598,N_3413);
nand U4541 (N_4541,N_3082,N_3417);
and U4542 (N_4542,N_3220,N_3797);
and U4543 (N_4543,N_3133,N_3661);
and U4544 (N_4544,N_3958,N_3770);
and U4545 (N_4545,N_3990,N_3449);
nand U4546 (N_4546,N_3300,N_3872);
or U4547 (N_4547,N_3816,N_3724);
and U4548 (N_4548,N_3323,N_3353);
or U4549 (N_4549,N_3535,N_3209);
nor U4550 (N_4550,N_3973,N_3381);
nor U4551 (N_4551,N_3412,N_3482);
nand U4552 (N_4552,N_3875,N_3381);
or U4553 (N_4553,N_3730,N_3147);
nor U4554 (N_4554,N_3402,N_3020);
and U4555 (N_4555,N_3494,N_3118);
nand U4556 (N_4556,N_3102,N_3571);
and U4557 (N_4557,N_3033,N_3690);
nand U4558 (N_4558,N_3835,N_3033);
and U4559 (N_4559,N_3454,N_3081);
nand U4560 (N_4560,N_3507,N_3024);
nor U4561 (N_4561,N_3168,N_3924);
nor U4562 (N_4562,N_3688,N_3629);
nor U4563 (N_4563,N_3280,N_3631);
nand U4564 (N_4564,N_3885,N_3606);
xor U4565 (N_4565,N_3409,N_3826);
nor U4566 (N_4566,N_3733,N_3380);
nand U4567 (N_4567,N_3160,N_3548);
nand U4568 (N_4568,N_3743,N_3088);
xnor U4569 (N_4569,N_3280,N_3057);
or U4570 (N_4570,N_3689,N_3010);
nand U4571 (N_4571,N_3944,N_3266);
and U4572 (N_4572,N_3104,N_3191);
xor U4573 (N_4573,N_3321,N_3965);
nor U4574 (N_4574,N_3450,N_3120);
and U4575 (N_4575,N_3892,N_3234);
nor U4576 (N_4576,N_3309,N_3270);
nand U4577 (N_4577,N_3959,N_3355);
and U4578 (N_4578,N_3652,N_3038);
and U4579 (N_4579,N_3308,N_3927);
and U4580 (N_4580,N_3162,N_3022);
or U4581 (N_4581,N_3905,N_3587);
or U4582 (N_4582,N_3498,N_3760);
nor U4583 (N_4583,N_3380,N_3771);
xor U4584 (N_4584,N_3323,N_3423);
or U4585 (N_4585,N_3612,N_3819);
nand U4586 (N_4586,N_3287,N_3854);
nand U4587 (N_4587,N_3103,N_3108);
nor U4588 (N_4588,N_3922,N_3635);
or U4589 (N_4589,N_3165,N_3295);
and U4590 (N_4590,N_3046,N_3796);
nand U4591 (N_4591,N_3602,N_3482);
xor U4592 (N_4592,N_3262,N_3076);
nor U4593 (N_4593,N_3969,N_3663);
nor U4594 (N_4594,N_3472,N_3029);
or U4595 (N_4595,N_3775,N_3518);
or U4596 (N_4596,N_3396,N_3385);
nand U4597 (N_4597,N_3597,N_3970);
or U4598 (N_4598,N_3471,N_3954);
nand U4599 (N_4599,N_3541,N_3454);
or U4600 (N_4600,N_3809,N_3938);
or U4601 (N_4601,N_3626,N_3464);
nor U4602 (N_4602,N_3834,N_3280);
and U4603 (N_4603,N_3572,N_3835);
nor U4604 (N_4604,N_3653,N_3552);
nor U4605 (N_4605,N_3699,N_3053);
and U4606 (N_4606,N_3690,N_3291);
nand U4607 (N_4607,N_3042,N_3635);
nor U4608 (N_4608,N_3405,N_3439);
xnor U4609 (N_4609,N_3428,N_3524);
and U4610 (N_4610,N_3193,N_3640);
and U4611 (N_4611,N_3939,N_3167);
or U4612 (N_4612,N_3589,N_3365);
xor U4613 (N_4613,N_3811,N_3651);
xnor U4614 (N_4614,N_3075,N_3488);
xnor U4615 (N_4615,N_3305,N_3166);
nand U4616 (N_4616,N_3254,N_3030);
nand U4617 (N_4617,N_3924,N_3413);
xnor U4618 (N_4618,N_3344,N_3917);
nand U4619 (N_4619,N_3575,N_3761);
and U4620 (N_4620,N_3192,N_3672);
nor U4621 (N_4621,N_3472,N_3415);
and U4622 (N_4622,N_3246,N_3948);
nor U4623 (N_4623,N_3945,N_3948);
nor U4624 (N_4624,N_3161,N_3275);
nand U4625 (N_4625,N_3007,N_3675);
or U4626 (N_4626,N_3736,N_3502);
and U4627 (N_4627,N_3589,N_3022);
nor U4628 (N_4628,N_3695,N_3110);
or U4629 (N_4629,N_3162,N_3246);
nand U4630 (N_4630,N_3609,N_3588);
xor U4631 (N_4631,N_3933,N_3394);
xnor U4632 (N_4632,N_3322,N_3957);
nand U4633 (N_4633,N_3653,N_3251);
nand U4634 (N_4634,N_3077,N_3829);
nor U4635 (N_4635,N_3242,N_3475);
nor U4636 (N_4636,N_3590,N_3367);
and U4637 (N_4637,N_3547,N_3510);
or U4638 (N_4638,N_3286,N_3689);
nor U4639 (N_4639,N_3602,N_3080);
or U4640 (N_4640,N_3048,N_3063);
nor U4641 (N_4641,N_3995,N_3498);
or U4642 (N_4642,N_3312,N_3379);
and U4643 (N_4643,N_3726,N_3509);
nand U4644 (N_4644,N_3003,N_3513);
nand U4645 (N_4645,N_3336,N_3246);
nand U4646 (N_4646,N_3121,N_3090);
xnor U4647 (N_4647,N_3710,N_3086);
or U4648 (N_4648,N_3669,N_3599);
nor U4649 (N_4649,N_3319,N_3669);
nand U4650 (N_4650,N_3974,N_3870);
nand U4651 (N_4651,N_3725,N_3675);
or U4652 (N_4652,N_3941,N_3666);
nor U4653 (N_4653,N_3076,N_3654);
or U4654 (N_4654,N_3854,N_3553);
or U4655 (N_4655,N_3501,N_3523);
nand U4656 (N_4656,N_3243,N_3844);
nand U4657 (N_4657,N_3824,N_3551);
xor U4658 (N_4658,N_3894,N_3302);
and U4659 (N_4659,N_3688,N_3576);
nor U4660 (N_4660,N_3324,N_3586);
and U4661 (N_4661,N_3868,N_3128);
nor U4662 (N_4662,N_3718,N_3821);
nor U4663 (N_4663,N_3171,N_3805);
nand U4664 (N_4664,N_3265,N_3959);
nor U4665 (N_4665,N_3173,N_3556);
nor U4666 (N_4666,N_3805,N_3790);
and U4667 (N_4667,N_3146,N_3387);
or U4668 (N_4668,N_3338,N_3517);
or U4669 (N_4669,N_3021,N_3776);
nor U4670 (N_4670,N_3235,N_3765);
or U4671 (N_4671,N_3275,N_3768);
nor U4672 (N_4672,N_3134,N_3645);
nand U4673 (N_4673,N_3019,N_3074);
nor U4674 (N_4674,N_3145,N_3946);
or U4675 (N_4675,N_3614,N_3303);
nor U4676 (N_4676,N_3153,N_3790);
nand U4677 (N_4677,N_3200,N_3170);
and U4678 (N_4678,N_3289,N_3350);
nand U4679 (N_4679,N_3726,N_3792);
nand U4680 (N_4680,N_3538,N_3805);
nor U4681 (N_4681,N_3565,N_3453);
or U4682 (N_4682,N_3926,N_3251);
and U4683 (N_4683,N_3581,N_3893);
nand U4684 (N_4684,N_3246,N_3464);
nor U4685 (N_4685,N_3846,N_3269);
nor U4686 (N_4686,N_3993,N_3544);
and U4687 (N_4687,N_3141,N_3635);
or U4688 (N_4688,N_3109,N_3787);
nor U4689 (N_4689,N_3392,N_3684);
nor U4690 (N_4690,N_3267,N_3680);
and U4691 (N_4691,N_3014,N_3895);
or U4692 (N_4692,N_3030,N_3182);
and U4693 (N_4693,N_3648,N_3687);
nor U4694 (N_4694,N_3330,N_3580);
nand U4695 (N_4695,N_3143,N_3318);
and U4696 (N_4696,N_3541,N_3041);
nand U4697 (N_4697,N_3144,N_3221);
and U4698 (N_4698,N_3676,N_3109);
and U4699 (N_4699,N_3627,N_3309);
and U4700 (N_4700,N_3371,N_3975);
xor U4701 (N_4701,N_3363,N_3228);
nand U4702 (N_4702,N_3282,N_3508);
and U4703 (N_4703,N_3395,N_3362);
xnor U4704 (N_4704,N_3641,N_3426);
nand U4705 (N_4705,N_3690,N_3027);
xnor U4706 (N_4706,N_3229,N_3825);
or U4707 (N_4707,N_3796,N_3816);
or U4708 (N_4708,N_3341,N_3120);
nor U4709 (N_4709,N_3524,N_3431);
and U4710 (N_4710,N_3802,N_3625);
or U4711 (N_4711,N_3039,N_3379);
nand U4712 (N_4712,N_3460,N_3912);
and U4713 (N_4713,N_3498,N_3240);
nand U4714 (N_4714,N_3749,N_3883);
or U4715 (N_4715,N_3908,N_3718);
nand U4716 (N_4716,N_3750,N_3551);
or U4717 (N_4717,N_3232,N_3587);
nor U4718 (N_4718,N_3840,N_3495);
nor U4719 (N_4719,N_3838,N_3494);
or U4720 (N_4720,N_3337,N_3150);
and U4721 (N_4721,N_3792,N_3205);
and U4722 (N_4722,N_3648,N_3144);
nand U4723 (N_4723,N_3699,N_3227);
and U4724 (N_4724,N_3642,N_3256);
nor U4725 (N_4725,N_3554,N_3759);
and U4726 (N_4726,N_3402,N_3059);
nor U4727 (N_4727,N_3672,N_3643);
nand U4728 (N_4728,N_3122,N_3053);
xnor U4729 (N_4729,N_3573,N_3142);
xnor U4730 (N_4730,N_3754,N_3675);
or U4731 (N_4731,N_3310,N_3788);
nor U4732 (N_4732,N_3061,N_3128);
and U4733 (N_4733,N_3706,N_3474);
nor U4734 (N_4734,N_3560,N_3081);
nand U4735 (N_4735,N_3418,N_3569);
or U4736 (N_4736,N_3548,N_3258);
nand U4737 (N_4737,N_3892,N_3998);
or U4738 (N_4738,N_3748,N_3986);
nor U4739 (N_4739,N_3496,N_3684);
and U4740 (N_4740,N_3698,N_3040);
nor U4741 (N_4741,N_3851,N_3501);
or U4742 (N_4742,N_3814,N_3367);
or U4743 (N_4743,N_3012,N_3903);
nand U4744 (N_4744,N_3160,N_3343);
nand U4745 (N_4745,N_3954,N_3713);
xnor U4746 (N_4746,N_3621,N_3506);
or U4747 (N_4747,N_3587,N_3147);
and U4748 (N_4748,N_3535,N_3501);
nand U4749 (N_4749,N_3498,N_3671);
or U4750 (N_4750,N_3571,N_3355);
nand U4751 (N_4751,N_3313,N_3252);
and U4752 (N_4752,N_3077,N_3592);
xnor U4753 (N_4753,N_3288,N_3592);
or U4754 (N_4754,N_3504,N_3014);
or U4755 (N_4755,N_3675,N_3663);
or U4756 (N_4756,N_3030,N_3358);
nand U4757 (N_4757,N_3217,N_3803);
or U4758 (N_4758,N_3615,N_3968);
and U4759 (N_4759,N_3372,N_3523);
nand U4760 (N_4760,N_3813,N_3617);
or U4761 (N_4761,N_3729,N_3693);
nand U4762 (N_4762,N_3192,N_3334);
nand U4763 (N_4763,N_3370,N_3401);
or U4764 (N_4764,N_3749,N_3965);
nor U4765 (N_4765,N_3353,N_3005);
and U4766 (N_4766,N_3187,N_3378);
xnor U4767 (N_4767,N_3103,N_3620);
nor U4768 (N_4768,N_3185,N_3094);
and U4769 (N_4769,N_3553,N_3450);
or U4770 (N_4770,N_3441,N_3389);
nand U4771 (N_4771,N_3692,N_3589);
nor U4772 (N_4772,N_3702,N_3469);
or U4773 (N_4773,N_3333,N_3251);
xnor U4774 (N_4774,N_3754,N_3083);
nand U4775 (N_4775,N_3142,N_3355);
and U4776 (N_4776,N_3429,N_3347);
xor U4777 (N_4777,N_3223,N_3825);
and U4778 (N_4778,N_3742,N_3593);
or U4779 (N_4779,N_3377,N_3365);
and U4780 (N_4780,N_3335,N_3540);
nor U4781 (N_4781,N_3076,N_3730);
nor U4782 (N_4782,N_3550,N_3299);
nand U4783 (N_4783,N_3398,N_3397);
nor U4784 (N_4784,N_3878,N_3990);
xor U4785 (N_4785,N_3596,N_3451);
and U4786 (N_4786,N_3318,N_3664);
nand U4787 (N_4787,N_3513,N_3096);
nor U4788 (N_4788,N_3369,N_3728);
or U4789 (N_4789,N_3055,N_3259);
nor U4790 (N_4790,N_3201,N_3227);
nand U4791 (N_4791,N_3572,N_3044);
and U4792 (N_4792,N_3240,N_3664);
or U4793 (N_4793,N_3463,N_3764);
and U4794 (N_4794,N_3524,N_3885);
nand U4795 (N_4795,N_3180,N_3698);
nor U4796 (N_4796,N_3574,N_3172);
and U4797 (N_4797,N_3264,N_3017);
and U4798 (N_4798,N_3915,N_3914);
nand U4799 (N_4799,N_3975,N_3640);
xor U4800 (N_4800,N_3902,N_3371);
xor U4801 (N_4801,N_3299,N_3665);
and U4802 (N_4802,N_3595,N_3878);
or U4803 (N_4803,N_3547,N_3270);
xnor U4804 (N_4804,N_3710,N_3701);
nand U4805 (N_4805,N_3583,N_3933);
nand U4806 (N_4806,N_3006,N_3791);
nand U4807 (N_4807,N_3105,N_3062);
or U4808 (N_4808,N_3460,N_3797);
nand U4809 (N_4809,N_3354,N_3397);
and U4810 (N_4810,N_3341,N_3246);
nor U4811 (N_4811,N_3671,N_3294);
and U4812 (N_4812,N_3823,N_3593);
and U4813 (N_4813,N_3119,N_3645);
or U4814 (N_4814,N_3188,N_3345);
and U4815 (N_4815,N_3066,N_3746);
or U4816 (N_4816,N_3580,N_3356);
nand U4817 (N_4817,N_3117,N_3679);
nand U4818 (N_4818,N_3504,N_3045);
and U4819 (N_4819,N_3619,N_3204);
or U4820 (N_4820,N_3462,N_3250);
and U4821 (N_4821,N_3216,N_3204);
and U4822 (N_4822,N_3087,N_3006);
xnor U4823 (N_4823,N_3833,N_3997);
nand U4824 (N_4824,N_3200,N_3871);
and U4825 (N_4825,N_3077,N_3456);
nand U4826 (N_4826,N_3756,N_3518);
nor U4827 (N_4827,N_3241,N_3146);
and U4828 (N_4828,N_3631,N_3731);
xnor U4829 (N_4829,N_3235,N_3979);
nand U4830 (N_4830,N_3181,N_3183);
nand U4831 (N_4831,N_3315,N_3874);
or U4832 (N_4832,N_3953,N_3209);
nand U4833 (N_4833,N_3317,N_3590);
and U4834 (N_4834,N_3803,N_3600);
nand U4835 (N_4835,N_3544,N_3724);
nor U4836 (N_4836,N_3626,N_3288);
nor U4837 (N_4837,N_3902,N_3150);
nand U4838 (N_4838,N_3212,N_3972);
xnor U4839 (N_4839,N_3894,N_3056);
nor U4840 (N_4840,N_3752,N_3249);
and U4841 (N_4841,N_3545,N_3493);
or U4842 (N_4842,N_3889,N_3350);
nand U4843 (N_4843,N_3882,N_3315);
nor U4844 (N_4844,N_3614,N_3318);
nor U4845 (N_4845,N_3485,N_3912);
xnor U4846 (N_4846,N_3965,N_3303);
or U4847 (N_4847,N_3578,N_3475);
xnor U4848 (N_4848,N_3527,N_3229);
nor U4849 (N_4849,N_3369,N_3989);
and U4850 (N_4850,N_3490,N_3685);
and U4851 (N_4851,N_3526,N_3776);
nand U4852 (N_4852,N_3996,N_3016);
nand U4853 (N_4853,N_3463,N_3672);
xor U4854 (N_4854,N_3670,N_3683);
nand U4855 (N_4855,N_3175,N_3685);
and U4856 (N_4856,N_3480,N_3881);
or U4857 (N_4857,N_3100,N_3722);
and U4858 (N_4858,N_3839,N_3235);
and U4859 (N_4859,N_3062,N_3243);
nor U4860 (N_4860,N_3461,N_3124);
nand U4861 (N_4861,N_3058,N_3834);
nand U4862 (N_4862,N_3221,N_3025);
or U4863 (N_4863,N_3120,N_3489);
and U4864 (N_4864,N_3974,N_3982);
nand U4865 (N_4865,N_3065,N_3693);
nand U4866 (N_4866,N_3348,N_3510);
and U4867 (N_4867,N_3553,N_3999);
nor U4868 (N_4868,N_3243,N_3509);
nor U4869 (N_4869,N_3845,N_3039);
and U4870 (N_4870,N_3083,N_3438);
nor U4871 (N_4871,N_3123,N_3459);
and U4872 (N_4872,N_3932,N_3336);
nor U4873 (N_4873,N_3211,N_3421);
nor U4874 (N_4874,N_3161,N_3651);
or U4875 (N_4875,N_3032,N_3888);
nor U4876 (N_4876,N_3724,N_3808);
or U4877 (N_4877,N_3538,N_3785);
nand U4878 (N_4878,N_3137,N_3006);
nor U4879 (N_4879,N_3873,N_3150);
nand U4880 (N_4880,N_3543,N_3853);
nand U4881 (N_4881,N_3497,N_3568);
and U4882 (N_4882,N_3276,N_3450);
nand U4883 (N_4883,N_3202,N_3049);
nand U4884 (N_4884,N_3476,N_3741);
nor U4885 (N_4885,N_3771,N_3297);
nor U4886 (N_4886,N_3160,N_3835);
or U4887 (N_4887,N_3505,N_3336);
nor U4888 (N_4888,N_3873,N_3663);
nand U4889 (N_4889,N_3878,N_3476);
or U4890 (N_4890,N_3914,N_3958);
xor U4891 (N_4891,N_3753,N_3949);
and U4892 (N_4892,N_3217,N_3543);
nor U4893 (N_4893,N_3412,N_3263);
and U4894 (N_4894,N_3720,N_3708);
and U4895 (N_4895,N_3931,N_3047);
or U4896 (N_4896,N_3360,N_3855);
xor U4897 (N_4897,N_3944,N_3303);
or U4898 (N_4898,N_3150,N_3448);
nor U4899 (N_4899,N_3449,N_3428);
or U4900 (N_4900,N_3610,N_3268);
or U4901 (N_4901,N_3689,N_3440);
nand U4902 (N_4902,N_3780,N_3776);
and U4903 (N_4903,N_3524,N_3928);
or U4904 (N_4904,N_3881,N_3671);
and U4905 (N_4905,N_3496,N_3098);
nor U4906 (N_4906,N_3110,N_3342);
and U4907 (N_4907,N_3883,N_3573);
or U4908 (N_4908,N_3050,N_3438);
and U4909 (N_4909,N_3750,N_3408);
xnor U4910 (N_4910,N_3729,N_3671);
nand U4911 (N_4911,N_3978,N_3340);
xnor U4912 (N_4912,N_3647,N_3757);
nand U4913 (N_4913,N_3436,N_3951);
or U4914 (N_4914,N_3768,N_3381);
and U4915 (N_4915,N_3244,N_3435);
and U4916 (N_4916,N_3409,N_3361);
nor U4917 (N_4917,N_3196,N_3195);
and U4918 (N_4918,N_3401,N_3130);
nand U4919 (N_4919,N_3999,N_3149);
or U4920 (N_4920,N_3547,N_3880);
nor U4921 (N_4921,N_3285,N_3182);
nor U4922 (N_4922,N_3250,N_3213);
nand U4923 (N_4923,N_3989,N_3256);
or U4924 (N_4924,N_3146,N_3525);
and U4925 (N_4925,N_3055,N_3934);
and U4926 (N_4926,N_3857,N_3364);
and U4927 (N_4927,N_3263,N_3130);
or U4928 (N_4928,N_3324,N_3674);
nand U4929 (N_4929,N_3046,N_3608);
nor U4930 (N_4930,N_3568,N_3379);
and U4931 (N_4931,N_3405,N_3566);
or U4932 (N_4932,N_3317,N_3509);
xnor U4933 (N_4933,N_3297,N_3089);
and U4934 (N_4934,N_3872,N_3317);
nor U4935 (N_4935,N_3461,N_3943);
nor U4936 (N_4936,N_3095,N_3915);
or U4937 (N_4937,N_3591,N_3238);
nand U4938 (N_4938,N_3219,N_3394);
and U4939 (N_4939,N_3684,N_3885);
or U4940 (N_4940,N_3082,N_3301);
nand U4941 (N_4941,N_3680,N_3985);
or U4942 (N_4942,N_3145,N_3012);
or U4943 (N_4943,N_3098,N_3520);
or U4944 (N_4944,N_3418,N_3814);
nand U4945 (N_4945,N_3001,N_3195);
or U4946 (N_4946,N_3334,N_3958);
nor U4947 (N_4947,N_3108,N_3728);
and U4948 (N_4948,N_3631,N_3011);
nand U4949 (N_4949,N_3615,N_3053);
nand U4950 (N_4950,N_3824,N_3778);
nor U4951 (N_4951,N_3003,N_3047);
nor U4952 (N_4952,N_3611,N_3581);
nand U4953 (N_4953,N_3272,N_3230);
and U4954 (N_4954,N_3886,N_3855);
nor U4955 (N_4955,N_3750,N_3077);
and U4956 (N_4956,N_3571,N_3418);
nor U4957 (N_4957,N_3454,N_3014);
and U4958 (N_4958,N_3895,N_3254);
nor U4959 (N_4959,N_3309,N_3407);
nand U4960 (N_4960,N_3223,N_3540);
or U4961 (N_4961,N_3983,N_3321);
nand U4962 (N_4962,N_3524,N_3404);
nor U4963 (N_4963,N_3027,N_3903);
nand U4964 (N_4964,N_3719,N_3648);
and U4965 (N_4965,N_3597,N_3979);
or U4966 (N_4966,N_3005,N_3624);
or U4967 (N_4967,N_3160,N_3824);
nor U4968 (N_4968,N_3511,N_3526);
nor U4969 (N_4969,N_3707,N_3058);
xor U4970 (N_4970,N_3439,N_3275);
nand U4971 (N_4971,N_3666,N_3516);
and U4972 (N_4972,N_3630,N_3971);
xnor U4973 (N_4973,N_3109,N_3455);
nor U4974 (N_4974,N_3038,N_3224);
or U4975 (N_4975,N_3196,N_3762);
nor U4976 (N_4976,N_3430,N_3222);
nand U4977 (N_4977,N_3054,N_3550);
or U4978 (N_4978,N_3630,N_3868);
and U4979 (N_4979,N_3136,N_3286);
xor U4980 (N_4980,N_3096,N_3132);
or U4981 (N_4981,N_3502,N_3537);
or U4982 (N_4982,N_3670,N_3473);
xor U4983 (N_4983,N_3227,N_3923);
and U4984 (N_4984,N_3673,N_3705);
nand U4985 (N_4985,N_3742,N_3201);
nor U4986 (N_4986,N_3357,N_3687);
or U4987 (N_4987,N_3729,N_3400);
or U4988 (N_4988,N_3793,N_3583);
nor U4989 (N_4989,N_3671,N_3847);
or U4990 (N_4990,N_3889,N_3568);
nand U4991 (N_4991,N_3016,N_3728);
or U4992 (N_4992,N_3253,N_3824);
xor U4993 (N_4993,N_3450,N_3934);
nand U4994 (N_4994,N_3110,N_3545);
and U4995 (N_4995,N_3381,N_3792);
nor U4996 (N_4996,N_3604,N_3494);
nand U4997 (N_4997,N_3780,N_3241);
or U4998 (N_4998,N_3778,N_3961);
or U4999 (N_4999,N_3532,N_3844);
and UO_0 (O_0,N_4515,N_4289);
and UO_1 (O_1,N_4909,N_4264);
xnor UO_2 (O_2,N_4036,N_4583);
and UO_3 (O_3,N_4979,N_4592);
and UO_4 (O_4,N_4285,N_4665);
or UO_5 (O_5,N_4989,N_4458);
or UO_6 (O_6,N_4559,N_4579);
and UO_7 (O_7,N_4806,N_4826);
and UO_8 (O_8,N_4914,N_4873);
nand UO_9 (O_9,N_4915,N_4197);
xor UO_10 (O_10,N_4783,N_4890);
or UO_11 (O_11,N_4723,N_4581);
xor UO_12 (O_12,N_4258,N_4772);
xor UO_13 (O_13,N_4596,N_4904);
nor UO_14 (O_14,N_4899,N_4934);
or UO_15 (O_15,N_4192,N_4278);
nand UO_16 (O_16,N_4548,N_4002);
or UO_17 (O_17,N_4427,N_4520);
nand UO_18 (O_18,N_4576,N_4460);
and UO_19 (O_19,N_4673,N_4729);
nand UO_20 (O_20,N_4813,N_4923);
nand UO_21 (O_21,N_4293,N_4660);
nor UO_22 (O_22,N_4620,N_4687);
or UO_23 (O_23,N_4283,N_4085);
xnor UO_24 (O_24,N_4249,N_4616);
xor UO_25 (O_25,N_4432,N_4602);
nor UO_26 (O_26,N_4091,N_4875);
xor UO_27 (O_27,N_4137,N_4752);
nor UO_28 (O_28,N_4812,N_4131);
xor UO_29 (O_29,N_4396,N_4566);
nor UO_30 (O_30,N_4822,N_4093);
xnor UO_31 (O_31,N_4896,N_4506);
or UO_32 (O_32,N_4181,N_4006);
and UO_33 (O_33,N_4417,N_4907);
nor UO_34 (O_34,N_4829,N_4717);
nand UO_35 (O_35,N_4646,N_4633);
nor UO_36 (O_36,N_4449,N_4951);
nand UO_37 (O_37,N_4864,N_4448);
nand UO_38 (O_38,N_4148,N_4632);
nand UO_39 (O_39,N_4836,N_4854);
and UO_40 (O_40,N_4861,N_4840);
nor UO_41 (O_41,N_4901,N_4946);
and UO_42 (O_42,N_4428,N_4378);
and UO_43 (O_43,N_4865,N_4852);
nand UO_44 (O_44,N_4132,N_4047);
nor UO_45 (O_45,N_4252,N_4498);
nand UO_46 (O_46,N_4344,N_4851);
or UO_47 (O_47,N_4297,N_4495);
nand UO_48 (O_48,N_4759,N_4100);
nand UO_49 (O_49,N_4941,N_4038);
nand UO_50 (O_50,N_4897,N_4929);
nor UO_51 (O_51,N_4442,N_4578);
or UO_52 (O_52,N_4163,N_4908);
or UO_53 (O_53,N_4310,N_4189);
nor UO_54 (O_54,N_4666,N_4327);
and UO_55 (O_55,N_4743,N_4236);
nor UO_56 (O_56,N_4201,N_4162);
or UO_57 (O_57,N_4701,N_4275);
nor UO_58 (O_58,N_4230,N_4168);
nor UO_59 (O_59,N_4755,N_4705);
nand UO_60 (O_60,N_4465,N_4124);
nor UO_61 (O_61,N_4221,N_4538);
nand UO_62 (O_62,N_4497,N_4404);
or UO_63 (O_63,N_4255,N_4203);
and UO_64 (O_64,N_4485,N_4195);
or UO_65 (O_65,N_4571,N_4756);
and UO_66 (O_66,N_4963,N_4645);
or UO_67 (O_67,N_4005,N_4069);
or UO_68 (O_68,N_4032,N_4695);
nand UO_69 (O_69,N_4993,N_4563);
nor UO_70 (O_70,N_4552,N_4707);
or UO_71 (O_71,N_4325,N_4688);
and UO_72 (O_72,N_4841,N_4985);
or UO_73 (O_73,N_4781,N_4346);
xor UO_74 (O_74,N_4526,N_4975);
or UO_75 (O_75,N_4459,N_4685);
or UO_76 (O_76,N_4519,N_4077);
or UO_77 (O_77,N_4614,N_4503);
or UO_78 (O_78,N_4347,N_4228);
nand UO_79 (O_79,N_4220,N_4775);
xor UO_80 (O_80,N_4965,N_4869);
nor UO_81 (O_81,N_4144,N_4142);
nand UO_82 (O_82,N_4892,N_4451);
or UO_83 (O_83,N_4016,N_4691);
or UO_84 (O_84,N_4700,N_4453);
xor UO_85 (O_85,N_4407,N_4948);
xnor UO_86 (O_86,N_4569,N_4523);
and UO_87 (O_87,N_4670,N_4867);
and UO_88 (O_88,N_4151,N_4245);
nand UO_89 (O_89,N_4480,N_4001);
or UO_90 (O_90,N_4223,N_4913);
and UO_91 (O_91,N_4547,N_4354);
nor UO_92 (O_92,N_4956,N_4356);
and UO_93 (O_93,N_4970,N_4490);
and UO_94 (O_94,N_4359,N_4092);
or UO_95 (O_95,N_4712,N_4771);
and UO_96 (O_96,N_4390,N_4521);
or UO_97 (O_97,N_4704,N_4291);
nand UO_98 (O_98,N_4227,N_4214);
nand UO_99 (O_99,N_4585,N_4218);
xnor UO_100 (O_100,N_4528,N_4368);
nor UO_101 (O_101,N_4727,N_4703);
and UO_102 (O_102,N_4338,N_4678);
nor UO_103 (O_103,N_4820,N_4351);
or UO_104 (O_104,N_4881,N_4080);
or UO_105 (O_105,N_4053,N_4997);
or UO_106 (O_106,N_4770,N_4933);
and UO_107 (O_107,N_4565,N_4430);
nor UO_108 (O_108,N_4676,N_4593);
xnor UO_109 (O_109,N_4714,N_4696);
nor UO_110 (O_110,N_4198,N_4161);
nand UO_111 (O_111,N_4641,N_4996);
xor UO_112 (O_112,N_4724,N_4054);
nand UO_113 (O_113,N_4482,N_4194);
nor UO_114 (O_114,N_4165,N_4467);
nand UO_115 (O_115,N_4323,N_4478);
nor UO_116 (O_116,N_4370,N_4824);
nor UO_117 (O_117,N_4030,N_4324);
nor UO_118 (O_118,N_4473,N_4987);
or UO_119 (O_119,N_4635,N_4487);
nor UO_120 (O_120,N_4363,N_4130);
nor UO_121 (O_121,N_4835,N_4008);
nand UO_122 (O_122,N_4493,N_4375);
nor UO_123 (O_123,N_4232,N_4023);
nor UO_124 (O_124,N_4697,N_4604);
nand UO_125 (O_125,N_4543,N_4170);
or UO_126 (O_126,N_4537,N_4573);
or UO_127 (O_127,N_4029,N_4922);
nor UO_128 (O_128,N_4044,N_4575);
and UO_129 (O_129,N_4436,N_4075);
nor UO_130 (O_130,N_4332,N_4631);
and UO_131 (O_131,N_4803,N_4988);
and UO_132 (O_132,N_4150,N_4022);
or UO_133 (O_133,N_4481,N_4174);
nand UO_134 (O_134,N_4784,N_4178);
nor UO_135 (O_135,N_4489,N_4135);
or UO_136 (O_136,N_4244,N_4730);
nand UO_137 (O_137,N_4968,N_4937);
nor UO_138 (O_138,N_4950,N_4874);
nand UO_139 (O_139,N_4582,N_4385);
xor UO_140 (O_140,N_4190,N_4990);
and UO_141 (O_141,N_4260,N_4280);
nand UO_142 (O_142,N_4684,N_4878);
or UO_143 (O_143,N_4516,N_4844);
and UO_144 (O_144,N_4982,N_4147);
nor UO_145 (O_145,N_4715,N_4474);
nand UO_146 (O_146,N_4850,N_4445);
xnor UO_147 (O_147,N_4401,N_4921);
or UO_148 (O_148,N_4207,N_4634);
nand UO_149 (O_149,N_4317,N_4898);
or UO_150 (O_150,N_4064,N_4452);
nor UO_151 (O_151,N_4846,N_4321);
and UO_152 (O_152,N_4042,N_4708);
nand UO_153 (O_153,N_4960,N_4469);
nor UO_154 (O_154,N_4247,N_4740);
nor UO_155 (O_155,N_4202,N_4827);
and UO_156 (O_156,N_4027,N_4362);
nor UO_157 (O_157,N_4377,N_4007);
or UO_158 (O_158,N_4647,N_4330);
nand UO_159 (O_159,N_4930,N_4859);
or UO_160 (O_160,N_4750,N_4216);
and UO_161 (O_161,N_4379,N_4919);
nor UO_162 (O_162,N_4425,N_4554);
or UO_163 (O_163,N_4862,N_4113);
nor UO_164 (O_164,N_4268,N_4828);
or UO_165 (O_165,N_4648,N_4574);
nand UO_166 (O_166,N_4818,N_4830);
xnor UO_167 (O_167,N_4590,N_4461);
nor UO_168 (O_168,N_4789,N_4629);
nor UO_169 (O_169,N_4991,N_4735);
and UO_170 (O_170,N_4880,N_4342);
nand UO_171 (O_171,N_4804,N_4464);
nand UO_172 (O_172,N_4035,N_4857);
and UO_173 (O_173,N_4761,N_4518);
nand UO_174 (O_174,N_4529,N_4782);
nand UO_175 (O_175,N_4295,N_4087);
xnor UO_176 (O_176,N_4580,N_4381);
and UO_177 (O_177,N_4718,N_4595);
nor UO_178 (O_178,N_4186,N_4954);
nand UO_179 (O_179,N_4553,N_4253);
nor UO_180 (O_180,N_4267,N_4671);
nor UO_181 (O_181,N_4541,N_4125);
and UO_182 (O_182,N_4738,N_4636);
nand UO_183 (O_183,N_4959,N_4057);
nor UO_184 (O_184,N_4380,N_4655);
or UO_185 (O_185,N_4078,N_4303);
or UO_186 (O_186,N_4305,N_4143);
nand UO_187 (O_187,N_4663,N_4773);
or UO_188 (O_188,N_4924,N_4763);
or UO_189 (O_189,N_4733,N_4664);
and UO_190 (O_190,N_4817,N_4618);
or UO_191 (O_191,N_4906,N_4339);
nor UO_192 (O_192,N_4004,N_4463);
and UO_193 (O_193,N_4051,N_4809);
nor UO_194 (O_194,N_4288,N_4188);
nor UO_195 (O_195,N_4502,N_4431);
or UO_196 (O_196,N_4702,N_4233);
nand UO_197 (O_197,N_4043,N_4849);
xnor UO_198 (O_198,N_4683,N_4643);
or UO_199 (O_199,N_4301,N_4208);
and UO_200 (O_200,N_4433,N_4597);
nand UO_201 (O_201,N_4807,N_4550);
or UO_202 (O_202,N_4888,N_4098);
nand UO_203 (O_203,N_4509,N_4248);
or UO_204 (O_204,N_4511,N_4096);
or UO_205 (O_205,N_4067,N_4600);
and UO_206 (O_206,N_4883,N_4911);
and UO_207 (O_207,N_4184,N_4879);
or UO_208 (O_208,N_4587,N_4172);
nand UO_209 (O_209,N_4331,N_4068);
nand UO_210 (O_210,N_4259,N_4101);
and UO_211 (O_211,N_4626,N_4483);
nand UO_212 (O_212,N_4367,N_4760);
xnor UO_213 (O_213,N_4508,N_4079);
and UO_214 (O_214,N_4577,N_4199);
and UO_215 (O_215,N_4556,N_4313);
nor UO_216 (O_216,N_4048,N_4839);
or UO_217 (O_217,N_4564,N_4667);
and UO_218 (O_218,N_4711,N_4816);
nand UO_219 (O_219,N_4065,N_4668);
nor UO_220 (O_220,N_4871,N_4681);
or UO_221 (O_221,N_4504,N_4779);
nor UO_222 (O_222,N_4468,N_4443);
and UO_223 (O_223,N_4139,N_4166);
xor UO_224 (O_224,N_4658,N_4061);
xnor UO_225 (O_225,N_4742,N_4319);
or UO_226 (O_226,N_4238,N_4967);
nand UO_227 (O_227,N_4369,N_4217);
and UO_228 (O_228,N_4121,N_4239);
and UO_229 (O_229,N_4376,N_4964);
or UO_230 (O_230,N_4066,N_4833);
or UO_231 (O_231,N_4336,N_4706);
or UO_232 (O_232,N_4505,N_4444);
nor UO_233 (O_233,N_4082,N_4603);
nand UO_234 (O_234,N_4307,N_4099);
xnor UO_235 (O_235,N_4383,N_4973);
nand UO_236 (O_236,N_4625,N_4877);
nor UO_237 (O_237,N_4455,N_4250);
and UO_238 (O_238,N_4847,N_4105);
nor UO_239 (O_239,N_4624,N_4978);
nor UO_240 (O_240,N_4391,N_4020);
nand UO_241 (O_241,N_4284,N_4457);
nand UO_242 (O_242,N_4389,N_4731);
nor UO_243 (O_243,N_4254,N_4741);
nand UO_244 (O_244,N_4224,N_4746);
and UO_245 (O_245,N_4825,N_4477);
nor UO_246 (O_246,N_4406,N_4212);
xor UO_247 (O_247,N_4891,N_4119);
nor UO_248 (O_248,N_4039,N_4501);
nand UO_249 (O_249,N_4397,N_4299);
xnor UO_250 (O_250,N_4675,N_4175);
or UO_251 (O_251,N_4357,N_4757);
nand UO_252 (O_252,N_4196,N_4074);
and UO_253 (O_253,N_4751,N_4187);
nor UO_254 (O_254,N_4126,N_4155);
or UO_255 (O_255,N_4104,N_4011);
or UO_256 (O_256,N_4415,N_4241);
or UO_257 (O_257,N_4765,N_4766);
xor UO_258 (O_258,N_4611,N_4103);
xnor UO_259 (O_259,N_4120,N_4679);
or UO_260 (O_260,N_4438,N_4606);
nand UO_261 (O_261,N_4315,N_4318);
or UO_262 (O_262,N_4387,N_4598);
nor UO_263 (O_263,N_4720,N_4621);
or UO_264 (O_264,N_4412,N_4279);
nand UO_265 (O_265,N_4586,N_4140);
and UO_266 (O_266,N_4429,N_4984);
nor UO_267 (O_267,N_4364,N_4456);
nor UO_268 (O_268,N_4605,N_4003);
and UO_269 (O_269,N_4447,N_4185);
nand UO_270 (O_270,N_4999,N_4118);
nand UO_271 (O_271,N_4215,N_4992);
or UO_272 (O_272,N_4010,N_4535);
xor UO_273 (O_273,N_4926,N_4333);
or UO_274 (O_274,N_4837,N_4622);
and UO_275 (O_275,N_4176,N_4395);
nor UO_276 (O_276,N_4117,N_4494);
nor UO_277 (O_277,N_4311,N_4567);
nand UO_278 (O_278,N_4209,N_4296);
and UO_279 (O_279,N_4152,N_4242);
nand UO_280 (O_280,N_4393,N_4127);
nor UO_281 (O_281,N_4097,N_4371);
or UO_282 (O_282,N_4774,N_4435);
xnor UO_283 (O_283,N_4328,N_4693);
nor UO_284 (O_284,N_4164,N_4949);
and UO_285 (O_285,N_4845,N_4419);
nor UO_286 (O_286,N_4955,N_4619);
or UO_287 (O_287,N_4698,N_4000);
or UO_288 (O_288,N_4158,N_4848);
nand UO_289 (O_289,N_4767,N_4562);
nand UO_290 (O_290,N_4601,N_4866);
and UO_291 (O_291,N_4843,N_4938);
xnor UO_292 (O_292,N_4800,N_4659);
nor UO_293 (O_293,N_4145,N_4046);
or UO_294 (O_294,N_4546,N_4037);
nor UO_295 (O_295,N_4111,N_4709);
nor UO_296 (O_296,N_4424,N_4470);
nor UO_297 (O_297,N_4925,N_4024);
nand UO_298 (O_298,N_4373,N_4366);
nor UO_299 (O_299,N_4094,N_4200);
xnor UO_300 (O_300,N_4270,N_4246);
nor UO_301 (O_301,N_4532,N_4302);
nor UO_302 (O_302,N_4551,N_4345);
xnor UO_303 (O_303,N_4682,N_4348);
nand UO_304 (O_304,N_4083,N_4617);
or UO_305 (O_305,N_4530,N_4527);
and UO_306 (O_306,N_4222,N_4609);
nor UO_307 (O_307,N_4167,N_4479);
nand UO_308 (O_308,N_4900,N_4271);
and UO_309 (O_309,N_4644,N_4748);
or UO_310 (O_310,N_4298,N_4725);
xnor UO_311 (O_311,N_4734,N_4441);
and UO_312 (O_312,N_4694,N_4669);
nand UO_313 (O_313,N_4420,N_4737);
and UO_314 (O_314,N_4749,N_4257);
xor UO_315 (O_315,N_4536,N_4049);
xnor UO_316 (O_316,N_4952,N_4801);
or UO_317 (O_317,N_4677,N_4388);
nand UO_318 (O_318,N_4823,N_4808);
nand UO_319 (O_319,N_4939,N_4014);
and UO_320 (O_320,N_4886,N_4889);
nor UO_321 (O_321,N_4572,N_4713);
nor UO_322 (O_322,N_4514,N_4558);
nand UO_323 (O_323,N_4986,N_4838);
nand UO_324 (O_324,N_4399,N_4692);
xor UO_325 (O_325,N_4744,N_4110);
nand UO_326 (O_326,N_4017,N_4510);
nor UO_327 (O_327,N_4607,N_4337);
or UO_328 (O_328,N_4762,N_4095);
or UO_329 (O_329,N_4674,N_4796);
or UO_330 (O_330,N_4365,N_4545);
xnor UO_331 (O_331,N_4034,N_4060);
or UO_332 (O_332,N_4795,N_4785);
nand UO_333 (O_333,N_4995,N_4885);
and UO_334 (O_334,N_4534,N_4780);
or UO_335 (O_335,N_4306,N_4699);
and UO_336 (O_336,N_4753,N_4764);
or UO_337 (O_337,N_4902,N_4832);
or UO_338 (O_338,N_4680,N_4831);
nor UO_339 (O_339,N_4472,N_4262);
nor UO_340 (O_340,N_4814,N_4608);
and UO_341 (O_341,N_4736,N_4895);
nand UO_342 (O_342,N_4903,N_4437);
nor UO_343 (O_343,N_4758,N_4936);
nor UO_344 (O_344,N_4326,N_4943);
nand UO_345 (O_345,N_4411,N_4540);
nor UO_346 (O_346,N_4918,N_4081);
and UO_347 (O_347,N_4128,N_4860);
and UO_348 (O_348,N_4791,N_4112);
nor UO_349 (O_349,N_4966,N_4916);
xnor UO_350 (O_350,N_4821,N_4355);
and UO_351 (O_351,N_4544,N_4205);
and UO_352 (O_352,N_4555,N_4882);
nand UO_353 (O_353,N_4454,N_4204);
nand UO_354 (O_354,N_4623,N_4334);
nand UO_355 (O_355,N_4234,N_4811);
and UO_356 (O_356,N_4870,N_4893);
nor UO_357 (O_357,N_4106,N_4776);
nor UO_358 (O_358,N_4123,N_4792);
and UO_359 (O_359,N_4513,N_4146);
xnor UO_360 (O_360,N_4969,N_4266);
and UO_361 (O_361,N_4059,N_4466);
or UO_362 (O_362,N_4721,N_4940);
nand UO_363 (O_363,N_4414,N_4193);
xnor UO_364 (O_364,N_4805,N_4863);
and UO_365 (O_365,N_4980,N_4052);
nand UO_366 (O_366,N_4072,N_4686);
or UO_367 (O_367,N_4599,N_4887);
and UO_368 (O_368,N_4810,N_4710);
nand UO_369 (O_369,N_4076,N_4570);
xor UO_370 (O_370,N_4722,N_4656);
xor UO_371 (O_371,N_4308,N_4329);
and UO_372 (O_372,N_4423,N_4793);
nor UO_373 (O_373,N_4942,N_4109);
xor UO_374 (O_374,N_4589,N_4434);
and UO_375 (O_375,N_4522,N_4213);
nor UO_376 (O_376,N_4386,N_4211);
nor UO_377 (O_377,N_4272,N_4834);
nand UO_378 (O_378,N_4855,N_4361);
nand UO_379 (O_379,N_4191,N_4349);
nand UO_380 (O_380,N_4690,N_4657);
and UO_381 (O_381,N_4019,N_4876);
and UO_382 (O_382,N_4013,N_4798);
and UO_383 (O_383,N_4180,N_4134);
nor UO_384 (O_384,N_4265,N_4507);
and UO_385 (O_385,N_4612,N_4856);
and UO_386 (O_386,N_4281,N_4591);
nor UO_387 (O_387,N_4372,N_4160);
nor UO_388 (O_388,N_4471,N_4440);
or UO_389 (O_389,N_4041,N_4932);
or UO_390 (O_390,N_4561,N_4450);
nand UO_391 (O_391,N_4944,N_4070);
nand UO_392 (O_392,N_4309,N_4484);
and UO_393 (O_393,N_4031,N_4133);
xor UO_394 (O_394,N_4630,N_4225);
nor UO_395 (O_395,N_4088,N_4475);
nor UO_396 (O_396,N_4304,N_4797);
nor UO_397 (O_397,N_4157,N_4947);
nor UO_398 (O_398,N_4116,N_4169);
or UO_399 (O_399,N_4953,N_4421);
nor UO_400 (O_400,N_4998,N_4894);
nand UO_401 (O_401,N_4108,N_4728);
xnor UO_402 (O_402,N_4353,N_4560);
nand UO_403 (O_403,N_4292,N_4261);
or UO_404 (O_404,N_4533,N_4251);
or UO_405 (O_405,N_4769,N_4154);
xor UO_406 (O_406,N_4492,N_4910);
nor UO_407 (O_407,N_4787,N_4408);
and UO_408 (O_408,N_4739,N_4413);
or UO_409 (O_409,N_4409,N_4322);
and UO_410 (O_410,N_4269,N_4488);
xor UO_411 (O_411,N_4149,N_4716);
xor UO_412 (O_412,N_4256,N_4958);
or UO_413 (O_413,N_4115,N_4063);
nor UO_414 (O_414,N_4439,N_4935);
nand UO_415 (O_415,N_4173,N_4177);
and UO_416 (O_416,N_4084,N_4962);
or UO_417 (O_417,N_4229,N_4786);
nand UO_418 (O_418,N_4777,N_4122);
and UO_419 (O_419,N_4352,N_4028);
or UO_420 (O_420,N_4405,N_4071);
and UO_421 (O_421,N_4138,N_4476);
and UO_422 (O_422,N_4983,N_4025);
xnor UO_423 (O_423,N_4961,N_4183);
or UO_424 (O_424,N_4652,N_4920);
and UO_425 (O_425,N_4613,N_4141);
xnor UO_426 (O_426,N_4219,N_4491);
or UO_427 (O_427,N_4858,N_4819);
nand UO_428 (O_428,N_4931,N_4206);
or UO_429 (O_429,N_4089,N_4237);
or UO_430 (O_430,N_4917,N_4642);
or UO_431 (O_431,N_4594,N_4568);
and UO_432 (O_432,N_4517,N_4410);
or UO_433 (O_433,N_4927,N_4732);
and UO_434 (O_434,N_4290,N_4073);
or UO_435 (O_435,N_4358,N_4335);
nand UO_436 (O_436,N_4977,N_4026);
nor UO_437 (O_437,N_4050,N_4426);
nor UO_438 (O_438,N_4058,N_4628);
and UO_439 (O_439,N_4945,N_4277);
nand UO_440 (O_440,N_4957,N_4136);
nor UO_441 (O_441,N_4588,N_4392);
and UO_442 (O_442,N_4790,N_4446);
nor UO_443 (O_443,N_4976,N_4639);
xor UO_444 (O_444,N_4649,N_4525);
xnor UO_445 (O_445,N_4654,N_4056);
nor UO_446 (O_446,N_4745,N_4418);
nor UO_447 (O_447,N_4314,N_4974);
nand UO_448 (O_448,N_4549,N_4129);
nand UO_449 (O_449,N_4416,N_4778);
or UO_450 (O_450,N_4815,N_4182);
or UO_451 (O_451,N_4341,N_4403);
or UO_452 (O_452,N_4086,N_4788);
nand UO_453 (O_453,N_4928,N_4971);
xor UO_454 (O_454,N_4640,N_4539);
or UO_455 (O_455,N_4055,N_4496);
or UO_456 (O_456,N_4524,N_4316);
nor UO_457 (O_457,N_4672,N_4726);
nor UO_458 (O_458,N_4114,N_4794);
nand UO_459 (O_459,N_4210,N_4320);
xnor UO_460 (O_460,N_4240,N_4462);
nor UO_461 (O_461,N_4040,N_4273);
nor UO_462 (O_462,N_4802,N_4153);
and UO_463 (O_463,N_4653,N_4179);
and UO_464 (O_464,N_4062,N_4662);
nor UO_465 (O_465,N_4235,N_4276);
nor UO_466 (O_466,N_4768,N_4799);
nor UO_467 (O_467,N_4542,N_4719);
nand UO_468 (O_468,N_4350,N_4499);
nand UO_469 (O_469,N_4243,N_4531);
or UO_470 (O_470,N_4102,N_4374);
nand UO_471 (O_471,N_4384,N_4584);
nand UO_472 (O_472,N_4312,N_4650);
nor UO_473 (O_473,N_4382,N_4012);
or UO_474 (O_474,N_4274,N_4360);
nand UO_475 (O_475,N_4045,N_4912);
or UO_476 (O_476,N_4300,N_4263);
nand UO_477 (O_477,N_4842,N_4868);
xnor UO_478 (O_478,N_4486,N_4905);
nand UO_479 (O_479,N_4398,N_4033);
nand UO_480 (O_480,N_4422,N_4400);
and UO_481 (O_481,N_4689,N_4394);
xor UO_482 (O_482,N_4021,N_4171);
nand UO_483 (O_483,N_4340,N_4615);
and UO_484 (O_484,N_4981,N_4015);
or UO_485 (O_485,N_4754,N_4286);
and UO_486 (O_486,N_4231,N_4972);
and UO_487 (O_487,N_4637,N_4638);
nand UO_488 (O_488,N_4107,N_4610);
nor UO_489 (O_489,N_4557,N_4402);
or UO_490 (O_490,N_4159,N_4294);
nor UO_491 (O_491,N_4872,N_4627);
and UO_492 (O_492,N_4156,N_4500);
and UO_493 (O_493,N_4090,N_4512);
nand UO_494 (O_494,N_4009,N_4661);
nor UO_495 (O_495,N_4853,N_4994);
xor UO_496 (O_496,N_4282,N_4226);
nand UO_497 (O_497,N_4343,N_4747);
xor UO_498 (O_498,N_4287,N_4018);
or UO_499 (O_499,N_4884,N_4651);
and UO_500 (O_500,N_4294,N_4778);
and UO_501 (O_501,N_4690,N_4215);
and UO_502 (O_502,N_4321,N_4490);
or UO_503 (O_503,N_4601,N_4315);
or UO_504 (O_504,N_4711,N_4059);
or UO_505 (O_505,N_4612,N_4419);
nor UO_506 (O_506,N_4518,N_4292);
nor UO_507 (O_507,N_4211,N_4653);
nand UO_508 (O_508,N_4221,N_4896);
nand UO_509 (O_509,N_4370,N_4700);
nand UO_510 (O_510,N_4609,N_4361);
nor UO_511 (O_511,N_4291,N_4934);
nor UO_512 (O_512,N_4035,N_4696);
and UO_513 (O_513,N_4925,N_4415);
and UO_514 (O_514,N_4324,N_4727);
nor UO_515 (O_515,N_4596,N_4309);
and UO_516 (O_516,N_4015,N_4765);
nand UO_517 (O_517,N_4049,N_4581);
nor UO_518 (O_518,N_4427,N_4765);
nor UO_519 (O_519,N_4298,N_4928);
xnor UO_520 (O_520,N_4019,N_4041);
nand UO_521 (O_521,N_4246,N_4505);
or UO_522 (O_522,N_4770,N_4684);
nand UO_523 (O_523,N_4249,N_4830);
and UO_524 (O_524,N_4700,N_4053);
and UO_525 (O_525,N_4979,N_4434);
and UO_526 (O_526,N_4630,N_4030);
nor UO_527 (O_527,N_4773,N_4280);
xnor UO_528 (O_528,N_4763,N_4486);
nand UO_529 (O_529,N_4503,N_4896);
or UO_530 (O_530,N_4916,N_4674);
and UO_531 (O_531,N_4482,N_4449);
xor UO_532 (O_532,N_4441,N_4985);
and UO_533 (O_533,N_4849,N_4998);
or UO_534 (O_534,N_4025,N_4853);
and UO_535 (O_535,N_4960,N_4360);
and UO_536 (O_536,N_4255,N_4855);
nor UO_537 (O_537,N_4021,N_4945);
or UO_538 (O_538,N_4822,N_4179);
and UO_539 (O_539,N_4572,N_4305);
or UO_540 (O_540,N_4567,N_4401);
xnor UO_541 (O_541,N_4438,N_4963);
nor UO_542 (O_542,N_4198,N_4961);
nor UO_543 (O_543,N_4807,N_4045);
xor UO_544 (O_544,N_4577,N_4660);
or UO_545 (O_545,N_4750,N_4301);
nor UO_546 (O_546,N_4646,N_4059);
nand UO_547 (O_547,N_4755,N_4012);
nand UO_548 (O_548,N_4353,N_4015);
and UO_549 (O_549,N_4241,N_4880);
or UO_550 (O_550,N_4510,N_4365);
nor UO_551 (O_551,N_4086,N_4413);
and UO_552 (O_552,N_4734,N_4670);
nor UO_553 (O_553,N_4997,N_4354);
xnor UO_554 (O_554,N_4292,N_4870);
nor UO_555 (O_555,N_4427,N_4826);
nor UO_556 (O_556,N_4186,N_4162);
nand UO_557 (O_557,N_4064,N_4275);
nand UO_558 (O_558,N_4313,N_4178);
nor UO_559 (O_559,N_4920,N_4357);
and UO_560 (O_560,N_4594,N_4004);
nor UO_561 (O_561,N_4501,N_4824);
or UO_562 (O_562,N_4636,N_4556);
xor UO_563 (O_563,N_4638,N_4196);
or UO_564 (O_564,N_4925,N_4233);
nand UO_565 (O_565,N_4047,N_4845);
xor UO_566 (O_566,N_4556,N_4517);
nand UO_567 (O_567,N_4646,N_4576);
xnor UO_568 (O_568,N_4520,N_4297);
nor UO_569 (O_569,N_4009,N_4298);
or UO_570 (O_570,N_4995,N_4936);
and UO_571 (O_571,N_4486,N_4411);
xor UO_572 (O_572,N_4937,N_4691);
nand UO_573 (O_573,N_4661,N_4669);
nor UO_574 (O_574,N_4703,N_4527);
nand UO_575 (O_575,N_4534,N_4367);
xor UO_576 (O_576,N_4936,N_4026);
and UO_577 (O_577,N_4637,N_4221);
nor UO_578 (O_578,N_4424,N_4116);
or UO_579 (O_579,N_4501,N_4448);
or UO_580 (O_580,N_4048,N_4357);
xnor UO_581 (O_581,N_4189,N_4836);
or UO_582 (O_582,N_4948,N_4048);
nand UO_583 (O_583,N_4161,N_4117);
xor UO_584 (O_584,N_4045,N_4939);
xor UO_585 (O_585,N_4299,N_4754);
nor UO_586 (O_586,N_4685,N_4675);
xnor UO_587 (O_587,N_4878,N_4569);
nor UO_588 (O_588,N_4023,N_4104);
nand UO_589 (O_589,N_4487,N_4007);
and UO_590 (O_590,N_4381,N_4795);
nand UO_591 (O_591,N_4108,N_4085);
nand UO_592 (O_592,N_4089,N_4121);
and UO_593 (O_593,N_4950,N_4247);
nor UO_594 (O_594,N_4016,N_4581);
nand UO_595 (O_595,N_4806,N_4831);
nor UO_596 (O_596,N_4145,N_4002);
or UO_597 (O_597,N_4281,N_4924);
and UO_598 (O_598,N_4677,N_4206);
nand UO_599 (O_599,N_4576,N_4891);
xor UO_600 (O_600,N_4389,N_4152);
nand UO_601 (O_601,N_4319,N_4250);
or UO_602 (O_602,N_4885,N_4111);
nor UO_603 (O_603,N_4226,N_4264);
nor UO_604 (O_604,N_4546,N_4665);
or UO_605 (O_605,N_4216,N_4556);
and UO_606 (O_606,N_4175,N_4265);
nor UO_607 (O_607,N_4495,N_4756);
or UO_608 (O_608,N_4862,N_4309);
or UO_609 (O_609,N_4104,N_4421);
and UO_610 (O_610,N_4331,N_4785);
xor UO_611 (O_611,N_4787,N_4521);
nand UO_612 (O_612,N_4795,N_4431);
xor UO_613 (O_613,N_4256,N_4576);
xor UO_614 (O_614,N_4238,N_4538);
nand UO_615 (O_615,N_4788,N_4363);
xor UO_616 (O_616,N_4356,N_4338);
and UO_617 (O_617,N_4718,N_4604);
nand UO_618 (O_618,N_4419,N_4069);
and UO_619 (O_619,N_4561,N_4992);
and UO_620 (O_620,N_4497,N_4284);
or UO_621 (O_621,N_4087,N_4548);
or UO_622 (O_622,N_4970,N_4752);
and UO_623 (O_623,N_4811,N_4024);
nor UO_624 (O_624,N_4999,N_4892);
xor UO_625 (O_625,N_4166,N_4730);
and UO_626 (O_626,N_4742,N_4151);
nor UO_627 (O_627,N_4735,N_4080);
xor UO_628 (O_628,N_4456,N_4996);
nand UO_629 (O_629,N_4164,N_4130);
and UO_630 (O_630,N_4538,N_4115);
nor UO_631 (O_631,N_4873,N_4092);
xnor UO_632 (O_632,N_4406,N_4720);
or UO_633 (O_633,N_4643,N_4948);
xor UO_634 (O_634,N_4615,N_4524);
and UO_635 (O_635,N_4856,N_4025);
nand UO_636 (O_636,N_4623,N_4012);
and UO_637 (O_637,N_4289,N_4425);
and UO_638 (O_638,N_4335,N_4015);
nand UO_639 (O_639,N_4340,N_4864);
nor UO_640 (O_640,N_4558,N_4167);
and UO_641 (O_641,N_4354,N_4243);
and UO_642 (O_642,N_4307,N_4174);
or UO_643 (O_643,N_4784,N_4874);
xnor UO_644 (O_644,N_4402,N_4642);
and UO_645 (O_645,N_4598,N_4753);
nand UO_646 (O_646,N_4828,N_4853);
and UO_647 (O_647,N_4620,N_4608);
xnor UO_648 (O_648,N_4469,N_4820);
or UO_649 (O_649,N_4329,N_4227);
or UO_650 (O_650,N_4331,N_4893);
and UO_651 (O_651,N_4269,N_4726);
nor UO_652 (O_652,N_4362,N_4975);
or UO_653 (O_653,N_4809,N_4638);
or UO_654 (O_654,N_4979,N_4843);
and UO_655 (O_655,N_4481,N_4032);
and UO_656 (O_656,N_4390,N_4882);
and UO_657 (O_657,N_4992,N_4639);
nor UO_658 (O_658,N_4065,N_4197);
and UO_659 (O_659,N_4529,N_4841);
nor UO_660 (O_660,N_4384,N_4754);
nand UO_661 (O_661,N_4675,N_4623);
and UO_662 (O_662,N_4896,N_4137);
or UO_663 (O_663,N_4325,N_4491);
nand UO_664 (O_664,N_4194,N_4570);
nor UO_665 (O_665,N_4924,N_4487);
nor UO_666 (O_666,N_4840,N_4182);
or UO_667 (O_667,N_4970,N_4047);
and UO_668 (O_668,N_4874,N_4548);
nor UO_669 (O_669,N_4027,N_4002);
and UO_670 (O_670,N_4956,N_4072);
and UO_671 (O_671,N_4481,N_4961);
or UO_672 (O_672,N_4481,N_4836);
nand UO_673 (O_673,N_4126,N_4271);
nand UO_674 (O_674,N_4557,N_4407);
and UO_675 (O_675,N_4605,N_4852);
xor UO_676 (O_676,N_4862,N_4476);
nand UO_677 (O_677,N_4894,N_4123);
and UO_678 (O_678,N_4298,N_4796);
nor UO_679 (O_679,N_4570,N_4168);
or UO_680 (O_680,N_4406,N_4392);
and UO_681 (O_681,N_4974,N_4206);
nor UO_682 (O_682,N_4890,N_4649);
nor UO_683 (O_683,N_4150,N_4194);
xor UO_684 (O_684,N_4550,N_4777);
xnor UO_685 (O_685,N_4581,N_4214);
and UO_686 (O_686,N_4190,N_4794);
nand UO_687 (O_687,N_4208,N_4178);
nor UO_688 (O_688,N_4448,N_4927);
or UO_689 (O_689,N_4955,N_4157);
nor UO_690 (O_690,N_4010,N_4973);
and UO_691 (O_691,N_4467,N_4074);
nand UO_692 (O_692,N_4210,N_4678);
and UO_693 (O_693,N_4515,N_4578);
or UO_694 (O_694,N_4476,N_4263);
nand UO_695 (O_695,N_4414,N_4012);
nand UO_696 (O_696,N_4273,N_4815);
nor UO_697 (O_697,N_4612,N_4695);
and UO_698 (O_698,N_4751,N_4239);
nor UO_699 (O_699,N_4820,N_4596);
and UO_700 (O_700,N_4532,N_4799);
and UO_701 (O_701,N_4937,N_4627);
nor UO_702 (O_702,N_4190,N_4354);
nor UO_703 (O_703,N_4889,N_4319);
or UO_704 (O_704,N_4541,N_4410);
nand UO_705 (O_705,N_4090,N_4927);
nand UO_706 (O_706,N_4617,N_4275);
nor UO_707 (O_707,N_4260,N_4774);
nor UO_708 (O_708,N_4807,N_4773);
and UO_709 (O_709,N_4689,N_4765);
and UO_710 (O_710,N_4676,N_4122);
nor UO_711 (O_711,N_4408,N_4132);
xor UO_712 (O_712,N_4821,N_4954);
nand UO_713 (O_713,N_4944,N_4305);
or UO_714 (O_714,N_4063,N_4471);
nor UO_715 (O_715,N_4796,N_4153);
and UO_716 (O_716,N_4361,N_4589);
xnor UO_717 (O_717,N_4007,N_4146);
nor UO_718 (O_718,N_4136,N_4203);
nand UO_719 (O_719,N_4658,N_4671);
or UO_720 (O_720,N_4732,N_4729);
or UO_721 (O_721,N_4365,N_4946);
or UO_722 (O_722,N_4037,N_4486);
or UO_723 (O_723,N_4935,N_4862);
or UO_724 (O_724,N_4360,N_4395);
and UO_725 (O_725,N_4866,N_4206);
and UO_726 (O_726,N_4941,N_4635);
or UO_727 (O_727,N_4462,N_4624);
nand UO_728 (O_728,N_4578,N_4316);
or UO_729 (O_729,N_4845,N_4918);
or UO_730 (O_730,N_4319,N_4675);
and UO_731 (O_731,N_4395,N_4096);
and UO_732 (O_732,N_4623,N_4430);
and UO_733 (O_733,N_4143,N_4948);
and UO_734 (O_734,N_4496,N_4100);
nand UO_735 (O_735,N_4533,N_4235);
and UO_736 (O_736,N_4750,N_4645);
or UO_737 (O_737,N_4043,N_4252);
and UO_738 (O_738,N_4496,N_4101);
and UO_739 (O_739,N_4501,N_4489);
nand UO_740 (O_740,N_4876,N_4053);
and UO_741 (O_741,N_4704,N_4764);
nor UO_742 (O_742,N_4296,N_4380);
or UO_743 (O_743,N_4140,N_4300);
and UO_744 (O_744,N_4151,N_4473);
xor UO_745 (O_745,N_4335,N_4347);
or UO_746 (O_746,N_4256,N_4544);
and UO_747 (O_747,N_4721,N_4690);
and UO_748 (O_748,N_4770,N_4441);
nor UO_749 (O_749,N_4789,N_4987);
nor UO_750 (O_750,N_4940,N_4144);
xor UO_751 (O_751,N_4361,N_4079);
nor UO_752 (O_752,N_4945,N_4133);
and UO_753 (O_753,N_4295,N_4861);
or UO_754 (O_754,N_4684,N_4239);
nor UO_755 (O_755,N_4648,N_4848);
and UO_756 (O_756,N_4816,N_4663);
or UO_757 (O_757,N_4744,N_4328);
nor UO_758 (O_758,N_4466,N_4970);
or UO_759 (O_759,N_4641,N_4369);
nand UO_760 (O_760,N_4849,N_4616);
nand UO_761 (O_761,N_4712,N_4182);
and UO_762 (O_762,N_4803,N_4034);
and UO_763 (O_763,N_4249,N_4122);
and UO_764 (O_764,N_4057,N_4105);
and UO_765 (O_765,N_4173,N_4418);
nand UO_766 (O_766,N_4536,N_4071);
xor UO_767 (O_767,N_4886,N_4572);
or UO_768 (O_768,N_4332,N_4441);
xnor UO_769 (O_769,N_4343,N_4188);
nand UO_770 (O_770,N_4107,N_4212);
nor UO_771 (O_771,N_4960,N_4504);
and UO_772 (O_772,N_4903,N_4570);
or UO_773 (O_773,N_4667,N_4556);
nor UO_774 (O_774,N_4902,N_4858);
and UO_775 (O_775,N_4292,N_4208);
nor UO_776 (O_776,N_4779,N_4034);
nor UO_777 (O_777,N_4812,N_4785);
or UO_778 (O_778,N_4136,N_4037);
nor UO_779 (O_779,N_4278,N_4216);
or UO_780 (O_780,N_4344,N_4076);
and UO_781 (O_781,N_4828,N_4631);
nand UO_782 (O_782,N_4161,N_4589);
nand UO_783 (O_783,N_4870,N_4626);
nand UO_784 (O_784,N_4935,N_4204);
and UO_785 (O_785,N_4278,N_4364);
nor UO_786 (O_786,N_4841,N_4731);
nor UO_787 (O_787,N_4621,N_4269);
nor UO_788 (O_788,N_4258,N_4589);
and UO_789 (O_789,N_4030,N_4878);
or UO_790 (O_790,N_4262,N_4481);
nand UO_791 (O_791,N_4691,N_4492);
or UO_792 (O_792,N_4373,N_4375);
or UO_793 (O_793,N_4820,N_4629);
and UO_794 (O_794,N_4654,N_4834);
and UO_795 (O_795,N_4784,N_4906);
or UO_796 (O_796,N_4370,N_4119);
or UO_797 (O_797,N_4833,N_4885);
nand UO_798 (O_798,N_4289,N_4326);
or UO_799 (O_799,N_4477,N_4931);
and UO_800 (O_800,N_4624,N_4108);
or UO_801 (O_801,N_4726,N_4081);
or UO_802 (O_802,N_4139,N_4181);
nand UO_803 (O_803,N_4964,N_4901);
or UO_804 (O_804,N_4713,N_4230);
xnor UO_805 (O_805,N_4892,N_4988);
or UO_806 (O_806,N_4229,N_4169);
and UO_807 (O_807,N_4997,N_4157);
or UO_808 (O_808,N_4687,N_4343);
or UO_809 (O_809,N_4640,N_4853);
nor UO_810 (O_810,N_4385,N_4451);
nor UO_811 (O_811,N_4062,N_4147);
and UO_812 (O_812,N_4690,N_4375);
nand UO_813 (O_813,N_4999,N_4104);
nand UO_814 (O_814,N_4446,N_4278);
nor UO_815 (O_815,N_4192,N_4324);
or UO_816 (O_816,N_4816,N_4420);
xor UO_817 (O_817,N_4717,N_4780);
or UO_818 (O_818,N_4006,N_4906);
nor UO_819 (O_819,N_4713,N_4507);
and UO_820 (O_820,N_4752,N_4720);
and UO_821 (O_821,N_4848,N_4179);
or UO_822 (O_822,N_4983,N_4708);
nand UO_823 (O_823,N_4098,N_4092);
or UO_824 (O_824,N_4083,N_4093);
nor UO_825 (O_825,N_4393,N_4099);
xnor UO_826 (O_826,N_4098,N_4209);
and UO_827 (O_827,N_4782,N_4626);
and UO_828 (O_828,N_4840,N_4662);
or UO_829 (O_829,N_4127,N_4532);
and UO_830 (O_830,N_4605,N_4749);
nor UO_831 (O_831,N_4976,N_4789);
nor UO_832 (O_832,N_4774,N_4390);
nand UO_833 (O_833,N_4250,N_4064);
nor UO_834 (O_834,N_4534,N_4098);
and UO_835 (O_835,N_4572,N_4692);
nor UO_836 (O_836,N_4605,N_4062);
and UO_837 (O_837,N_4595,N_4857);
and UO_838 (O_838,N_4241,N_4705);
xnor UO_839 (O_839,N_4145,N_4878);
nor UO_840 (O_840,N_4589,N_4053);
nand UO_841 (O_841,N_4030,N_4685);
and UO_842 (O_842,N_4619,N_4535);
nor UO_843 (O_843,N_4509,N_4198);
nor UO_844 (O_844,N_4305,N_4384);
and UO_845 (O_845,N_4972,N_4388);
and UO_846 (O_846,N_4987,N_4947);
xnor UO_847 (O_847,N_4190,N_4337);
and UO_848 (O_848,N_4216,N_4391);
nor UO_849 (O_849,N_4433,N_4527);
nand UO_850 (O_850,N_4487,N_4112);
nand UO_851 (O_851,N_4102,N_4474);
nand UO_852 (O_852,N_4352,N_4089);
or UO_853 (O_853,N_4413,N_4446);
or UO_854 (O_854,N_4757,N_4071);
and UO_855 (O_855,N_4788,N_4726);
nor UO_856 (O_856,N_4332,N_4088);
nor UO_857 (O_857,N_4439,N_4583);
or UO_858 (O_858,N_4495,N_4288);
xnor UO_859 (O_859,N_4658,N_4548);
or UO_860 (O_860,N_4283,N_4628);
nor UO_861 (O_861,N_4841,N_4109);
and UO_862 (O_862,N_4246,N_4020);
and UO_863 (O_863,N_4580,N_4105);
nor UO_864 (O_864,N_4827,N_4765);
nor UO_865 (O_865,N_4792,N_4631);
and UO_866 (O_866,N_4214,N_4960);
or UO_867 (O_867,N_4231,N_4079);
or UO_868 (O_868,N_4583,N_4507);
or UO_869 (O_869,N_4120,N_4304);
or UO_870 (O_870,N_4975,N_4833);
nor UO_871 (O_871,N_4115,N_4459);
or UO_872 (O_872,N_4039,N_4657);
and UO_873 (O_873,N_4392,N_4399);
and UO_874 (O_874,N_4888,N_4111);
and UO_875 (O_875,N_4095,N_4078);
nand UO_876 (O_876,N_4958,N_4580);
or UO_877 (O_877,N_4051,N_4212);
and UO_878 (O_878,N_4126,N_4284);
nand UO_879 (O_879,N_4358,N_4675);
nand UO_880 (O_880,N_4468,N_4804);
nor UO_881 (O_881,N_4979,N_4409);
and UO_882 (O_882,N_4385,N_4752);
nand UO_883 (O_883,N_4156,N_4395);
or UO_884 (O_884,N_4588,N_4496);
xnor UO_885 (O_885,N_4805,N_4590);
nand UO_886 (O_886,N_4084,N_4760);
and UO_887 (O_887,N_4031,N_4659);
nand UO_888 (O_888,N_4100,N_4763);
nor UO_889 (O_889,N_4067,N_4604);
nand UO_890 (O_890,N_4958,N_4057);
nor UO_891 (O_891,N_4782,N_4254);
or UO_892 (O_892,N_4661,N_4298);
and UO_893 (O_893,N_4828,N_4658);
nand UO_894 (O_894,N_4504,N_4595);
or UO_895 (O_895,N_4075,N_4528);
or UO_896 (O_896,N_4892,N_4237);
and UO_897 (O_897,N_4870,N_4455);
nand UO_898 (O_898,N_4346,N_4656);
or UO_899 (O_899,N_4345,N_4965);
xnor UO_900 (O_900,N_4136,N_4342);
nand UO_901 (O_901,N_4477,N_4039);
nor UO_902 (O_902,N_4486,N_4261);
or UO_903 (O_903,N_4981,N_4283);
and UO_904 (O_904,N_4937,N_4256);
and UO_905 (O_905,N_4724,N_4524);
or UO_906 (O_906,N_4647,N_4162);
nor UO_907 (O_907,N_4268,N_4911);
nand UO_908 (O_908,N_4503,N_4909);
or UO_909 (O_909,N_4420,N_4406);
and UO_910 (O_910,N_4421,N_4668);
or UO_911 (O_911,N_4486,N_4009);
or UO_912 (O_912,N_4534,N_4455);
or UO_913 (O_913,N_4391,N_4161);
nor UO_914 (O_914,N_4201,N_4688);
and UO_915 (O_915,N_4513,N_4585);
or UO_916 (O_916,N_4309,N_4288);
and UO_917 (O_917,N_4699,N_4730);
nor UO_918 (O_918,N_4071,N_4019);
nor UO_919 (O_919,N_4227,N_4711);
nand UO_920 (O_920,N_4541,N_4606);
nor UO_921 (O_921,N_4665,N_4406);
nor UO_922 (O_922,N_4335,N_4102);
nor UO_923 (O_923,N_4559,N_4556);
or UO_924 (O_924,N_4867,N_4953);
nand UO_925 (O_925,N_4996,N_4568);
nor UO_926 (O_926,N_4811,N_4599);
xor UO_927 (O_927,N_4758,N_4287);
nor UO_928 (O_928,N_4418,N_4649);
or UO_929 (O_929,N_4988,N_4032);
and UO_930 (O_930,N_4081,N_4730);
or UO_931 (O_931,N_4541,N_4360);
or UO_932 (O_932,N_4292,N_4483);
or UO_933 (O_933,N_4535,N_4356);
or UO_934 (O_934,N_4444,N_4724);
nor UO_935 (O_935,N_4539,N_4604);
or UO_936 (O_936,N_4723,N_4100);
nand UO_937 (O_937,N_4250,N_4982);
and UO_938 (O_938,N_4095,N_4190);
or UO_939 (O_939,N_4090,N_4486);
nor UO_940 (O_940,N_4101,N_4784);
xor UO_941 (O_941,N_4230,N_4792);
and UO_942 (O_942,N_4079,N_4127);
or UO_943 (O_943,N_4235,N_4162);
or UO_944 (O_944,N_4235,N_4161);
xor UO_945 (O_945,N_4834,N_4694);
or UO_946 (O_946,N_4090,N_4800);
or UO_947 (O_947,N_4509,N_4883);
xor UO_948 (O_948,N_4511,N_4240);
xnor UO_949 (O_949,N_4413,N_4914);
xor UO_950 (O_950,N_4742,N_4473);
and UO_951 (O_951,N_4892,N_4442);
and UO_952 (O_952,N_4312,N_4786);
xnor UO_953 (O_953,N_4234,N_4906);
or UO_954 (O_954,N_4892,N_4533);
xor UO_955 (O_955,N_4417,N_4340);
and UO_956 (O_956,N_4697,N_4922);
and UO_957 (O_957,N_4022,N_4255);
and UO_958 (O_958,N_4076,N_4441);
nand UO_959 (O_959,N_4422,N_4233);
and UO_960 (O_960,N_4232,N_4142);
or UO_961 (O_961,N_4626,N_4072);
nand UO_962 (O_962,N_4620,N_4406);
nand UO_963 (O_963,N_4712,N_4095);
and UO_964 (O_964,N_4349,N_4509);
nand UO_965 (O_965,N_4000,N_4663);
or UO_966 (O_966,N_4332,N_4894);
and UO_967 (O_967,N_4572,N_4559);
nor UO_968 (O_968,N_4279,N_4341);
or UO_969 (O_969,N_4647,N_4135);
or UO_970 (O_970,N_4993,N_4334);
or UO_971 (O_971,N_4863,N_4613);
nand UO_972 (O_972,N_4518,N_4662);
nor UO_973 (O_973,N_4495,N_4028);
or UO_974 (O_974,N_4969,N_4561);
nand UO_975 (O_975,N_4619,N_4257);
nand UO_976 (O_976,N_4604,N_4939);
nor UO_977 (O_977,N_4527,N_4847);
nor UO_978 (O_978,N_4192,N_4015);
and UO_979 (O_979,N_4253,N_4879);
and UO_980 (O_980,N_4420,N_4937);
and UO_981 (O_981,N_4500,N_4995);
and UO_982 (O_982,N_4400,N_4002);
nand UO_983 (O_983,N_4188,N_4115);
nor UO_984 (O_984,N_4588,N_4063);
xnor UO_985 (O_985,N_4976,N_4756);
or UO_986 (O_986,N_4050,N_4802);
nand UO_987 (O_987,N_4850,N_4549);
xnor UO_988 (O_988,N_4715,N_4956);
nor UO_989 (O_989,N_4495,N_4070);
nand UO_990 (O_990,N_4440,N_4664);
and UO_991 (O_991,N_4898,N_4987);
or UO_992 (O_992,N_4697,N_4260);
nor UO_993 (O_993,N_4121,N_4409);
or UO_994 (O_994,N_4734,N_4400);
nor UO_995 (O_995,N_4494,N_4734);
nand UO_996 (O_996,N_4843,N_4755);
and UO_997 (O_997,N_4681,N_4773);
nand UO_998 (O_998,N_4226,N_4846);
nand UO_999 (O_999,N_4949,N_4209);
endmodule