module basic_750_5000_1000_10_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_441,In_654);
and U1 (N_1,In_424,In_144);
and U2 (N_2,In_474,In_621);
nand U3 (N_3,In_187,In_664);
nand U4 (N_4,In_205,In_562);
or U5 (N_5,In_475,In_128);
nor U6 (N_6,In_423,In_302);
and U7 (N_7,In_135,In_356);
nor U8 (N_8,In_100,In_466);
or U9 (N_9,In_733,In_702);
and U10 (N_10,In_172,In_674);
nor U11 (N_11,In_617,In_668);
and U12 (N_12,In_241,In_207);
nand U13 (N_13,In_609,In_666);
nor U14 (N_14,In_595,In_245);
nor U15 (N_15,In_583,In_578);
and U16 (N_16,In_684,In_122);
nand U17 (N_17,In_107,In_274);
and U18 (N_18,In_115,In_27);
or U19 (N_19,In_159,In_382);
nand U20 (N_20,In_734,In_735);
nand U21 (N_21,In_171,In_535);
nor U22 (N_22,In_141,In_667);
and U23 (N_23,In_66,In_426);
and U24 (N_24,In_386,In_142);
or U25 (N_25,In_532,In_322);
nand U26 (N_26,In_297,In_43);
or U27 (N_27,In_248,In_581);
and U28 (N_28,In_83,In_251);
and U29 (N_29,In_231,In_148);
or U30 (N_30,In_299,In_565);
nand U31 (N_31,In_346,In_476);
or U32 (N_32,In_606,In_634);
and U33 (N_33,In_449,In_513);
nor U34 (N_34,In_269,In_74);
and U35 (N_35,In_61,In_614);
and U36 (N_36,In_727,In_95);
and U37 (N_37,In_511,In_427);
and U38 (N_38,In_58,In_292);
nand U39 (N_39,In_619,In_71);
nor U40 (N_40,In_3,In_25);
nor U41 (N_41,In_549,In_166);
nand U42 (N_42,In_226,In_362);
nand U43 (N_43,In_678,In_216);
and U44 (N_44,In_252,In_652);
or U45 (N_45,In_452,In_94);
nor U46 (N_46,In_536,In_429);
and U47 (N_47,In_594,In_335);
or U48 (N_48,In_454,In_214);
nor U49 (N_49,In_92,In_432);
and U50 (N_50,In_331,In_194);
and U51 (N_51,In_742,In_316);
nand U52 (N_52,In_747,In_604);
nand U53 (N_53,In_105,In_30);
nor U54 (N_54,In_255,In_208);
nand U55 (N_55,In_264,In_648);
nand U56 (N_56,In_84,In_661);
nand U57 (N_57,In_591,In_448);
nor U58 (N_58,In_360,In_109);
and U59 (N_59,In_163,In_39);
and U60 (N_60,In_85,In_601);
and U61 (N_61,In_101,In_263);
nor U62 (N_62,In_314,In_398);
nor U63 (N_63,In_552,In_239);
xnor U64 (N_64,In_640,In_183);
nand U65 (N_65,In_701,In_64);
nand U66 (N_66,In_36,In_193);
nand U67 (N_67,In_695,In_313);
and U68 (N_68,In_519,In_537);
nand U69 (N_69,In_560,In_384);
nand U70 (N_70,In_390,In_342);
nor U71 (N_71,In_479,In_660);
xnor U72 (N_72,In_553,In_143);
nand U73 (N_73,In_87,In_202);
nand U74 (N_74,In_21,In_180);
nand U75 (N_75,In_259,In_206);
nand U76 (N_76,In_410,In_718);
nor U77 (N_77,In_308,In_315);
and U78 (N_78,In_372,In_408);
nor U79 (N_79,In_28,In_98);
nand U80 (N_80,In_195,In_744);
nor U81 (N_81,In_662,In_675);
nor U82 (N_82,In_131,In_147);
nand U83 (N_83,In_364,In_355);
or U84 (N_84,In_749,In_374);
and U85 (N_85,In_284,In_289);
nand U86 (N_86,In_442,In_499);
nor U87 (N_87,In_687,In_124);
nor U88 (N_88,In_732,In_280);
nor U89 (N_89,In_510,In_444);
or U90 (N_90,In_602,In_104);
and U91 (N_91,In_724,In_254);
nand U92 (N_92,In_544,In_305);
and U93 (N_93,In_86,In_430);
and U94 (N_94,In_572,In_670);
nor U95 (N_95,In_433,In_75);
nor U96 (N_96,In_9,In_389);
or U97 (N_97,In_458,In_35);
nor U98 (N_98,In_65,In_230);
xnor U99 (N_99,In_392,In_638);
nor U100 (N_100,In_170,In_707);
or U101 (N_101,In_396,In_420);
or U102 (N_102,In_45,In_484);
or U103 (N_103,In_385,In_469);
or U104 (N_104,In_567,In_130);
nor U105 (N_105,In_542,In_233);
and U106 (N_106,In_406,In_19);
nand U107 (N_107,In_76,In_298);
nand U108 (N_108,In_459,In_34);
or U109 (N_109,In_689,In_137);
nand U110 (N_110,In_691,In_505);
or U111 (N_111,In_78,In_268);
or U112 (N_112,In_447,In_464);
or U113 (N_113,In_696,In_63);
nand U114 (N_114,In_743,In_278);
or U115 (N_115,In_373,In_630);
nor U116 (N_116,In_598,In_51);
nand U117 (N_117,In_445,In_577);
nand U118 (N_118,In_134,In_303);
nor U119 (N_119,In_222,In_157);
nand U120 (N_120,In_411,In_726);
nand U121 (N_121,In_24,In_82);
nand U122 (N_122,In_324,In_326);
and U123 (N_123,In_132,In_688);
or U124 (N_124,In_29,In_267);
nand U125 (N_125,In_38,In_629);
or U126 (N_126,In_12,In_234);
and U127 (N_127,In_174,In_319);
nand U128 (N_128,In_57,In_462);
nor U129 (N_129,In_185,In_123);
nor U130 (N_130,In_439,In_482);
or U131 (N_131,In_164,In_238);
or U132 (N_132,In_561,In_497);
nor U133 (N_133,In_490,In_540);
nor U134 (N_134,In_498,In_329);
or U135 (N_135,In_261,In_515);
and U136 (N_136,In_327,In_626);
nand U137 (N_137,In_470,In_271);
and U138 (N_138,In_4,In_196);
nor U139 (N_139,In_120,In_73);
or U140 (N_140,In_333,In_600);
or U141 (N_141,In_375,In_70);
and U142 (N_142,In_473,In_112);
or U143 (N_143,In_745,In_69);
nor U144 (N_144,In_547,In_309);
nor U145 (N_145,In_677,In_291);
xor U146 (N_146,In_179,In_443);
nand U147 (N_147,In_173,In_161);
nand U148 (N_148,In_41,In_113);
and U149 (N_149,In_8,In_68);
and U150 (N_150,In_698,In_203);
or U151 (N_151,In_740,In_610);
nand U152 (N_152,In_438,In_463);
nor U153 (N_153,In_79,In_690);
nor U154 (N_154,In_242,In_527);
nand U155 (N_155,In_573,In_188);
and U156 (N_156,In_275,In_627);
nand U157 (N_157,In_225,In_388);
and U158 (N_158,In_672,In_383);
and U159 (N_159,In_489,In_359);
nand U160 (N_160,In_538,In_720);
or U161 (N_161,In_746,In_541);
and U162 (N_162,In_571,In_88);
nor U163 (N_163,In_312,In_425);
or U164 (N_164,In_223,In_415);
and U165 (N_165,In_421,In_692);
and U166 (N_166,In_340,In_414);
nor U167 (N_167,In_184,In_31);
nand U168 (N_168,In_713,In_201);
or U169 (N_169,In_647,In_471);
nand U170 (N_170,In_217,In_545);
or U171 (N_171,In_32,In_270);
or U172 (N_172,In_686,In_114);
and U173 (N_173,In_468,In_62);
nor U174 (N_174,In_26,In_139);
and U175 (N_175,In_300,In_256);
nor U176 (N_176,In_108,In_546);
nand U177 (N_177,In_265,In_198);
and U178 (N_178,In_91,In_697);
or U179 (N_179,In_282,In_221);
nand U180 (N_180,In_244,In_635);
and U181 (N_181,In_150,In_646);
or U182 (N_182,In_523,In_461);
or U183 (N_183,In_149,In_487);
and U184 (N_184,In_628,In_199);
or U185 (N_185,In_491,In_60);
or U186 (N_186,In_422,In_262);
and U187 (N_187,In_368,In_190);
nor U188 (N_188,In_50,In_435);
and U189 (N_189,In_710,In_357);
or U190 (N_190,In_679,In_518);
or U191 (N_191,In_77,In_323);
nand U192 (N_192,In_126,In_676);
and U193 (N_193,In_683,In_637);
or U194 (N_194,In_237,In_493);
or U195 (N_195,In_402,In_22);
or U196 (N_196,In_15,In_680);
or U197 (N_197,In_644,In_236);
nor U198 (N_198,In_555,In_228);
and U199 (N_199,In_310,In_731);
or U200 (N_200,In_328,In_723);
nand U201 (N_201,In_266,In_46);
xor U202 (N_202,In_11,In_729);
nand U203 (N_203,In_558,In_153);
nand U204 (N_204,In_419,In_528);
nand U205 (N_205,In_703,In_494);
or U206 (N_206,In_119,In_370);
or U207 (N_207,In_394,In_343);
and U208 (N_208,In_492,In_559);
nor U209 (N_209,In_706,In_645);
nor U210 (N_210,In_719,In_611);
nand U211 (N_211,In_453,In_397);
nand U212 (N_212,In_632,In_440);
and U213 (N_213,In_520,In_240);
and U214 (N_214,In_564,In_568);
xor U215 (N_215,In_334,In_283);
nor U216 (N_216,In_377,In_344);
or U217 (N_217,In_566,In_349);
nand U218 (N_218,In_365,In_550);
nor U219 (N_219,In_13,In_465);
or U220 (N_220,In_127,In_55);
nand U221 (N_221,In_514,In_133);
or U222 (N_222,In_1,In_579);
nand U223 (N_223,In_138,In_279);
nand U224 (N_224,In_665,In_249);
or U225 (N_225,In_739,In_320);
and U226 (N_226,In_529,In_605);
nand U227 (N_227,In_431,In_507);
and U228 (N_228,In_158,In_533);
or U229 (N_229,In_250,In_176);
nand U230 (N_230,In_56,In_480);
or U231 (N_231,In_705,In_146);
nand U232 (N_232,In_508,In_590);
nand U233 (N_233,In_6,In_220);
nand U234 (N_234,In_737,In_363);
nor U235 (N_235,In_391,In_294);
or U236 (N_236,In_296,In_556);
nand U237 (N_237,In_592,In_227);
nand U238 (N_238,In_403,In_496);
nand U239 (N_239,In_636,In_721);
xor U240 (N_240,In_409,In_53);
or U241 (N_241,In_44,In_257);
nor U242 (N_242,In_512,In_593);
or U243 (N_243,In_286,In_204);
nor U244 (N_244,In_67,In_694);
nor U245 (N_245,In_699,In_129);
nor U246 (N_246,In_106,In_273);
nand U247 (N_247,In_481,In_0);
nand U248 (N_248,In_526,In_521);
nand U249 (N_249,In_615,In_277);
nor U250 (N_250,In_612,In_393);
or U251 (N_251,In_708,In_118);
and U252 (N_252,In_387,In_318);
and U253 (N_253,In_418,In_378);
and U254 (N_254,In_395,In_99);
and U255 (N_255,In_716,In_584);
nand U256 (N_256,In_81,In_290);
nand U257 (N_257,In_301,In_658);
and U258 (N_258,In_502,In_500);
nor U259 (N_259,In_140,In_486);
and U260 (N_260,In_243,In_209);
and U261 (N_261,In_437,In_399);
or U262 (N_262,In_693,In_625);
or U263 (N_263,In_436,In_20);
nand U264 (N_264,In_178,In_715);
or U265 (N_265,In_748,In_369);
nand U266 (N_266,In_455,In_434);
or U267 (N_267,In_16,In_192);
or U268 (N_268,In_506,In_597);
nor U269 (N_269,In_211,In_253);
and U270 (N_270,In_14,In_407);
or U271 (N_271,In_175,In_288);
and U272 (N_272,In_599,In_416);
and U273 (N_273,In_371,In_111);
nand U274 (N_274,In_162,In_376);
or U275 (N_275,In_451,In_714);
and U276 (N_276,In_224,In_557);
nand U277 (N_277,In_405,In_154);
nor U278 (N_278,In_307,In_186);
and U279 (N_279,In_167,In_285);
nor U280 (N_280,In_657,In_712);
nand U281 (N_281,In_582,In_446);
and U282 (N_282,In_235,In_151);
nand U283 (N_283,In_522,In_304);
nand U284 (N_284,In_563,In_93);
or U285 (N_285,In_367,In_295);
and U286 (N_286,In_350,In_306);
nand U287 (N_287,In_125,In_197);
or U288 (N_288,In_608,In_649);
or U289 (N_289,In_650,In_229);
nand U290 (N_290,In_642,In_246);
and U291 (N_291,In_495,In_345);
nand U292 (N_292,In_293,In_603);
nor U293 (N_293,In_671,In_110);
and U294 (N_294,In_352,In_40);
nor U295 (N_295,In_189,In_478);
or U296 (N_296,In_358,In_155);
and U297 (N_297,In_450,In_413);
and U298 (N_298,In_219,In_589);
and U299 (N_299,In_49,In_607);
and U300 (N_300,In_210,In_741);
and U301 (N_301,In_539,In_90);
nor U302 (N_302,In_7,In_400);
nor U303 (N_303,In_457,In_191);
nand U304 (N_304,In_639,In_738);
or U305 (N_305,In_258,In_704);
nor U306 (N_306,In_287,In_18);
nand U307 (N_307,In_417,In_669);
nand U308 (N_308,In_483,In_655);
or U309 (N_309,In_569,In_48);
and U310 (N_310,In_682,In_169);
nor U311 (N_311,In_624,In_23);
or U312 (N_312,In_103,In_136);
nand U313 (N_313,In_530,In_213);
and U314 (N_314,In_276,In_631);
or U315 (N_315,In_663,In_548);
or U316 (N_316,In_722,In_700);
and U317 (N_317,In_348,In_353);
xnor U318 (N_318,In_47,In_485);
and U319 (N_319,In_576,In_570);
nand U320 (N_320,In_218,In_354);
nor U321 (N_321,In_260,In_232);
or U322 (N_322,In_428,In_351);
nor U323 (N_323,In_97,In_456);
and U324 (N_324,In_89,In_311);
and U325 (N_325,In_551,In_156);
nor U326 (N_326,In_717,In_622);
nand U327 (N_327,In_531,In_200);
nor U328 (N_328,In_633,In_10);
nor U329 (N_329,In_380,In_339);
or U330 (N_330,In_586,In_325);
or U331 (N_331,In_33,In_623);
xnor U332 (N_332,In_80,In_341);
and U333 (N_333,In_580,In_534);
and U334 (N_334,In_59,In_477);
or U335 (N_335,In_121,In_587);
or U336 (N_336,In_616,In_596);
and U337 (N_337,In_585,In_117);
nand U338 (N_338,In_96,In_711);
and U339 (N_339,In_182,In_177);
and U340 (N_340,In_338,In_525);
nor U341 (N_341,In_503,In_575);
nand U342 (N_342,In_467,In_736);
nor U343 (N_343,In_160,In_347);
or U344 (N_344,In_332,In_643);
nand U345 (N_345,In_728,In_17);
nor U346 (N_346,In_412,In_651);
nand U347 (N_347,In_379,In_2);
or U348 (N_348,In_181,In_488);
and U349 (N_349,In_653,In_366);
or U350 (N_350,In_381,In_401);
and U351 (N_351,In_212,In_618);
or U352 (N_352,In_543,In_509);
or U353 (N_353,In_152,In_247);
and U354 (N_354,In_54,In_52);
nor U355 (N_355,In_102,In_725);
or U356 (N_356,In_361,In_681);
and U357 (N_357,In_472,In_516);
or U358 (N_358,In_709,In_336);
and U359 (N_359,In_501,In_321);
xnor U360 (N_360,In_337,In_116);
nor U361 (N_361,In_168,In_404);
and U362 (N_362,In_145,In_517);
or U363 (N_363,In_165,In_317);
nand U364 (N_364,In_5,In_215);
or U365 (N_365,In_72,In_588);
nor U366 (N_366,In_37,In_554);
nand U367 (N_367,In_574,In_504);
nand U368 (N_368,In_42,In_685);
or U369 (N_369,In_659,In_272);
nor U370 (N_370,In_730,In_613);
and U371 (N_371,In_673,In_524);
nor U372 (N_372,In_656,In_281);
nand U373 (N_373,In_330,In_641);
and U374 (N_374,In_620,In_460);
nand U375 (N_375,In_191,In_310);
nor U376 (N_376,In_143,In_697);
nor U377 (N_377,In_411,In_713);
or U378 (N_378,In_746,In_47);
nand U379 (N_379,In_666,In_232);
nor U380 (N_380,In_86,In_552);
and U381 (N_381,In_454,In_701);
or U382 (N_382,In_622,In_89);
nand U383 (N_383,In_412,In_688);
nor U384 (N_384,In_92,In_346);
nor U385 (N_385,In_381,In_672);
or U386 (N_386,In_255,In_245);
and U387 (N_387,In_211,In_183);
and U388 (N_388,In_251,In_719);
or U389 (N_389,In_195,In_197);
or U390 (N_390,In_163,In_66);
nor U391 (N_391,In_690,In_361);
nor U392 (N_392,In_428,In_432);
nor U393 (N_393,In_568,In_683);
nor U394 (N_394,In_704,In_583);
nor U395 (N_395,In_358,In_578);
nand U396 (N_396,In_727,In_550);
nor U397 (N_397,In_404,In_439);
nand U398 (N_398,In_706,In_704);
nand U399 (N_399,In_67,In_718);
nand U400 (N_400,In_416,In_137);
and U401 (N_401,In_433,In_21);
xnor U402 (N_402,In_685,In_288);
nor U403 (N_403,In_722,In_509);
nand U404 (N_404,In_711,In_233);
and U405 (N_405,In_113,In_225);
and U406 (N_406,In_715,In_284);
nor U407 (N_407,In_629,In_361);
nor U408 (N_408,In_138,In_155);
nor U409 (N_409,In_518,In_27);
and U410 (N_410,In_394,In_558);
or U411 (N_411,In_265,In_70);
and U412 (N_412,In_52,In_214);
nor U413 (N_413,In_631,In_735);
or U414 (N_414,In_26,In_578);
or U415 (N_415,In_53,In_506);
and U416 (N_416,In_693,In_220);
or U417 (N_417,In_510,In_570);
and U418 (N_418,In_680,In_166);
or U419 (N_419,In_582,In_597);
and U420 (N_420,In_535,In_684);
nand U421 (N_421,In_306,In_172);
or U422 (N_422,In_662,In_19);
nor U423 (N_423,In_288,In_419);
nand U424 (N_424,In_442,In_659);
nand U425 (N_425,In_639,In_171);
and U426 (N_426,In_677,In_462);
or U427 (N_427,In_97,In_483);
nor U428 (N_428,In_570,In_124);
nor U429 (N_429,In_364,In_701);
and U430 (N_430,In_548,In_717);
nor U431 (N_431,In_61,In_294);
or U432 (N_432,In_528,In_500);
or U433 (N_433,In_280,In_355);
nor U434 (N_434,In_668,In_329);
or U435 (N_435,In_288,In_97);
nor U436 (N_436,In_537,In_267);
nor U437 (N_437,In_221,In_239);
xor U438 (N_438,In_495,In_123);
and U439 (N_439,In_18,In_266);
and U440 (N_440,In_716,In_432);
nand U441 (N_441,In_529,In_198);
and U442 (N_442,In_422,In_483);
and U443 (N_443,In_698,In_662);
and U444 (N_444,In_411,In_663);
xnor U445 (N_445,In_625,In_286);
and U446 (N_446,In_436,In_124);
nand U447 (N_447,In_187,In_330);
and U448 (N_448,In_613,In_169);
nand U449 (N_449,In_282,In_716);
nand U450 (N_450,In_286,In_50);
or U451 (N_451,In_31,In_134);
nand U452 (N_452,In_645,In_314);
and U453 (N_453,In_192,In_427);
xnor U454 (N_454,In_483,In_334);
and U455 (N_455,In_6,In_358);
or U456 (N_456,In_625,In_405);
or U457 (N_457,In_724,In_494);
nand U458 (N_458,In_13,In_421);
nand U459 (N_459,In_55,In_247);
nor U460 (N_460,In_656,In_1);
or U461 (N_461,In_699,In_7);
nor U462 (N_462,In_55,In_695);
nor U463 (N_463,In_140,In_593);
and U464 (N_464,In_213,In_108);
and U465 (N_465,In_589,In_432);
nor U466 (N_466,In_130,In_75);
nor U467 (N_467,In_49,In_521);
or U468 (N_468,In_185,In_515);
nand U469 (N_469,In_219,In_448);
nand U470 (N_470,In_332,In_39);
nor U471 (N_471,In_495,In_202);
or U472 (N_472,In_189,In_597);
nor U473 (N_473,In_316,In_591);
nor U474 (N_474,In_331,In_554);
nand U475 (N_475,In_339,In_425);
or U476 (N_476,In_381,In_572);
nand U477 (N_477,In_542,In_396);
or U478 (N_478,In_205,In_85);
nand U479 (N_479,In_61,In_113);
nor U480 (N_480,In_558,In_292);
or U481 (N_481,In_577,In_532);
nand U482 (N_482,In_273,In_534);
nand U483 (N_483,In_733,In_599);
and U484 (N_484,In_677,In_499);
nor U485 (N_485,In_25,In_301);
xor U486 (N_486,In_294,In_573);
or U487 (N_487,In_225,In_631);
nor U488 (N_488,In_690,In_214);
or U489 (N_489,In_470,In_418);
and U490 (N_490,In_112,In_706);
nor U491 (N_491,In_357,In_370);
nand U492 (N_492,In_197,In_727);
and U493 (N_493,In_131,In_412);
nand U494 (N_494,In_406,In_651);
nand U495 (N_495,In_282,In_525);
and U496 (N_496,In_537,In_351);
or U497 (N_497,In_647,In_94);
and U498 (N_498,In_157,In_18);
and U499 (N_499,In_624,In_492);
nand U500 (N_500,N_430,N_471);
nand U501 (N_501,N_329,N_289);
and U502 (N_502,N_168,N_438);
and U503 (N_503,N_424,N_335);
and U504 (N_504,N_97,N_345);
or U505 (N_505,N_298,N_328);
and U506 (N_506,N_91,N_326);
nand U507 (N_507,N_419,N_316);
nand U508 (N_508,N_140,N_337);
nand U509 (N_509,N_384,N_201);
or U510 (N_510,N_407,N_92);
and U511 (N_511,N_295,N_347);
and U512 (N_512,N_404,N_374);
or U513 (N_513,N_477,N_36);
nor U514 (N_514,N_302,N_322);
and U515 (N_515,N_285,N_400);
or U516 (N_516,N_320,N_389);
nor U517 (N_517,N_34,N_358);
and U518 (N_518,N_78,N_21);
or U519 (N_519,N_169,N_309);
and U520 (N_520,N_236,N_213);
nor U521 (N_521,N_293,N_120);
and U522 (N_522,N_139,N_3);
or U523 (N_523,N_11,N_283);
and U524 (N_524,N_25,N_127);
and U525 (N_525,N_472,N_207);
nand U526 (N_526,N_95,N_223);
nor U527 (N_527,N_147,N_451);
or U528 (N_528,N_495,N_107);
or U529 (N_529,N_184,N_216);
and U530 (N_530,N_167,N_24);
and U531 (N_531,N_143,N_432);
and U532 (N_532,N_177,N_359);
nor U533 (N_533,N_490,N_195);
nor U534 (N_534,N_254,N_173);
and U535 (N_535,N_277,N_255);
and U536 (N_536,N_257,N_376);
or U537 (N_537,N_391,N_408);
nand U538 (N_538,N_245,N_398);
or U539 (N_539,N_193,N_148);
nand U540 (N_540,N_416,N_146);
or U541 (N_541,N_48,N_80);
or U542 (N_542,N_464,N_74);
or U543 (N_543,N_222,N_450);
and U544 (N_544,N_403,N_2);
or U545 (N_545,N_175,N_69);
nor U546 (N_546,N_433,N_323);
nor U547 (N_547,N_394,N_484);
or U548 (N_548,N_83,N_275);
or U549 (N_549,N_145,N_237);
nand U550 (N_550,N_434,N_33);
and U551 (N_551,N_138,N_333);
or U552 (N_552,N_470,N_230);
or U553 (N_553,N_116,N_395);
and U554 (N_554,N_258,N_38);
nand U555 (N_555,N_281,N_498);
xnor U556 (N_556,N_499,N_387);
nand U557 (N_557,N_410,N_284);
or U558 (N_558,N_288,N_153);
and U559 (N_559,N_462,N_104);
or U560 (N_560,N_194,N_378);
or U561 (N_561,N_212,N_312);
nand U562 (N_562,N_105,N_160);
or U563 (N_563,N_415,N_436);
or U564 (N_564,N_343,N_87);
or U565 (N_565,N_411,N_109);
nand U566 (N_566,N_493,N_456);
nand U567 (N_567,N_414,N_150);
or U568 (N_568,N_20,N_152);
nand U569 (N_569,N_181,N_227);
or U570 (N_570,N_6,N_55);
nor U571 (N_571,N_297,N_70);
nand U572 (N_572,N_242,N_31);
nor U573 (N_573,N_413,N_474);
nor U574 (N_574,N_187,N_57);
and U575 (N_575,N_304,N_392);
nand U576 (N_576,N_4,N_26);
nand U577 (N_577,N_52,N_369);
or U578 (N_578,N_496,N_64);
nor U579 (N_579,N_355,N_292);
nor U580 (N_580,N_8,N_278);
or U581 (N_581,N_235,N_303);
nor U582 (N_582,N_14,N_294);
and U583 (N_583,N_136,N_249);
nand U584 (N_584,N_202,N_30);
nor U585 (N_585,N_75,N_122);
or U586 (N_586,N_142,N_252);
nor U587 (N_587,N_179,N_115);
nor U588 (N_588,N_367,N_307);
or U589 (N_589,N_190,N_117);
nor U590 (N_590,N_112,N_94);
or U591 (N_591,N_199,N_126);
and U592 (N_592,N_189,N_290);
or U593 (N_593,N_267,N_132);
nand U594 (N_594,N_98,N_204);
xor U595 (N_595,N_17,N_100);
nor U596 (N_596,N_185,N_421);
nand U597 (N_597,N_10,N_487);
and U598 (N_598,N_377,N_176);
nor U599 (N_599,N_89,N_274);
or U600 (N_600,N_338,N_197);
nand U601 (N_601,N_50,N_271);
nor U602 (N_602,N_119,N_68);
nand U603 (N_603,N_82,N_299);
or U604 (N_604,N_319,N_330);
nand U605 (N_605,N_71,N_76);
and U606 (N_606,N_427,N_318);
nand U607 (N_607,N_219,N_183);
or U608 (N_608,N_114,N_226);
and U609 (N_609,N_485,N_366);
nand U610 (N_610,N_476,N_422);
and U611 (N_611,N_396,N_15);
nand U612 (N_612,N_262,N_130);
nor U613 (N_613,N_467,N_386);
and U614 (N_614,N_110,N_27);
nand U615 (N_615,N_247,N_124);
and U616 (N_616,N_270,N_453);
nand U617 (N_617,N_269,N_444);
or U618 (N_618,N_129,N_291);
nor U619 (N_619,N_233,N_339);
or U620 (N_620,N_435,N_348);
and U621 (N_621,N_23,N_469);
and U622 (N_622,N_344,N_29);
and U623 (N_623,N_45,N_7);
nand U624 (N_624,N_399,N_253);
nand U625 (N_625,N_118,N_39);
and U626 (N_626,N_310,N_443);
nor U627 (N_627,N_191,N_131);
and U628 (N_628,N_93,N_231);
xor U629 (N_629,N_43,N_418);
or U630 (N_630,N_198,N_84);
nor U631 (N_631,N_238,N_186);
or U632 (N_632,N_441,N_221);
nand U633 (N_633,N_113,N_217);
or U634 (N_634,N_426,N_159);
nor U635 (N_635,N_458,N_103);
nand U636 (N_636,N_321,N_282);
nor U637 (N_637,N_172,N_448);
nor U638 (N_638,N_67,N_459);
nor U639 (N_639,N_352,N_158);
nand U640 (N_640,N_16,N_287);
nor U641 (N_641,N_357,N_300);
nand U642 (N_642,N_360,N_261);
nand U643 (N_643,N_61,N_431);
or U644 (N_644,N_311,N_215);
nand U645 (N_645,N_224,N_273);
nor U646 (N_646,N_121,N_455);
nor U647 (N_647,N_156,N_388);
nor U648 (N_648,N_86,N_225);
and U649 (N_649,N_51,N_232);
nor U650 (N_650,N_406,N_340);
and U651 (N_651,N_439,N_135);
nand U652 (N_652,N_268,N_354);
or U653 (N_653,N_99,N_266);
nand U654 (N_654,N_494,N_341);
or U655 (N_655,N_144,N_308);
or U656 (N_656,N_58,N_417);
or U657 (N_657,N_218,N_88);
or U658 (N_658,N_383,N_314);
nor U659 (N_659,N_149,N_250);
nand U660 (N_660,N_390,N_41);
or U661 (N_661,N_361,N_196);
nand U662 (N_662,N_209,N_37);
nor U663 (N_663,N_137,N_449);
nand U664 (N_664,N_382,N_47);
or U665 (N_665,N_368,N_350);
nand U666 (N_666,N_381,N_62);
and U667 (N_667,N_35,N_380);
nor U668 (N_668,N_125,N_461);
nor U669 (N_669,N_220,N_446);
nand U670 (N_670,N_286,N_200);
nor U671 (N_671,N_73,N_151);
nand U672 (N_672,N_351,N_210);
nand U673 (N_673,N_452,N_85);
and U674 (N_674,N_49,N_272);
and U675 (N_675,N_486,N_171);
and U676 (N_676,N_346,N_342);
and U677 (N_677,N_134,N_332);
nor U678 (N_678,N_362,N_141);
nand U679 (N_679,N_248,N_428);
nand U680 (N_680,N_90,N_405);
nor U681 (N_681,N_211,N_128);
and U682 (N_682,N_240,N_473);
nor U683 (N_683,N_180,N_28);
nand U684 (N_684,N_460,N_402);
nand U685 (N_685,N_466,N_178);
nand U686 (N_686,N_166,N_246);
and U687 (N_687,N_445,N_203);
nor U688 (N_688,N_489,N_315);
nand U689 (N_689,N_425,N_457);
nor U690 (N_690,N_206,N_106);
and U691 (N_691,N_325,N_440);
or U692 (N_692,N_163,N_256);
and U693 (N_693,N_53,N_108);
and U694 (N_694,N_96,N_483);
and U695 (N_695,N_56,N_44);
or U696 (N_696,N_491,N_488);
nand U697 (N_697,N_264,N_372);
and U698 (N_698,N_482,N_259);
nor U699 (N_699,N_497,N_81);
nand U700 (N_700,N_324,N_492);
xnor U701 (N_701,N_463,N_157);
or U702 (N_702,N_479,N_327);
or U703 (N_703,N_363,N_412);
nand U704 (N_704,N_401,N_155);
nor U705 (N_705,N_437,N_364);
xor U706 (N_706,N_385,N_454);
and U707 (N_707,N_214,N_111);
and U708 (N_708,N_243,N_468);
or U709 (N_709,N_123,N_208);
nand U710 (N_710,N_13,N_60);
nand U711 (N_711,N_46,N_18);
or U712 (N_712,N_162,N_371);
and U713 (N_713,N_164,N_32);
nand U714 (N_714,N_409,N_475);
and U715 (N_715,N_22,N_301);
and U716 (N_716,N_481,N_5);
and U717 (N_717,N_228,N_188);
and U718 (N_718,N_77,N_279);
nor U719 (N_719,N_478,N_192);
nor U720 (N_720,N_66,N_244);
nor U721 (N_721,N_251,N_154);
nor U722 (N_722,N_349,N_260);
nand U723 (N_723,N_379,N_65);
nand U724 (N_724,N_19,N_42);
and U725 (N_725,N_265,N_0);
and U726 (N_726,N_165,N_465);
and U727 (N_727,N_375,N_420);
and U728 (N_728,N_280,N_353);
or U729 (N_729,N_40,N_161);
nand U730 (N_730,N_317,N_423);
nor U731 (N_731,N_239,N_170);
or U732 (N_732,N_429,N_305);
and U733 (N_733,N_336,N_447);
nand U734 (N_734,N_63,N_370);
nor U735 (N_735,N_182,N_442);
nor U736 (N_736,N_306,N_331);
nor U737 (N_737,N_59,N_296);
and U738 (N_738,N_9,N_365);
nor U739 (N_739,N_480,N_356);
nand U740 (N_740,N_276,N_133);
nor U741 (N_741,N_12,N_101);
nand U742 (N_742,N_79,N_72);
nor U743 (N_743,N_241,N_174);
nor U744 (N_744,N_334,N_205);
nor U745 (N_745,N_397,N_229);
nand U746 (N_746,N_313,N_1);
nor U747 (N_747,N_54,N_373);
and U748 (N_748,N_234,N_393);
nor U749 (N_749,N_263,N_102);
or U750 (N_750,N_81,N_480);
and U751 (N_751,N_66,N_21);
and U752 (N_752,N_352,N_247);
and U753 (N_753,N_204,N_306);
nor U754 (N_754,N_442,N_157);
nand U755 (N_755,N_230,N_227);
nor U756 (N_756,N_256,N_413);
or U757 (N_757,N_379,N_181);
nor U758 (N_758,N_149,N_402);
nor U759 (N_759,N_328,N_303);
or U760 (N_760,N_78,N_279);
or U761 (N_761,N_347,N_19);
nand U762 (N_762,N_84,N_95);
and U763 (N_763,N_59,N_217);
and U764 (N_764,N_359,N_169);
nand U765 (N_765,N_135,N_85);
or U766 (N_766,N_450,N_81);
nor U767 (N_767,N_248,N_427);
and U768 (N_768,N_223,N_84);
and U769 (N_769,N_195,N_307);
nand U770 (N_770,N_311,N_431);
nand U771 (N_771,N_106,N_103);
nand U772 (N_772,N_41,N_314);
and U773 (N_773,N_350,N_73);
or U774 (N_774,N_471,N_154);
or U775 (N_775,N_358,N_490);
or U776 (N_776,N_428,N_448);
nand U777 (N_777,N_325,N_308);
and U778 (N_778,N_186,N_442);
or U779 (N_779,N_488,N_183);
and U780 (N_780,N_259,N_186);
nor U781 (N_781,N_78,N_205);
or U782 (N_782,N_464,N_157);
nor U783 (N_783,N_489,N_403);
nand U784 (N_784,N_305,N_21);
and U785 (N_785,N_462,N_391);
or U786 (N_786,N_375,N_437);
or U787 (N_787,N_379,N_474);
or U788 (N_788,N_56,N_117);
nand U789 (N_789,N_348,N_170);
or U790 (N_790,N_18,N_485);
nor U791 (N_791,N_426,N_92);
nor U792 (N_792,N_255,N_301);
nand U793 (N_793,N_92,N_6);
nand U794 (N_794,N_195,N_350);
or U795 (N_795,N_428,N_110);
nor U796 (N_796,N_65,N_327);
nand U797 (N_797,N_5,N_190);
and U798 (N_798,N_440,N_282);
and U799 (N_799,N_466,N_85);
or U800 (N_800,N_227,N_334);
nand U801 (N_801,N_225,N_105);
and U802 (N_802,N_376,N_343);
or U803 (N_803,N_176,N_71);
and U804 (N_804,N_93,N_292);
or U805 (N_805,N_326,N_163);
nand U806 (N_806,N_211,N_493);
nor U807 (N_807,N_227,N_25);
and U808 (N_808,N_33,N_26);
and U809 (N_809,N_295,N_328);
nand U810 (N_810,N_308,N_135);
and U811 (N_811,N_92,N_493);
nor U812 (N_812,N_23,N_293);
nand U813 (N_813,N_24,N_49);
and U814 (N_814,N_178,N_218);
nor U815 (N_815,N_210,N_371);
and U816 (N_816,N_47,N_139);
nand U817 (N_817,N_299,N_387);
nand U818 (N_818,N_357,N_421);
nor U819 (N_819,N_398,N_348);
nor U820 (N_820,N_182,N_282);
nor U821 (N_821,N_127,N_97);
and U822 (N_822,N_7,N_179);
nor U823 (N_823,N_341,N_210);
nand U824 (N_824,N_210,N_228);
and U825 (N_825,N_171,N_397);
and U826 (N_826,N_216,N_173);
nor U827 (N_827,N_110,N_395);
nor U828 (N_828,N_232,N_225);
nor U829 (N_829,N_161,N_274);
and U830 (N_830,N_69,N_446);
and U831 (N_831,N_457,N_489);
and U832 (N_832,N_406,N_46);
and U833 (N_833,N_461,N_361);
and U834 (N_834,N_75,N_94);
and U835 (N_835,N_6,N_328);
or U836 (N_836,N_224,N_20);
or U837 (N_837,N_237,N_472);
nor U838 (N_838,N_245,N_177);
and U839 (N_839,N_420,N_391);
nor U840 (N_840,N_287,N_224);
nor U841 (N_841,N_249,N_451);
or U842 (N_842,N_265,N_248);
and U843 (N_843,N_9,N_363);
and U844 (N_844,N_429,N_53);
and U845 (N_845,N_196,N_37);
and U846 (N_846,N_345,N_411);
nand U847 (N_847,N_27,N_2);
nor U848 (N_848,N_167,N_236);
and U849 (N_849,N_297,N_121);
nand U850 (N_850,N_5,N_239);
nand U851 (N_851,N_298,N_89);
nand U852 (N_852,N_494,N_7);
nor U853 (N_853,N_340,N_161);
nand U854 (N_854,N_411,N_171);
and U855 (N_855,N_485,N_50);
or U856 (N_856,N_273,N_301);
nand U857 (N_857,N_439,N_134);
or U858 (N_858,N_442,N_410);
and U859 (N_859,N_48,N_209);
or U860 (N_860,N_490,N_375);
nor U861 (N_861,N_226,N_281);
or U862 (N_862,N_5,N_142);
nand U863 (N_863,N_489,N_5);
nand U864 (N_864,N_303,N_369);
and U865 (N_865,N_156,N_325);
nor U866 (N_866,N_123,N_57);
and U867 (N_867,N_40,N_167);
and U868 (N_868,N_468,N_184);
nand U869 (N_869,N_441,N_391);
and U870 (N_870,N_343,N_404);
or U871 (N_871,N_425,N_111);
nand U872 (N_872,N_114,N_308);
and U873 (N_873,N_362,N_215);
or U874 (N_874,N_409,N_89);
or U875 (N_875,N_112,N_91);
nand U876 (N_876,N_171,N_430);
nand U877 (N_877,N_247,N_75);
and U878 (N_878,N_246,N_187);
nor U879 (N_879,N_387,N_254);
nand U880 (N_880,N_417,N_47);
or U881 (N_881,N_472,N_61);
nor U882 (N_882,N_47,N_157);
or U883 (N_883,N_318,N_350);
or U884 (N_884,N_240,N_29);
or U885 (N_885,N_153,N_405);
or U886 (N_886,N_166,N_281);
nand U887 (N_887,N_367,N_39);
nor U888 (N_888,N_193,N_39);
nor U889 (N_889,N_119,N_275);
nand U890 (N_890,N_466,N_203);
nor U891 (N_891,N_241,N_159);
or U892 (N_892,N_77,N_378);
or U893 (N_893,N_332,N_187);
or U894 (N_894,N_291,N_57);
and U895 (N_895,N_250,N_239);
and U896 (N_896,N_23,N_489);
or U897 (N_897,N_471,N_463);
or U898 (N_898,N_130,N_100);
and U899 (N_899,N_147,N_432);
or U900 (N_900,N_387,N_105);
and U901 (N_901,N_112,N_312);
nor U902 (N_902,N_436,N_211);
and U903 (N_903,N_53,N_126);
and U904 (N_904,N_123,N_399);
nand U905 (N_905,N_283,N_271);
or U906 (N_906,N_114,N_262);
nor U907 (N_907,N_267,N_475);
nor U908 (N_908,N_139,N_182);
and U909 (N_909,N_358,N_71);
nor U910 (N_910,N_413,N_348);
nor U911 (N_911,N_282,N_207);
nor U912 (N_912,N_319,N_178);
or U913 (N_913,N_416,N_279);
nor U914 (N_914,N_310,N_217);
nand U915 (N_915,N_353,N_46);
nor U916 (N_916,N_89,N_457);
and U917 (N_917,N_10,N_175);
nand U918 (N_918,N_23,N_388);
and U919 (N_919,N_285,N_362);
nand U920 (N_920,N_257,N_74);
nor U921 (N_921,N_163,N_0);
nor U922 (N_922,N_167,N_470);
nor U923 (N_923,N_425,N_166);
nand U924 (N_924,N_251,N_10);
nor U925 (N_925,N_174,N_179);
nor U926 (N_926,N_139,N_364);
and U927 (N_927,N_222,N_55);
nor U928 (N_928,N_283,N_267);
nor U929 (N_929,N_229,N_21);
nand U930 (N_930,N_178,N_226);
or U931 (N_931,N_192,N_51);
nor U932 (N_932,N_295,N_472);
and U933 (N_933,N_340,N_238);
nor U934 (N_934,N_153,N_385);
and U935 (N_935,N_150,N_308);
nand U936 (N_936,N_99,N_405);
and U937 (N_937,N_412,N_457);
nand U938 (N_938,N_405,N_372);
and U939 (N_939,N_259,N_417);
nor U940 (N_940,N_147,N_431);
and U941 (N_941,N_331,N_189);
nand U942 (N_942,N_460,N_395);
or U943 (N_943,N_361,N_303);
or U944 (N_944,N_239,N_235);
or U945 (N_945,N_76,N_362);
nor U946 (N_946,N_156,N_173);
and U947 (N_947,N_256,N_4);
or U948 (N_948,N_327,N_455);
and U949 (N_949,N_151,N_406);
and U950 (N_950,N_166,N_189);
nand U951 (N_951,N_107,N_99);
and U952 (N_952,N_204,N_89);
nand U953 (N_953,N_399,N_186);
and U954 (N_954,N_314,N_130);
nor U955 (N_955,N_119,N_81);
and U956 (N_956,N_118,N_302);
or U957 (N_957,N_320,N_248);
or U958 (N_958,N_125,N_188);
nor U959 (N_959,N_380,N_76);
nor U960 (N_960,N_51,N_362);
or U961 (N_961,N_95,N_163);
nor U962 (N_962,N_423,N_466);
or U963 (N_963,N_52,N_366);
nand U964 (N_964,N_269,N_3);
nand U965 (N_965,N_304,N_72);
and U966 (N_966,N_66,N_123);
or U967 (N_967,N_356,N_198);
and U968 (N_968,N_121,N_167);
or U969 (N_969,N_429,N_33);
nor U970 (N_970,N_288,N_129);
nor U971 (N_971,N_90,N_154);
nand U972 (N_972,N_15,N_151);
or U973 (N_973,N_390,N_59);
nand U974 (N_974,N_302,N_194);
and U975 (N_975,N_16,N_186);
or U976 (N_976,N_90,N_345);
nand U977 (N_977,N_355,N_196);
and U978 (N_978,N_29,N_453);
nor U979 (N_979,N_356,N_316);
nor U980 (N_980,N_449,N_125);
nor U981 (N_981,N_346,N_110);
nor U982 (N_982,N_249,N_125);
or U983 (N_983,N_329,N_436);
nor U984 (N_984,N_214,N_388);
or U985 (N_985,N_95,N_425);
and U986 (N_986,N_152,N_469);
or U987 (N_987,N_282,N_461);
and U988 (N_988,N_96,N_130);
nand U989 (N_989,N_392,N_219);
and U990 (N_990,N_20,N_276);
and U991 (N_991,N_210,N_48);
nor U992 (N_992,N_83,N_13);
or U993 (N_993,N_186,N_329);
and U994 (N_994,N_279,N_256);
and U995 (N_995,N_295,N_344);
nand U996 (N_996,N_490,N_404);
xor U997 (N_997,N_441,N_8);
or U998 (N_998,N_68,N_475);
nand U999 (N_999,N_170,N_326);
nand U1000 (N_1000,N_702,N_543);
nand U1001 (N_1001,N_792,N_859);
and U1002 (N_1002,N_576,N_993);
nor U1003 (N_1003,N_961,N_989);
or U1004 (N_1004,N_670,N_645);
or U1005 (N_1005,N_669,N_967);
or U1006 (N_1006,N_869,N_529);
xnor U1007 (N_1007,N_725,N_506);
and U1008 (N_1008,N_971,N_690);
and U1009 (N_1009,N_912,N_538);
and U1010 (N_1010,N_577,N_819);
or U1011 (N_1011,N_911,N_829);
and U1012 (N_1012,N_635,N_696);
and U1013 (N_1013,N_867,N_977);
or U1014 (N_1014,N_826,N_633);
nor U1015 (N_1015,N_882,N_655);
and U1016 (N_1016,N_668,N_803);
nand U1017 (N_1017,N_515,N_871);
and U1018 (N_1018,N_663,N_774);
and U1019 (N_1019,N_592,N_621);
nor U1020 (N_1020,N_748,N_895);
nor U1021 (N_1021,N_862,N_717);
nand U1022 (N_1022,N_501,N_959);
nand U1023 (N_1023,N_892,N_806);
or U1024 (N_1024,N_901,N_958);
nand U1025 (N_1025,N_606,N_764);
nor U1026 (N_1026,N_990,N_904);
nor U1027 (N_1027,N_540,N_768);
and U1028 (N_1028,N_557,N_916);
nor U1029 (N_1029,N_816,N_639);
or U1030 (N_1030,N_897,N_986);
or U1031 (N_1031,N_523,N_595);
nand U1032 (N_1032,N_842,N_855);
or U1033 (N_1033,N_505,N_646);
and U1034 (N_1034,N_902,N_787);
or U1035 (N_1035,N_783,N_561);
and U1036 (N_1036,N_952,N_599);
nand U1037 (N_1037,N_770,N_628);
nand U1038 (N_1038,N_604,N_714);
and U1039 (N_1039,N_603,N_607);
and U1040 (N_1040,N_512,N_778);
and U1041 (N_1041,N_636,N_907);
or U1042 (N_1042,N_718,N_611);
or U1043 (N_1043,N_522,N_514);
nor U1044 (N_1044,N_638,N_550);
nor U1045 (N_1045,N_531,N_622);
nand U1046 (N_1046,N_831,N_894);
nand U1047 (N_1047,N_558,N_818);
nor U1048 (N_1048,N_874,N_526);
nor U1049 (N_1049,N_572,N_503);
nand U1050 (N_1050,N_728,N_813);
nand U1051 (N_1051,N_692,N_528);
nand U1052 (N_1052,N_846,N_931);
nand U1053 (N_1053,N_652,N_739);
or U1054 (N_1054,N_651,N_548);
nand U1055 (N_1055,N_891,N_566);
and U1056 (N_1056,N_962,N_624);
nor U1057 (N_1057,N_588,N_996);
nand U1058 (N_1058,N_922,N_502);
or U1059 (N_1059,N_972,N_785);
nor U1060 (N_1060,N_811,N_684);
nor U1061 (N_1061,N_755,N_649);
and U1062 (N_1062,N_618,N_913);
or U1063 (N_1063,N_758,N_975);
or U1064 (N_1064,N_847,N_659);
and U1065 (N_1065,N_613,N_845);
nand U1066 (N_1066,N_637,N_695);
nor U1067 (N_1067,N_948,N_941);
or U1068 (N_1068,N_798,N_693);
nand U1069 (N_1069,N_769,N_940);
nand U1070 (N_1070,N_982,N_697);
nand U1071 (N_1071,N_954,N_620);
and U1072 (N_1072,N_598,N_716);
or U1073 (N_1073,N_736,N_957);
or U1074 (N_1074,N_662,N_753);
and U1075 (N_1075,N_915,N_925);
or U1076 (N_1076,N_590,N_623);
nor U1077 (N_1077,N_887,N_699);
nor U1078 (N_1078,N_995,N_625);
or U1079 (N_1079,N_927,N_614);
nand U1080 (N_1080,N_876,N_596);
nor U1081 (N_1081,N_556,N_641);
or U1082 (N_1082,N_609,N_861);
or U1083 (N_1083,N_804,N_893);
or U1084 (N_1084,N_738,N_926);
nand U1085 (N_1085,N_551,N_744);
nor U1086 (N_1086,N_541,N_726);
nand U1087 (N_1087,N_994,N_791);
or U1088 (N_1088,N_704,N_667);
or U1089 (N_1089,N_732,N_762);
or U1090 (N_1090,N_851,N_708);
nand U1091 (N_1091,N_909,N_838);
and U1092 (N_1092,N_722,N_681);
and U1093 (N_1093,N_835,N_767);
xor U1094 (N_1094,N_568,N_873);
nand U1095 (N_1095,N_733,N_786);
nor U1096 (N_1096,N_661,N_581);
nor U1097 (N_1097,N_875,N_780);
or U1098 (N_1098,N_878,N_741);
nor U1099 (N_1099,N_565,N_809);
nor U1100 (N_1100,N_886,N_700);
nand U1101 (N_1101,N_573,N_689);
or U1102 (N_1102,N_510,N_934);
or U1103 (N_1103,N_965,N_602);
and U1104 (N_1104,N_881,N_998);
nor U1105 (N_1105,N_898,N_850);
or U1106 (N_1106,N_937,N_766);
xor U1107 (N_1107,N_953,N_589);
nand U1108 (N_1108,N_919,N_761);
nand U1109 (N_1109,N_719,N_591);
or U1110 (N_1110,N_923,N_519);
or U1111 (N_1111,N_802,N_539);
nand U1112 (N_1112,N_720,N_513);
nand U1113 (N_1113,N_585,N_883);
nand U1114 (N_1114,N_735,N_688);
and U1115 (N_1115,N_924,N_676);
nor U1116 (N_1116,N_933,N_921);
nor U1117 (N_1117,N_644,N_509);
nor U1118 (N_1118,N_932,N_777);
nand U1119 (N_1119,N_698,N_547);
nand U1120 (N_1120,N_964,N_563);
and U1121 (N_1121,N_530,N_711);
nor U1122 (N_1122,N_782,N_908);
or U1123 (N_1123,N_605,N_760);
or U1124 (N_1124,N_889,N_945);
nor U1125 (N_1125,N_827,N_794);
nor U1126 (N_1126,N_640,N_685);
or U1127 (N_1127,N_671,N_910);
nor U1128 (N_1128,N_852,N_991);
nand U1129 (N_1129,N_552,N_853);
nor U1130 (N_1130,N_920,N_918);
nor U1131 (N_1131,N_928,N_799);
nor U1132 (N_1132,N_935,N_631);
nand U1133 (N_1133,N_678,N_749);
and U1134 (N_1134,N_537,N_772);
nand U1135 (N_1135,N_517,N_946);
nor U1136 (N_1136,N_754,N_675);
and U1137 (N_1137,N_981,N_617);
or U1138 (N_1138,N_694,N_658);
nor U1139 (N_1139,N_858,N_788);
nor U1140 (N_1140,N_992,N_983);
or U1141 (N_1141,N_656,N_860);
nor U1142 (N_1142,N_820,N_864);
nand U1143 (N_1143,N_507,N_730);
and U1144 (N_1144,N_943,N_843);
and U1145 (N_1145,N_709,N_665);
nand U1146 (N_1146,N_840,N_721);
and U1147 (N_1147,N_610,N_579);
nor U1148 (N_1148,N_757,N_527);
or U1149 (N_1149,N_564,N_608);
or U1150 (N_1150,N_976,N_747);
or U1151 (N_1151,N_936,N_666);
or U1152 (N_1152,N_823,N_980);
xnor U1153 (N_1153,N_546,N_734);
or U1154 (N_1154,N_906,N_657);
nor U1155 (N_1155,N_955,N_844);
nand U1156 (N_1156,N_900,N_963);
or U1157 (N_1157,N_567,N_533);
or U1158 (N_1158,N_839,N_830);
nand U1159 (N_1159,N_516,N_751);
nand U1160 (N_1160,N_880,N_903);
nor U1161 (N_1161,N_575,N_879);
or U1162 (N_1162,N_808,N_797);
or U1163 (N_1163,N_759,N_524);
or U1164 (N_1164,N_706,N_834);
or U1165 (N_1165,N_703,N_594);
nor U1166 (N_1166,N_745,N_687);
nand U1167 (N_1167,N_781,N_868);
and U1168 (N_1168,N_817,N_586);
xnor U1169 (N_1169,N_511,N_815);
nor U1170 (N_1170,N_833,N_544);
or U1171 (N_1171,N_885,N_612);
or U1172 (N_1172,N_653,N_899);
or U1173 (N_1173,N_984,N_956);
or U1174 (N_1174,N_500,N_997);
or U1175 (N_1175,N_619,N_508);
nor U1176 (N_1176,N_583,N_518);
or U1177 (N_1177,N_571,N_947);
nor U1178 (N_1178,N_789,N_584);
nor U1179 (N_1179,N_627,N_828);
and U1180 (N_1180,N_740,N_987);
nand U1181 (N_1181,N_715,N_731);
nor U1182 (N_1182,N_863,N_822);
or U1183 (N_1183,N_950,N_939);
nand U1184 (N_1184,N_999,N_705);
or U1185 (N_1185,N_532,N_870);
nand U1186 (N_1186,N_836,N_679);
nor U1187 (N_1187,N_857,N_710);
nand U1188 (N_1188,N_807,N_535);
nor U1189 (N_1189,N_872,N_654);
or U1190 (N_1190,N_773,N_629);
or U1191 (N_1191,N_888,N_854);
or U1192 (N_1192,N_877,N_542);
and U1193 (N_1193,N_865,N_812);
nor U1194 (N_1194,N_553,N_691);
nor U1195 (N_1195,N_974,N_559);
nor U1196 (N_1196,N_848,N_580);
and U1197 (N_1197,N_555,N_856);
and U1198 (N_1198,N_793,N_930);
nand U1199 (N_1199,N_712,N_632);
xor U1200 (N_1200,N_779,N_832);
or U1201 (N_1201,N_536,N_988);
nand U1202 (N_1202,N_884,N_985);
or U1203 (N_1203,N_944,N_682);
nor U1204 (N_1204,N_578,N_680);
and U1205 (N_1205,N_549,N_771);
nand U1206 (N_1206,N_801,N_570);
and U1207 (N_1207,N_756,N_562);
nor U1208 (N_1208,N_973,N_713);
and U1209 (N_1209,N_587,N_765);
nor U1210 (N_1210,N_582,N_866);
nor U1211 (N_1211,N_784,N_978);
or U1212 (N_1212,N_890,N_742);
and U1213 (N_1213,N_821,N_724);
nand U1214 (N_1214,N_660,N_960);
or U1215 (N_1215,N_616,N_743);
and U1216 (N_1216,N_630,N_634);
nor U1217 (N_1217,N_574,N_942);
nor U1218 (N_1218,N_917,N_569);
nand U1219 (N_1219,N_929,N_648);
nand U1220 (N_1220,N_729,N_746);
nand U1221 (N_1221,N_825,N_969);
nand U1222 (N_1222,N_914,N_800);
or U1223 (N_1223,N_642,N_723);
and U1224 (N_1224,N_905,N_970);
or U1225 (N_1225,N_534,N_968);
nor U1226 (N_1226,N_979,N_615);
and U1227 (N_1227,N_677,N_643);
or U1228 (N_1228,N_837,N_790);
xnor U1229 (N_1229,N_707,N_966);
or U1230 (N_1230,N_737,N_664);
or U1231 (N_1231,N_949,N_849);
and U1232 (N_1232,N_686,N_683);
nand U1233 (N_1233,N_701,N_597);
or U1234 (N_1234,N_727,N_841);
nor U1235 (N_1235,N_896,N_795);
and U1236 (N_1236,N_814,N_951);
and U1237 (N_1237,N_520,N_824);
and U1238 (N_1238,N_750,N_545);
nor U1239 (N_1239,N_796,N_504);
and U1240 (N_1240,N_560,N_805);
or U1241 (N_1241,N_593,N_938);
or U1242 (N_1242,N_672,N_601);
xor U1243 (N_1243,N_776,N_650);
nand U1244 (N_1244,N_600,N_673);
nand U1245 (N_1245,N_810,N_752);
nor U1246 (N_1246,N_763,N_554);
and U1247 (N_1247,N_674,N_647);
nor U1248 (N_1248,N_521,N_626);
or U1249 (N_1249,N_775,N_525);
nor U1250 (N_1250,N_907,N_675);
and U1251 (N_1251,N_908,N_791);
nor U1252 (N_1252,N_549,N_506);
nand U1253 (N_1253,N_772,N_942);
or U1254 (N_1254,N_650,N_644);
nand U1255 (N_1255,N_979,N_983);
nand U1256 (N_1256,N_867,N_964);
or U1257 (N_1257,N_929,N_565);
and U1258 (N_1258,N_741,N_633);
and U1259 (N_1259,N_723,N_777);
nor U1260 (N_1260,N_962,N_976);
or U1261 (N_1261,N_731,N_908);
nor U1262 (N_1262,N_720,N_504);
nand U1263 (N_1263,N_830,N_688);
nor U1264 (N_1264,N_891,N_843);
or U1265 (N_1265,N_850,N_981);
nand U1266 (N_1266,N_647,N_524);
nand U1267 (N_1267,N_925,N_710);
or U1268 (N_1268,N_905,N_922);
nand U1269 (N_1269,N_535,N_924);
nor U1270 (N_1270,N_951,N_907);
and U1271 (N_1271,N_844,N_530);
nand U1272 (N_1272,N_809,N_581);
nor U1273 (N_1273,N_785,N_738);
or U1274 (N_1274,N_612,N_593);
or U1275 (N_1275,N_724,N_937);
and U1276 (N_1276,N_672,N_972);
nand U1277 (N_1277,N_873,N_737);
xnor U1278 (N_1278,N_617,N_777);
nand U1279 (N_1279,N_567,N_780);
nand U1280 (N_1280,N_666,N_657);
and U1281 (N_1281,N_564,N_755);
nor U1282 (N_1282,N_635,N_629);
and U1283 (N_1283,N_919,N_548);
nor U1284 (N_1284,N_742,N_760);
nand U1285 (N_1285,N_948,N_759);
or U1286 (N_1286,N_916,N_707);
nand U1287 (N_1287,N_713,N_505);
or U1288 (N_1288,N_563,N_858);
nand U1289 (N_1289,N_746,N_534);
or U1290 (N_1290,N_930,N_863);
or U1291 (N_1291,N_906,N_815);
and U1292 (N_1292,N_994,N_665);
nand U1293 (N_1293,N_814,N_610);
nand U1294 (N_1294,N_913,N_577);
and U1295 (N_1295,N_838,N_610);
nor U1296 (N_1296,N_990,N_697);
or U1297 (N_1297,N_887,N_774);
or U1298 (N_1298,N_906,N_879);
or U1299 (N_1299,N_780,N_502);
nor U1300 (N_1300,N_708,N_516);
and U1301 (N_1301,N_822,N_657);
nor U1302 (N_1302,N_529,N_826);
or U1303 (N_1303,N_744,N_910);
nand U1304 (N_1304,N_863,N_887);
or U1305 (N_1305,N_963,N_594);
or U1306 (N_1306,N_536,N_646);
nand U1307 (N_1307,N_803,N_674);
nor U1308 (N_1308,N_912,N_616);
nor U1309 (N_1309,N_673,N_584);
or U1310 (N_1310,N_975,N_649);
or U1311 (N_1311,N_530,N_818);
and U1312 (N_1312,N_745,N_781);
or U1313 (N_1313,N_632,N_560);
and U1314 (N_1314,N_698,N_578);
nor U1315 (N_1315,N_847,N_915);
and U1316 (N_1316,N_683,N_736);
or U1317 (N_1317,N_891,N_705);
nor U1318 (N_1318,N_599,N_640);
nand U1319 (N_1319,N_700,N_575);
or U1320 (N_1320,N_664,N_713);
and U1321 (N_1321,N_564,N_815);
or U1322 (N_1322,N_774,N_920);
nand U1323 (N_1323,N_533,N_760);
nor U1324 (N_1324,N_951,N_975);
or U1325 (N_1325,N_956,N_830);
nor U1326 (N_1326,N_982,N_602);
or U1327 (N_1327,N_682,N_587);
nor U1328 (N_1328,N_507,N_686);
nor U1329 (N_1329,N_904,N_891);
nor U1330 (N_1330,N_561,N_911);
nand U1331 (N_1331,N_958,N_776);
and U1332 (N_1332,N_516,N_611);
nand U1333 (N_1333,N_929,N_895);
or U1334 (N_1334,N_791,N_817);
nor U1335 (N_1335,N_673,N_755);
nor U1336 (N_1336,N_917,N_942);
or U1337 (N_1337,N_843,N_530);
nor U1338 (N_1338,N_627,N_646);
and U1339 (N_1339,N_698,N_507);
nor U1340 (N_1340,N_765,N_549);
or U1341 (N_1341,N_779,N_606);
nor U1342 (N_1342,N_850,N_864);
and U1343 (N_1343,N_980,N_615);
nor U1344 (N_1344,N_769,N_689);
and U1345 (N_1345,N_600,N_564);
and U1346 (N_1346,N_800,N_582);
or U1347 (N_1347,N_547,N_609);
or U1348 (N_1348,N_661,N_844);
or U1349 (N_1349,N_931,N_691);
or U1350 (N_1350,N_633,N_976);
or U1351 (N_1351,N_922,N_562);
nor U1352 (N_1352,N_765,N_537);
nand U1353 (N_1353,N_634,N_757);
nor U1354 (N_1354,N_864,N_872);
or U1355 (N_1355,N_861,N_741);
nand U1356 (N_1356,N_859,N_786);
nor U1357 (N_1357,N_958,N_855);
or U1358 (N_1358,N_542,N_731);
and U1359 (N_1359,N_571,N_853);
nor U1360 (N_1360,N_574,N_756);
nand U1361 (N_1361,N_610,N_620);
nand U1362 (N_1362,N_987,N_884);
nor U1363 (N_1363,N_685,N_655);
and U1364 (N_1364,N_833,N_545);
nor U1365 (N_1365,N_876,N_577);
or U1366 (N_1366,N_690,N_965);
and U1367 (N_1367,N_895,N_922);
or U1368 (N_1368,N_908,N_995);
and U1369 (N_1369,N_629,N_520);
nor U1370 (N_1370,N_554,N_690);
nor U1371 (N_1371,N_869,N_985);
or U1372 (N_1372,N_936,N_591);
nor U1373 (N_1373,N_813,N_602);
nor U1374 (N_1374,N_814,N_716);
nand U1375 (N_1375,N_707,N_676);
nand U1376 (N_1376,N_948,N_937);
nor U1377 (N_1377,N_833,N_977);
nand U1378 (N_1378,N_731,N_957);
and U1379 (N_1379,N_525,N_994);
and U1380 (N_1380,N_893,N_903);
nand U1381 (N_1381,N_727,N_708);
and U1382 (N_1382,N_941,N_515);
nor U1383 (N_1383,N_879,N_672);
or U1384 (N_1384,N_840,N_741);
and U1385 (N_1385,N_519,N_836);
and U1386 (N_1386,N_524,N_574);
nand U1387 (N_1387,N_836,N_999);
nand U1388 (N_1388,N_654,N_967);
or U1389 (N_1389,N_706,N_841);
and U1390 (N_1390,N_609,N_863);
or U1391 (N_1391,N_614,N_693);
and U1392 (N_1392,N_508,N_609);
or U1393 (N_1393,N_893,N_644);
nor U1394 (N_1394,N_504,N_753);
or U1395 (N_1395,N_819,N_933);
or U1396 (N_1396,N_764,N_797);
nor U1397 (N_1397,N_929,N_826);
nand U1398 (N_1398,N_978,N_757);
nand U1399 (N_1399,N_828,N_585);
nor U1400 (N_1400,N_529,N_805);
or U1401 (N_1401,N_699,N_621);
nor U1402 (N_1402,N_539,N_875);
nand U1403 (N_1403,N_847,N_592);
nor U1404 (N_1404,N_774,N_839);
nor U1405 (N_1405,N_905,N_982);
or U1406 (N_1406,N_517,N_799);
nor U1407 (N_1407,N_743,N_593);
and U1408 (N_1408,N_714,N_902);
and U1409 (N_1409,N_709,N_588);
nand U1410 (N_1410,N_648,N_677);
and U1411 (N_1411,N_563,N_703);
nor U1412 (N_1412,N_805,N_956);
and U1413 (N_1413,N_911,N_598);
nor U1414 (N_1414,N_987,N_599);
or U1415 (N_1415,N_815,N_637);
or U1416 (N_1416,N_869,N_691);
or U1417 (N_1417,N_796,N_974);
nor U1418 (N_1418,N_751,N_589);
nor U1419 (N_1419,N_872,N_531);
or U1420 (N_1420,N_985,N_909);
or U1421 (N_1421,N_507,N_575);
nor U1422 (N_1422,N_665,N_576);
nand U1423 (N_1423,N_585,N_542);
or U1424 (N_1424,N_873,N_933);
nand U1425 (N_1425,N_600,N_684);
and U1426 (N_1426,N_684,N_858);
nor U1427 (N_1427,N_864,N_785);
and U1428 (N_1428,N_652,N_767);
and U1429 (N_1429,N_951,N_891);
nor U1430 (N_1430,N_917,N_975);
nor U1431 (N_1431,N_858,N_680);
and U1432 (N_1432,N_842,N_882);
nor U1433 (N_1433,N_999,N_915);
nand U1434 (N_1434,N_530,N_583);
and U1435 (N_1435,N_983,N_546);
nand U1436 (N_1436,N_505,N_884);
and U1437 (N_1437,N_663,N_821);
nand U1438 (N_1438,N_638,N_869);
or U1439 (N_1439,N_595,N_978);
and U1440 (N_1440,N_835,N_754);
nand U1441 (N_1441,N_552,N_681);
and U1442 (N_1442,N_532,N_777);
or U1443 (N_1443,N_957,N_826);
or U1444 (N_1444,N_921,N_703);
nor U1445 (N_1445,N_540,N_681);
nor U1446 (N_1446,N_854,N_760);
nor U1447 (N_1447,N_787,N_954);
or U1448 (N_1448,N_891,N_940);
and U1449 (N_1449,N_827,N_577);
nand U1450 (N_1450,N_842,N_553);
and U1451 (N_1451,N_605,N_767);
nor U1452 (N_1452,N_944,N_824);
or U1453 (N_1453,N_503,N_606);
nand U1454 (N_1454,N_634,N_719);
or U1455 (N_1455,N_869,N_635);
nor U1456 (N_1456,N_982,N_961);
and U1457 (N_1457,N_796,N_526);
or U1458 (N_1458,N_955,N_670);
nor U1459 (N_1459,N_675,N_965);
nand U1460 (N_1460,N_864,N_570);
nand U1461 (N_1461,N_698,N_920);
nor U1462 (N_1462,N_822,N_903);
or U1463 (N_1463,N_890,N_886);
nand U1464 (N_1464,N_706,N_700);
xnor U1465 (N_1465,N_693,N_820);
and U1466 (N_1466,N_943,N_748);
nand U1467 (N_1467,N_815,N_862);
and U1468 (N_1468,N_592,N_657);
nand U1469 (N_1469,N_812,N_984);
and U1470 (N_1470,N_949,N_581);
nor U1471 (N_1471,N_545,N_534);
and U1472 (N_1472,N_504,N_553);
nand U1473 (N_1473,N_537,N_900);
nand U1474 (N_1474,N_949,N_667);
nand U1475 (N_1475,N_545,N_967);
nand U1476 (N_1476,N_637,N_769);
and U1477 (N_1477,N_611,N_777);
nand U1478 (N_1478,N_579,N_895);
and U1479 (N_1479,N_755,N_550);
or U1480 (N_1480,N_806,N_783);
nor U1481 (N_1481,N_709,N_862);
nor U1482 (N_1482,N_715,N_668);
nand U1483 (N_1483,N_719,N_844);
nand U1484 (N_1484,N_648,N_573);
nand U1485 (N_1485,N_923,N_998);
and U1486 (N_1486,N_621,N_862);
nand U1487 (N_1487,N_878,N_854);
nand U1488 (N_1488,N_598,N_736);
nand U1489 (N_1489,N_827,N_563);
nor U1490 (N_1490,N_672,N_565);
or U1491 (N_1491,N_518,N_579);
and U1492 (N_1492,N_601,N_965);
nor U1493 (N_1493,N_626,N_869);
nor U1494 (N_1494,N_500,N_894);
or U1495 (N_1495,N_565,N_521);
or U1496 (N_1496,N_576,N_669);
nand U1497 (N_1497,N_768,N_650);
and U1498 (N_1498,N_531,N_845);
nor U1499 (N_1499,N_994,N_870);
nor U1500 (N_1500,N_1285,N_1092);
nor U1501 (N_1501,N_1404,N_1495);
nand U1502 (N_1502,N_1327,N_1170);
and U1503 (N_1503,N_1376,N_1298);
nor U1504 (N_1504,N_1009,N_1146);
nor U1505 (N_1505,N_1482,N_1111);
or U1506 (N_1506,N_1183,N_1228);
or U1507 (N_1507,N_1022,N_1154);
or U1508 (N_1508,N_1319,N_1302);
nand U1509 (N_1509,N_1441,N_1421);
nand U1510 (N_1510,N_1379,N_1165);
and U1511 (N_1511,N_1270,N_1024);
and U1512 (N_1512,N_1335,N_1210);
nand U1513 (N_1513,N_1093,N_1251);
and U1514 (N_1514,N_1247,N_1004);
nor U1515 (N_1515,N_1095,N_1209);
nand U1516 (N_1516,N_1366,N_1365);
or U1517 (N_1517,N_1063,N_1011);
nor U1518 (N_1518,N_1419,N_1296);
and U1519 (N_1519,N_1345,N_1295);
and U1520 (N_1520,N_1412,N_1467);
and U1521 (N_1521,N_1294,N_1279);
nand U1522 (N_1522,N_1289,N_1081);
and U1523 (N_1523,N_1307,N_1152);
and U1524 (N_1524,N_1336,N_1357);
nand U1525 (N_1525,N_1292,N_1189);
nand U1526 (N_1526,N_1089,N_1044);
or U1527 (N_1527,N_1072,N_1498);
or U1528 (N_1528,N_1206,N_1016);
nand U1529 (N_1529,N_1389,N_1130);
nand U1530 (N_1530,N_1108,N_1394);
and U1531 (N_1531,N_1264,N_1329);
nor U1532 (N_1532,N_1242,N_1418);
or U1533 (N_1533,N_1179,N_1401);
nand U1534 (N_1534,N_1400,N_1036);
or U1535 (N_1535,N_1184,N_1139);
nor U1536 (N_1536,N_1017,N_1299);
nor U1537 (N_1537,N_1356,N_1040);
nand U1538 (N_1538,N_1133,N_1315);
or U1539 (N_1539,N_1118,N_1432);
and U1540 (N_1540,N_1191,N_1196);
and U1541 (N_1541,N_1186,N_1002);
nor U1542 (N_1542,N_1159,N_1455);
and U1543 (N_1543,N_1318,N_1180);
or U1544 (N_1544,N_1403,N_1476);
and U1545 (N_1545,N_1045,N_1144);
and U1546 (N_1546,N_1042,N_1230);
nor U1547 (N_1547,N_1381,N_1190);
nand U1548 (N_1548,N_1123,N_1488);
or U1549 (N_1549,N_1034,N_1140);
nand U1550 (N_1550,N_1005,N_1491);
xor U1551 (N_1551,N_1342,N_1128);
nand U1552 (N_1552,N_1220,N_1258);
nand U1553 (N_1553,N_1200,N_1372);
and U1554 (N_1554,N_1428,N_1126);
or U1555 (N_1555,N_1167,N_1338);
nor U1556 (N_1556,N_1271,N_1399);
nand U1557 (N_1557,N_1217,N_1424);
or U1558 (N_1558,N_1352,N_1173);
nor U1559 (N_1559,N_1290,N_1347);
nor U1560 (N_1560,N_1127,N_1323);
nor U1561 (N_1561,N_1354,N_1281);
or U1562 (N_1562,N_1324,N_1348);
nor U1563 (N_1563,N_1208,N_1020);
nor U1564 (N_1564,N_1331,N_1231);
nor U1565 (N_1565,N_1332,N_1142);
or U1566 (N_1566,N_1253,N_1479);
nand U1567 (N_1567,N_1411,N_1023);
nor U1568 (N_1568,N_1246,N_1070);
nor U1569 (N_1569,N_1109,N_1141);
nor U1570 (N_1570,N_1280,N_1459);
and U1571 (N_1571,N_1326,N_1098);
and U1572 (N_1572,N_1143,N_1273);
and U1573 (N_1573,N_1337,N_1090);
or U1574 (N_1574,N_1346,N_1069);
and U1575 (N_1575,N_1349,N_1333);
or U1576 (N_1576,N_1041,N_1188);
and U1577 (N_1577,N_1057,N_1019);
nor U1578 (N_1578,N_1388,N_1390);
nand U1579 (N_1579,N_1135,N_1368);
nor U1580 (N_1580,N_1275,N_1132);
xor U1581 (N_1581,N_1313,N_1344);
nand U1582 (N_1582,N_1480,N_1074);
nor U1583 (N_1583,N_1218,N_1269);
and U1584 (N_1584,N_1107,N_1169);
or U1585 (N_1585,N_1028,N_1465);
nor U1586 (N_1586,N_1448,N_1305);
and U1587 (N_1587,N_1048,N_1484);
nor U1588 (N_1588,N_1182,N_1216);
nor U1589 (N_1589,N_1075,N_1151);
nand U1590 (N_1590,N_1496,N_1406);
or U1591 (N_1591,N_1021,N_1248);
or U1592 (N_1592,N_1413,N_1393);
nand U1593 (N_1593,N_1014,N_1160);
or U1594 (N_1594,N_1261,N_1447);
or U1595 (N_1595,N_1314,N_1158);
and U1596 (N_1596,N_1065,N_1157);
nand U1597 (N_1597,N_1362,N_1079);
nor U1598 (N_1598,N_1262,N_1436);
or U1599 (N_1599,N_1047,N_1461);
and U1600 (N_1600,N_1174,N_1266);
nor U1601 (N_1601,N_1103,N_1457);
and U1602 (N_1602,N_1168,N_1468);
and U1603 (N_1603,N_1355,N_1437);
nand U1604 (N_1604,N_1172,N_1256);
nand U1605 (N_1605,N_1229,N_1369);
or U1606 (N_1606,N_1238,N_1147);
nand U1607 (N_1607,N_1440,N_1083);
and U1608 (N_1608,N_1101,N_1297);
nor U1609 (N_1609,N_1472,N_1375);
nor U1610 (N_1610,N_1477,N_1417);
or U1611 (N_1611,N_1010,N_1061);
or U1612 (N_1612,N_1257,N_1115);
and U1613 (N_1613,N_1078,N_1199);
and U1614 (N_1614,N_1304,N_1100);
or U1615 (N_1615,N_1192,N_1420);
or U1616 (N_1616,N_1322,N_1265);
or U1617 (N_1617,N_1385,N_1384);
or U1618 (N_1618,N_1463,N_1032);
and U1619 (N_1619,N_1125,N_1122);
nand U1620 (N_1620,N_1058,N_1303);
nand U1621 (N_1621,N_1250,N_1177);
or U1622 (N_1622,N_1382,N_1232);
nor U1623 (N_1623,N_1148,N_1263);
nor U1624 (N_1624,N_1233,N_1489);
nor U1625 (N_1625,N_1052,N_1490);
nand U1626 (N_1626,N_1360,N_1031);
or U1627 (N_1627,N_1202,N_1235);
and U1628 (N_1628,N_1328,N_1056);
nand U1629 (N_1629,N_1306,N_1176);
or U1630 (N_1630,N_1452,N_1236);
or U1631 (N_1631,N_1062,N_1082);
nand U1632 (N_1632,N_1293,N_1300);
and U1633 (N_1633,N_1311,N_1071);
nand U1634 (N_1634,N_1383,N_1097);
nand U1635 (N_1635,N_1155,N_1156);
nor U1636 (N_1636,N_1254,N_1214);
nand U1637 (N_1637,N_1013,N_1112);
or U1638 (N_1638,N_1361,N_1429);
and U1639 (N_1639,N_1374,N_1096);
and U1640 (N_1640,N_1007,N_1053);
and U1641 (N_1641,N_1149,N_1037);
or U1642 (N_1642,N_1325,N_1162);
nor U1643 (N_1643,N_1185,N_1066);
nor U1644 (N_1644,N_1046,N_1422);
nor U1645 (N_1645,N_1334,N_1012);
and U1646 (N_1646,N_1282,N_1198);
or U1647 (N_1647,N_1391,N_1138);
or U1648 (N_1648,N_1226,N_1284);
nor U1649 (N_1649,N_1387,N_1317);
or U1650 (N_1650,N_1478,N_1094);
or U1651 (N_1651,N_1105,N_1060);
and U1652 (N_1652,N_1438,N_1493);
or U1653 (N_1653,N_1102,N_1373);
or U1654 (N_1654,N_1030,N_1224);
and U1655 (N_1655,N_1458,N_1405);
nand U1656 (N_1656,N_1131,N_1163);
nand U1657 (N_1657,N_1470,N_1129);
and U1658 (N_1658,N_1364,N_1240);
nand U1659 (N_1659,N_1464,N_1410);
nand U1660 (N_1660,N_1055,N_1225);
or U1661 (N_1661,N_1310,N_1178);
nor U1662 (N_1662,N_1085,N_1194);
nand U1663 (N_1663,N_1309,N_1219);
and U1664 (N_1664,N_1234,N_1260);
or U1665 (N_1665,N_1175,N_1187);
and U1666 (N_1666,N_1466,N_1475);
and U1667 (N_1667,N_1207,N_1088);
nand U1668 (N_1668,N_1245,N_1205);
and U1669 (N_1669,N_1409,N_1025);
nor U1670 (N_1670,N_1408,N_1227);
nand U1671 (N_1671,N_1378,N_1171);
and U1672 (N_1672,N_1425,N_1018);
or U1673 (N_1673,N_1116,N_1396);
or U1674 (N_1674,N_1287,N_1267);
or U1675 (N_1675,N_1320,N_1445);
nor U1676 (N_1676,N_1039,N_1215);
nand U1677 (N_1677,N_1166,N_1439);
nor U1678 (N_1678,N_1099,N_1255);
nor U1679 (N_1679,N_1164,N_1276);
and U1680 (N_1680,N_1402,N_1145);
nor U1681 (N_1681,N_1259,N_1221);
and U1682 (N_1682,N_1433,N_1414);
nor U1683 (N_1683,N_1456,N_1239);
or U1684 (N_1684,N_1029,N_1443);
nand U1685 (N_1685,N_1435,N_1080);
nor U1686 (N_1686,N_1150,N_1343);
or U1687 (N_1687,N_1134,N_1213);
nor U1688 (N_1688,N_1211,N_1444);
and U1689 (N_1689,N_1043,N_1054);
nor U1690 (N_1690,N_1446,N_1237);
nor U1691 (N_1691,N_1084,N_1120);
nand U1692 (N_1692,N_1241,N_1434);
or U1693 (N_1693,N_1137,N_1398);
nand U1694 (N_1694,N_1487,N_1450);
nand U1695 (N_1695,N_1492,N_1380);
or U1696 (N_1696,N_1386,N_1283);
and U1697 (N_1697,N_1316,N_1462);
nand U1698 (N_1698,N_1153,N_1113);
nand U1699 (N_1699,N_1124,N_1330);
nor U1700 (N_1700,N_1119,N_1026);
or U1701 (N_1701,N_1321,N_1415);
nor U1702 (N_1702,N_1181,N_1268);
nand U1703 (N_1703,N_1367,N_1272);
and U1704 (N_1704,N_1033,N_1243);
and U1705 (N_1705,N_1474,N_1106);
or U1706 (N_1706,N_1370,N_1006);
nand U1707 (N_1707,N_1000,N_1486);
nor U1708 (N_1708,N_1121,N_1288);
and U1709 (N_1709,N_1201,N_1442);
or U1710 (N_1710,N_1301,N_1104);
nand U1711 (N_1711,N_1204,N_1223);
or U1712 (N_1712,N_1453,N_1049);
and U1713 (N_1713,N_1073,N_1001);
nor U1714 (N_1714,N_1312,N_1067);
or U1715 (N_1715,N_1091,N_1449);
nor U1716 (N_1716,N_1212,N_1471);
and U1717 (N_1717,N_1249,N_1483);
or U1718 (N_1718,N_1340,N_1497);
and U1719 (N_1719,N_1371,N_1499);
nor U1720 (N_1720,N_1423,N_1114);
and U1721 (N_1721,N_1222,N_1278);
nand U1722 (N_1722,N_1451,N_1274);
or U1723 (N_1723,N_1161,N_1117);
or U1724 (N_1724,N_1460,N_1363);
or U1725 (N_1725,N_1392,N_1350);
and U1726 (N_1726,N_1416,N_1469);
or U1727 (N_1727,N_1252,N_1038);
or U1728 (N_1728,N_1473,N_1485);
nor U1729 (N_1729,N_1397,N_1203);
nor U1730 (N_1730,N_1426,N_1430);
nand U1731 (N_1731,N_1351,N_1064);
and U1732 (N_1732,N_1286,N_1087);
or U1733 (N_1733,N_1431,N_1077);
or U1734 (N_1734,N_1377,N_1277);
and U1735 (N_1735,N_1197,N_1136);
or U1736 (N_1736,N_1308,N_1051);
or U1737 (N_1737,N_1050,N_1481);
xnor U1738 (N_1738,N_1027,N_1015);
nand U1739 (N_1739,N_1068,N_1059);
nand U1740 (N_1740,N_1086,N_1291);
or U1741 (N_1741,N_1193,N_1494);
nor U1742 (N_1742,N_1358,N_1003);
nand U1743 (N_1743,N_1407,N_1035);
nor U1744 (N_1744,N_1427,N_1339);
and U1745 (N_1745,N_1195,N_1395);
and U1746 (N_1746,N_1353,N_1454);
or U1747 (N_1747,N_1008,N_1076);
and U1748 (N_1748,N_1244,N_1110);
nand U1749 (N_1749,N_1359,N_1341);
or U1750 (N_1750,N_1414,N_1208);
nor U1751 (N_1751,N_1196,N_1285);
nand U1752 (N_1752,N_1337,N_1414);
and U1753 (N_1753,N_1089,N_1457);
and U1754 (N_1754,N_1187,N_1415);
nor U1755 (N_1755,N_1377,N_1030);
nor U1756 (N_1756,N_1244,N_1418);
and U1757 (N_1757,N_1035,N_1181);
and U1758 (N_1758,N_1246,N_1237);
nand U1759 (N_1759,N_1175,N_1107);
and U1760 (N_1760,N_1325,N_1399);
or U1761 (N_1761,N_1319,N_1068);
and U1762 (N_1762,N_1197,N_1480);
and U1763 (N_1763,N_1037,N_1147);
or U1764 (N_1764,N_1481,N_1374);
nor U1765 (N_1765,N_1326,N_1070);
or U1766 (N_1766,N_1492,N_1327);
and U1767 (N_1767,N_1218,N_1133);
xor U1768 (N_1768,N_1063,N_1139);
nand U1769 (N_1769,N_1474,N_1191);
nor U1770 (N_1770,N_1390,N_1242);
and U1771 (N_1771,N_1229,N_1487);
or U1772 (N_1772,N_1189,N_1206);
and U1773 (N_1773,N_1084,N_1271);
nor U1774 (N_1774,N_1284,N_1306);
and U1775 (N_1775,N_1381,N_1302);
and U1776 (N_1776,N_1335,N_1482);
and U1777 (N_1777,N_1113,N_1220);
and U1778 (N_1778,N_1249,N_1335);
nand U1779 (N_1779,N_1096,N_1071);
nand U1780 (N_1780,N_1476,N_1450);
nand U1781 (N_1781,N_1254,N_1422);
and U1782 (N_1782,N_1280,N_1083);
nor U1783 (N_1783,N_1260,N_1303);
and U1784 (N_1784,N_1229,N_1436);
nor U1785 (N_1785,N_1363,N_1091);
and U1786 (N_1786,N_1149,N_1319);
and U1787 (N_1787,N_1180,N_1191);
nand U1788 (N_1788,N_1214,N_1029);
nor U1789 (N_1789,N_1019,N_1402);
nor U1790 (N_1790,N_1058,N_1145);
nand U1791 (N_1791,N_1161,N_1375);
nor U1792 (N_1792,N_1265,N_1077);
nor U1793 (N_1793,N_1462,N_1324);
nor U1794 (N_1794,N_1139,N_1194);
nand U1795 (N_1795,N_1241,N_1336);
nor U1796 (N_1796,N_1276,N_1064);
nand U1797 (N_1797,N_1076,N_1315);
and U1798 (N_1798,N_1141,N_1483);
or U1799 (N_1799,N_1409,N_1097);
or U1800 (N_1800,N_1462,N_1105);
and U1801 (N_1801,N_1049,N_1340);
nand U1802 (N_1802,N_1058,N_1293);
nor U1803 (N_1803,N_1023,N_1107);
nand U1804 (N_1804,N_1041,N_1199);
or U1805 (N_1805,N_1486,N_1084);
nand U1806 (N_1806,N_1371,N_1208);
nor U1807 (N_1807,N_1497,N_1476);
and U1808 (N_1808,N_1293,N_1089);
nand U1809 (N_1809,N_1179,N_1075);
or U1810 (N_1810,N_1353,N_1153);
or U1811 (N_1811,N_1207,N_1467);
nor U1812 (N_1812,N_1271,N_1015);
or U1813 (N_1813,N_1329,N_1151);
and U1814 (N_1814,N_1066,N_1358);
nor U1815 (N_1815,N_1057,N_1116);
nand U1816 (N_1816,N_1256,N_1175);
or U1817 (N_1817,N_1223,N_1124);
nand U1818 (N_1818,N_1158,N_1037);
or U1819 (N_1819,N_1029,N_1445);
or U1820 (N_1820,N_1263,N_1229);
xor U1821 (N_1821,N_1167,N_1180);
nand U1822 (N_1822,N_1211,N_1341);
nand U1823 (N_1823,N_1302,N_1284);
nor U1824 (N_1824,N_1354,N_1041);
or U1825 (N_1825,N_1123,N_1004);
nor U1826 (N_1826,N_1136,N_1293);
nor U1827 (N_1827,N_1003,N_1497);
nor U1828 (N_1828,N_1376,N_1332);
nand U1829 (N_1829,N_1407,N_1006);
or U1830 (N_1830,N_1264,N_1144);
nand U1831 (N_1831,N_1325,N_1465);
nand U1832 (N_1832,N_1464,N_1319);
and U1833 (N_1833,N_1418,N_1073);
or U1834 (N_1834,N_1373,N_1439);
and U1835 (N_1835,N_1244,N_1162);
nor U1836 (N_1836,N_1491,N_1201);
and U1837 (N_1837,N_1127,N_1376);
nand U1838 (N_1838,N_1087,N_1274);
nand U1839 (N_1839,N_1117,N_1184);
or U1840 (N_1840,N_1006,N_1046);
nand U1841 (N_1841,N_1177,N_1240);
or U1842 (N_1842,N_1061,N_1331);
nor U1843 (N_1843,N_1202,N_1497);
xnor U1844 (N_1844,N_1056,N_1290);
and U1845 (N_1845,N_1084,N_1218);
nand U1846 (N_1846,N_1387,N_1159);
nand U1847 (N_1847,N_1269,N_1349);
nor U1848 (N_1848,N_1371,N_1435);
or U1849 (N_1849,N_1397,N_1323);
nand U1850 (N_1850,N_1012,N_1397);
or U1851 (N_1851,N_1418,N_1236);
and U1852 (N_1852,N_1274,N_1147);
or U1853 (N_1853,N_1395,N_1255);
nand U1854 (N_1854,N_1405,N_1485);
nand U1855 (N_1855,N_1407,N_1336);
nand U1856 (N_1856,N_1049,N_1184);
nor U1857 (N_1857,N_1026,N_1359);
and U1858 (N_1858,N_1044,N_1088);
nand U1859 (N_1859,N_1354,N_1369);
and U1860 (N_1860,N_1220,N_1061);
nor U1861 (N_1861,N_1347,N_1123);
nand U1862 (N_1862,N_1166,N_1278);
or U1863 (N_1863,N_1472,N_1293);
or U1864 (N_1864,N_1071,N_1195);
nand U1865 (N_1865,N_1189,N_1086);
nor U1866 (N_1866,N_1356,N_1226);
nor U1867 (N_1867,N_1070,N_1451);
and U1868 (N_1868,N_1076,N_1326);
nor U1869 (N_1869,N_1006,N_1166);
nor U1870 (N_1870,N_1180,N_1095);
and U1871 (N_1871,N_1245,N_1497);
nor U1872 (N_1872,N_1499,N_1004);
nor U1873 (N_1873,N_1190,N_1108);
or U1874 (N_1874,N_1327,N_1168);
or U1875 (N_1875,N_1002,N_1317);
nand U1876 (N_1876,N_1304,N_1034);
nor U1877 (N_1877,N_1245,N_1188);
or U1878 (N_1878,N_1357,N_1054);
or U1879 (N_1879,N_1075,N_1069);
and U1880 (N_1880,N_1470,N_1240);
nand U1881 (N_1881,N_1219,N_1099);
nand U1882 (N_1882,N_1376,N_1257);
or U1883 (N_1883,N_1372,N_1445);
or U1884 (N_1884,N_1135,N_1318);
or U1885 (N_1885,N_1484,N_1078);
nand U1886 (N_1886,N_1434,N_1196);
or U1887 (N_1887,N_1285,N_1159);
or U1888 (N_1888,N_1494,N_1470);
or U1889 (N_1889,N_1180,N_1230);
nand U1890 (N_1890,N_1144,N_1178);
nand U1891 (N_1891,N_1157,N_1101);
or U1892 (N_1892,N_1074,N_1418);
nor U1893 (N_1893,N_1084,N_1452);
or U1894 (N_1894,N_1386,N_1469);
nor U1895 (N_1895,N_1384,N_1165);
nor U1896 (N_1896,N_1141,N_1428);
or U1897 (N_1897,N_1436,N_1246);
nor U1898 (N_1898,N_1039,N_1473);
or U1899 (N_1899,N_1328,N_1441);
nor U1900 (N_1900,N_1340,N_1469);
or U1901 (N_1901,N_1065,N_1410);
or U1902 (N_1902,N_1283,N_1199);
or U1903 (N_1903,N_1027,N_1310);
nor U1904 (N_1904,N_1062,N_1492);
and U1905 (N_1905,N_1396,N_1264);
nor U1906 (N_1906,N_1460,N_1088);
nand U1907 (N_1907,N_1396,N_1164);
or U1908 (N_1908,N_1179,N_1127);
and U1909 (N_1909,N_1154,N_1095);
or U1910 (N_1910,N_1096,N_1264);
or U1911 (N_1911,N_1299,N_1250);
nand U1912 (N_1912,N_1343,N_1415);
and U1913 (N_1913,N_1015,N_1474);
nor U1914 (N_1914,N_1493,N_1461);
or U1915 (N_1915,N_1216,N_1047);
and U1916 (N_1916,N_1374,N_1209);
and U1917 (N_1917,N_1132,N_1343);
and U1918 (N_1918,N_1499,N_1176);
nand U1919 (N_1919,N_1485,N_1461);
and U1920 (N_1920,N_1427,N_1372);
nand U1921 (N_1921,N_1245,N_1248);
and U1922 (N_1922,N_1028,N_1324);
and U1923 (N_1923,N_1183,N_1159);
or U1924 (N_1924,N_1378,N_1321);
nand U1925 (N_1925,N_1115,N_1047);
nand U1926 (N_1926,N_1068,N_1439);
or U1927 (N_1927,N_1301,N_1034);
and U1928 (N_1928,N_1450,N_1115);
nor U1929 (N_1929,N_1034,N_1106);
or U1930 (N_1930,N_1461,N_1368);
or U1931 (N_1931,N_1399,N_1348);
nor U1932 (N_1932,N_1022,N_1425);
and U1933 (N_1933,N_1413,N_1197);
nor U1934 (N_1934,N_1344,N_1138);
nor U1935 (N_1935,N_1168,N_1306);
and U1936 (N_1936,N_1105,N_1430);
and U1937 (N_1937,N_1031,N_1480);
nand U1938 (N_1938,N_1142,N_1206);
or U1939 (N_1939,N_1095,N_1101);
nand U1940 (N_1940,N_1345,N_1476);
or U1941 (N_1941,N_1320,N_1230);
nand U1942 (N_1942,N_1336,N_1014);
or U1943 (N_1943,N_1359,N_1107);
nor U1944 (N_1944,N_1201,N_1296);
nand U1945 (N_1945,N_1303,N_1181);
nor U1946 (N_1946,N_1143,N_1359);
nand U1947 (N_1947,N_1015,N_1167);
nor U1948 (N_1948,N_1376,N_1190);
nor U1949 (N_1949,N_1039,N_1034);
or U1950 (N_1950,N_1080,N_1284);
nand U1951 (N_1951,N_1086,N_1102);
or U1952 (N_1952,N_1030,N_1336);
or U1953 (N_1953,N_1461,N_1481);
or U1954 (N_1954,N_1098,N_1020);
nor U1955 (N_1955,N_1263,N_1413);
nor U1956 (N_1956,N_1285,N_1400);
or U1957 (N_1957,N_1438,N_1100);
or U1958 (N_1958,N_1135,N_1418);
nand U1959 (N_1959,N_1172,N_1085);
and U1960 (N_1960,N_1209,N_1445);
and U1961 (N_1961,N_1195,N_1181);
nand U1962 (N_1962,N_1187,N_1088);
or U1963 (N_1963,N_1184,N_1202);
nor U1964 (N_1964,N_1419,N_1366);
nor U1965 (N_1965,N_1340,N_1084);
or U1966 (N_1966,N_1225,N_1167);
or U1967 (N_1967,N_1160,N_1020);
nor U1968 (N_1968,N_1445,N_1367);
nor U1969 (N_1969,N_1171,N_1350);
and U1970 (N_1970,N_1273,N_1123);
nor U1971 (N_1971,N_1440,N_1415);
nor U1972 (N_1972,N_1217,N_1089);
and U1973 (N_1973,N_1210,N_1277);
or U1974 (N_1974,N_1056,N_1186);
and U1975 (N_1975,N_1011,N_1031);
and U1976 (N_1976,N_1172,N_1066);
and U1977 (N_1977,N_1109,N_1162);
nand U1978 (N_1978,N_1167,N_1071);
or U1979 (N_1979,N_1245,N_1368);
or U1980 (N_1980,N_1045,N_1033);
nor U1981 (N_1981,N_1057,N_1268);
and U1982 (N_1982,N_1286,N_1031);
nand U1983 (N_1983,N_1344,N_1239);
and U1984 (N_1984,N_1413,N_1301);
and U1985 (N_1985,N_1299,N_1451);
nand U1986 (N_1986,N_1047,N_1260);
or U1987 (N_1987,N_1256,N_1079);
and U1988 (N_1988,N_1203,N_1005);
or U1989 (N_1989,N_1165,N_1336);
nor U1990 (N_1990,N_1210,N_1497);
and U1991 (N_1991,N_1056,N_1456);
nand U1992 (N_1992,N_1150,N_1479);
nor U1993 (N_1993,N_1188,N_1329);
nor U1994 (N_1994,N_1128,N_1294);
nand U1995 (N_1995,N_1068,N_1169);
nand U1996 (N_1996,N_1089,N_1123);
nor U1997 (N_1997,N_1497,N_1261);
nand U1998 (N_1998,N_1474,N_1160);
and U1999 (N_1999,N_1162,N_1232);
nand U2000 (N_2000,N_1512,N_1501);
nor U2001 (N_2001,N_1636,N_1643);
and U2002 (N_2002,N_1879,N_1586);
or U2003 (N_2003,N_1579,N_1925);
and U2004 (N_2004,N_1670,N_1793);
and U2005 (N_2005,N_1701,N_1769);
and U2006 (N_2006,N_1943,N_1807);
and U2007 (N_2007,N_1800,N_1983);
nand U2008 (N_2008,N_1536,N_1936);
and U2009 (N_2009,N_1808,N_1559);
and U2010 (N_2010,N_1573,N_1693);
or U2011 (N_2011,N_1588,N_1647);
or U2012 (N_2012,N_1702,N_1872);
or U2013 (N_2013,N_1682,N_1641);
nand U2014 (N_2014,N_1650,N_1757);
nand U2015 (N_2015,N_1881,N_1821);
or U2016 (N_2016,N_1746,N_1562);
nand U2017 (N_2017,N_1803,N_1520);
nand U2018 (N_2018,N_1662,N_1846);
nand U2019 (N_2019,N_1933,N_1502);
or U2020 (N_2020,N_1699,N_1843);
nand U2021 (N_2021,N_1624,N_1784);
or U2022 (N_2022,N_1873,N_1566);
or U2023 (N_2023,N_1688,N_1868);
or U2024 (N_2024,N_1811,N_1564);
and U2025 (N_2025,N_1584,N_1594);
and U2026 (N_2026,N_1984,N_1759);
xor U2027 (N_2027,N_1836,N_1550);
nor U2028 (N_2028,N_1547,N_1833);
or U2029 (N_2029,N_1503,N_1906);
nand U2030 (N_2030,N_1995,N_1866);
nand U2031 (N_2031,N_1830,N_1639);
or U2032 (N_2032,N_1590,N_1954);
or U2033 (N_2033,N_1595,N_1894);
nor U2034 (N_2034,N_1867,N_1953);
or U2035 (N_2035,N_1883,N_1511);
nand U2036 (N_2036,N_1999,N_1542);
and U2037 (N_2037,N_1780,N_1727);
nand U2038 (N_2038,N_1823,N_1797);
and U2039 (N_2039,N_1993,N_1937);
nor U2040 (N_2040,N_1805,N_1630);
nor U2041 (N_2041,N_1723,N_1761);
or U2042 (N_2042,N_1616,N_1825);
or U2043 (N_2043,N_1987,N_1838);
or U2044 (N_2044,N_1979,N_1749);
nand U2045 (N_2045,N_1645,N_1801);
or U2046 (N_2046,N_1692,N_1721);
nor U2047 (N_2047,N_1596,N_1978);
and U2048 (N_2048,N_1629,N_1728);
and U2049 (N_2049,N_1621,N_1895);
and U2050 (N_2050,N_1648,N_1826);
nor U2051 (N_2051,N_1915,N_1926);
nor U2052 (N_2052,N_1612,N_1950);
or U2053 (N_2053,N_1664,N_1877);
nand U2054 (N_2054,N_1582,N_1909);
and U2055 (N_2055,N_1585,N_1975);
or U2056 (N_2056,N_1663,N_1745);
nor U2057 (N_2057,N_1534,N_1944);
or U2058 (N_2058,N_1768,N_1908);
or U2059 (N_2059,N_1731,N_1526);
nor U2060 (N_2060,N_1565,N_1638);
or U2061 (N_2061,N_1733,N_1765);
nand U2062 (N_2062,N_1659,N_1694);
nand U2063 (N_2063,N_1913,N_1608);
nand U2064 (N_2064,N_1890,N_1507);
nand U2065 (N_2065,N_1996,N_1802);
and U2066 (N_2066,N_1773,N_1781);
nand U2067 (N_2067,N_1934,N_1697);
nor U2068 (N_2068,N_1907,N_1851);
nor U2069 (N_2069,N_1666,N_1574);
nor U2070 (N_2070,N_1703,N_1985);
and U2071 (N_2071,N_1632,N_1790);
nor U2072 (N_2072,N_1841,N_1887);
nand U2073 (N_2073,N_1537,N_1738);
and U2074 (N_2074,N_1555,N_1528);
nor U2075 (N_2075,N_1637,N_1928);
nand U2076 (N_2076,N_1712,N_1857);
nor U2077 (N_2077,N_1615,N_1634);
xnor U2078 (N_2078,N_1726,N_1794);
or U2079 (N_2079,N_1543,N_1569);
and U2080 (N_2080,N_1820,N_1893);
or U2081 (N_2081,N_1661,N_1519);
nand U2082 (N_2082,N_1902,N_1905);
and U2083 (N_2083,N_1891,N_1530);
nor U2084 (N_2084,N_1976,N_1743);
and U2085 (N_2085,N_1609,N_1763);
nor U2086 (N_2086,N_1742,N_1824);
nand U2087 (N_2087,N_1737,N_1837);
nand U2088 (N_2088,N_1911,N_1762);
nor U2089 (N_2089,N_1782,N_1923);
and U2090 (N_2090,N_1581,N_1626);
nor U2091 (N_2091,N_1657,N_1690);
nand U2092 (N_2092,N_1809,N_1912);
or U2093 (N_2093,N_1709,N_1561);
nor U2094 (N_2094,N_1989,N_1842);
nand U2095 (N_2095,N_1618,N_1916);
or U2096 (N_2096,N_1570,N_1577);
and U2097 (N_2097,N_1901,N_1527);
or U2098 (N_2098,N_1601,N_1567);
nor U2099 (N_2099,N_1540,N_1840);
nor U2100 (N_2100,N_1655,N_1558);
nand U2101 (N_2101,N_1829,N_1865);
or U2102 (N_2102,N_1597,N_1521);
nor U2103 (N_2103,N_1929,N_1600);
and U2104 (N_2104,N_1997,N_1750);
and U2105 (N_2105,N_1982,N_1844);
or U2106 (N_2106,N_1967,N_1892);
or U2107 (N_2107,N_1516,N_1853);
or U2108 (N_2108,N_1785,N_1869);
nand U2109 (N_2109,N_1810,N_1796);
and U2110 (N_2110,N_1651,N_1748);
or U2111 (N_2111,N_1652,N_1658);
nand U2112 (N_2112,N_1506,N_1930);
nor U2113 (N_2113,N_1505,N_1948);
or U2114 (N_2114,N_1560,N_1813);
nor U2115 (N_2115,N_1741,N_1740);
or U2116 (N_2116,N_1961,N_1628);
and U2117 (N_2117,N_1729,N_1681);
and U2118 (N_2118,N_1646,N_1792);
nand U2119 (N_2119,N_1849,N_1756);
and U2120 (N_2120,N_1962,N_1683);
and U2121 (N_2121,N_1988,N_1971);
or U2122 (N_2122,N_1860,N_1932);
or U2123 (N_2123,N_1722,N_1940);
or U2124 (N_2124,N_1724,N_1777);
and U2125 (N_2125,N_1691,N_1899);
or U2126 (N_2126,N_1964,N_1848);
and U2127 (N_2127,N_1551,N_1568);
and U2128 (N_2128,N_1856,N_1735);
or U2129 (N_2129,N_1958,N_1714);
nor U2130 (N_2130,N_1938,N_1922);
nor U2131 (N_2131,N_1960,N_1529);
and U2132 (N_2132,N_1587,N_1939);
and U2133 (N_2133,N_1970,N_1998);
or U2134 (N_2134,N_1678,N_1610);
nand U2135 (N_2135,N_1719,N_1606);
or U2136 (N_2136,N_1992,N_1607);
or U2137 (N_2137,N_1968,N_1994);
and U2138 (N_2138,N_1775,N_1900);
nand U2139 (N_2139,N_1675,N_1705);
and U2140 (N_2140,N_1966,N_1704);
or U2141 (N_2141,N_1734,N_1642);
and U2142 (N_2142,N_1716,N_1708);
nor U2143 (N_2143,N_1942,N_1973);
or U2144 (N_2144,N_1563,N_1889);
or U2145 (N_2145,N_1874,N_1772);
nor U2146 (N_2146,N_1752,N_1770);
nand U2147 (N_2147,N_1556,N_1924);
nand U2148 (N_2148,N_1766,N_1665);
or U2149 (N_2149,N_1834,N_1653);
nand U2150 (N_2150,N_1700,N_1611);
or U2151 (N_2151,N_1622,N_1832);
or U2152 (N_2152,N_1671,N_1518);
and U2153 (N_2153,N_1522,N_1798);
and U2154 (N_2154,N_1715,N_1620);
or U2155 (N_2155,N_1863,N_1605);
and U2156 (N_2156,N_1875,N_1941);
and U2157 (N_2157,N_1888,N_1686);
or U2158 (N_2158,N_1687,N_1847);
nand U2159 (N_2159,N_1839,N_1627);
nand U2160 (N_2160,N_1783,N_1977);
and U2161 (N_2161,N_1965,N_1854);
or U2162 (N_2162,N_1771,N_1539);
nand U2163 (N_2163,N_1580,N_1515);
or U2164 (N_2164,N_1812,N_1956);
nand U2165 (N_2165,N_1774,N_1730);
xor U2166 (N_2166,N_1592,N_1764);
and U2167 (N_2167,N_1500,N_1882);
nand U2168 (N_2168,N_1602,N_1710);
nor U2169 (N_2169,N_1633,N_1747);
nor U2170 (N_2170,N_1921,N_1945);
nor U2171 (N_2171,N_1946,N_1835);
or U2172 (N_2172,N_1695,N_1754);
nor U2173 (N_2173,N_1786,N_1986);
nor U2174 (N_2174,N_1778,N_1957);
or U2175 (N_2175,N_1787,N_1649);
xor U2176 (N_2176,N_1862,N_1679);
and U2177 (N_2177,N_1598,N_1583);
or U2178 (N_2178,N_1919,N_1935);
nand U2179 (N_2179,N_1546,N_1532);
and U2180 (N_2180,N_1673,N_1917);
nand U2181 (N_2181,N_1739,N_1514);
nor U2182 (N_2182,N_1791,N_1914);
and U2183 (N_2183,N_1955,N_1903);
and U2184 (N_2184,N_1549,N_1969);
or U2185 (N_2185,N_1885,N_1725);
and U2186 (N_2186,N_1776,N_1918);
nor U2187 (N_2187,N_1852,N_1816);
or U2188 (N_2188,N_1572,N_1508);
or U2189 (N_2189,N_1613,N_1713);
and U2190 (N_2190,N_1603,N_1804);
and U2191 (N_2191,N_1717,N_1544);
nor U2192 (N_2192,N_1656,N_1760);
nor U2193 (N_2193,N_1677,N_1896);
nand U2194 (N_2194,N_1654,N_1980);
and U2195 (N_2195,N_1698,N_1758);
or U2196 (N_2196,N_1513,N_1861);
or U2197 (N_2197,N_1541,N_1554);
and U2198 (N_2198,N_1755,N_1814);
and U2199 (N_2199,N_1795,N_1689);
nor U2200 (N_2200,N_1864,N_1711);
nand U2201 (N_2201,N_1720,N_1667);
nor U2202 (N_2202,N_1949,N_1631);
or U2203 (N_2203,N_1952,N_1974);
nand U2204 (N_2204,N_1817,N_1831);
or U2205 (N_2205,N_1523,N_1990);
and U2206 (N_2206,N_1676,N_1828);
nand U2207 (N_2207,N_1669,N_1951);
nand U2208 (N_2208,N_1707,N_1927);
nor U2209 (N_2209,N_1684,N_1880);
nor U2210 (N_2210,N_1789,N_1644);
nor U2211 (N_2211,N_1640,N_1668);
nor U2212 (N_2212,N_1672,N_1576);
or U2213 (N_2213,N_1845,N_1753);
or U2214 (N_2214,N_1876,N_1571);
or U2215 (N_2215,N_1799,N_1991);
nand U2216 (N_2216,N_1859,N_1827);
nand U2217 (N_2217,N_1878,N_1545);
nand U2218 (N_2218,N_1972,N_1718);
and U2219 (N_2219,N_1910,N_1660);
nor U2220 (N_2220,N_1931,N_1779);
nand U2221 (N_2221,N_1619,N_1504);
or U2222 (N_2222,N_1591,N_1674);
nor U2223 (N_2223,N_1818,N_1815);
nor U2224 (N_2224,N_1788,N_1806);
or U2225 (N_2225,N_1870,N_1947);
and U2226 (N_2226,N_1578,N_1517);
nor U2227 (N_2227,N_1819,N_1524);
or U2228 (N_2228,N_1920,N_1886);
nand U2229 (N_2229,N_1552,N_1538);
or U2230 (N_2230,N_1736,N_1589);
nor U2231 (N_2231,N_1963,N_1625);
nand U2232 (N_2232,N_1680,N_1751);
or U2233 (N_2233,N_1533,N_1593);
or U2234 (N_2234,N_1897,N_1696);
nand U2235 (N_2235,N_1904,N_1604);
nand U2236 (N_2236,N_1557,N_1525);
and U2237 (N_2237,N_1531,N_1884);
nand U2238 (N_2238,N_1685,N_1535);
and U2239 (N_2239,N_1744,N_1732);
nand U2240 (N_2240,N_1898,N_1767);
and U2241 (N_2241,N_1850,N_1871);
or U2242 (N_2242,N_1855,N_1623);
and U2243 (N_2243,N_1553,N_1981);
or U2244 (N_2244,N_1614,N_1822);
xnor U2245 (N_2245,N_1635,N_1706);
and U2246 (N_2246,N_1575,N_1858);
and U2247 (N_2247,N_1599,N_1509);
and U2248 (N_2248,N_1617,N_1959);
xnor U2249 (N_2249,N_1510,N_1548);
nand U2250 (N_2250,N_1919,N_1739);
and U2251 (N_2251,N_1587,N_1869);
nand U2252 (N_2252,N_1995,N_1909);
nand U2253 (N_2253,N_1890,N_1797);
and U2254 (N_2254,N_1665,N_1660);
and U2255 (N_2255,N_1811,N_1931);
nor U2256 (N_2256,N_1890,N_1786);
nand U2257 (N_2257,N_1772,N_1866);
or U2258 (N_2258,N_1770,N_1838);
nor U2259 (N_2259,N_1801,N_1676);
or U2260 (N_2260,N_1797,N_1540);
and U2261 (N_2261,N_1785,N_1501);
nor U2262 (N_2262,N_1959,N_1589);
or U2263 (N_2263,N_1633,N_1573);
or U2264 (N_2264,N_1729,N_1641);
and U2265 (N_2265,N_1661,N_1755);
xnor U2266 (N_2266,N_1836,N_1536);
and U2267 (N_2267,N_1939,N_1647);
nand U2268 (N_2268,N_1860,N_1963);
nor U2269 (N_2269,N_1537,N_1924);
nand U2270 (N_2270,N_1658,N_1832);
nor U2271 (N_2271,N_1737,N_1648);
or U2272 (N_2272,N_1967,N_1609);
or U2273 (N_2273,N_1770,N_1802);
and U2274 (N_2274,N_1596,N_1760);
or U2275 (N_2275,N_1773,N_1512);
or U2276 (N_2276,N_1826,N_1877);
nand U2277 (N_2277,N_1508,N_1953);
or U2278 (N_2278,N_1706,N_1634);
and U2279 (N_2279,N_1885,N_1645);
xor U2280 (N_2280,N_1614,N_1814);
nor U2281 (N_2281,N_1953,N_1956);
nand U2282 (N_2282,N_1738,N_1728);
nor U2283 (N_2283,N_1729,N_1776);
nand U2284 (N_2284,N_1510,N_1935);
nand U2285 (N_2285,N_1977,N_1769);
nand U2286 (N_2286,N_1550,N_1953);
nand U2287 (N_2287,N_1645,N_1970);
and U2288 (N_2288,N_1856,N_1968);
and U2289 (N_2289,N_1842,N_1786);
nand U2290 (N_2290,N_1874,N_1586);
nand U2291 (N_2291,N_1813,N_1505);
nor U2292 (N_2292,N_1575,N_1850);
or U2293 (N_2293,N_1793,N_1846);
nand U2294 (N_2294,N_1722,N_1534);
or U2295 (N_2295,N_1918,N_1824);
nor U2296 (N_2296,N_1536,N_1581);
nor U2297 (N_2297,N_1979,N_1847);
or U2298 (N_2298,N_1586,N_1835);
nand U2299 (N_2299,N_1826,N_1597);
nor U2300 (N_2300,N_1835,N_1593);
nor U2301 (N_2301,N_1961,N_1886);
nor U2302 (N_2302,N_1506,N_1843);
nand U2303 (N_2303,N_1932,N_1823);
and U2304 (N_2304,N_1723,N_1655);
nor U2305 (N_2305,N_1554,N_1913);
nor U2306 (N_2306,N_1866,N_1953);
nand U2307 (N_2307,N_1736,N_1603);
and U2308 (N_2308,N_1648,N_1549);
nand U2309 (N_2309,N_1502,N_1665);
and U2310 (N_2310,N_1953,N_1618);
or U2311 (N_2311,N_1863,N_1530);
nor U2312 (N_2312,N_1894,N_1991);
and U2313 (N_2313,N_1566,N_1524);
nand U2314 (N_2314,N_1916,N_1840);
or U2315 (N_2315,N_1587,N_1668);
nand U2316 (N_2316,N_1989,N_1869);
and U2317 (N_2317,N_1957,N_1557);
or U2318 (N_2318,N_1842,N_1879);
and U2319 (N_2319,N_1912,N_1975);
nand U2320 (N_2320,N_1598,N_1631);
nor U2321 (N_2321,N_1864,N_1628);
nor U2322 (N_2322,N_1601,N_1962);
and U2323 (N_2323,N_1521,N_1612);
or U2324 (N_2324,N_1596,N_1817);
and U2325 (N_2325,N_1525,N_1884);
nor U2326 (N_2326,N_1955,N_1747);
and U2327 (N_2327,N_1947,N_1583);
or U2328 (N_2328,N_1841,N_1715);
nand U2329 (N_2329,N_1656,N_1687);
nand U2330 (N_2330,N_1916,N_1918);
or U2331 (N_2331,N_1638,N_1768);
nor U2332 (N_2332,N_1919,N_1565);
or U2333 (N_2333,N_1737,N_1639);
nor U2334 (N_2334,N_1952,N_1710);
or U2335 (N_2335,N_1670,N_1931);
nand U2336 (N_2336,N_1755,N_1627);
and U2337 (N_2337,N_1707,N_1680);
nor U2338 (N_2338,N_1641,N_1615);
and U2339 (N_2339,N_1769,N_1641);
and U2340 (N_2340,N_1791,N_1821);
nand U2341 (N_2341,N_1942,N_1833);
or U2342 (N_2342,N_1761,N_1886);
nor U2343 (N_2343,N_1558,N_1870);
and U2344 (N_2344,N_1862,N_1826);
nand U2345 (N_2345,N_1572,N_1553);
nand U2346 (N_2346,N_1872,N_1791);
or U2347 (N_2347,N_1701,N_1560);
nand U2348 (N_2348,N_1782,N_1878);
nor U2349 (N_2349,N_1803,N_1808);
nor U2350 (N_2350,N_1872,N_1551);
and U2351 (N_2351,N_1707,N_1535);
and U2352 (N_2352,N_1831,N_1758);
and U2353 (N_2353,N_1518,N_1565);
nand U2354 (N_2354,N_1563,N_1734);
and U2355 (N_2355,N_1817,N_1550);
nand U2356 (N_2356,N_1689,N_1891);
nor U2357 (N_2357,N_1811,N_1688);
and U2358 (N_2358,N_1679,N_1932);
nor U2359 (N_2359,N_1725,N_1662);
nand U2360 (N_2360,N_1780,N_1567);
nor U2361 (N_2361,N_1928,N_1754);
nand U2362 (N_2362,N_1862,N_1577);
nand U2363 (N_2363,N_1956,N_1796);
and U2364 (N_2364,N_1641,N_1857);
nor U2365 (N_2365,N_1700,N_1584);
and U2366 (N_2366,N_1762,N_1648);
or U2367 (N_2367,N_1854,N_1801);
nor U2368 (N_2368,N_1518,N_1785);
or U2369 (N_2369,N_1829,N_1906);
nor U2370 (N_2370,N_1635,N_1916);
nor U2371 (N_2371,N_1786,N_1866);
nand U2372 (N_2372,N_1925,N_1769);
nand U2373 (N_2373,N_1607,N_1854);
nand U2374 (N_2374,N_1731,N_1574);
nand U2375 (N_2375,N_1651,N_1948);
or U2376 (N_2376,N_1962,N_1525);
nand U2377 (N_2377,N_1639,N_1891);
nor U2378 (N_2378,N_1591,N_1770);
or U2379 (N_2379,N_1869,N_1968);
nand U2380 (N_2380,N_1695,N_1726);
and U2381 (N_2381,N_1927,N_1895);
nor U2382 (N_2382,N_1615,N_1986);
or U2383 (N_2383,N_1554,N_1701);
nand U2384 (N_2384,N_1626,N_1586);
nand U2385 (N_2385,N_1532,N_1888);
nor U2386 (N_2386,N_1892,N_1765);
or U2387 (N_2387,N_1646,N_1643);
nand U2388 (N_2388,N_1517,N_1998);
nor U2389 (N_2389,N_1594,N_1977);
nand U2390 (N_2390,N_1836,N_1735);
nor U2391 (N_2391,N_1846,N_1710);
nand U2392 (N_2392,N_1957,N_1623);
nand U2393 (N_2393,N_1827,N_1759);
nor U2394 (N_2394,N_1901,N_1556);
and U2395 (N_2395,N_1956,N_1512);
and U2396 (N_2396,N_1844,N_1851);
and U2397 (N_2397,N_1766,N_1736);
and U2398 (N_2398,N_1556,N_1813);
or U2399 (N_2399,N_1904,N_1662);
and U2400 (N_2400,N_1976,N_1689);
or U2401 (N_2401,N_1572,N_1883);
nand U2402 (N_2402,N_1648,N_1760);
nor U2403 (N_2403,N_1527,N_1670);
nand U2404 (N_2404,N_1797,N_1967);
or U2405 (N_2405,N_1613,N_1528);
and U2406 (N_2406,N_1943,N_1590);
or U2407 (N_2407,N_1731,N_1806);
or U2408 (N_2408,N_1985,N_1768);
or U2409 (N_2409,N_1911,N_1613);
and U2410 (N_2410,N_1850,N_1584);
or U2411 (N_2411,N_1676,N_1798);
nor U2412 (N_2412,N_1686,N_1919);
nor U2413 (N_2413,N_1572,N_1828);
and U2414 (N_2414,N_1997,N_1747);
nand U2415 (N_2415,N_1790,N_1641);
nand U2416 (N_2416,N_1732,N_1620);
and U2417 (N_2417,N_1873,N_1557);
and U2418 (N_2418,N_1854,N_1833);
or U2419 (N_2419,N_1833,N_1645);
or U2420 (N_2420,N_1866,N_1823);
nand U2421 (N_2421,N_1539,N_1733);
nand U2422 (N_2422,N_1814,N_1745);
nor U2423 (N_2423,N_1633,N_1602);
and U2424 (N_2424,N_1910,N_1621);
nor U2425 (N_2425,N_1580,N_1677);
or U2426 (N_2426,N_1628,N_1792);
nor U2427 (N_2427,N_1737,N_1982);
and U2428 (N_2428,N_1922,N_1608);
and U2429 (N_2429,N_1569,N_1809);
or U2430 (N_2430,N_1692,N_1795);
nor U2431 (N_2431,N_1581,N_1690);
or U2432 (N_2432,N_1707,N_1759);
or U2433 (N_2433,N_1757,N_1836);
or U2434 (N_2434,N_1808,N_1753);
nand U2435 (N_2435,N_1815,N_1543);
nor U2436 (N_2436,N_1999,N_1611);
nand U2437 (N_2437,N_1792,N_1854);
and U2438 (N_2438,N_1918,N_1576);
or U2439 (N_2439,N_1833,N_1954);
nor U2440 (N_2440,N_1905,N_1626);
xor U2441 (N_2441,N_1901,N_1660);
nor U2442 (N_2442,N_1703,N_1590);
or U2443 (N_2443,N_1844,N_1526);
nand U2444 (N_2444,N_1541,N_1581);
or U2445 (N_2445,N_1895,N_1711);
and U2446 (N_2446,N_1656,N_1878);
nand U2447 (N_2447,N_1731,N_1596);
and U2448 (N_2448,N_1678,N_1898);
nand U2449 (N_2449,N_1532,N_1867);
and U2450 (N_2450,N_1897,N_1823);
nand U2451 (N_2451,N_1699,N_1826);
nor U2452 (N_2452,N_1959,N_1862);
and U2453 (N_2453,N_1559,N_1903);
or U2454 (N_2454,N_1610,N_1613);
nor U2455 (N_2455,N_1944,N_1945);
nand U2456 (N_2456,N_1796,N_1688);
nor U2457 (N_2457,N_1761,N_1635);
nand U2458 (N_2458,N_1804,N_1755);
nand U2459 (N_2459,N_1837,N_1792);
nand U2460 (N_2460,N_1622,N_1643);
nand U2461 (N_2461,N_1712,N_1655);
nor U2462 (N_2462,N_1840,N_1675);
nor U2463 (N_2463,N_1926,N_1505);
or U2464 (N_2464,N_1785,N_1875);
and U2465 (N_2465,N_1727,N_1615);
nor U2466 (N_2466,N_1829,N_1723);
nand U2467 (N_2467,N_1633,N_1687);
nor U2468 (N_2468,N_1710,N_1707);
nand U2469 (N_2469,N_1687,N_1703);
and U2470 (N_2470,N_1970,N_1684);
nand U2471 (N_2471,N_1840,N_1894);
and U2472 (N_2472,N_1629,N_1662);
or U2473 (N_2473,N_1929,N_1554);
or U2474 (N_2474,N_1632,N_1773);
or U2475 (N_2475,N_1944,N_1747);
nand U2476 (N_2476,N_1629,N_1993);
or U2477 (N_2477,N_1638,N_1744);
or U2478 (N_2478,N_1803,N_1960);
and U2479 (N_2479,N_1888,N_1544);
or U2480 (N_2480,N_1506,N_1918);
and U2481 (N_2481,N_1870,N_1523);
and U2482 (N_2482,N_1808,N_1556);
or U2483 (N_2483,N_1626,N_1616);
or U2484 (N_2484,N_1813,N_1914);
nor U2485 (N_2485,N_1773,N_1880);
or U2486 (N_2486,N_1853,N_1777);
and U2487 (N_2487,N_1879,N_1802);
nor U2488 (N_2488,N_1946,N_1621);
or U2489 (N_2489,N_1605,N_1890);
or U2490 (N_2490,N_1655,N_1835);
or U2491 (N_2491,N_1675,N_1566);
nor U2492 (N_2492,N_1785,N_1653);
and U2493 (N_2493,N_1663,N_1696);
nand U2494 (N_2494,N_1948,N_1807);
xnor U2495 (N_2495,N_1644,N_1590);
and U2496 (N_2496,N_1520,N_1831);
and U2497 (N_2497,N_1833,N_1632);
or U2498 (N_2498,N_1769,N_1880);
or U2499 (N_2499,N_1766,N_1690);
nor U2500 (N_2500,N_2398,N_2494);
xnor U2501 (N_2501,N_2059,N_2286);
nand U2502 (N_2502,N_2143,N_2264);
and U2503 (N_2503,N_2141,N_2316);
and U2504 (N_2504,N_2047,N_2228);
or U2505 (N_2505,N_2462,N_2038);
nand U2506 (N_2506,N_2114,N_2474);
and U2507 (N_2507,N_2050,N_2176);
xor U2508 (N_2508,N_2083,N_2188);
and U2509 (N_2509,N_2233,N_2307);
nor U2510 (N_2510,N_2285,N_2111);
nor U2511 (N_2511,N_2464,N_2475);
and U2512 (N_2512,N_2063,N_2287);
and U2513 (N_2513,N_2385,N_2219);
or U2514 (N_2514,N_2397,N_2218);
nand U2515 (N_2515,N_2488,N_2422);
nand U2516 (N_2516,N_2117,N_2189);
nand U2517 (N_2517,N_2186,N_2262);
or U2518 (N_2518,N_2314,N_2357);
and U2519 (N_2519,N_2402,N_2377);
nor U2520 (N_2520,N_2208,N_2267);
or U2521 (N_2521,N_2336,N_2042);
and U2522 (N_2522,N_2044,N_2294);
and U2523 (N_2523,N_2325,N_2106);
or U2524 (N_2524,N_2386,N_2115);
and U2525 (N_2525,N_2376,N_2012);
nor U2526 (N_2526,N_2322,N_2053);
nor U2527 (N_2527,N_2400,N_2079);
nor U2528 (N_2528,N_2473,N_2088);
nand U2529 (N_2529,N_2452,N_2399);
xnor U2530 (N_2530,N_2362,N_2209);
xor U2531 (N_2531,N_2436,N_2277);
nand U2532 (N_2532,N_2230,N_2102);
nor U2533 (N_2533,N_2035,N_2393);
and U2534 (N_2534,N_2305,N_2387);
nand U2535 (N_2535,N_2247,N_2346);
and U2536 (N_2536,N_2283,N_2270);
or U2537 (N_2537,N_2185,N_2232);
or U2538 (N_2538,N_2345,N_2451);
nand U2539 (N_2539,N_2168,N_2371);
or U2540 (N_2540,N_2253,N_2204);
and U2541 (N_2541,N_2093,N_2197);
or U2542 (N_2542,N_2401,N_2472);
nor U2543 (N_2543,N_2309,N_2036);
nor U2544 (N_2544,N_2011,N_2368);
nor U2545 (N_2545,N_2434,N_2476);
and U2546 (N_2546,N_2173,N_2203);
and U2547 (N_2547,N_2131,N_2238);
nand U2548 (N_2548,N_2082,N_2146);
nor U2549 (N_2549,N_2084,N_2340);
and U2550 (N_2550,N_2181,N_2463);
or U2551 (N_2551,N_2034,N_2221);
and U2552 (N_2552,N_2183,N_2407);
and U2553 (N_2553,N_2388,N_2123);
nand U2554 (N_2554,N_2069,N_2259);
nor U2555 (N_2555,N_2236,N_2423);
or U2556 (N_2556,N_2070,N_2097);
nor U2557 (N_2557,N_2160,N_2443);
or U2558 (N_2558,N_2220,N_2394);
nand U2559 (N_2559,N_2136,N_2212);
nor U2560 (N_2560,N_2293,N_2354);
nand U2561 (N_2561,N_2017,N_2284);
nand U2562 (N_2562,N_2075,N_2095);
or U2563 (N_2563,N_2049,N_2105);
and U2564 (N_2564,N_2409,N_2348);
nand U2565 (N_2565,N_2190,N_2458);
xnor U2566 (N_2566,N_2216,N_2091);
or U2567 (N_2567,N_2299,N_2447);
nand U2568 (N_2568,N_2437,N_2078);
and U2569 (N_2569,N_2275,N_2032);
nand U2570 (N_2570,N_2415,N_2000);
nand U2571 (N_2571,N_2297,N_2318);
nor U2572 (N_2572,N_2470,N_2425);
and U2573 (N_2573,N_2308,N_2243);
nand U2574 (N_2574,N_2483,N_2057);
nand U2575 (N_2575,N_2090,N_2410);
nor U2576 (N_2576,N_2298,N_2266);
nand U2577 (N_2577,N_2113,N_2302);
nor U2578 (N_2578,N_2353,N_2380);
and U2579 (N_2579,N_2107,N_2058);
or U2580 (N_2580,N_2338,N_2015);
and U2581 (N_2581,N_2331,N_2004);
and U2582 (N_2582,N_2389,N_2237);
or U2583 (N_2583,N_2223,N_2485);
and U2584 (N_2584,N_2092,N_2229);
and U2585 (N_2585,N_2184,N_2144);
and U2586 (N_2586,N_2125,N_2450);
or U2587 (N_2587,N_2002,N_2198);
nor U2588 (N_2588,N_2326,N_2449);
or U2589 (N_2589,N_2067,N_2039);
nand U2590 (N_2590,N_2043,N_2076);
nand U2591 (N_2591,N_2295,N_2022);
and U2592 (N_2592,N_2211,N_2148);
and U2593 (N_2593,N_2018,N_2135);
or U2594 (N_2594,N_2177,N_2033);
nor U2595 (N_2595,N_2440,N_2482);
nor U2596 (N_2596,N_2013,N_2352);
nor U2597 (N_2597,N_2477,N_2147);
or U2598 (N_2598,N_2260,N_2263);
and U2599 (N_2599,N_2414,N_2214);
nand U2600 (N_2600,N_2174,N_2094);
or U2601 (N_2601,N_2241,N_2031);
nor U2602 (N_2602,N_2142,N_2210);
or U2603 (N_2603,N_2392,N_2225);
or U2604 (N_2604,N_2378,N_2244);
nand U2605 (N_2605,N_2341,N_2065);
or U2606 (N_2606,N_2048,N_2427);
nand U2607 (N_2607,N_2312,N_2311);
or U2608 (N_2608,N_2444,N_2453);
or U2609 (N_2609,N_2213,N_2104);
nand U2610 (N_2610,N_2467,N_2372);
and U2611 (N_2611,N_2124,N_2207);
nand U2612 (N_2612,N_2412,N_2342);
or U2613 (N_2613,N_2037,N_2226);
nor U2614 (N_2614,N_2152,N_2460);
nor U2615 (N_2615,N_2491,N_2480);
nor U2616 (N_2616,N_2112,N_2315);
and U2617 (N_2617,N_2138,N_2156);
and U2618 (N_2618,N_2003,N_2461);
and U2619 (N_2619,N_2149,N_2347);
xnor U2620 (N_2620,N_2193,N_2364);
nand U2621 (N_2621,N_2014,N_2154);
or U2622 (N_2622,N_2206,N_2187);
or U2623 (N_2623,N_2391,N_2010);
nand U2624 (N_2624,N_2195,N_2465);
or U2625 (N_2625,N_2040,N_2441);
or U2626 (N_2626,N_2413,N_2296);
or U2627 (N_2627,N_2484,N_2481);
or U2628 (N_2628,N_2426,N_2313);
nor U2629 (N_2629,N_2051,N_2055);
nor U2630 (N_2630,N_2435,N_2269);
or U2631 (N_2631,N_2019,N_2157);
nor U2632 (N_2632,N_2418,N_2486);
nand U2633 (N_2633,N_2265,N_2268);
or U2634 (N_2634,N_2317,N_2170);
nand U2635 (N_2635,N_2356,N_2257);
nor U2636 (N_2636,N_2217,N_2324);
or U2637 (N_2637,N_2344,N_2430);
or U2638 (N_2638,N_2224,N_2278);
nor U2639 (N_2639,N_2116,N_2360);
and U2640 (N_2640,N_2479,N_2246);
nand U2641 (N_2641,N_2381,N_2273);
and U2642 (N_2642,N_2321,N_2178);
nor U2643 (N_2643,N_2457,N_2099);
nor U2644 (N_2644,N_2245,N_2098);
and U2645 (N_2645,N_2439,N_2350);
nand U2646 (N_2646,N_2056,N_2454);
nand U2647 (N_2647,N_2054,N_2169);
nand U2648 (N_2648,N_2007,N_2172);
and U2649 (N_2649,N_2145,N_2100);
and U2650 (N_2650,N_2367,N_2122);
and U2651 (N_2651,N_2096,N_2199);
nor U2652 (N_2652,N_2175,N_2406);
nand U2653 (N_2653,N_2066,N_2041);
nor U2654 (N_2654,N_2155,N_2163);
nand U2655 (N_2655,N_2196,N_2490);
or U2656 (N_2656,N_2194,N_2395);
nand U2657 (N_2657,N_2129,N_2432);
and U2658 (N_2658,N_2251,N_2256);
or U2659 (N_2659,N_2153,N_2016);
nor U2660 (N_2660,N_2408,N_2358);
and U2661 (N_2661,N_2008,N_2180);
or U2662 (N_2662,N_2110,N_2165);
or U2663 (N_2663,N_2499,N_2121);
nand U2664 (N_2664,N_2020,N_2234);
nor U2665 (N_2665,N_2349,N_2061);
nand U2666 (N_2666,N_2201,N_2127);
nand U2667 (N_2667,N_2329,N_2289);
nor U2668 (N_2668,N_2300,N_2366);
and U2669 (N_2669,N_2151,N_2081);
nand U2670 (N_2670,N_2001,N_2108);
nand U2671 (N_2671,N_2379,N_2416);
and U2672 (N_2672,N_2179,N_2159);
nand U2673 (N_2673,N_2009,N_2323);
nor U2674 (N_2674,N_2327,N_2139);
and U2675 (N_2675,N_2133,N_2292);
nor U2676 (N_2676,N_2134,N_2428);
nand U2677 (N_2677,N_2077,N_2478);
nand U2678 (N_2678,N_2369,N_2337);
nand U2679 (N_2679,N_2074,N_2024);
nor U2680 (N_2680,N_2046,N_2351);
xor U2681 (N_2681,N_2445,N_2085);
xor U2682 (N_2682,N_2469,N_2227);
nor U2683 (N_2683,N_2442,N_2384);
xor U2684 (N_2684,N_2021,N_2330);
nand U2685 (N_2685,N_2334,N_2242);
nand U2686 (N_2686,N_2304,N_2261);
or U2687 (N_2687,N_2150,N_2167);
nand U2688 (N_2688,N_2468,N_2373);
or U2689 (N_2689,N_2332,N_2489);
and U2690 (N_2690,N_2252,N_2166);
nand U2691 (N_2691,N_2333,N_2493);
and U2692 (N_2692,N_2086,N_2320);
and U2693 (N_2693,N_2071,N_2029);
nand U2694 (N_2694,N_2140,N_2158);
nand U2695 (N_2695,N_2382,N_2404);
nand U2696 (N_2696,N_2306,N_2433);
or U2697 (N_2697,N_2192,N_2466);
nor U2698 (N_2698,N_2310,N_2006);
and U2699 (N_2699,N_2103,N_2281);
or U2700 (N_2700,N_2126,N_2487);
or U2701 (N_2701,N_2420,N_2355);
and U2702 (N_2702,N_2130,N_2471);
nor U2703 (N_2703,N_2164,N_2424);
or U2704 (N_2704,N_2446,N_2301);
or U2705 (N_2705,N_2411,N_2249);
nand U2706 (N_2706,N_2492,N_2374);
or U2707 (N_2707,N_2419,N_2182);
nor U2708 (N_2708,N_2254,N_2335);
and U2709 (N_2709,N_2248,N_2025);
and U2710 (N_2710,N_2137,N_2162);
nor U2711 (N_2711,N_2101,N_2459);
nor U2712 (N_2712,N_2359,N_2279);
nand U2713 (N_2713,N_2403,N_2250);
and U2714 (N_2714,N_2343,N_2319);
and U2715 (N_2715,N_2365,N_2240);
nor U2716 (N_2716,N_2222,N_2089);
nor U2717 (N_2717,N_2235,N_2073);
and U2718 (N_2718,N_2291,N_2421);
or U2719 (N_2719,N_2231,N_2087);
and U2720 (N_2720,N_2200,N_2361);
or U2721 (N_2721,N_2328,N_2438);
nor U2722 (N_2722,N_2498,N_2191);
nand U2723 (N_2723,N_2288,N_2495);
nor U2724 (N_2724,N_2429,N_2271);
nor U2725 (N_2725,N_2405,N_2128);
and U2726 (N_2726,N_2072,N_2202);
and U2727 (N_2727,N_2026,N_2496);
or U2728 (N_2728,N_2052,N_2119);
nand U2729 (N_2729,N_2161,N_2456);
nand U2730 (N_2730,N_2120,N_2045);
and U2731 (N_2731,N_2258,N_2396);
or U2732 (N_2732,N_2363,N_2370);
and U2733 (N_2733,N_2431,N_2109);
nor U2734 (N_2734,N_2455,N_2027);
nor U2735 (N_2735,N_2030,N_2303);
and U2736 (N_2736,N_2171,N_2239);
nand U2737 (N_2737,N_2080,N_2448);
or U2738 (N_2738,N_2282,N_2023);
nand U2739 (N_2739,N_2255,N_2375);
nor U2740 (N_2740,N_2497,N_2005);
and U2741 (N_2741,N_2383,N_2276);
and U2742 (N_2742,N_2390,N_2064);
and U2743 (N_2743,N_2068,N_2280);
and U2744 (N_2744,N_2272,N_2290);
nand U2745 (N_2745,N_2205,N_2417);
and U2746 (N_2746,N_2060,N_2274);
and U2747 (N_2747,N_2132,N_2215);
nand U2748 (N_2748,N_2062,N_2028);
nor U2749 (N_2749,N_2339,N_2118);
nor U2750 (N_2750,N_2023,N_2144);
or U2751 (N_2751,N_2339,N_2145);
nor U2752 (N_2752,N_2008,N_2093);
or U2753 (N_2753,N_2326,N_2450);
nand U2754 (N_2754,N_2431,N_2382);
or U2755 (N_2755,N_2130,N_2183);
nand U2756 (N_2756,N_2061,N_2411);
nand U2757 (N_2757,N_2315,N_2192);
or U2758 (N_2758,N_2214,N_2298);
and U2759 (N_2759,N_2309,N_2024);
nand U2760 (N_2760,N_2021,N_2049);
or U2761 (N_2761,N_2220,N_2403);
nor U2762 (N_2762,N_2407,N_2486);
or U2763 (N_2763,N_2418,N_2227);
and U2764 (N_2764,N_2188,N_2003);
and U2765 (N_2765,N_2479,N_2424);
nor U2766 (N_2766,N_2481,N_2483);
nand U2767 (N_2767,N_2160,N_2371);
xor U2768 (N_2768,N_2066,N_2459);
and U2769 (N_2769,N_2353,N_2130);
or U2770 (N_2770,N_2411,N_2351);
and U2771 (N_2771,N_2282,N_2206);
nor U2772 (N_2772,N_2119,N_2110);
or U2773 (N_2773,N_2199,N_2446);
and U2774 (N_2774,N_2151,N_2126);
and U2775 (N_2775,N_2393,N_2353);
nand U2776 (N_2776,N_2281,N_2243);
nor U2777 (N_2777,N_2084,N_2137);
or U2778 (N_2778,N_2068,N_2006);
and U2779 (N_2779,N_2429,N_2233);
nand U2780 (N_2780,N_2410,N_2307);
or U2781 (N_2781,N_2490,N_2241);
nand U2782 (N_2782,N_2488,N_2326);
nand U2783 (N_2783,N_2389,N_2204);
and U2784 (N_2784,N_2210,N_2261);
or U2785 (N_2785,N_2239,N_2004);
nand U2786 (N_2786,N_2046,N_2114);
and U2787 (N_2787,N_2180,N_2271);
nand U2788 (N_2788,N_2350,N_2381);
nor U2789 (N_2789,N_2066,N_2385);
or U2790 (N_2790,N_2268,N_2019);
or U2791 (N_2791,N_2342,N_2392);
nand U2792 (N_2792,N_2314,N_2046);
nor U2793 (N_2793,N_2391,N_2041);
and U2794 (N_2794,N_2305,N_2275);
nor U2795 (N_2795,N_2040,N_2395);
or U2796 (N_2796,N_2099,N_2088);
and U2797 (N_2797,N_2064,N_2037);
and U2798 (N_2798,N_2211,N_2015);
or U2799 (N_2799,N_2246,N_2315);
and U2800 (N_2800,N_2145,N_2032);
and U2801 (N_2801,N_2343,N_2051);
and U2802 (N_2802,N_2078,N_2446);
nand U2803 (N_2803,N_2220,N_2152);
nand U2804 (N_2804,N_2193,N_2293);
and U2805 (N_2805,N_2241,N_2228);
and U2806 (N_2806,N_2434,N_2141);
and U2807 (N_2807,N_2253,N_2232);
or U2808 (N_2808,N_2111,N_2487);
or U2809 (N_2809,N_2069,N_2436);
and U2810 (N_2810,N_2161,N_2248);
or U2811 (N_2811,N_2131,N_2186);
xor U2812 (N_2812,N_2364,N_2480);
nand U2813 (N_2813,N_2392,N_2099);
and U2814 (N_2814,N_2368,N_2294);
nor U2815 (N_2815,N_2332,N_2303);
nand U2816 (N_2816,N_2019,N_2280);
nor U2817 (N_2817,N_2404,N_2222);
nor U2818 (N_2818,N_2103,N_2238);
or U2819 (N_2819,N_2108,N_2174);
or U2820 (N_2820,N_2247,N_2470);
nor U2821 (N_2821,N_2003,N_2363);
and U2822 (N_2822,N_2080,N_2139);
or U2823 (N_2823,N_2437,N_2461);
and U2824 (N_2824,N_2047,N_2238);
and U2825 (N_2825,N_2089,N_2161);
or U2826 (N_2826,N_2182,N_2068);
nor U2827 (N_2827,N_2252,N_2251);
or U2828 (N_2828,N_2444,N_2400);
and U2829 (N_2829,N_2195,N_2189);
and U2830 (N_2830,N_2357,N_2049);
nand U2831 (N_2831,N_2102,N_2333);
nand U2832 (N_2832,N_2409,N_2410);
nor U2833 (N_2833,N_2235,N_2130);
or U2834 (N_2834,N_2002,N_2195);
nand U2835 (N_2835,N_2457,N_2388);
and U2836 (N_2836,N_2136,N_2424);
and U2837 (N_2837,N_2411,N_2039);
nor U2838 (N_2838,N_2348,N_2335);
or U2839 (N_2839,N_2112,N_2466);
or U2840 (N_2840,N_2484,N_2198);
or U2841 (N_2841,N_2121,N_2297);
nand U2842 (N_2842,N_2290,N_2009);
nand U2843 (N_2843,N_2106,N_2039);
and U2844 (N_2844,N_2266,N_2303);
and U2845 (N_2845,N_2061,N_2164);
nand U2846 (N_2846,N_2287,N_2397);
nor U2847 (N_2847,N_2098,N_2359);
xnor U2848 (N_2848,N_2205,N_2073);
nor U2849 (N_2849,N_2037,N_2332);
and U2850 (N_2850,N_2406,N_2307);
or U2851 (N_2851,N_2372,N_2218);
nor U2852 (N_2852,N_2379,N_2205);
nor U2853 (N_2853,N_2388,N_2137);
or U2854 (N_2854,N_2008,N_2248);
or U2855 (N_2855,N_2329,N_2248);
or U2856 (N_2856,N_2496,N_2265);
nand U2857 (N_2857,N_2233,N_2384);
or U2858 (N_2858,N_2288,N_2189);
nor U2859 (N_2859,N_2219,N_2049);
or U2860 (N_2860,N_2389,N_2246);
nand U2861 (N_2861,N_2310,N_2371);
and U2862 (N_2862,N_2457,N_2287);
nor U2863 (N_2863,N_2236,N_2318);
and U2864 (N_2864,N_2146,N_2430);
or U2865 (N_2865,N_2467,N_2213);
nand U2866 (N_2866,N_2442,N_2495);
and U2867 (N_2867,N_2309,N_2087);
or U2868 (N_2868,N_2109,N_2089);
and U2869 (N_2869,N_2102,N_2128);
nand U2870 (N_2870,N_2294,N_2205);
and U2871 (N_2871,N_2078,N_2342);
nand U2872 (N_2872,N_2375,N_2209);
or U2873 (N_2873,N_2271,N_2473);
or U2874 (N_2874,N_2122,N_2029);
or U2875 (N_2875,N_2494,N_2469);
nor U2876 (N_2876,N_2317,N_2345);
and U2877 (N_2877,N_2012,N_2303);
nand U2878 (N_2878,N_2231,N_2405);
nand U2879 (N_2879,N_2383,N_2416);
nand U2880 (N_2880,N_2030,N_2436);
nand U2881 (N_2881,N_2182,N_2103);
and U2882 (N_2882,N_2181,N_2242);
or U2883 (N_2883,N_2190,N_2170);
nor U2884 (N_2884,N_2491,N_2449);
nor U2885 (N_2885,N_2306,N_2160);
nand U2886 (N_2886,N_2064,N_2399);
and U2887 (N_2887,N_2444,N_2017);
and U2888 (N_2888,N_2057,N_2235);
or U2889 (N_2889,N_2261,N_2442);
xnor U2890 (N_2890,N_2110,N_2062);
or U2891 (N_2891,N_2359,N_2204);
or U2892 (N_2892,N_2101,N_2135);
and U2893 (N_2893,N_2436,N_2181);
and U2894 (N_2894,N_2206,N_2407);
or U2895 (N_2895,N_2054,N_2251);
or U2896 (N_2896,N_2425,N_2319);
nor U2897 (N_2897,N_2021,N_2358);
or U2898 (N_2898,N_2108,N_2185);
and U2899 (N_2899,N_2488,N_2049);
or U2900 (N_2900,N_2056,N_2331);
nor U2901 (N_2901,N_2473,N_2018);
nand U2902 (N_2902,N_2396,N_2150);
nor U2903 (N_2903,N_2244,N_2329);
and U2904 (N_2904,N_2383,N_2286);
nor U2905 (N_2905,N_2313,N_2403);
nand U2906 (N_2906,N_2258,N_2451);
or U2907 (N_2907,N_2166,N_2220);
and U2908 (N_2908,N_2027,N_2029);
and U2909 (N_2909,N_2184,N_2127);
or U2910 (N_2910,N_2321,N_2003);
nand U2911 (N_2911,N_2001,N_2355);
and U2912 (N_2912,N_2129,N_2372);
and U2913 (N_2913,N_2023,N_2086);
nand U2914 (N_2914,N_2050,N_2367);
and U2915 (N_2915,N_2200,N_2164);
and U2916 (N_2916,N_2085,N_2223);
or U2917 (N_2917,N_2303,N_2478);
nand U2918 (N_2918,N_2292,N_2440);
nand U2919 (N_2919,N_2172,N_2474);
nand U2920 (N_2920,N_2299,N_2339);
or U2921 (N_2921,N_2251,N_2366);
nand U2922 (N_2922,N_2471,N_2298);
nand U2923 (N_2923,N_2098,N_2287);
and U2924 (N_2924,N_2484,N_2474);
and U2925 (N_2925,N_2255,N_2061);
nor U2926 (N_2926,N_2123,N_2111);
or U2927 (N_2927,N_2385,N_2298);
nor U2928 (N_2928,N_2466,N_2327);
and U2929 (N_2929,N_2475,N_2008);
nand U2930 (N_2930,N_2302,N_2181);
nand U2931 (N_2931,N_2286,N_2241);
or U2932 (N_2932,N_2010,N_2446);
or U2933 (N_2933,N_2193,N_2016);
nor U2934 (N_2934,N_2124,N_2078);
or U2935 (N_2935,N_2398,N_2013);
and U2936 (N_2936,N_2083,N_2185);
or U2937 (N_2937,N_2200,N_2010);
nand U2938 (N_2938,N_2379,N_2372);
or U2939 (N_2939,N_2370,N_2453);
nor U2940 (N_2940,N_2140,N_2336);
xor U2941 (N_2941,N_2204,N_2395);
xor U2942 (N_2942,N_2051,N_2011);
and U2943 (N_2943,N_2234,N_2493);
nor U2944 (N_2944,N_2018,N_2348);
and U2945 (N_2945,N_2345,N_2336);
nor U2946 (N_2946,N_2133,N_2294);
or U2947 (N_2947,N_2109,N_2249);
nor U2948 (N_2948,N_2175,N_2171);
nand U2949 (N_2949,N_2104,N_2303);
and U2950 (N_2950,N_2004,N_2347);
nand U2951 (N_2951,N_2241,N_2264);
nor U2952 (N_2952,N_2339,N_2076);
and U2953 (N_2953,N_2044,N_2370);
nor U2954 (N_2954,N_2216,N_2407);
and U2955 (N_2955,N_2201,N_2162);
nand U2956 (N_2956,N_2162,N_2092);
nor U2957 (N_2957,N_2109,N_2073);
nand U2958 (N_2958,N_2294,N_2381);
nand U2959 (N_2959,N_2460,N_2081);
or U2960 (N_2960,N_2009,N_2165);
and U2961 (N_2961,N_2019,N_2481);
nand U2962 (N_2962,N_2077,N_2307);
nand U2963 (N_2963,N_2472,N_2281);
nand U2964 (N_2964,N_2143,N_2410);
nand U2965 (N_2965,N_2185,N_2417);
nor U2966 (N_2966,N_2396,N_2091);
or U2967 (N_2967,N_2337,N_2170);
and U2968 (N_2968,N_2310,N_2272);
or U2969 (N_2969,N_2223,N_2288);
nand U2970 (N_2970,N_2257,N_2160);
nand U2971 (N_2971,N_2257,N_2091);
and U2972 (N_2972,N_2064,N_2295);
nor U2973 (N_2973,N_2009,N_2052);
or U2974 (N_2974,N_2110,N_2016);
or U2975 (N_2975,N_2456,N_2286);
nand U2976 (N_2976,N_2111,N_2211);
nor U2977 (N_2977,N_2146,N_2041);
or U2978 (N_2978,N_2457,N_2209);
or U2979 (N_2979,N_2140,N_2329);
or U2980 (N_2980,N_2102,N_2219);
and U2981 (N_2981,N_2006,N_2191);
nor U2982 (N_2982,N_2478,N_2165);
nor U2983 (N_2983,N_2375,N_2269);
or U2984 (N_2984,N_2186,N_2022);
xnor U2985 (N_2985,N_2166,N_2245);
nand U2986 (N_2986,N_2396,N_2040);
and U2987 (N_2987,N_2291,N_2282);
and U2988 (N_2988,N_2168,N_2394);
or U2989 (N_2989,N_2406,N_2088);
nand U2990 (N_2990,N_2395,N_2076);
nor U2991 (N_2991,N_2225,N_2309);
or U2992 (N_2992,N_2141,N_2440);
and U2993 (N_2993,N_2316,N_2143);
or U2994 (N_2994,N_2416,N_2147);
and U2995 (N_2995,N_2054,N_2351);
and U2996 (N_2996,N_2271,N_2106);
nand U2997 (N_2997,N_2431,N_2025);
nor U2998 (N_2998,N_2091,N_2486);
xnor U2999 (N_2999,N_2298,N_2294);
and U3000 (N_3000,N_2777,N_2548);
and U3001 (N_3001,N_2900,N_2963);
xor U3002 (N_3002,N_2671,N_2753);
and U3003 (N_3003,N_2829,N_2999);
nor U3004 (N_3004,N_2534,N_2692);
nor U3005 (N_3005,N_2870,N_2518);
nand U3006 (N_3006,N_2970,N_2511);
nand U3007 (N_3007,N_2883,N_2683);
or U3008 (N_3008,N_2682,N_2556);
or U3009 (N_3009,N_2551,N_2721);
nor U3010 (N_3010,N_2539,N_2737);
nand U3011 (N_3011,N_2642,N_2506);
or U3012 (N_3012,N_2908,N_2543);
or U3013 (N_3013,N_2526,N_2693);
nand U3014 (N_3014,N_2756,N_2665);
or U3015 (N_3015,N_2815,N_2795);
and U3016 (N_3016,N_2869,N_2765);
and U3017 (N_3017,N_2858,N_2610);
xor U3018 (N_3018,N_2647,N_2750);
or U3019 (N_3019,N_2638,N_2819);
and U3020 (N_3020,N_2565,N_2961);
nand U3021 (N_3021,N_2586,N_2615);
or U3022 (N_3022,N_2987,N_2505);
and U3023 (N_3023,N_2764,N_2664);
nor U3024 (N_3024,N_2790,N_2824);
and U3025 (N_3025,N_2997,N_2748);
or U3026 (N_3026,N_2798,N_2724);
nand U3027 (N_3027,N_2668,N_2516);
and U3028 (N_3028,N_2532,N_2677);
and U3029 (N_3029,N_2949,N_2744);
and U3030 (N_3030,N_2743,N_2656);
nor U3031 (N_3031,N_2923,N_2805);
or U3032 (N_3032,N_2713,N_2901);
nand U3033 (N_3033,N_2742,N_2546);
nand U3034 (N_3034,N_2995,N_2857);
and U3035 (N_3035,N_2754,N_2891);
or U3036 (N_3036,N_2809,N_2818);
nor U3037 (N_3037,N_2909,N_2731);
and U3038 (N_3038,N_2928,N_2855);
or U3039 (N_3039,N_2527,N_2609);
or U3040 (N_3040,N_2813,N_2884);
nand U3041 (N_3041,N_2710,N_2956);
nand U3042 (N_3042,N_2968,N_2902);
nor U3043 (N_3043,N_2852,N_2853);
nand U3044 (N_3044,N_2559,N_2567);
nor U3045 (N_3045,N_2926,N_2655);
or U3046 (N_3046,N_2627,N_2689);
or U3047 (N_3047,N_2550,N_2931);
nand U3048 (N_3048,N_2581,N_2728);
nand U3049 (N_3049,N_2604,N_2579);
and U3050 (N_3050,N_2585,N_2629);
or U3051 (N_3051,N_2593,N_2797);
nor U3052 (N_3052,N_2603,N_2502);
or U3053 (N_3053,N_2879,N_2538);
or U3054 (N_3054,N_2739,N_2924);
or U3055 (N_3055,N_2760,N_2523);
or U3056 (N_3056,N_2938,N_2957);
and U3057 (N_3057,N_2821,N_2934);
nand U3058 (N_3058,N_2566,N_2962);
nand U3059 (N_3059,N_2597,N_2633);
nand U3060 (N_3060,N_2769,N_2907);
or U3061 (N_3061,N_2639,N_2948);
nor U3062 (N_3062,N_2835,N_2899);
or U3063 (N_3063,N_2568,N_2555);
or U3064 (N_3064,N_2872,N_2787);
and U3065 (N_3065,N_2802,N_2998);
nand U3066 (N_3066,N_2904,N_2657);
or U3067 (N_3067,N_2670,N_2807);
nor U3068 (N_3068,N_2833,N_2770);
nand U3069 (N_3069,N_2861,N_2732);
and U3070 (N_3070,N_2828,N_2782);
nor U3071 (N_3071,N_2822,N_2911);
nand U3072 (N_3072,N_2827,N_2906);
and U3073 (N_3073,N_2868,N_2529);
nor U3074 (N_3074,N_2594,N_2661);
or U3075 (N_3075,N_2783,N_2605);
nand U3076 (N_3076,N_2607,N_2560);
nand U3077 (N_3077,N_2952,N_2501);
nand U3078 (N_3078,N_2662,N_2613);
or U3079 (N_3079,N_2549,N_2836);
nor U3080 (N_3080,N_2755,N_2576);
and U3081 (N_3081,N_2838,N_2940);
or U3082 (N_3082,N_2658,N_2981);
or U3083 (N_3083,N_2542,N_2706);
or U3084 (N_3084,N_2977,N_2942);
or U3085 (N_3085,N_2601,N_2767);
nand U3086 (N_3086,N_2722,N_2793);
and U3087 (N_3087,N_2641,N_2735);
nand U3088 (N_3088,N_2915,N_2863);
or U3089 (N_3089,N_2707,N_2619);
nand U3090 (N_3090,N_2644,N_2704);
nor U3091 (N_3091,N_2975,N_2740);
nand U3092 (N_3092,N_2958,N_2719);
and U3093 (N_3093,N_2686,N_2696);
or U3094 (N_3094,N_2986,N_2898);
or U3095 (N_3095,N_2843,N_2877);
or U3096 (N_3096,N_2894,N_2602);
xnor U3097 (N_3097,N_2687,N_2826);
or U3098 (N_3098,N_2561,N_2959);
nor U3099 (N_3099,N_2606,N_2889);
and U3100 (N_3100,N_2752,N_2660);
nand U3101 (N_3101,N_2648,N_2955);
nand U3102 (N_3102,N_2759,N_2984);
nor U3103 (N_3103,N_2749,N_2508);
nand U3104 (N_3104,N_2530,N_2563);
and U3105 (N_3105,N_2745,N_2634);
nor U3106 (N_3106,N_2751,N_2834);
nand U3107 (N_3107,N_2705,N_2544);
nor U3108 (N_3108,N_2941,N_2669);
and U3109 (N_3109,N_2831,N_2932);
or U3110 (N_3110,N_2637,N_2645);
nor U3111 (N_3111,N_2935,N_2509);
nand U3112 (N_3112,N_2564,N_2982);
nor U3113 (N_3113,N_2659,N_2865);
and U3114 (N_3114,N_2874,N_2771);
nor U3115 (N_3115,N_2845,N_2587);
nand U3116 (N_3116,N_2575,N_2806);
or U3117 (N_3117,N_2896,N_2557);
nor U3118 (N_3118,N_2810,N_2608);
or U3119 (N_3119,N_2700,N_2875);
or U3120 (N_3120,N_2703,N_2685);
or U3121 (N_3121,N_2763,N_2800);
nor U3122 (N_3122,N_2622,N_2712);
xor U3123 (N_3123,N_2730,N_2903);
and U3124 (N_3124,N_2667,N_2890);
and U3125 (N_3125,N_2631,N_2570);
and U3126 (N_3126,N_2988,N_2572);
or U3127 (N_3127,N_2723,N_2596);
or U3128 (N_3128,N_2734,N_2794);
nor U3129 (N_3129,N_2533,N_2621);
nand U3130 (N_3130,N_2599,N_2515);
nor U3131 (N_3131,N_2729,N_2580);
nand U3132 (N_3132,N_2673,N_2913);
nand U3133 (N_3133,N_2577,N_2727);
nand U3134 (N_3134,N_2878,N_2573);
nor U3135 (N_3135,N_2578,N_2820);
or U3136 (N_3136,N_2880,N_2652);
nor U3137 (N_3137,N_2611,N_2620);
or U3138 (N_3138,N_2983,N_2781);
and U3139 (N_3139,N_2702,N_2676);
nand U3140 (N_3140,N_2552,N_2985);
and U3141 (N_3141,N_2646,N_2851);
nand U3142 (N_3142,N_2953,N_2943);
and U3143 (N_3143,N_2640,N_2757);
and U3144 (N_3144,N_2643,N_2929);
nor U3145 (N_3145,N_2974,N_2690);
nor U3146 (N_3146,N_2967,N_2849);
or U3147 (N_3147,N_2892,N_2814);
nand U3148 (N_3148,N_2583,N_2680);
or U3149 (N_3149,N_2914,N_2918);
nor U3150 (N_3150,N_2698,N_2993);
and U3151 (N_3151,N_2947,N_2653);
and U3152 (N_3152,N_2830,N_2871);
nor U3153 (N_3153,N_2626,N_2916);
and U3154 (N_3154,N_2775,N_2888);
or U3155 (N_3155,N_2697,N_2589);
nor U3156 (N_3156,N_2558,N_2684);
and U3157 (N_3157,N_2571,N_2945);
nand U3158 (N_3158,N_2545,N_2796);
nor U3159 (N_3159,N_2972,N_2786);
nor U3160 (N_3160,N_2925,N_2715);
nand U3161 (N_3161,N_2873,N_2514);
nor U3162 (N_3162,N_2950,N_2996);
and U3163 (N_3163,N_2741,N_2688);
nand U3164 (N_3164,N_2854,N_2699);
nor U3165 (N_3165,N_2582,N_2649);
nand U3166 (N_3166,N_2847,N_2841);
or U3167 (N_3167,N_2994,N_2960);
and U3168 (N_3168,N_2716,N_2618);
or U3169 (N_3169,N_2776,N_2848);
nor U3170 (N_3170,N_2992,N_2537);
nor U3171 (N_3171,N_2635,N_2939);
or U3172 (N_3172,N_2791,N_2973);
and U3173 (N_3173,N_2708,N_2825);
or U3174 (N_3174,N_2823,N_2976);
nand U3175 (N_3175,N_2636,N_2524);
xnor U3176 (N_3176,N_2864,N_2584);
nor U3177 (N_3177,N_2691,N_2846);
or U3178 (N_3178,N_2844,N_2562);
and U3179 (N_3179,N_2746,N_2917);
nand U3180 (N_3180,N_2991,N_2927);
nand U3181 (N_3181,N_2630,N_2905);
and U3182 (N_3182,N_2886,N_2598);
nor U3183 (N_3183,N_2758,N_2885);
and U3184 (N_3184,N_2614,N_2535);
and U3185 (N_3185,N_2531,N_2522);
xor U3186 (N_3186,N_2859,N_2681);
or U3187 (N_3187,N_2651,N_2921);
or U3188 (N_3188,N_2574,N_2547);
or U3189 (N_3189,N_2674,N_2937);
nand U3190 (N_3190,N_2517,N_2979);
and U3191 (N_3191,N_2540,N_2792);
nor U3192 (N_3192,N_2964,N_2816);
and U3193 (N_3193,N_2591,N_2966);
or U3194 (N_3194,N_2897,N_2616);
and U3195 (N_3195,N_2788,N_2808);
nand U3196 (N_3196,N_2612,N_2856);
nand U3197 (N_3197,N_2837,N_2553);
and U3198 (N_3198,N_2528,N_2842);
and U3199 (N_3199,N_2701,N_2801);
nor U3200 (N_3200,N_2720,N_2588);
nor U3201 (N_3201,N_2774,N_2717);
or U3202 (N_3202,N_2711,N_2628);
nand U3203 (N_3203,N_2772,N_2840);
or U3204 (N_3204,N_2910,N_2590);
nor U3205 (N_3205,N_2541,N_2980);
nand U3206 (N_3206,N_2778,N_2920);
nand U3207 (N_3207,N_2866,N_2679);
nor U3208 (N_3208,N_2632,N_2784);
nor U3209 (N_3209,N_2512,N_2922);
nor U3210 (N_3210,N_2850,N_2832);
nor U3211 (N_3211,N_2503,N_2990);
or U3212 (N_3212,N_2623,N_2695);
nor U3213 (N_3213,N_2675,N_2978);
nand U3214 (N_3214,N_2663,N_2617);
and U3215 (N_3215,N_2860,N_2747);
or U3216 (N_3216,N_2803,N_2694);
nor U3217 (N_3217,N_2804,N_2881);
nand U3218 (N_3218,N_2507,N_2882);
nand U3219 (N_3219,N_2650,N_2504);
and U3220 (N_3220,N_2733,N_2600);
nand U3221 (N_3221,N_2785,N_2519);
nand U3222 (N_3222,N_2789,N_2965);
nor U3223 (N_3223,N_2624,N_2933);
nor U3224 (N_3224,N_2989,N_2817);
and U3225 (N_3225,N_2736,N_2500);
and U3226 (N_3226,N_2766,N_2761);
nor U3227 (N_3227,N_2862,N_2672);
nand U3228 (N_3228,N_2520,N_2811);
nand U3229 (N_3229,N_2887,N_2536);
nand U3230 (N_3230,N_2554,N_2678);
or U3231 (N_3231,N_2510,N_2919);
nor U3232 (N_3232,N_2595,N_2625);
nor U3233 (N_3233,N_2944,N_2930);
nand U3234 (N_3234,N_2971,N_2936);
or U3235 (N_3235,N_2654,N_2521);
or U3236 (N_3236,N_2780,N_2954);
nor U3237 (N_3237,N_2569,N_2709);
nand U3238 (N_3238,N_2799,N_2592);
and U3239 (N_3239,N_2839,N_2912);
and U3240 (N_3240,N_2876,N_2525);
nand U3241 (N_3241,N_2779,N_2762);
or U3242 (N_3242,N_2812,N_2895);
nand U3243 (N_3243,N_2726,N_2768);
nor U3244 (N_3244,N_2773,N_2951);
nor U3245 (N_3245,N_2867,N_2666);
and U3246 (N_3246,N_2714,N_2725);
nor U3247 (N_3247,N_2513,N_2946);
and U3248 (N_3248,N_2893,N_2718);
and U3249 (N_3249,N_2738,N_2969);
or U3250 (N_3250,N_2794,N_2776);
and U3251 (N_3251,N_2939,N_2593);
and U3252 (N_3252,N_2593,N_2500);
and U3253 (N_3253,N_2835,N_2607);
nor U3254 (N_3254,N_2774,N_2557);
nor U3255 (N_3255,N_2897,N_2829);
nor U3256 (N_3256,N_2890,N_2788);
nor U3257 (N_3257,N_2807,N_2596);
nor U3258 (N_3258,N_2820,N_2966);
nor U3259 (N_3259,N_2677,N_2880);
nor U3260 (N_3260,N_2633,N_2772);
or U3261 (N_3261,N_2507,N_2627);
or U3262 (N_3262,N_2868,N_2946);
nand U3263 (N_3263,N_2811,N_2808);
or U3264 (N_3264,N_2599,N_2955);
nor U3265 (N_3265,N_2873,N_2669);
and U3266 (N_3266,N_2793,N_2586);
nor U3267 (N_3267,N_2835,N_2834);
nor U3268 (N_3268,N_2623,N_2923);
nor U3269 (N_3269,N_2876,N_2637);
nand U3270 (N_3270,N_2555,N_2957);
nor U3271 (N_3271,N_2969,N_2789);
nand U3272 (N_3272,N_2621,N_2687);
and U3273 (N_3273,N_2937,N_2627);
and U3274 (N_3274,N_2791,N_2553);
nand U3275 (N_3275,N_2635,N_2751);
nand U3276 (N_3276,N_2942,N_2782);
or U3277 (N_3277,N_2980,N_2593);
or U3278 (N_3278,N_2838,N_2586);
and U3279 (N_3279,N_2565,N_2778);
and U3280 (N_3280,N_2600,N_2942);
xor U3281 (N_3281,N_2892,N_2738);
or U3282 (N_3282,N_2942,N_2744);
nand U3283 (N_3283,N_2952,N_2899);
xnor U3284 (N_3284,N_2679,N_2807);
or U3285 (N_3285,N_2603,N_2539);
and U3286 (N_3286,N_2565,N_2962);
and U3287 (N_3287,N_2974,N_2665);
nor U3288 (N_3288,N_2508,N_2668);
or U3289 (N_3289,N_2938,N_2862);
and U3290 (N_3290,N_2959,N_2941);
or U3291 (N_3291,N_2971,N_2839);
nor U3292 (N_3292,N_2733,N_2761);
nor U3293 (N_3293,N_2626,N_2817);
and U3294 (N_3294,N_2619,N_2539);
or U3295 (N_3295,N_2786,N_2695);
or U3296 (N_3296,N_2652,N_2940);
nor U3297 (N_3297,N_2624,N_2785);
and U3298 (N_3298,N_2870,N_2780);
nor U3299 (N_3299,N_2597,N_2961);
nand U3300 (N_3300,N_2578,N_2961);
and U3301 (N_3301,N_2983,N_2952);
or U3302 (N_3302,N_2994,N_2959);
nand U3303 (N_3303,N_2702,N_2535);
or U3304 (N_3304,N_2703,N_2864);
or U3305 (N_3305,N_2527,N_2706);
nand U3306 (N_3306,N_2886,N_2546);
nand U3307 (N_3307,N_2964,N_2719);
nand U3308 (N_3308,N_2911,N_2971);
nor U3309 (N_3309,N_2551,N_2539);
or U3310 (N_3310,N_2522,N_2954);
and U3311 (N_3311,N_2516,N_2545);
nand U3312 (N_3312,N_2786,N_2597);
nand U3313 (N_3313,N_2877,N_2572);
nor U3314 (N_3314,N_2643,N_2649);
or U3315 (N_3315,N_2883,N_2687);
nor U3316 (N_3316,N_2741,N_2511);
or U3317 (N_3317,N_2609,N_2709);
nor U3318 (N_3318,N_2589,N_2648);
and U3319 (N_3319,N_2861,N_2899);
and U3320 (N_3320,N_2533,N_2818);
nand U3321 (N_3321,N_2703,N_2705);
nand U3322 (N_3322,N_2674,N_2617);
nor U3323 (N_3323,N_2923,N_2516);
and U3324 (N_3324,N_2991,N_2896);
nand U3325 (N_3325,N_2938,N_2889);
and U3326 (N_3326,N_2865,N_2884);
or U3327 (N_3327,N_2932,N_2719);
nand U3328 (N_3328,N_2758,N_2634);
or U3329 (N_3329,N_2744,N_2785);
nand U3330 (N_3330,N_2532,N_2771);
and U3331 (N_3331,N_2613,N_2501);
or U3332 (N_3332,N_2754,N_2513);
nor U3333 (N_3333,N_2596,N_2726);
nand U3334 (N_3334,N_2949,N_2988);
or U3335 (N_3335,N_2896,N_2830);
or U3336 (N_3336,N_2887,N_2976);
nand U3337 (N_3337,N_2923,N_2607);
nor U3338 (N_3338,N_2570,N_2818);
nor U3339 (N_3339,N_2892,N_2931);
or U3340 (N_3340,N_2747,N_2548);
and U3341 (N_3341,N_2773,N_2668);
and U3342 (N_3342,N_2573,N_2908);
nand U3343 (N_3343,N_2502,N_2818);
nand U3344 (N_3344,N_2817,N_2528);
nand U3345 (N_3345,N_2986,N_2867);
nand U3346 (N_3346,N_2793,N_2644);
nand U3347 (N_3347,N_2983,N_2736);
or U3348 (N_3348,N_2718,N_2930);
nand U3349 (N_3349,N_2955,N_2888);
nand U3350 (N_3350,N_2897,N_2899);
or U3351 (N_3351,N_2527,N_2512);
or U3352 (N_3352,N_2604,N_2874);
or U3353 (N_3353,N_2969,N_2821);
or U3354 (N_3354,N_2714,N_2915);
nor U3355 (N_3355,N_2522,N_2500);
nand U3356 (N_3356,N_2909,N_2727);
and U3357 (N_3357,N_2574,N_2720);
nor U3358 (N_3358,N_2780,N_2583);
nor U3359 (N_3359,N_2957,N_2604);
or U3360 (N_3360,N_2727,N_2633);
nand U3361 (N_3361,N_2878,N_2662);
nand U3362 (N_3362,N_2909,N_2918);
nor U3363 (N_3363,N_2530,N_2540);
or U3364 (N_3364,N_2601,N_2973);
nand U3365 (N_3365,N_2829,N_2736);
or U3366 (N_3366,N_2924,N_2838);
and U3367 (N_3367,N_2587,N_2860);
or U3368 (N_3368,N_2798,N_2568);
and U3369 (N_3369,N_2585,N_2775);
or U3370 (N_3370,N_2826,N_2870);
and U3371 (N_3371,N_2724,N_2947);
and U3372 (N_3372,N_2802,N_2573);
and U3373 (N_3373,N_2817,N_2820);
nand U3374 (N_3374,N_2877,N_2781);
and U3375 (N_3375,N_2580,N_2652);
nand U3376 (N_3376,N_2806,N_2588);
nor U3377 (N_3377,N_2597,N_2739);
and U3378 (N_3378,N_2660,N_2926);
and U3379 (N_3379,N_2700,N_2976);
nand U3380 (N_3380,N_2764,N_2680);
or U3381 (N_3381,N_2677,N_2984);
or U3382 (N_3382,N_2881,N_2843);
or U3383 (N_3383,N_2806,N_2886);
and U3384 (N_3384,N_2731,N_2984);
and U3385 (N_3385,N_2988,N_2990);
and U3386 (N_3386,N_2858,N_2714);
and U3387 (N_3387,N_2558,N_2854);
and U3388 (N_3388,N_2722,N_2544);
and U3389 (N_3389,N_2936,N_2991);
nor U3390 (N_3390,N_2546,N_2585);
nand U3391 (N_3391,N_2915,N_2558);
or U3392 (N_3392,N_2820,N_2976);
nand U3393 (N_3393,N_2583,N_2534);
or U3394 (N_3394,N_2705,N_2894);
and U3395 (N_3395,N_2507,N_2819);
and U3396 (N_3396,N_2707,N_2628);
or U3397 (N_3397,N_2871,N_2506);
nor U3398 (N_3398,N_2805,N_2853);
nand U3399 (N_3399,N_2561,N_2654);
and U3400 (N_3400,N_2975,N_2755);
or U3401 (N_3401,N_2851,N_2570);
nand U3402 (N_3402,N_2987,N_2848);
or U3403 (N_3403,N_2772,N_2930);
and U3404 (N_3404,N_2593,N_2528);
and U3405 (N_3405,N_2821,N_2650);
nor U3406 (N_3406,N_2957,N_2688);
or U3407 (N_3407,N_2824,N_2832);
or U3408 (N_3408,N_2943,N_2659);
xor U3409 (N_3409,N_2963,N_2638);
nand U3410 (N_3410,N_2677,N_2535);
nand U3411 (N_3411,N_2802,N_2800);
nor U3412 (N_3412,N_2565,N_2568);
nor U3413 (N_3413,N_2927,N_2660);
or U3414 (N_3414,N_2987,N_2867);
or U3415 (N_3415,N_2740,N_2515);
nand U3416 (N_3416,N_2666,N_2869);
nor U3417 (N_3417,N_2753,N_2963);
or U3418 (N_3418,N_2682,N_2618);
and U3419 (N_3419,N_2821,N_2713);
and U3420 (N_3420,N_2783,N_2679);
nand U3421 (N_3421,N_2900,N_2856);
or U3422 (N_3422,N_2539,N_2925);
and U3423 (N_3423,N_2954,N_2971);
and U3424 (N_3424,N_2892,N_2964);
nand U3425 (N_3425,N_2766,N_2774);
or U3426 (N_3426,N_2910,N_2891);
nand U3427 (N_3427,N_2537,N_2585);
and U3428 (N_3428,N_2758,N_2734);
or U3429 (N_3429,N_2602,N_2560);
and U3430 (N_3430,N_2572,N_2518);
or U3431 (N_3431,N_2566,N_2764);
nand U3432 (N_3432,N_2848,N_2678);
nand U3433 (N_3433,N_2882,N_2856);
nor U3434 (N_3434,N_2685,N_2538);
nor U3435 (N_3435,N_2656,N_2883);
nor U3436 (N_3436,N_2838,N_2720);
and U3437 (N_3437,N_2711,N_2876);
nor U3438 (N_3438,N_2639,N_2554);
nor U3439 (N_3439,N_2948,N_2519);
nor U3440 (N_3440,N_2802,N_2746);
nand U3441 (N_3441,N_2771,N_2941);
nor U3442 (N_3442,N_2587,N_2673);
and U3443 (N_3443,N_2808,N_2688);
nor U3444 (N_3444,N_2782,N_2644);
or U3445 (N_3445,N_2747,N_2631);
or U3446 (N_3446,N_2969,N_2924);
xor U3447 (N_3447,N_2892,N_2990);
nor U3448 (N_3448,N_2982,N_2782);
or U3449 (N_3449,N_2609,N_2846);
and U3450 (N_3450,N_2851,N_2516);
nand U3451 (N_3451,N_2859,N_2770);
nand U3452 (N_3452,N_2910,N_2818);
nor U3453 (N_3453,N_2760,N_2733);
or U3454 (N_3454,N_2710,N_2762);
nand U3455 (N_3455,N_2599,N_2526);
nand U3456 (N_3456,N_2810,N_2513);
or U3457 (N_3457,N_2759,N_2880);
or U3458 (N_3458,N_2645,N_2619);
nand U3459 (N_3459,N_2608,N_2986);
nand U3460 (N_3460,N_2549,N_2542);
nand U3461 (N_3461,N_2967,N_2546);
nand U3462 (N_3462,N_2904,N_2954);
and U3463 (N_3463,N_2775,N_2958);
and U3464 (N_3464,N_2806,N_2876);
and U3465 (N_3465,N_2936,N_2981);
or U3466 (N_3466,N_2651,N_2702);
or U3467 (N_3467,N_2535,N_2760);
nor U3468 (N_3468,N_2529,N_2501);
and U3469 (N_3469,N_2924,N_2760);
or U3470 (N_3470,N_2638,N_2719);
or U3471 (N_3471,N_2508,N_2929);
and U3472 (N_3472,N_2616,N_2895);
and U3473 (N_3473,N_2641,N_2726);
and U3474 (N_3474,N_2654,N_2756);
nand U3475 (N_3475,N_2649,N_2682);
or U3476 (N_3476,N_2894,N_2814);
and U3477 (N_3477,N_2603,N_2571);
and U3478 (N_3478,N_2787,N_2648);
nand U3479 (N_3479,N_2913,N_2868);
nor U3480 (N_3480,N_2938,N_2650);
nor U3481 (N_3481,N_2946,N_2659);
nand U3482 (N_3482,N_2989,N_2879);
and U3483 (N_3483,N_2957,N_2659);
nor U3484 (N_3484,N_2649,N_2901);
or U3485 (N_3485,N_2571,N_2773);
or U3486 (N_3486,N_2974,N_2751);
and U3487 (N_3487,N_2517,N_2922);
and U3488 (N_3488,N_2958,N_2808);
nor U3489 (N_3489,N_2701,N_2915);
and U3490 (N_3490,N_2609,N_2572);
nor U3491 (N_3491,N_2919,N_2953);
or U3492 (N_3492,N_2763,N_2872);
and U3493 (N_3493,N_2781,N_2890);
nand U3494 (N_3494,N_2816,N_2593);
or U3495 (N_3495,N_2718,N_2564);
nor U3496 (N_3496,N_2674,N_2514);
nor U3497 (N_3497,N_2573,N_2997);
nor U3498 (N_3498,N_2973,N_2762);
nand U3499 (N_3499,N_2989,N_2963);
nor U3500 (N_3500,N_3083,N_3472);
and U3501 (N_3501,N_3096,N_3322);
or U3502 (N_3502,N_3396,N_3140);
or U3503 (N_3503,N_3289,N_3249);
and U3504 (N_3504,N_3199,N_3226);
and U3505 (N_3505,N_3086,N_3484);
and U3506 (N_3506,N_3463,N_3369);
or U3507 (N_3507,N_3332,N_3297);
nor U3508 (N_3508,N_3153,N_3216);
or U3509 (N_3509,N_3097,N_3033);
and U3510 (N_3510,N_3327,N_3209);
nand U3511 (N_3511,N_3161,N_3459);
nand U3512 (N_3512,N_3383,N_3326);
nor U3513 (N_3513,N_3169,N_3093);
and U3514 (N_3514,N_3107,N_3349);
nand U3515 (N_3515,N_3134,N_3353);
and U3516 (N_3516,N_3448,N_3423);
nor U3517 (N_3517,N_3218,N_3208);
nor U3518 (N_3518,N_3432,N_3178);
nand U3519 (N_3519,N_3317,N_3422);
or U3520 (N_3520,N_3409,N_3241);
and U3521 (N_3521,N_3010,N_3379);
nand U3522 (N_3522,N_3110,N_3399);
or U3523 (N_3523,N_3125,N_3386);
and U3524 (N_3524,N_3136,N_3228);
nor U3525 (N_3525,N_3024,N_3334);
nor U3526 (N_3526,N_3306,N_3478);
nand U3527 (N_3527,N_3293,N_3382);
nand U3528 (N_3528,N_3048,N_3047);
and U3529 (N_3529,N_3470,N_3286);
and U3530 (N_3530,N_3115,N_3407);
and U3531 (N_3531,N_3489,N_3338);
or U3532 (N_3532,N_3028,N_3112);
nand U3533 (N_3533,N_3066,N_3159);
or U3534 (N_3534,N_3363,N_3356);
and U3535 (N_3535,N_3064,N_3273);
nor U3536 (N_3536,N_3251,N_3189);
or U3537 (N_3537,N_3416,N_3256);
and U3538 (N_3538,N_3079,N_3271);
nand U3539 (N_3539,N_3468,N_3390);
and U3540 (N_3540,N_3045,N_3281);
nand U3541 (N_3541,N_3277,N_3344);
and U3542 (N_3542,N_3258,N_3185);
nor U3543 (N_3543,N_3290,N_3425);
nor U3544 (N_3544,N_3156,N_3476);
and U3545 (N_3545,N_3205,N_3458);
or U3546 (N_3546,N_3405,N_3137);
or U3547 (N_3547,N_3479,N_3165);
and U3548 (N_3548,N_3133,N_3167);
or U3549 (N_3549,N_3378,N_3352);
nor U3550 (N_3550,N_3291,N_3447);
nor U3551 (N_3551,N_3138,N_3487);
nand U3552 (N_3552,N_3375,N_3454);
and U3553 (N_3553,N_3203,N_3032);
nand U3554 (N_3554,N_3320,N_3077);
nor U3555 (N_3555,N_3410,N_3401);
and U3556 (N_3556,N_3460,N_3308);
and U3557 (N_3557,N_3295,N_3151);
nand U3558 (N_3558,N_3054,N_3359);
and U3559 (N_3559,N_3044,N_3452);
nand U3560 (N_3560,N_3239,N_3019);
and U3561 (N_3561,N_3182,N_3337);
nand U3562 (N_3562,N_3069,N_3051);
or U3563 (N_3563,N_3393,N_3157);
and U3564 (N_3564,N_3309,N_3466);
nor U3565 (N_3565,N_3365,N_3127);
or U3566 (N_3566,N_3074,N_3380);
and U3567 (N_3567,N_3457,N_3003);
and U3568 (N_3568,N_3229,N_3499);
nand U3569 (N_3569,N_3296,N_3259);
nand U3570 (N_3570,N_3341,N_3419);
or U3571 (N_3571,N_3040,N_3105);
nor U3572 (N_3572,N_3493,N_3202);
and U3573 (N_3573,N_3328,N_3148);
or U3574 (N_3574,N_3065,N_3438);
nor U3575 (N_3575,N_3494,N_3404);
or U3576 (N_3576,N_3323,N_3307);
and U3577 (N_3577,N_3408,N_3310);
and U3578 (N_3578,N_3444,N_3374);
and U3579 (N_3579,N_3158,N_3449);
and U3580 (N_3580,N_3222,N_3418);
nor U3581 (N_3581,N_3498,N_3397);
nor U3582 (N_3582,N_3465,N_3053);
or U3583 (N_3583,N_3160,N_3321);
nand U3584 (N_3584,N_3362,N_3385);
nor U3585 (N_3585,N_3100,N_3283);
xnor U3586 (N_3586,N_3084,N_3442);
and U3587 (N_3587,N_3145,N_3340);
nor U3588 (N_3588,N_3435,N_3485);
nand U3589 (N_3589,N_3453,N_3068);
and U3590 (N_3590,N_3123,N_3347);
nor U3591 (N_3591,N_3016,N_3211);
or U3592 (N_3592,N_3031,N_3020);
nand U3593 (N_3593,N_3215,N_3173);
and U3594 (N_3594,N_3139,N_3312);
nand U3595 (N_3595,N_3092,N_3242);
nand U3596 (N_3596,N_3023,N_3276);
nand U3597 (N_3597,N_3035,N_3262);
nor U3598 (N_3598,N_3298,N_3431);
and U3599 (N_3599,N_3441,N_3147);
nand U3600 (N_3600,N_3163,N_3225);
and U3601 (N_3601,N_3252,N_3475);
and U3602 (N_3602,N_3060,N_3000);
nor U3603 (N_3603,N_3018,N_3324);
nor U3604 (N_3604,N_3261,N_3427);
nand U3605 (N_3605,N_3184,N_3109);
or U3606 (N_3606,N_3041,N_3474);
nor U3607 (N_3607,N_3336,N_3377);
and U3608 (N_3608,N_3471,N_3067);
or U3609 (N_3609,N_3063,N_3392);
nor U3610 (N_3610,N_3398,N_3126);
nand U3611 (N_3611,N_3168,N_3257);
and U3612 (N_3612,N_3196,N_3154);
nor U3613 (N_3613,N_3164,N_3070);
nand U3614 (N_3614,N_3265,N_3090);
nand U3615 (N_3615,N_3267,N_3223);
nand U3616 (N_3616,N_3001,N_3176);
nand U3617 (N_3617,N_3469,N_3017);
nand U3618 (N_3618,N_3464,N_3181);
and U3619 (N_3619,N_3108,N_3269);
or U3620 (N_3620,N_3114,N_3013);
or U3621 (N_3621,N_3279,N_3400);
and U3622 (N_3622,N_3039,N_3142);
nand U3623 (N_3623,N_3049,N_3302);
nor U3624 (N_3624,N_3343,N_3346);
nor U3625 (N_3625,N_3195,N_3091);
and U3626 (N_3626,N_3339,N_3437);
nor U3627 (N_3627,N_3434,N_3099);
or U3628 (N_3628,N_3219,N_3094);
or U3629 (N_3629,N_3187,N_3274);
and U3630 (N_3630,N_3482,N_3025);
or U3631 (N_3631,N_3287,N_3233);
nand U3632 (N_3632,N_3191,N_3333);
or U3633 (N_3633,N_3119,N_3214);
nor U3634 (N_3634,N_3008,N_3062);
nand U3635 (N_3635,N_3106,N_3305);
nor U3636 (N_3636,N_3120,N_3073);
or U3637 (N_3637,N_3411,N_3245);
nor U3638 (N_3638,N_3388,N_3179);
and U3639 (N_3639,N_3301,N_3480);
nor U3640 (N_3640,N_3194,N_3244);
or U3641 (N_3641,N_3027,N_3481);
nor U3642 (N_3642,N_3117,N_3367);
nand U3643 (N_3643,N_3443,N_3072);
and U3644 (N_3644,N_3381,N_3313);
nand U3645 (N_3645,N_3373,N_3204);
nand U3646 (N_3646,N_3217,N_3304);
nand U3647 (N_3647,N_3162,N_3420);
nand U3648 (N_3648,N_3387,N_3350);
and U3649 (N_3649,N_3080,N_3183);
and U3650 (N_3650,N_3180,N_3315);
nand U3651 (N_3651,N_3104,N_3030);
nand U3652 (N_3652,N_3103,N_3456);
and U3653 (N_3653,N_3206,N_3050);
or U3654 (N_3654,N_3412,N_3220);
or U3655 (N_3655,N_3288,N_3490);
and U3656 (N_3656,N_3175,N_3192);
and U3657 (N_3657,N_3232,N_3371);
nand U3658 (N_3658,N_3372,N_3348);
nand U3659 (N_3659,N_3282,N_3243);
or U3660 (N_3660,N_3467,N_3171);
and U3661 (N_3661,N_3015,N_3085);
and U3662 (N_3662,N_3095,N_3294);
nand U3663 (N_3663,N_3012,N_3076);
or U3664 (N_3664,N_3057,N_3201);
nor U3665 (N_3665,N_3329,N_3473);
nand U3666 (N_3666,N_3190,N_3237);
nor U3667 (N_3667,N_3355,N_3235);
nand U3668 (N_3668,N_3200,N_3414);
or U3669 (N_3669,N_3426,N_3146);
and U3670 (N_3670,N_3394,N_3421);
nor U3671 (N_3671,N_3234,N_3224);
nand U3672 (N_3672,N_3495,N_3428);
or U3673 (N_3673,N_3089,N_3197);
or U3674 (N_3674,N_3342,N_3132);
nand U3675 (N_3675,N_3250,N_3406);
nor U3676 (N_3676,N_3005,N_3056);
nor U3677 (N_3677,N_3491,N_3166);
or U3678 (N_3678,N_3430,N_3022);
nand U3679 (N_3679,N_3461,N_3021);
nand U3680 (N_3680,N_3477,N_3462);
nor U3681 (N_3681,N_3402,N_3360);
nor U3682 (N_3682,N_3436,N_3036);
nor U3683 (N_3683,N_3247,N_3177);
or U3684 (N_3684,N_3303,N_3038);
and U3685 (N_3685,N_3129,N_3121);
nand U3686 (N_3686,N_3314,N_3455);
and U3687 (N_3687,N_3440,N_3330);
nand U3688 (N_3688,N_3488,N_3088);
nand U3689 (N_3689,N_3292,N_3246);
and U3690 (N_3690,N_3345,N_3361);
or U3691 (N_3691,N_3155,N_3497);
nor U3692 (N_3692,N_3450,N_3486);
or U3693 (N_3693,N_3354,N_3364);
or U3694 (N_3694,N_3004,N_3144);
nor U3695 (N_3695,N_3284,N_3300);
nand U3696 (N_3696,N_3207,N_3268);
and U3697 (N_3697,N_3055,N_3034);
or U3698 (N_3698,N_3266,N_3058);
nand U3699 (N_3699,N_3483,N_3111);
or U3700 (N_3700,N_3141,N_3122);
or U3701 (N_3701,N_3335,N_3270);
nand U3702 (N_3702,N_3445,N_3078);
nor U3703 (N_3703,N_3007,N_3188);
or U3704 (N_3704,N_3029,N_3150);
or U3705 (N_3705,N_3213,N_3116);
or U3706 (N_3706,N_3172,N_3113);
or U3707 (N_3707,N_3370,N_3319);
nand U3708 (N_3708,N_3130,N_3240);
nand U3709 (N_3709,N_3316,N_3143);
or U3710 (N_3710,N_3135,N_3238);
and U3711 (N_3711,N_3037,N_3014);
nor U3712 (N_3712,N_3061,N_3451);
or U3713 (N_3713,N_3009,N_3087);
or U3714 (N_3714,N_3311,N_3230);
or U3715 (N_3715,N_3102,N_3391);
nor U3716 (N_3716,N_3075,N_3255);
and U3717 (N_3717,N_3006,N_3026);
or U3718 (N_3718,N_3263,N_3118);
nor U3719 (N_3719,N_3059,N_3221);
nor U3720 (N_3720,N_3248,N_3433);
nand U3721 (N_3721,N_3264,N_3376);
nand U3722 (N_3722,N_3081,N_3318);
nor U3723 (N_3723,N_3212,N_3042);
and U3724 (N_3724,N_3071,N_3128);
and U3725 (N_3725,N_3424,N_3043);
and U3726 (N_3726,N_3131,N_3124);
or U3727 (N_3727,N_3253,N_3358);
nor U3728 (N_3728,N_3272,N_3101);
nor U3729 (N_3729,N_3210,N_3439);
nor U3730 (N_3730,N_3198,N_3429);
nand U3731 (N_3731,N_3152,N_3325);
nand U3732 (N_3732,N_3231,N_3351);
nor U3733 (N_3733,N_3193,N_3413);
nand U3734 (N_3734,N_3174,N_3299);
and U3735 (N_3735,N_3275,N_3260);
or U3736 (N_3736,N_3227,N_3331);
nor U3737 (N_3737,N_3011,N_3492);
or U3738 (N_3738,N_3278,N_3446);
and U3739 (N_3739,N_3186,N_3170);
nand U3740 (N_3740,N_3357,N_3002);
and U3741 (N_3741,N_3254,N_3285);
nor U3742 (N_3742,N_3384,N_3052);
nor U3743 (N_3743,N_3395,N_3496);
nand U3744 (N_3744,N_3046,N_3366);
or U3745 (N_3745,N_3417,N_3403);
nor U3746 (N_3746,N_3236,N_3098);
or U3747 (N_3747,N_3149,N_3082);
or U3748 (N_3748,N_3280,N_3389);
nor U3749 (N_3749,N_3368,N_3415);
nor U3750 (N_3750,N_3395,N_3003);
nand U3751 (N_3751,N_3031,N_3185);
and U3752 (N_3752,N_3322,N_3377);
nand U3753 (N_3753,N_3027,N_3480);
or U3754 (N_3754,N_3252,N_3424);
and U3755 (N_3755,N_3135,N_3397);
nor U3756 (N_3756,N_3347,N_3192);
nand U3757 (N_3757,N_3116,N_3091);
nand U3758 (N_3758,N_3368,N_3210);
nand U3759 (N_3759,N_3140,N_3032);
and U3760 (N_3760,N_3209,N_3240);
or U3761 (N_3761,N_3356,N_3444);
or U3762 (N_3762,N_3150,N_3366);
nor U3763 (N_3763,N_3246,N_3235);
or U3764 (N_3764,N_3409,N_3030);
nand U3765 (N_3765,N_3433,N_3151);
and U3766 (N_3766,N_3333,N_3067);
nand U3767 (N_3767,N_3422,N_3367);
and U3768 (N_3768,N_3404,N_3001);
nor U3769 (N_3769,N_3194,N_3371);
nor U3770 (N_3770,N_3037,N_3138);
nor U3771 (N_3771,N_3323,N_3495);
nor U3772 (N_3772,N_3462,N_3258);
nor U3773 (N_3773,N_3472,N_3095);
nand U3774 (N_3774,N_3375,N_3447);
and U3775 (N_3775,N_3113,N_3137);
nand U3776 (N_3776,N_3059,N_3296);
and U3777 (N_3777,N_3272,N_3244);
nand U3778 (N_3778,N_3002,N_3289);
and U3779 (N_3779,N_3027,N_3489);
nand U3780 (N_3780,N_3243,N_3131);
or U3781 (N_3781,N_3153,N_3118);
nor U3782 (N_3782,N_3448,N_3066);
nor U3783 (N_3783,N_3364,N_3400);
nand U3784 (N_3784,N_3339,N_3211);
nand U3785 (N_3785,N_3430,N_3338);
or U3786 (N_3786,N_3320,N_3225);
or U3787 (N_3787,N_3256,N_3313);
and U3788 (N_3788,N_3219,N_3265);
or U3789 (N_3789,N_3155,N_3344);
nand U3790 (N_3790,N_3455,N_3268);
nand U3791 (N_3791,N_3140,N_3483);
nor U3792 (N_3792,N_3296,N_3126);
and U3793 (N_3793,N_3431,N_3073);
or U3794 (N_3794,N_3338,N_3286);
or U3795 (N_3795,N_3235,N_3372);
nor U3796 (N_3796,N_3280,N_3008);
or U3797 (N_3797,N_3380,N_3236);
and U3798 (N_3798,N_3350,N_3265);
or U3799 (N_3799,N_3047,N_3230);
or U3800 (N_3800,N_3134,N_3050);
nor U3801 (N_3801,N_3252,N_3426);
and U3802 (N_3802,N_3081,N_3434);
xnor U3803 (N_3803,N_3007,N_3225);
and U3804 (N_3804,N_3073,N_3399);
nand U3805 (N_3805,N_3027,N_3273);
and U3806 (N_3806,N_3347,N_3054);
nand U3807 (N_3807,N_3310,N_3430);
nand U3808 (N_3808,N_3346,N_3265);
and U3809 (N_3809,N_3017,N_3219);
nor U3810 (N_3810,N_3213,N_3020);
and U3811 (N_3811,N_3098,N_3457);
nand U3812 (N_3812,N_3062,N_3309);
nor U3813 (N_3813,N_3092,N_3152);
or U3814 (N_3814,N_3131,N_3479);
or U3815 (N_3815,N_3202,N_3067);
nand U3816 (N_3816,N_3010,N_3115);
nor U3817 (N_3817,N_3188,N_3396);
nand U3818 (N_3818,N_3089,N_3097);
or U3819 (N_3819,N_3193,N_3154);
nor U3820 (N_3820,N_3262,N_3022);
nor U3821 (N_3821,N_3282,N_3378);
or U3822 (N_3822,N_3057,N_3360);
and U3823 (N_3823,N_3491,N_3382);
and U3824 (N_3824,N_3325,N_3479);
or U3825 (N_3825,N_3410,N_3168);
nand U3826 (N_3826,N_3046,N_3228);
and U3827 (N_3827,N_3018,N_3417);
or U3828 (N_3828,N_3127,N_3061);
nor U3829 (N_3829,N_3332,N_3268);
or U3830 (N_3830,N_3347,N_3285);
or U3831 (N_3831,N_3121,N_3441);
nor U3832 (N_3832,N_3053,N_3343);
nor U3833 (N_3833,N_3075,N_3183);
and U3834 (N_3834,N_3356,N_3225);
or U3835 (N_3835,N_3125,N_3048);
or U3836 (N_3836,N_3407,N_3498);
or U3837 (N_3837,N_3260,N_3407);
nor U3838 (N_3838,N_3358,N_3474);
nand U3839 (N_3839,N_3478,N_3268);
nor U3840 (N_3840,N_3351,N_3455);
and U3841 (N_3841,N_3437,N_3343);
nor U3842 (N_3842,N_3334,N_3340);
nand U3843 (N_3843,N_3061,N_3093);
nand U3844 (N_3844,N_3048,N_3325);
nand U3845 (N_3845,N_3442,N_3446);
and U3846 (N_3846,N_3175,N_3239);
nor U3847 (N_3847,N_3143,N_3400);
nand U3848 (N_3848,N_3472,N_3168);
nor U3849 (N_3849,N_3245,N_3051);
or U3850 (N_3850,N_3021,N_3118);
or U3851 (N_3851,N_3450,N_3217);
or U3852 (N_3852,N_3333,N_3153);
and U3853 (N_3853,N_3449,N_3138);
nor U3854 (N_3854,N_3262,N_3039);
nor U3855 (N_3855,N_3177,N_3368);
nor U3856 (N_3856,N_3012,N_3329);
nand U3857 (N_3857,N_3488,N_3136);
or U3858 (N_3858,N_3112,N_3271);
nand U3859 (N_3859,N_3223,N_3214);
and U3860 (N_3860,N_3147,N_3347);
nand U3861 (N_3861,N_3232,N_3071);
and U3862 (N_3862,N_3228,N_3095);
or U3863 (N_3863,N_3243,N_3409);
and U3864 (N_3864,N_3309,N_3175);
nor U3865 (N_3865,N_3472,N_3455);
or U3866 (N_3866,N_3227,N_3224);
or U3867 (N_3867,N_3244,N_3306);
or U3868 (N_3868,N_3353,N_3096);
or U3869 (N_3869,N_3459,N_3050);
nor U3870 (N_3870,N_3163,N_3243);
or U3871 (N_3871,N_3321,N_3296);
nor U3872 (N_3872,N_3432,N_3170);
nor U3873 (N_3873,N_3215,N_3119);
and U3874 (N_3874,N_3422,N_3020);
nor U3875 (N_3875,N_3354,N_3290);
nand U3876 (N_3876,N_3034,N_3091);
or U3877 (N_3877,N_3400,N_3415);
nor U3878 (N_3878,N_3265,N_3082);
and U3879 (N_3879,N_3332,N_3190);
nand U3880 (N_3880,N_3392,N_3417);
nor U3881 (N_3881,N_3472,N_3066);
or U3882 (N_3882,N_3192,N_3099);
or U3883 (N_3883,N_3325,N_3476);
nor U3884 (N_3884,N_3468,N_3274);
and U3885 (N_3885,N_3360,N_3340);
nor U3886 (N_3886,N_3219,N_3245);
nor U3887 (N_3887,N_3181,N_3306);
nor U3888 (N_3888,N_3460,N_3160);
or U3889 (N_3889,N_3402,N_3264);
nand U3890 (N_3890,N_3186,N_3309);
nor U3891 (N_3891,N_3190,N_3157);
and U3892 (N_3892,N_3363,N_3228);
and U3893 (N_3893,N_3482,N_3289);
or U3894 (N_3894,N_3327,N_3340);
or U3895 (N_3895,N_3182,N_3232);
nor U3896 (N_3896,N_3056,N_3121);
or U3897 (N_3897,N_3378,N_3425);
nand U3898 (N_3898,N_3402,N_3277);
nand U3899 (N_3899,N_3464,N_3224);
and U3900 (N_3900,N_3271,N_3423);
nor U3901 (N_3901,N_3102,N_3455);
and U3902 (N_3902,N_3454,N_3366);
or U3903 (N_3903,N_3232,N_3283);
or U3904 (N_3904,N_3449,N_3248);
nand U3905 (N_3905,N_3404,N_3490);
or U3906 (N_3906,N_3459,N_3334);
or U3907 (N_3907,N_3301,N_3145);
nand U3908 (N_3908,N_3334,N_3321);
or U3909 (N_3909,N_3182,N_3043);
and U3910 (N_3910,N_3109,N_3252);
and U3911 (N_3911,N_3400,N_3138);
nor U3912 (N_3912,N_3257,N_3361);
nor U3913 (N_3913,N_3378,N_3210);
and U3914 (N_3914,N_3124,N_3152);
or U3915 (N_3915,N_3479,N_3466);
or U3916 (N_3916,N_3356,N_3468);
nor U3917 (N_3917,N_3475,N_3270);
or U3918 (N_3918,N_3163,N_3308);
or U3919 (N_3919,N_3429,N_3499);
and U3920 (N_3920,N_3058,N_3101);
nand U3921 (N_3921,N_3139,N_3478);
nand U3922 (N_3922,N_3446,N_3315);
and U3923 (N_3923,N_3378,N_3384);
and U3924 (N_3924,N_3490,N_3287);
nand U3925 (N_3925,N_3222,N_3452);
and U3926 (N_3926,N_3361,N_3451);
or U3927 (N_3927,N_3119,N_3385);
or U3928 (N_3928,N_3248,N_3343);
or U3929 (N_3929,N_3270,N_3309);
and U3930 (N_3930,N_3403,N_3318);
or U3931 (N_3931,N_3083,N_3172);
or U3932 (N_3932,N_3149,N_3087);
nor U3933 (N_3933,N_3153,N_3460);
nand U3934 (N_3934,N_3196,N_3276);
or U3935 (N_3935,N_3364,N_3374);
nor U3936 (N_3936,N_3115,N_3059);
nor U3937 (N_3937,N_3255,N_3191);
and U3938 (N_3938,N_3164,N_3441);
and U3939 (N_3939,N_3347,N_3256);
nand U3940 (N_3940,N_3241,N_3337);
nor U3941 (N_3941,N_3454,N_3327);
and U3942 (N_3942,N_3453,N_3274);
and U3943 (N_3943,N_3041,N_3388);
nand U3944 (N_3944,N_3366,N_3096);
or U3945 (N_3945,N_3115,N_3074);
or U3946 (N_3946,N_3375,N_3040);
nand U3947 (N_3947,N_3403,N_3401);
nand U3948 (N_3948,N_3015,N_3247);
nand U3949 (N_3949,N_3247,N_3209);
nand U3950 (N_3950,N_3089,N_3359);
nor U3951 (N_3951,N_3463,N_3122);
nand U3952 (N_3952,N_3439,N_3170);
nor U3953 (N_3953,N_3497,N_3180);
and U3954 (N_3954,N_3132,N_3365);
or U3955 (N_3955,N_3337,N_3101);
or U3956 (N_3956,N_3278,N_3295);
nand U3957 (N_3957,N_3397,N_3307);
and U3958 (N_3958,N_3204,N_3199);
or U3959 (N_3959,N_3160,N_3238);
nand U3960 (N_3960,N_3221,N_3331);
nand U3961 (N_3961,N_3051,N_3103);
or U3962 (N_3962,N_3397,N_3139);
and U3963 (N_3963,N_3178,N_3254);
and U3964 (N_3964,N_3200,N_3182);
and U3965 (N_3965,N_3314,N_3186);
nor U3966 (N_3966,N_3018,N_3203);
or U3967 (N_3967,N_3442,N_3400);
nand U3968 (N_3968,N_3005,N_3044);
or U3969 (N_3969,N_3284,N_3389);
and U3970 (N_3970,N_3242,N_3398);
or U3971 (N_3971,N_3494,N_3018);
nand U3972 (N_3972,N_3349,N_3493);
nor U3973 (N_3973,N_3135,N_3060);
nand U3974 (N_3974,N_3023,N_3387);
and U3975 (N_3975,N_3083,N_3070);
and U3976 (N_3976,N_3397,N_3383);
nand U3977 (N_3977,N_3204,N_3120);
nand U3978 (N_3978,N_3485,N_3121);
nand U3979 (N_3979,N_3217,N_3482);
or U3980 (N_3980,N_3141,N_3139);
or U3981 (N_3981,N_3372,N_3101);
and U3982 (N_3982,N_3212,N_3405);
or U3983 (N_3983,N_3094,N_3474);
nor U3984 (N_3984,N_3427,N_3120);
nand U3985 (N_3985,N_3057,N_3358);
and U3986 (N_3986,N_3006,N_3124);
or U3987 (N_3987,N_3206,N_3032);
nor U3988 (N_3988,N_3157,N_3216);
nand U3989 (N_3989,N_3415,N_3153);
nor U3990 (N_3990,N_3177,N_3174);
nand U3991 (N_3991,N_3248,N_3471);
or U3992 (N_3992,N_3249,N_3035);
or U3993 (N_3993,N_3361,N_3232);
or U3994 (N_3994,N_3477,N_3384);
and U3995 (N_3995,N_3200,N_3430);
nor U3996 (N_3996,N_3492,N_3067);
and U3997 (N_3997,N_3150,N_3495);
and U3998 (N_3998,N_3274,N_3061);
nor U3999 (N_3999,N_3211,N_3340);
nand U4000 (N_4000,N_3863,N_3645);
nand U4001 (N_4001,N_3699,N_3789);
nor U4002 (N_4002,N_3716,N_3772);
nor U4003 (N_4003,N_3788,N_3638);
nand U4004 (N_4004,N_3726,N_3949);
and U4005 (N_4005,N_3641,N_3874);
and U4006 (N_4006,N_3795,N_3833);
nand U4007 (N_4007,N_3852,N_3545);
nand U4008 (N_4008,N_3862,N_3991);
and U4009 (N_4009,N_3929,N_3786);
nor U4010 (N_4010,N_3683,N_3878);
or U4011 (N_4011,N_3958,N_3625);
or U4012 (N_4012,N_3662,N_3721);
or U4013 (N_4013,N_3696,N_3647);
or U4014 (N_4014,N_3681,N_3692);
nor U4015 (N_4015,N_3679,N_3698);
nor U4016 (N_4016,N_3654,N_3834);
or U4017 (N_4017,N_3604,N_3741);
nand U4018 (N_4018,N_3501,N_3932);
or U4019 (N_4019,N_3558,N_3888);
or U4020 (N_4020,N_3573,N_3898);
nand U4021 (N_4021,N_3818,N_3694);
and U4022 (N_4022,N_3970,N_3646);
and U4023 (N_4023,N_3785,N_3589);
nand U4024 (N_4024,N_3961,N_3986);
nor U4025 (N_4025,N_3596,N_3639);
nand U4026 (N_4026,N_3658,N_3881);
and U4027 (N_4027,N_3511,N_3619);
or U4028 (N_4028,N_3842,N_3736);
or U4029 (N_4029,N_3931,N_3676);
and U4030 (N_4030,N_3876,N_3928);
and U4031 (N_4031,N_3959,N_3934);
nand U4032 (N_4032,N_3925,N_3762);
and U4033 (N_4033,N_3602,N_3983);
nand U4034 (N_4034,N_3856,N_3951);
nor U4035 (N_4035,N_3728,N_3743);
nand U4036 (N_4036,N_3980,N_3627);
nand U4037 (N_4037,N_3629,N_3872);
nor U4038 (N_4038,N_3583,N_3776);
nand U4039 (N_4039,N_3615,N_3671);
or U4040 (N_4040,N_3582,N_3996);
and U4041 (N_4041,N_3708,N_3797);
or U4042 (N_4042,N_3841,N_3550);
nand U4043 (N_4043,N_3590,N_3712);
nor U4044 (N_4044,N_3591,N_3967);
nand U4045 (N_4045,N_3952,N_3960);
nand U4046 (N_4046,N_3910,N_3992);
nor U4047 (N_4047,N_3865,N_3626);
or U4048 (N_4048,N_3606,N_3846);
or U4049 (N_4049,N_3636,N_3853);
and U4050 (N_4050,N_3567,N_3701);
nand U4051 (N_4051,N_3551,N_3571);
nand U4052 (N_4052,N_3611,N_3840);
nor U4053 (N_4053,N_3924,N_3977);
nand U4054 (N_4054,N_3587,N_3782);
and U4055 (N_4055,N_3908,N_3754);
and U4056 (N_4056,N_3635,N_3526);
xnor U4057 (N_4057,N_3897,N_3819);
nand U4058 (N_4058,N_3826,N_3978);
and U4059 (N_4059,N_3889,N_3631);
or U4060 (N_4060,N_3505,N_3588);
nand U4061 (N_4061,N_3825,N_3945);
nand U4062 (N_4062,N_3560,N_3612);
nand U4063 (N_4063,N_3578,N_3901);
and U4064 (N_4064,N_3987,N_3643);
or U4065 (N_4065,N_3745,N_3665);
and U4066 (N_4066,N_3860,N_3637);
nand U4067 (N_4067,N_3542,N_3974);
and U4068 (N_4068,N_3870,N_3737);
or U4069 (N_4069,N_3927,N_3500);
nor U4070 (N_4070,N_3514,N_3890);
nand U4071 (N_4071,N_3779,N_3892);
nand U4072 (N_4072,N_3668,N_3807);
nand U4073 (N_4073,N_3933,N_3957);
and U4074 (N_4074,N_3656,N_3963);
nor U4075 (N_4075,N_3584,N_3792);
or U4076 (N_4076,N_3747,N_3954);
nor U4077 (N_4077,N_3534,N_3948);
and U4078 (N_4078,N_3719,N_3537);
nor U4079 (N_4079,N_3577,N_3766);
or U4080 (N_4080,N_3985,N_3733);
and U4081 (N_4081,N_3599,N_3815);
and U4082 (N_4082,N_3975,N_3669);
or U4083 (N_4083,N_3735,N_3902);
and U4084 (N_4084,N_3520,N_3845);
nand U4085 (N_4085,N_3761,N_3835);
nand U4086 (N_4086,N_3667,N_3969);
nor U4087 (N_4087,N_3940,N_3912);
nand U4088 (N_4088,N_3794,N_3999);
and U4089 (N_4089,N_3718,N_3953);
or U4090 (N_4090,N_3546,N_3919);
nand U4091 (N_4091,N_3621,N_3697);
nand U4092 (N_4092,N_3793,N_3880);
or U4093 (N_4093,N_3995,N_3572);
or U4094 (N_4094,N_3784,N_3555);
nand U4095 (N_4095,N_3877,N_3704);
nor U4096 (N_4096,N_3956,N_3642);
or U4097 (N_4097,N_3528,N_3564);
or U4098 (N_4098,N_3670,N_3661);
nor U4099 (N_4099,N_3757,N_3682);
nand U4100 (N_4100,N_3773,N_3968);
or U4101 (N_4101,N_3805,N_3905);
or U4102 (N_4102,N_3962,N_3946);
or U4103 (N_4103,N_3966,N_3802);
nor U4104 (N_4104,N_3937,N_3755);
and U4105 (N_4105,N_3724,N_3965);
nand U4106 (N_4106,N_3552,N_3891);
nand U4107 (N_4107,N_3557,N_3509);
or U4108 (N_4108,N_3610,N_3715);
nor U4109 (N_4109,N_3767,N_3817);
or U4110 (N_4110,N_3541,N_3864);
nand U4111 (N_4111,N_3738,N_3909);
and U4112 (N_4112,N_3828,N_3801);
nand U4113 (N_4113,N_3886,N_3579);
nand U4114 (N_4114,N_3812,N_3559);
or U4115 (N_4115,N_3700,N_3765);
xnor U4116 (N_4116,N_3866,N_3950);
nor U4117 (N_4117,N_3790,N_3838);
nand U4118 (N_4118,N_3673,N_3502);
nor U4119 (N_4119,N_3508,N_3750);
or U4120 (N_4120,N_3632,N_3556);
and U4121 (N_4121,N_3561,N_3764);
and U4122 (N_4122,N_3533,N_3608);
nand U4123 (N_4123,N_3717,N_3981);
or U4124 (N_4124,N_3839,N_3749);
nor U4125 (N_4125,N_3798,N_3522);
nand U4126 (N_4126,N_3706,N_3650);
nand U4127 (N_4127,N_3814,N_3796);
or U4128 (N_4128,N_3525,N_3729);
nand U4129 (N_4129,N_3744,N_3623);
nand U4130 (N_4130,N_3693,N_3770);
nor U4131 (N_4131,N_3823,N_3622);
or U4132 (N_4132,N_3585,N_3594);
and U4133 (N_4133,N_3707,N_3593);
and U4134 (N_4134,N_3914,N_3563);
nand U4135 (N_4135,N_3988,N_3820);
and U4136 (N_4136,N_3844,N_3882);
or U4137 (N_4137,N_3690,N_3907);
nand U4138 (N_4138,N_3935,N_3849);
or U4139 (N_4139,N_3680,N_3565);
and U4140 (N_4140,N_3603,N_3574);
nand U4141 (N_4141,N_3851,N_3936);
and U4142 (N_4142,N_3710,N_3506);
nand U4143 (N_4143,N_3711,N_3854);
and U4144 (N_4144,N_3722,N_3648);
nor U4145 (N_4145,N_3628,N_3781);
or U4146 (N_4146,N_3768,N_3869);
nor U4147 (N_4147,N_3678,N_3887);
or U4148 (N_4148,N_3831,N_3758);
nand U4149 (N_4149,N_3672,N_3518);
nand U4150 (N_4150,N_3899,N_3994);
nand U4151 (N_4151,N_3517,N_3944);
nor U4152 (N_4152,N_3879,N_3512);
nand U4153 (N_4153,N_3677,N_3685);
and U4154 (N_4154,N_3895,N_3600);
nand U4155 (N_4155,N_3822,N_3867);
or U4156 (N_4156,N_3529,N_3884);
nor U4157 (N_4157,N_3868,N_3725);
or U4158 (N_4158,N_3896,N_3739);
and U4159 (N_4159,N_3943,N_3618);
nor U4160 (N_4160,N_3675,N_3893);
or U4161 (N_4161,N_3799,N_3535);
nand U4162 (N_4162,N_3503,N_3539);
nor U4163 (N_4163,N_3947,N_3740);
and U4164 (N_4164,N_3855,N_3971);
or U4165 (N_4165,N_3544,N_3836);
nor U4166 (N_4166,N_3955,N_3832);
nor U4167 (N_4167,N_3979,N_3777);
and U4168 (N_4168,N_3997,N_3581);
nand U4169 (N_4169,N_3808,N_3727);
nand U4170 (N_4170,N_3664,N_3605);
or U4171 (N_4171,N_3911,N_3806);
nor U4172 (N_4172,N_3549,N_3554);
and U4173 (N_4173,N_3920,N_3527);
and U4174 (N_4174,N_3989,N_3649);
and U4175 (N_4175,N_3538,N_3595);
and U4176 (N_4176,N_3663,N_3837);
and U4177 (N_4177,N_3810,N_3686);
and U4178 (N_4178,N_3515,N_3939);
or U4179 (N_4179,N_3926,N_3900);
nand U4180 (N_4180,N_3660,N_3616);
and U4181 (N_4181,N_3922,N_3830);
and U4182 (N_4182,N_3703,N_3580);
and U4183 (N_4183,N_3548,N_3875);
nand U4184 (N_4184,N_3921,N_3657);
nor U4185 (N_4185,N_3859,N_3873);
nand U4186 (N_4186,N_3732,N_3783);
or U4187 (N_4187,N_3684,N_3614);
and U4188 (N_4188,N_3871,N_3941);
nor U4189 (N_4189,N_3586,N_3553);
xor U4190 (N_4190,N_3655,N_3547);
nor U4191 (N_4191,N_3811,N_3714);
or U4192 (N_4192,N_3674,N_3913);
or U4193 (N_4193,N_3780,N_3569);
or U4194 (N_4194,N_3705,N_3894);
or U4195 (N_4195,N_3816,N_3752);
and U4196 (N_4196,N_3575,N_3513);
and U4197 (N_4197,N_3976,N_3702);
and U4198 (N_4198,N_3742,N_3769);
nor U4199 (N_4199,N_3510,N_3659);
nand U4200 (N_4200,N_3691,N_3519);
or U4201 (N_4201,N_3803,N_3938);
nor U4202 (N_4202,N_3843,N_3653);
and U4203 (N_4203,N_3568,N_3923);
or U4204 (N_4204,N_3883,N_3906);
nand U4205 (N_4205,N_3601,N_3751);
nor U4206 (N_4206,N_3917,N_3562);
and U4207 (N_4207,N_3760,N_3756);
or U4208 (N_4208,N_3688,N_3827);
nand U4209 (N_4209,N_3570,N_3734);
nor U4210 (N_4210,N_3720,N_3847);
or U4211 (N_4211,N_3613,N_3532);
and U4212 (N_4212,N_3516,N_3543);
and U4213 (N_4213,N_3930,N_3530);
or U4214 (N_4214,N_3885,N_3504);
and U4215 (N_4215,N_3652,N_3630);
xnor U4216 (N_4216,N_3998,N_3759);
or U4217 (N_4217,N_3774,N_3771);
and U4218 (N_4218,N_3848,N_3644);
or U4219 (N_4219,N_3521,N_3531);
and U4220 (N_4220,N_3857,N_3540);
nor U4221 (N_4221,N_3993,N_3990);
nor U4222 (N_4222,N_3607,N_3982);
nor U4223 (N_4223,N_3634,N_3566);
and U4224 (N_4224,N_3746,N_3904);
nand U4225 (N_4225,N_3813,N_3984);
or U4226 (N_4226,N_3972,N_3791);
nor U4227 (N_4227,N_3809,N_3731);
and U4228 (N_4228,N_3964,N_3903);
nand U4229 (N_4229,N_3689,N_3651);
nor U4230 (N_4230,N_3730,N_3824);
and U4231 (N_4231,N_3536,N_3597);
xnor U4232 (N_4232,N_3800,N_3861);
and U4233 (N_4233,N_3804,N_3723);
and U4234 (N_4234,N_3748,N_3576);
nand U4235 (N_4235,N_3915,N_3787);
nor U4236 (N_4236,N_3617,N_3507);
nand U4237 (N_4237,N_3592,N_3609);
and U4238 (N_4238,N_3858,N_3753);
and U4239 (N_4239,N_3942,N_3775);
nand U4240 (N_4240,N_3687,N_3973);
nor U4241 (N_4241,N_3598,N_3695);
and U4242 (N_4242,N_3829,N_3778);
nand U4243 (N_4243,N_3666,N_3850);
or U4244 (N_4244,N_3709,N_3763);
nor U4245 (N_4245,N_3918,N_3524);
or U4246 (N_4246,N_3523,N_3821);
or U4247 (N_4247,N_3640,N_3624);
or U4248 (N_4248,N_3633,N_3713);
or U4249 (N_4249,N_3916,N_3620);
or U4250 (N_4250,N_3930,N_3708);
nand U4251 (N_4251,N_3597,N_3607);
or U4252 (N_4252,N_3595,N_3953);
nor U4253 (N_4253,N_3765,N_3856);
or U4254 (N_4254,N_3592,N_3741);
nor U4255 (N_4255,N_3783,N_3622);
nor U4256 (N_4256,N_3699,N_3996);
nor U4257 (N_4257,N_3818,N_3681);
nand U4258 (N_4258,N_3751,N_3692);
nor U4259 (N_4259,N_3667,N_3795);
or U4260 (N_4260,N_3686,N_3526);
nor U4261 (N_4261,N_3625,N_3801);
nand U4262 (N_4262,N_3880,N_3843);
nand U4263 (N_4263,N_3903,N_3738);
or U4264 (N_4264,N_3793,N_3835);
or U4265 (N_4265,N_3508,N_3728);
nor U4266 (N_4266,N_3816,N_3554);
or U4267 (N_4267,N_3558,N_3894);
nand U4268 (N_4268,N_3753,N_3850);
nand U4269 (N_4269,N_3840,N_3524);
or U4270 (N_4270,N_3990,N_3516);
or U4271 (N_4271,N_3630,N_3786);
and U4272 (N_4272,N_3738,N_3601);
nand U4273 (N_4273,N_3910,N_3836);
nor U4274 (N_4274,N_3807,N_3780);
or U4275 (N_4275,N_3974,N_3955);
nand U4276 (N_4276,N_3645,N_3840);
or U4277 (N_4277,N_3544,N_3918);
and U4278 (N_4278,N_3959,N_3876);
nor U4279 (N_4279,N_3903,N_3850);
nand U4280 (N_4280,N_3969,N_3662);
or U4281 (N_4281,N_3909,N_3529);
nor U4282 (N_4282,N_3916,N_3685);
nand U4283 (N_4283,N_3996,N_3564);
nor U4284 (N_4284,N_3922,N_3508);
or U4285 (N_4285,N_3741,N_3936);
and U4286 (N_4286,N_3587,N_3603);
and U4287 (N_4287,N_3540,N_3536);
nand U4288 (N_4288,N_3941,N_3528);
or U4289 (N_4289,N_3881,N_3524);
nor U4290 (N_4290,N_3631,N_3719);
nand U4291 (N_4291,N_3820,N_3511);
or U4292 (N_4292,N_3909,N_3986);
and U4293 (N_4293,N_3770,N_3667);
nor U4294 (N_4294,N_3793,N_3952);
or U4295 (N_4295,N_3549,N_3961);
and U4296 (N_4296,N_3780,N_3607);
nor U4297 (N_4297,N_3709,N_3940);
and U4298 (N_4298,N_3733,N_3641);
nor U4299 (N_4299,N_3918,N_3936);
nand U4300 (N_4300,N_3553,N_3776);
or U4301 (N_4301,N_3703,N_3915);
and U4302 (N_4302,N_3996,N_3617);
xor U4303 (N_4303,N_3522,N_3708);
nor U4304 (N_4304,N_3571,N_3930);
nand U4305 (N_4305,N_3684,N_3575);
or U4306 (N_4306,N_3945,N_3539);
nor U4307 (N_4307,N_3973,N_3987);
nand U4308 (N_4308,N_3985,N_3932);
nor U4309 (N_4309,N_3526,N_3856);
nand U4310 (N_4310,N_3665,N_3681);
nor U4311 (N_4311,N_3897,N_3787);
nand U4312 (N_4312,N_3722,N_3945);
nand U4313 (N_4313,N_3822,N_3804);
and U4314 (N_4314,N_3600,N_3786);
or U4315 (N_4315,N_3690,N_3612);
nor U4316 (N_4316,N_3950,N_3843);
or U4317 (N_4317,N_3996,N_3920);
or U4318 (N_4318,N_3510,N_3937);
or U4319 (N_4319,N_3599,N_3933);
or U4320 (N_4320,N_3628,N_3506);
and U4321 (N_4321,N_3816,N_3642);
or U4322 (N_4322,N_3716,N_3755);
or U4323 (N_4323,N_3952,N_3867);
nand U4324 (N_4324,N_3683,N_3917);
nand U4325 (N_4325,N_3893,N_3533);
nor U4326 (N_4326,N_3595,N_3945);
or U4327 (N_4327,N_3865,N_3819);
and U4328 (N_4328,N_3529,N_3946);
and U4329 (N_4329,N_3998,N_3904);
nand U4330 (N_4330,N_3768,N_3791);
and U4331 (N_4331,N_3690,N_3617);
nor U4332 (N_4332,N_3625,N_3795);
and U4333 (N_4333,N_3539,N_3831);
or U4334 (N_4334,N_3879,N_3579);
or U4335 (N_4335,N_3876,N_3735);
and U4336 (N_4336,N_3750,N_3560);
and U4337 (N_4337,N_3506,N_3502);
xnor U4338 (N_4338,N_3744,N_3986);
nor U4339 (N_4339,N_3766,N_3956);
nor U4340 (N_4340,N_3593,N_3889);
or U4341 (N_4341,N_3770,N_3885);
nand U4342 (N_4342,N_3717,N_3528);
and U4343 (N_4343,N_3885,N_3641);
nand U4344 (N_4344,N_3877,N_3565);
nor U4345 (N_4345,N_3571,N_3904);
nor U4346 (N_4346,N_3754,N_3618);
nand U4347 (N_4347,N_3983,N_3780);
nand U4348 (N_4348,N_3755,N_3512);
nand U4349 (N_4349,N_3600,N_3923);
and U4350 (N_4350,N_3987,N_3869);
nand U4351 (N_4351,N_3685,N_3520);
xor U4352 (N_4352,N_3815,N_3675);
and U4353 (N_4353,N_3854,N_3776);
and U4354 (N_4354,N_3550,N_3825);
nand U4355 (N_4355,N_3894,N_3648);
nor U4356 (N_4356,N_3948,N_3905);
and U4357 (N_4357,N_3752,N_3961);
nand U4358 (N_4358,N_3993,N_3792);
and U4359 (N_4359,N_3531,N_3760);
or U4360 (N_4360,N_3583,N_3690);
or U4361 (N_4361,N_3821,N_3696);
or U4362 (N_4362,N_3638,N_3504);
nand U4363 (N_4363,N_3612,N_3762);
or U4364 (N_4364,N_3508,N_3762);
or U4365 (N_4365,N_3599,N_3822);
and U4366 (N_4366,N_3856,N_3515);
or U4367 (N_4367,N_3623,N_3906);
nand U4368 (N_4368,N_3723,N_3926);
nor U4369 (N_4369,N_3811,N_3799);
nor U4370 (N_4370,N_3833,N_3733);
nand U4371 (N_4371,N_3593,N_3695);
or U4372 (N_4372,N_3767,N_3838);
nor U4373 (N_4373,N_3540,N_3571);
nand U4374 (N_4374,N_3852,N_3858);
and U4375 (N_4375,N_3537,N_3751);
nor U4376 (N_4376,N_3697,N_3908);
nor U4377 (N_4377,N_3874,N_3553);
and U4378 (N_4378,N_3620,N_3597);
nand U4379 (N_4379,N_3567,N_3537);
nand U4380 (N_4380,N_3769,N_3654);
nor U4381 (N_4381,N_3919,N_3699);
nor U4382 (N_4382,N_3981,N_3651);
nor U4383 (N_4383,N_3784,N_3615);
nand U4384 (N_4384,N_3653,N_3508);
nor U4385 (N_4385,N_3962,N_3905);
nor U4386 (N_4386,N_3802,N_3637);
and U4387 (N_4387,N_3643,N_3877);
nor U4388 (N_4388,N_3859,N_3882);
or U4389 (N_4389,N_3651,N_3708);
or U4390 (N_4390,N_3900,N_3589);
nand U4391 (N_4391,N_3831,N_3597);
nand U4392 (N_4392,N_3971,N_3821);
or U4393 (N_4393,N_3509,N_3647);
nor U4394 (N_4394,N_3505,N_3755);
and U4395 (N_4395,N_3545,N_3862);
or U4396 (N_4396,N_3695,N_3508);
or U4397 (N_4397,N_3864,N_3860);
or U4398 (N_4398,N_3993,N_3795);
and U4399 (N_4399,N_3911,N_3656);
nor U4400 (N_4400,N_3852,N_3622);
nand U4401 (N_4401,N_3620,N_3660);
nand U4402 (N_4402,N_3997,N_3605);
or U4403 (N_4403,N_3592,N_3562);
or U4404 (N_4404,N_3517,N_3722);
nor U4405 (N_4405,N_3516,N_3585);
and U4406 (N_4406,N_3547,N_3666);
nor U4407 (N_4407,N_3560,N_3980);
nor U4408 (N_4408,N_3987,N_3959);
nor U4409 (N_4409,N_3621,N_3848);
nor U4410 (N_4410,N_3506,N_3771);
or U4411 (N_4411,N_3817,N_3900);
and U4412 (N_4412,N_3750,N_3777);
or U4413 (N_4413,N_3878,N_3571);
nor U4414 (N_4414,N_3972,N_3536);
and U4415 (N_4415,N_3753,N_3825);
nand U4416 (N_4416,N_3578,N_3761);
nand U4417 (N_4417,N_3559,N_3866);
nor U4418 (N_4418,N_3581,N_3506);
nand U4419 (N_4419,N_3528,N_3577);
nand U4420 (N_4420,N_3916,N_3608);
nand U4421 (N_4421,N_3643,N_3576);
nand U4422 (N_4422,N_3858,N_3888);
or U4423 (N_4423,N_3884,N_3767);
nand U4424 (N_4424,N_3691,N_3614);
nor U4425 (N_4425,N_3535,N_3991);
nor U4426 (N_4426,N_3763,N_3710);
and U4427 (N_4427,N_3786,N_3800);
nand U4428 (N_4428,N_3676,N_3608);
and U4429 (N_4429,N_3762,N_3837);
nand U4430 (N_4430,N_3559,N_3892);
or U4431 (N_4431,N_3953,N_3652);
nor U4432 (N_4432,N_3671,N_3736);
and U4433 (N_4433,N_3703,N_3581);
and U4434 (N_4434,N_3981,N_3663);
or U4435 (N_4435,N_3595,N_3964);
or U4436 (N_4436,N_3670,N_3781);
nand U4437 (N_4437,N_3894,N_3937);
nand U4438 (N_4438,N_3695,N_3817);
nor U4439 (N_4439,N_3903,N_3896);
or U4440 (N_4440,N_3956,N_3844);
nor U4441 (N_4441,N_3877,N_3872);
nor U4442 (N_4442,N_3823,N_3715);
and U4443 (N_4443,N_3971,N_3765);
or U4444 (N_4444,N_3945,N_3789);
nor U4445 (N_4445,N_3644,N_3841);
nor U4446 (N_4446,N_3814,N_3778);
or U4447 (N_4447,N_3641,N_3558);
and U4448 (N_4448,N_3974,N_3945);
nor U4449 (N_4449,N_3951,N_3899);
or U4450 (N_4450,N_3529,N_3587);
and U4451 (N_4451,N_3866,N_3670);
nor U4452 (N_4452,N_3520,N_3765);
nor U4453 (N_4453,N_3981,N_3858);
nor U4454 (N_4454,N_3586,N_3517);
and U4455 (N_4455,N_3762,N_3666);
nand U4456 (N_4456,N_3582,N_3838);
and U4457 (N_4457,N_3534,N_3698);
or U4458 (N_4458,N_3674,N_3805);
nand U4459 (N_4459,N_3679,N_3875);
and U4460 (N_4460,N_3699,N_3816);
and U4461 (N_4461,N_3963,N_3819);
nand U4462 (N_4462,N_3837,N_3773);
and U4463 (N_4463,N_3840,N_3624);
and U4464 (N_4464,N_3548,N_3800);
and U4465 (N_4465,N_3670,N_3934);
or U4466 (N_4466,N_3708,N_3965);
nand U4467 (N_4467,N_3502,N_3973);
nor U4468 (N_4468,N_3743,N_3636);
nand U4469 (N_4469,N_3867,N_3660);
and U4470 (N_4470,N_3787,N_3731);
and U4471 (N_4471,N_3714,N_3650);
xor U4472 (N_4472,N_3613,N_3654);
nand U4473 (N_4473,N_3932,N_3945);
and U4474 (N_4474,N_3790,N_3921);
or U4475 (N_4475,N_3540,N_3650);
and U4476 (N_4476,N_3750,N_3711);
nor U4477 (N_4477,N_3541,N_3975);
nand U4478 (N_4478,N_3707,N_3588);
nand U4479 (N_4479,N_3724,N_3575);
xor U4480 (N_4480,N_3605,N_3809);
nand U4481 (N_4481,N_3665,N_3530);
and U4482 (N_4482,N_3504,N_3511);
and U4483 (N_4483,N_3898,N_3788);
nor U4484 (N_4484,N_3663,N_3561);
nor U4485 (N_4485,N_3773,N_3766);
or U4486 (N_4486,N_3968,N_3948);
and U4487 (N_4487,N_3919,N_3743);
nor U4488 (N_4488,N_3735,N_3835);
nor U4489 (N_4489,N_3653,N_3826);
nand U4490 (N_4490,N_3688,N_3595);
and U4491 (N_4491,N_3587,N_3996);
nor U4492 (N_4492,N_3947,N_3651);
or U4493 (N_4493,N_3837,N_3590);
and U4494 (N_4494,N_3590,N_3655);
or U4495 (N_4495,N_3641,N_3710);
nor U4496 (N_4496,N_3759,N_3563);
and U4497 (N_4497,N_3591,N_3722);
nor U4498 (N_4498,N_3751,N_3796);
nand U4499 (N_4499,N_3667,N_3772);
and U4500 (N_4500,N_4319,N_4383);
nor U4501 (N_4501,N_4478,N_4302);
nor U4502 (N_4502,N_4473,N_4039);
nand U4503 (N_4503,N_4176,N_4119);
or U4504 (N_4504,N_4173,N_4469);
nor U4505 (N_4505,N_4028,N_4390);
nand U4506 (N_4506,N_4282,N_4378);
nand U4507 (N_4507,N_4144,N_4297);
or U4508 (N_4508,N_4356,N_4274);
and U4509 (N_4509,N_4163,N_4171);
nor U4510 (N_4510,N_4277,N_4232);
nand U4511 (N_4511,N_4299,N_4472);
nor U4512 (N_4512,N_4262,N_4010);
and U4513 (N_4513,N_4270,N_4480);
nor U4514 (N_4514,N_4229,N_4191);
and U4515 (N_4515,N_4419,N_4209);
nor U4516 (N_4516,N_4219,N_4036);
or U4517 (N_4517,N_4303,N_4442);
and U4518 (N_4518,N_4353,N_4427);
nand U4519 (N_4519,N_4037,N_4438);
nand U4520 (N_4520,N_4100,N_4338);
and U4521 (N_4521,N_4159,N_4058);
nor U4522 (N_4522,N_4385,N_4214);
nor U4523 (N_4523,N_4175,N_4285);
or U4524 (N_4524,N_4174,N_4321);
or U4525 (N_4525,N_4309,N_4283);
nand U4526 (N_4526,N_4448,N_4399);
and U4527 (N_4527,N_4167,N_4308);
or U4528 (N_4528,N_4123,N_4458);
nand U4529 (N_4529,N_4375,N_4252);
or U4530 (N_4530,N_4397,N_4327);
and U4531 (N_4531,N_4437,N_4064);
or U4532 (N_4532,N_4475,N_4195);
nor U4533 (N_4533,N_4244,N_4294);
or U4534 (N_4534,N_4067,N_4073);
and U4535 (N_4535,N_4426,N_4150);
nand U4536 (N_4536,N_4396,N_4454);
nand U4537 (N_4537,N_4237,N_4117);
or U4538 (N_4538,N_4009,N_4449);
or U4539 (N_4539,N_4253,N_4323);
nand U4540 (N_4540,N_4223,N_4366);
nand U4541 (N_4541,N_4372,N_4129);
nor U4542 (N_4542,N_4069,N_4351);
nor U4543 (N_4543,N_4025,N_4127);
nor U4544 (N_4544,N_4125,N_4359);
and U4545 (N_4545,N_4062,N_4160);
nand U4546 (N_4546,N_4398,N_4026);
nand U4547 (N_4547,N_4441,N_4381);
nand U4548 (N_4548,N_4003,N_4030);
and U4549 (N_4549,N_4393,N_4379);
nor U4550 (N_4550,N_4417,N_4189);
or U4551 (N_4551,N_4004,N_4373);
nor U4552 (N_4552,N_4406,N_4422);
and U4553 (N_4553,N_4466,N_4235);
or U4554 (N_4554,N_4497,N_4126);
and U4555 (N_4555,N_4492,N_4247);
or U4556 (N_4556,N_4094,N_4170);
and U4557 (N_4557,N_4272,N_4263);
nand U4558 (N_4558,N_4459,N_4217);
and U4559 (N_4559,N_4413,N_4177);
and U4560 (N_4560,N_4462,N_4114);
nand U4561 (N_4561,N_4330,N_4290);
and U4562 (N_4562,N_4334,N_4249);
nand U4563 (N_4563,N_4401,N_4298);
and U4564 (N_4564,N_4429,N_4121);
nand U4565 (N_4565,N_4395,N_4460);
nor U4566 (N_4566,N_4193,N_4051);
nor U4567 (N_4567,N_4246,N_4345);
nor U4568 (N_4568,N_4444,N_4452);
or U4569 (N_4569,N_4013,N_4499);
nor U4570 (N_4570,N_4254,N_4428);
nand U4571 (N_4571,N_4485,N_4260);
and U4572 (N_4572,N_4352,N_4233);
and U4573 (N_4573,N_4464,N_4491);
nor U4574 (N_4574,N_4280,N_4151);
nor U4575 (N_4575,N_4342,N_4139);
nor U4576 (N_4576,N_4349,N_4197);
nand U4577 (N_4577,N_4425,N_4494);
nand U4578 (N_4578,N_4227,N_4423);
or U4579 (N_4579,N_4453,N_4243);
and U4580 (N_4580,N_4387,N_4434);
nor U4581 (N_4581,N_4134,N_4063);
and U4582 (N_4582,N_4465,N_4137);
or U4583 (N_4583,N_4082,N_4386);
nand U4584 (N_4584,N_4412,N_4200);
or U4585 (N_4585,N_4113,N_4258);
and U4586 (N_4586,N_4220,N_4410);
nand U4587 (N_4587,N_4456,N_4078);
nor U4588 (N_4588,N_4455,N_4043);
and U4589 (N_4589,N_4482,N_4157);
nand U4590 (N_4590,N_4055,N_4088);
or U4591 (N_4591,N_4124,N_4207);
nand U4592 (N_4592,N_4420,N_4259);
nand U4593 (N_4593,N_4289,N_4221);
and U4594 (N_4594,N_4486,N_4084);
nand U4595 (N_4595,N_4218,N_4181);
nand U4596 (N_4596,N_4414,N_4291);
nor U4597 (N_4597,N_4196,N_4186);
and U4598 (N_4598,N_4314,N_4089);
nor U4599 (N_4599,N_4045,N_4066);
and U4600 (N_4600,N_4182,N_4484);
nand U4601 (N_4601,N_4098,N_4076);
or U4602 (N_4602,N_4116,N_4046);
nor U4603 (N_4603,N_4267,N_4156);
nor U4604 (N_4604,N_4436,N_4421);
and U4605 (N_4605,N_4047,N_4060);
and U4606 (N_4606,N_4012,N_4257);
and U4607 (N_4607,N_4268,N_4476);
nor U4608 (N_4608,N_4337,N_4205);
or U4609 (N_4609,N_4305,N_4131);
or U4610 (N_4610,N_4279,N_4145);
and U4611 (N_4611,N_4198,N_4471);
and U4612 (N_4612,N_4130,N_4498);
nand U4613 (N_4613,N_4435,N_4049);
nor U4614 (N_4614,N_4147,N_4087);
nand U4615 (N_4615,N_4408,N_4018);
nor U4616 (N_4616,N_4143,N_4095);
nor U4617 (N_4617,N_4059,N_4006);
and U4618 (N_4618,N_4324,N_4029);
or U4619 (N_4619,N_4447,N_4365);
nand U4620 (N_4620,N_4377,N_4360);
or U4621 (N_4621,N_4122,N_4287);
nand U4622 (N_4622,N_4140,N_4072);
and U4623 (N_4623,N_4384,N_4281);
and U4624 (N_4624,N_4407,N_4310);
nor U4625 (N_4625,N_4344,N_4483);
or U4626 (N_4626,N_4264,N_4265);
nand U4627 (N_4627,N_4015,N_4431);
and U4628 (N_4628,N_4216,N_4370);
or U4629 (N_4629,N_4135,N_4346);
nand U4630 (N_4630,N_4011,N_4208);
and U4631 (N_4631,N_4261,N_4248);
nor U4632 (N_4632,N_4206,N_4023);
nor U4633 (N_4633,N_4090,N_4236);
and U4634 (N_4634,N_4403,N_4457);
and U4635 (N_4635,N_4065,N_4038);
nor U4636 (N_4636,N_4154,N_4101);
nand U4637 (N_4637,N_4112,N_4179);
nand U4638 (N_4638,N_4409,N_4042);
nor U4639 (N_4639,N_4284,N_4192);
nor U4640 (N_4640,N_4041,N_4091);
and U4641 (N_4641,N_4416,N_4008);
and U4642 (N_4642,N_4450,N_4120);
nor U4643 (N_4643,N_4363,N_4085);
nor U4644 (N_4644,N_4424,N_4071);
or U4645 (N_4645,N_4228,N_4418);
nand U4646 (N_4646,N_4230,N_4096);
nand U4647 (N_4647,N_4354,N_4312);
or U4648 (N_4648,N_4276,N_4273);
nor U4649 (N_4649,N_4343,N_4389);
or U4650 (N_4650,N_4070,N_4374);
nand U4651 (N_4651,N_4231,N_4307);
nor U4652 (N_4652,N_4148,N_4295);
nor U4653 (N_4653,N_4439,N_4316);
nor U4654 (N_4654,N_4180,N_4487);
and U4655 (N_4655,N_4380,N_4024);
nor U4656 (N_4656,N_4361,N_4052);
and U4657 (N_4657,N_4190,N_4315);
nand U4658 (N_4658,N_4007,N_4187);
or U4659 (N_4659,N_4204,N_4057);
nor U4660 (N_4660,N_4490,N_4102);
nor U4661 (N_4661,N_4250,N_4288);
nand U4662 (N_4662,N_4463,N_4111);
nor U4663 (N_4663,N_4222,N_4357);
or U4664 (N_4664,N_4239,N_4162);
nor U4665 (N_4665,N_4251,N_4077);
nor U4666 (N_4666,N_4341,N_4443);
and U4667 (N_4667,N_4301,N_4211);
nor U4668 (N_4668,N_4155,N_4014);
nor U4669 (N_4669,N_4245,N_4234);
or U4670 (N_4670,N_4040,N_4000);
or U4671 (N_4671,N_4031,N_4056);
or U4672 (N_4672,N_4099,N_4355);
and U4673 (N_4673,N_4371,N_4138);
and U4674 (N_4674,N_4415,N_4496);
nor U4675 (N_4675,N_4210,N_4165);
and U4676 (N_4676,N_4002,N_4027);
and U4677 (N_4677,N_4325,N_4440);
and U4678 (N_4678,N_4061,N_4376);
and U4679 (N_4679,N_4255,N_4118);
and U4680 (N_4680,N_4278,N_4106);
or U4681 (N_4681,N_4035,N_4226);
and U4682 (N_4682,N_4184,N_4053);
or U4683 (N_4683,N_4021,N_4347);
or U4684 (N_4684,N_4275,N_4430);
nor U4685 (N_4685,N_4050,N_4362);
nor U4686 (N_4686,N_4172,N_4202);
or U4687 (N_4687,N_4199,N_4132);
nor U4688 (N_4688,N_4411,N_4400);
or U4689 (N_4689,N_4242,N_4017);
or U4690 (N_4690,N_4185,N_4477);
nand U4691 (N_4691,N_4079,N_4183);
nand U4692 (N_4692,N_4001,N_4313);
or U4693 (N_4693,N_4212,N_4488);
or U4694 (N_4694,N_4367,N_4339);
and U4695 (N_4695,N_4153,N_4080);
nor U4696 (N_4696,N_4368,N_4493);
xnor U4697 (N_4697,N_4340,N_4161);
or U4698 (N_4698,N_4016,N_4225);
nand U4699 (N_4699,N_4203,N_4188);
nand U4700 (N_4700,N_4468,N_4097);
or U4701 (N_4701,N_4110,N_4022);
or U4702 (N_4702,N_4318,N_4388);
and U4703 (N_4703,N_4481,N_4292);
nand U4704 (N_4704,N_4364,N_4109);
or U4705 (N_4705,N_4446,N_4320);
nor U4706 (N_4706,N_4020,N_4152);
nand U4707 (N_4707,N_4083,N_4240);
and U4708 (N_4708,N_4166,N_4201);
and U4709 (N_4709,N_4093,N_4034);
and U4710 (N_4710,N_4104,N_4107);
nor U4711 (N_4711,N_4271,N_4391);
and U4712 (N_4712,N_4048,N_4329);
or U4713 (N_4713,N_4108,N_4433);
and U4714 (N_4714,N_4470,N_4479);
and U4715 (N_4715,N_4495,N_4194);
nand U4716 (N_4716,N_4461,N_4044);
and U4717 (N_4717,N_4333,N_4300);
and U4718 (N_4718,N_4335,N_4326);
or U4719 (N_4719,N_4404,N_4358);
nor U4720 (N_4720,N_4103,N_4405);
and U4721 (N_4721,N_4322,N_4266);
or U4722 (N_4722,N_4142,N_4467);
or U4723 (N_4723,N_4074,N_4336);
nand U4724 (N_4724,N_4328,N_4054);
nor U4725 (N_4725,N_4033,N_4402);
nor U4726 (N_4726,N_4178,N_4394);
and U4727 (N_4727,N_4164,N_4128);
nand U4728 (N_4728,N_4304,N_4158);
or U4729 (N_4729,N_4141,N_4105);
and U4730 (N_4730,N_4115,N_4296);
xor U4731 (N_4731,N_4317,N_4451);
nand U4732 (N_4732,N_4331,N_4215);
or U4733 (N_4733,N_4256,N_4432);
and U4734 (N_4734,N_4311,N_4382);
nor U4735 (N_4735,N_4032,N_4241);
nor U4736 (N_4736,N_4092,N_4075);
and U4737 (N_4737,N_4306,N_4369);
or U4738 (N_4738,N_4238,N_4474);
and U4739 (N_4739,N_4168,N_4133);
nand U4740 (N_4740,N_4286,N_4392);
and U4741 (N_4741,N_4149,N_4136);
nor U4742 (N_4742,N_4068,N_4269);
nor U4743 (N_4743,N_4489,N_4224);
or U4744 (N_4744,N_4086,N_4213);
nand U4745 (N_4745,N_4169,N_4146);
or U4746 (N_4746,N_4445,N_4019);
nor U4747 (N_4747,N_4348,N_4081);
nor U4748 (N_4748,N_4332,N_4293);
nand U4749 (N_4749,N_4350,N_4005);
or U4750 (N_4750,N_4479,N_4155);
nor U4751 (N_4751,N_4330,N_4001);
nor U4752 (N_4752,N_4402,N_4019);
and U4753 (N_4753,N_4266,N_4149);
or U4754 (N_4754,N_4483,N_4448);
nor U4755 (N_4755,N_4252,N_4240);
or U4756 (N_4756,N_4489,N_4495);
nand U4757 (N_4757,N_4019,N_4038);
nand U4758 (N_4758,N_4164,N_4043);
nand U4759 (N_4759,N_4163,N_4141);
and U4760 (N_4760,N_4013,N_4321);
or U4761 (N_4761,N_4338,N_4031);
or U4762 (N_4762,N_4354,N_4256);
and U4763 (N_4763,N_4450,N_4086);
nand U4764 (N_4764,N_4273,N_4479);
nand U4765 (N_4765,N_4429,N_4426);
nand U4766 (N_4766,N_4139,N_4086);
and U4767 (N_4767,N_4448,N_4179);
or U4768 (N_4768,N_4231,N_4392);
nand U4769 (N_4769,N_4118,N_4157);
nand U4770 (N_4770,N_4133,N_4420);
or U4771 (N_4771,N_4447,N_4050);
and U4772 (N_4772,N_4073,N_4489);
nor U4773 (N_4773,N_4045,N_4096);
nor U4774 (N_4774,N_4081,N_4294);
nor U4775 (N_4775,N_4033,N_4449);
nand U4776 (N_4776,N_4354,N_4305);
nor U4777 (N_4777,N_4364,N_4352);
or U4778 (N_4778,N_4386,N_4354);
and U4779 (N_4779,N_4048,N_4482);
nand U4780 (N_4780,N_4201,N_4493);
and U4781 (N_4781,N_4429,N_4059);
and U4782 (N_4782,N_4298,N_4373);
or U4783 (N_4783,N_4242,N_4331);
nand U4784 (N_4784,N_4095,N_4005);
or U4785 (N_4785,N_4473,N_4186);
nand U4786 (N_4786,N_4305,N_4172);
and U4787 (N_4787,N_4292,N_4230);
nand U4788 (N_4788,N_4083,N_4029);
and U4789 (N_4789,N_4071,N_4342);
nor U4790 (N_4790,N_4370,N_4419);
nand U4791 (N_4791,N_4000,N_4200);
or U4792 (N_4792,N_4163,N_4009);
nand U4793 (N_4793,N_4480,N_4090);
and U4794 (N_4794,N_4036,N_4059);
nand U4795 (N_4795,N_4407,N_4324);
nand U4796 (N_4796,N_4269,N_4366);
and U4797 (N_4797,N_4281,N_4129);
nand U4798 (N_4798,N_4456,N_4132);
and U4799 (N_4799,N_4371,N_4432);
xor U4800 (N_4800,N_4225,N_4490);
nor U4801 (N_4801,N_4312,N_4263);
nand U4802 (N_4802,N_4466,N_4285);
nor U4803 (N_4803,N_4388,N_4094);
nand U4804 (N_4804,N_4498,N_4203);
nand U4805 (N_4805,N_4420,N_4352);
nor U4806 (N_4806,N_4209,N_4096);
and U4807 (N_4807,N_4396,N_4324);
nand U4808 (N_4808,N_4376,N_4059);
or U4809 (N_4809,N_4397,N_4334);
nand U4810 (N_4810,N_4259,N_4102);
nor U4811 (N_4811,N_4453,N_4494);
and U4812 (N_4812,N_4017,N_4433);
nor U4813 (N_4813,N_4192,N_4457);
or U4814 (N_4814,N_4027,N_4397);
or U4815 (N_4815,N_4414,N_4258);
nand U4816 (N_4816,N_4496,N_4435);
and U4817 (N_4817,N_4118,N_4252);
nand U4818 (N_4818,N_4460,N_4282);
nand U4819 (N_4819,N_4292,N_4456);
nand U4820 (N_4820,N_4023,N_4108);
and U4821 (N_4821,N_4199,N_4253);
nand U4822 (N_4822,N_4273,N_4476);
nand U4823 (N_4823,N_4312,N_4211);
nand U4824 (N_4824,N_4114,N_4427);
nand U4825 (N_4825,N_4060,N_4110);
and U4826 (N_4826,N_4443,N_4456);
nand U4827 (N_4827,N_4088,N_4353);
or U4828 (N_4828,N_4317,N_4434);
or U4829 (N_4829,N_4180,N_4135);
nand U4830 (N_4830,N_4219,N_4450);
nand U4831 (N_4831,N_4401,N_4165);
nand U4832 (N_4832,N_4124,N_4413);
nand U4833 (N_4833,N_4206,N_4314);
or U4834 (N_4834,N_4226,N_4038);
and U4835 (N_4835,N_4044,N_4065);
nor U4836 (N_4836,N_4294,N_4264);
nor U4837 (N_4837,N_4417,N_4264);
xnor U4838 (N_4838,N_4418,N_4336);
nor U4839 (N_4839,N_4278,N_4326);
and U4840 (N_4840,N_4385,N_4421);
or U4841 (N_4841,N_4310,N_4361);
nand U4842 (N_4842,N_4391,N_4178);
and U4843 (N_4843,N_4432,N_4081);
nor U4844 (N_4844,N_4447,N_4157);
and U4845 (N_4845,N_4317,N_4245);
nand U4846 (N_4846,N_4388,N_4070);
nand U4847 (N_4847,N_4230,N_4413);
or U4848 (N_4848,N_4172,N_4149);
nor U4849 (N_4849,N_4197,N_4250);
and U4850 (N_4850,N_4132,N_4461);
nor U4851 (N_4851,N_4433,N_4456);
and U4852 (N_4852,N_4012,N_4177);
nand U4853 (N_4853,N_4057,N_4041);
or U4854 (N_4854,N_4012,N_4150);
and U4855 (N_4855,N_4409,N_4101);
nor U4856 (N_4856,N_4295,N_4260);
or U4857 (N_4857,N_4321,N_4012);
nor U4858 (N_4858,N_4311,N_4437);
nor U4859 (N_4859,N_4104,N_4174);
or U4860 (N_4860,N_4452,N_4274);
nand U4861 (N_4861,N_4037,N_4248);
nor U4862 (N_4862,N_4151,N_4361);
nand U4863 (N_4863,N_4191,N_4112);
nand U4864 (N_4864,N_4053,N_4163);
or U4865 (N_4865,N_4034,N_4486);
nand U4866 (N_4866,N_4268,N_4211);
or U4867 (N_4867,N_4179,N_4143);
and U4868 (N_4868,N_4170,N_4302);
or U4869 (N_4869,N_4026,N_4042);
and U4870 (N_4870,N_4426,N_4273);
nor U4871 (N_4871,N_4144,N_4399);
xnor U4872 (N_4872,N_4163,N_4069);
or U4873 (N_4873,N_4452,N_4455);
nor U4874 (N_4874,N_4133,N_4145);
nand U4875 (N_4875,N_4348,N_4002);
or U4876 (N_4876,N_4479,N_4233);
or U4877 (N_4877,N_4193,N_4095);
nand U4878 (N_4878,N_4244,N_4150);
and U4879 (N_4879,N_4320,N_4250);
or U4880 (N_4880,N_4449,N_4120);
or U4881 (N_4881,N_4363,N_4233);
nand U4882 (N_4882,N_4468,N_4332);
nor U4883 (N_4883,N_4007,N_4108);
or U4884 (N_4884,N_4499,N_4131);
and U4885 (N_4885,N_4451,N_4205);
nor U4886 (N_4886,N_4297,N_4475);
and U4887 (N_4887,N_4395,N_4306);
nor U4888 (N_4888,N_4092,N_4174);
nand U4889 (N_4889,N_4376,N_4399);
and U4890 (N_4890,N_4193,N_4031);
nor U4891 (N_4891,N_4395,N_4299);
nor U4892 (N_4892,N_4221,N_4317);
or U4893 (N_4893,N_4459,N_4040);
nand U4894 (N_4894,N_4066,N_4299);
nor U4895 (N_4895,N_4264,N_4346);
nor U4896 (N_4896,N_4133,N_4405);
nor U4897 (N_4897,N_4180,N_4303);
or U4898 (N_4898,N_4076,N_4234);
nor U4899 (N_4899,N_4342,N_4131);
and U4900 (N_4900,N_4054,N_4343);
nor U4901 (N_4901,N_4077,N_4023);
or U4902 (N_4902,N_4404,N_4457);
nand U4903 (N_4903,N_4225,N_4209);
and U4904 (N_4904,N_4345,N_4316);
and U4905 (N_4905,N_4320,N_4211);
and U4906 (N_4906,N_4088,N_4329);
or U4907 (N_4907,N_4101,N_4137);
nor U4908 (N_4908,N_4276,N_4293);
nor U4909 (N_4909,N_4109,N_4158);
and U4910 (N_4910,N_4143,N_4174);
or U4911 (N_4911,N_4101,N_4050);
and U4912 (N_4912,N_4436,N_4298);
or U4913 (N_4913,N_4386,N_4296);
nor U4914 (N_4914,N_4135,N_4395);
nor U4915 (N_4915,N_4420,N_4387);
or U4916 (N_4916,N_4299,N_4244);
nand U4917 (N_4917,N_4077,N_4253);
nand U4918 (N_4918,N_4153,N_4247);
and U4919 (N_4919,N_4356,N_4449);
and U4920 (N_4920,N_4208,N_4366);
nor U4921 (N_4921,N_4356,N_4498);
and U4922 (N_4922,N_4280,N_4241);
nand U4923 (N_4923,N_4252,N_4479);
or U4924 (N_4924,N_4422,N_4471);
and U4925 (N_4925,N_4099,N_4497);
and U4926 (N_4926,N_4099,N_4260);
nand U4927 (N_4927,N_4181,N_4183);
nor U4928 (N_4928,N_4064,N_4255);
nor U4929 (N_4929,N_4160,N_4273);
or U4930 (N_4930,N_4066,N_4487);
or U4931 (N_4931,N_4474,N_4166);
nand U4932 (N_4932,N_4427,N_4084);
nor U4933 (N_4933,N_4145,N_4296);
nor U4934 (N_4934,N_4297,N_4403);
nor U4935 (N_4935,N_4475,N_4256);
and U4936 (N_4936,N_4001,N_4146);
or U4937 (N_4937,N_4055,N_4370);
nand U4938 (N_4938,N_4050,N_4266);
xnor U4939 (N_4939,N_4112,N_4133);
nor U4940 (N_4940,N_4291,N_4249);
nor U4941 (N_4941,N_4295,N_4098);
and U4942 (N_4942,N_4452,N_4174);
or U4943 (N_4943,N_4005,N_4261);
and U4944 (N_4944,N_4237,N_4160);
nor U4945 (N_4945,N_4170,N_4008);
or U4946 (N_4946,N_4455,N_4494);
nand U4947 (N_4947,N_4108,N_4088);
nor U4948 (N_4948,N_4336,N_4013);
nand U4949 (N_4949,N_4098,N_4182);
or U4950 (N_4950,N_4079,N_4056);
or U4951 (N_4951,N_4018,N_4472);
nand U4952 (N_4952,N_4484,N_4074);
and U4953 (N_4953,N_4045,N_4063);
nand U4954 (N_4954,N_4496,N_4030);
and U4955 (N_4955,N_4403,N_4075);
or U4956 (N_4956,N_4427,N_4346);
nor U4957 (N_4957,N_4138,N_4411);
nor U4958 (N_4958,N_4482,N_4348);
or U4959 (N_4959,N_4417,N_4158);
nor U4960 (N_4960,N_4365,N_4234);
nand U4961 (N_4961,N_4149,N_4040);
nor U4962 (N_4962,N_4086,N_4460);
nand U4963 (N_4963,N_4218,N_4111);
or U4964 (N_4964,N_4232,N_4152);
nand U4965 (N_4965,N_4021,N_4014);
nand U4966 (N_4966,N_4026,N_4013);
nand U4967 (N_4967,N_4243,N_4456);
nand U4968 (N_4968,N_4343,N_4042);
and U4969 (N_4969,N_4418,N_4066);
nor U4970 (N_4970,N_4125,N_4104);
or U4971 (N_4971,N_4076,N_4358);
nor U4972 (N_4972,N_4069,N_4321);
nand U4973 (N_4973,N_4256,N_4084);
or U4974 (N_4974,N_4470,N_4239);
or U4975 (N_4975,N_4062,N_4012);
nor U4976 (N_4976,N_4494,N_4094);
nor U4977 (N_4977,N_4117,N_4321);
nand U4978 (N_4978,N_4141,N_4042);
nor U4979 (N_4979,N_4472,N_4465);
nand U4980 (N_4980,N_4373,N_4429);
and U4981 (N_4981,N_4393,N_4204);
nor U4982 (N_4982,N_4104,N_4170);
nor U4983 (N_4983,N_4207,N_4358);
and U4984 (N_4984,N_4025,N_4350);
nand U4985 (N_4985,N_4000,N_4449);
or U4986 (N_4986,N_4238,N_4413);
nor U4987 (N_4987,N_4460,N_4391);
or U4988 (N_4988,N_4374,N_4340);
nor U4989 (N_4989,N_4037,N_4061);
or U4990 (N_4990,N_4364,N_4041);
nand U4991 (N_4991,N_4385,N_4313);
nand U4992 (N_4992,N_4007,N_4206);
nor U4993 (N_4993,N_4215,N_4378);
or U4994 (N_4994,N_4281,N_4440);
and U4995 (N_4995,N_4272,N_4136);
and U4996 (N_4996,N_4109,N_4007);
nor U4997 (N_4997,N_4177,N_4383);
and U4998 (N_4998,N_4367,N_4337);
nor U4999 (N_4999,N_4475,N_4315);
or UO_0 (O_0,N_4782,N_4693);
and UO_1 (O_1,N_4646,N_4953);
or UO_2 (O_2,N_4839,N_4948);
nor UO_3 (O_3,N_4518,N_4589);
nand UO_4 (O_4,N_4949,N_4701);
nand UO_5 (O_5,N_4581,N_4885);
and UO_6 (O_6,N_4835,N_4863);
and UO_7 (O_7,N_4592,N_4741);
or UO_8 (O_8,N_4696,N_4932);
or UO_9 (O_9,N_4896,N_4884);
xor UO_10 (O_10,N_4785,N_4814);
or UO_11 (O_11,N_4593,N_4858);
and UO_12 (O_12,N_4594,N_4915);
nand UO_13 (O_13,N_4645,N_4945);
or UO_14 (O_14,N_4745,N_4742);
nor UO_15 (O_15,N_4638,N_4935);
nand UO_16 (O_16,N_4985,N_4982);
nor UO_17 (O_17,N_4610,N_4973);
or UO_18 (O_18,N_4889,N_4801);
nand UO_19 (O_19,N_4923,N_4715);
and UO_20 (O_20,N_4941,N_4606);
and UO_21 (O_21,N_4961,N_4723);
nand UO_22 (O_22,N_4721,N_4841);
nand UO_23 (O_23,N_4920,N_4684);
nor UO_24 (O_24,N_4629,N_4548);
and UO_25 (O_25,N_4910,N_4636);
and UO_26 (O_26,N_4672,N_4882);
nand UO_27 (O_27,N_4978,N_4979);
nor UO_28 (O_28,N_4955,N_4981);
nand UO_29 (O_29,N_4768,N_4544);
or UO_30 (O_30,N_4698,N_4853);
nand UO_31 (O_31,N_4634,N_4954);
nor UO_32 (O_32,N_4632,N_4644);
or UO_33 (O_33,N_4854,N_4588);
or UO_34 (O_34,N_4622,N_4895);
or UO_35 (O_35,N_4578,N_4522);
and UO_36 (O_36,N_4685,N_4603);
and UO_37 (O_37,N_4909,N_4731);
and UO_38 (O_38,N_4877,N_4591);
or UO_39 (O_39,N_4675,N_4735);
nor UO_40 (O_40,N_4535,N_4780);
or UO_41 (O_41,N_4905,N_4706);
nor UO_42 (O_42,N_4859,N_4984);
and UO_43 (O_43,N_4612,N_4605);
nor UO_44 (O_44,N_4702,N_4778);
or UO_45 (O_45,N_4756,N_4989);
or UO_46 (O_46,N_4775,N_4971);
nor UO_47 (O_47,N_4597,N_4680);
nand UO_48 (O_48,N_4669,N_4720);
or UO_49 (O_49,N_4911,N_4837);
nand UO_50 (O_50,N_4618,N_4657);
nand UO_51 (O_51,N_4747,N_4537);
nand UO_52 (O_52,N_4627,N_4808);
or UO_53 (O_53,N_4571,N_4554);
and UO_54 (O_54,N_4956,N_4994);
nor UO_55 (O_55,N_4664,N_4963);
nor UO_56 (O_56,N_4958,N_4766);
nand UO_57 (O_57,N_4861,N_4927);
nand UO_58 (O_58,N_4972,N_4687);
nor UO_59 (O_59,N_4743,N_4897);
nor UO_60 (O_60,N_4648,N_4857);
nor UO_61 (O_61,N_4810,N_4803);
or UO_62 (O_62,N_4543,N_4912);
and UO_63 (O_63,N_4846,N_4893);
nor UO_64 (O_64,N_4812,N_4553);
or UO_65 (O_65,N_4767,N_4898);
nand UO_66 (O_66,N_4582,N_4616);
nand UO_67 (O_67,N_4848,N_4661);
or UO_68 (O_68,N_4565,N_4748);
nor UO_69 (O_69,N_4811,N_4545);
xor UO_70 (O_70,N_4786,N_4541);
or UO_71 (O_71,N_4671,N_4866);
nand UO_72 (O_72,N_4755,N_4753);
nand UO_73 (O_73,N_4650,N_4950);
nand UO_74 (O_74,N_4531,N_4916);
or UO_75 (O_75,N_4962,N_4681);
nand UO_76 (O_76,N_4906,N_4815);
nand UO_77 (O_77,N_4779,N_4770);
nand UO_78 (O_78,N_4580,N_4868);
nand UO_79 (O_79,N_4992,N_4821);
and UO_80 (O_80,N_4934,N_4507);
or UO_81 (O_81,N_4843,N_4744);
nor UO_82 (O_82,N_4523,N_4538);
nor UO_83 (O_83,N_4660,N_4959);
and UO_84 (O_84,N_4809,N_4516);
xor UO_85 (O_85,N_4967,N_4558);
nor UO_86 (O_86,N_4716,N_4668);
and UO_87 (O_87,N_4718,N_4805);
or UO_88 (O_88,N_4762,N_4600);
or UO_89 (O_89,N_4734,N_4506);
nand UO_90 (O_90,N_4813,N_4752);
nand UO_91 (O_91,N_4609,N_4659);
nand UO_92 (O_92,N_4828,N_4595);
and UO_93 (O_93,N_4737,N_4783);
nand UO_94 (O_94,N_4562,N_4880);
nor UO_95 (O_95,N_4765,N_4662);
nand UO_96 (O_96,N_4514,N_4700);
nand UO_97 (O_97,N_4789,N_4567);
and UO_98 (O_98,N_4900,N_4840);
or UO_99 (O_99,N_4930,N_4947);
nor UO_100 (O_100,N_4501,N_4724);
nand UO_101 (O_101,N_4879,N_4823);
and UO_102 (O_102,N_4802,N_4599);
and UO_103 (O_103,N_4876,N_4960);
nand UO_104 (O_104,N_4856,N_4620);
nand UO_105 (O_105,N_4824,N_4980);
and UO_106 (O_106,N_4590,N_4793);
nor UO_107 (O_107,N_4736,N_4740);
nand UO_108 (O_108,N_4678,N_4710);
or UO_109 (O_109,N_4628,N_4951);
nand UO_110 (O_110,N_4561,N_4936);
and UO_111 (O_111,N_4851,N_4942);
nand UO_112 (O_112,N_4804,N_4692);
and UO_113 (O_113,N_4864,N_4583);
or UO_114 (O_114,N_4642,N_4845);
and UO_115 (O_115,N_4750,N_4826);
and UO_116 (O_116,N_4707,N_4625);
or UO_117 (O_117,N_4760,N_4933);
or UO_118 (O_118,N_4695,N_4873);
or UO_119 (O_119,N_4509,N_4820);
nand UO_120 (O_120,N_4795,N_4774);
nand UO_121 (O_121,N_4528,N_4704);
and UO_122 (O_122,N_4919,N_4536);
and UO_123 (O_123,N_4502,N_4844);
or UO_124 (O_124,N_4635,N_4943);
or UO_125 (O_125,N_4623,N_4777);
nand UO_126 (O_126,N_4519,N_4639);
and UO_127 (O_127,N_4727,N_4568);
and UO_128 (O_128,N_4527,N_4990);
nand UO_129 (O_129,N_4656,N_4913);
nor UO_130 (O_130,N_4862,N_4987);
or UO_131 (O_131,N_4673,N_4529);
nand UO_132 (O_132,N_4914,N_4974);
nand UO_133 (O_133,N_4799,N_4559);
and UO_134 (O_134,N_4577,N_4574);
and UO_135 (O_135,N_4572,N_4907);
nand UO_136 (O_136,N_4686,N_4887);
and UO_137 (O_137,N_4834,N_4924);
or UO_138 (O_138,N_4511,N_4938);
nand UO_139 (O_139,N_4998,N_4886);
nand UO_140 (O_140,N_4641,N_4613);
or UO_141 (O_141,N_4878,N_4822);
and UO_142 (O_142,N_4763,N_4643);
nor UO_143 (O_143,N_4991,N_4560);
nand UO_144 (O_144,N_4689,N_4533);
nand UO_145 (O_145,N_4557,N_4831);
or UO_146 (O_146,N_4520,N_4530);
nand UO_147 (O_147,N_4792,N_4807);
nand UO_148 (O_148,N_4626,N_4794);
or UO_149 (O_149,N_4546,N_4649);
or UO_150 (O_150,N_4798,N_4827);
nor UO_151 (O_151,N_4607,N_4819);
and UO_152 (O_152,N_4637,N_4739);
nor UO_153 (O_153,N_4892,N_4573);
and UO_154 (O_154,N_4764,N_4564);
nor UO_155 (O_155,N_4719,N_4711);
nor UO_156 (O_156,N_4587,N_4615);
nand UO_157 (O_157,N_4504,N_4881);
and UO_158 (O_158,N_4838,N_4703);
xor UO_159 (O_159,N_4630,N_4797);
nor UO_160 (O_160,N_4926,N_4850);
nor UO_161 (O_161,N_4539,N_4852);
nand UO_162 (O_162,N_4829,N_4633);
or UO_163 (O_163,N_4904,N_4771);
and UO_164 (O_164,N_4818,N_4966);
and UO_165 (O_165,N_4601,N_4705);
nand UO_166 (O_166,N_4849,N_4526);
nor UO_167 (O_167,N_4749,N_4901);
nor UO_168 (O_168,N_4697,N_4517);
and UO_169 (O_169,N_4883,N_4902);
and UO_170 (O_170,N_4655,N_4776);
or UO_171 (O_171,N_4746,N_4722);
and UO_172 (O_172,N_4570,N_4510);
nand UO_173 (O_173,N_4865,N_4617);
or UO_174 (O_174,N_4796,N_4872);
or UO_175 (O_175,N_4658,N_4917);
or UO_176 (O_176,N_4817,N_4759);
or UO_177 (O_177,N_4874,N_4946);
nand UO_178 (O_178,N_4758,N_4891);
or UO_179 (O_179,N_4761,N_4908);
nor UO_180 (O_180,N_4997,N_4729);
and UO_181 (O_181,N_4683,N_4717);
and UO_182 (O_182,N_4732,N_4647);
or UO_183 (O_183,N_4550,N_4787);
nand UO_184 (O_184,N_4993,N_4624);
or UO_185 (O_185,N_4754,N_4791);
nand UO_186 (O_186,N_4772,N_4730);
nor UO_187 (O_187,N_4503,N_4556);
and UO_188 (O_188,N_4922,N_4944);
or UO_189 (O_189,N_4757,N_4604);
and UO_190 (O_190,N_4965,N_4769);
or UO_191 (O_191,N_4585,N_4842);
nand UO_192 (O_192,N_4690,N_4576);
nor UO_193 (O_193,N_4894,N_4569);
nand UO_194 (O_194,N_4800,N_4988);
nor UO_195 (O_195,N_4726,N_4832);
nand UO_196 (O_196,N_4670,N_4547);
nor UO_197 (O_197,N_4552,N_4855);
and UO_198 (O_198,N_4712,N_4867);
and UO_199 (O_199,N_4733,N_4970);
nor UO_200 (O_200,N_4555,N_4999);
and UO_201 (O_201,N_4875,N_4709);
or UO_202 (O_202,N_4534,N_4977);
nand UO_203 (O_203,N_4964,N_4521);
and UO_204 (O_204,N_4666,N_4513);
or UO_205 (O_205,N_4563,N_4677);
or UO_206 (O_206,N_4738,N_4929);
nor UO_207 (O_207,N_4586,N_4674);
nand UO_208 (O_208,N_4512,N_4694);
nor UO_209 (O_209,N_4596,N_4957);
and UO_210 (O_210,N_4871,N_4784);
and UO_211 (O_211,N_4983,N_4751);
and UO_212 (O_212,N_4676,N_4614);
or UO_213 (O_213,N_4725,N_4969);
nor UO_214 (O_214,N_4975,N_4781);
nor UO_215 (O_215,N_4621,N_4691);
or UO_216 (O_216,N_4825,N_4699);
or UO_217 (O_217,N_4714,N_4816);
or UO_218 (O_218,N_4663,N_4654);
or UO_219 (O_219,N_4939,N_4566);
xor UO_220 (O_220,N_4995,N_4652);
nor UO_221 (O_221,N_4602,N_4903);
and UO_222 (O_222,N_4640,N_4688);
or UO_223 (O_223,N_4833,N_4505);
and UO_224 (O_224,N_4925,N_4870);
nor UO_225 (O_225,N_4525,N_4682);
nand UO_226 (O_226,N_4500,N_4899);
and UO_227 (O_227,N_4708,N_4551);
or UO_228 (O_228,N_4611,N_4524);
nand UO_229 (O_229,N_4540,N_4542);
nor UO_230 (O_230,N_4836,N_4788);
and UO_231 (O_231,N_4619,N_4830);
or UO_232 (O_232,N_4773,N_4532);
nor UO_233 (O_233,N_4790,N_4549);
and UO_234 (O_234,N_4986,N_4921);
or UO_235 (O_235,N_4890,N_4847);
and UO_236 (O_236,N_4679,N_4508);
or UO_237 (O_237,N_4968,N_4918);
and UO_238 (O_238,N_4728,N_4515);
and UO_239 (O_239,N_4928,N_4631);
nand UO_240 (O_240,N_4667,N_4869);
nand UO_241 (O_241,N_4931,N_4665);
nand UO_242 (O_242,N_4584,N_4976);
nand UO_243 (O_243,N_4713,N_4937);
and UO_244 (O_244,N_4579,N_4888);
nor UO_245 (O_245,N_4598,N_4575);
nor UO_246 (O_246,N_4940,N_4651);
and UO_247 (O_247,N_4653,N_4860);
and UO_248 (O_248,N_4806,N_4996);
nand UO_249 (O_249,N_4608,N_4952);
nand UO_250 (O_250,N_4659,N_4736);
nor UO_251 (O_251,N_4748,N_4596);
nand UO_252 (O_252,N_4544,N_4580);
nand UO_253 (O_253,N_4879,N_4583);
nand UO_254 (O_254,N_4930,N_4844);
and UO_255 (O_255,N_4990,N_4501);
nor UO_256 (O_256,N_4827,N_4716);
or UO_257 (O_257,N_4794,N_4750);
nor UO_258 (O_258,N_4522,N_4796);
or UO_259 (O_259,N_4724,N_4682);
nand UO_260 (O_260,N_4846,N_4675);
nand UO_261 (O_261,N_4654,N_4729);
nand UO_262 (O_262,N_4512,N_4962);
or UO_263 (O_263,N_4798,N_4978);
nand UO_264 (O_264,N_4975,N_4849);
nand UO_265 (O_265,N_4823,N_4501);
and UO_266 (O_266,N_4922,N_4645);
or UO_267 (O_267,N_4839,N_4900);
and UO_268 (O_268,N_4504,N_4519);
and UO_269 (O_269,N_4586,N_4940);
nor UO_270 (O_270,N_4751,N_4556);
nor UO_271 (O_271,N_4988,N_4908);
and UO_272 (O_272,N_4507,N_4692);
and UO_273 (O_273,N_4802,N_4591);
and UO_274 (O_274,N_4927,N_4699);
nand UO_275 (O_275,N_4508,N_4759);
or UO_276 (O_276,N_4638,N_4585);
and UO_277 (O_277,N_4949,N_4733);
or UO_278 (O_278,N_4739,N_4723);
and UO_279 (O_279,N_4800,N_4978);
nand UO_280 (O_280,N_4611,N_4688);
nand UO_281 (O_281,N_4703,N_4713);
nand UO_282 (O_282,N_4584,N_4774);
or UO_283 (O_283,N_4608,N_4667);
and UO_284 (O_284,N_4757,N_4821);
or UO_285 (O_285,N_4817,N_4907);
and UO_286 (O_286,N_4680,N_4690);
or UO_287 (O_287,N_4502,N_4984);
or UO_288 (O_288,N_4804,N_4799);
or UO_289 (O_289,N_4603,N_4756);
nor UO_290 (O_290,N_4771,N_4621);
and UO_291 (O_291,N_4895,N_4974);
and UO_292 (O_292,N_4568,N_4625);
nor UO_293 (O_293,N_4710,N_4783);
and UO_294 (O_294,N_4694,N_4858);
nor UO_295 (O_295,N_4766,N_4811);
nand UO_296 (O_296,N_4752,N_4606);
or UO_297 (O_297,N_4809,N_4757);
or UO_298 (O_298,N_4871,N_4692);
and UO_299 (O_299,N_4550,N_4844);
nor UO_300 (O_300,N_4598,N_4596);
and UO_301 (O_301,N_4921,N_4942);
nor UO_302 (O_302,N_4868,N_4792);
nor UO_303 (O_303,N_4917,N_4896);
or UO_304 (O_304,N_4534,N_4624);
nand UO_305 (O_305,N_4672,N_4782);
and UO_306 (O_306,N_4961,N_4553);
nand UO_307 (O_307,N_4689,N_4710);
nor UO_308 (O_308,N_4679,N_4756);
or UO_309 (O_309,N_4992,N_4899);
or UO_310 (O_310,N_4710,N_4872);
nor UO_311 (O_311,N_4673,N_4570);
and UO_312 (O_312,N_4894,N_4952);
nor UO_313 (O_313,N_4753,N_4877);
nor UO_314 (O_314,N_4559,N_4937);
or UO_315 (O_315,N_4755,N_4775);
or UO_316 (O_316,N_4971,N_4779);
and UO_317 (O_317,N_4563,N_4541);
nor UO_318 (O_318,N_4601,N_4570);
and UO_319 (O_319,N_4650,N_4608);
or UO_320 (O_320,N_4791,N_4591);
and UO_321 (O_321,N_4984,N_4819);
nand UO_322 (O_322,N_4510,N_4908);
nand UO_323 (O_323,N_4781,N_4639);
nand UO_324 (O_324,N_4670,N_4858);
nor UO_325 (O_325,N_4805,N_4844);
and UO_326 (O_326,N_4997,N_4902);
nor UO_327 (O_327,N_4739,N_4954);
or UO_328 (O_328,N_4682,N_4683);
and UO_329 (O_329,N_4766,N_4728);
nand UO_330 (O_330,N_4847,N_4817);
nand UO_331 (O_331,N_4863,N_4759);
nand UO_332 (O_332,N_4693,N_4760);
nor UO_333 (O_333,N_4588,N_4836);
nand UO_334 (O_334,N_4728,N_4966);
or UO_335 (O_335,N_4973,N_4538);
or UO_336 (O_336,N_4785,N_4890);
nor UO_337 (O_337,N_4971,N_4803);
or UO_338 (O_338,N_4870,N_4835);
nand UO_339 (O_339,N_4768,N_4526);
and UO_340 (O_340,N_4924,N_4830);
nor UO_341 (O_341,N_4715,N_4516);
nor UO_342 (O_342,N_4543,N_4723);
or UO_343 (O_343,N_4635,N_4740);
nor UO_344 (O_344,N_4719,N_4907);
nor UO_345 (O_345,N_4592,N_4979);
nor UO_346 (O_346,N_4856,N_4948);
nand UO_347 (O_347,N_4595,N_4931);
and UO_348 (O_348,N_4694,N_4725);
nand UO_349 (O_349,N_4657,N_4663);
and UO_350 (O_350,N_4839,N_4560);
and UO_351 (O_351,N_4843,N_4696);
nand UO_352 (O_352,N_4980,N_4807);
or UO_353 (O_353,N_4588,N_4555);
xor UO_354 (O_354,N_4822,N_4519);
nor UO_355 (O_355,N_4521,N_4890);
or UO_356 (O_356,N_4874,N_4895);
or UO_357 (O_357,N_4690,N_4580);
nand UO_358 (O_358,N_4501,N_4713);
nand UO_359 (O_359,N_4877,N_4775);
and UO_360 (O_360,N_4662,N_4892);
and UO_361 (O_361,N_4906,N_4638);
nand UO_362 (O_362,N_4858,N_4798);
nand UO_363 (O_363,N_4664,N_4989);
and UO_364 (O_364,N_4625,N_4827);
nand UO_365 (O_365,N_4756,N_4544);
nor UO_366 (O_366,N_4539,N_4789);
or UO_367 (O_367,N_4963,N_4634);
and UO_368 (O_368,N_4565,N_4903);
or UO_369 (O_369,N_4554,N_4507);
nand UO_370 (O_370,N_4978,N_4658);
nand UO_371 (O_371,N_4959,N_4659);
and UO_372 (O_372,N_4616,N_4791);
and UO_373 (O_373,N_4808,N_4994);
or UO_374 (O_374,N_4720,N_4989);
and UO_375 (O_375,N_4968,N_4826);
nor UO_376 (O_376,N_4596,N_4529);
and UO_377 (O_377,N_4766,N_4608);
nor UO_378 (O_378,N_4676,N_4816);
or UO_379 (O_379,N_4990,N_4807);
nor UO_380 (O_380,N_4854,N_4870);
nand UO_381 (O_381,N_4648,N_4657);
nor UO_382 (O_382,N_4889,N_4827);
nor UO_383 (O_383,N_4630,N_4647);
nor UO_384 (O_384,N_4726,N_4751);
or UO_385 (O_385,N_4870,N_4648);
or UO_386 (O_386,N_4531,N_4500);
nor UO_387 (O_387,N_4561,N_4532);
or UO_388 (O_388,N_4687,N_4731);
and UO_389 (O_389,N_4594,N_4925);
nor UO_390 (O_390,N_4851,N_4863);
or UO_391 (O_391,N_4666,N_4916);
nor UO_392 (O_392,N_4966,N_4950);
nor UO_393 (O_393,N_4699,N_4834);
nor UO_394 (O_394,N_4598,N_4537);
or UO_395 (O_395,N_4707,N_4572);
nand UO_396 (O_396,N_4931,N_4740);
and UO_397 (O_397,N_4970,N_4714);
or UO_398 (O_398,N_4919,N_4955);
nor UO_399 (O_399,N_4977,N_4908);
nor UO_400 (O_400,N_4617,N_4924);
or UO_401 (O_401,N_4956,N_4550);
and UO_402 (O_402,N_4885,N_4988);
nor UO_403 (O_403,N_4741,N_4887);
and UO_404 (O_404,N_4983,N_4871);
nand UO_405 (O_405,N_4593,N_4610);
or UO_406 (O_406,N_4874,N_4720);
nand UO_407 (O_407,N_4706,N_4946);
nand UO_408 (O_408,N_4587,N_4715);
nand UO_409 (O_409,N_4554,N_4760);
nor UO_410 (O_410,N_4579,N_4683);
and UO_411 (O_411,N_4537,N_4613);
nor UO_412 (O_412,N_4763,N_4908);
and UO_413 (O_413,N_4533,N_4717);
nand UO_414 (O_414,N_4637,N_4860);
nand UO_415 (O_415,N_4828,N_4621);
and UO_416 (O_416,N_4548,N_4589);
nor UO_417 (O_417,N_4997,N_4726);
or UO_418 (O_418,N_4816,N_4869);
nor UO_419 (O_419,N_4644,N_4675);
nor UO_420 (O_420,N_4849,N_4642);
and UO_421 (O_421,N_4706,N_4916);
nor UO_422 (O_422,N_4789,N_4505);
or UO_423 (O_423,N_4941,N_4848);
and UO_424 (O_424,N_4530,N_4558);
nand UO_425 (O_425,N_4656,N_4848);
and UO_426 (O_426,N_4835,N_4670);
and UO_427 (O_427,N_4750,N_4515);
nor UO_428 (O_428,N_4716,N_4675);
and UO_429 (O_429,N_4723,N_4888);
nor UO_430 (O_430,N_4619,N_4597);
and UO_431 (O_431,N_4725,N_4783);
or UO_432 (O_432,N_4962,N_4798);
and UO_433 (O_433,N_4731,N_4915);
nor UO_434 (O_434,N_4505,N_4915);
nor UO_435 (O_435,N_4940,N_4579);
or UO_436 (O_436,N_4887,N_4629);
nor UO_437 (O_437,N_4677,N_4939);
nand UO_438 (O_438,N_4900,N_4825);
and UO_439 (O_439,N_4729,N_4951);
nor UO_440 (O_440,N_4886,N_4733);
or UO_441 (O_441,N_4930,N_4566);
or UO_442 (O_442,N_4992,N_4758);
nand UO_443 (O_443,N_4919,N_4800);
and UO_444 (O_444,N_4950,N_4663);
or UO_445 (O_445,N_4520,N_4592);
nand UO_446 (O_446,N_4810,N_4522);
nand UO_447 (O_447,N_4942,N_4989);
or UO_448 (O_448,N_4784,N_4523);
nand UO_449 (O_449,N_4727,N_4541);
or UO_450 (O_450,N_4569,N_4645);
and UO_451 (O_451,N_4683,N_4845);
or UO_452 (O_452,N_4655,N_4986);
or UO_453 (O_453,N_4577,N_4534);
nor UO_454 (O_454,N_4782,N_4661);
nand UO_455 (O_455,N_4957,N_4760);
nand UO_456 (O_456,N_4750,N_4874);
and UO_457 (O_457,N_4744,N_4760);
and UO_458 (O_458,N_4565,N_4713);
nor UO_459 (O_459,N_4947,N_4884);
nor UO_460 (O_460,N_4512,N_4578);
or UO_461 (O_461,N_4739,N_4525);
nor UO_462 (O_462,N_4508,N_4580);
nor UO_463 (O_463,N_4705,N_4837);
or UO_464 (O_464,N_4768,N_4842);
nor UO_465 (O_465,N_4819,N_4529);
and UO_466 (O_466,N_4968,N_4706);
nor UO_467 (O_467,N_4533,N_4939);
nand UO_468 (O_468,N_4671,N_4592);
nand UO_469 (O_469,N_4575,N_4521);
nor UO_470 (O_470,N_4745,N_4667);
nand UO_471 (O_471,N_4691,N_4832);
nor UO_472 (O_472,N_4918,N_4979);
and UO_473 (O_473,N_4838,N_4766);
nand UO_474 (O_474,N_4951,N_4639);
or UO_475 (O_475,N_4904,N_4970);
or UO_476 (O_476,N_4838,N_4769);
or UO_477 (O_477,N_4676,N_4952);
nand UO_478 (O_478,N_4955,N_4877);
nand UO_479 (O_479,N_4665,N_4791);
nand UO_480 (O_480,N_4849,N_4617);
and UO_481 (O_481,N_4513,N_4680);
xor UO_482 (O_482,N_4688,N_4683);
or UO_483 (O_483,N_4991,N_4788);
nor UO_484 (O_484,N_4695,N_4546);
and UO_485 (O_485,N_4600,N_4986);
nor UO_486 (O_486,N_4787,N_4523);
nand UO_487 (O_487,N_4844,N_4656);
nand UO_488 (O_488,N_4772,N_4816);
nand UO_489 (O_489,N_4619,N_4717);
and UO_490 (O_490,N_4964,N_4793);
nor UO_491 (O_491,N_4568,N_4511);
xor UO_492 (O_492,N_4501,N_4750);
nor UO_493 (O_493,N_4571,N_4730);
nand UO_494 (O_494,N_4659,N_4860);
nor UO_495 (O_495,N_4949,N_4593);
and UO_496 (O_496,N_4955,N_4528);
and UO_497 (O_497,N_4993,N_4714);
or UO_498 (O_498,N_4619,N_4515);
or UO_499 (O_499,N_4876,N_4698);
and UO_500 (O_500,N_4651,N_4723);
nor UO_501 (O_501,N_4860,N_4780);
nor UO_502 (O_502,N_4511,N_4811);
nand UO_503 (O_503,N_4864,N_4767);
or UO_504 (O_504,N_4738,N_4648);
nand UO_505 (O_505,N_4785,N_4816);
and UO_506 (O_506,N_4871,N_4969);
nand UO_507 (O_507,N_4874,N_4734);
or UO_508 (O_508,N_4543,N_4803);
and UO_509 (O_509,N_4929,N_4961);
nand UO_510 (O_510,N_4699,N_4637);
and UO_511 (O_511,N_4866,N_4619);
and UO_512 (O_512,N_4992,N_4857);
nor UO_513 (O_513,N_4849,N_4993);
nor UO_514 (O_514,N_4532,N_4898);
and UO_515 (O_515,N_4617,N_4843);
or UO_516 (O_516,N_4603,N_4845);
or UO_517 (O_517,N_4686,N_4575);
nand UO_518 (O_518,N_4898,N_4885);
or UO_519 (O_519,N_4803,N_4763);
and UO_520 (O_520,N_4823,N_4857);
nand UO_521 (O_521,N_4785,N_4545);
nand UO_522 (O_522,N_4774,N_4571);
and UO_523 (O_523,N_4899,N_4767);
and UO_524 (O_524,N_4936,N_4943);
nand UO_525 (O_525,N_4770,N_4660);
and UO_526 (O_526,N_4907,N_4687);
or UO_527 (O_527,N_4918,N_4727);
and UO_528 (O_528,N_4832,N_4839);
or UO_529 (O_529,N_4758,N_4606);
and UO_530 (O_530,N_4648,N_4515);
or UO_531 (O_531,N_4782,N_4692);
xor UO_532 (O_532,N_4683,N_4788);
and UO_533 (O_533,N_4894,N_4857);
nand UO_534 (O_534,N_4857,N_4839);
nand UO_535 (O_535,N_4990,N_4993);
and UO_536 (O_536,N_4519,N_4705);
and UO_537 (O_537,N_4894,N_4743);
and UO_538 (O_538,N_4865,N_4641);
nor UO_539 (O_539,N_4674,N_4649);
nor UO_540 (O_540,N_4691,N_4565);
or UO_541 (O_541,N_4895,N_4634);
and UO_542 (O_542,N_4579,N_4892);
nor UO_543 (O_543,N_4973,N_4951);
nand UO_544 (O_544,N_4962,N_4813);
nand UO_545 (O_545,N_4685,N_4562);
or UO_546 (O_546,N_4712,N_4588);
xor UO_547 (O_547,N_4948,N_4705);
nor UO_548 (O_548,N_4885,N_4517);
nand UO_549 (O_549,N_4657,N_4590);
nor UO_550 (O_550,N_4902,N_4867);
nor UO_551 (O_551,N_4606,N_4578);
and UO_552 (O_552,N_4716,N_4705);
or UO_553 (O_553,N_4770,N_4758);
and UO_554 (O_554,N_4546,N_4857);
and UO_555 (O_555,N_4652,N_4872);
and UO_556 (O_556,N_4667,N_4623);
or UO_557 (O_557,N_4676,N_4582);
and UO_558 (O_558,N_4784,N_4664);
xor UO_559 (O_559,N_4906,N_4759);
and UO_560 (O_560,N_4887,N_4791);
and UO_561 (O_561,N_4812,N_4687);
and UO_562 (O_562,N_4592,N_4759);
nor UO_563 (O_563,N_4753,N_4793);
nand UO_564 (O_564,N_4651,N_4551);
nor UO_565 (O_565,N_4937,N_4888);
nor UO_566 (O_566,N_4627,N_4816);
nor UO_567 (O_567,N_4886,N_4570);
nand UO_568 (O_568,N_4929,N_4649);
nor UO_569 (O_569,N_4968,N_4546);
xnor UO_570 (O_570,N_4558,N_4759);
nand UO_571 (O_571,N_4703,N_4601);
and UO_572 (O_572,N_4901,N_4745);
or UO_573 (O_573,N_4650,N_4820);
nor UO_574 (O_574,N_4923,N_4619);
or UO_575 (O_575,N_4502,N_4511);
or UO_576 (O_576,N_4841,N_4757);
or UO_577 (O_577,N_4751,N_4854);
nand UO_578 (O_578,N_4695,N_4595);
nor UO_579 (O_579,N_4800,N_4632);
or UO_580 (O_580,N_4980,N_4958);
nor UO_581 (O_581,N_4578,N_4917);
and UO_582 (O_582,N_4730,N_4703);
nor UO_583 (O_583,N_4504,N_4623);
or UO_584 (O_584,N_4861,N_4922);
nor UO_585 (O_585,N_4746,N_4858);
and UO_586 (O_586,N_4616,N_4641);
and UO_587 (O_587,N_4710,N_4865);
or UO_588 (O_588,N_4638,N_4940);
and UO_589 (O_589,N_4689,N_4632);
nor UO_590 (O_590,N_4667,N_4961);
nor UO_591 (O_591,N_4911,N_4603);
and UO_592 (O_592,N_4818,N_4598);
and UO_593 (O_593,N_4764,N_4955);
nand UO_594 (O_594,N_4806,N_4812);
or UO_595 (O_595,N_4836,N_4540);
or UO_596 (O_596,N_4955,N_4815);
xnor UO_597 (O_597,N_4548,N_4721);
nor UO_598 (O_598,N_4918,N_4553);
and UO_599 (O_599,N_4822,N_4778);
or UO_600 (O_600,N_4617,N_4625);
nor UO_601 (O_601,N_4672,N_4776);
nor UO_602 (O_602,N_4502,N_4509);
and UO_603 (O_603,N_4534,N_4877);
or UO_604 (O_604,N_4979,N_4851);
and UO_605 (O_605,N_4982,N_4913);
nor UO_606 (O_606,N_4677,N_4628);
nand UO_607 (O_607,N_4776,N_4757);
nand UO_608 (O_608,N_4896,N_4961);
or UO_609 (O_609,N_4926,N_4643);
or UO_610 (O_610,N_4570,N_4954);
nor UO_611 (O_611,N_4604,N_4723);
and UO_612 (O_612,N_4999,N_4745);
and UO_613 (O_613,N_4853,N_4585);
nor UO_614 (O_614,N_4586,N_4613);
nor UO_615 (O_615,N_4877,N_4970);
and UO_616 (O_616,N_4909,N_4640);
nor UO_617 (O_617,N_4883,N_4983);
or UO_618 (O_618,N_4952,N_4949);
nand UO_619 (O_619,N_4594,N_4889);
nand UO_620 (O_620,N_4857,N_4841);
and UO_621 (O_621,N_4968,N_4930);
or UO_622 (O_622,N_4895,N_4754);
nand UO_623 (O_623,N_4650,N_4675);
nand UO_624 (O_624,N_4757,N_4606);
and UO_625 (O_625,N_4886,N_4775);
nand UO_626 (O_626,N_4717,N_4753);
nor UO_627 (O_627,N_4701,N_4574);
or UO_628 (O_628,N_4636,N_4925);
or UO_629 (O_629,N_4886,N_4629);
nand UO_630 (O_630,N_4731,N_4604);
nor UO_631 (O_631,N_4525,N_4600);
nand UO_632 (O_632,N_4890,N_4946);
nand UO_633 (O_633,N_4656,N_4985);
and UO_634 (O_634,N_4797,N_4794);
or UO_635 (O_635,N_4669,N_4690);
or UO_636 (O_636,N_4802,N_4644);
nand UO_637 (O_637,N_4846,N_4548);
or UO_638 (O_638,N_4708,N_4505);
nor UO_639 (O_639,N_4738,N_4538);
nand UO_640 (O_640,N_4587,N_4954);
nor UO_641 (O_641,N_4767,N_4970);
and UO_642 (O_642,N_4522,N_4516);
nor UO_643 (O_643,N_4500,N_4864);
or UO_644 (O_644,N_4509,N_4713);
nor UO_645 (O_645,N_4876,N_4790);
or UO_646 (O_646,N_4899,N_4917);
nand UO_647 (O_647,N_4847,N_4996);
and UO_648 (O_648,N_4516,N_4848);
and UO_649 (O_649,N_4909,N_4957);
and UO_650 (O_650,N_4736,N_4658);
nand UO_651 (O_651,N_4654,N_4631);
nor UO_652 (O_652,N_4945,N_4807);
and UO_653 (O_653,N_4770,N_4573);
and UO_654 (O_654,N_4691,N_4763);
and UO_655 (O_655,N_4796,N_4715);
and UO_656 (O_656,N_4965,N_4910);
nand UO_657 (O_657,N_4857,N_4988);
and UO_658 (O_658,N_4985,N_4801);
and UO_659 (O_659,N_4925,N_4689);
or UO_660 (O_660,N_4521,N_4775);
nand UO_661 (O_661,N_4740,N_4862);
and UO_662 (O_662,N_4947,N_4612);
or UO_663 (O_663,N_4535,N_4822);
and UO_664 (O_664,N_4958,N_4788);
nand UO_665 (O_665,N_4584,N_4560);
and UO_666 (O_666,N_4549,N_4718);
nand UO_667 (O_667,N_4731,N_4703);
nand UO_668 (O_668,N_4992,N_4960);
or UO_669 (O_669,N_4810,N_4811);
nor UO_670 (O_670,N_4642,N_4923);
or UO_671 (O_671,N_4875,N_4669);
or UO_672 (O_672,N_4536,N_4920);
and UO_673 (O_673,N_4562,N_4635);
nor UO_674 (O_674,N_4886,N_4566);
nor UO_675 (O_675,N_4793,N_4669);
nand UO_676 (O_676,N_4607,N_4674);
nor UO_677 (O_677,N_4876,N_4704);
and UO_678 (O_678,N_4715,N_4504);
nand UO_679 (O_679,N_4541,N_4893);
nor UO_680 (O_680,N_4804,N_4511);
nor UO_681 (O_681,N_4523,N_4626);
nand UO_682 (O_682,N_4966,N_4605);
nor UO_683 (O_683,N_4786,N_4564);
nor UO_684 (O_684,N_4816,N_4866);
nand UO_685 (O_685,N_4939,N_4760);
nor UO_686 (O_686,N_4852,N_4574);
nand UO_687 (O_687,N_4631,N_4553);
nand UO_688 (O_688,N_4753,N_4952);
nor UO_689 (O_689,N_4567,N_4858);
or UO_690 (O_690,N_4637,N_4988);
or UO_691 (O_691,N_4774,N_4854);
or UO_692 (O_692,N_4837,N_4619);
nor UO_693 (O_693,N_4599,N_4744);
and UO_694 (O_694,N_4719,N_4853);
nand UO_695 (O_695,N_4664,N_4795);
and UO_696 (O_696,N_4774,N_4824);
nand UO_697 (O_697,N_4824,N_4942);
nand UO_698 (O_698,N_4628,N_4949);
and UO_699 (O_699,N_4716,N_4802);
nor UO_700 (O_700,N_4968,N_4825);
nor UO_701 (O_701,N_4936,N_4749);
nor UO_702 (O_702,N_4992,N_4564);
or UO_703 (O_703,N_4850,N_4613);
and UO_704 (O_704,N_4986,N_4525);
nand UO_705 (O_705,N_4714,N_4530);
and UO_706 (O_706,N_4827,N_4738);
nor UO_707 (O_707,N_4506,N_4829);
nand UO_708 (O_708,N_4644,N_4638);
nand UO_709 (O_709,N_4828,N_4607);
or UO_710 (O_710,N_4570,N_4537);
and UO_711 (O_711,N_4953,N_4737);
and UO_712 (O_712,N_4633,N_4641);
and UO_713 (O_713,N_4855,N_4940);
xnor UO_714 (O_714,N_4845,N_4733);
nor UO_715 (O_715,N_4858,N_4718);
nor UO_716 (O_716,N_4907,N_4835);
or UO_717 (O_717,N_4579,N_4978);
or UO_718 (O_718,N_4643,N_4558);
or UO_719 (O_719,N_4824,N_4528);
nor UO_720 (O_720,N_4590,N_4519);
nand UO_721 (O_721,N_4724,N_4802);
or UO_722 (O_722,N_4825,N_4866);
nor UO_723 (O_723,N_4571,N_4867);
nand UO_724 (O_724,N_4724,N_4618);
or UO_725 (O_725,N_4760,N_4839);
or UO_726 (O_726,N_4555,N_4844);
or UO_727 (O_727,N_4640,N_4953);
nor UO_728 (O_728,N_4628,N_4914);
and UO_729 (O_729,N_4856,N_4651);
nor UO_730 (O_730,N_4709,N_4842);
nand UO_731 (O_731,N_4798,N_4650);
or UO_732 (O_732,N_4965,N_4843);
or UO_733 (O_733,N_4714,N_4704);
and UO_734 (O_734,N_4817,N_4756);
or UO_735 (O_735,N_4892,N_4696);
nand UO_736 (O_736,N_4911,N_4696);
nand UO_737 (O_737,N_4900,N_4647);
nand UO_738 (O_738,N_4600,N_4804);
nand UO_739 (O_739,N_4708,N_4754);
and UO_740 (O_740,N_4658,N_4867);
or UO_741 (O_741,N_4847,N_4792);
and UO_742 (O_742,N_4897,N_4535);
nand UO_743 (O_743,N_4997,N_4701);
or UO_744 (O_744,N_4639,N_4555);
nor UO_745 (O_745,N_4748,N_4881);
or UO_746 (O_746,N_4828,N_4918);
nand UO_747 (O_747,N_4962,N_4968);
and UO_748 (O_748,N_4856,N_4765);
nor UO_749 (O_749,N_4810,N_4645);
and UO_750 (O_750,N_4525,N_4653);
and UO_751 (O_751,N_4707,N_4743);
and UO_752 (O_752,N_4719,N_4977);
nor UO_753 (O_753,N_4872,N_4563);
nand UO_754 (O_754,N_4506,N_4732);
and UO_755 (O_755,N_4909,N_4910);
and UO_756 (O_756,N_4981,N_4803);
and UO_757 (O_757,N_4609,N_4685);
nand UO_758 (O_758,N_4925,N_4928);
nand UO_759 (O_759,N_4924,N_4887);
nand UO_760 (O_760,N_4955,N_4735);
nor UO_761 (O_761,N_4773,N_4722);
or UO_762 (O_762,N_4977,N_4847);
nand UO_763 (O_763,N_4951,N_4629);
and UO_764 (O_764,N_4694,N_4879);
or UO_765 (O_765,N_4854,N_4717);
nor UO_766 (O_766,N_4783,N_4941);
and UO_767 (O_767,N_4805,N_4776);
and UO_768 (O_768,N_4816,N_4847);
nand UO_769 (O_769,N_4674,N_4779);
and UO_770 (O_770,N_4506,N_4662);
and UO_771 (O_771,N_4557,N_4592);
nand UO_772 (O_772,N_4687,N_4523);
or UO_773 (O_773,N_4673,N_4738);
nor UO_774 (O_774,N_4946,N_4545);
nor UO_775 (O_775,N_4696,N_4868);
or UO_776 (O_776,N_4950,N_4644);
nor UO_777 (O_777,N_4633,N_4797);
nand UO_778 (O_778,N_4839,N_4996);
nor UO_779 (O_779,N_4737,N_4593);
and UO_780 (O_780,N_4702,N_4502);
and UO_781 (O_781,N_4992,N_4618);
or UO_782 (O_782,N_4779,N_4584);
or UO_783 (O_783,N_4523,N_4842);
and UO_784 (O_784,N_4866,N_4817);
or UO_785 (O_785,N_4524,N_4739);
or UO_786 (O_786,N_4978,N_4544);
or UO_787 (O_787,N_4545,N_4633);
and UO_788 (O_788,N_4541,N_4866);
and UO_789 (O_789,N_4798,N_4608);
nand UO_790 (O_790,N_4701,N_4794);
nand UO_791 (O_791,N_4824,N_4737);
nor UO_792 (O_792,N_4854,N_4541);
nand UO_793 (O_793,N_4908,N_4767);
or UO_794 (O_794,N_4595,N_4932);
xor UO_795 (O_795,N_4987,N_4636);
nor UO_796 (O_796,N_4830,N_4677);
and UO_797 (O_797,N_4880,N_4696);
nand UO_798 (O_798,N_4631,N_4813);
nor UO_799 (O_799,N_4672,N_4935);
nand UO_800 (O_800,N_4992,N_4910);
and UO_801 (O_801,N_4865,N_4824);
nand UO_802 (O_802,N_4825,N_4975);
or UO_803 (O_803,N_4959,N_4736);
and UO_804 (O_804,N_4728,N_4676);
and UO_805 (O_805,N_4660,N_4505);
and UO_806 (O_806,N_4837,N_4820);
and UO_807 (O_807,N_4604,N_4634);
nand UO_808 (O_808,N_4601,N_4921);
nor UO_809 (O_809,N_4580,N_4990);
and UO_810 (O_810,N_4886,N_4659);
or UO_811 (O_811,N_4574,N_4588);
nor UO_812 (O_812,N_4788,N_4678);
or UO_813 (O_813,N_4834,N_4525);
and UO_814 (O_814,N_4585,N_4682);
nor UO_815 (O_815,N_4857,N_4550);
and UO_816 (O_816,N_4722,N_4988);
and UO_817 (O_817,N_4832,N_4862);
or UO_818 (O_818,N_4576,N_4905);
or UO_819 (O_819,N_4591,N_4946);
and UO_820 (O_820,N_4969,N_4529);
or UO_821 (O_821,N_4785,N_4651);
or UO_822 (O_822,N_4910,N_4969);
and UO_823 (O_823,N_4560,N_4668);
xor UO_824 (O_824,N_4697,N_4938);
nand UO_825 (O_825,N_4574,N_4866);
nor UO_826 (O_826,N_4714,N_4735);
or UO_827 (O_827,N_4666,N_4862);
and UO_828 (O_828,N_4769,N_4981);
or UO_829 (O_829,N_4922,N_4990);
and UO_830 (O_830,N_4713,N_4651);
or UO_831 (O_831,N_4895,N_4594);
or UO_832 (O_832,N_4807,N_4970);
and UO_833 (O_833,N_4715,N_4999);
or UO_834 (O_834,N_4609,N_4569);
or UO_835 (O_835,N_4655,N_4519);
and UO_836 (O_836,N_4981,N_4520);
nand UO_837 (O_837,N_4613,N_4880);
nand UO_838 (O_838,N_4770,N_4874);
and UO_839 (O_839,N_4679,N_4643);
and UO_840 (O_840,N_4924,N_4991);
nor UO_841 (O_841,N_4913,N_4690);
and UO_842 (O_842,N_4993,N_4994);
and UO_843 (O_843,N_4961,N_4867);
nor UO_844 (O_844,N_4517,N_4596);
nand UO_845 (O_845,N_4983,N_4902);
or UO_846 (O_846,N_4951,N_4592);
xnor UO_847 (O_847,N_4736,N_4817);
or UO_848 (O_848,N_4530,N_4928);
or UO_849 (O_849,N_4722,N_4804);
nor UO_850 (O_850,N_4964,N_4627);
nand UO_851 (O_851,N_4554,N_4612);
nor UO_852 (O_852,N_4978,N_4587);
nand UO_853 (O_853,N_4611,N_4824);
and UO_854 (O_854,N_4907,N_4708);
nand UO_855 (O_855,N_4890,N_4705);
and UO_856 (O_856,N_4505,N_4859);
nand UO_857 (O_857,N_4595,N_4709);
nor UO_858 (O_858,N_4820,N_4781);
and UO_859 (O_859,N_4518,N_4670);
nor UO_860 (O_860,N_4537,N_4604);
and UO_861 (O_861,N_4507,N_4586);
or UO_862 (O_862,N_4909,N_4890);
nor UO_863 (O_863,N_4935,N_4633);
and UO_864 (O_864,N_4901,N_4741);
and UO_865 (O_865,N_4659,N_4537);
nand UO_866 (O_866,N_4690,N_4937);
or UO_867 (O_867,N_4863,N_4899);
and UO_868 (O_868,N_4586,N_4601);
nor UO_869 (O_869,N_4968,N_4654);
and UO_870 (O_870,N_4623,N_4723);
and UO_871 (O_871,N_4860,N_4579);
and UO_872 (O_872,N_4523,N_4525);
and UO_873 (O_873,N_4969,N_4516);
and UO_874 (O_874,N_4947,N_4846);
nor UO_875 (O_875,N_4767,N_4740);
or UO_876 (O_876,N_4961,N_4710);
and UO_877 (O_877,N_4996,N_4897);
or UO_878 (O_878,N_4619,N_4604);
nor UO_879 (O_879,N_4824,N_4567);
nor UO_880 (O_880,N_4633,N_4976);
and UO_881 (O_881,N_4970,N_4863);
or UO_882 (O_882,N_4714,N_4619);
and UO_883 (O_883,N_4591,N_4948);
nand UO_884 (O_884,N_4907,N_4988);
nand UO_885 (O_885,N_4544,N_4822);
nor UO_886 (O_886,N_4811,N_4532);
or UO_887 (O_887,N_4975,N_4816);
nand UO_888 (O_888,N_4832,N_4889);
and UO_889 (O_889,N_4917,N_4600);
or UO_890 (O_890,N_4516,N_4656);
nand UO_891 (O_891,N_4808,N_4706);
or UO_892 (O_892,N_4598,N_4613);
and UO_893 (O_893,N_4516,N_4696);
and UO_894 (O_894,N_4532,N_4518);
and UO_895 (O_895,N_4883,N_4674);
or UO_896 (O_896,N_4702,N_4903);
or UO_897 (O_897,N_4893,N_4544);
nand UO_898 (O_898,N_4717,N_4950);
and UO_899 (O_899,N_4550,N_4780);
nor UO_900 (O_900,N_4841,N_4719);
nand UO_901 (O_901,N_4755,N_4981);
and UO_902 (O_902,N_4564,N_4780);
and UO_903 (O_903,N_4761,N_4772);
and UO_904 (O_904,N_4853,N_4848);
and UO_905 (O_905,N_4526,N_4908);
xnor UO_906 (O_906,N_4680,N_4849);
nor UO_907 (O_907,N_4891,N_4612);
nand UO_908 (O_908,N_4520,N_4873);
nor UO_909 (O_909,N_4719,N_4509);
or UO_910 (O_910,N_4948,N_4579);
nor UO_911 (O_911,N_4658,N_4769);
nor UO_912 (O_912,N_4715,N_4823);
nand UO_913 (O_913,N_4820,N_4660);
nor UO_914 (O_914,N_4556,N_4579);
nor UO_915 (O_915,N_4982,N_4670);
and UO_916 (O_916,N_4855,N_4617);
nand UO_917 (O_917,N_4894,N_4631);
and UO_918 (O_918,N_4562,N_4971);
nand UO_919 (O_919,N_4621,N_4902);
nor UO_920 (O_920,N_4647,N_4984);
nand UO_921 (O_921,N_4776,N_4685);
nor UO_922 (O_922,N_4681,N_4724);
nor UO_923 (O_923,N_4885,N_4691);
or UO_924 (O_924,N_4537,N_4993);
nand UO_925 (O_925,N_4597,N_4555);
xnor UO_926 (O_926,N_4978,N_4535);
or UO_927 (O_927,N_4711,N_4808);
nor UO_928 (O_928,N_4637,N_4968);
or UO_929 (O_929,N_4627,N_4874);
nand UO_930 (O_930,N_4587,N_4620);
or UO_931 (O_931,N_4962,N_4916);
nor UO_932 (O_932,N_4632,N_4928);
nand UO_933 (O_933,N_4690,N_4772);
xnor UO_934 (O_934,N_4781,N_4878);
or UO_935 (O_935,N_4994,N_4586);
and UO_936 (O_936,N_4632,N_4634);
nand UO_937 (O_937,N_4595,N_4794);
and UO_938 (O_938,N_4978,N_4816);
nor UO_939 (O_939,N_4961,N_4573);
nor UO_940 (O_940,N_4895,N_4913);
and UO_941 (O_941,N_4696,N_4735);
nand UO_942 (O_942,N_4609,N_4605);
or UO_943 (O_943,N_4959,N_4760);
or UO_944 (O_944,N_4643,N_4849);
nand UO_945 (O_945,N_4699,N_4933);
nor UO_946 (O_946,N_4888,N_4797);
nor UO_947 (O_947,N_4669,N_4859);
nand UO_948 (O_948,N_4612,N_4509);
or UO_949 (O_949,N_4960,N_4845);
or UO_950 (O_950,N_4769,N_4652);
or UO_951 (O_951,N_4726,N_4725);
or UO_952 (O_952,N_4842,N_4672);
and UO_953 (O_953,N_4933,N_4549);
or UO_954 (O_954,N_4607,N_4848);
nand UO_955 (O_955,N_4840,N_4556);
or UO_956 (O_956,N_4623,N_4960);
nor UO_957 (O_957,N_4760,N_4600);
nand UO_958 (O_958,N_4522,N_4908);
or UO_959 (O_959,N_4988,N_4514);
nor UO_960 (O_960,N_4973,N_4905);
and UO_961 (O_961,N_4994,N_4745);
nor UO_962 (O_962,N_4941,N_4578);
and UO_963 (O_963,N_4584,N_4763);
nand UO_964 (O_964,N_4820,N_4605);
and UO_965 (O_965,N_4505,N_4956);
nand UO_966 (O_966,N_4833,N_4681);
and UO_967 (O_967,N_4801,N_4906);
and UO_968 (O_968,N_4887,N_4735);
or UO_969 (O_969,N_4553,N_4847);
nand UO_970 (O_970,N_4913,N_4890);
nand UO_971 (O_971,N_4633,N_4827);
or UO_972 (O_972,N_4755,N_4512);
or UO_973 (O_973,N_4695,N_4995);
or UO_974 (O_974,N_4961,N_4663);
or UO_975 (O_975,N_4770,N_4968);
nand UO_976 (O_976,N_4990,N_4666);
xnor UO_977 (O_977,N_4689,N_4542);
nand UO_978 (O_978,N_4714,N_4847);
nand UO_979 (O_979,N_4621,N_4901);
xnor UO_980 (O_980,N_4850,N_4631);
nand UO_981 (O_981,N_4830,N_4844);
or UO_982 (O_982,N_4609,N_4752);
nand UO_983 (O_983,N_4735,N_4573);
nand UO_984 (O_984,N_4978,N_4963);
nand UO_985 (O_985,N_4565,N_4752);
or UO_986 (O_986,N_4583,N_4716);
or UO_987 (O_987,N_4503,N_4755);
nand UO_988 (O_988,N_4733,N_4860);
nor UO_989 (O_989,N_4625,N_4521);
and UO_990 (O_990,N_4695,N_4981);
or UO_991 (O_991,N_4699,N_4986);
nand UO_992 (O_992,N_4647,N_4997);
nor UO_993 (O_993,N_4608,N_4727);
nand UO_994 (O_994,N_4707,N_4872);
and UO_995 (O_995,N_4836,N_4625);
nor UO_996 (O_996,N_4807,N_4628);
nor UO_997 (O_997,N_4701,N_4815);
nand UO_998 (O_998,N_4721,N_4798);
nor UO_999 (O_999,N_4869,N_4728);
endmodule