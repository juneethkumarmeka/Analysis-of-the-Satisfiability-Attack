module basic_3000_30000_3500_6_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_1103,In_302);
xor U1 (N_1,In_1130,In_88);
xnor U2 (N_2,In_1305,In_674);
nand U3 (N_3,In_1864,In_1137);
nand U4 (N_4,In_233,In_2677);
xor U5 (N_5,In_1334,In_1272);
xor U6 (N_6,In_1476,In_1671);
xnor U7 (N_7,In_1067,In_700);
nand U8 (N_8,In_2949,In_643);
and U9 (N_9,In_2828,In_703);
or U10 (N_10,In_2843,In_1095);
xor U11 (N_11,In_765,In_1405);
and U12 (N_12,In_1695,In_1750);
nor U13 (N_13,In_1174,In_437);
and U14 (N_14,In_2608,In_203);
or U15 (N_15,In_2972,In_460);
nor U16 (N_16,In_319,In_1599);
nand U17 (N_17,In_656,In_2381);
or U18 (N_18,In_1669,In_1071);
nor U19 (N_19,In_267,In_1717);
xnor U20 (N_20,In_1815,In_673);
nand U21 (N_21,In_1893,In_1374);
or U22 (N_22,In_2286,In_2890);
and U23 (N_23,In_124,In_2570);
xor U24 (N_24,In_2299,In_2601);
xnor U25 (N_25,In_1625,In_954);
xor U26 (N_26,In_178,In_1868);
nor U27 (N_27,In_10,In_2503);
nand U28 (N_28,In_1425,In_2938);
or U29 (N_29,In_556,In_2384);
nand U30 (N_30,In_62,In_2144);
nand U31 (N_31,In_611,In_2595);
xor U32 (N_32,In_2597,In_2529);
nand U33 (N_33,In_2180,In_895);
nand U34 (N_34,In_2347,In_1110);
nand U35 (N_35,In_839,In_518);
or U36 (N_36,In_8,In_352);
and U37 (N_37,In_2399,In_2365);
nor U38 (N_38,In_2305,In_446);
nor U39 (N_39,In_2551,In_949);
nand U40 (N_40,In_472,In_1404);
nor U41 (N_41,In_2770,In_2190);
nand U42 (N_42,In_2835,In_2408);
xor U43 (N_43,In_392,In_741);
xnor U44 (N_44,In_2525,In_1445);
xnor U45 (N_45,In_1696,In_59);
or U46 (N_46,In_917,In_2829);
xor U47 (N_47,In_2308,In_763);
nand U48 (N_48,In_279,In_347);
nor U49 (N_49,In_862,In_1951);
or U50 (N_50,In_2557,In_465);
or U51 (N_51,In_1031,In_2338);
xnor U52 (N_52,In_2398,In_589);
nand U53 (N_53,In_1099,In_2075);
nand U54 (N_54,In_2039,In_2096);
xor U55 (N_55,In_2255,In_1654);
or U56 (N_56,In_2052,In_1954);
nor U57 (N_57,In_2623,In_141);
nor U58 (N_58,In_2173,In_2790);
nand U59 (N_59,In_1459,In_381);
or U60 (N_60,In_1899,In_550);
nor U61 (N_61,In_1813,In_2030);
nor U62 (N_62,In_2893,In_1752);
and U63 (N_63,In_1348,In_992);
nand U64 (N_64,In_308,In_1724);
nand U65 (N_65,In_2647,In_2650);
xor U66 (N_66,In_2705,In_2625);
xor U67 (N_67,In_2146,In_1441);
nand U68 (N_68,In_822,In_1610);
nor U69 (N_69,In_2488,In_265);
xnor U70 (N_70,In_1368,In_587);
xor U71 (N_71,In_2068,In_2813);
nor U72 (N_72,In_600,In_2497);
nor U73 (N_73,In_94,In_2020);
xnor U74 (N_74,In_758,In_2065);
nor U75 (N_75,In_2543,In_582);
and U76 (N_76,In_543,In_1213);
nor U77 (N_77,In_1340,In_2581);
and U78 (N_78,In_1367,In_2248);
nand U79 (N_79,In_1656,In_1915);
or U80 (N_80,In_2285,In_2249);
and U81 (N_81,In_49,In_2087);
or U82 (N_82,In_1351,In_216);
nand U83 (N_83,In_775,In_1366);
or U84 (N_84,In_1082,In_2711);
xnor U85 (N_85,In_2322,In_2434);
nand U86 (N_86,In_492,In_2694);
nand U87 (N_87,In_1331,In_2059);
nand U88 (N_88,In_1207,In_1420);
nand U89 (N_89,In_853,In_1451);
or U90 (N_90,In_383,In_1276);
nor U91 (N_91,In_752,In_2196);
xnor U92 (N_92,In_2135,In_2638);
nor U93 (N_93,In_647,In_940);
and U94 (N_94,In_2022,In_1081);
and U95 (N_95,In_2532,In_1212);
or U96 (N_96,In_1831,In_2914);
or U97 (N_97,In_274,In_1215);
nor U98 (N_98,In_266,In_2303);
nand U99 (N_99,In_264,In_2066);
xnor U100 (N_100,In_478,In_2763);
nand U101 (N_101,In_1784,In_1021);
nand U102 (N_102,In_715,In_619);
nor U103 (N_103,In_1707,In_1527);
or U104 (N_104,In_2147,In_400);
or U105 (N_105,In_2811,In_1265);
and U106 (N_106,In_1162,In_2117);
and U107 (N_107,In_2072,In_299);
nor U108 (N_108,In_711,In_2684);
and U109 (N_109,In_2743,In_2159);
or U110 (N_110,In_1824,In_1539);
or U111 (N_111,In_67,In_1297);
or U112 (N_112,In_2375,In_2453);
or U113 (N_113,In_1995,In_1820);
or U114 (N_114,In_1538,In_2069);
xnor U115 (N_115,In_125,In_2254);
xor U116 (N_116,In_236,In_237);
or U117 (N_117,In_2247,In_37);
and U118 (N_118,In_2427,In_982);
nor U119 (N_119,In_1719,In_666);
nor U120 (N_120,In_2028,In_2928);
or U121 (N_121,In_2917,In_2686);
and U122 (N_122,In_1238,In_1950);
and U123 (N_123,In_527,In_1470);
nor U124 (N_124,In_2726,In_1833);
nor U125 (N_125,In_1809,In_2221);
xnor U126 (N_126,In_2079,In_507);
nor U127 (N_127,In_2007,In_20);
and U128 (N_128,In_635,In_486);
and U129 (N_129,In_1423,In_2413);
or U130 (N_130,In_2493,In_2432);
and U131 (N_131,In_730,In_2518);
and U132 (N_132,In_753,In_959);
nand U133 (N_133,In_45,In_2231);
nor U134 (N_134,In_658,In_257);
nand U135 (N_135,In_130,In_1579);
nand U136 (N_136,In_1972,In_1490);
or U137 (N_137,In_1729,In_719);
or U138 (N_138,In_1085,In_1027);
nor U139 (N_139,In_935,In_2903);
nor U140 (N_140,In_2293,In_2386);
xnor U141 (N_141,In_733,In_1450);
nor U142 (N_142,In_2900,In_2553);
nor U143 (N_143,In_1063,In_732);
or U144 (N_144,In_2202,In_334);
or U145 (N_145,In_2415,In_2867);
xor U146 (N_146,In_2219,In_2420);
nand U147 (N_147,In_1391,In_2130);
and U148 (N_148,In_2354,In_688);
nand U149 (N_149,In_293,In_761);
xor U150 (N_150,In_642,In_2586);
or U151 (N_151,In_1121,In_1894);
or U152 (N_152,In_1512,In_2986);
nor U153 (N_153,In_2626,In_2641);
xor U154 (N_154,In_1294,In_490);
and U155 (N_155,In_2954,In_814);
xnor U156 (N_156,In_1416,In_512);
xnor U157 (N_157,In_2545,In_2667);
nand U158 (N_158,In_1034,In_2590);
nand U159 (N_159,In_1756,In_1901);
nand U160 (N_160,In_2778,In_2437);
nor U161 (N_161,In_450,In_1100);
or U162 (N_162,In_2664,In_411);
nand U163 (N_163,In_2931,In_2081);
xnor U164 (N_164,In_2137,In_1258);
or U165 (N_165,In_2213,In_1937);
and U166 (N_166,In_397,In_2418);
nor U167 (N_167,In_1264,In_425);
nor U168 (N_168,In_426,In_180);
or U169 (N_169,In_2780,In_629);
xor U170 (N_170,In_2655,In_722);
and U171 (N_171,In_154,In_2609);
and U172 (N_172,In_342,In_2592);
nor U173 (N_173,In_2878,In_1716);
and U174 (N_174,In_821,In_1353);
xnor U175 (N_175,In_2017,In_813);
or U176 (N_176,In_2212,In_2192);
or U177 (N_177,In_2058,In_706);
xnor U178 (N_178,In_239,In_942);
nor U179 (N_179,In_598,In_1038);
nand U180 (N_180,In_1902,In_1505);
and U181 (N_181,In_2492,In_2730);
nor U182 (N_182,In_655,In_1545);
or U183 (N_183,In_2268,In_213);
or U184 (N_184,In_312,In_1898);
and U185 (N_185,In_1659,In_468);
or U186 (N_186,In_2636,In_2681);
nand U187 (N_187,In_1112,In_2319);
nor U188 (N_188,In_315,In_2663);
nand U189 (N_189,In_607,In_454);
nand U190 (N_190,In_2669,In_1332);
nor U191 (N_191,In_859,In_770);
and U192 (N_192,In_2339,In_2490);
and U193 (N_193,In_354,In_2163);
nand U194 (N_194,In_2732,In_146);
and U195 (N_195,In_691,In_287);
xor U196 (N_196,In_845,In_1515);
nand U197 (N_197,In_1997,In_1280);
or U198 (N_198,In_742,In_2206);
or U199 (N_199,In_2011,In_2891);
nand U200 (N_200,In_885,In_1436);
nand U201 (N_201,In_890,In_1380);
nor U202 (N_202,In_2548,In_2393);
or U203 (N_203,In_2719,In_1727);
nor U204 (N_204,In_491,In_2980);
and U205 (N_205,In_2531,In_905);
and U206 (N_206,In_1573,In_1770);
nor U207 (N_207,In_1637,In_2818);
xor U208 (N_208,In_269,In_441);
nor U209 (N_209,In_429,In_1442);
and U210 (N_210,In_1775,In_82);
nor U211 (N_211,In_760,In_2031);
or U212 (N_212,In_2985,In_2652);
nor U213 (N_213,In_2907,In_173);
nand U214 (N_214,In_2912,In_965);
xor U215 (N_215,In_2430,In_1589);
nand U216 (N_216,In_2544,In_440);
or U217 (N_217,In_1127,In_2654);
or U218 (N_218,In_38,In_762);
nor U219 (N_219,In_345,In_477);
nor U220 (N_220,In_1285,In_224);
xnor U221 (N_221,In_1065,In_1411);
nand U222 (N_222,In_1010,In_150);
and U223 (N_223,In_1473,In_1392);
xor U224 (N_224,In_1347,In_2982);
xor U225 (N_225,In_1266,In_1487);
xnor U226 (N_226,In_2808,In_1356);
nand U227 (N_227,In_2474,In_1938);
or U228 (N_228,In_604,In_1106);
nand U229 (N_229,In_744,In_1399);
or U230 (N_230,In_1867,In_1861);
nor U231 (N_231,In_1734,In_2209);
or U232 (N_232,In_2389,In_1157);
xor U233 (N_233,In_71,In_1428);
and U234 (N_234,In_689,In_579);
or U235 (N_235,In_152,In_1923);
nor U236 (N_236,In_128,In_2043);
or U237 (N_237,In_1313,In_209);
and U238 (N_238,In_356,In_1378);
or U239 (N_239,In_1605,In_2807);
and U240 (N_240,In_2046,In_1224);
nor U241 (N_241,In_1042,In_1237);
nand U242 (N_242,In_404,In_2649);
or U243 (N_243,In_801,In_363);
and U244 (N_244,In_520,In_2123);
nand U245 (N_245,In_242,In_2617);
nor U246 (N_246,In_1373,In_2336);
and U247 (N_247,In_2707,In_2584);
nor U248 (N_248,In_538,In_2416);
xor U249 (N_249,In_1216,In_676);
nand U250 (N_250,In_2971,In_1714);
nand U251 (N_251,In_375,In_1419);
and U252 (N_252,In_1241,In_780);
nor U253 (N_253,In_1461,In_1591);
and U254 (N_254,In_1713,In_2542);
nand U255 (N_255,In_338,In_1381);
nor U256 (N_256,In_2361,In_1536);
and U257 (N_257,In_1751,In_1803);
nor U258 (N_258,In_561,In_2576);
and U259 (N_259,In_792,In_155);
nand U260 (N_260,In_876,In_2675);
nand U261 (N_261,In_1726,In_1246);
xor U262 (N_262,In_899,In_2312);
xor U263 (N_263,In_68,In_2100);
or U264 (N_264,In_1846,In_2252);
xnor U265 (N_265,In_2331,In_2197);
and U266 (N_266,In_416,In_2603);
nor U267 (N_267,In_1664,In_2676);
nor U268 (N_268,In_2325,In_2659);
xor U269 (N_269,In_84,In_2124);
or U270 (N_270,In_2793,In_2051);
and U271 (N_271,In_1288,In_2155);
nand U272 (N_272,In_1931,In_1608);
nand U273 (N_273,In_1706,In_716);
nand U274 (N_274,In_2118,In_2988);
xor U275 (N_275,In_808,In_2296);
nor U276 (N_276,In_1830,In_951);
nor U277 (N_277,In_843,In_2919);
or U278 (N_278,In_101,In_880);
and U279 (N_279,In_343,In_421);
or U280 (N_280,In_869,In_1074);
and U281 (N_281,In_2307,In_1330);
or U282 (N_282,In_927,In_2379);
xor U283 (N_283,In_1084,In_728);
nand U284 (N_284,In_2761,In_2396);
and U285 (N_285,In_893,In_1444);
xnor U286 (N_286,In_1218,In_1692);
or U287 (N_287,In_2332,In_612);
or U288 (N_288,In_2152,In_2480);
nor U289 (N_289,In_1778,In_2442);
or U290 (N_290,In_2195,In_424);
or U291 (N_291,In_262,In_1182);
xor U292 (N_292,In_234,In_361);
nor U293 (N_293,In_2512,In_2624);
or U294 (N_294,In_2351,In_672);
xnor U295 (N_295,In_721,In_2070);
and U296 (N_296,In_2318,In_235);
xor U297 (N_297,In_480,In_73);
and U298 (N_298,In_1032,In_794);
and U299 (N_299,In_840,In_2089);
nand U300 (N_300,In_273,In_535);
nor U301 (N_301,In_1779,In_2539);
nand U302 (N_302,In_1811,In_566);
nor U303 (N_303,In_1007,In_495);
xnor U304 (N_304,In_963,In_1501);
nand U305 (N_305,In_637,In_1994);
and U306 (N_306,In_2400,In_1583);
and U307 (N_307,In_2585,In_1971);
nand U308 (N_308,In_2611,In_922);
xor U309 (N_309,In_1616,In_986);
or U310 (N_310,In_405,In_777);
xnor U311 (N_311,In_9,In_1662);
and U312 (N_312,In_1295,In_1959);
and U313 (N_313,In_1427,In_2614);
nor U314 (N_314,In_1666,In_1834);
nor U315 (N_315,In_1148,In_452);
nor U316 (N_316,In_1204,In_2168);
or U317 (N_317,In_458,In_292);
nand U318 (N_318,In_466,In_55);
and U319 (N_319,In_372,In_524);
nor U320 (N_320,In_937,In_2661);
or U321 (N_321,In_2547,In_2259);
or U322 (N_322,In_1509,In_628);
nand U323 (N_323,In_1787,In_1448);
and U324 (N_324,In_2869,In_737);
or U325 (N_325,In_2153,In_1271);
nor U326 (N_326,In_2847,In_1982);
xnor U327 (N_327,In_896,In_812);
xnor U328 (N_328,In_1299,In_2897);
or U329 (N_329,In_1647,In_272);
nor U330 (N_330,In_2409,In_1167);
nand U331 (N_331,In_1836,In_904);
xnor U332 (N_332,In_36,In_1467);
or U333 (N_333,In_289,In_314);
or U334 (N_334,In_2290,In_1617);
nand U335 (N_335,In_2363,In_43);
xnor U336 (N_336,In_2945,In_1242);
xor U337 (N_337,In_2796,In_1256);
nand U338 (N_338,In_2443,In_1140);
or U339 (N_339,In_955,In_2662);
and U340 (N_340,In_1688,In_2693);
nand U341 (N_341,In_2034,In_410);
nor U342 (N_342,In_1134,In_177);
nand U343 (N_343,In_1362,In_493);
xor U344 (N_344,In_303,In_26);
and U345 (N_345,In_734,In_2883);
xnor U346 (N_346,In_573,In_1650);
nand U347 (N_347,In_710,In_591);
nor U348 (N_348,In_1475,In_1233);
xor U349 (N_349,In_1025,In_34);
nand U350 (N_350,In_2166,In_1731);
nand U351 (N_351,In_1682,In_1906);
and U352 (N_352,In_2772,In_121);
or U353 (N_353,In_2,In_2837);
xor U354 (N_354,In_2356,In_1194);
or U355 (N_355,In_47,In_608);
and U356 (N_356,In_1414,In_1989);
nor U357 (N_357,In_181,In_1072);
or U358 (N_358,In_2154,In_1684);
or U359 (N_359,In_1595,In_2558);
or U360 (N_360,In_855,In_888);
nor U361 (N_361,In_849,In_2513);
nor U362 (N_362,In_1456,In_2447);
xnor U363 (N_363,In_2700,In_976);
or U364 (N_364,In_1240,In_1003);
or U365 (N_365,In_541,In_2734);
xnor U366 (N_366,In_500,In_2327);
and U367 (N_367,In_1766,In_2181);
nor U368 (N_368,In_727,In_355);
xor U369 (N_369,In_1581,In_2775);
nand U370 (N_370,In_2479,In_2905);
nor U371 (N_371,In_66,In_2412);
and U372 (N_372,In_1320,In_1138);
and U373 (N_373,In_1364,In_1553);
xnor U374 (N_374,In_403,In_2865);
and U375 (N_375,In_2721,In_240);
nor U376 (N_376,In_1466,In_1486);
or U377 (N_377,In_1452,In_1765);
or U378 (N_378,In_2037,In_337);
xor U379 (N_379,In_1286,In_1917);
xnor U380 (N_380,In_1843,In_2631);
nand U381 (N_381,In_1761,In_1985);
or U382 (N_382,In_726,In_1057);
and U383 (N_383,In_610,In_2041);
or U384 (N_384,In_2616,In_2600);
and U385 (N_385,In_805,In_2064);
and U386 (N_386,In_969,In_532);
xor U387 (N_387,In_552,In_1872);
or U388 (N_388,In_2768,In_48);
and U389 (N_389,In_766,In_2445);
or U390 (N_390,In_2174,In_1646);
and U391 (N_391,In_983,In_1909);
nand U392 (N_392,In_448,In_2784);
xnor U393 (N_393,In_2606,In_2459);
xor U394 (N_394,In_897,In_431);
nand U395 (N_395,In_936,In_14);
xor U396 (N_396,In_1986,In_2035);
nor U397 (N_397,In_2767,In_2728);
nand U398 (N_398,In_2217,In_669);
nor U399 (N_399,In_1432,In_774);
or U400 (N_400,In_903,In_340);
and U401 (N_401,In_1739,In_134);
nand U402 (N_402,In_2871,In_276);
nand U403 (N_403,In_2541,In_799);
and U404 (N_404,In_683,In_1339);
xor U405 (N_405,In_1667,In_1676);
and U406 (N_406,In_1054,In_2692);
xor U407 (N_407,In_449,In_1422);
xor U408 (N_408,In_2833,In_168);
nand U409 (N_409,In_510,In_1284);
nand U410 (N_410,In_326,In_975);
nor U411 (N_411,In_40,In_623);
nor U412 (N_412,In_436,In_838);
and U413 (N_413,In_1806,In_990);
nor U414 (N_414,In_804,In_2569);
nor U415 (N_415,In_2108,In_968);
nor U416 (N_416,In_1131,In_2657);
and U417 (N_417,In_2111,In_2788);
nor U418 (N_418,In_2080,In_1564);
and U419 (N_419,In_588,In_2527);
or U420 (N_420,In_1172,In_1567);
and U421 (N_421,In_164,In_2673);
nor U422 (N_422,In_2171,In_1609);
or U423 (N_423,In_1960,In_2487);
or U424 (N_424,In_185,In_2520);
nor U425 (N_425,In_2560,In_1160);
xnor U426 (N_426,In_2282,In_147);
xor U427 (N_427,In_2628,In_2754);
nand U428 (N_428,In_1168,In_2397);
nand U429 (N_429,In_1144,In_1449);
xnor U430 (N_430,In_1125,In_606);
and U431 (N_431,In_1088,In_2874);
and U432 (N_432,In_2568,In_1471);
nor U433 (N_433,In_694,In_2549);
and U434 (N_434,In_1886,In_1772);
nand U435 (N_435,In_1703,In_748);
or U436 (N_436,In_2882,In_2436);
xor U437 (N_437,In_1962,In_2151);
or U438 (N_438,In_978,In_1788);
nand U439 (N_439,In_2446,In_1838);
xor U440 (N_440,In_2324,In_2297);
or U441 (N_441,In_533,In_2403);
nor U442 (N_442,In_1687,In_2464);
xnor U443 (N_443,In_542,In_2745);
nor U444 (N_444,In_1665,In_382);
xor U445 (N_445,In_2918,In_2984);
and U446 (N_446,In_1698,In_1773);
xnor U447 (N_447,In_483,In_1139);
xor U448 (N_448,In_707,In_2751);
nand U449 (N_449,In_1958,In_172);
and U450 (N_450,In_1730,In_580);
nand U451 (N_451,In_2302,In_2263);
and U452 (N_452,In_296,In_1346);
and U453 (N_453,In_2564,In_907);
nor U454 (N_454,In_2696,In_1774);
or U455 (N_455,In_2467,In_2469);
and U456 (N_456,In_832,In_1415);
nand U457 (N_457,In_1375,In_238);
nand U458 (N_458,In_860,In_1376);
nand U459 (N_459,In_1040,In_1789);
nor U460 (N_460,In_2500,In_2183);
and U461 (N_461,In_1749,In_1763);
nand U462 (N_462,In_671,In_1225);
and U463 (N_463,In_2272,In_609);
and U464 (N_464,In_1437,In_1303);
nor U465 (N_465,In_2378,In_574);
nor U466 (N_466,In_1944,In_453);
xnor U467 (N_467,In_988,In_39);
or U468 (N_468,In_2593,In_2736);
or U469 (N_469,In_1529,In_634);
nor U470 (N_470,In_116,In_2757);
and U471 (N_471,In_2857,In_900);
nand U472 (N_472,In_2161,In_439);
nand U473 (N_473,In_166,In_1455);
xor U474 (N_474,In_1556,In_2326);
and U475 (N_475,In_504,In_362);
nor U476 (N_476,In_102,In_2368);
xnor U477 (N_477,In_2310,In_1019);
or U478 (N_478,In_914,In_259);
nor U479 (N_479,In_1094,In_547);
or U480 (N_480,In_2010,In_2888);
xor U481 (N_481,In_868,In_2947);
or U482 (N_482,In_1498,In_681);
nand U483 (N_483,In_2177,In_377);
nand U484 (N_484,In_455,In_2227);
and U485 (N_485,In_329,In_2777);
nand U486 (N_486,In_675,In_19);
xnor U487 (N_487,In_746,In_1936);
nor U488 (N_488,In_331,In_2634);
nand U489 (N_489,In_2789,In_1736);
nor U490 (N_490,In_2766,In_93);
nor U491 (N_491,In_408,In_2067);
and U492 (N_492,In_2695,In_962);
nand U493 (N_493,In_738,In_1741);
and U494 (N_494,In_517,In_755);
or U495 (N_495,In_616,In_1606);
nand U496 (N_496,In_2280,In_2517);
nor U497 (N_497,In_160,In_2910);
nor U498 (N_498,In_1478,In_882);
nand U499 (N_499,In_1016,In_2717);
or U500 (N_500,In_2762,In_2765);
xnor U501 (N_501,In_638,In_374);
and U502 (N_502,In_1919,In_1642);
nor U503 (N_503,In_1558,In_2642);
or U504 (N_504,In_2672,In_2463);
nor U505 (N_505,In_140,In_2261);
xor U506 (N_506,In_2205,In_153);
nor U507 (N_507,In_1117,In_1163);
nand U508 (N_508,In_2240,In_162);
or U509 (N_509,In_863,In_1897);
or U510 (N_510,In_546,In_2709);
and U511 (N_511,In_1250,In_225);
xor U512 (N_512,In_2771,In_2916);
nand U513 (N_513,In_1342,In_2019);
nand U514 (N_514,In_1661,In_2831);
xnor U515 (N_515,In_1814,In_593);
or U516 (N_516,In_709,In_1333);
xor U517 (N_517,In_462,In_1178);
and U518 (N_518,In_723,In_136);
and U519 (N_519,In_641,In_27);
or U520 (N_520,In_1626,In_925);
nand U521 (N_521,In_555,In_2352);
nand U522 (N_522,In_2781,In_1062);
xnor U523 (N_523,In_2264,In_2401);
nor U524 (N_524,In_435,In_231);
nand U525 (N_525,In_2870,In_1022);
xor U526 (N_526,In_994,In_2349);
nor U527 (N_527,In_1802,In_2279);
nand U528 (N_528,In_1191,In_2242);
nand U529 (N_529,In_270,In_365);
or U530 (N_530,In_930,In_1298);
or U531 (N_531,In_1500,In_1945);
nor U532 (N_532,In_2507,In_973);
or U533 (N_533,In_1977,In_1781);
nand U534 (N_534,In_984,In_196);
nand U535 (N_535,In_827,In_878);
nand U536 (N_536,In_2208,In_889);
or U537 (N_537,In_2643,In_2328);
xnor U538 (N_538,In_2203,In_194);
nand U539 (N_539,In_934,In_228);
and U540 (N_540,In_2357,In_784);
and U541 (N_541,In_2758,In_2605);
nor U542 (N_542,In_519,In_1879);
or U543 (N_543,In_2801,In_654);
nand U544 (N_544,In_2128,In_1387);
or U545 (N_545,In_522,In_1060);
xor U546 (N_546,In_2102,In_795);
nand U547 (N_547,In_779,In_815);
and U548 (N_548,In_12,In_847);
nand U549 (N_549,In_2995,In_2139);
or U550 (N_550,In_679,In_278);
or U551 (N_551,In_2805,In_44);
xor U552 (N_552,In_956,In_1747);
or U553 (N_553,In_1884,In_2404);
or U554 (N_554,In_2246,In_2275);
or U555 (N_555,In_2633,In_2157);
nand U556 (N_556,In_1245,In_2506);
xor U557 (N_557,In_2392,In_2731);
nor U558 (N_558,In_2262,In_1098);
nand U559 (N_559,In_170,In_2794);
xor U560 (N_560,In_1169,In_25);
or U561 (N_561,In_1544,In_1321);
and U562 (N_562,In_1327,In_143);
or U563 (N_563,In_506,In_1324);
xnor U564 (N_564,In_2391,In_2976);
nand U565 (N_565,In_360,In_2935);
nand U566 (N_566,In_2082,In_1370);
or U567 (N_567,In_924,In_702);
nor U568 (N_568,In_2690,In_1156);
xnor U569 (N_569,In_651,In_1315);
nand U570 (N_570,In_1151,In_2567);
xnor U571 (N_571,In_2563,In_1211);
xnor U572 (N_572,In_18,In_396);
and U573 (N_573,In_1360,In_1383);
or U574 (N_574,In_2360,In_767);
nor U575 (N_575,In_2504,In_1794);
nand U576 (N_576,In_1685,In_2946);
nand U577 (N_577,In_1289,In_2622);
nand U578 (N_578,In_2314,In_980);
and U579 (N_579,In_250,In_2025);
and U580 (N_580,In_1396,In_1070);
xnor U581 (N_581,In_2237,In_1639);
or U582 (N_582,In_176,In_2704);
xnor U583 (N_583,In_1371,In_2635);
nor U584 (N_584,In_1119,In_445);
or U585 (N_585,In_1548,In_1967);
xnor U586 (N_586,In_52,In_1796);
xor U587 (N_587,In_2637,In_479);
and U588 (N_588,In_1102,In_966);
xnor U589 (N_589,In_2791,In_1394);
nor U590 (N_590,In_515,In_926);
xnor U591 (N_591,In_1300,In_2288);
nor U592 (N_592,In_2926,In_2708);
and U593 (N_593,In_1050,In_2298);
or U594 (N_594,In_1552,In_2466);
xor U595 (N_595,In_443,In_1504);
and U596 (N_596,In_1197,In_1928);
and U597 (N_597,In_2160,In_2451);
nor U598 (N_598,In_2598,In_1503);
nor U599 (N_599,In_2619,In_2555);
and U600 (N_600,In_244,In_782);
and U601 (N_601,In_2932,In_2243);
or U602 (N_602,In_985,In_2534);
xor U603 (N_603,In_2653,In_595);
and U604 (N_604,In_1840,In_1652);
or U605 (N_605,In_1575,In_605);
and U606 (N_606,In_1798,In_2738);
nor U607 (N_607,In_644,In_138);
nand U608 (N_608,In_1384,In_1469);
and U609 (N_609,In_592,In_2103);
or U610 (N_610,In_1780,In_1924);
nand U611 (N_611,In_1598,In_1184);
xor U612 (N_612,In_2271,In_1708);
and U613 (N_613,In_1497,In_563);
nand U614 (N_614,In_1574,In_1769);
nor U615 (N_615,In_594,In_6);
or U616 (N_616,In_1629,In_2521);
or U617 (N_617,In_1488,In_695);
or U618 (N_618,In_1472,In_1516);
nand U619 (N_619,In_1485,In_2364);
and U620 (N_620,In_2747,In_652);
and U621 (N_621,In_1217,In_2253);
nand U622 (N_622,In_1274,In_1171);
nand U623 (N_623,In_1494,In_1092);
nor U624 (N_624,In_1657,In_1302);
nor U625 (N_625,In_632,In_2105);
and U626 (N_626,In_251,In_2987);
xnor U627 (N_627,In_1029,In_2367);
nor U628 (N_628,In_816,In_1325);
or U629 (N_629,In_1066,In_457);
nor U630 (N_630,In_2267,In_2956);
and U631 (N_631,In_1413,In_2741);
or U632 (N_632,In_1329,In_1004);
xor U633 (N_633,In_85,In_1720);
and U634 (N_634,In_2536,In_385);
or U635 (N_635,In_1128,In_406);
xor U636 (N_636,In_696,In_835);
nor U637 (N_637,In_2222,In_2714);
nand U638 (N_638,In_1464,In_461);
nand U639 (N_639,In_96,In_2604);
or U640 (N_640,In_2106,In_911);
xor U641 (N_641,In_2341,In_2908);
nor U642 (N_642,In_718,In_1525);
or U643 (N_643,In_317,In_328);
nand U644 (N_644,In_2126,In_389);
or U645 (N_645,In_1587,In_2792);
and U646 (N_646,In_1903,In_2856);
nor U647 (N_647,In_1069,In_1998);
or U648 (N_648,In_1263,In_1075);
nor U649 (N_649,In_569,In_258);
or U650 (N_650,In_1221,In_750);
and U651 (N_651,In_1046,In_2930);
and U652 (N_652,In_2448,In_2109);
nand U653 (N_653,In_1491,In_2462);
nand U654 (N_654,In_1733,In_1849);
and U655 (N_655,In_1341,In_2806);
xnor U656 (N_656,In_713,In_1322);
and U657 (N_657,In_1463,In_91);
nor U658 (N_658,In_1856,In_1115);
nor U659 (N_659,In_2773,In_29);
and U660 (N_660,In_2143,In_1812);
and U661 (N_661,In_1513,In_7);
and U662 (N_662,In_996,In_1317);
or U663 (N_663,In_2377,In_2110);
and U664 (N_664,In_1379,In_2454);
nor U665 (N_665,In_1259,In_705);
nand U666 (N_666,In_1835,In_1651);
xnor U667 (N_667,In_2967,In_295);
and U668 (N_668,In_2658,In_1920);
xnor U669 (N_669,In_1877,In_229);
nand U670 (N_670,In_2583,In_2114);
xor U671 (N_671,In_223,In_902);
xor U672 (N_672,In_212,In_2578);
and U673 (N_673,In_2994,In_2526);
and U674 (N_674,In_2428,In_1807);
and U675 (N_675,In_2148,In_1435);
and U676 (N_676,In_387,In_525);
nand U677 (N_677,In_2550,In_280);
nor U678 (N_678,In_261,In_947);
xor U679 (N_679,In_2720,In_1753);
nand U680 (N_680,In_987,In_2084);
and U681 (N_681,In_1551,In_712);
nand U682 (N_682,In_2483,In_106);
nor U683 (N_683,In_2277,In_2851);
nor U684 (N_684,In_1875,In_1621);
and U685 (N_685,In_2607,In_2425);
or U686 (N_686,In_2473,In_516);
nor U687 (N_687,In_2371,In_2340);
or U688 (N_688,In_841,In_2858);
nand U689 (N_689,In_2989,In_469);
or U690 (N_690,In_2422,In_215);
nand U691 (N_691,In_2444,In_2933);
nand U692 (N_692,In_1623,In_294);
nor U693 (N_693,In_699,In_1890);
xnor U694 (N_694,In_539,In_1175);
and U695 (N_695,In_2687,In_1592);
xor U696 (N_696,In_1999,In_2224);
nor U697 (N_697,In_1196,In_1369);
or U698 (N_698,In_1424,In_2150);
nor U699 (N_699,In_2716,In_2841);
nand U700 (N_700,In_1232,In_599);
nand U701 (N_701,In_576,In_484);
nand U702 (N_702,In_1743,In_70);
nand U703 (N_703,In_2922,In_368);
nand U704 (N_704,In_2678,In_1632);
xnor U705 (N_705,In_2178,In_2911);
or U706 (N_706,In_206,In_977);
xnor U707 (N_707,In_2848,In_1805);
and U708 (N_708,In_803,In_2862);
or U709 (N_709,In_529,In_2689);
and U710 (N_710,In_2394,In_1479);
and U711 (N_711,In_423,In_2899);
or U712 (N_712,In_811,In_2724);
nand U713 (N_713,In_2697,In_1510);
nand U714 (N_714,In_2969,In_2044);
nand U715 (N_715,In_2281,In_313);
or U716 (N_716,In_1358,In_1418);
nand U717 (N_717,In_46,In_1561);
xnor U718 (N_718,In_1619,In_2001);
and U719 (N_719,In_135,In_1458);
or U720 (N_720,In_333,In_81);
xnor U721 (N_721,In_2236,In_182);
nand U722 (N_722,In_456,In_13);
xnor U723 (N_723,In_2729,In_1895);
nor U724 (N_724,In_2942,In_2991);
nand U725 (N_725,In_1711,In_1883);
or U726 (N_726,In_1597,In_2119);
nand U727 (N_727,In_1746,In_1946);
nand U728 (N_728,In_1648,In_2410);
or U729 (N_729,In_1602,In_2104);
and U730 (N_730,In_1568,In_222);
nand U731 (N_731,In_615,In_2062);
or U732 (N_732,In_2572,In_724);
nor U733 (N_733,In_1164,In_2172);
or U734 (N_734,In_2362,In_2559);
nand U735 (N_735,In_256,In_2134);
and U736 (N_736,In_2132,In_1810);
or U737 (N_737,In_0,In_514);
nor U738 (N_738,In_1208,In_1935);
and U739 (N_739,In_1712,In_2185);
nor U740 (N_740,In_558,In_1326);
and U741 (N_741,In_1825,In_304);
xnor U742 (N_742,In_1354,In_1201);
and U743 (N_743,In_2235,In_489);
xor U744 (N_744,In_661,In_2121);
nor U745 (N_745,In_434,In_564);
and U746 (N_746,In_2329,In_2691);
or U747 (N_747,In_41,In_825);
nand U748 (N_748,In_625,In_2049);
xnor U749 (N_749,In_1077,In_548);
or U750 (N_750,In_1912,In_757);
nor U751 (N_751,In_2973,In_2193);
xor U752 (N_752,In_2682,In_471);
xor U753 (N_753,In_1760,In_99);
and U754 (N_754,In_1737,In_2960);
xnor U755 (N_755,In_1978,In_818);
xnor U756 (N_756,In_508,In_2670);
nand U757 (N_757,In_2300,In_952);
nand U758 (N_758,In_1433,In_1521);
and U759 (N_759,In_1359,In_2433);
xor U760 (N_760,In_111,In_2421);
and U761 (N_761,In_791,In_571);
or U762 (N_762,In_1892,In_78);
nand U763 (N_763,In_1528,In_657);
or U764 (N_764,In_131,In_1293);
xnor U765 (N_765,In_1231,In_1001);
and U766 (N_766,In_488,In_682);
xor U767 (N_767,In_2779,In_739);
or U768 (N_768,In_2029,In_1291);
or U769 (N_769,In_2959,In_1876);
nor U770 (N_770,In_2239,In_2861);
nor U771 (N_771,In_2125,In_2390);
xor U772 (N_772,In_1845,In_2216);
xnor U773 (N_773,In_2824,In_898);
or U774 (N_774,In_824,In_1878);
xnor U775 (N_775,In_783,In_2348);
or U776 (N_776,In_1732,In_1030);
or U777 (N_777,In_1382,In_219);
nor U778 (N_778,In_798,In_427);
nand U779 (N_779,In_1547,In_370);
nand U780 (N_780,In_1489,In_16);
or U781 (N_781,In_1555,In_1202);
or U782 (N_782,In_523,In_1990);
nand U783 (N_783,In_171,In_1135);
nand U784 (N_784,In_887,In_2260);
and U785 (N_785,In_1600,In_1948);
nand U786 (N_786,In_1554,In_2735);
or U787 (N_787,In_1930,In_115);
or U788 (N_788,In_1058,In_1588);
or U789 (N_789,In_31,In_1888);
nor U790 (N_790,In_1992,In_1220);
xnor U791 (N_791,In_1988,In_369);
xnor U792 (N_792,In_1636,In_2278);
nand U793 (N_793,In_2099,In_2860);
or U794 (N_794,In_394,In_2815);
nand U795 (N_795,In_2826,In_2191);
and U796 (N_796,In_447,In_1957);
or U797 (N_797,In_1822,In_2725);
nand U798 (N_798,In_2674,In_2840);
xor U799 (N_799,In_894,In_2149);
nand U800 (N_800,In_2232,In_2798);
and U801 (N_801,In_793,In_2287);
and U802 (N_802,In_833,In_2940);
xnor U803 (N_803,In_1818,In_1014);
and U804 (N_804,In_1519,In_2998);
nor U805 (N_805,In_754,In_459);
or U806 (N_806,In_1275,In_2014);
and U807 (N_807,In_1312,In_2510);
or U808 (N_808,In_1190,In_2685);
xnor U809 (N_809,In_2701,In_1421);
or U810 (N_810,In_2978,In_2184);
xor U811 (N_811,In_866,In_2122);
nor U812 (N_812,In_2683,In_220);
nor U813 (N_813,In_1693,In_127);
and U814 (N_814,In_83,In_2167);
or U815 (N_815,In_1570,In_2760);
nand U816 (N_816,In_175,In_1572);
and U817 (N_817,In_5,In_944);
nand U818 (N_818,In_1023,In_1975);
nand U819 (N_819,In_584,In_2120);
or U820 (N_820,In_2892,In_2875);
xor U821 (N_821,In_1680,In_2962);
or U822 (N_822,In_56,In_1198);
and U823 (N_823,In_613,In_912);
nand U824 (N_824,In_1839,In_772);
or U825 (N_825,In_602,In_2501);
nand U826 (N_826,In_2929,In_2533);
and U827 (N_827,In_881,In_2621);
and U828 (N_828,In_149,In_200);
and U829 (N_829,In_1804,In_2465);
nor U830 (N_830,In_1816,In_35);
nand U831 (N_831,In_1101,In_1120);
nand U832 (N_832,In_2086,In_1388);
or U833 (N_833,In_487,In_193);
or U834 (N_834,In_2993,In_778);
nor U835 (N_835,In_69,In_823);
xnor U836 (N_836,In_1881,In_1372);
xor U837 (N_837,In_1782,In_2859);
nand U838 (N_838,In_864,In_191);
nor U839 (N_839,In_1543,In_4);
nor U840 (N_840,In_2509,In_1277);
xnor U841 (N_841,In_2395,In_663);
or U842 (N_842,In_837,In_2999);
nand U843 (N_843,In_386,In_2854);
xnor U844 (N_844,In_418,In_1799);
and U845 (N_845,In_2823,In_2665);
or U846 (N_846,In_1974,In_1735);
xnor U847 (N_847,In_2737,In_614);
or U848 (N_848,In_995,In_2015);
or U849 (N_849,In_2966,In_156);
and U850 (N_850,In_660,In_1790);
or U851 (N_851,In_2101,In_1133);
or U852 (N_852,In_2485,In_554);
nor U853 (N_853,In_1848,In_243);
xnor U854 (N_854,In_1439,In_189);
and U855 (N_855,In_2244,In_24);
nor U856 (N_856,In_2230,In_1273);
or U857 (N_857,In_2450,In_1826);
nand U858 (N_858,In_2358,In_117);
nor U859 (N_859,In_2723,In_1002);
and U860 (N_860,In_1453,In_1700);
nand U861 (N_861,In_1122,In_494);
and U862 (N_862,In_2964,In_1701);
xor U863 (N_863,In_501,In_179);
or U864 (N_864,In_943,In_1244);
xnor U865 (N_865,In_1083,In_201);
xor U866 (N_866,In_1116,In_1847);
nand U867 (N_867,In_90,In_1304);
nor U868 (N_868,In_161,In_2898);
nor U869 (N_869,In_2756,In_2496);
or U870 (N_870,In_1882,In_2407);
and U871 (N_871,In_1604,In_407);
xnor U872 (N_872,In_1970,In_1352);
nor U873 (N_873,In_2582,In_92);
nand U874 (N_874,In_974,In_1511);
xnor U875 (N_875,In_2481,In_2145);
or U876 (N_876,In_2838,In_476);
nor U877 (N_877,In_1188,In_2097);
or U878 (N_878,In_534,In_1859);
nand U879 (N_879,In_2060,In_945);
nand U880 (N_880,In_2975,In_2524);
nand U881 (N_881,In_348,In_2951);
nor U882 (N_882,In_1535,In_485);
nand U883 (N_883,In_2546,In_1389);
nor U884 (N_884,In_1800,In_100);
nand U885 (N_885,In_169,In_1296);
nor U886 (N_886,In_2269,In_2000);
xnor U887 (N_887,In_961,In_359);
or U888 (N_888,In_391,In_2535);
nor U889 (N_889,In_1896,In_167);
or U890 (N_890,In_2925,In_502);
nand U891 (N_891,In_249,In_1618);
or U892 (N_892,In_2834,In_2164);
nor U893 (N_893,In_1150,In_2884);
nor U894 (N_894,In_1757,In_1740);
and U895 (N_895,In_1939,In_2304);
and U896 (N_896,In_2799,In_119);
and U897 (N_897,In_163,In_971);
nand U898 (N_898,In_433,In_2992);
nor U899 (N_899,In_2016,In_2405);
nor U900 (N_900,In_2957,In_2250);
or U901 (N_901,In_670,In_879);
xor U902 (N_902,In_846,In_848);
or U903 (N_903,In_322,In_697);
nand U904 (N_904,In_2055,In_1793);
nor U905 (N_905,In_2955,In_624);
xor U906 (N_906,In_1087,In_1316);
and U907 (N_907,In_1355,In_717);
and U908 (N_908,In_2226,In_1499);
and U909 (N_909,In_388,In_2894);
or U910 (N_910,In_357,In_87);
xnor U911 (N_911,In_1653,In_1801);
nor U912 (N_912,In_2599,In_151);
nor U913 (N_913,In_1710,In_678);
and U914 (N_914,In_1518,In_1699);
and U915 (N_915,In_241,In_1533);
xor U916 (N_916,In_810,In_1307);
nor U917 (N_917,In_2040,In_1443);
and U918 (N_918,In_378,In_1484);
nor U919 (N_919,In_475,In_339);
nor U920 (N_920,In_581,In_2478);
nor U921 (N_921,In_2344,In_1097);
nand U922 (N_922,In_1012,In_1481);
nor U923 (N_923,In_690,In_749);
or U924 (N_924,In_1855,In_1438);
or U925 (N_925,In_497,In_2374);
xor U926 (N_926,In_271,In_941);
or U927 (N_927,In_553,In_578);
nor U928 (N_928,In_2449,In_1968);
xor U929 (N_929,In_950,In_2981);
nand U930 (N_930,In_77,In_2804);
nor U931 (N_931,In_1718,In_2618);
nor U932 (N_932,In_1921,In_1979);
and U933 (N_933,In_2225,In_1440);
or U934 (N_934,In_23,In_1235);
nor U935 (N_935,In_2113,In_2886);
xor U936 (N_936,In_1267,In_1308);
nand U937 (N_937,In_2257,In_1385);
and U938 (N_938,In_2739,In_2822);
xor U939 (N_939,In_1219,In_2943);
nand U940 (N_940,In_2005,In_2063);
or U941 (N_941,In_1715,In_1622);
and U942 (N_942,In_64,In_2977);
nand U943 (N_943,In_1205,In_2472);
nor U944 (N_944,In_310,In_931);
xnor U945 (N_945,In_998,In_2194);
or U946 (N_946,In_2388,In_1223);
xor U947 (N_947,In_1603,In_2632);
xor U948 (N_948,In_2411,In_2317);
or U949 (N_949,In_2850,In_1254);
and U950 (N_950,In_1914,In_2864);
and U951 (N_951,In_2333,In_139);
nor U952 (N_952,In_1247,In_1209);
xnor U953 (N_953,In_2270,In_2301);
xnor U954 (N_954,In_1949,In_1055);
xor U955 (N_955,In_2812,In_2629);
or U956 (N_956,In_759,In_1335);
or U957 (N_957,In_865,In_412);
and U958 (N_958,In_526,In_2012);
and U959 (N_959,In_159,In_60);
or U960 (N_960,In_28,In_393);
and U961 (N_961,In_1261,In_373);
nor U962 (N_962,In_1153,In_1113);
xor U963 (N_963,In_1562,In_33);
xor U964 (N_964,In_2952,In_1786);
nand U965 (N_965,In_390,In_126);
or U966 (N_966,In_350,In_419);
xnor U967 (N_967,In_2141,In_283);
and U968 (N_968,In_2337,In_790);
xnor U969 (N_969,In_1887,In_745);
and U970 (N_970,In_1563,In_2881);
and U971 (N_971,In_275,In_2680);
and U972 (N_972,In_1908,In_531);
and U973 (N_973,In_2440,In_1922);
or U974 (N_974,In_2241,In_1199);
and U975 (N_975,In_79,In_2215);
or U976 (N_976,In_2198,In_1668);
or U977 (N_977,In_263,In_2846);
xnor U978 (N_978,In_2372,In_195);
xor U979 (N_979,In_1507,In_1725);
or U980 (N_980,In_428,In_1431);
nor U981 (N_981,In_764,In_95);
nor U982 (N_982,In_1214,In_735);
nand U983 (N_983,In_2078,In_2438);
xor U984 (N_984,In_929,In_110);
and U985 (N_985,In_1549,In_247);
or U986 (N_986,In_1582,In_402);
or U987 (N_987,In_1837,In_1287);
or U988 (N_988,In_1226,In_2038);
nor U989 (N_989,In_1996,In_1262);
and U990 (N_990,In_1702,In_1910);
nand U991 (N_991,In_2668,In_300);
or U992 (N_992,In_910,In_2816);
and U993 (N_993,In_2306,In_1336);
xnor U994 (N_994,In_1180,In_1557);
nand U995 (N_995,In_2295,In_2742);
or U996 (N_996,In_1195,In_1620);
nor U997 (N_997,In_1314,In_1343);
nor U998 (N_998,In_1791,In_1251);
and U999 (N_999,In_551,In_2523);
xnor U1000 (N_1000,In_22,In_1635);
nand U1001 (N_1001,In_1679,In_1566);
xnor U1002 (N_1002,In_1984,In_307);
and U1003 (N_1003,In_2071,In_2107);
nand U1004 (N_1004,In_1056,In_659);
and U1005 (N_1005,In_1086,In_2266);
nand U1006 (N_1006,In_1141,In_560);
nor U1007 (N_1007,In_1964,In_731);
nor U1008 (N_1008,In_2054,In_2927);
xor U1009 (N_1009,In_596,In_2343);
and U1010 (N_1010,In_2915,In_2651);
or U1011 (N_1011,In_1474,In_645);
nand U1012 (N_1012,In_1446,In_80);
or U1013 (N_1013,In_145,In_1674);
nor U1014 (N_1014,In_1234,In_1916);
nand U1015 (N_1015,In_1146,In_451);
nor U1016 (N_1016,In_2832,In_1540);
nor U1017 (N_1017,In_2284,In_1638);
nand U1018 (N_1018,In_1795,In_1863);
nor U1019 (N_1019,In_586,In_2115);
nor U1020 (N_1020,In_1797,In_204);
or U1021 (N_1021,In_65,In_686);
and U1022 (N_1022,In_1577,In_851);
nor U1023 (N_1023,In_640,In_463);
nand U1024 (N_1024,In_2032,In_1857);
xor U1025 (N_1025,In_633,In_957);
nand U1026 (N_1026,In_920,In_2283);
or U1027 (N_1027,In_646,In_2494);
nand U1028 (N_1028,In_1940,In_2877);
nand U1029 (N_1029,In_444,In_877);
nor U1030 (N_1030,In_2528,In_202);
and U1031 (N_1031,In_928,In_1744);
nand U1032 (N_1032,In_2414,In_1541);
or U1033 (N_1033,In_1123,In_2554);
nand U1034 (N_1034,In_693,In_1565);
and U1035 (N_1035,In_1108,In_1585);
and U1036 (N_1036,In_2800,In_2321);
xor U1037 (N_1037,In_2047,In_54);
nor U1038 (N_1038,In_2204,In_2671);
xor U1039 (N_1039,In_2924,In_2162);
xor U1040 (N_1040,In_1059,In_1611);
nor U1041 (N_1041,In_2983,In_1187);
nand U1042 (N_1042,In_438,In_1268);
or U1043 (N_1043,In_1673,In_2188);
xor U1044 (N_1044,In_1520,In_2703);
nand U1045 (N_1045,In_2825,In_2223);
nand U1046 (N_1046,In_2715,In_1677);
and U1047 (N_1047,In_630,In_2733);
and U1048 (N_1048,In_2782,In_708);
nor U1049 (N_1049,In_2074,In_1832);
and U1050 (N_1050,In_1311,In_2787);
or U1051 (N_1051,In_1492,In_817);
nor U1052 (N_1052,In_2958,In_1319);
and U1053 (N_1053,In_1865,In_401);
or U1054 (N_1054,In_2138,In_528);
nand U1055 (N_1055,In_1255,In_188);
nor U1056 (N_1056,In_442,In_133);
or U1057 (N_1057,In_1641,In_1973);
and U1058 (N_1058,In_2355,In_316);
nor U1059 (N_1059,In_2913,In_1078);
nand U1060 (N_1060,In_123,In_874);
nand U1061 (N_1061,In_1738,In_309);
nand U1062 (N_1062,In_1559,In_2229);
and U1063 (N_1063,In_2868,In_1111);
nand U1064 (N_1064,In_1454,In_967);
nand U1065 (N_1065,In_565,In_2896);
nor U1066 (N_1066,In_1309,In_1417);
xor U1067 (N_1067,In_1363,In_1393);
and U1068 (N_1068,In_1956,In_1686);
xnor U1069 (N_1069,In_1395,In_207);
nor U1070 (N_1070,In_2744,In_2920);
and U1071 (N_1071,In_245,In_1155);
nand U1072 (N_1072,In_785,In_467);
nor U1073 (N_1073,In_2091,In_2639);
or U1074 (N_1074,In_1053,In_836);
and U1075 (N_1075,In_2602,In_2330);
nor U1076 (N_1076,In_1965,In_118);
or U1077 (N_1077,In_1546,In_1093);
or U1078 (N_1078,In_2797,In_677);
nand U1079 (N_1079,In_826,In_1200);
nor U1080 (N_1080,In_964,In_2366);
nor U1081 (N_1081,In_1124,In_2003);
nand U1082 (N_1082,In_2698,In_1026);
xor U1083 (N_1083,In_1037,In_1593);
and U1084 (N_1084,In_2666,In_2090);
and U1085 (N_1085,In_2713,In_1993);
xor U1086 (N_1086,In_1522,In_2127);
or U1087 (N_1087,In_2165,In_687);
or U1088 (N_1088,In_120,In_2470);
nand U1089 (N_1089,In_1306,In_2176);
nand U1090 (N_1090,In_2979,In_165);
or U1091 (N_1091,In_1869,In_585);
nor U1092 (N_1092,In_2323,In_1292);
nand U1093 (N_1093,In_1278,In_570);
xor U1094 (N_1094,In_736,In_174);
nand U1095 (N_1095,In_74,In_1966);
nor U1096 (N_1096,In_1870,In_1927);
or U1097 (N_1097,In_970,In_568);
nor U1098 (N_1098,In_417,In_2810);
xnor U1099 (N_1099,In_415,In_1282);
nand U1100 (N_1100,In_1118,In_297);
xnor U1101 (N_1101,In_884,In_208);
nand U1102 (N_1102,In_2382,In_939);
nor U1103 (N_1103,In_2589,In_725);
nand U1104 (N_1104,In_829,In_1495);
nand U1105 (N_1105,In_1043,In_621);
nor U1106 (N_1106,In_740,In_1808);
or U1107 (N_1107,In_2061,In_701);
and U1108 (N_1108,In_2562,In_395);
xor U1109 (N_1109,In_1206,In_2710);
xor U1110 (N_1110,In_618,In_1033);
or U1111 (N_1111,In_626,In_991);
and U1112 (N_1112,In_1596,In_1073);
and U1113 (N_1113,In_802,In_993);
nand U1114 (N_1114,In_704,In_2627);
and U1115 (N_1115,In_1854,In_1655);
nand U1116 (N_1116,In_305,In_1203);
nor U1117 (N_1117,In_1694,In_1980);
or U1118 (N_1118,In_1407,In_199);
and U1119 (N_1119,In_1612,In_1943);
xor U1120 (N_1120,In_2571,In_773);
or U1121 (N_1121,In_2458,In_834);
nor U1122 (N_1122,In_575,In_1578);
nor U1123 (N_1123,In_1722,In_1390);
xor U1124 (N_1124,In_807,In_2640);
nand U1125 (N_1125,In_1477,In_311);
nand U1126 (N_1126,In_2056,In_298);
nand U1127 (N_1127,In_2785,In_981);
xor U1128 (N_1128,In_197,In_1858);
nand U1129 (N_1129,In_2702,In_114);
nor U1130 (N_1130,In_2990,In_72);
nand U1131 (N_1131,In_2251,In_2484);
xnor U1132 (N_1132,In_157,In_2245);
nor U1133 (N_1133,In_11,In_1096);
and U1134 (N_1134,In_1526,In_1482);
xnor U1135 (N_1135,In_1560,In_1228);
and U1136 (N_1136,In_364,In_537);
xnor U1137 (N_1137,In_1705,In_2895);
nor U1138 (N_1138,In_2042,In_2577);
nor U1139 (N_1139,In_2182,In_2809);
nor U1140 (N_1140,In_325,In_2140);
or U1141 (N_1141,In_1842,In_2921);
or U1142 (N_1142,In_1193,In_2345);
nor U1143 (N_1143,In_2876,In_1177);
and U1144 (N_1144,In_858,In_1721);
nand U1145 (N_1145,In_1143,In_1523);
xor U1146 (N_1146,In_2836,In_1104);
and U1147 (N_1147,In_603,In_1406);
nor U1148 (N_1148,In_1015,In_857);
xnor U1149 (N_1149,In_1542,In_1227);
or U1150 (N_1150,In_2200,In_2961);
nor U1151 (N_1151,In_2256,In_2759);
or U1152 (N_1152,In_617,In_1408);
nand U1153 (N_1153,In_572,In_470);
xnor U1154 (N_1154,In_2027,In_284);
nor U1155 (N_1155,In_1281,In_482);
xnor U1156 (N_1156,In_367,In_2175);
nor U1157 (N_1157,In_1483,In_89);
nor U1158 (N_1158,In_1496,In_2423);
and U1159 (N_1159,In_137,In_1640);
nor U1160 (N_1160,In_2749,In_2538);
nor U1161 (N_1161,In_870,In_2289);
nor U1162 (N_1162,In_1052,In_1580);
or U1163 (N_1163,In_2786,In_2852);
and U1164 (N_1164,In_776,In_414);
xnor U1165 (N_1165,In_2839,In_1270);
or U1166 (N_1166,In_2769,In_781);
nand U1167 (N_1167,In_873,In_1181);
xnor U1168 (N_1168,In_2498,In_2024);
nor U1169 (N_1169,In_2522,In_2116);
nand U1170 (N_1170,In_1827,In_198);
xnor U1171 (N_1171,In_2904,In_2426);
or U1172 (N_1172,In_2033,In_1709);
and U1173 (N_1173,In_1987,In_1828);
and U1174 (N_1174,In_379,In_1697);
nand U1175 (N_1175,In_2948,In_75);
nor U1176 (N_1176,In_349,In_290);
nand U1177 (N_1177,In_1821,In_892);
nor U1178 (N_1178,In_1792,In_1222);
xor U1179 (N_1179,In_1627,In_714);
xor U1180 (N_1180,In_913,In_1165);
or U1181 (N_1181,In_1633,In_505);
and U1182 (N_1182,In_972,In_398);
nand U1183 (N_1183,In_1853,In_1402);
nor U1184 (N_1184,In_2187,In_509);
or U1185 (N_1185,In_86,In_2755);
nand U1186 (N_1186,In_1105,In_230);
nand U1187 (N_1187,In_1248,In_1068);
and U1188 (N_1188,In_1913,In_1290);
nor U1189 (N_1189,In_1257,In_1126);
xor U1190 (N_1190,In_2018,In_1844);
nand U1191 (N_1191,In_650,In_1550);
nor U1192 (N_1192,In_2457,In_856);
xnor U1193 (N_1193,In_1337,In_530);
xnor U1194 (N_1194,In_1345,In_2863);
or U1195 (N_1195,In_1907,In_1186);
xor U1196 (N_1196,In_2587,In_1767);
nand U1197 (N_1197,In_513,In_2098);
nor U1198 (N_1198,In_1776,In_1457);
xor U1199 (N_1199,In_2088,In_2872);
nor U1200 (N_1200,In_2906,In_1690);
nor U1201 (N_1201,In_2515,In_2189);
or U1202 (N_1202,In_1983,In_1091);
nor U1203 (N_1203,In_2879,In_844);
and U1204 (N_1204,In_2294,In_1447);
or U1205 (N_1205,In_1279,In_50);
and U1206 (N_1206,In_226,In_1537);
or U1207 (N_1207,In_2819,In_2941);
nor U1208 (N_1208,In_420,In_2646);
or U1209 (N_1209,In_1576,In_214);
nor U1210 (N_1210,In_909,In_631);
nand U1211 (N_1211,In_921,In_756);
nor U1212 (N_1212,In_2342,In_2077);
nor U1213 (N_1213,In_2316,In_210);
nor U1214 (N_1214,In_1723,In_32);
xor U1215 (N_1215,In_831,In_187);
nand U1216 (N_1216,In_1013,In_1745);
xnor U1217 (N_1217,In_1614,In_97);
xnor U1218 (N_1218,In_376,In_2456);
xnor U1219 (N_1219,In_720,In_729);
nand U1220 (N_1220,In_109,In_2873);
and U1221 (N_1221,In_1061,In_1955);
or U1222 (N_1222,In_1754,In_2346);
or U1223 (N_1223,In_217,In_1426);
xor U1224 (N_1224,In_1183,In_1783);
xnor U1225 (N_1225,In_2901,In_2475);
or U1226 (N_1226,In_1941,In_1107);
nor U1227 (N_1227,In_2142,In_498);
nor U1228 (N_1228,In_366,In_301);
or U1229 (N_1229,In_2350,In_320);
or U1230 (N_1230,In_923,In_1961);
and U1231 (N_1231,In_2417,In_2218);
or U1232 (N_1232,In_1643,In_1409);
and U1233 (N_1233,In_2845,In_2889);
or U1234 (N_1234,In_2435,In_246);
and U1235 (N_1235,In_2620,In_15);
nand U1236 (N_1236,In_2923,In_2746);
nand U1237 (N_1237,In_2802,In_2095);
nand U1238 (N_1238,In_1981,In_432);
and U1239 (N_1239,In_21,In_2579);
xnor U1240 (N_1240,In_2199,In_2291);
nor U1241 (N_1241,In_107,In_590);
xor U1242 (N_1242,In_2276,In_2013);
xnor U1243 (N_1243,In_1764,In_2530);
and U1244 (N_1244,In_2511,In_1158);
or U1245 (N_1245,In_2612,In_1166);
and U1246 (N_1246,In_1301,In_1873);
nor U1247 (N_1247,In_2455,In_286);
nand U1248 (N_1248,In_2776,In_916);
and U1249 (N_1249,In_2207,In_1586);
or U1250 (N_1250,In_960,In_1819);
or U1251 (N_1251,In_653,In_933);
nor U1252 (N_1252,In_3,In_1338);
or U1253 (N_1253,In_1051,In_1283);
nor U1254 (N_1254,In_2827,In_743);
nor U1255 (N_1255,In_1594,In_380);
xor U1256 (N_1256,In_649,In_1953);
nor U1257 (N_1257,In_148,In_2094);
or U1258 (N_1258,In_2369,In_1925);
and U1259 (N_1259,In_1260,In_2591);
xor U1260 (N_1260,In_1852,In_2002);
or U1261 (N_1261,In_1465,In_1976);
xor U1262 (N_1262,In_248,In_277);
or U1263 (N_1263,In_1349,In_953);
and U1264 (N_1264,In_57,In_1506);
nor U1265 (N_1265,In_2615,In_1243);
nor U1266 (N_1266,In_1430,In_2537);
xnor U1267 (N_1267,In_2566,In_2238);
nand U1268 (N_1268,In_2073,In_620);
nor U1269 (N_1269,In_2718,In_2050);
or U1270 (N_1270,In_2439,In_806);
nor U1271 (N_1271,In_2486,In_2740);
xor U1272 (N_1272,In_2750,In_2476);
nand U1273 (N_1273,In_1036,In_1136);
xnor U1274 (N_1274,In_2580,In_211);
xor U1275 (N_1275,In_908,In_144);
nor U1276 (N_1276,In_1401,In_2934);
nor U1277 (N_1277,In_2093,In_2334);
and U1278 (N_1278,In_1350,In_1011);
nand U1279 (N_1279,In_1249,In_58);
xor U1280 (N_1280,In_282,In_636);
or U1281 (N_1281,In_1493,In_2201);
xor U1282 (N_1282,In_800,In_1889);
xor U1283 (N_1283,In_1880,In_2214);
or U1284 (N_1284,In_105,In_2573);
nand U1285 (N_1285,In_1185,In_751);
xor U1286 (N_1286,In_2380,In_2383);
and U1287 (N_1287,In_891,In_1429);
nor U1288 (N_1288,In_989,In_540);
nor U1289 (N_1289,In_2909,In_1584);
xor U1290 (N_1290,In_371,In_1142);
nand U1291 (N_1291,In_1344,In_2023);
and U1292 (N_1292,In_842,In_218);
and U1293 (N_1293,In_1681,In_1942);
nor U1294 (N_1294,In_1018,In_1900);
xnor U1295 (N_1295,In_2359,In_2429);
xor U1296 (N_1296,In_2048,In_2596);
or U1297 (N_1297,In_1017,In_1785);
xor U1298 (N_1298,In_549,In_1891);
and U1299 (N_1299,In_854,In_627);
xor U1300 (N_1300,In_2575,In_2489);
or U1301 (N_1301,In_353,In_1569);
and U1302 (N_1302,In_597,In_63);
or U1303 (N_1303,In_1129,In_330);
xnor U1304 (N_1304,In_562,In_2588);
xor U1305 (N_1305,In_1850,In_2508);
nor U1306 (N_1306,In_769,In_1020);
xnor U1307 (N_1307,In_183,In_1871);
and U1308 (N_1308,In_1,In_2335);
or U1309 (N_1309,In_2170,In_2169);
and U1310 (N_1310,In_1851,In_1607);
and U1311 (N_1311,In_2460,In_1829);
nand U1312 (N_1312,In_1468,In_192);
nand U1313 (N_1313,In_103,In_1532);
xnor U1314 (N_1314,In_932,In_1934);
nand U1315 (N_1315,In_281,In_1514);
and U1316 (N_1316,In_2402,In_788);
and U1317 (N_1317,In_2131,In_98);
or U1318 (N_1318,In_2053,In_2471);
nor U1319 (N_1319,In_2519,In_664);
xnor U1320 (N_1320,In_1253,In_1841);
and U1321 (N_1321,In_42,In_1502);
nor U1322 (N_1322,In_828,In_2753);
nor U1323 (N_1323,In_747,In_948);
xnor U1324 (N_1324,In_958,In_336);
xor U1325 (N_1325,In_1089,In_2441);
nor U1326 (N_1326,In_883,In_324);
nand U1327 (N_1327,In_1768,In_1047);
nor U1328 (N_1328,In_1660,In_2679);
xor U1329 (N_1329,In_2495,In_1008);
xor U1330 (N_1330,In_680,In_1252);
and U1331 (N_1331,In_850,In_61);
and U1332 (N_1332,In_684,In_1310);
xor U1333 (N_1333,In_2083,In_1357);
or U1334 (N_1334,In_1678,In_2129);
or U1335 (N_1335,In_2706,In_1009);
xor U1336 (N_1336,In_1365,In_1039);
nor U1337 (N_1337,In_1410,In_2830);
nand U1338 (N_1338,In_1918,In_1149);
xor U1339 (N_1339,In_1817,In_536);
nand U1340 (N_1340,In_2803,In_2468);
nand U1341 (N_1341,In_2820,In_2158);
xor U1342 (N_1342,In_1176,In_158);
nor U1343 (N_1343,In_830,In_2057);
or U1344 (N_1344,In_1041,In_1777);
nor U1345 (N_1345,In_1035,In_2419);
and U1346 (N_1346,In_2210,In_1114);
xor U1347 (N_1347,In_999,In_577);
or U1348 (N_1348,In_186,In_1132);
nand U1349 (N_1349,In_2866,In_2309);
nor U1350 (N_1350,In_819,In_2265);
nor U1351 (N_1351,In_648,In_17);
and U1352 (N_1352,In_667,In_499);
nor U1353 (N_1353,In_2311,In_254);
nand U1354 (N_1354,In_901,In_544);
or U1355 (N_1355,In_1239,In_918);
and U1356 (N_1356,In_872,In_2502);
nand U1357 (N_1357,In_318,In_1534);
and U1358 (N_1358,In_768,In_1189);
nor U1359 (N_1359,In_496,In_2844);
or U1360 (N_1360,In_665,In_685);
and U1361 (N_1361,In_2997,In_2610);
nor U1362 (N_1362,In_1759,In_1480);
and U1363 (N_1363,In_1675,In_1210);
or U1364 (N_1364,In_2482,In_1170);
and U1365 (N_1365,In_786,In_129);
nor U1366 (N_1366,In_521,In_2594);
and U1367 (N_1367,In_2320,In_797);
or U1368 (N_1368,In_2186,In_2234);
or U1369 (N_1369,In_1874,In_1823);
or U1370 (N_1370,In_2274,In_142);
or U1371 (N_1371,In_1462,In_2688);
or U1372 (N_1372,In_464,In_1628);
and U1373 (N_1373,In_1152,In_2648);
nand U1374 (N_1374,In_2036,In_787);
xnor U1375 (N_1375,In_2968,In_2764);
nor U1376 (N_1376,In_1860,In_1090);
and U1377 (N_1377,In_1400,In_2026);
nor U1378 (N_1378,In_1905,In_2376);
nor U1379 (N_1379,In_2461,In_2561);
and U1380 (N_1380,In_327,In_1904);
or U1381 (N_1381,In_285,In_1229);
or U1382 (N_1382,In_1179,In_915);
and U1383 (N_1383,In_1590,In_232);
and U1384 (N_1384,In_875,In_559);
nor U1385 (N_1385,In_871,In_2752);
or U1386 (N_1386,In_2009,In_1173);
xnor U1387 (N_1387,In_2880,In_1269);
and U1388 (N_1388,In_2431,In_268);
nor U1389 (N_1389,In_698,In_30);
xor U1390 (N_1390,In_1508,In_252);
xor U1391 (N_1391,In_1672,In_2045);
xnor U1392 (N_1392,In_2965,In_1006);
nor U1393 (N_1393,In_511,In_2814);
nor U1394 (N_1394,In_2853,In_1236);
and U1395 (N_1395,In_2774,In_2491);
and U1396 (N_1396,In_1434,In_2373);
nand U1397 (N_1397,In_399,In_1683);
xor U1398 (N_1398,In_422,In_205);
nor U1399 (N_1399,In_1969,In_1748);
nor U1400 (N_1400,In_323,In_335);
xnor U1401 (N_1401,In_1323,In_2179);
or U1402 (N_1402,In_2939,In_2887);
nand U1403 (N_1403,In_122,In_2092);
nor U1404 (N_1404,In_321,In_1076);
nand U1405 (N_1405,In_1531,In_2885);
xor U1406 (N_1406,In_2211,In_1079);
nor U1407 (N_1407,In_2660,In_771);
xor U1408 (N_1408,In_2228,In_2970);
xor U1409 (N_1409,In_1028,In_2849);
or U1410 (N_1410,In_1911,In_1460);
nand U1411 (N_1411,In_2021,In_1049);
nand U1412 (N_1412,In_2821,In_384);
nor U1413 (N_1413,In_430,In_2699);
nor U1414 (N_1414,In_2076,In_1742);
nor U1415 (N_1415,In_1154,In_1991);
nand U1416 (N_1416,In_2514,In_1403);
nand U1417 (N_1417,In_867,In_332);
nand U1418 (N_1418,In_2817,In_288);
nor U1419 (N_1419,In_2313,In_2936);
and U1420 (N_1420,In_2552,In_1230);
and U1421 (N_1421,In_2004,In_2644);
or U1422 (N_1422,In_622,In_1634);
nand U1423 (N_1423,In_796,In_1398);
xnor U1424 (N_1424,In_1758,In_809);
nor U1425 (N_1425,In_1885,In_2950);
and U1426 (N_1426,In_2424,In_474);
nor U1427 (N_1427,In_938,In_2565);
xor U1428 (N_1428,In_906,In_1947);
xor U1429 (N_1429,In_1929,In_919);
nor U1430 (N_1430,In_1524,In_51);
nand U1431 (N_1431,In_503,In_1963);
xnor U1432 (N_1432,In_1630,In_2963);
nand U1433 (N_1433,In_1147,In_2855);
xnor U1434 (N_1434,In_2353,In_291);
nor U1435 (N_1435,In_1658,In_2540);
nor U1436 (N_1436,In_1064,In_1530);
nor U1437 (N_1437,In_2258,In_473);
nand U1438 (N_1438,In_1663,In_221);
or U1439 (N_1439,In_2477,In_1645);
or U1440 (N_1440,In_2133,In_1192);
or U1441 (N_1441,In_1644,In_2974);
nand U1442 (N_1442,In_260,In_1601);
nand U1443 (N_1443,In_346,In_2233);
nand U1444 (N_1444,In_2516,In_1159);
and U1445 (N_1445,In_1728,In_2452);
nand U1446 (N_1446,In_190,In_2499);
nand U1447 (N_1447,In_2937,In_1318);
and U1448 (N_1448,In_1361,In_132);
or U1449 (N_1449,In_1771,In_852);
or U1450 (N_1450,In_1000,In_2630);
xor U1451 (N_1451,In_2953,In_2795);
or U1452 (N_1452,In_1005,In_1689);
or U1453 (N_1453,In_2112,In_2996);
xnor U1454 (N_1454,In_2748,In_112);
and U1455 (N_1455,In_1386,In_1161);
xnor U1456 (N_1456,In_358,In_481);
nor U1457 (N_1457,In_113,In_545);
and U1458 (N_1458,In_979,In_1517);
and U1459 (N_1459,In_1613,In_1571);
or U1460 (N_1460,In_2006,In_1670);
and U1461 (N_1461,In_2085,In_2220);
xor U1462 (N_1462,In_861,In_108);
or U1463 (N_1463,In_227,In_1145);
nor U1464 (N_1464,In_1932,In_2842);
xnor U1465 (N_1465,In_946,In_1109);
nor U1466 (N_1466,In_2505,In_2574);
xor U1467 (N_1467,In_557,In_1704);
nor U1468 (N_1468,In_2292,In_351);
nand U1469 (N_1469,In_668,In_1048);
xnor U1470 (N_1470,In_2406,In_1866);
or U1471 (N_1471,In_341,In_692);
nand U1472 (N_1472,In_1691,In_2902);
or U1473 (N_1473,In_1377,In_1926);
nor U1474 (N_1474,In_1045,In_253);
and U1475 (N_1475,In_662,In_76);
nor U1476 (N_1476,In_2613,In_1080);
or U1477 (N_1477,In_2136,In_2315);
xnor U1478 (N_1478,In_2156,In_1615);
nand U1479 (N_1479,In_567,In_1044);
nor U1480 (N_1480,In_1024,In_306);
and U1481 (N_1481,In_2370,In_409);
nor U1482 (N_1482,In_2273,In_583);
nor U1483 (N_1483,In_1631,In_2008);
or U1484 (N_1484,In_2722,In_2944);
or U1485 (N_1485,In_1762,In_1624);
or U1486 (N_1486,In_1649,In_255);
xor U1487 (N_1487,In_2783,In_2727);
nor U1488 (N_1488,In_601,In_2387);
and U1489 (N_1489,In_2712,In_789);
nand U1490 (N_1490,In_886,In_2556);
and U1491 (N_1491,In_639,In_1933);
nor U1492 (N_1492,In_1397,In_104);
and U1493 (N_1493,In_997,In_2385);
nor U1494 (N_1494,In_820,In_2645);
and U1495 (N_1495,In_2656,In_1328);
nor U1496 (N_1496,In_184,In_344);
nand U1497 (N_1497,In_53,In_1862);
nor U1498 (N_1498,In_1412,In_1755);
or U1499 (N_1499,In_413,In_1952);
xnor U1500 (N_1500,In_2673,In_2451);
nand U1501 (N_1501,In_1767,In_385);
nand U1502 (N_1502,In_1521,In_2810);
nand U1503 (N_1503,In_2452,In_1873);
nor U1504 (N_1504,In_1890,In_1106);
nand U1505 (N_1505,In_1617,In_1982);
and U1506 (N_1506,In_16,In_2864);
or U1507 (N_1507,In_1249,In_2089);
and U1508 (N_1508,In_571,In_1202);
or U1509 (N_1509,In_428,In_103);
nand U1510 (N_1510,In_592,In_1780);
xor U1511 (N_1511,In_401,In_121);
nand U1512 (N_1512,In_1636,In_1916);
nand U1513 (N_1513,In_2189,In_2906);
nand U1514 (N_1514,In_1145,In_1150);
or U1515 (N_1515,In_696,In_1458);
nand U1516 (N_1516,In_2930,In_1655);
xor U1517 (N_1517,In_565,In_2);
or U1518 (N_1518,In_1654,In_1062);
nor U1519 (N_1519,In_2272,In_861);
nand U1520 (N_1520,In_2620,In_1209);
nand U1521 (N_1521,In_27,In_256);
and U1522 (N_1522,In_353,In_1387);
xnor U1523 (N_1523,In_290,In_1111);
xor U1524 (N_1524,In_1694,In_124);
nor U1525 (N_1525,In_952,In_2742);
and U1526 (N_1526,In_2167,In_1527);
nor U1527 (N_1527,In_1777,In_1065);
xnor U1528 (N_1528,In_2100,In_614);
xnor U1529 (N_1529,In_2765,In_303);
and U1530 (N_1530,In_2496,In_1336);
nor U1531 (N_1531,In_2743,In_347);
and U1532 (N_1532,In_1400,In_1573);
or U1533 (N_1533,In_1770,In_1252);
nor U1534 (N_1534,In_844,In_2197);
nor U1535 (N_1535,In_1275,In_797);
or U1536 (N_1536,In_1748,In_496);
and U1537 (N_1537,In_1077,In_1640);
xor U1538 (N_1538,In_2518,In_1948);
nor U1539 (N_1539,In_2937,In_832);
or U1540 (N_1540,In_563,In_1036);
xnor U1541 (N_1541,In_2668,In_107);
and U1542 (N_1542,In_966,In_2677);
nor U1543 (N_1543,In_1034,In_2968);
or U1544 (N_1544,In_2049,In_1379);
nand U1545 (N_1545,In_608,In_2160);
nand U1546 (N_1546,In_1838,In_605);
nor U1547 (N_1547,In_2488,In_777);
nand U1548 (N_1548,In_398,In_838);
nor U1549 (N_1549,In_1924,In_397);
and U1550 (N_1550,In_2575,In_2615);
or U1551 (N_1551,In_145,In_2640);
xnor U1552 (N_1552,In_2193,In_411);
nor U1553 (N_1553,In_692,In_2668);
nand U1554 (N_1554,In_1045,In_2866);
and U1555 (N_1555,In_364,In_237);
or U1556 (N_1556,In_1724,In_590);
nor U1557 (N_1557,In_478,In_1798);
or U1558 (N_1558,In_983,In_2456);
nand U1559 (N_1559,In_805,In_2834);
and U1560 (N_1560,In_1326,In_1879);
nand U1561 (N_1561,In_2299,In_1634);
nand U1562 (N_1562,In_1369,In_2467);
nand U1563 (N_1563,In_645,In_1110);
nor U1564 (N_1564,In_2165,In_2571);
or U1565 (N_1565,In_1,In_904);
and U1566 (N_1566,In_684,In_2173);
and U1567 (N_1567,In_2974,In_599);
xor U1568 (N_1568,In_2016,In_2178);
nand U1569 (N_1569,In_986,In_2837);
nand U1570 (N_1570,In_870,In_1213);
nor U1571 (N_1571,In_2950,In_1735);
xor U1572 (N_1572,In_1339,In_312);
and U1573 (N_1573,In_1434,In_562);
and U1574 (N_1574,In_485,In_363);
or U1575 (N_1575,In_2720,In_2288);
nor U1576 (N_1576,In_1466,In_1293);
nor U1577 (N_1577,In_2549,In_903);
nand U1578 (N_1578,In_628,In_2039);
nand U1579 (N_1579,In_1705,In_2859);
nor U1580 (N_1580,In_1090,In_370);
xnor U1581 (N_1581,In_1991,In_2476);
or U1582 (N_1582,In_1710,In_2610);
nand U1583 (N_1583,In_34,In_2819);
and U1584 (N_1584,In_1844,In_597);
or U1585 (N_1585,In_1290,In_187);
nor U1586 (N_1586,In_458,In_1346);
nand U1587 (N_1587,In_360,In_2635);
and U1588 (N_1588,In_2105,In_407);
or U1589 (N_1589,In_2301,In_2855);
and U1590 (N_1590,In_2015,In_1512);
and U1591 (N_1591,In_2758,In_792);
nor U1592 (N_1592,In_558,In_1896);
or U1593 (N_1593,In_2007,In_150);
and U1594 (N_1594,In_2198,In_1136);
nand U1595 (N_1595,In_447,In_2618);
nor U1596 (N_1596,In_2652,In_277);
xor U1597 (N_1597,In_1238,In_1313);
nand U1598 (N_1598,In_460,In_2994);
nand U1599 (N_1599,In_1540,In_2208);
nor U1600 (N_1600,In_807,In_1818);
and U1601 (N_1601,In_1664,In_1603);
and U1602 (N_1602,In_409,In_2210);
nand U1603 (N_1603,In_2519,In_449);
or U1604 (N_1604,In_42,In_765);
nand U1605 (N_1605,In_2948,In_2142);
or U1606 (N_1606,In_1201,In_254);
nor U1607 (N_1607,In_67,In_2311);
and U1608 (N_1608,In_1875,In_589);
and U1609 (N_1609,In_2793,In_923);
nor U1610 (N_1610,In_1180,In_1338);
nor U1611 (N_1611,In_489,In_2682);
and U1612 (N_1612,In_1256,In_1007);
xor U1613 (N_1613,In_598,In_2540);
xnor U1614 (N_1614,In_923,In_759);
nor U1615 (N_1615,In_2367,In_2986);
xnor U1616 (N_1616,In_890,In_335);
nand U1617 (N_1617,In_937,In_193);
or U1618 (N_1618,In_1611,In_584);
nor U1619 (N_1619,In_209,In_444);
nor U1620 (N_1620,In_118,In_2196);
or U1621 (N_1621,In_1257,In_2520);
or U1622 (N_1622,In_2714,In_1106);
or U1623 (N_1623,In_1438,In_2833);
xnor U1624 (N_1624,In_1724,In_794);
or U1625 (N_1625,In_1154,In_127);
and U1626 (N_1626,In_1116,In_1465);
or U1627 (N_1627,In_637,In_2358);
and U1628 (N_1628,In_2193,In_1467);
nand U1629 (N_1629,In_314,In_1990);
or U1630 (N_1630,In_533,In_2855);
nand U1631 (N_1631,In_1297,In_565);
nand U1632 (N_1632,In_942,In_2567);
xor U1633 (N_1633,In_143,In_2400);
and U1634 (N_1634,In_468,In_2311);
or U1635 (N_1635,In_1980,In_2933);
nor U1636 (N_1636,In_444,In_956);
nor U1637 (N_1637,In_2658,In_669);
and U1638 (N_1638,In_982,In_2666);
and U1639 (N_1639,In_945,In_2166);
xor U1640 (N_1640,In_883,In_2808);
and U1641 (N_1641,In_1515,In_495);
and U1642 (N_1642,In_836,In_1448);
and U1643 (N_1643,In_651,In_2045);
or U1644 (N_1644,In_470,In_1912);
nand U1645 (N_1645,In_297,In_1261);
and U1646 (N_1646,In_2268,In_533);
or U1647 (N_1647,In_722,In_1497);
xor U1648 (N_1648,In_1618,In_754);
or U1649 (N_1649,In_1723,In_2036);
nor U1650 (N_1650,In_2113,In_1894);
nand U1651 (N_1651,In_1921,In_1901);
nand U1652 (N_1652,In_921,In_994);
nand U1653 (N_1653,In_904,In_2856);
xnor U1654 (N_1654,In_1497,In_2261);
and U1655 (N_1655,In_1341,In_233);
xor U1656 (N_1656,In_1975,In_2144);
nor U1657 (N_1657,In_1221,In_1070);
nand U1658 (N_1658,In_2859,In_757);
xor U1659 (N_1659,In_2773,In_1037);
or U1660 (N_1660,In_1701,In_1043);
xnor U1661 (N_1661,In_2363,In_1104);
xor U1662 (N_1662,In_463,In_546);
nor U1663 (N_1663,In_626,In_966);
xnor U1664 (N_1664,In_334,In_1026);
nor U1665 (N_1665,In_2466,In_2221);
or U1666 (N_1666,In_2496,In_1941);
and U1667 (N_1667,In_1861,In_1142);
nor U1668 (N_1668,In_1971,In_2224);
xnor U1669 (N_1669,In_2837,In_1218);
xnor U1670 (N_1670,In_733,In_2414);
nand U1671 (N_1671,In_1377,In_2301);
or U1672 (N_1672,In_1584,In_2461);
nor U1673 (N_1673,In_2740,In_2756);
and U1674 (N_1674,In_2601,In_2823);
nor U1675 (N_1675,In_353,In_1126);
or U1676 (N_1676,In_1249,In_2991);
or U1677 (N_1677,In_2935,In_1514);
nor U1678 (N_1678,In_2092,In_1918);
and U1679 (N_1679,In_565,In_2756);
nor U1680 (N_1680,In_2883,In_987);
or U1681 (N_1681,In_730,In_919);
and U1682 (N_1682,In_1161,In_2585);
nand U1683 (N_1683,In_1430,In_2777);
nand U1684 (N_1684,In_1547,In_2629);
xor U1685 (N_1685,In_1172,In_1294);
or U1686 (N_1686,In_2371,In_1977);
or U1687 (N_1687,In_1341,In_1893);
xor U1688 (N_1688,In_1398,In_116);
xnor U1689 (N_1689,In_2579,In_436);
and U1690 (N_1690,In_729,In_1204);
and U1691 (N_1691,In_1442,In_556);
and U1692 (N_1692,In_2026,In_647);
nor U1693 (N_1693,In_996,In_1380);
xnor U1694 (N_1694,In_1061,In_1682);
or U1695 (N_1695,In_2597,In_967);
nor U1696 (N_1696,In_133,In_2840);
and U1697 (N_1697,In_1341,In_45);
and U1698 (N_1698,In_989,In_390);
xnor U1699 (N_1699,In_1856,In_1970);
xor U1700 (N_1700,In_2476,In_160);
or U1701 (N_1701,In_2785,In_313);
or U1702 (N_1702,In_684,In_1155);
nand U1703 (N_1703,In_2829,In_1654);
or U1704 (N_1704,In_2933,In_2337);
nand U1705 (N_1705,In_2990,In_283);
or U1706 (N_1706,In_2815,In_2867);
xor U1707 (N_1707,In_35,In_1412);
and U1708 (N_1708,In_1316,In_2015);
nor U1709 (N_1709,In_2373,In_1022);
nand U1710 (N_1710,In_1723,In_645);
and U1711 (N_1711,In_576,In_1373);
nand U1712 (N_1712,In_1372,In_210);
nand U1713 (N_1713,In_1925,In_610);
nor U1714 (N_1714,In_163,In_2877);
or U1715 (N_1715,In_594,In_1121);
nor U1716 (N_1716,In_1272,In_2372);
or U1717 (N_1717,In_986,In_439);
nor U1718 (N_1718,In_2279,In_815);
nand U1719 (N_1719,In_2902,In_1634);
and U1720 (N_1720,In_1114,In_2305);
nor U1721 (N_1721,In_2208,In_1182);
and U1722 (N_1722,In_680,In_922);
or U1723 (N_1723,In_2028,In_591);
and U1724 (N_1724,In_2478,In_254);
nor U1725 (N_1725,In_55,In_2744);
xor U1726 (N_1726,In_1747,In_2467);
nor U1727 (N_1727,In_1985,In_446);
nand U1728 (N_1728,In_1235,In_404);
nor U1729 (N_1729,In_1364,In_784);
xnor U1730 (N_1730,In_152,In_1670);
nand U1731 (N_1731,In_1114,In_1506);
or U1732 (N_1732,In_138,In_2314);
nor U1733 (N_1733,In_493,In_1979);
or U1734 (N_1734,In_2526,In_1338);
xnor U1735 (N_1735,In_390,In_1189);
and U1736 (N_1736,In_210,In_1337);
or U1737 (N_1737,In_60,In_1245);
nand U1738 (N_1738,In_349,In_1536);
or U1739 (N_1739,In_33,In_2756);
or U1740 (N_1740,In_2713,In_1572);
and U1741 (N_1741,In_228,In_511);
or U1742 (N_1742,In_2645,In_2502);
and U1743 (N_1743,In_726,In_2609);
xnor U1744 (N_1744,In_82,In_1980);
or U1745 (N_1745,In_2019,In_669);
xor U1746 (N_1746,In_2797,In_1572);
or U1747 (N_1747,In_1940,In_628);
xor U1748 (N_1748,In_1360,In_2626);
nor U1749 (N_1749,In_1542,In_2848);
nand U1750 (N_1750,In_2227,In_712);
or U1751 (N_1751,In_1997,In_1277);
or U1752 (N_1752,In_1158,In_577);
nor U1753 (N_1753,In_2132,In_2688);
xnor U1754 (N_1754,In_2363,In_2429);
nor U1755 (N_1755,In_781,In_2864);
or U1756 (N_1756,In_2434,In_541);
nor U1757 (N_1757,In_2668,In_1158);
and U1758 (N_1758,In_2398,In_2819);
and U1759 (N_1759,In_2119,In_849);
or U1760 (N_1760,In_2898,In_1483);
nand U1761 (N_1761,In_1863,In_1804);
nand U1762 (N_1762,In_1141,In_1922);
xor U1763 (N_1763,In_1869,In_1353);
nor U1764 (N_1764,In_2848,In_1214);
nand U1765 (N_1765,In_2928,In_755);
nand U1766 (N_1766,In_869,In_2335);
xnor U1767 (N_1767,In_2849,In_1336);
xor U1768 (N_1768,In_2113,In_1078);
xnor U1769 (N_1769,In_1631,In_1054);
nor U1770 (N_1770,In_1257,In_499);
or U1771 (N_1771,In_2534,In_1710);
nand U1772 (N_1772,In_738,In_1628);
nor U1773 (N_1773,In_476,In_1798);
and U1774 (N_1774,In_1118,In_2205);
xor U1775 (N_1775,In_1969,In_151);
nand U1776 (N_1776,In_763,In_2166);
nor U1777 (N_1777,In_1973,In_2610);
xor U1778 (N_1778,In_683,In_2437);
xnor U1779 (N_1779,In_1035,In_1960);
xnor U1780 (N_1780,In_2876,In_1638);
nand U1781 (N_1781,In_446,In_267);
nand U1782 (N_1782,In_1344,In_1746);
nor U1783 (N_1783,In_1564,In_1020);
nor U1784 (N_1784,In_2295,In_762);
xnor U1785 (N_1785,In_1412,In_2527);
nor U1786 (N_1786,In_2786,In_2316);
nor U1787 (N_1787,In_2323,In_1362);
and U1788 (N_1788,In_1249,In_1032);
xnor U1789 (N_1789,In_2910,In_29);
nor U1790 (N_1790,In_2071,In_178);
nand U1791 (N_1791,In_1575,In_1124);
nand U1792 (N_1792,In_2991,In_2971);
and U1793 (N_1793,In_2116,In_2817);
and U1794 (N_1794,In_1026,In_2014);
nor U1795 (N_1795,In_288,In_2025);
xor U1796 (N_1796,In_21,In_1906);
xor U1797 (N_1797,In_1755,In_699);
nand U1798 (N_1798,In_808,In_2086);
and U1799 (N_1799,In_824,In_2712);
xnor U1800 (N_1800,In_2132,In_579);
xnor U1801 (N_1801,In_1790,In_164);
xor U1802 (N_1802,In_1959,In_344);
nor U1803 (N_1803,In_878,In_2436);
and U1804 (N_1804,In_878,In_582);
or U1805 (N_1805,In_2577,In_1099);
nor U1806 (N_1806,In_1064,In_2473);
and U1807 (N_1807,In_380,In_586);
xnor U1808 (N_1808,In_1929,In_2315);
nor U1809 (N_1809,In_886,In_1576);
nor U1810 (N_1810,In_1099,In_1467);
xor U1811 (N_1811,In_1795,In_1048);
and U1812 (N_1812,In_2316,In_1710);
nand U1813 (N_1813,In_248,In_1066);
nor U1814 (N_1814,In_341,In_1271);
nand U1815 (N_1815,In_1926,In_954);
nand U1816 (N_1816,In_2951,In_19);
xor U1817 (N_1817,In_2090,In_700);
and U1818 (N_1818,In_2669,In_1026);
xnor U1819 (N_1819,In_930,In_1775);
or U1820 (N_1820,In_237,In_1177);
or U1821 (N_1821,In_2274,In_1176);
or U1822 (N_1822,In_2964,In_1299);
or U1823 (N_1823,In_1884,In_248);
nand U1824 (N_1824,In_580,In_652);
xor U1825 (N_1825,In_444,In_825);
nor U1826 (N_1826,In_2258,In_2410);
nor U1827 (N_1827,In_563,In_2652);
xor U1828 (N_1828,In_2130,In_2958);
nor U1829 (N_1829,In_346,In_2708);
and U1830 (N_1830,In_897,In_2914);
nor U1831 (N_1831,In_274,In_65);
xnor U1832 (N_1832,In_2959,In_70);
and U1833 (N_1833,In_2923,In_2197);
nor U1834 (N_1834,In_1250,In_157);
nand U1835 (N_1835,In_1545,In_650);
or U1836 (N_1836,In_906,In_1501);
nand U1837 (N_1837,In_2250,In_101);
or U1838 (N_1838,In_2387,In_2099);
xor U1839 (N_1839,In_717,In_665);
nor U1840 (N_1840,In_1830,In_826);
nand U1841 (N_1841,In_2167,In_2532);
and U1842 (N_1842,In_2601,In_1449);
xor U1843 (N_1843,In_409,In_2076);
or U1844 (N_1844,In_1974,In_1844);
nor U1845 (N_1845,In_616,In_1948);
nand U1846 (N_1846,In_1084,In_78);
nand U1847 (N_1847,In_500,In_1936);
nor U1848 (N_1848,In_713,In_2758);
xor U1849 (N_1849,In_1296,In_254);
nand U1850 (N_1850,In_2100,In_900);
and U1851 (N_1851,In_2696,In_2608);
nor U1852 (N_1852,In_1565,In_1836);
xnor U1853 (N_1853,In_2142,In_290);
and U1854 (N_1854,In_738,In_1543);
nor U1855 (N_1855,In_756,In_1416);
and U1856 (N_1856,In_2187,In_1289);
or U1857 (N_1857,In_1340,In_1158);
and U1858 (N_1858,In_1683,In_2520);
and U1859 (N_1859,In_9,In_800);
xnor U1860 (N_1860,In_1794,In_35);
nor U1861 (N_1861,In_486,In_662);
and U1862 (N_1862,In_2314,In_2219);
nand U1863 (N_1863,In_1144,In_1254);
nand U1864 (N_1864,In_1300,In_1261);
nor U1865 (N_1865,In_640,In_845);
xnor U1866 (N_1866,In_2218,In_2206);
xnor U1867 (N_1867,In_2675,In_2310);
xor U1868 (N_1868,In_1395,In_846);
nand U1869 (N_1869,In_1635,In_2205);
xnor U1870 (N_1870,In_2206,In_2397);
or U1871 (N_1871,In_1014,In_2812);
or U1872 (N_1872,In_1586,In_2816);
nor U1873 (N_1873,In_683,In_1105);
or U1874 (N_1874,In_2900,In_2678);
nand U1875 (N_1875,In_1117,In_1124);
or U1876 (N_1876,In_2828,In_1351);
and U1877 (N_1877,In_1463,In_1644);
nand U1878 (N_1878,In_200,In_2441);
nand U1879 (N_1879,In_2172,In_1261);
and U1880 (N_1880,In_694,In_289);
nor U1881 (N_1881,In_1294,In_1833);
or U1882 (N_1882,In_298,In_1646);
or U1883 (N_1883,In_1163,In_1302);
nor U1884 (N_1884,In_1583,In_1580);
or U1885 (N_1885,In_2280,In_2571);
nand U1886 (N_1886,In_1709,In_2068);
nor U1887 (N_1887,In_995,In_868);
and U1888 (N_1888,In_345,In_296);
and U1889 (N_1889,In_1468,In_1879);
xnor U1890 (N_1890,In_2728,In_1007);
and U1891 (N_1891,In_2534,In_1068);
and U1892 (N_1892,In_2287,In_2561);
or U1893 (N_1893,In_1943,In_2215);
nor U1894 (N_1894,In_86,In_1298);
xnor U1895 (N_1895,In_2359,In_2719);
nand U1896 (N_1896,In_2237,In_2393);
xnor U1897 (N_1897,In_869,In_1360);
xor U1898 (N_1898,In_2408,In_2480);
xnor U1899 (N_1899,In_1864,In_1115);
nand U1900 (N_1900,In_708,In_2260);
xnor U1901 (N_1901,In_2089,In_729);
nor U1902 (N_1902,In_337,In_610);
and U1903 (N_1903,In_1392,In_456);
or U1904 (N_1904,In_2227,In_2311);
xor U1905 (N_1905,In_560,In_804);
nand U1906 (N_1906,In_1643,In_895);
nand U1907 (N_1907,In_872,In_1391);
or U1908 (N_1908,In_1141,In_2822);
and U1909 (N_1909,In_885,In_1274);
nand U1910 (N_1910,In_1413,In_1529);
nor U1911 (N_1911,In_891,In_2608);
and U1912 (N_1912,In_1257,In_677);
or U1913 (N_1913,In_1399,In_2098);
xor U1914 (N_1914,In_723,In_1425);
nand U1915 (N_1915,In_2350,In_2268);
nor U1916 (N_1916,In_2881,In_446);
or U1917 (N_1917,In_2846,In_2035);
nor U1918 (N_1918,In_2032,In_1268);
nand U1919 (N_1919,In_1974,In_786);
and U1920 (N_1920,In_628,In_2195);
nor U1921 (N_1921,In_1673,In_1620);
xnor U1922 (N_1922,In_481,In_1113);
nand U1923 (N_1923,In_2932,In_1031);
and U1924 (N_1924,In_1725,In_952);
and U1925 (N_1925,In_675,In_902);
xor U1926 (N_1926,In_1502,In_1258);
nand U1927 (N_1927,In_2795,In_1372);
xnor U1928 (N_1928,In_293,In_1821);
nor U1929 (N_1929,In_1545,In_2449);
nand U1930 (N_1930,In_1481,In_1602);
xor U1931 (N_1931,In_841,In_683);
or U1932 (N_1932,In_1120,In_2442);
and U1933 (N_1933,In_805,In_161);
nor U1934 (N_1934,In_1979,In_1790);
nand U1935 (N_1935,In_2442,In_1983);
xor U1936 (N_1936,In_768,In_283);
or U1937 (N_1937,In_1017,In_2176);
xor U1938 (N_1938,In_147,In_1466);
nand U1939 (N_1939,In_49,In_144);
xor U1940 (N_1940,In_1306,In_2806);
or U1941 (N_1941,In_2871,In_816);
xnor U1942 (N_1942,In_1811,In_208);
xor U1943 (N_1943,In_610,In_2668);
nand U1944 (N_1944,In_904,In_91);
nand U1945 (N_1945,In_2869,In_855);
xnor U1946 (N_1946,In_2963,In_126);
and U1947 (N_1947,In_681,In_1901);
nand U1948 (N_1948,In_1517,In_820);
xor U1949 (N_1949,In_896,In_530);
nand U1950 (N_1950,In_2551,In_2358);
nor U1951 (N_1951,In_2300,In_1307);
nor U1952 (N_1952,In_1849,In_863);
xnor U1953 (N_1953,In_360,In_348);
nor U1954 (N_1954,In_575,In_2519);
nor U1955 (N_1955,In_42,In_2836);
nor U1956 (N_1956,In_815,In_1709);
or U1957 (N_1957,In_1998,In_2190);
or U1958 (N_1958,In_225,In_39);
nor U1959 (N_1959,In_2734,In_2910);
xnor U1960 (N_1960,In_2026,In_2037);
and U1961 (N_1961,In_1967,In_1879);
and U1962 (N_1962,In_2083,In_2682);
xnor U1963 (N_1963,In_2524,In_928);
or U1964 (N_1964,In_1927,In_368);
xor U1965 (N_1965,In_1715,In_1155);
xnor U1966 (N_1966,In_2450,In_1611);
or U1967 (N_1967,In_845,In_433);
xnor U1968 (N_1968,In_2738,In_2448);
nor U1969 (N_1969,In_951,In_1604);
xnor U1970 (N_1970,In_421,In_1773);
and U1971 (N_1971,In_1291,In_884);
nand U1972 (N_1972,In_682,In_1579);
nor U1973 (N_1973,In_1280,In_731);
nor U1974 (N_1974,In_2167,In_2673);
and U1975 (N_1975,In_447,In_1914);
xor U1976 (N_1976,In_1160,In_260);
and U1977 (N_1977,In_670,In_2310);
and U1978 (N_1978,In_2499,In_1944);
or U1979 (N_1979,In_2437,In_1276);
or U1980 (N_1980,In_2893,In_1730);
xor U1981 (N_1981,In_1366,In_2912);
nor U1982 (N_1982,In_587,In_1316);
and U1983 (N_1983,In_1518,In_1961);
nand U1984 (N_1984,In_1012,In_96);
and U1985 (N_1985,In_2724,In_316);
or U1986 (N_1986,In_2809,In_1339);
xnor U1987 (N_1987,In_2782,In_917);
nand U1988 (N_1988,In_2120,In_1382);
nor U1989 (N_1989,In_2526,In_1098);
or U1990 (N_1990,In_1122,In_2666);
and U1991 (N_1991,In_943,In_2425);
xnor U1992 (N_1992,In_575,In_1917);
nor U1993 (N_1993,In_79,In_2152);
nand U1994 (N_1994,In_1531,In_2322);
and U1995 (N_1995,In_412,In_298);
xnor U1996 (N_1996,In_2374,In_1064);
xnor U1997 (N_1997,In_1414,In_2180);
nor U1998 (N_1998,In_2657,In_1936);
or U1999 (N_1999,In_1474,In_2833);
and U2000 (N_2000,In_2044,In_1029);
nor U2001 (N_2001,In_2095,In_764);
or U2002 (N_2002,In_482,In_1749);
nand U2003 (N_2003,In_1700,In_592);
and U2004 (N_2004,In_85,In_2079);
or U2005 (N_2005,In_996,In_1175);
nand U2006 (N_2006,In_624,In_1595);
xnor U2007 (N_2007,In_1893,In_1364);
nor U2008 (N_2008,In_643,In_1818);
or U2009 (N_2009,In_1444,In_910);
or U2010 (N_2010,In_2021,In_1186);
xnor U2011 (N_2011,In_2964,In_863);
nor U2012 (N_2012,In_2082,In_1135);
xnor U2013 (N_2013,In_2104,In_910);
nor U2014 (N_2014,In_1833,In_697);
nor U2015 (N_2015,In_1440,In_992);
or U2016 (N_2016,In_1518,In_1846);
nand U2017 (N_2017,In_1785,In_963);
and U2018 (N_2018,In_233,In_2314);
and U2019 (N_2019,In_197,In_1464);
or U2020 (N_2020,In_2729,In_1408);
nor U2021 (N_2021,In_2943,In_1444);
or U2022 (N_2022,In_1659,In_1730);
and U2023 (N_2023,In_2511,In_1393);
nor U2024 (N_2024,In_2210,In_1540);
and U2025 (N_2025,In_99,In_4);
and U2026 (N_2026,In_2337,In_594);
and U2027 (N_2027,In_329,In_1040);
xor U2028 (N_2028,In_548,In_2456);
xnor U2029 (N_2029,In_2780,In_2269);
nor U2030 (N_2030,In_2500,In_2649);
xor U2031 (N_2031,In_475,In_1713);
xor U2032 (N_2032,In_2143,In_1588);
and U2033 (N_2033,In_1961,In_1630);
or U2034 (N_2034,In_2388,In_917);
nand U2035 (N_2035,In_1492,In_50);
nand U2036 (N_2036,In_2172,In_1177);
nor U2037 (N_2037,In_2337,In_2905);
or U2038 (N_2038,In_1241,In_294);
nand U2039 (N_2039,In_1557,In_2974);
xnor U2040 (N_2040,In_2254,In_1612);
nor U2041 (N_2041,In_2335,In_668);
and U2042 (N_2042,In_1244,In_1441);
or U2043 (N_2043,In_1888,In_2296);
nand U2044 (N_2044,In_1075,In_2369);
nand U2045 (N_2045,In_880,In_1669);
or U2046 (N_2046,In_554,In_2927);
and U2047 (N_2047,In_70,In_2137);
nand U2048 (N_2048,In_754,In_750);
nand U2049 (N_2049,In_1532,In_2394);
and U2050 (N_2050,In_182,In_2233);
and U2051 (N_2051,In_88,In_1112);
or U2052 (N_2052,In_186,In_2590);
and U2053 (N_2053,In_765,In_525);
nor U2054 (N_2054,In_256,In_2495);
xor U2055 (N_2055,In_2256,In_2444);
or U2056 (N_2056,In_783,In_996);
xnor U2057 (N_2057,In_487,In_2754);
and U2058 (N_2058,In_2643,In_1855);
nor U2059 (N_2059,In_1965,In_1763);
nor U2060 (N_2060,In_71,In_2267);
and U2061 (N_2061,In_2373,In_2173);
nand U2062 (N_2062,In_1113,In_1294);
or U2063 (N_2063,In_362,In_2523);
and U2064 (N_2064,In_2844,In_1451);
nor U2065 (N_2065,In_2022,In_1811);
or U2066 (N_2066,In_715,In_1691);
or U2067 (N_2067,In_2208,In_1014);
nand U2068 (N_2068,In_107,In_914);
xnor U2069 (N_2069,In_2256,In_1374);
nand U2070 (N_2070,In_2231,In_809);
xnor U2071 (N_2071,In_2849,In_1842);
nand U2072 (N_2072,In_912,In_245);
or U2073 (N_2073,In_2966,In_1596);
xor U2074 (N_2074,In_166,In_1813);
nor U2075 (N_2075,In_683,In_89);
nand U2076 (N_2076,In_1115,In_2565);
xnor U2077 (N_2077,In_823,In_58);
nor U2078 (N_2078,In_2838,In_2631);
or U2079 (N_2079,In_2574,In_355);
xor U2080 (N_2080,In_736,In_1566);
and U2081 (N_2081,In_798,In_566);
or U2082 (N_2082,In_2335,In_1266);
nor U2083 (N_2083,In_453,In_728);
or U2084 (N_2084,In_2855,In_2515);
xor U2085 (N_2085,In_149,In_352);
and U2086 (N_2086,In_238,In_2687);
or U2087 (N_2087,In_872,In_2295);
nand U2088 (N_2088,In_70,In_2733);
or U2089 (N_2089,In_1190,In_1832);
and U2090 (N_2090,In_1413,In_1965);
or U2091 (N_2091,In_2954,In_93);
nand U2092 (N_2092,In_195,In_546);
nor U2093 (N_2093,In_628,In_993);
or U2094 (N_2094,In_1145,In_193);
nand U2095 (N_2095,In_2896,In_1660);
nor U2096 (N_2096,In_2949,In_2448);
xor U2097 (N_2097,In_2595,In_1176);
and U2098 (N_2098,In_208,In_589);
xor U2099 (N_2099,In_1639,In_230);
nand U2100 (N_2100,In_501,In_2073);
or U2101 (N_2101,In_2058,In_436);
and U2102 (N_2102,In_298,In_1560);
or U2103 (N_2103,In_2003,In_2860);
and U2104 (N_2104,In_2646,In_862);
nand U2105 (N_2105,In_1293,In_1532);
nor U2106 (N_2106,In_104,In_142);
nand U2107 (N_2107,In_2958,In_1248);
or U2108 (N_2108,In_2277,In_1491);
xor U2109 (N_2109,In_1229,In_1177);
nor U2110 (N_2110,In_2191,In_2738);
nand U2111 (N_2111,In_1542,In_137);
nor U2112 (N_2112,In_2217,In_2341);
nand U2113 (N_2113,In_245,In_2657);
nand U2114 (N_2114,In_264,In_416);
xnor U2115 (N_2115,In_1749,In_1450);
xnor U2116 (N_2116,In_178,In_110);
and U2117 (N_2117,In_787,In_1223);
nand U2118 (N_2118,In_172,In_2902);
nand U2119 (N_2119,In_290,In_738);
xor U2120 (N_2120,In_2508,In_1253);
nand U2121 (N_2121,In_197,In_1897);
xor U2122 (N_2122,In_2848,In_2266);
or U2123 (N_2123,In_1410,In_996);
nor U2124 (N_2124,In_2359,In_1847);
or U2125 (N_2125,In_2711,In_2703);
nand U2126 (N_2126,In_394,In_2504);
nor U2127 (N_2127,In_2426,In_2645);
or U2128 (N_2128,In_1128,In_2175);
or U2129 (N_2129,In_2136,In_645);
and U2130 (N_2130,In_1646,In_2716);
and U2131 (N_2131,In_139,In_1983);
and U2132 (N_2132,In_1435,In_1663);
nand U2133 (N_2133,In_1316,In_1883);
nand U2134 (N_2134,In_1993,In_1528);
and U2135 (N_2135,In_2674,In_106);
and U2136 (N_2136,In_2900,In_2687);
or U2137 (N_2137,In_979,In_456);
nand U2138 (N_2138,In_659,In_807);
nand U2139 (N_2139,In_2744,In_2069);
xor U2140 (N_2140,In_2896,In_1488);
nor U2141 (N_2141,In_182,In_2684);
and U2142 (N_2142,In_2770,In_2698);
nand U2143 (N_2143,In_399,In_1168);
and U2144 (N_2144,In_958,In_619);
nor U2145 (N_2145,In_290,In_2062);
xor U2146 (N_2146,In_2661,In_636);
nand U2147 (N_2147,In_1378,In_738);
and U2148 (N_2148,In_2700,In_2802);
nor U2149 (N_2149,In_1856,In_793);
xnor U2150 (N_2150,In_2273,In_1284);
nor U2151 (N_2151,In_703,In_113);
xor U2152 (N_2152,In_2314,In_523);
xor U2153 (N_2153,In_1250,In_715);
and U2154 (N_2154,In_2958,In_2248);
nand U2155 (N_2155,In_1533,In_1008);
or U2156 (N_2156,In_134,In_177);
and U2157 (N_2157,In_2471,In_1065);
or U2158 (N_2158,In_2398,In_1747);
xnor U2159 (N_2159,In_683,In_2258);
or U2160 (N_2160,In_568,In_2160);
or U2161 (N_2161,In_400,In_1702);
nor U2162 (N_2162,In_1662,In_177);
nor U2163 (N_2163,In_1136,In_498);
xnor U2164 (N_2164,In_239,In_230);
and U2165 (N_2165,In_2072,In_2931);
nand U2166 (N_2166,In_1125,In_747);
xnor U2167 (N_2167,In_2401,In_1709);
or U2168 (N_2168,In_772,In_880);
and U2169 (N_2169,In_1022,In_527);
or U2170 (N_2170,In_823,In_2679);
or U2171 (N_2171,In_161,In_2695);
and U2172 (N_2172,In_446,In_541);
xor U2173 (N_2173,In_811,In_1838);
nor U2174 (N_2174,In_2405,In_1111);
and U2175 (N_2175,In_2264,In_1221);
nand U2176 (N_2176,In_1813,In_1446);
and U2177 (N_2177,In_1815,In_774);
and U2178 (N_2178,In_2703,In_2538);
nor U2179 (N_2179,In_367,In_801);
and U2180 (N_2180,In_318,In_1943);
or U2181 (N_2181,In_2243,In_1574);
or U2182 (N_2182,In_2829,In_2039);
or U2183 (N_2183,In_1508,In_1387);
and U2184 (N_2184,In_951,In_712);
and U2185 (N_2185,In_1136,In_2581);
and U2186 (N_2186,In_2377,In_1661);
nand U2187 (N_2187,In_1745,In_37);
xnor U2188 (N_2188,In_322,In_2578);
nor U2189 (N_2189,In_1436,In_1665);
xnor U2190 (N_2190,In_2774,In_1712);
xor U2191 (N_2191,In_1801,In_1977);
nor U2192 (N_2192,In_324,In_122);
nand U2193 (N_2193,In_598,In_827);
nand U2194 (N_2194,In_532,In_334);
and U2195 (N_2195,In_298,In_680);
or U2196 (N_2196,In_13,In_305);
nand U2197 (N_2197,In_249,In_184);
or U2198 (N_2198,In_2368,In_160);
or U2199 (N_2199,In_113,In_2158);
or U2200 (N_2200,In_2670,In_1);
and U2201 (N_2201,In_1865,In_1638);
nor U2202 (N_2202,In_2665,In_13);
and U2203 (N_2203,In_959,In_2272);
nor U2204 (N_2204,In_474,In_2944);
nor U2205 (N_2205,In_1304,In_519);
and U2206 (N_2206,In_2092,In_1624);
xnor U2207 (N_2207,In_1535,In_2278);
nor U2208 (N_2208,In_258,In_1005);
nor U2209 (N_2209,In_1903,In_2189);
nor U2210 (N_2210,In_109,In_40);
or U2211 (N_2211,In_81,In_592);
xor U2212 (N_2212,In_1056,In_2434);
nor U2213 (N_2213,In_452,In_2371);
xor U2214 (N_2214,In_1472,In_14);
or U2215 (N_2215,In_2921,In_2875);
xnor U2216 (N_2216,In_1139,In_2752);
and U2217 (N_2217,In_1768,In_1554);
xor U2218 (N_2218,In_2608,In_2395);
or U2219 (N_2219,In_2405,In_1797);
nand U2220 (N_2220,In_2261,In_607);
and U2221 (N_2221,In_369,In_1476);
or U2222 (N_2222,In_2318,In_2702);
nand U2223 (N_2223,In_2166,In_2782);
or U2224 (N_2224,In_197,In_491);
or U2225 (N_2225,In_2202,In_776);
nand U2226 (N_2226,In_2306,In_400);
nor U2227 (N_2227,In_1135,In_119);
or U2228 (N_2228,In_2531,In_1061);
and U2229 (N_2229,In_1166,In_2683);
nand U2230 (N_2230,In_502,In_658);
nor U2231 (N_2231,In_2800,In_892);
xnor U2232 (N_2232,In_1685,In_1487);
nand U2233 (N_2233,In_2639,In_660);
xor U2234 (N_2234,In_1916,In_977);
nor U2235 (N_2235,In_2028,In_1573);
or U2236 (N_2236,In_664,In_2961);
nand U2237 (N_2237,In_593,In_723);
xor U2238 (N_2238,In_2410,In_8);
nand U2239 (N_2239,In_782,In_641);
and U2240 (N_2240,In_381,In_1577);
and U2241 (N_2241,In_1982,In_1151);
and U2242 (N_2242,In_929,In_2948);
or U2243 (N_2243,In_5,In_1475);
nand U2244 (N_2244,In_2844,In_353);
or U2245 (N_2245,In_1776,In_877);
nand U2246 (N_2246,In_2170,In_1454);
and U2247 (N_2247,In_2075,In_1605);
xor U2248 (N_2248,In_1545,In_284);
nor U2249 (N_2249,In_1177,In_1206);
nand U2250 (N_2250,In_753,In_1682);
nor U2251 (N_2251,In_1391,In_2124);
xor U2252 (N_2252,In_2645,In_1194);
xor U2253 (N_2253,In_151,In_1517);
nor U2254 (N_2254,In_100,In_1291);
nand U2255 (N_2255,In_1897,In_441);
nor U2256 (N_2256,In_170,In_2174);
or U2257 (N_2257,In_1377,In_687);
nor U2258 (N_2258,In_1043,In_454);
nand U2259 (N_2259,In_118,In_2107);
xor U2260 (N_2260,In_84,In_922);
nor U2261 (N_2261,In_2719,In_2756);
or U2262 (N_2262,In_2011,In_2094);
or U2263 (N_2263,In_2303,In_872);
nand U2264 (N_2264,In_1808,In_1446);
nor U2265 (N_2265,In_740,In_89);
and U2266 (N_2266,In_1756,In_2749);
nor U2267 (N_2267,In_93,In_2951);
nor U2268 (N_2268,In_2795,In_1959);
and U2269 (N_2269,In_2520,In_330);
xor U2270 (N_2270,In_137,In_0);
or U2271 (N_2271,In_1185,In_756);
or U2272 (N_2272,In_2755,In_1588);
xnor U2273 (N_2273,In_518,In_2233);
nor U2274 (N_2274,In_2083,In_2770);
xor U2275 (N_2275,In_1001,In_2651);
xnor U2276 (N_2276,In_444,In_2763);
and U2277 (N_2277,In_2309,In_1026);
nor U2278 (N_2278,In_2219,In_1926);
nand U2279 (N_2279,In_2212,In_2994);
or U2280 (N_2280,In_1575,In_2540);
nor U2281 (N_2281,In_595,In_2593);
or U2282 (N_2282,In_2046,In_412);
or U2283 (N_2283,In_2491,In_919);
xnor U2284 (N_2284,In_2799,In_1170);
nand U2285 (N_2285,In_1800,In_2643);
nand U2286 (N_2286,In_1573,In_2033);
xnor U2287 (N_2287,In_2109,In_2394);
nand U2288 (N_2288,In_1898,In_587);
and U2289 (N_2289,In_1321,In_1225);
nand U2290 (N_2290,In_2957,In_141);
nor U2291 (N_2291,In_2908,In_1823);
and U2292 (N_2292,In_1953,In_277);
xnor U2293 (N_2293,In_2982,In_954);
xnor U2294 (N_2294,In_1014,In_597);
and U2295 (N_2295,In_2178,In_1805);
xnor U2296 (N_2296,In_1317,In_1717);
nand U2297 (N_2297,In_2298,In_756);
nand U2298 (N_2298,In_327,In_72);
nor U2299 (N_2299,In_2855,In_2173);
and U2300 (N_2300,In_579,In_961);
or U2301 (N_2301,In_1956,In_149);
and U2302 (N_2302,In_904,In_2004);
nand U2303 (N_2303,In_140,In_1563);
nor U2304 (N_2304,In_135,In_1804);
nor U2305 (N_2305,In_2128,In_2287);
and U2306 (N_2306,In_827,In_403);
nor U2307 (N_2307,In_296,In_589);
nor U2308 (N_2308,In_1998,In_859);
nand U2309 (N_2309,In_1847,In_1709);
nor U2310 (N_2310,In_2152,In_102);
or U2311 (N_2311,In_1559,In_284);
and U2312 (N_2312,In_1792,In_2134);
and U2313 (N_2313,In_2429,In_2285);
xnor U2314 (N_2314,In_1864,In_549);
or U2315 (N_2315,In_927,In_229);
nand U2316 (N_2316,In_851,In_487);
nand U2317 (N_2317,In_1845,In_1228);
and U2318 (N_2318,In_1957,In_1263);
or U2319 (N_2319,In_298,In_2979);
xnor U2320 (N_2320,In_963,In_2180);
nand U2321 (N_2321,In_1186,In_1368);
xor U2322 (N_2322,In_431,In_611);
and U2323 (N_2323,In_1620,In_2757);
xnor U2324 (N_2324,In_2691,In_933);
or U2325 (N_2325,In_2955,In_1316);
xor U2326 (N_2326,In_776,In_1565);
or U2327 (N_2327,In_1285,In_2319);
nand U2328 (N_2328,In_1502,In_2042);
xnor U2329 (N_2329,In_2527,In_2697);
or U2330 (N_2330,In_250,In_2347);
or U2331 (N_2331,In_1483,In_1137);
or U2332 (N_2332,In_461,In_273);
nand U2333 (N_2333,In_687,In_875);
nor U2334 (N_2334,In_1169,In_1916);
xor U2335 (N_2335,In_2183,In_1202);
nand U2336 (N_2336,In_969,In_1407);
and U2337 (N_2337,In_2217,In_609);
nand U2338 (N_2338,In_2883,In_1976);
or U2339 (N_2339,In_1830,In_1079);
or U2340 (N_2340,In_1351,In_1067);
nand U2341 (N_2341,In_2893,In_1293);
nand U2342 (N_2342,In_2991,In_382);
and U2343 (N_2343,In_1553,In_1430);
xor U2344 (N_2344,In_2755,In_1663);
xor U2345 (N_2345,In_2286,In_1892);
xor U2346 (N_2346,In_1929,In_1163);
and U2347 (N_2347,In_265,In_34);
nor U2348 (N_2348,In_2565,In_1136);
nand U2349 (N_2349,In_1896,In_1851);
and U2350 (N_2350,In_2987,In_716);
nor U2351 (N_2351,In_2892,In_784);
xnor U2352 (N_2352,In_1511,In_267);
nand U2353 (N_2353,In_2029,In_107);
and U2354 (N_2354,In_2272,In_2215);
nor U2355 (N_2355,In_2678,In_322);
and U2356 (N_2356,In_2387,In_53);
nand U2357 (N_2357,In_2951,In_1523);
nand U2358 (N_2358,In_26,In_1432);
nand U2359 (N_2359,In_180,In_560);
xnor U2360 (N_2360,In_1191,In_1180);
nand U2361 (N_2361,In_2467,In_2536);
nor U2362 (N_2362,In_88,In_31);
xnor U2363 (N_2363,In_260,In_2448);
nor U2364 (N_2364,In_24,In_7);
xnor U2365 (N_2365,In_2669,In_733);
xnor U2366 (N_2366,In_2102,In_2972);
or U2367 (N_2367,In_2237,In_1008);
or U2368 (N_2368,In_427,In_1244);
and U2369 (N_2369,In_2160,In_1212);
and U2370 (N_2370,In_1430,In_1893);
or U2371 (N_2371,In_377,In_1358);
nand U2372 (N_2372,In_762,In_469);
xor U2373 (N_2373,In_685,In_2489);
xor U2374 (N_2374,In_955,In_1398);
xor U2375 (N_2375,In_2877,In_1368);
or U2376 (N_2376,In_1074,In_76);
or U2377 (N_2377,In_2577,In_1792);
or U2378 (N_2378,In_2538,In_138);
nand U2379 (N_2379,In_2709,In_895);
and U2380 (N_2380,In_2452,In_2536);
nand U2381 (N_2381,In_2238,In_1126);
and U2382 (N_2382,In_1264,In_1305);
nor U2383 (N_2383,In_1399,In_542);
nor U2384 (N_2384,In_717,In_1029);
nor U2385 (N_2385,In_955,In_2745);
and U2386 (N_2386,In_516,In_1160);
nand U2387 (N_2387,In_2662,In_610);
or U2388 (N_2388,In_857,In_2354);
nor U2389 (N_2389,In_25,In_725);
nand U2390 (N_2390,In_369,In_268);
nor U2391 (N_2391,In_376,In_2720);
xnor U2392 (N_2392,In_239,In_2773);
nand U2393 (N_2393,In_2736,In_1777);
nor U2394 (N_2394,In_677,In_834);
and U2395 (N_2395,In_314,In_1657);
xor U2396 (N_2396,In_2968,In_1601);
xnor U2397 (N_2397,In_2553,In_199);
and U2398 (N_2398,In_2525,In_2316);
or U2399 (N_2399,In_152,In_982);
nor U2400 (N_2400,In_834,In_1453);
and U2401 (N_2401,In_588,In_2299);
nor U2402 (N_2402,In_955,In_2706);
or U2403 (N_2403,In_2176,In_2472);
or U2404 (N_2404,In_2610,In_835);
nand U2405 (N_2405,In_2419,In_1652);
xnor U2406 (N_2406,In_2308,In_751);
xor U2407 (N_2407,In_685,In_1757);
xor U2408 (N_2408,In_1885,In_1489);
xor U2409 (N_2409,In_771,In_2568);
nand U2410 (N_2410,In_1964,In_77);
or U2411 (N_2411,In_1427,In_2791);
nor U2412 (N_2412,In_1679,In_514);
nand U2413 (N_2413,In_2771,In_1196);
nor U2414 (N_2414,In_163,In_577);
nand U2415 (N_2415,In_1854,In_1013);
xnor U2416 (N_2416,In_737,In_2348);
xnor U2417 (N_2417,In_766,In_402);
xor U2418 (N_2418,In_494,In_1358);
or U2419 (N_2419,In_572,In_2978);
or U2420 (N_2420,In_629,In_1847);
nand U2421 (N_2421,In_2509,In_2971);
nand U2422 (N_2422,In_2389,In_1663);
nand U2423 (N_2423,In_2498,In_2974);
or U2424 (N_2424,In_146,In_1485);
nor U2425 (N_2425,In_1716,In_129);
and U2426 (N_2426,In_853,In_919);
or U2427 (N_2427,In_380,In_2823);
nand U2428 (N_2428,In_2802,In_2321);
xnor U2429 (N_2429,In_2972,In_427);
or U2430 (N_2430,In_503,In_1984);
and U2431 (N_2431,In_2963,In_2224);
and U2432 (N_2432,In_1080,In_441);
or U2433 (N_2433,In_288,In_2781);
or U2434 (N_2434,In_2079,In_1097);
xor U2435 (N_2435,In_2615,In_2251);
nand U2436 (N_2436,In_9,In_60);
or U2437 (N_2437,In_2288,In_866);
xnor U2438 (N_2438,In_1008,In_3);
nor U2439 (N_2439,In_1113,In_1542);
and U2440 (N_2440,In_2701,In_335);
nand U2441 (N_2441,In_1318,In_1666);
nor U2442 (N_2442,In_2611,In_1331);
and U2443 (N_2443,In_529,In_2768);
nor U2444 (N_2444,In_980,In_1373);
xnor U2445 (N_2445,In_2068,In_741);
and U2446 (N_2446,In_1754,In_17);
xnor U2447 (N_2447,In_2317,In_1735);
xor U2448 (N_2448,In_1393,In_355);
or U2449 (N_2449,In_1556,In_2349);
xnor U2450 (N_2450,In_171,In_403);
and U2451 (N_2451,In_1489,In_556);
nor U2452 (N_2452,In_299,In_908);
and U2453 (N_2453,In_1874,In_1713);
nand U2454 (N_2454,In_1666,In_2679);
nor U2455 (N_2455,In_1196,In_2559);
nand U2456 (N_2456,In_372,In_718);
or U2457 (N_2457,In_2041,In_2260);
nor U2458 (N_2458,In_133,In_230);
nand U2459 (N_2459,In_1200,In_1790);
xor U2460 (N_2460,In_1560,In_2688);
and U2461 (N_2461,In_2532,In_2485);
xnor U2462 (N_2462,In_89,In_1213);
or U2463 (N_2463,In_367,In_1363);
or U2464 (N_2464,In_1262,In_2773);
and U2465 (N_2465,In_40,In_1377);
nand U2466 (N_2466,In_2899,In_2037);
nand U2467 (N_2467,In_1231,In_258);
nor U2468 (N_2468,In_1740,In_1440);
nand U2469 (N_2469,In_1159,In_321);
nand U2470 (N_2470,In_1928,In_796);
and U2471 (N_2471,In_776,In_1682);
and U2472 (N_2472,In_1922,In_2513);
or U2473 (N_2473,In_2262,In_2002);
nor U2474 (N_2474,In_2704,In_2636);
nor U2475 (N_2475,In_1945,In_2019);
xor U2476 (N_2476,In_2088,In_1784);
or U2477 (N_2477,In_567,In_284);
xor U2478 (N_2478,In_2418,In_283);
or U2479 (N_2479,In_995,In_829);
and U2480 (N_2480,In_415,In_1130);
nand U2481 (N_2481,In_2144,In_504);
xor U2482 (N_2482,In_2821,In_2168);
nand U2483 (N_2483,In_1210,In_2562);
nand U2484 (N_2484,In_1558,In_14);
or U2485 (N_2485,In_1823,In_2880);
xnor U2486 (N_2486,In_2060,In_552);
nand U2487 (N_2487,In_2161,In_1568);
nand U2488 (N_2488,In_1607,In_973);
xnor U2489 (N_2489,In_786,In_326);
nand U2490 (N_2490,In_2890,In_2334);
and U2491 (N_2491,In_271,In_546);
or U2492 (N_2492,In_98,In_446);
nor U2493 (N_2493,In_2317,In_444);
and U2494 (N_2494,In_137,In_75);
nand U2495 (N_2495,In_1889,In_947);
nor U2496 (N_2496,In_206,In_896);
and U2497 (N_2497,In_1092,In_2044);
nor U2498 (N_2498,In_421,In_557);
or U2499 (N_2499,In_585,In_2019);
nor U2500 (N_2500,In_1233,In_178);
or U2501 (N_2501,In_1750,In_1641);
or U2502 (N_2502,In_193,In_2090);
nor U2503 (N_2503,In_1268,In_2658);
and U2504 (N_2504,In_2460,In_1513);
nand U2505 (N_2505,In_333,In_1189);
or U2506 (N_2506,In_2929,In_1944);
and U2507 (N_2507,In_782,In_2880);
or U2508 (N_2508,In_884,In_2499);
nor U2509 (N_2509,In_1895,In_1257);
or U2510 (N_2510,In_894,In_1016);
nor U2511 (N_2511,In_1721,In_1300);
nor U2512 (N_2512,In_2794,In_2911);
and U2513 (N_2513,In_547,In_789);
xor U2514 (N_2514,In_2389,In_2366);
or U2515 (N_2515,In_2808,In_1745);
nand U2516 (N_2516,In_2724,In_354);
or U2517 (N_2517,In_2427,In_2912);
xnor U2518 (N_2518,In_1164,In_2848);
or U2519 (N_2519,In_1809,In_541);
nand U2520 (N_2520,In_576,In_649);
or U2521 (N_2521,In_794,In_1368);
nand U2522 (N_2522,In_504,In_838);
xnor U2523 (N_2523,In_2543,In_2590);
and U2524 (N_2524,In_2377,In_2796);
nand U2525 (N_2525,In_2513,In_29);
or U2526 (N_2526,In_1494,In_2986);
nor U2527 (N_2527,In_1454,In_2000);
nand U2528 (N_2528,In_2305,In_1186);
nor U2529 (N_2529,In_1275,In_2609);
xnor U2530 (N_2530,In_1608,In_957);
nor U2531 (N_2531,In_2276,In_1357);
nand U2532 (N_2532,In_1074,In_2313);
xor U2533 (N_2533,In_2253,In_1818);
and U2534 (N_2534,In_2224,In_1940);
xor U2535 (N_2535,In_1267,In_2906);
or U2536 (N_2536,In_1820,In_486);
xor U2537 (N_2537,In_2232,In_2332);
nand U2538 (N_2538,In_738,In_2003);
and U2539 (N_2539,In_763,In_2635);
xnor U2540 (N_2540,In_2188,In_387);
and U2541 (N_2541,In_1476,In_1017);
nor U2542 (N_2542,In_1439,In_2353);
xnor U2543 (N_2543,In_2882,In_788);
and U2544 (N_2544,In_1142,In_1683);
nor U2545 (N_2545,In_1206,In_2336);
nor U2546 (N_2546,In_2627,In_1794);
or U2547 (N_2547,In_1258,In_1520);
or U2548 (N_2548,In_871,In_152);
xor U2549 (N_2549,In_134,In_2151);
nand U2550 (N_2550,In_1396,In_1480);
or U2551 (N_2551,In_1165,In_416);
or U2552 (N_2552,In_457,In_1778);
xor U2553 (N_2553,In_2236,In_760);
and U2554 (N_2554,In_2487,In_1521);
nand U2555 (N_2555,In_2994,In_2974);
nand U2556 (N_2556,In_1736,In_1250);
and U2557 (N_2557,In_973,In_72);
or U2558 (N_2558,In_1086,In_2872);
nor U2559 (N_2559,In_1368,In_334);
or U2560 (N_2560,In_433,In_242);
nor U2561 (N_2561,In_797,In_1555);
or U2562 (N_2562,In_931,In_2447);
and U2563 (N_2563,In_2633,In_692);
or U2564 (N_2564,In_2194,In_2971);
nor U2565 (N_2565,In_1941,In_1542);
xnor U2566 (N_2566,In_1872,In_27);
and U2567 (N_2567,In_301,In_867);
nand U2568 (N_2568,In_1845,In_1421);
and U2569 (N_2569,In_2552,In_1523);
nand U2570 (N_2570,In_1307,In_440);
or U2571 (N_2571,In_1774,In_908);
nor U2572 (N_2572,In_2766,In_2844);
xnor U2573 (N_2573,In_2618,In_954);
nand U2574 (N_2574,In_1575,In_1184);
nand U2575 (N_2575,In_415,In_1765);
and U2576 (N_2576,In_1886,In_338);
or U2577 (N_2577,In_991,In_1834);
or U2578 (N_2578,In_2856,In_2953);
nor U2579 (N_2579,In_207,In_1806);
nor U2580 (N_2580,In_2767,In_349);
nand U2581 (N_2581,In_2521,In_1651);
and U2582 (N_2582,In_2673,In_496);
and U2583 (N_2583,In_1314,In_607);
and U2584 (N_2584,In_2802,In_1510);
xnor U2585 (N_2585,In_2277,In_783);
and U2586 (N_2586,In_950,In_494);
nand U2587 (N_2587,In_949,In_772);
or U2588 (N_2588,In_638,In_2484);
nand U2589 (N_2589,In_2869,In_2710);
xnor U2590 (N_2590,In_1281,In_1445);
xor U2591 (N_2591,In_1601,In_2917);
nor U2592 (N_2592,In_2952,In_1624);
nand U2593 (N_2593,In_1493,In_2774);
and U2594 (N_2594,In_1022,In_448);
or U2595 (N_2595,In_1087,In_2422);
or U2596 (N_2596,In_679,In_1150);
xnor U2597 (N_2597,In_2752,In_2433);
and U2598 (N_2598,In_2277,In_1435);
nor U2599 (N_2599,In_2454,In_2918);
or U2600 (N_2600,In_2322,In_633);
nor U2601 (N_2601,In_740,In_1199);
nor U2602 (N_2602,In_2864,In_2952);
or U2603 (N_2603,In_1382,In_1958);
and U2604 (N_2604,In_1564,In_63);
nor U2605 (N_2605,In_2907,In_579);
and U2606 (N_2606,In_2643,In_19);
and U2607 (N_2607,In_2662,In_1958);
nand U2608 (N_2608,In_1806,In_1501);
nand U2609 (N_2609,In_2383,In_1321);
xnor U2610 (N_2610,In_955,In_834);
xor U2611 (N_2611,In_408,In_544);
nor U2612 (N_2612,In_432,In_2739);
or U2613 (N_2613,In_994,In_2219);
or U2614 (N_2614,In_1085,In_2652);
and U2615 (N_2615,In_1563,In_86);
or U2616 (N_2616,In_2073,In_2483);
xnor U2617 (N_2617,In_2609,In_1953);
xnor U2618 (N_2618,In_967,In_2602);
nor U2619 (N_2619,In_1754,In_2812);
nor U2620 (N_2620,In_2467,In_778);
or U2621 (N_2621,In_2854,In_1426);
and U2622 (N_2622,In_34,In_476);
nand U2623 (N_2623,In_1695,In_1807);
nor U2624 (N_2624,In_2148,In_2784);
or U2625 (N_2625,In_1419,In_2500);
and U2626 (N_2626,In_2660,In_2262);
or U2627 (N_2627,In_2267,In_2417);
nand U2628 (N_2628,In_1868,In_1849);
nor U2629 (N_2629,In_2372,In_398);
xor U2630 (N_2630,In_2072,In_377);
nand U2631 (N_2631,In_1661,In_2444);
xnor U2632 (N_2632,In_2286,In_2368);
xor U2633 (N_2633,In_2797,In_2681);
or U2634 (N_2634,In_1194,In_2037);
nand U2635 (N_2635,In_1949,In_1347);
or U2636 (N_2636,In_2453,In_2285);
xnor U2637 (N_2637,In_1130,In_330);
or U2638 (N_2638,In_1862,In_1956);
nand U2639 (N_2639,In_2640,In_886);
or U2640 (N_2640,In_28,In_1069);
nand U2641 (N_2641,In_2783,In_1748);
nand U2642 (N_2642,In_1975,In_1728);
nor U2643 (N_2643,In_2140,In_1296);
and U2644 (N_2644,In_1849,In_1139);
nand U2645 (N_2645,In_2886,In_1763);
nor U2646 (N_2646,In_2311,In_249);
nor U2647 (N_2647,In_2673,In_2244);
nor U2648 (N_2648,In_672,In_866);
nand U2649 (N_2649,In_1231,In_2896);
and U2650 (N_2650,In_150,In_2417);
or U2651 (N_2651,In_2097,In_1798);
nand U2652 (N_2652,In_1253,In_2248);
or U2653 (N_2653,In_2286,In_553);
and U2654 (N_2654,In_1704,In_508);
nor U2655 (N_2655,In_2278,In_2450);
nor U2656 (N_2656,In_2096,In_613);
and U2657 (N_2657,In_1100,In_1477);
nor U2658 (N_2658,In_2960,In_2891);
nor U2659 (N_2659,In_284,In_801);
nor U2660 (N_2660,In_1303,In_2106);
or U2661 (N_2661,In_1005,In_1129);
nand U2662 (N_2662,In_1758,In_192);
or U2663 (N_2663,In_1787,In_2095);
xor U2664 (N_2664,In_2130,In_1684);
and U2665 (N_2665,In_2474,In_1995);
xor U2666 (N_2666,In_324,In_1506);
nand U2667 (N_2667,In_414,In_1798);
and U2668 (N_2668,In_805,In_217);
or U2669 (N_2669,In_2707,In_1433);
nor U2670 (N_2670,In_1926,In_1892);
and U2671 (N_2671,In_2272,In_2497);
xnor U2672 (N_2672,In_1629,In_2218);
xor U2673 (N_2673,In_1911,In_481);
nor U2674 (N_2674,In_2823,In_2339);
and U2675 (N_2675,In_1416,In_2459);
and U2676 (N_2676,In_2297,In_538);
and U2677 (N_2677,In_2395,In_1446);
xor U2678 (N_2678,In_621,In_1111);
nand U2679 (N_2679,In_2593,In_1427);
xnor U2680 (N_2680,In_1156,In_1044);
or U2681 (N_2681,In_675,In_2092);
xnor U2682 (N_2682,In_2908,In_2928);
nor U2683 (N_2683,In_1686,In_2968);
nand U2684 (N_2684,In_1670,In_1266);
or U2685 (N_2685,In_2923,In_2760);
and U2686 (N_2686,In_800,In_356);
xor U2687 (N_2687,In_6,In_658);
and U2688 (N_2688,In_598,In_157);
and U2689 (N_2689,In_824,In_2513);
or U2690 (N_2690,In_260,In_2141);
nand U2691 (N_2691,In_1532,In_1620);
or U2692 (N_2692,In_2370,In_1455);
xor U2693 (N_2693,In_702,In_2995);
xnor U2694 (N_2694,In_1744,In_309);
xnor U2695 (N_2695,In_656,In_2552);
nand U2696 (N_2696,In_1179,In_2994);
nor U2697 (N_2697,In_1222,In_1698);
and U2698 (N_2698,In_1259,In_954);
or U2699 (N_2699,In_2141,In_929);
nor U2700 (N_2700,In_1931,In_2417);
nand U2701 (N_2701,In_1860,In_2950);
nor U2702 (N_2702,In_2891,In_2557);
and U2703 (N_2703,In_2071,In_1826);
and U2704 (N_2704,In_993,In_1459);
xnor U2705 (N_2705,In_965,In_1866);
and U2706 (N_2706,In_2935,In_1895);
nor U2707 (N_2707,In_2459,In_556);
nor U2708 (N_2708,In_2407,In_1332);
and U2709 (N_2709,In_294,In_101);
and U2710 (N_2710,In_826,In_2865);
and U2711 (N_2711,In_915,In_2226);
and U2712 (N_2712,In_999,In_1038);
nand U2713 (N_2713,In_1867,In_1284);
nand U2714 (N_2714,In_1252,In_565);
xor U2715 (N_2715,In_179,In_2465);
nand U2716 (N_2716,In_705,In_906);
xnor U2717 (N_2717,In_1377,In_177);
nor U2718 (N_2718,In_2861,In_1550);
and U2719 (N_2719,In_740,In_1081);
xnor U2720 (N_2720,In_2175,In_1728);
nand U2721 (N_2721,In_781,In_1284);
and U2722 (N_2722,In_1393,In_2120);
xor U2723 (N_2723,In_2068,In_996);
or U2724 (N_2724,In_2478,In_31);
nand U2725 (N_2725,In_1952,In_1717);
nand U2726 (N_2726,In_327,In_1003);
and U2727 (N_2727,In_1521,In_861);
and U2728 (N_2728,In_123,In_2777);
or U2729 (N_2729,In_282,In_1428);
or U2730 (N_2730,In_1481,In_2679);
nor U2731 (N_2731,In_2080,In_1770);
and U2732 (N_2732,In_676,In_915);
nor U2733 (N_2733,In_1779,In_2056);
or U2734 (N_2734,In_1538,In_2878);
nor U2735 (N_2735,In_1716,In_2406);
nor U2736 (N_2736,In_401,In_2729);
nand U2737 (N_2737,In_2681,In_1549);
or U2738 (N_2738,In_2794,In_1323);
xnor U2739 (N_2739,In_2108,In_1878);
or U2740 (N_2740,In_2923,In_717);
nand U2741 (N_2741,In_2635,In_2894);
xor U2742 (N_2742,In_1847,In_1729);
nor U2743 (N_2743,In_1587,In_1956);
and U2744 (N_2744,In_2317,In_501);
or U2745 (N_2745,In_2619,In_249);
and U2746 (N_2746,In_2772,In_2069);
or U2747 (N_2747,In_209,In_2034);
and U2748 (N_2748,In_88,In_2640);
nor U2749 (N_2749,In_833,In_1733);
or U2750 (N_2750,In_1430,In_439);
nand U2751 (N_2751,In_447,In_2932);
and U2752 (N_2752,In_2186,In_963);
and U2753 (N_2753,In_1016,In_1902);
xnor U2754 (N_2754,In_1112,In_2211);
nor U2755 (N_2755,In_1563,In_159);
nand U2756 (N_2756,In_152,In_1591);
and U2757 (N_2757,In_2639,In_1325);
nand U2758 (N_2758,In_1519,In_187);
and U2759 (N_2759,In_1915,In_1756);
nand U2760 (N_2760,In_1333,In_1514);
and U2761 (N_2761,In_739,In_2067);
nor U2762 (N_2762,In_963,In_799);
nor U2763 (N_2763,In_1398,In_830);
xnor U2764 (N_2764,In_2478,In_1837);
or U2765 (N_2765,In_870,In_1060);
or U2766 (N_2766,In_1217,In_608);
xnor U2767 (N_2767,In_1226,In_2078);
nand U2768 (N_2768,In_2598,In_1690);
nor U2769 (N_2769,In_956,In_1277);
nor U2770 (N_2770,In_1178,In_952);
or U2771 (N_2771,In_129,In_818);
xor U2772 (N_2772,In_693,In_2886);
nand U2773 (N_2773,In_1721,In_2367);
and U2774 (N_2774,In_670,In_1609);
nand U2775 (N_2775,In_314,In_1097);
nand U2776 (N_2776,In_2491,In_1031);
xnor U2777 (N_2777,In_2330,In_870);
and U2778 (N_2778,In_731,In_293);
nand U2779 (N_2779,In_1117,In_2868);
or U2780 (N_2780,In_2516,In_2805);
xnor U2781 (N_2781,In_1609,In_1901);
xnor U2782 (N_2782,In_2899,In_1188);
xor U2783 (N_2783,In_1011,In_2560);
nor U2784 (N_2784,In_607,In_534);
nor U2785 (N_2785,In_1762,In_664);
or U2786 (N_2786,In_1196,In_2811);
and U2787 (N_2787,In_833,In_244);
and U2788 (N_2788,In_1761,In_2162);
and U2789 (N_2789,In_2665,In_837);
nor U2790 (N_2790,In_2096,In_1537);
and U2791 (N_2791,In_775,In_1491);
nor U2792 (N_2792,In_799,In_2972);
nand U2793 (N_2793,In_167,In_160);
or U2794 (N_2794,In_493,In_1463);
nor U2795 (N_2795,In_1124,In_1509);
nor U2796 (N_2796,In_870,In_2139);
nand U2797 (N_2797,In_183,In_1105);
nor U2798 (N_2798,In_228,In_1065);
nand U2799 (N_2799,In_1824,In_1412);
xnor U2800 (N_2800,In_1599,In_2680);
xnor U2801 (N_2801,In_1097,In_232);
or U2802 (N_2802,In_1742,In_131);
xor U2803 (N_2803,In_2023,In_1170);
nor U2804 (N_2804,In_2963,In_1882);
or U2805 (N_2805,In_1587,In_1855);
and U2806 (N_2806,In_2206,In_951);
or U2807 (N_2807,In_455,In_1316);
and U2808 (N_2808,In_525,In_981);
and U2809 (N_2809,In_1240,In_1295);
nor U2810 (N_2810,In_1871,In_852);
nand U2811 (N_2811,In_2026,In_2680);
xnor U2812 (N_2812,In_2665,In_1782);
and U2813 (N_2813,In_1983,In_1167);
nor U2814 (N_2814,In_534,In_363);
and U2815 (N_2815,In_1318,In_489);
nor U2816 (N_2816,In_201,In_439);
nand U2817 (N_2817,In_2562,In_655);
and U2818 (N_2818,In_1745,In_2160);
and U2819 (N_2819,In_494,In_2654);
or U2820 (N_2820,In_255,In_1014);
and U2821 (N_2821,In_274,In_2608);
nor U2822 (N_2822,In_1938,In_2243);
xor U2823 (N_2823,In_2202,In_1261);
or U2824 (N_2824,In_2895,In_2953);
or U2825 (N_2825,In_1024,In_1879);
nand U2826 (N_2826,In_792,In_2737);
or U2827 (N_2827,In_2499,In_618);
or U2828 (N_2828,In_2417,In_1343);
and U2829 (N_2829,In_254,In_2172);
xor U2830 (N_2830,In_759,In_207);
xnor U2831 (N_2831,In_885,In_191);
or U2832 (N_2832,In_820,In_508);
or U2833 (N_2833,In_743,In_798);
or U2834 (N_2834,In_1575,In_2068);
nor U2835 (N_2835,In_419,In_1257);
nand U2836 (N_2836,In_501,In_882);
or U2837 (N_2837,In_344,In_1676);
and U2838 (N_2838,In_1134,In_2145);
or U2839 (N_2839,In_71,In_2112);
xor U2840 (N_2840,In_600,In_421);
xnor U2841 (N_2841,In_2630,In_511);
nand U2842 (N_2842,In_728,In_670);
xnor U2843 (N_2843,In_888,In_316);
and U2844 (N_2844,In_10,In_2452);
xor U2845 (N_2845,In_1242,In_140);
nor U2846 (N_2846,In_2190,In_2042);
and U2847 (N_2847,In_1755,In_2416);
nand U2848 (N_2848,In_2079,In_584);
xnor U2849 (N_2849,In_404,In_1208);
nor U2850 (N_2850,In_875,In_1789);
xor U2851 (N_2851,In_176,In_2662);
xnor U2852 (N_2852,In_2904,In_2824);
xnor U2853 (N_2853,In_2815,In_1358);
and U2854 (N_2854,In_1362,In_2761);
or U2855 (N_2855,In_1794,In_2757);
or U2856 (N_2856,In_954,In_658);
nand U2857 (N_2857,In_1036,In_770);
nor U2858 (N_2858,In_2543,In_660);
xnor U2859 (N_2859,In_1457,In_1368);
nand U2860 (N_2860,In_1768,In_2097);
nor U2861 (N_2861,In_2231,In_2886);
or U2862 (N_2862,In_1769,In_2951);
nand U2863 (N_2863,In_8,In_1810);
xor U2864 (N_2864,In_465,In_463);
nor U2865 (N_2865,In_1951,In_1460);
or U2866 (N_2866,In_292,In_172);
nand U2867 (N_2867,In_2976,In_2347);
nand U2868 (N_2868,In_697,In_1912);
nor U2869 (N_2869,In_1362,In_1221);
nand U2870 (N_2870,In_815,In_1872);
nor U2871 (N_2871,In_2818,In_2812);
xnor U2872 (N_2872,In_1639,In_939);
xnor U2873 (N_2873,In_2954,In_1297);
xnor U2874 (N_2874,In_1932,In_2486);
nor U2875 (N_2875,In_2024,In_582);
nor U2876 (N_2876,In_1923,In_1809);
or U2877 (N_2877,In_2213,In_1996);
xnor U2878 (N_2878,In_1127,In_2251);
xnor U2879 (N_2879,In_489,In_1741);
xnor U2880 (N_2880,In_1497,In_2950);
or U2881 (N_2881,In_89,In_1890);
or U2882 (N_2882,In_1128,In_1892);
or U2883 (N_2883,In_1689,In_804);
and U2884 (N_2884,In_763,In_425);
nor U2885 (N_2885,In_1799,In_1227);
nor U2886 (N_2886,In_2440,In_1082);
and U2887 (N_2887,In_680,In_752);
xnor U2888 (N_2888,In_2604,In_1823);
and U2889 (N_2889,In_2277,In_2576);
nand U2890 (N_2890,In_1000,In_1946);
nor U2891 (N_2891,In_774,In_471);
nand U2892 (N_2892,In_718,In_333);
xnor U2893 (N_2893,In_1436,In_70);
nand U2894 (N_2894,In_118,In_1278);
nand U2895 (N_2895,In_451,In_2452);
nor U2896 (N_2896,In_1117,In_1329);
and U2897 (N_2897,In_1395,In_539);
or U2898 (N_2898,In_275,In_779);
nand U2899 (N_2899,In_1922,In_2582);
or U2900 (N_2900,In_2668,In_2057);
and U2901 (N_2901,In_2610,In_653);
or U2902 (N_2902,In_2861,In_1996);
nor U2903 (N_2903,In_2679,In_885);
nand U2904 (N_2904,In_1922,In_1456);
nor U2905 (N_2905,In_1873,In_2537);
nand U2906 (N_2906,In_131,In_2749);
and U2907 (N_2907,In_1593,In_2770);
nand U2908 (N_2908,In_1480,In_1060);
and U2909 (N_2909,In_1564,In_1328);
and U2910 (N_2910,In_64,In_2408);
nand U2911 (N_2911,In_647,In_322);
nor U2912 (N_2912,In_2553,In_1716);
nand U2913 (N_2913,In_1852,In_2740);
xor U2914 (N_2914,In_2970,In_2316);
and U2915 (N_2915,In_2895,In_2584);
or U2916 (N_2916,In_2639,In_1414);
nand U2917 (N_2917,In_2600,In_2681);
xor U2918 (N_2918,In_2821,In_2029);
xor U2919 (N_2919,In_1966,In_2687);
nand U2920 (N_2920,In_260,In_544);
or U2921 (N_2921,In_990,In_1507);
and U2922 (N_2922,In_854,In_1893);
xor U2923 (N_2923,In_2097,In_167);
nor U2924 (N_2924,In_1637,In_1673);
nor U2925 (N_2925,In_2684,In_1927);
and U2926 (N_2926,In_2457,In_543);
and U2927 (N_2927,In_1176,In_2187);
nand U2928 (N_2928,In_1750,In_515);
or U2929 (N_2929,In_398,In_700);
and U2930 (N_2930,In_2554,In_2630);
xnor U2931 (N_2931,In_385,In_1325);
or U2932 (N_2932,In_1963,In_2657);
xor U2933 (N_2933,In_1765,In_422);
or U2934 (N_2934,In_2874,In_2941);
nor U2935 (N_2935,In_2117,In_2009);
or U2936 (N_2936,In_255,In_836);
nor U2937 (N_2937,In_2349,In_2229);
xnor U2938 (N_2938,In_57,In_320);
xor U2939 (N_2939,In_98,In_571);
and U2940 (N_2940,In_71,In_446);
or U2941 (N_2941,In_207,In_549);
or U2942 (N_2942,In_708,In_1194);
nand U2943 (N_2943,In_1568,In_2658);
or U2944 (N_2944,In_1079,In_2662);
nor U2945 (N_2945,In_1430,In_1521);
xnor U2946 (N_2946,In_2953,In_638);
and U2947 (N_2947,In_2494,In_535);
xnor U2948 (N_2948,In_1378,In_2074);
nor U2949 (N_2949,In_990,In_2556);
or U2950 (N_2950,In_1702,In_1991);
or U2951 (N_2951,In_2772,In_1711);
or U2952 (N_2952,In_2404,In_2691);
nor U2953 (N_2953,In_1053,In_2649);
nor U2954 (N_2954,In_725,In_1884);
nand U2955 (N_2955,In_2087,In_1482);
and U2956 (N_2956,In_656,In_2724);
nor U2957 (N_2957,In_1217,In_2647);
nand U2958 (N_2958,In_1033,In_1136);
nor U2959 (N_2959,In_586,In_2387);
nor U2960 (N_2960,In_1505,In_2306);
and U2961 (N_2961,In_2116,In_2752);
or U2962 (N_2962,In_1448,In_2601);
nand U2963 (N_2963,In_531,In_2522);
xor U2964 (N_2964,In_337,In_1820);
and U2965 (N_2965,In_1451,In_2516);
or U2966 (N_2966,In_2762,In_1965);
and U2967 (N_2967,In_1531,In_679);
or U2968 (N_2968,In_219,In_1344);
nand U2969 (N_2969,In_339,In_23);
nor U2970 (N_2970,In_275,In_2514);
nand U2971 (N_2971,In_543,In_1221);
xor U2972 (N_2972,In_2567,In_2639);
nor U2973 (N_2973,In_126,In_1587);
nand U2974 (N_2974,In_2593,In_2144);
nor U2975 (N_2975,In_2334,In_2999);
or U2976 (N_2976,In_1378,In_1168);
xnor U2977 (N_2977,In_172,In_1778);
nor U2978 (N_2978,In_1933,In_2658);
xor U2979 (N_2979,In_1204,In_262);
nand U2980 (N_2980,In_877,In_2698);
and U2981 (N_2981,In_1999,In_2599);
nand U2982 (N_2982,In_2683,In_2105);
or U2983 (N_2983,In_659,In_1467);
nand U2984 (N_2984,In_1779,In_1674);
or U2985 (N_2985,In_1174,In_2132);
or U2986 (N_2986,In_2999,In_2868);
and U2987 (N_2987,In_346,In_216);
xor U2988 (N_2988,In_2089,In_657);
xnor U2989 (N_2989,In_1097,In_2523);
xor U2990 (N_2990,In_1170,In_1328);
nand U2991 (N_2991,In_2478,In_434);
nand U2992 (N_2992,In_367,In_610);
nor U2993 (N_2993,In_957,In_253);
nor U2994 (N_2994,In_762,In_1878);
xor U2995 (N_2995,In_1080,In_1656);
nor U2996 (N_2996,In_979,In_1667);
xnor U2997 (N_2997,In_1080,In_1829);
and U2998 (N_2998,In_102,In_1617);
or U2999 (N_2999,In_616,In_1253);
nand U3000 (N_3000,In_586,In_1801);
xnor U3001 (N_3001,In_1441,In_155);
nor U3002 (N_3002,In_1668,In_2640);
nand U3003 (N_3003,In_2968,In_2106);
and U3004 (N_3004,In_1527,In_27);
and U3005 (N_3005,In_724,In_2316);
nand U3006 (N_3006,In_871,In_2699);
nand U3007 (N_3007,In_2779,In_1761);
or U3008 (N_3008,In_597,In_548);
and U3009 (N_3009,In_2366,In_630);
xor U3010 (N_3010,In_1652,In_1999);
and U3011 (N_3011,In_1923,In_1082);
or U3012 (N_3012,In_2532,In_944);
and U3013 (N_3013,In_2676,In_2420);
nand U3014 (N_3014,In_654,In_658);
nand U3015 (N_3015,In_2314,In_2902);
nor U3016 (N_3016,In_2507,In_2827);
nor U3017 (N_3017,In_48,In_1237);
xor U3018 (N_3018,In_2118,In_2322);
and U3019 (N_3019,In_1830,In_799);
and U3020 (N_3020,In_1965,In_755);
xnor U3021 (N_3021,In_392,In_1443);
and U3022 (N_3022,In_2759,In_2245);
or U3023 (N_3023,In_2085,In_1911);
nand U3024 (N_3024,In_476,In_801);
or U3025 (N_3025,In_993,In_2394);
nand U3026 (N_3026,In_1315,In_1454);
xor U3027 (N_3027,In_12,In_2221);
xor U3028 (N_3028,In_1183,In_332);
nor U3029 (N_3029,In_2264,In_1709);
nand U3030 (N_3030,In_2804,In_11);
xnor U3031 (N_3031,In_2096,In_2590);
nand U3032 (N_3032,In_942,In_2409);
xor U3033 (N_3033,In_1794,In_193);
and U3034 (N_3034,In_504,In_954);
nand U3035 (N_3035,In_569,In_1372);
nor U3036 (N_3036,In_1091,In_2907);
and U3037 (N_3037,In_1700,In_942);
xor U3038 (N_3038,In_2216,In_1467);
or U3039 (N_3039,In_2180,In_2087);
xor U3040 (N_3040,In_2715,In_1263);
and U3041 (N_3041,In_982,In_1341);
xnor U3042 (N_3042,In_673,In_690);
nand U3043 (N_3043,In_2110,In_2836);
and U3044 (N_3044,In_2942,In_920);
nor U3045 (N_3045,In_2490,In_2907);
or U3046 (N_3046,In_2149,In_2341);
or U3047 (N_3047,In_730,In_2357);
xor U3048 (N_3048,In_2932,In_44);
nand U3049 (N_3049,In_1348,In_2230);
xnor U3050 (N_3050,In_2126,In_2153);
xnor U3051 (N_3051,In_2343,In_1709);
nor U3052 (N_3052,In_289,In_193);
xor U3053 (N_3053,In_1198,In_1595);
nand U3054 (N_3054,In_2407,In_859);
nor U3055 (N_3055,In_1796,In_1752);
nor U3056 (N_3056,In_2461,In_1881);
or U3057 (N_3057,In_179,In_2311);
or U3058 (N_3058,In_2944,In_2697);
nand U3059 (N_3059,In_1813,In_378);
or U3060 (N_3060,In_1010,In_1138);
nor U3061 (N_3061,In_520,In_1561);
and U3062 (N_3062,In_2267,In_1685);
xor U3063 (N_3063,In_197,In_2631);
nor U3064 (N_3064,In_2350,In_525);
xor U3065 (N_3065,In_1935,In_407);
nand U3066 (N_3066,In_2102,In_253);
nand U3067 (N_3067,In_302,In_244);
nand U3068 (N_3068,In_174,In_2292);
nor U3069 (N_3069,In_2795,In_2532);
and U3070 (N_3070,In_689,In_2676);
xnor U3071 (N_3071,In_529,In_2342);
nor U3072 (N_3072,In_2363,In_951);
nor U3073 (N_3073,In_2846,In_2958);
nand U3074 (N_3074,In_2488,In_615);
and U3075 (N_3075,In_1997,In_66);
or U3076 (N_3076,In_1169,In_2398);
nor U3077 (N_3077,In_2294,In_321);
nor U3078 (N_3078,In_840,In_2638);
xnor U3079 (N_3079,In_2751,In_1724);
or U3080 (N_3080,In_391,In_14);
or U3081 (N_3081,In_556,In_259);
xnor U3082 (N_3082,In_2098,In_1299);
and U3083 (N_3083,In_2636,In_2264);
nor U3084 (N_3084,In_2842,In_735);
xnor U3085 (N_3085,In_1270,In_1784);
and U3086 (N_3086,In_162,In_1991);
or U3087 (N_3087,In_2680,In_1678);
and U3088 (N_3088,In_205,In_2801);
or U3089 (N_3089,In_926,In_2386);
xor U3090 (N_3090,In_1923,In_1751);
or U3091 (N_3091,In_1948,In_2073);
nand U3092 (N_3092,In_387,In_1807);
nand U3093 (N_3093,In_2793,In_2384);
xnor U3094 (N_3094,In_903,In_2771);
nand U3095 (N_3095,In_1893,In_165);
xnor U3096 (N_3096,In_383,In_1028);
xnor U3097 (N_3097,In_1843,In_1363);
xnor U3098 (N_3098,In_2671,In_690);
nand U3099 (N_3099,In_1513,In_1958);
xor U3100 (N_3100,In_1669,In_1154);
or U3101 (N_3101,In_685,In_2876);
or U3102 (N_3102,In_2235,In_472);
nand U3103 (N_3103,In_2862,In_1325);
or U3104 (N_3104,In_1699,In_991);
or U3105 (N_3105,In_2253,In_2184);
and U3106 (N_3106,In_934,In_46);
or U3107 (N_3107,In_2844,In_198);
or U3108 (N_3108,In_2234,In_1813);
or U3109 (N_3109,In_529,In_1602);
and U3110 (N_3110,In_2457,In_239);
nand U3111 (N_3111,In_2311,In_2835);
or U3112 (N_3112,In_2792,In_808);
and U3113 (N_3113,In_806,In_2406);
and U3114 (N_3114,In_1585,In_862);
or U3115 (N_3115,In_2569,In_1667);
nor U3116 (N_3116,In_592,In_1299);
xor U3117 (N_3117,In_1561,In_580);
and U3118 (N_3118,In_1628,In_843);
or U3119 (N_3119,In_1303,In_466);
nor U3120 (N_3120,In_2940,In_2388);
or U3121 (N_3121,In_1406,In_1948);
xnor U3122 (N_3122,In_2561,In_2458);
xor U3123 (N_3123,In_2890,In_2651);
nand U3124 (N_3124,In_1869,In_1714);
xor U3125 (N_3125,In_2402,In_1472);
nor U3126 (N_3126,In_1885,In_1612);
xnor U3127 (N_3127,In_1928,In_180);
xor U3128 (N_3128,In_2314,In_1060);
nor U3129 (N_3129,In_2944,In_1687);
and U3130 (N_3130,In_439,In_616);
or U3131 (N_3131,In_1347,In_2330);
xor U3132 (N_3132,In_831,In_1615);
nor U3133 (N_3133,In_198,In_1551);
xnor U3134 (N_3134,In_1070,In_2937);
and U3135 (N_3135,In_6,In_1125);
nand U3136 (N_3136,In_830,In_1961);
xor U3137 (N_3137,In_2654,In_1772);
xor U3138 (N_3138,In_2278,In_2030);
or U3139 (N_3139,In_631,In_1310);
nor U3140 (N_3140,In_1035,In_2527);
or U3141 (N_3141,In_8,In_252);
and U3142 (N_3142,In_967,In_14);
or U3143 (N_3143,In_273,In_1485);
nand U3144 (N_3144,In_2315,In_1236);
nand U3145 (N_3145,In_2321,In_2987);
nor U3146 (N_3146,In_1059,In_1296);
xor U3147 (N_3147,In_928,In_1965);
nand U3148 (N_3148,In_1578,In_1069);
nor U3149 (N_3149,In_429,In_2303);
nand U3150 (N_3150,In_2133,In_1872);
xnor U3151 (N_3151,In_1856,In_1566);
xnor U3152 (N_3152,In_2285,In_377);
and U3153 (N_3153,In_2449,In_329);
or U3154 (N_3154,In_1667,In_675);
xor U3155 (N_3155,In_1986,In_470);
nor U3156 (N_3156,In_1391,In_934);
or U3157 (N_3157,In_1065,In_2772);
nor U3158 (N_3158,In_940,In_1658);
nor U3159 (N_3159,In_1234,In_672);
nor U3160 (N_3160,In_2101,In_1649);
nor U3161 (N_3161,In_1431,In_2907);
nor U3162 (N_3162,In_2536,In_1430);
nor U3163 (N_3163,In_923,In_832);
or U3164 (N_3164,In_2187,In_1756);
or U3165 (N_3165,In_1669,In_1960);
and U3166 (N_3166,In_1736,In_887);
or U3167 (N_3167,In_225,In_1662);
nor U3168 (N_3168,In_2816,In_1782);
or U3169 (N_3169,In_208,In_2504);
nand U3170 (N_3170,In_1013,In_631);
xor U3171 (N_3171,In_2069,In_421);
xor U3172 (N_3172,In_2057,In_1641);
and U3173 (N_3173,In_1947,In_458);
xnor U3174 (N_3174,In_138,In_2956);
or U3175 (N_3175,In_1573,In_1623);
xnor U3176 (N_3176,In_1565,In_1085);
xor U3177 (N_3177,In_2639,In_132);
and U3178 (N_3178,In_2452,In_1686);
nor U3179 (N_3179,In_2046,In_2277);
nor U3180 (N_3180,In_90,In_2475);
or U3181 (N_3181,In_709,In_2403);
and U3182 (N_3182,In_255,In_1613);
and U3183 (N_3183,In_763,In_2894);
nor U3184 (N_3184,In_1730,In_285);
nand U3185 (N_3185,In_470,In_2392);
or U3186 (N_3186,In_1119,In_1690);
or U3187 (N_3187,In_2951,In_2611);
or U3188 (N_3188,In_340,In_1108);
xnor U3189 (N_3189,In_14,In_1722);
and U3190 (N_3190,In_2031,In_288);
and U3191 (N_3191,In_1784,In_165);
nand U3192 (N_3192,In_2139,In_1265);
nor U3193 (N_3193,In_962,In_269);
nor U3194 (N_3194,In_1344,In_456);
xnor U3195 (N_3195,In_603,In_1731);
and U3196 (N_3196,In_1681,In_1792);
and U3197 (N_3197,In_1968,In_2841);
nand U3198 (N_3198,In_1097,In_1111);
nor U3199 (N_3199,In_1475,In_1054);
or U3200 (N_3200,In_2738,In_711);
or U3201 (N_3201,In_1809,In_1617);
and U3202 (N_3202,In_731,In_2037);
xor U3203 (N_3203,In_1220,In_2010);
or U3204 (N_3204,In_555,In_367);
and U3205 (N_3205,In_928,In_995);
and U3206 (N_3206,In_2619,In_1195);
nand U3207 (N_3207,In_2261,In_2195);
nand U3208 (N_3208,In_2272,In_2011);
nand U3209 (N_3209,In_2953,In_870);
or U3210 (N_3210,In_2673,In_2892);
nor U3211 (N_3211,In_1022,In_2680);
and U3212 (N_3212,In_901,In_1077);
nand U3213 (N_3213,In_942,In_1405);
nor U3214 (N_3214,In_2461,In_1387);
nand U3215 (N_3215,In_2263,In_2204);
and U3216 (N_3216,In_2980,In_1459);
xor U3217 (N_3217,In_424,In_1658);
or U3218 (N_3218,In_831,In_1023);
xor U3219 (N_3219,In_953,In_2457);
xor U3220 (N_3220,In_1357,In_236);
xnor U3221 (N_3221,In_2689,In_2521);
nand U3222 (N_3222,In_1019,In_1947);
nor U3223 (N_3223,In_1760,In_1243);
nand U3224 (N_3224,In_2834,In_1134);
xor U3225 (N_3225,In_848,In_1642);
or U3226 (N_3226,In_2912,In_2176);
xor U3227 (N_3227,In_1850,In_939);
and U3228 (N_3228,In_2145,In_1761);
and U3229 (N_3229,In_592,In_2670);
xnor U3230 (N_3230,In_379,In_2705);
xnor U3231 (N_3231,In_1227,In_2303);
and U3232 (N_3232,In_126,In_563);
xnor U3233 (N_3233,In_717,In_2337);
xnor U3234 (N_3234,In_2201,In_1424);
and U3235 (N_3235,In_1951,In_2899);
or U3236 (N_3236,In_1315,In_2144);
nand U3237 (N_3237,In_2151,In_1011);
and U3238 (N_3238,In_2661,In_961);
nand U3239 (N_3239,In_2860,In_1942);
xnor U3240 (N_3240,In_1039,In_2092);
nor U3241 (N_3241,In_2187,In_2516);
xor U3242 (N_3242,In_2330,In_1920);
xor U3243 (N_3243,In_1706,In_48);
and U3244 (N_3244,In_1503,In_1361);
nor U3245 (N_3245,In_1625,In_968);
and U3246 (N_3246,In_2194,In_369);
or U3247 (N_3247,In_494,In_848);
and U3248 (N_3248,In_2357,In_2614);
and U3249 (N_3249,In_800,In_1714);
xor U3250 (N_3250,In_2126,In_2520);
and U3251 (N_3251,In_2255,In_2177);
nor U3252 (N_3252,In_2426,In_581);
nand U3253 (N_3253,In_1160,In_466);
nor U3254 (N_3254,In_2719,In_2551);
and U3255 (N_3255,In_2976,In_2523);
and U3256 (N_3256,In_2845,In_80);
and U3257 (N_3257,In_771,In_2516);
nor U3258 (N_3258,In_1527,In_1997);
nor U3259 (N_3259,In_1407,In_2576);
nand U3260 (N_3260,In_1271,In_1676);
and U3261 (N_3261,In_772,In_1969);
xnor U3262 (N_3262,In_2912,In_2180);
nand U3263 (N_3263,In_982,In_2616);
xor U3264 (N_3264,In_2980,In_98);
nand U3265 (N_3265,In_1364,In_917);
nor U3266 (N_3266,In_437,In_2770);
nor U3267 (N_3267,In_1077,In_2640);
and U3268 (N_3268,In_546,In_640);
and U3269 (N_3269,In_807,In_223);
or U3270 (N_3270,In_2375,In_2942);
and U3271 (N_3271,In_1177,In_2301);
and U3272 (N_3272,In_2669,In_1040);
or U3273 (N_3273,In_2424,In_64);
nor U3274 (N_3274,In_1635,In_1174);
and U3275 (N_3275,In_1849,In_993);
xnor U3276 (N_3276,In_2252,In_1091);
nor U3277 (N_3277,In_2017,In_2717);
nand U3278 (N_3278,In_2830,In_448);
and U3279 (N_3279,In_1114,In_109);
or U3280 (N_3280,In_1695,In_2866);
nor U3281 (N_3281,In_2490,In_93);
or U3282 (N_3282,In_644,In_1242);
or U3283 (N_3283,In_396,In_2175);
nand U3284 (N_3284,In_1090,In_2704);
nand U3285 (N_3285,In_2640,In_1983);
nor U3286 (N_3286,In_2148,In_1304);
xor U3287 (N_3287,In_2359,In_2015);
or U3288 (N_3288,In_642,In_1570);
or U3289 (N_3289,In_1095,In_1971);
and U3290 (N_3290,In_1508,In_862);
nor U3291 (N_3291,In_2489,In_2585);
and U3292 (N_3292,In_1361,In_2139);
or U3293 (N_3293,In_1259,In_538);
nand U3294 (N_3294,In_1591,In_1268);
and U3295 (N_3295,In_1033,In_2586);
or U3296 (N_3296,In_2728,In_824);
nand U3297 (N_3297,In_2548,In_1587);
or U3298 (N_3298,In_866,In_1368);
and U3299 (N_3299,In_175,In_478);
nor U3300 (N_3300,In_1358,In_199);
and U3301 (N_3301,In_1485,In_1265);
xnor U3302 (N_3302,In_396,In_498);
xnor U3303 (N_3303,In_2707,In_776);
nor U3304 (N_3304,In_149,In_734);
xor U3305 (N_3305,In_2842,In_2771);
xnor U3306 (N_3306,In_2231,In_1679);
and U3307 (N_3307,In_2375,In_892);
and U3308 (N_3308,In_269,In_2840);
xor U3309 (N_3309,In_695,In_2304);
nor U3310 (N_3310,In_1659,In_1944);
and U3311 (N_3311,In_1006,In_1796);
nand U3312 (N_3312,In_1993,In_2358);
and U3313 (N_3313,In_2669,In_1554);
nor U3314 (N_3314,In_1060,In_2739);
nor U3315 (N_3315,In_2614,In_216);
or U3316 (N_3316,In_1424,In_37);
xnor U3317 (N_3317,In_1894,In_1019);
and U3318 (N_3318,In_1284,In_873);
nand U3319 (N_3319,In_774,In_982);
xor U3320 (N_3320,In_598,In_953);
and U3321 (N_3321,In_2737,In_28);
or U3322 (N_3322,In_2701,In_1294);
and U3323 (N_3323,In_777,In_158);
nand U3324 (N_3324,In_590,In_238);
nor U3325 (N_3325,In_1289,In_1923);
or U3326 (N_3326,In_73,In_1275);
xor U3327 (N_3327,In_1342,In_653);
and U3328 (N_3328,In_2152,In_2659);
nand U3329 (N_3329,In_1660,In_1329);
nor U3330 (N_3330,In_2295,In_2643);
or U3331 (N_3331,In_2568,In_2426);
or U3332 (N_3332,In_2631,In_2281);
or U3333 (N_3333,In_1010,In_1931);
and U3334 (N_3334,In_1374,In_954);
nor U3335 (N_3335,In_616,In_2589);
nor U3336 (N_3336,In_1484,In_1829);
nor U3337 (N_3337,In_1893,In_691);
xor U3338 (N_3338,In_974,In_2401);
or U3339 (N_3339,In_2007,In_2417);
and U3340 (N_3340,In_586,In_79);
or U3341 (N_3341,In_1610,In_1646);
nor U3342 (N_3342,In_1090,In_2039);
nand U3343 (N_3343,In_586,In_1529);
and U3344 (N_3344,In_1008,In_2122);
nand U3345 (N_3345,In_262,In_1846);
xnor U3346 (N_3346,In_1774,In_2455);
nand U3347 (N_3347,In_1960,In_496);
nor U3348 (N_3348,In_2596,In_154);
nor U3349 (N_3349,In_1571,In_1913);
nand U3350 (N_3350,In_1471,In_2430);
xnor U3351 (N_3351,In_1844,In_1007);
nand U3352 (N_3352,In_158,In_992);
and U3353 (N_3353,In_2550,In_2873);
or U3354 (N_3354,In_1414,In_536);
or U3355 (N_3355,In_2440,In_2128);
xor U3356 (N_3356,In_1844,In_449);
xor U3357 (N_3357,In_965,In_1933);
nand U3358 (N_3358,In_524,In_1250);
nor U3359 (N_3359,In_2431,In_1548);
nor U3360 (N_3360,In_1840,In_1523);
nor U3361 (N_3361,In_2199,In_1834);
nand U3362 (N_3362,In_2601,In_2998);
and U3363 (N_3363,In_0,In_2234);
or U3364 (N_3364,In_1837,In_167);
xor U3365 (N_3365,In_925,In_2578);
and U3366 (N_3366,In_1545,In_405);
or U3367 (N_3367,In_2894,In_2419);
nand U3368 (N_3368,In_545,In_1601);
nor U3369 (N_3369,In_200,In_1270);
nor U3370 (N_3370,In_2316,In_214);
nor U3371 (N_3371,In_747,In_2668);
xnor U3372 (N_3372,In_87,In_2318);
xnor U3373 (N_3373,In_2144,In_2715);
xor U3374 (N_3374,In_577,In_1069);
or U3375 (N_3375,In_2961,In_788);
and U3376 (N_3376,In_640,In_419);
and U3377 (N_3377,In_2242,In_1793);
xor U3378 (N_3378,In_486,In_234);
xnor U3379 (N_3379,In_37,In_2803);
nor U3380 (N_3380,In_1672,In_1892);
xor U3381 (N_3381,In_2023,In_2715);
xnor U3382 (N_3382,In_647,In_1313);
and U3383 (N_3383,In_2845,In_2412);
or U3384 (N_3384,In_1062,In_2263);
or U3385 (N_3385,In_2841,In_65);
xor U3386 (N_3386,In_266,In_1934);
or U3387 (N_3387,In_1932,In_339);
nor U3388 (N_3388,In_2941,In_460);
nand U3389 (N_3389,In_56,In_2193);
nor U3390 (N_3390,In_934,In_1783);
xor U3391 (N_3391,In_1631,In_2423);
xor U3392 (N_3392,In_141,In_259);
xnor U3393 (N_3393,In_2185,In_2038);
xnor U3394 (N_3394,In_1501,In_61);
xnor U3395 (N_3395,In_2763,In_1152);
nor U3396 (N_3396,In_2526,In_458);
or U3397 (N_3397,In_916,In_2533);
or U3398 (N_3398,In_1702,In_1155);
nor U3399 (N_3399,In_2574,In_1981);
or U3400 (N_3400,In_2698,In_403);
and U3401 (N_3401,In_189,In_2858);
and U3402 (N_3402,In_229,In_257);
xor U3403 (N_3403,In_1614,In_2894);
and U3404 (N_3404,In_2629,In_334);
xor U3405 (N_3405,In_629,In_1525);
xor U3406 (N_3406,In_481,In_523);
xnor U3407 (N_3407,In_1780,In_213);
or U3408 (N_3408,In_2500,In_256);
xor U3409 (N_3409,In_1658,In_2953);
nand U3410 (N_3410,In_1035,In_2896);
and U3411 (N_3411,In_8,In_889);
or U3412 (N_3412,In_2794,In_700);
xor U3413 (N_3413,In_985,In_2984);
nor U3414 (N_3414,In_529,In_1109);
nand U3415 (N_3415,In_777,In_2542);
or U3416 (N_3416,In_255,In_1516);
or U3417 (N_3417,In_1639,In_1570);
and U3418 (N_3418,In_448,In_2148);
nand U3419 (N_3419,In_29,In_1794);
and U3420 (N_3420,In_34,In_2868);
and U3421 (N_3421,In_1334,In_2885);
xor U3422 (N_3422,In_1979,In_573);
and U3423 (N_3423,In_2522,In_1529);
nor U3424 (N_3424,In_2336,In_1858);
and U3425 (N_3425,In_2149,In_942);
nor U3426 (N_3426,In_689,In_979);
xnor U3427 (N_3427,In_2943,In_2114);
nor U3428 (N_3428,In_2713,In_283);
or U3429 (N_3429,In_2216,In_2872);
and U3430 (N_3430,In_552,In_586);
or U3431 (N_3431,In_1319,In_726);
xor U3432 (N_3432,In_2332,In_2677);
nand U3433 (N_3433,In_1388,In_2206);
or U3434 (N_3434,In_1999,In_658);
and U3435 (N_3435,In_1720,In_2946);
nand U3436 (N_3436,In_161,In_1483);
nand U3437 (N_3437,In_544,In_768);
nand U3438 (N_3438,In_432,In_2446);
nand U3439 (N_3439,In_1589,In_2526);
and U3440 (N_3440,In_2771,In_1422);
xor U3441 (N_3441,In_1890,In_1730);
or U3442 (N_3442,In_686,In_320);
and U3443 (N_3443,In_583,In_288);
and U3444 (N_3444,In_676,In_316);
and U3445 (N_3445,In_2628,In_503);
nor U3446 (N_3446,In_2312,In_884);
xnor U3447 (N_3447,In_2750,In_2680);
nor U3448 (N_3448,In_805,In_1367);
or U3449 (N_3449,In_740,In_2126);
or U3450 (N_3450,In_326,In_2396);
and U3451 (N_3451,In_565,In_354);
nor U3452 (N_3452,In_2948,In_1697);
or U3453 (N_3453,In_643,In_653);
nand U3454 (N_3454,In_1091,In_1373);
nor U3455 (N_3455,In_1414,In_2710);
and U3456 (N_3456,In_796,In_2347);
and U3457 (N_3457,In_1540,In_2013);
and U3458 (N_3458,In_2355,In_249);
or U3459 (N_3459,In_1677,In_2436);
xor U3460 (N_3460,In_2763,In_2605);
or U3461 (N_3461,In_2238,In_2404);
and U3462 (N_3462,In_162,In_2986);
nor U3463 (N_3463,In_2488,In_254);
xnor U3464 (N_3464,In_960,In_1929);
and U3465 (N_3465,In_1806,In_2938);
nand U3466 (N_3466,In_2823,In_1618);
or U3467 (N_3467,In_433,In_1593);
and U3468 (N_3468,In_2839,In_521);
or U3469 (N_3469,In_2290,In_2317);
and U3470 (N_3470,In_1690,In_1428);
xnor U3471 (N_3471,In_906,In_2226);
or U3472 (N_3472,In_1936,In_2255);
and U3473 (N_3473,In_133,In_425);
or U3474 (N_3474,In_1918,In_838);
nor U3475 (N_3475,In_1215,In_2073);
or U3476 (N_3476,In_2720,In_553);
xnor U3477 (N_3477,In_54,In_1963);
nor U3478 (N_3478,In_210,In_2505);
xor U3479 (N_3479,In_2515,In_1084);
nor U3480 (N_3480,In_2439,In_89);
or U3481 (N_3481,In_1175,In_590);
or U3482 (N_3482,In_441,In_415);
nor U3483 (N_3483,In_2904,In_288);
and U3484 (N_3484,In_1741,In_479);
nand U3485 (N_3485,In_462,In_88);
nor U3486 (N_3486,In_1984,In_570);
nor U3487 (N_3487,In_1078,In_712);
or U3488 (N_3488,In_2008,In_1638);
nand U3489 (N_3489,In_711,In_1370);
nand U3490 (N_3490,In_680,In_762);
nand U3491 (N_3491,In_1454,In_289);
nand U3492 (N_3492,In_2865,In_1651);
nand U3493 (N_3493,In_1281,In_368);
nor U3494 (N_3494,In_2896,In_1623);
and U3495 (N_3495,In_2063,In_843);
or U3496 (N_3496,In_1568,In_2993);
xor U3497 (N_3497,In_1629,In_337);
nand U3498 (N_3498,In_437,In_1103);
xnor U3499 (N_3499,In_1646,In_1781);
and U3500 (N_3500,In_1015,In_520);
nor U3501 (N_3501,In_1677,In_113);
nand U3502 (N_3502,In_1642,In_2150);
nor U3503 (N_3503,In_2558,In_320);
xor U3504 (N_3504,In_1297,In_858);
xor U3505 (N_3505,In_1125,In_2106);
or U3506 (N_3506,In_165,In_1761);
and U3507 (N_3507,In_2158,In_2951);
nor U3508 (N_3508,In_2279,In_2180);
xor U3509 (N_3509,In_950,In_5);
nand U3510 (N_3510,In_2286,In_2956);
nor U3511 (N_3511,In_2378,In_1963);
nand U3512 (N_3512,In_1398,In_1620);
or U3513 (N_3513,In_736,In_1580);
or U3514 (N_3514,In_2456,In_2486);
and U3515 (N_3515,In_10,In_1479);
nand U3516 (N_3516,In_1723,In_2186);
and U3517 (N_3517,In_488,In_1116);
nand U3518 (N_3518,In_2233,In_1328);
xor U3519 (N_3519,In_2136,In_683);
xnor U3520 (N_3520,In_348,In_1442);
nor U3521 (N_3521,In_1145,In_1267);
or U3522 (N_3522,In_1715,In_277);
and U3523 (N_3523,In_368,In_2423);
xnor U3524 (N_3524,In_1180,In_2371);
xor U3525 (N_3525,In_580,In_961);
or U3526 (N_3526,In_1986,In_1559);
nor U3527 (N_3527,In_1176,In_1634);
xnor U3528 (N_3528,In_2607,In_631);
xor U3529 (N_3529,In_1116,In_894);
nand U3530 (N_3530,In_2569,In_2388);
nand U3531 (N_3531,In_1374,In_1867);
nand U3532 (N_3532,In_809,In_795);
nand U3533 (N_3533,In_4,In_2581);
and U3534 (N_3534,In_2166,In_422);
nor U3535 (N_3535,In_1148,In_2770);
and U3536 (N_3536,In_1980,In_1105);
nand U3537 (N_3537,In_2630,In_1092);
nand U3538 (N_3538,In_2914,In_495);
xnor U3539 (N_3539,In_1485,In_179);
and U3540 (N_3540,In_493,In_853);
and U3541 (N_3541,In_523,In_914);
xnor U3542 (N_3542,In_2266,In_1683);
nand U3543 (N_3543,In_53,In_1239);
and U3544 (N_3544,In_887,In_2722);
nor U3545 (N_3545,In_1293,In_1588);
xor U3546 (N_3546,In_45,In_2224);
or U3547 (N_3547,In_2932,In_1643);
nand U3548 (N_3548,In_925,In_843);
nor U3549 (N_3549,In_653,In_2589);
nand U3550 (N_3550,In_1428,In_77);
and U3551 (N_3551,In_23,In_2105);
nor U3552 (N_3552,In_742,In_769);
and U3553 (N_3553,In_1507,In_314);
or U3554 (N_3554,In_575,In_2399);
or U3555 (N_3555,In_1075,In_2184);
or U3556 (N_3556,In_434,In_1965);
nand U3557 (N_3557,In_2270,In_2714);
nor U3558 (N_3558,In_305,In_1496);
and U3559 (N_3559,In_659,In_2302);
xor U3560 (N_3560,In_963,In_576);
and U3561 (N_3561,In_1949,In_108);
nor U3562 (N_3562,In_2069,In_2622);
or U3563 (N_3563,In_2567,In_2745);
or U3564 (N_3564,In_263,In_2740);
xnor U3565 (N_3565,In_426,In_742);
nand U3566 (N_3566,In_293,In_78);
and U3567 (N_3567,In_506,In_2273);
and U3568 (N_3568,In_2510,In_1502);
or U3569 (N_3569,In_1665,In_2497);
or U3570 (N_3570,In_2102,In_154);
and U3571 (N_3571,In_1085,In_1399);
xnor U3572 (N_3572,In_1760,In_2332);
xor U3573 (N_3573,In_2641,In_1511);
nand U3574 (N_3574,In_826,In_16);
xnor U3575 (N_3575,In_1817,In_1162);
nand U3576 (N_3576,In_469,In_324);
and U3577 (N_3577,In_1167,In_1660);
or U3578 (N_3578,In_292,In_1106);
xor U3579 (N_3579,In_2752,In_2999);
xor U3580 (N_3580,In_2344,In_1383);
xor U3581 (N_3581,In_1325,In_694);
or U3582 (N_3582,In_2039,In_2506);
nand U3583 (N_3583,In_2079,In_1739);
and U3584 (N_3584,In_1334,In_631);
and U3585 (N_3585,In_2059,In_577);
and U3586 (N_3586,In_1912,In_834);
or U3587 (N_3587,In_265,In_2986);
nor U3588 (N_3588,In_448,In_2284);
or U3589 (N_3589,In_1836,In_1068);
xor U3590 (N_3590,In_1195,In_1426);
and U3591 (N_3591,In_1788,In_2853);
nand U3592 (N_3592,In_1750,In_950);
and U3593 (N_3593,In_2761,In_1160);
nand U3594 (N_3594,In_1562,In_1109);
nand U3595 (N_3595,In_944,In_2781);
or U3596 (N_3596,In_535,In_1724);
nor U3597 (N_3597,In_1166,In_243);
xor U3598 (N_3598,In_632,In_2843);
xor U3599 (N_3599,In_2361,In_404);
nor U3600 (N_3600,In_1809,In_1233);
or U3601 (N_3601,In_2233,In_1642);
nor U3602 (N_3602,In_2765,In_709);
or U3603 (N_3603,In_2072,In_2308);
xor U3604 (N_3604,In_2727,In_2193);
xnor U3605 (N_3605,In_1053,In_560);
nand U3606 (N_3606,In_310,In_1180);
nand U3607 (N_3607,In_2406,In_897);
nand U3608 (N_3608,In_1975,In_1664);
xnor U3609 (N_3609,In_529,In_2851);
nand U3610 (N_3610,In_1069,In_306);
xor U3611 (N_3611,In_2893,In_755);
or U3612 (N_3612,In_2512,In_1455);
nand U3613 (N_3613,In_733,In_923);
nand U3614 (N_3614,In_2233,In_2299);
and U3615 (N_3615,In_603,In_371);
and U3616 (N_3616,In_2790,In_465);
or U3617 (N_3617,In_2043,In_1744);
and U3618 (N_3618,In_962,In_2682);
nor U3619 (N_3619,In_2000,In_739);
or U3620 (N_3620,In_1995,In_2448);
xor U3621 (N_3621,In_984,In_2108);
xor U3622 (N_3622,In_1415,In_1992);
nand U3623 (N_3623,In_1635,In_1444);
nand U3624 (N_3624,In_251,In_1243);
nand U3625 (N_3625,In_2081,In_2548);
or U3626 (N_3626,In_61,In_1886);
and U3627 (N_3627,In_1778,In_2026);
nor U3628 (N_3628,In_1441,In_1374);
nor U3629 (N_3629,In_2978,In_1724);
and U3630 (N_3630,In_2149,In_2436);
nand U3631 (N_3631,In_2833,In_993);
nand U3632 (N_3632,In_574,In_2585);
nor U3633 (N_3633,In_1232,In_61);
or U3634 (N_3634,In_195,In_754);
nand U3635 (N_3635,In_893,In_1874);
and U3636 (N_3636,In_650,In_800);
or U3637 (N_3637,In_1282,In_1475);
and U3638 (N_3638,In_2428,In_1943);
nor U3639 (N_3639,In_2394,In_524);
or U3640 (N_3640,In_472,In_1165);
nor U3641 (N_3641,In_448,In_2837);
xnor U3642 (N_3642,In_1918,In_1296);
xor U3643 (N_3643,In_1966,In_2189);
nor U3644 (N_3644,In_2106,In_934);
or U3645 (N_3645,In_1258,In_113);
nand U3646 (N_3646,In_2560,In_1591);
nand U3647 (N_3647,In_2220,In_422);
nor U3648 (N_3648,In_846,In_296);
nand U3649 (N_3649,In_1284,In_2631);
and U3650 (N_3650,In_1834,In_394);
nor U3651 (N_3651,In_1992,In_1181);
and U3652 (N_3652,In_523,In_2693);
and U3653 (N_3653,In_1226,In_2581);
and U3654 (N_3654,In_2368,In_866);
nand U3655 (N_3655,In_2211,In_400);
nand U3656 (N_3656,In_1822,In_177);
nor U3657 (N_3657,In_1974,In_2347);
and U3658 (N_3658,In_566,In_91);
nand U3659 (N_3659,In_1205,In_1845);
nand U3660 (N_3660,In_2688,In_344);
nand U3661 (N_3661,In_2239,In_850);
nor U3662 (N_3662,In_2680,In_132);
nand U3663 (N_3663,In_2819,In_1319);
xor U3664 (N_3664,In_2165,In_861);
nor U3665 (N_3665,In_1670,In_206);
xor U3666 (N_3666,In_588,In_2971);
nand U3667 (N_3667,In_2919,In_1350);
xnor U3668 (N_3668,In_1743,In_1027);
xnor U3669 (N_3669,In_271,In_2785);
nand U3670 (N_3670,In_80,In_1690);
nor U3671 (N_3671,In_704,In_1884);
xnor U3672 (N_3672,In_676,In_541);
or U3673 (N_3673,In_2447,In_1486);
or U3674 (N_3674,In_2178,In_2257);
nor U3675 (N_3675,In_2938,In_2559);
or U3676 (N_3676,In_1542,In_1258);
nor U3677 (N_3677,In_2376,In_2056);
nor U3678 (N_3678,In_1953,In_2082);
and U3679 (N_3679,In_2126,In_318);
nand U3680 (N_3680,In_2921,In_771);
and U3681 (N_3681,In_526,In_453);
nand U3682 (N_3682,In_1049,In_792);
xor U3683 (N_3683,In_2608,In_2155);
and U3684 (N_3684,In_622,In_1348);
nor U3685 (N_3685,In_2911,In_769);
or U3686 (N_3686,In_2199,In_2678);
nand U3687 (N_3687,In_536,In_272);
nand U3688 (N_3688,In_978,In_984);
nand U3689 (N_3689,In_1041,In_431);
xor U3690 (N_3690,In_2185,In_443);
nor U3691 (N_3691,In_2363,In_2592);
and U3692 (N_3692,In_259,In_515);
xor U3693 (N_3693,In_2828,In_1582);
and U3694 (N_3694,In_1811,In_2503);
nand U3695 (N_3695,In_2667,In_1799);
and U3696 (N_3696,In_2335,In_299);
nand U3697 (N_3697,In_1620,In_2413);
or U3698 (N_3698,In_976,In_1531);
nand U3699 (N_3699,In_81,In_303);
nand U3700 (N_3700,In_828,In_445);
or U3701 (N_3701,In_398,In_2630);
and U3702 (N_3702,In_1110,In_1941);
or U3703 (N_3703,In_1047,In_2438);
xor U3704 (N_3704,In_2489,In_375);
or U3705 (N_3705,In_2787,In_1010);
nand U3706 (N_3706,In_2623,In_668);
nand U3707 (N_3707,In_983,In_432);
nor U3708 (N_3708,In_837,In_1913);
and U3709 (N_3709,In_1611,In_156);
or U3710 (N_3710,In_1511,In_548);
or U3711 (N_3711,In_2683,In_664);
nand U3712 (N_3712,In_919,In_1790);
nand U3713 (N_3713,In_1268,In_1704);
xor U3714 (N_3714,In_986,In_1055);
xor U3715 (N_3715,In_2973,In_1536);
nand U3716 (N_3716,In_987,In_1362);
nand U3717 (N_3717,In_112,In_559);
nor U3718 (N_3718,In_752,In_2061);
nor U3719 (N_3719,In_2297,In_1452);
nor U3720 (N_3720,In_2262,In_599);
and U3721 (N_3721,In_1121,In_1702);
xor U3722 (N_3722,In_147,In_1055);
and U3723 (N_3723,In_1554,In_1804);
or U3724 (N_3724,In_711,In_4);
nor U3725 (N_3725,In_1632,In_1947);
xor U3726 (N_3726,In_1902,In_441);
nor U3727 (N_3727,In_863,In_1314);
nand U3728 (N_3728,In_793,In_2957);
nor U3729 (N_3729,In_339,In_781);
and U3730 (N_3730,In_1168,In_1776);
or U3731 (N_3731,In_1132,In_1947);
nand U3732 (N_3732,In_27,In_799);
and U3733 (N_3733,In_2411,In_1106);
nand U3734 (N_3734,In_781,In_9);
xnor U3735 (N_3735,In_2859,In_1627);
and U3736 (N_3736,In_2794,In_892);
xor U3737 (N_3737,In_500,In_2801);
nand U3738 (N_3738,In_2977,In_476);
or U3739 (N_3739,In_2624,In_2731);
and U3740 (N_3740,In_68,In_1756);
xor U3741 (N_3741,In_56,In_1390);
nor U3742 (N_3742,In_1339,In_2409);
or U3743 (N_3743,In_718,In_454);
or U3744 (N_3744,In_480,In_936);
xor U3745 (N_3745,In_1105,In_1731);
and U3746 (N_3746,In_1289,In_174);
and U3747 (N_3747,In_2504,In_1195);
or U3748 (N_3748,In_2361,In_193);
nand U3749 (N_3749,In_1941,In_1896);
nand U3750 (N_3750,In_889,In_2264);
xor U3751 (N_3751,In_1484,In_1317);
or U3752 (N_3752,In_996,In_2339);
or U3753 (N_3753,In_204,In_1855);
nor U3754 (N_3754,In_2518,In_249);
nand U3755 (N_3755,In_171,In_2902);
nand U3756 (N_3756,In_17,In_820);
or U3757 (N_3757,In_2724,In_107);
xor U3758 (N_3758,In_2969,In_1916);
nand U3759 (N_3759,In_1637,In_2246);
nand U3760 (N_3760,In_2368,In_1191);
nand U3761 (N_3761,In_2014,In_2788);
nand U3762 (N_3762,In_1117,In_1114);
xor U3763 (N_3763,In_97,In_2068);
xor U3764 (N_3764,In_123,In_209);
or U3765 (N_3765,In_2999,In_894);
nor U3766 (N_3766,In_873,In_2256);
nor U3767 (N_3767,In_1694,In_1038);
and U3768 (N_3768,In_1086,In_2761);
xnor U3769 (N_3769,In_2228,In_923);
nand U3770 (N_3770,In_53,In_1579);
nor U3771 (N_3771,In_2192,In_2514);
nand U3772 (N_3772,In_125,In_2711);
or U3773 (N_3773,In_2416,In_1276);
nand U3774 (N_3774,In_1166,In_1219);
nand U3775 (N_3775,In_2838,In_1870);
or U3776 (N_3776,In_1304,In_1128);
or U3777 (N_3777,In_893,In_877);
nor U3778 (N_3778,In_539,In_1695);
xor U3779 (N_3779,In_1499,In_2889);
nand U3780 (N_3780,In_1759,In_864);
nand U3781 (N_3781,In_1024,In_2143);
xnor U3782 (N_3782,In_426,In_280);
xor U3783 (N_3783,In_564,In_2784);
nand U3784 (N_3784,In_167,In_1398);
and U3785 (N_3785,In_1003,In_1467);
and U3786 (N_3786,In_405,In_590);
or U3787 (N_3787,In_1164,In_385);
xor U3788 (N_3788,In_2589,In_734);
nor U3789 (N_3789,In_30,In_788);
nor U3790 (N_3790,In_413,In_2255);
nor U3791 (N_3791,In_1303,In_2197);
and U3792 (N_3792,In_1283,In_2270);
or U3793 (N_3793,In_2630,In_2478);
or U3794 (N_3794,In_286,In_2984);
nand U3795 (N_3795,In_1264,In_2693);
or U3796 (N_3796,In_875,In_1839);
nor U3797 (N_3797,In_1770,In_2598);
xor U3798 (N_3798,In_1550,In_2780);
nand U3799 (N_3799,In_1627,In_748);
nor U3800 (N_3800,In_1062,In_1012);
nor U3801 (N_3801,In_225,In_2264);
or U3802 (N_3802,In_930,In_797);
and U3803 (N_3803,In_1301,In_2115);
or U3804 (N_3804,In_2211,In_168);
nand U3805 (N_3805,In_2582,In_2156);
nor U3806 (N_3806,In_303,In_695);
xnor U3807 (N_3807,In_1652,In_648);
nand U3808 (N_3808,In_2363,In_501);
nand U3809 (N_3809,In_2352,In_1523);
nor U3810 (N_3810,In_1552,In_502);
nand U3811 (N_3811,In_2436,In_2938);
xnor U3812 (N_3812,In_1160,In_2627);
xor U3813 (N_3813,In_78,In_1523);
and U3814 (N_3814,In_613,In_974);
nand U3815 (N_3815,In_2084,In_791);
xor U3816 (N_3816,In_1861,In_325);
nor U3817 (N_3817,In_1971,In_2575);
xor U3818 (N_3818,In_945,In_1728);
nor U3819 (N_3819,In_453,In_405);
xor U3820 (N_3820,In_626,In_1074);
nand U3821 (N_3821,In_648,In_2794);
xnor U3822 (N_3822,In_1777,In_2772);
nor U3823 (N_3823,In_676,In_988);
or U3824 (N_3824,In_516,In_215);
or U3825 (N_3825,In_2022,In_2368);
xor U3826 (N_3826,In_2945,In_507);
and U3827 (N_3827,In_451,In_2436);
nand U3828 (N_3828,In_2944,In_1243);
and U3829 (N_3829,In_2962,In_423);
xnor U3830 (N_3830,In_2073,In_2295);
nand U3831 (N_3831,In_2109,In_1883);
nand U3832 (N_3832,In_1240,In_747);
xor U3833 (N_3833,In_1870,In_1133);
nand U3834 (N_3834,In_2948,In_1062);
nand U3835 (N_3835,In_1444,In_1918);
nor U3836 (N_3836,In_1417,In_175);
nor U3837 (N_3837,In_1000,In_95);
nor U3838 (N_3838,In_133,In_794);
xnor U3839 (N_3839,In_670,In_1452);
xnor U3840 (N_3840,In_2267,In_1976);
nand U3841 (N_3841,In_367,In_2283);
xor U3842 (N_3842,In_1038,In_2978);
nor U3843 (N_3843,In_1563,In_1245);
nand U3844 (N_3844,In_911,In_1458);
xnor U3845 (N_3845,In_1092,In_2887);
nor U3846 (N_3846,In_2249,In_381);
xor U3847 (N_3847,In_2341,In_1753);
xor U3848 (N_3848,In_2858,In_1824);
nand U3849 (N_3849,In_855,In_1203);
or U3850 (N_3850,In_225,In_1347);
xor U3851 (N_3851,In_2050,In_2547);
or U3852 (N_3852,In_2034,In_2708);
nor U3853 (N_3853,In_1719,In_2766);
nand U3854 (N_3854,In_2016,In_1548);
nor U3855 (N_3855,In_2919,In_1659);
or U3856 (N_3856,In_453,In_1128);
nand U3857 (N_3857,In_1374,In_2992);
nor U3858 (N_3858,In_2524,In_1196);
nor U3859 (N_3859,In_2885,In_2889);
nor U3860 (N_3860,In_1244,In_90);
nor U3861 (N_3861,In_243,In_2365);
xor U3862 (N_3862,In_2727,In_2869);
and U3863 (N_3863,In_334,In_2289);
and U3864 (N_3864,In_2467,In_1280);
xor U3865 (N_3865,In_469,In_2969);
nand U3866 (N_3866,In_283,In_2940);
xnor U3867 (N_3867,In_62,In_2202);
and U3868 (N_3868,In_397,In_514);
xor U3869 (N_3869,In_741,In_542);
and U3870 (N_3870,In_258,In_1018);
nor U3871 (N_3871,In_2204,In_1654);
and U3872 (N_3872,In_2715,In_2846);
xnor U3873 (N_3873,In_326,In_2982);
xnor U3874 (N_3874,In_2321,In_1541);
nor U3875 (N_3875,In_2255,In_2126);
and U3876 (N_3876,In_458,In_2322);
xor U3877 (N_3877,In_1527,In_711);
or U3878 (N_3878,In_1708,In_1778);
nand U3879 (N_3879,In_930,In_1491);
nor U3880 (N_3880,In_860,In_2565);
nor U3881 (N_3881,In_1460,In_1958);
xor U3882 (N_3882,In_920,In_1617);
xor U3883 (N_3883,In_2097,In_501);
or U3884 (N_3884,In_785,In_145);
or U3885 (N_3885,In_1049,In_0);
nand U3886 (N_3886,In_1187,In_481);
and U3887 (N_3887,In_64,In_2457);
nor U3888 (N_3888,In_1948,In_611);
or U3889 (N_3889,In_697,In_2858);
nand U3890 (N_3890,In_2429,In_576);
xnor U3891 (N_3891,In_2493,In_1725);
and U3892 (N_3892,In_2755,In_2401);
or U3893 (N_3893,In_777,In_913);
xor U3894 (N_3894,In_2883,In_678);
and U3895 (N_3895,In_569,In_241);
or U3896 (N_3896,In_2987,In_1312);
xor U3897 (N_3897,In_2713,In_1012);
xor U3898 (N_3898,In_2358,In_2198);
nand U3899 (N_3899,In_1939,In_2943);
xor U3900 (N_3900,In_1215,In_1873);
nand U3901 (N_3901,In_2505,In_2659);
nand U3902 (N_3902,In_1850,In_2792);
or U3903 (N_3903,In_2291,In_1502);
or U3904 (N_3904,In_1503,In_2174);
xnor U3905 (N_3905,In_1716,In_1685);
nor U3906 (N_3906,In_612,In_2339);
and U3907 (N_3907,In_1080,In_1010);
nand U3908 (N_3908,In_2987,In_1595);
nand U3909 (N_3909,In_2705,In_1882);
or U3910 (N_3910,In_2210,In_1191);
xor U3911 (N_3911,In_737,In_918);
nor U3912 (N_3912,In_1002,In_923);
nor U3913 (N_3913,In_2263,In_2840);
and U3914 (N_3914,In_1305,In_1186);
and U3915 (N_3915,In_617,In_1395);
or U3916 (N_3916,In_1058,In_326);
or U3917 (N_3917,In_995,In_2078);
or U3918 (N_3918,In_35,In_854);
xor U3919 (N_3919,In_941,In_130);
xnor U3920 (N_3920,In_1763,In_2724);
and U3921 (N_3921,In_148,In_111);
xnor U3922 (N_3922,In_1445,In_2701);
nand U3923 (N_3923,In_500,In_2944);
nor U3924 (N_3924,In_1624,In_1599);
nor U3925 (N_3925,In_1092,In_110);
xnor U3926 (N_3926,In_2566,In_2280);
nand U3927 (N_3927,In_1717,In_20);
or U3928 (N_3928,In_1200,In_2894);
nor U3929 (N_3929,In_181,In_109);
nand U3930 (N_3930,In_2969,In_1401);
nand U3931 (N_3931,In_1898,In_1216);
nand U3932 (N_3932,In_1711,In_21);
xor U3933 (N_3933,In_1082,In_1771);
nor U3934 (N_3934,In_400,In_2457);
xor U3935 (N_3935,In_2760,In_906);
nand U3936 (N_3936,In_1446,In_2533);
or U3937 (N_3937,In_68,In_325);
and U3938 (N_3938,In_1174,In_2508);
nor U3939 (N_3939,In_2306,In_2541);
xnor U3940 (N_3940,In_577,In_1806);
nand U3941 (N_3941,In_1683,In_714);
nand U3942 (N_3942,In_1872,In_179);
or U3943 (N_3943,In_2736,In_2375);
and U3944 (N_3944,In_1958,In_576);
xor U3945 (N_3945,In_1456,In_472);
nor U3946 (N_3946,In_311,In_649);
nand U3947 (N_3947,In_1391,In_2610);
and U3948 (N_3948,In_952,In_1803);
nor U3949 (N_3949,In_2281,In_2029);
nand U3950 (N_3950,In_1934,In_397);
nand U3951 (N_3951,In_2305,In_1042);
and U3952 (N_3952,In_1769,In_304);
nand U3953 (N_3953,In_2889,In_1448);
nor U3954 (N_3954,In_1793,In_853);
and U3955 (N_3955,In_746,In_251);
and U3956 (N_3956,In_973,In_1622);
nor U3957 (N_3957,In_2969,In_1481);
xnor U3958 (N_3958,In_63,In_2980);
nand U3959 (N_3959,In_1636,In_1792);
nor U3960 (N_3960,In_1275,In_630);
or U3961 (N_3961,In_2585,In_2093);
nor U3962 (N_3962,In_272,In_1470);
nor U3963 (N_3963,In_906,In_1073);
and U3964 (N_3964,In_1049,In_613);
or U3965 (N_3965,In_1652,In_2125);
xnor U3966 (N_3966,In_1575,In_773);
nand U3967 (N_3967,In_6,In_61);
or U3968 (N_3968,In_1811,In_471);
and U3969 (N_3969,In_1864,In_2251);
and U3970 (N_3970,In_320,In_496);
nand U3971 (N_3971,In_39,In_2203);
nor U3972 (N_3972,In_35,In_1582);
nor U3973 (N_3973,In_2181,In_760);
and U3974 (N_3974,In_1920,In_2720);
nand U3975 (N_3975,In_745,In_915);
xor U3976 (N_3976,In_1939,In_887);
nor U3977 (N_3977,In_2552,In_2214);
nand U3978 (N_3978,In_1757,In_122);
and U3979 (N_3979,In_1579,In_1003);
nor U3980 (N_3980,In_2697,In_1901);
nand U3981 (N_3981,In_1507,In_1101);
xor U3982 (N_3982,In_1373,In_259);
or U3983 (N_3983,In_1145,In_457);
nand U3984 (N_3984,In_2259,In_454);
nor U3985 (N_3985,In_1974,In_810);
and U3986 (N_3986,In_1854,In_2788);
nor U3987 (N_3987,In_2674,In_2364);
and U3988 (N_3988,In_1719,In_872);
or U3989 (N_3989,In_2135,In_481);
xor U3990 (N_3990,In_70,In_380);
and U3991 (N_3991,In_1022,In_2270);
xor U3992 (N_3992,In_417,In_1551);
and U3993 (N_3993,In_2527,In_988);
xor U3994 (N_3994,In_1356,In_808);
xor U3995 (N_3995,In_1215,In_500);
nor U3996 (N_3996,In_2980,In_2698);
xor U3997 (N_3997,In_856,In_2372);
or U3998 (N_3998,In_2311,In_2303);
nand U3999 (N_3999,In_1322,In_1363);
and U4000 (N_4000,In_2954,In_1922);
or U4001 (N_4001,In_1749,In_306);
or U4002 (N_4002,In_1897,In_2136);
nand U4003 (N_4003,In_1592,In_2292);
nor U4004 (N_4004,In_2612,In_2635);
or U4005 (N_4005,In_2818,In_267);
nand U4006 (N_4006,In_32,In_1047);
or U4007 (N_4007,In_6,In_1953);
or U4008 (N_4008,In_1333,In_1788);
nor U4009 (N_4009,In_422,In_1449);
or U4010 (N_4010,In_1839,In_19);
and U4011 (N_4011,In_372,In_488);
or U4012 (N_4012,In_2982,In_397);
xnor U4013 (N_4013,In_1883,In_2947);
xor U4014 (N_4014,In_2745,In_2884);
or U4015 (N_4015,In_17,In_83);
nand U4016 (N_4016,In_1935,In_510);
nor U4017 (N_4017,In_1059,In_972);
nor U4018 (N_4018,In_525,In_1585);
nand U4019 (N_4019,In_1817,In_1461);
nand U4020 (N_4020,In_52,In_2648);
nor U4021 (N_4021,In_2419,In_1399);
or U4022 (N_4022,In_2684,In_1795);
and U4023 (N_4023,In_49,In_2168);
or U4024 (N_4024,In_1347,In_100);
nor U4025 (N_4025,In_619,In_443);
xor U4026 (N_4026,In_2478,In_11);
nor U4027 (N_4027,In_132,In_2807);
nor U4028 (N_4028,In_1189,In_1519);
nand U4029 (N_4029,In_2606,In_2785);
nor U4030 (N_4030,In_2445,In_8);
nor U4031 (N_4031,In_960,In_376);
and U4032 (N_4032,In_1321,In_1784);
xnor U4033 (N_4033,In_2357,In_557);
and U4034 (N_4034,In_2240,In_294);
nand U4035 (N_4035,In_418,In_386);
nor U4036 (N_4036,In_980,In_2097);
and U4037 (N_4037,In_2504,In_575);
or U4038 (N_4038,In_2027,In_2023);
and U4039 (N_4039,In_129,In_2303);
nor U4040 (N_4040,In_2147,In_1245);
and U4041 (N_4041,In_2815,In_1203);
nor U4042 (N_4042,In_2706,In_2810);
or U4043 (N_4043,In_1317,In_2049);
nor U4044 (N_4044,In_1245,In_210);
and U4045 (N_4045,In_1094,In_176);
nor U4046 (N_4046,In_178,In_1345);
or U4047 (N_4047,In_2446,In_2787);
nor U4048 (N_4048,In_2012,In_396);
and U4049 (N_4049,In_1019,In_2167);
or U4050 (N_4050,In_539,In_1203);
and U4051 (N_4051,In_1077,In_2462);
xnor U4052 (N_4052,In_922,In_2459);
xor U4053 (N_4053,In_2251,In_2203);
nor U4054 (N_4054,In_780,In_274);
nor U4055 (N_4055,In_12,In_356);
nor U4056 (N_4056,In_2172,In_22);
or U4057 (N_4057,In_320,In_2614);
nor U4058 (N_4058,In_254,In_2443);
nor U4059 (N_4059,In_575,In_2052);
and U4060 (N_4060,In_617,In_1588);
and U4061 (N_4061,In_2246,In_1653);
nor U4062 (N_4062,In_1893,In_2148);
or U4063 (N_4063,In_749,In_2120);
xnor U4064 (N_4064,In_190,In_2464);
nand U4065 (N_4065,In_2617,In_418);
and U4066 (N_4066,In_2540,In_451);
nor U4067 (N_4067,In_664,In_278);
xor U4068 (N_4068,In_1613,In_1205);
or U4069 (N_4069,In_2856,In_2923);
nor U4070 (N_4070,In_1006,In_141);
and U4071 (N_4071,In_449,In_220);
and U4072 (N_4072,In_2723,In_1855);
or U4073 (N_4073,In_2282,In_1933);
and U4074 (N_4074,In_2206,In_1348);
nand U4075 (N_4075,In_2712,In_2765);
nand U4076 (N_4076,In_2217,In_947);
nor U4077 (N_4077,In_1055,In_2545);
or U4078 (N_4078,In_342,In_2281);
or U4079 (N_4079,In_121,In_484);
nor U4080 (N_4080,In_1696,In_1443);
nand U4081 (N_4081,In_1449,In_1408);
and U4082 (N_4082,In_940,In_402);
nand U4083 (N_4083,In_1851,In_42);
and U4084 (N_4084,In_1122,In_2849);
or U4085 (N_4085,In_2374,In_2856);
or U4086 (N_4086,In_2505,In_170);
and U4087 (N_4087,In_1597,In_1113);
or U4088 (N_4088,In_718,In_1138);
xor U4089 (N_4089,In_1082,In_660);
and U4090 (N_4090,In_1943,In_2711);
or U4091 (N_4091,In_1433,In_2782);
nand U4092 (N_4092,In_2912,In_2567);
xnor U4093 (N_4093,In_2995,In_2737);
or U4094 (N_4094,In_2035,In_1376);
and U4095 (N_4095,In_1604,In_1148);
nand U4096 (N_4096,In_1800,In_1537);
nor U4097 (N_4097,In_597,In_1313);
or U4098 (N_4098,In_2959,In_899);
nor U4099 (N_4099,In_2416,In_20);
nand U4100 (N_4100,In_1554,In_1043);
and U4101 (N_4101,In_121,In_2879);
nand U4102 (N_4102,In_1974,In_275);
nand U4103 (N_4103,In_1545,In_246);
nor U4104 (N_4104,In_2429,In_279);
xor U4105 (N_4105,In_2326,In_674);
and U4106 (N_4106,In_2808,In_2860);
and U4107 (N_4107,In_931,In_60);
nor U4108 (N_4108,In_2917,In_2439);
and U4109 (N_4109,In_89,In_1642);
or U4110 (N_4110,In_2231,In_761);
or U4111 (N_4111,In_2910,In_2669);
nor U4112 (N_4112,In_2146,In_1855);
nor U4113 (N_4113,In_590,In_2589);
xor U4114 (N_4114,In_626,In_2402);
nor U4115 (N_4115,In_28,In_307);
nand U4116 (N_4116,In_1177,In_2831);
and U4117 (N_4117,In_234,In_1978);
or U4118 (N_4118,In_1038,In_13);
or U4119 (N_4119,In_578,In_1371);
or U4120 (N_4120,In_66,In_2994);
or U4121 (N_4121,In_2655,In_629);
and U4122 (N_4122,In_1808,In_2656);
or U4123 (N_4123,In_340,In_2752);
and U4124 (N_4124,In_1067,In_1531);
nor U4125 (N_4125,In_1691,In_496);
and U4126 (N_4126,In_2757,In_69);
nand U4127 (N_4127,In_670,In_1144);
and U4128 (N_4128,In_1316,In_2071);
nand U4129 (N_4129,In_1330,In_1141);
nand U4130 (N_4130,In_24,In_116);
xor U4131 (N_4131,In_935,In_499);
or U4132 (N_4132,In_2010,In_467);
and U4133 (N_4133,In_2889,In_1699);
xnor U4134 (N_4134,In_2462,In_982);
nand U4135 (N_4135,In_2204,In_623);
xor U4136 (N_4136,In_2077,In_97);
xnor U4137 (N_4137,In_2247,In_2958);
xnor U4138 (N_4138,In_843,In_1706);
or U4139 (N_4139,In_381,In_2578);
and U4140 (N_4140,In_353,In_1326);
or U4141 (N_4141,In_891,In_2212);
nand U4142 (N_4142,In_567,In_2277);
or U4143 (N_4143,In_365,In_1257);
nand U4144 (N_4144,In_1889,In_1583);
and U4145 (N_4145,In_997,In_967);
or U4146 (N_4146,In_2741,In_1355);
xor U4147 (N_4147,In_2182,In_1107);
nor U4148 (N_4148,In_2351,In_2190);
nand U4149 (N_4149,In_178,In_2125);
nand U4150 (N_4150,In_2473,In_173);
nor U4151 (N_4151,In_1746,In_446);
or U4152 (N_4152,In_420,In_2209);
or U4153 (N_4153,In_1872,In_1645);
or U4154 (N_4154,In_1142,In_1015);
nor U4155 (N_4155,In_1408,In_437);
and U4156 (N_4156,In_1385,In_964);
or U4157 (N_4157,In_7,In_352);
xor U4158 (N_4158,In_338,In_979);
nand U4159 (N_4159,In_704,In_1408);
or U4160 (N_4160,In_618,In_1313);
nor U4161 (N_4161,In_203,In_2753);
and U4162 (N_4162,In_1670,In_1960);
xnor U4163 (N_4163,In_2194,In_302);
nor U4164 (N_4164,In_660,In_1746);
nand U4165 (N_4165,In_2338,In_291);
xor U4166 (N_4166,In_1966,In_2139);
or U4167 (N_4167,In_120,In_405);
and U4168 (N_4168,In_2366,In_1628);
nand U4169 (N_4169,In_1407,In_1500);
xnor U4170 (N_4170,In_2703,In_833);
or U4171 (N_4171,In_826,In_2799);
or U4172 (N_4172,In_945,In_2952);
nand U4173 (N_4173,In_2540,In_2334);
and U4174 (N_4174,In_2258,In_1578);
or U4175 (N_4175,In_1452,In_1825);
and U4176 (N_4176,In_90,In_322);
or U4177 (N_4177,In_2151,In_2806);
xnor U4178 (N_4178,In_2945,In_729);
xnor U4179 (N_4179,In_344,In_2250);
xor U4180 (N_4180,In_2972,In_1332);
nor U4181 (N_4181,In_2773,In_719);
nor U4182 (N_4182,In_469,In_1701);
and U4183 (N_4183,In_456,In_744);
and U4184 (N_4184,In_2272,In_2176);
nor U4185 (N_4185,In_2481,In_1739);
xnor U4186 (N_4186,In_2300,In_2757);
xnor U4187 (N_4187,In_715,In_1698);
and U4188 (N_4188,In_2407,In_2426);
or U4189 (N_4189,In_1726,In_2148);
nand U4190 (N_4190,In_1285,In_354);
or U4191 (N_4191,In_2421,In_848);
xor U4192 (N_4192,In_2503,In_1767);
xnor U4193 (N_4193,In_2501,In_1891);
xnor U4194 (N_4194,In_1184,In_2477);
nand U4195 (N_4195,In_2761,In_1124);
nor U4196 (N_4196,In_605,In_2110);
and U4197 (N_4197,In_1703,In_1637);
or U4198 (N_4198,In_112,In_927);
nor U4199 (N_4199,In_126,In_2540);
or U4200 (N_4200,In_90,In_1829);
nand U4201 (N_4201,In_2638,In_551);
nand U4202 (N_4202,In_2677,In_644);
nor U4203 (N_4203,In_1272,In_2619);
and U4204 (N_4204,In_666,In_1375);
and U4205 (N_4205,In_2938,In_430);
or U4206 (N_4206,In_1978,In_1032);
and U4207 (N_4207,In_2128,In_724);
xor U4208 (N_4208,In_2297,In_357);
nand U4209 (N_4209,In_2447,In_258);
and U4210 (N_4210,In_2243,In_589);
and U4211 (N_4211,In_1134,In_858);
nand U4212 (N_4212,In_402,In_1904);
xor U4213 (N_4213,In_2355,In_1445);
and U4214 (N_4214,In_1509,In_1715);
and U4215 (N_4215,In_2789,In_2179);
nand U4216 (N_4216,In_327,In_2709);
and U4217 (N_4217,In_1660,In_2429);
nor U4218 (N_4218,In_2061,In_160);
nor U4219 (N_4219,In_1672,In_532);
nand U4220 (N_4220,In_1160,In_1919);
nand U4221 (N_4221,In_1577,In_1181);
and U4222 (N_4222,In_1843,In_2568);
or U4223 (N_4223,In_769,In_1188);
and U4224 (N_4224,In_104,In_2262);
or U4225 (N_4225,In_922,In_2874);
nand U4226 (N_4226,In_152,In_2010);
nor U4227 (N_4227,In_746,In_1148);
and U4228 (N_4228,In_2011,In_2706);
or U4229 (N_4229,In_2362,In_2075);
xnor U4230 (N_4230,In_2042,In_346);
nand U4231 (N_4231,In_1907,In_2918);
xnor U4232 (N_4232,In_1940,In_872);
and U4233 (N_4233,In_2469,In_2583);
xnor U4234 (N_4234,In_833,In_2630);
xor U4235 (N_4235,In_674,In_1688);
and U4236 (N_4236,In_288,In_1629);
and U4237 (N_4237,In_2647,In_2485);
and U4238 (N_4238,In_2506,In_2896);
nand U4239 (N_4239,In_743,In_1477);
and U4240 (N_4240,In_2407,In_2601);
nand U4241 (N_4241,In_479,In_640);
or U4242 (N_4242,In_1446,In_1532);
xor U4243 (N_4243,In_2793,In_1814);
or U4244 (N_4244,In_2444,In_2072);
nand U4245 (N_4245,In_194,In_794);
nor U4246 (N_4246,In_1526,In_763);
nor U4247 (N_4247,In_67,In_984);
and U4248 (N_4248,In_880,In_1575);
xnor U4249 (N_4249,In_683,In_10);
or U4250 (N_4250,In_1074,In_1503);
or U4251 (N_4251,In_74,In_1537);
xnor U4252 (N_4252,In_1911,In_2833);
xnor U4253 (N_4253,In_1798,In_1475);
xor U4254 (N_4254,In_555,In_2837);
xor U4255 (N_4255,In_2684,In_895);
nor U4256 (N_4256,In_1042,In_145);
xor U4257 (N_4257,In_478,In_507);
nor U4258 (N_4258,In_1295,In_1426);
xnor U4259 (N_4259,In_571,In_1761);
and U4260 (N_4260,In_1062,In_1162);
and U4261 (N_4261,In_1769,In_416);
nor U4262 (N_4262,In_1176,In_1135);
and U4263 (N_4263,In_1466,In_843);
nand U4264 (N_4264,In_2601,In_1526);
or U4265 (N_4265,In_1111,In_956);
xnor U4266 (N_4266,In_465,In_397);
and U4267 (N_4267,In_102,In_2125);
nand U4268 (N_4268,In_2893,In_1453);
and U4269 (N_4269,In_2214,In_1456);
or U4270 (N_4270,In_582,In_2513);
nor U4271 (N_4271,In_2381,In_2498);
xor U4272 (N_4272,In_1134,In_217);
xnor U4273 (N_4273,In_1655,In_821);
xor U4274 (N_4274,In_1218,In_2623);
nor U4275 (N_4275,In_2646,In_1513);
nor U4276 (N_4276,In_1866,In_2835);
or U4277 (N_4277,In_1764,In_378);
or U4278 (N_4278,In_2063,In_1218);
nand U4279 (N_4279,In_13,In_563);
or U4280 (N_4280,In_2554,In_2886);
xor U4281 (N_4281,In_738,In_2097);
nand U4282 (N_4282,In_2966,In_2482);
or U4283 (N_4283,In_2808,In_2657);
and U4284 (N_4284,In_1370,In_2313);
nand U4285 (N_4285,In_1122,In_1267);
nor U4286 (N_4286,In_1992,In_55);
and U4287 (N_4287,In_2170,In_82);
xnor U4288 (N_4288,In_169,In_2656);
xnor U4289 (N_4289,In_2501,In_877);
and U4290 (N_4290,In_1820,In_1325);
nor U4291 (N_4291,In_1589,In_2036);
xnor U4292 (N_4292,In_2070,In_2802);
nor U4293 (N_4293,In_1596,In_1721);
and U4294 (N_4294,In_949,In_809);
and U4295 (N_4295,In_2371,In_2488);
or U4296 (N_4296,In_752,In_2658);
nand U4297 (N_4297,In_2993,In_2005);
nor U4298 (N_4298,In_2040,In_252);
and U4299 (N_4299,In_2,In_1312);
xor U4300 (N_4300,In_985,In_2806);
or U4301 (N_4301,In_2973,In_1369);
nor U4302 (N_4302,In_1434,In_664);
xnor U4303 (N_4303,In_1255,In_2476);
and U4304 (N_4304,In_1565,In_2985);
nor U4305 (N_4305,In_805,In_338);
nor U4306 (N_4306,In_2847,In_2284);
or U4307 (N_4307,In_2416,In_1149);
or U4308 (N_4308,In_2714,In_884);
and U4309 (N_4309,In_871,In_179);
or U4310 (N_4310,In_745,In_5);
xnor U4311 (N_4311,In_2404,In_1504);
xnor U4312 (N_4312,In_2224,In_100);
xor U4313 (N_4313,In_2945,In_699);
or U4314 (N_4314,In_519,In_577);
xor U4315 (N_4315,In_1615,In_1579);
and U4316 (N_4316,In_1184,In_2274);
nand U4317 (N_4317,In_417,In_2509);
and U4318 (N_4318,In_1764,In_2195);
and U4319 (N_4319,In_1383,In_1572);
nor U4320 (N_4320,In_1096,In_1737);
xor U4321 (N_4321,In_2510,In_130);
or U4322 (N_4322,In_1477,In_1506);
nand U4323 (N_4323,In_1299,In_20);
xor U4324 (N_4324,In_1001,In_1390);
xor U4325 (N_4325,In_2651,In_1315);
nand U4326 (N_4326,In_3,In_1865);
or U4327 (N_4327,In_30,In_1204);
xnor U4328 (N_4328,In_31,In_1829);
nor U4329 (N_4329,In_2167,In_2216);
nor U4330 (N_4330,In_2644,In_2913);
nand U4331 (N_4331,In_2912,In_2723);
xnor U4332 (N_4332,In_1555,In_821);
and U4333 (N_4333,In_1694,In_20);
and U4334 (N_4334,In_186,In_1466);
nor U4335 (N_4335,In_1577,In_1740);
nand U4336 (N_4336,In_170,In_2374);
nand U4337 (N_4337,In_2360,In_2904);
or U4338 (N_4338,In_1008,In_2933);
nand U4339 (N_4339,In_1208,In_752);
xnor U4340 (N_4340,In_917,In_2970);
nor U4341 (N_4341,In_1699,In_118);
xor U4342 (N_4342,In_2810,In_2374);
xor U4343 (N_4343,In_1627,In_2634);
or U4344 (N_4344,In_1188,In_1340);
xor U4345 (N_4345,In_237,In_2965);
and U4346 (N_4346,In_214,In_588);
and U4347 (N_4347,In_984,In_2064);
nand U4348 (N_4348,In_174,In_2161);
nor U4349 (N_4349,In_102,In_1072);
or U4350 (N_4350,In_2826,In_2117);
or U4351 (N_4351,In_2880,In_2368);
nor U4352 (N_4352,In_1770,In_160);
and U4353 (N_4353,In_1539,In_1796);
xnor U4354 (N_4354,In_757,In_2327);
xnor U4355 (N_4355,In_1304,In_1992);
nand U4356 (N_4356,In_2329,In_115);
and U4357 (N_4357,In_1515,In_2174);
and U4358 (N_4358,In_2138,In_723);
nand U4359 (N_4359,In_2274,In_970);
nor U4360 (N_4360,In_2414,In_2610);
nor U4361 (N_4361,In_2318,In_1067);
and U4362 (N_4362,In_1177,In_916);
nor U4363 (N_4363,In_1106,In_1563);
and U4364 (N_4364,In_409,In_548);
nand U4365 (N_4365,In_2141,In_1139);
and U4366 (N_4366,In_579,In_1237);
nor U4367 (N_4367,In_2455,In_637);
xor U4368 (N_4368,In_2036,In_2081);
nor U4369 (N_4369,In_1929,In_836);
and U4370 (N_4370,In_1408,In_2078);
nor U4371 (N_4371,In_1175,In_2337);
xnor U4372 (N_4372,In_37,In_310);
and U4373 (N_4373,In_1125,In_1958);
and U4374 (N_4374,In_2908,In_1306);
and U4375 (N_4375,In_662,In_2590);
nor U4376 (N_4376,In_773,In_527);
and U4377 (N_4377,In_2266,In_2723);
xnor U4378 (N_4378,In_485,In_2644);
and U4379 (N_4379,In_952,In_2512);
and U4380 (N_4380,In_2505,In_1139);
and U4381 (N_4381,In_2976,In_2907);
nand U4382 (N_4382,In_1368,In_483);
nand U4383 (N_4383,In_2356,In_483);
xor U4384 (N_4384,In_733,In_1604);
xor U4385 (N_4385,In_1759,In_1101);
and U4386 (N_4386,In_1092,In_609);
and U4387 (N_4387,In_629,In_96);
xor U4388 (N_4388,In_1091,In_599);
xnor U4389 (N_4389,In_1603,In_2101);
nand U4390 (N_4390,In_2817,In_2727);
or U4391 (N_4391,In_1446,In_2976);
nand U4392 (N_4392,In_1323,In_1026);
and U4393 (N_4393,In_125,In_275);
nor U4394 (N_4394,In_1632,In_1516);
and U4395 (N_4395,In_2852,In_2757);
nor U4396 (N_4396,In_2679,In_1893);
and U4397 (N_4397,In_1899,In_2461);
nor U4398 (N_4398,In_156,In_691);
xnor U4399 (N_4399,In_1689,In_2248);
nand U4400 (N_4400,In_2966,In_2550);
and U4401 (N_4401,In_2946,In_1601);
nor U4402 (N_4402,In_1781,In_2265);
nor U4403 (N_4403,In_2006,In_2051);
nor U4404 (N_4404,In_1455,In_2073);
nor U4405 (N_4405,In_2123,In_1871);
and U4406 (N_4406,In_839,In_602);
or U4407 (N_4407,In_2544,In_2783);
and U4408 (N_4408,In_1910,In_1068);
nor U4409 (N_4409,In_1043,In_1244);
and U4410 (N_4410,In_961,In_181);
nor U4411 (N_4411,In_551,In_1056);
nor U4412 (N_4412,In_661,In_2837);
or U4413 (N_4413,In_1101,In_2014);
nor U4414 (N_4414,In_1054,In_2497);
nand U4415 (N_4415,In_2480,In_1045);
nand U4416 (N_4416,In_153,In_1556);
and U4417 (N_4417,In_1028,In_2357);
or U4418 (N_4418,In_72,In_222);
or U4419 (N_4419,In_527,In_1532);
nor U4420 (N_4420,In_1548,In_791);
nor U4421 (N_4421,In_961,In_2598);
nand U4422 (N_4422,In_832,In_2528);
or U4423 (N_4423,In_2894,In_1130);
nand U4424 (N_4424,In_1393,In_431);
xor U4425 (N_4425,In_227,In_981);
nand U4426 (N_4426,In_199,In_2776);
nor U4427 (N_4427,In_1291,In_2503);
nor U4428 (N_4428,In_1394,In_2229);
or U4429 (N_4429,In_1696,In_471);
or U4430 (N_4430,In_1068,In_731);
and U4431 (N_4431,In_93,In_2787);
nand U4432 (N_4432,In_354,In_2526);
nor U4433 (N_4433,In_1090,In_2374);
or U4434 (N_4434,In_2654,In_459);
or U4435 (N_4435,In_2245,In_2285);
and U4436 (N_4436,In_2045,In_1022);
or U4437 (N_4437,In_2891,In_852);
and U4438 (N_4438,In_252,In_2832);
and U4439 (N_4439,In_384,In_2327);
xor U4440 (N_4440,In_2602,In_1480);
or U4441 (N_4441,In_1901,In_2749);
xnor U4442 (N_4442,In_46,In_1877);
or U4443 (N_4443,In_2778,In_1574);
and U4444 (N_4444,In_2889,In_2824);
or U4445 (N_4445,In_988,In_699);
and U4446 (N_4446,In_1321,In_660);
nor U4447 (N_4447,In_1312,In_199);
xor U4448 (N_4448,In_2254,In_295);
or U4449 (N_4449,In_731,In_510);
nand U4450 (N_4450,In_1162,In_2226);
nor U4451 (N_4451,In_1575,In_2614);
nand U4452 (N_4452,In_855,In_1560);
xnor U4453 (N_4453,In_1489,In_141);
nor U4454 (N_4454,In_2908,In_873);
nand U4455 (N_4455,In_365,In_314);
or U4456 (N_4456,In_1602,In_1890);
and U4457 (N_4457,In_484,In_2308);
or U4458 (N_4458,In_411,In_2760);
or U4459 (N_4459,In_1813,In_1120);
and U4460 (N_4460,In_2960,In_2516);
xnor U4461 (N_4461,In_824,In_2945);
nand U4462 (N_4462,In_366,In_37);
or U4463 (N_4463,In_2334,In_447);
xor U4464 (N_4464,In_571,In_1847);
nor U4465 (N_4465,In_2094,In_1216);
xnor U4466 (N_4466,In_597,In_2182);
or U4467 (N_4467,In_927,In_2585);
xnor U4468 (N_4468,In_1735,In_1317);
and U4469 (N_4469,In_1501,In_2314);
and U4470 (N_4470,In_1117,In_1797);
nand U4471 (N_4471,In_1516,In_2691);
xor U4472 (N_4472,In_2116,In_988);
and U4473 (N_4473,In_638,In_229);
nand U4474 (N_4474,In_1219,In_2380);
and U4475 (N_4475,In_1811,In_1176);
nor U4476 (N_4476,In_2834,In_2415);
or U4477 (N_4477,In_2283,In_2744);
xor U4478 (N_4478,In_153,In_2112);
or U4479 (N_4479,In_1285,In_762);
nor U4480 (N_4480,In_460,In_968);
and U4481 (N_4481,In_193,In_775);
nand U4482 (N_4482,In_327,In_2206);
and U4483 (N_4483,In_573,In_772);
nor U4484 (N_4484,In_2752,In_1965);
xor U4485 (N_4485,In_1824,In_266);
nor U4486 (N_4486,In_816,In_747);
nand U4487 (N_4487,In_661,In_886);
and U4488 (N_4488,In_185,In_1207);
xnor U4489 (N_4489,In_2680,In_774);
or U4490 (N_4490,In_352,In_215);
xnor U4491 (N_4491,In_2645,In_2699);
and U4492 (N_4492,In_287,In_894);
nor U4493 (N_4493,In_1369,In_2949);
xnor U4494 (N_4494,In_1450,In_101);
nor U4495 (N_4495,In_2666,In_1657);
xor U4496 (N_4496,In_2428,In_2589);
xor U4497 (N_4497,In_2566,In_1804);
or U4498 (N_4498,In_2106,In_2950);
and U4499 (N_4499,In_1819,In_2623);
nor U4500 (N_4500,In_1947,In_1897);
and U4501 (N_4501,In_946,In_2250);
nor U4502 (N_4502,In_1158,In_802);
or U4503 (N_4503,In_2533,In_983);
nor U4504 (N_4504,In_2223,In_569);
or U4505 (N_4505,In_309,In_2262);
xnor U4506 (N_4506,In_2641,In_2575);
xor U4507 (N_4507,In_832,In_431);
and U4508 (N_4508,In_1923,In_448);
xnor U4509 (N_4509,In_1723,In_2626);
xnor U4510 (N_4510,In_2876,In_257);
nand U4511 (N_4511,In_784,In_177);
nand U4512 (N_4512,In_123,In_2395);
and U4513 (N_4513,In_1692,In_669);
and U4514 (N_4514,In_478,In_2272);
xnor U4515 (N_4515,In_2793,In_2404);
nor U4516 (N_4516,In_807,In_805);
and U4517 (N_4517,In_2213,In_2356);
xor U4518 (N_4518,In_496,In_1352);
or U4519 (N_4519,In_2381,In_1074);
and U4520 (N_4520,In_2184,In_762);
xnor U4521 (N_4521,In_1608,In_1969);
and U4522 (N_4522,In_1934,In_383);
nand U4523 (N_4523,In_2944,In_149);
nor U4524 (N_4524,In_705,In_2226);
and U4525 (N_4525,In_397,In_2712);
and U4526 (N_4526,In_624,In_242);
xnor U4527 (N_4527,In_1008,In_2438);
nor U4528 (N_4528,In_1564,In_2869);
xnor U4529 (N_4529,In_2470,In_861);
and U4530 (N_4530,In_1789,In_1897);
nand U4531 (N_4531,In_492,In_346);
nand U4532 (N_4532,In_2427,In_351);
or U4533 (N_4533,In_556,In_365);
or U4534 (N_4534,In_115,In_784);
nor U4535 (N_4535,In_2200,In_1277);
nor U4536 (N_4536,In_1490,In_2761);
xnor U4537 (N_4537,In_935,In_1663);
or U4538 (N_4538,In_1580,In_1784);
nand U4539 (N_4539,In_1458,In_828);
nor U4540 (N_4540,In_570,In_1938);
xnor U4541 (N_4541,In_1980,In_60);
nand U4542 (N_4542,In_1522,In_1091);
xnor U4543 (N_4543,In_2681,In_1419);
xnor U4544 (N_4544,In_2436,In_2855);
nor U4545 (N_4545,In_2414,In_1401);
and U4546 (N_4546,In_286,In_424);
and U4547 (N_4547,In_1205,In_1748);
and U4548 (N_4548,In_1643,In_1429);
nand U4549 (N_4549,In_1101,In_2159);
and U4550 (N_4550,In_2343,In_1224);
xnor U4551 (N_4551,In_2246,In_612);
and U4552 (N_4552,In_845,In_2593);
nor U4553 (N_4553,In_361,In_724);
or U4554 (N_4554,In_2686,In_1820);
xnor U4555 (N_4555,In_2008,In_2729);
nand U4556 (N_4556,In_2239,In_1579);
nand U4557 (N_4557,In_47,In_1202);
or U4558 (N_4558,In_2706,In_1691);
nor U4559 (N_4559,In_2369,In_1868);
and U4560 (N_4560,In_2901,In_2867);
and U4561 (N_4561,In_1695,In_434);
nor U4562 (N_4562,In_194,In_124);
nor U4563 (N_4563,In_1470,In_2371);
and U4564 (N_4564,In_2124,In_993);
xor U4565 (N_4565,In_452,In_1377);
xnor U4566 (N_4566,In_2302,In_2321);
or U4567 (N_4567,In_2049,In_2600);
nand U4568 (N_4568,In_2286,In_1380);
nand U4569 (N_4569,In_2243,In_1886);
nand U4570 (N_4570,In_2553,In_1321);
and U4571 (N_4571,In_402,In_583);
and U4572 (N_4572,In_489,In_25);
nand U4573 (N_4573,In_2356,In_1753);
or U4574 (N_4574,In_1397,In_2720);
or U4575 (N_4575,In_756,In_1806);
xor U4576 (N_4576,In_55,In_351);
or U4577 (N_4577,In_663,In_2993);
xor U4578 (N_4578,In_175,In_991);
or U4579 (N_4579,In_360,In_227);
and U4580 (N_4580,In_1060,In_2524);
nand U4581 (N_4581,In_1354,In_55);
xor U4582 (N_4582,In_197,In_936);
nand U4583 (N_4583,In_2859,In_637);
and U4584 (N_4584,In_1106,In_1085);
nor U4585 (N_4585,In_888,In_2304);
xor U4586 (N_4586,In_1705,In_243);
and U4587 (N_4587,In_1976,In_512);
and U4588 (N_4588,In_2504,In_2317);
nor U4589 (N_4589,In_744,In_477);
and U4590 (N_4590,In_2763,In_2483);
xnor U4591 (N_4591,In_1917,In_970);
xor U4592 (N_4592,In_1736,In_2509);
nor U4593 (N_4593,In_1728,In_2420);
and U4594 (N_4594,In_2248,In_1742);
and U4595 (N_4595,In_34,In_729);
or U4596 (N_4596,In_643,In_1449);
nor U4597 (N_4597,In_1275,In_2194);
and U4598 (N_4598,In_2314,In_2557);
and U4599 (N_4599,In_51,In_2755);
xor U4600 (N_4600,In_1013,In_1220);
xor U4601 (N_4601,In_360,In_1834);
xnor U4602 (N_4602,In_1092,In_1483);
and U4603 (N_4603,In_1690,In_1374);
xnor U4604 (N_4604,In_1841,In_2730);
or U4605 (N_4605,In_2691,In_2982);
xor U4606 (N_4606,In_1950,In_1158);
nand U4607 (N_4607,In_2487,In_888);
or U4608 (N_4608,In_1129,In_2122);
and U4609 (N_4609,In_2461,In_2780);
xnor U4610 (N_4610,In_619,In_1824);
or U4611 (N_4611,In_1581,In_1979);
or U4612 (N_4612,In_1415,In_752);
and U4613 (N_4613,In_1075,In_953);
nand U4614 (N_4614,In_2634,In_2789);
or U4615 (N_4615,In_331,In_2500);
nor U4616 (N_4616,In_815,In_975);
and U4617 (N_4617,In_2833,In_2495);
nand U4618 (N_4618,In_1235,In_678);
or U4619 (N_4619,In_567,In_2239);
and U4620 (N_4620,In_2472,In_640);
or U4621 (N_4621,In_557,In_2744);
nor U4622 (N_4622,In_2400,In_339);
nor U4623 (N_4623,In_2443,In_544);
xnor U4624 (N_4624,In_837,In_2146);
nand U4625 (N_4625,In_1557,In_2379);
and U4626 (N_4626,In_2152,In_89);
xnor U4627 (N_4627,In_2384,In_90);
nand U4628 (N_4628,In_625,In_2498);
and U4629 (N_4629,In_982,In_153);
and U4630 (N_4630,In_618,In_2277);
nand U4631 (N_4631,In_704,In_646);
nand U4632 (N_4632,In_953,In_2584);
xnor U4633 (N_4633,In_945,In_251);
nand U4634 (N_4634,In_1402,In_1717);
nand U4635 (N_4635,In_2111,In_1333);
nor U4636 (N_4636,In_914,In_2484);
nor U4637 (N_4637,In_1115,In_937);
or U4638 (N_4638,In_2946,In_1789);
nor U4639 (N_4639,In_794,In_2294);
or U4640 (N_4640,In_1806,In_2166);
or U4641 (N_4641,In_92,In_1125);
xor U4642 (N_4642,In_329,In_405);
xor U4643 (N_4643,In_255,In_2285);
nor U4644 (N_4644,In_1411,In_2355);
and U4645 (N_4645,In_2348,In_344);
nand U4646 (N_4646,In_1749,In_144);
nor U4647 (N_4647,In_2064,In_220);
nand U4648 (N_4648,In_1146,In_2621);
and U4649 (N_4649,In_1457,In_1562);
nor U4650 (N_4650,In_29,In_1300);
and U4651 (N_4651,In_1707,In_2438);
or U4652 (N_4652,In_20,In_1075);
nand U4653 (N_4653,In_992,In_2813);
or U4654 (N_4654,In_294,In_2832);
nor U4655 (N_4655,In_2671,In_1631);
and U4656 (N_4656,In_1538,In_1702);
nand U4657 (N_4657,In_502,In_314);
or U4658 (N_4658,In_308,In_1219);
nand U4659 (N_4659,In_642,In_1156);
and U4660 (N_4660,In_994,In_1211);
or U4661 (N_4661,In_1741,In_153);
nand U4662 (N_4662,In_2824,In_718);
nand U4663 (N_4663,In_2801,In_461);
nand U4664 (N_4664,In_1824,In_2541);
or U4665 (N_4665,In_571,In_2222);
nand U4666 (N_4666,In_1999,In_992);
nor U4667 (N_4667,In_1782,In_2240);
nor U4668 (N_4668,In_1247,In_1847);
nor U4669 (N_4669,In_2205,In_1522);
nor U4670 (N_4670,In_2183,In_2786);
or U4671 (N_4671,In_1341,In_2378);
or U4672 (N_4672,In_773,In_1408);
and U4673 (N_4673,In_2938,In_1860);
or U4674 (N_4674,In_494,In_1256);
nor U4675 (N_4675,In_890,In_2335);
xor U4676 (N_4676,In_1032,In_439);
nand U4677 (N_4677,In_503,In_2400);
nand U4678 (N_4678,In_2053,In_1951);
xor U4679 (N_4679,In_306,In_2407);
nand U4680 (N_4680,In_576,In_738);
xor U4681 (N_4681,In_331,In_2426);
or U4682 (N_4682,In_1639,In_652);
xnor U4683 (N_4683,In_2755,In_210);
and U4684 (N_4684,In_1293,In_317);
nand U4685 (N_4685,In_1702,In_1835);
or U4686 (N_4686,In_1781,In_2539);
nor U4687 (N_4687,In_1347,In_2677);
nand U4688 (N_4688,In_193,In_2244);
and U4689 (N_4689,In_1748,In_1244);
xor U4690 (N_4690,In_1711,In_2122);
xnor U4691 (N_4691,In_174,In_1525);
nor U4692 (N_4692,In_190,In_401);
xor U4693 (N_4693,In_2235,In_2930);
nor U4694 (N_4694,In_2692,In_840);
nor U4695 (N_4695,In_1143,In_2304);
nor U4696 (N_4696,In_152,In_6);
xnor U4697 (N_4697,In_2079,In_1183);
or U4698 (N_4698,In_2928,In_2892);
and U4699 (N_4699,In_1130,In_1394);
and U4700 (N_4700,In_573,In_2382);
or U4701 (N_4701,In_1953,In_1805);
xnor U4702 (N_4702,In_2289,In_1230);
nand U4703 (N_4703,In_2852,In_902);
or U4704 (N_4704,In_1966,In_1244);
or U4705 (N_4705,In_2890,In_2052);
nor U4706 (N_4706,In_534,In_701);
nor U4707 (N_4707,In_1653,In_2257);
nand U4708 (N_4708,In_1791,In_3);
and U4709 (N_4709,In_649,In_587);
nor U4710 (N_4710,In_1476,In_110);
xor U4711 (N_4711,In_1284,In_542);
xor U4712 (N_4712,In_384,In_556);
xor U4713 (N_4713,In_549,In_553);
nand U4714 (N_4714,In_519,In_2390);
or U4715 (N_4715,In_1568,In_1065);
and U4716 (N_4716,In_154,In_139);
and U4717 (N_4717,In_2141,In_196);
nand U4718 (N_4718,In_2223,In_1354);
xor U4719 (N_4719,In_2637,In_2028);
xor U4720 (N_4720,In_68,In_1970);
nand U4721 (N_4721,In_2767,In_270);
nor U4722 (N_4722,In_136,In_2297);
or U4723 (N_4723,In_1245,In_570);
nand U4724 (N_4724,In_1193,In_738);
nand U4725 (N_4725,In_2395,In_1631);
xnor U4726 (N_4726,In_1834,In_23);
xor U4727 (N_4727,In_2930,In_691);
or U4728 (N_4728,In_148,In_436);
and U4729 (N_4729,In_1102,In_2066);
xnor U4730 (N_4730,In_1777,In_2665);
xor U4731 (N_4731,In_2215,In_375);
xnor U4732 (N_4732,In_2838,In_429);
and U4733 (N_4733,In_2261,In_2471);
nand U4734 (N_4734,In_2286,In_98);
nand U4735 (N_4735,In_2114,In_1297);
nand U4736 (N_4736,In_39,In_1608);
nor U4737 (N_4737,In_1303,In_1013);
nand U4738 (N_4738,In_2742,In_550);
xnor U4739 (N_4739,In_1737,In_1612);
and U4740 (N_4740,In_1650,In_1837);
nor U4741 (N_4741,In_821,In_814);
xnor U4742 (N_4742,In_1478,In_1449);
xor U4743 (N_4743,In_1469,In_2828);
nor U4744 (N_4744,In_2389,In_2819);
and U4745 (N_4745,In_2432,In_501);
and U4746 (N_4746,In_2452,In_773);
xor U4747 (N_4747,In_1162,In_9);
nand U4748 (N_4748,In_1734,In_2447);
nor U4749 (N_4749,In_2108,In_420);
xnor U4750 (N_4750,In_528,In_224);
nor U4751 (N_4751,In_672,In_245);
nor U4752 (N_4752,In_2456,In_2668);
and U4753 (N_4753,In_1375,In_1282);
and U4754 (N_4754,In_82,In_2317);
and U4755 (N_4755,In_2844,In_244);
nor U4756 (N_4756,In_2246,In_1651);
or U4757 (N_4757,In_85,In_1883);
nand U4758 (N_4758,In_629,In_2090);
nand U4759 (N_4759,In_2180,In_2051);
and U4760 (N_4760,In_137,In_2106);
nand U4761 (N_4761,In_1547,In_951);
nand U4762 (N_4762,In_2132,In_307);
or U4763 (N_4763,In_1473,In_2102);
and U4764 (N_4764,In_125,In_2636);
or U4765 (N_4765,In_207,In_1716);
or U4766 (N_4766,In_1704,In_521);
xor U4767 (N_4767,In_2173,In_1226);
xnor U4768 (N_4768,In_2042,In_368);
nor U4769 (N_4769,In_2703,In_2567);
or U4770 (N_4770,In_1615,In_1609);
nand U4771 (N_4771,In_833,In_1283);
or U4772 (N_4772,In_2484,In_2791);
nor U4773 (N_4773,In_1116,In_1050);
or U4774 (N_4774,In_1755,In_1097);
xor U4775 (N_4775,In_2322,In_584);
or U4776 (N_4776,In_2189,In_332);
or U4777 (N_4777,In_512,In_911);
nor U4778 (N_4778,In_759,In_1990);
or U4779 (N_4779,In_879,In_1181);
xnor U4780 (N_4780,In_2131,In_900);
nor U4781 (N_4781,In_2393,In_620);
nor U4782 (N_4782,In_741,In_1915);
nand U4783 (N_4783,In_905,In_1367);
or U4784 (N_4784,In_386,In_2568);
nor U4785 (N_4785,In_2671,In_1449);
nand U4786 (N_4786,In_2887,In_282);
nor U4787 (N_4787,In_2410,In_1307);
nor U4788 (N_4788,In_2201,In_580);
xnor U4789 (N_4789,In_2293,In_330);
nand U4790 (N_4790,In_27,In_973);
xnor U4791 (N_4791,In_976,In_1352);
nor U4792 (N_4792,In_87,In_1357);
or U4793 (N_4793,In_1160,In_1517);
nor U4794 (N_4794,In_2183,In_1662);
nor U4795 (N_4795,In_391,In_590);
nor U4796 (N_4796,In_2024,In_970);
nor U4797 (N_4797,In_2226,In_2392);
and U4798 (N_4798,In_1722,In_1856);
or U4799 (N_4799,In_2387,In_764);
or U4800 (N_4800,In_1704,In_1306);
nor U4801 (N_4801,In_1557,In_1628);
nand U4802 (N_4802,In_262,In_331);
xor U4803 (N_4803,In_2566,In_1447);
or U4804 (N_4804,In_641,In_2919);
nand U4805 (N_4805,In_2591,In_354);
nand U4806 (N_4806,In_1361,In_1142);
or U4807 (N_4807,In_477,In_1037);
and U4808 (N_4808,In_2436,In_1703);
nor U4809 (N_4809,In_2168,In_1659);
nor U4810 (N_4810,In_801,In_605);
and U4811 (N_4811,In_29,In_2479);
and U4812 (N_4812,In_363,In_1146);
xor U4813 (N_4813,In_828,In_673);
or U4814 (N_4814,In_1488,In_2792);
or U4815 (N_4815,In_1234,In_2508);
nand U4816 (N_4816,In_549,In_512);
nand U4817 (N_4817,In_693,In_469);
nand U4818 (N_4818,In_2172,In_474);
and U4819 (N_4819,In_2369,In_256);
or U4820 (N_4820,In_1348,In_1073);
nor U4821 (N_4821,In_2719,In_1322);
nand U4822 (N_4822,In_1625,In_2195);
or U4823 (N_4823,In_1343,In_2354);
nor U4824 (N_4824,In_1999,In_346);
and U4825 (N_4825,In_1723,In_1797);
and U4826 (N_4826,In_640,In_2623);
and U4827 (N_4827,In_611,In_1613);
nor U4828 (N_4828,In_556,In_2173);
nand U4829 (N_4829,In_2460,In_561);
or U4830 (N_4830,In_1772,In_1044);
nand U4831 (N_4831,In_183,In_11);
xor U4832 (N_4832,In_330,In_1631);
nor U4833 (N_4833,In_5,In_2787);
xnor U4834 (N_4834,In_2018,In_2036);
xnor U4835 (N_4835,In_1609,In_2667);
and U4836 (N_4836,In_2538,In_2558);
nand U4837 (N_4837,In_1231,In_23);
xor U4838 (N_4838,In_675,In_1518);
nor U4839 (N_4839,In_713,In_2692);
and U4840 (N_4840,In_840,In_160);
nor U4841 (N_4841,In_542,In_128);
and U4842 (N_4842,In_1685,In_1589);
nand U4843 (N_4843,In_1946,In_1839);
nand U4844 (N_4844,In_1533,In_2784);
nand U4845 (N_4845,In_2095,In_848);
and U4846 (N_4846,In_1647,In_2790);
nand U4847 (N_4847,In_804,In_1405);
nor U4848 (N_4848,In_1547,In_636);
and U4849 (N_4849,In_584,In_1900);
or U4850 (N_4850,In_1497,In_2457);
nand U4851 (N_4851,In_1985,In_329);
nor U4852 (N_4852,In_1617,In_2108);
and U4853 (N_4853,In_1861,In_2338);
or U4854 (N_4854,In_1691,In_2530);
and U4855 (N_4855,In_1466,In_577);
nor U4856 (N_4856,In_994,In_2018);
and U4857 (N_4857,In_957,In_2605);
nand U4858 (N_4858,In_1432,In_1986);
xor U4859 (N_4859,In_1267,In_2010);
and U4860 (N_4860,In_2003,In_1053);
and U4861 (N_4861,In_817,In_2344);
nand U4862 (N_4862,In_1178,In_1456);
and U4863 (N_4863,In_1859,In_1031);
or U4864 (N_4864,In_410,In_453);
and U4865 (N_4865,In_1345,In_844);
xor U4866 (N_4866,In_996,In_255);
or U4867 (N_4867,In_857,In_770);
xnor U4868 (N_4868,In_400,In_2521);
and U4869 (N_4869,In_1818,In_2699);
nor U4870 (N_4870,In_2493,In_1925);
or U4871 (N_4871,In_2672,In_491);
xnor U4872 (N_4872,In_1408,In_1061);
and U4873 (N_4873,In_154,In_76);
nand U4874 (N_4874,In_1242,In_1477);
xnor U4875 (N_4875,In_2628,In_2294);
nand U4876 (N_4876,In_918,In_1859);
nor U4877 (N_4877,In_543,In_1045);
and U4878 (N_4878,In_366,In_1350);
or U4879 (N_4879,In_2497,In_86);
nor U4880 (N_4880,In_1033,In_2976);
or U4881 (N_4881,In_2029,In_934);
or U4882 (N_4882,In_1959,In_2800);
xor U4883 (N_4883,In_1844,In_2290);
or U4884 (N_4884,In_44,In_2970);
xor U4885 (N_4885,In_722,In_2630);
or U4886 (N_4886,In_582,In_1367);
or U4887 (N_4887,In_1955,In_1382);
and U4888 (N_4888,In_584,In_58);
xor U4889 (N_4889,In_24,In_2933);
or U4890 (N_4890,In_2398,In_948);
nor U4891 (N_4891,In_2797,In_795);
xnor U4892 (N_4892,In_1306,In_2759);
nor U4893 (N_4893,In_452,In_327);
or U4894 (N_4894,In_108,In_971);
and U4895 (N_4895,In_1859,In_2126);
and U4896 (N_4896,In_2950,In_570);
nand U4897 (N_4897,In_2556,In_568);
nor U4898 (N_4898,In_2007,In_1937);
or U4899 (N_4899,In_2480,In_2801);
nand U4900 (N_4900,In_2145,In_1564);
nor U4901 (N_4901,In_1258,In_2904);
nor U4902 (N_4902,In_2875,In_934);
and U4903 (N_4903,In_842,In_768);
xnor U4904 (N_4904,In_1813,In_364);
or U4905 (N_4905,In_1503,In_1129);
or U4906 (N_4906,In_1179,In_1895);
or U4907 (N_4907,In_1994,In_1211);
nand U4908 (N_4908,In_606,In_2850);
nand U4909 (N_4909,In_2744,In_1539);
nand U4910 (N_4910,In_140,In_2042);
nand U4911 (N_4911,In_375,In_971);
and U4912 (N_4912,In_1671,In_2833);
and U4913 (N_4913,In_40,In_897);
and U4914 (N_4914,In_934,In_190);
xnor U4915 (N_4915,In_546,In_1378);
nor U4916 (N_4916,In_2192,In_2218);
xnor U4917 (N_4917,In_814,In_1556);
xor U4918 (N_4918,In_43,In_2268);
and U4919 (N_4919,In_2476,In_1507);
or U4920 (N_4920,In_50,In_1538);
xor U4921 (N_4921,In_2317,In_537);
and U4922 (N_4922,In_636,In_1749);
or U4923 (N_4923,In_1776,In_518);
nor U4924 (N_4924,In_1043,In_2130);
and U4925 (N_4925,In_1904,In_349);
or U4926 (N_4926,In_2587,In_1157);
nor U4927 (N_4927,In_2077,In_1522);
nor U4928 (N_4928,In_401,In_1143);
or U4929 (N_4929,In_1524,In_1149);
nor U4930 (N_4930,In_1959,In_2628);
nor U4931 (N_4931,In_1484,In_1700);
nand U4932 (N_4932,In_1465,In_294);
nand U4933 (N_4933,In_198,In_1748);
and U4934 (N_4934,In_2232,In_1762);
nand U4935 (N_4935,In_662,In_1659);
nor U4936 (N_4936,In_2017,In_2468);
nor U4937 (N_4937,In_1383,In_637);
nor U4938 (N_4938,In_2512,In_1793);
and U4939 (N_4939,In_639,In_1862);
and U4940 (N_4940,In_1029,In_2893);
and U4941 (N_4941,In_2118,In_2934);
xor U4942 (N_4942,In_2131,In_2818);
or U4943 (N_4943,In_2239,In_1641);
and U4944 (N_4944,In_2859,In_292);
nand U4945 (N_4945,In_440,In_2900);
and U4946 (N_4946,In_2230,In_2099);
nand U4947 (N_4947,In_392,In_2189);
nor U4948 (N_4948,In_1788,In_2373);
and U4949 (N_4949,In_2760,In_1411);
and U4950 (N_4950,In_2887,In_2534);
and U4951 (N_4951,In_2233,In_980);
nand U4952 (N_4952,In_1226,In_959);
or U4953 (N_4953,In_2191,In_2119);
or U4954 (N_4954,In_2232,In_930);
and U4955 (N_4955,In_1094,In_2402);
xnor U4956 (N_4956,In_1028,In_1060);
xor U4957 (N_4957,In_2816,In_189);
or U4958 (N_4958,In_2989,In_1384);
and U4959 (N_4959,In_2425,In_2036);
and U4960 (N_4960,In_2838,In_30);
and U4961 (N_4961,In_1727,In_748);
or U4962 (N_4962,In_1853,In_1481);
and U4963 (N_4963,In_1663,In_1914);
nor U4964 (N_4964,In_1433,In_1476);
or U4965 (N_4965,In_2187,In_1361);
nand U4966 (N_4966,In_1083,In_2628);
xnor U4967 (N_4967,In_1871,In_190);
nor U4968 (N_4968,In_1304,In_1433);
nand U4969 (N_4969,In_790,In_353);
or U4970 (N_4970,In_2408,In_2930);
nor U4971 (N_4971,In_387,In_692);
or U4972 (N_4972,In_1081,In_796);
and U4973 (N_4973,In_2016,In_2962);
and U4974 (N_4974,In_1001,In_751);
xor U4975 (N_4975,In_1530,In_1332);
xor U4976 (N_4976,In_1727,In_2845);
xnor U4977 (N_4977,In_612,In_2969);
or U4978 (N_4978,In_640,In_285);
or U4979 (N_4979,In_2600,In_571);
nand U4980 (N_4980,In_1997,In_2684);
xnor U4981 (N_4981,In_469,In_893);
or U4982 (N_4982,In_1304,In_662);
or U4983 (N_4983,In_847,In_621);
nor U4984 (N_4984,In_97,In_1692);
nor U4985 (N_4985,In_1265,In_911);
xnor U4986 (N_4986,In_445,In_806);
nor U4987 (N_4987,In_80,In_1102);
nor U4988 (N_4988,In_1600,In_655);
nand U4989 (N_4989,In_2502,In_2305);
or U4990 (N_4990,In_1157,In_2510);
nand U4991 (N_4991,In_2593,In_814);
nand U4992 (N_4992,In_1243,In_1437);
and U4993 (N_4993,In_379,In_866);
and U4994 (N_4994,In_3,In_2228);
and U4995 (N_4995,In_1641,In_781);
or U4996 (N_4996,In_599,In_909);
and U4997 (N_4997,In_2311,In_668);
xnor U4998 (N_4998,In_1334,In_1760);
or U4999 (N_4999,In_942,In_300);
nand U5000 (N_5000,N_583,N_812);
and U5001 (N_5001,N_3824,N_4764);
nor U5002 (N_5002,N_908,N_2859);
or U5003 (N_5003,N_1649,N_3188);
or U5004 (N_5004,N_471,N_4649);
or U5005 (N_5005,N_342,N_3379);
and U5006 (N_5006,N_4920,N_599);
xnor U5007 (N_5007,N_1576,N_2854);
nor U5008 (N_5008,N_4289,N_232);
nand U5009 (N_5009,N_434,N_1998);
and U5010 (N_5010,N_3167,N_754);
nor U5011 (N_5011,N_4219,N_3994);
nor U5012 (N_5012,N_4724,N_1197);
or U5013 (N_5013,N_3268,N_3323);
nor U5014 (N_5014,N_3898,N_4576);
xor U5015 (N_5015,N_2210,N_3484);
nor U5016 (N_5016,N_94,N_2561);
nor U5017 (N_5017,N_4389,N_4507);
nand U5018 (N_5018,N_1131,N_3461);
or U5019 (N_5019,N_4470,N_4010);
or U5020 (N_5020,N_2282,N_4012);
xor U5021 (N_5021,N_1714,N_2898);
nand U5022 (N_5022,N_3077,N_1697);
or U5023 (N_5023,N_938,N_2646);
xor U5024 (N_5024,N_1170,N_40);
or U5025 (N_5025,N_2619,N_4222);
nand U5026 (N_5026,N_454,N_4917);
nand U5027 (N_5027,N_3131,N_1051);
xor U5028 (N_5028,N_4819,N_2693);
or U5029 (N_5029,N_3711,N_1348);
and U5030 (N_5030,N_2221,N_1160);
or U5031 (N_5031,N_1600,N_4338);
xor U5032 (N_5032,N_3515,N_4652);
xnor U5033 (N_5033,N_2392,N_2625);
or U5034 (N_5034,N_3799,N_2275);
and U5035 (N_5035,N_4272,N_4947);
nand U5036 (N_5036,N_621,N_2658);
and U5037 (N_5037,N_2986,N_1428);
xor U5038 (N_5038,N_3511,N_2167);
or U5039 (N_5039,N_3840,N_3398);
xnor U5040 (N_5040,N_1320,N_4036);
and U5041 (N_5041,N_3069,N_3298);
and U5042 (N_5042,N_2756,N_1311);
or U5043 (N_5043,N_4069,N_969);
nand U5044 (N_5044,N_1662,N_474);
or U5045 (N_5045,N_4665,N_3970);
or U5046 (N_5046,N_245,N_2074);
nor U5047 (N_5047,N_1945,N_2034);
nor U5048 (N_5048,N_395,N_2029);
nor U5049 (N_5049,N_1145,N_2610);
nand U5050 (N_5050,N_4377,N_1106);
nor U5051 (N_5051,N_4633,N_93);
nand U5052 (N_5052,N_3943,N_2445);
and U5053 (N_5053,N_674,N_4335);
nand U5054 (N_5054,N_1818,N_48);
nor U5055 (N_5055,N_1217,N_548);
nand U5056 (N_5056,N_1684,N_1836);
nand U5057 (N_5057,N_296,N_64);
and U5058 (N_5058,N_3396,N_1720);
and U5059 (N_5059,N_1400,N_1349);
and U5060 (N_5060,N_4963,N_2021);
xnor U5061 (N_5061,N_1833,N_1553);
nand U5062 (N_5062,N_3636,N_473);
nand U5063 (N_5063,N_121,N_1515);
or U5064 (N_5064,N_4136,N_2052);
or U5065 (N_5065,N_4570,N_1177);
nor U5066 (N_5066,N_3063,N_2801);
nand U5067 (N_5067,N_4580,N_1538);
nand U5068 (N_5068,N_2541,N_1977);
xnor U5069 (N_5069,N_2968,N_1883);
nor U5070 (N_5070,N_338,N_785);
nand U5071 (N_5071,N_402,N_1816);
xor U5072 (N_5072,N_1847,N_562);
and U5073 (N_5073,N_3614,N_3562);
nand U5074 (N_5074,N_3776,N_4726);
xnor U5075 (N_5075,N_3561,N_2039);
and U5076 (N_5076,N_2344,N_2516);
nor U5077 (N_5077,N_4096,N_704);
nor U5078 (N_5078,N_4479,N_3748);
nor U5079 (N_5079,N_2082,N_2791);
nor U5080 (N_5080,N_1689,N_3767);
xnor U5081 (N_5081,N_1931,N_1245);
nor U5082 (N_5082,N_2355,N_4591);
and U5083 (N_5083,N_227,N_192);
or U5084 (N_5084,N_1295,N_2284);
nand U5085 (N_5085,N_1050,N_4748);
or U5086 (N_5086,N_1656,N_580);
or U5087 (N_5087,N_2691,N_375);
xnor U5088 (N_5088,N_687,N_3201);
nand U5089 (N_5089,N_2790,N_2844);
xnor U5090 (N_5090,N_696,N_4380);
xor U5091 (N_5091,N_4695,N_551);
xnor U5092 (N_5092,N_3107,N_1301);
and U5093 (N_5093,N_2003,N_4303);
xnor U5094 (N_5094,N_3883,N_4004);
or U5095 (N_5095,N_3966,N_3411);
nor U5096 (N_5096,N_675,N_3982);
xnor U5097 (N_5097,N_4405,N_107);
and U5098 (N_5098,N_3645,N_2218);
xnor U5099 (N_5099,N_678,N_377);
nand U5100 (N_5100,N_881,N_462);
nand U5101 (N_5101,N_55,N_1156);
nand U5102 (N_5102,N_1746,N_1770);
nor U5103 (N_5103,N_4935,N_4539);
or U5104 (N_5104,N_3090,N_3231);
and U5105 (N_5105,N_4631,N_4880);
nor U5106 (N_5106,N_4934,N_1469);
and U5107 (N_5107,N_1278,N_1627);
nand U5108 (N_5108,N_733,N_482);
and U5109 (N_5109,N_4108,N_4533);
and U5110 (N_5110,N_447,N_2489);
nor U5111 (N_5111,N_1372,N_4195);
nor U5112 (N_5112,N_824,N_2199);
nor U5113 (N_5113,N_2297,N_1316);
and U5114 (N_5114,N_3370,N_1915);
nand U5115 (N_5115,N_2931,N_470);
nor U5116 (N_5116,N_265,N_3859);
xor U5117 (N_5117,N_1364,N_398);
and U5118 (N_5118,N_3083,N_489);
or U5119 (N_5119,N_2660,N_2747);
nand U5120 (N_5120,N_1060,N_1448);
nand U5121 (N_5121,N_651,N_1205);
nor U5122 (N_5122,N_4171,N_2925);
or U5123 (N_5123,N_3429,N_4813);
xnor U5124 (N_5124,N_953,N_3691);
nand U5125 (N_5125,N_4116,N_4605);
nor U5126 (N_5126,N_1404,N_579);
nand U5127 (N_5127,N_4566,N_3774);
nor U5128 (N_5128,N_1834,N_3794);
nand U5129 (N_5129,N_4721,N_4937);
nor U5130 (N_5130,N_1323,N_1298);
nor U5131 (N_5131,N_4121,N_3642);
xor U5132 (N_5132,N_4766,N_176);
nand U5133 (N_5133,N_1195,N_4913);
or U5134 (N_5134,N_1228,N_1490);
and U5135 (N_5135,N_4824,N_1992);
nor U5136 (N_5136,N_1505,N_1957);
nand U5137 (N_5137,N_3375,N_2554);
or U5138 (N_5138,N_3655,N_4158);
or U5139 (N_5139,N_4231,N_4246);
or U5140 (N_5140,N_3708,N_3560);
nor U5141 (N_5141,N_1378,N_2110);
xnor U5142 (N_5142,N_4024,N_528);
nor U5143 (N_5143,N_1613,N_4878);
or U5144 (N_5144,N_4543,N_541);
and U5145 (N_5145,N_1263,N_4157);
nor U5146 (N_5146,N_3670,N_2696);
nand U5147 (N_5147,N_2111,N_4581);
or U5148 (N_5148,N_381,N_2534);
or U5149 (N_5149,N_3781,N_1483);
nor U5150 (N_5150,N_1109,N_2500);
nor U5151 (N_5151,N_3504,N_119);
and U5152 (N_5152,N_3246,N_122);
or U5153 (N_5153,N_4446,N_2088);
nor U5154 (N_5154,N_3110,N_1086);
xor U5155 (N_5155,N_2817,N_2623);
and U5156 (N_5156,N_2170,N_2136);
xnor U5157 (N_5157,N_2182,N_3101);
nor U5158 (N_5158,N_3959,N_83);
or U5159 (N_5159,N_1875,N_131);
xnor U5160 (N_5160,N_775,N_4471);
or U5161 (N_5161,N_4911,N_4867);
or U5162 (N_5162,N_2771,N_2874);
or U5163 (N_5163,N_3972,N_3444);
or U5164 (N_5164,N_3307,N_1650);
xnor U5165 (N_5165,N_2853,N_1068);
and U5166 (N_5166,N_2682,N_3261);
nand U5167 (N_5167,N_3588,N_2954);
xor U5168 (N_5168,N_1517,N_335);
and U5169 (N_5169,N_1528,N_1560);
nor U5170 (N_5170,N_4902,N_2031);
nor U5171 (N_5171,N_4129,N_568);
nor U5172 (N_5172,N_590,N_2257);
and U5173 (N_5173,N_3577,N_2592);
xnor U5174 (N_5174,N_2286,N_1657);
nor U5175 (N_5175,N_4145,N_2905);
or U5176 (N_5176,N_2922,N_1822);
xnor U5177 (N_5177,N_4894,N_201);
or U5178 (N_5178,N_166,N_1933);
or U5179 (N_5179,N_1531,N_2155);
xnor U5180 (N_5180,N_2796,N_393);
or U5181 (N_5181,N_4704,N_3873);
nor U5182 (N_5182,N_4297,N_2615);
or U5183 (N_5183,N_4249,N_4943);
xor U5184 (N_5184,N_1212,N_2292);
xor U5185 (N_5185,N_1007,N_1853);
xnor U5186 (N_5186,N_3028,N_3076);
and U5187 (N_5187,N_1595,N_2187);
nor U5188 (N_5188,N_3773,N_4350);
nor U5189 (N_5189,N_526,N_382);
or U5190 (N_5190,N_1111,N_1837);
or U5191 (N_5191,N_4213,N_2066);
or U5192 (N_5192,N_206,N_3423);
and U5193 (N_5193,N_4737,N_445);
and U5194 (N_5194,N_1722,N_4861);
xnor U5195 (N_5195,N_936,N_2409);
xnor U5196 (N_5196,N_628,N_1710);
nand U5197 (N_5197,N_4945,N_118);
or U5198 (N_5198,N_3027,N_4968);
and U5199 (N_5199,N_3317,N_70);
nor U5200 (N_5200,N_2628,N_1139);
and U5201 (N_5201,N_2985,N_1831);
and U5202 (N_5202,N_3432,N_1824);
or U5203 (N_5203,N_4628,N_67);
nand U5204 (N_5204,N_4032,N_3762);
nand U5205 (N_5205,N_2429,N_2805);
nand U5206 (N_5206,N_198,N_1715);
nor U5207 (N_5207,N_4607,N_1376);
xnor U5208 (N_5208,N_3803,N_1488);
xnor U5209 (N_5209,N_1030,N_4042);
nor U5210 (N_5210,N_2010,N_175);
and U5211 (N_5211,N_3908,N_495);
and U5212 (N_5212,N_2733,N_1984);
nand U5213 (N_5213,N_1209,N_808);
nand U5214 (N_5214,N_1427,N_700);
and U5215 (N_5215,N_1440,N_1046);
nand U5216 (N_5216,N_3666,N_2472);
nor U5217 (N_5217,N_468,N_417);
nand U5218 (N_5218,N_2982,N_184);
nand U5219 (N_5219,N_1288,N_1201);
nor U5220 (N_5220,N_4199,N_2131);
and U5221 (N_5221,N_2401,N_3372);
or U5222 (N_5222,N_337,N_1609);
and U5223 (N_5223,N_4435,N_2171);
xor U5224 (N_5224,N_1959,N_3173);
nand U5225 (N_5225,N_3732,N_5);
nor U5226 (N_5226,N_303,N_2462);
and U5227 (N_5227,N_3291,N_4731);
xnor U5228 (N_5228,N_738,N_1669);
nand U5229 (N_5229,N_848,N_2381);
nand U5230 (N_5230,N_2024,N_889);
or U5231 (N_5231,N_2928,N_346);
xnor U5232 (N_5232,N_2942,N_4821);
and U5233 (N_5233,N_4608,N_4065);
xor U5234 (N_5234,N_1247,N_3009);
nor U5235 (N_5235,N_174,N_2588);
xnor U5236 (N_5236,N_1069,N_3166);
xnor U5237 (N_5237,N_777,N_2871);
nand U5238 (N_5238,N_4260,N_3595);
xnor U5239 (N_5239,N_2018,N_319);
nand U5240 (N_5240,N_62,N_4982);
nor U5241 (N_5241,N_3255,N_2882);
and U5242 (N_5242,N_1183,N_3071);
nor U5243 (N_5243,N_4162,N_2914);
nand U5244 (N_5244,N_1099,N_2255);
nor U5245 (N_5245,N_2271,N_4210);
or U5246 (N_5246,N_69,N_3106);
and U5247 (N_5247,N_4225,N_1127);
nor U5248 (N_5248,N_1732,N_4701);
and U5249 (N_5249,N_3386,N_2644);
nor U5250 (N_5250,N_1660,N_2886);
nand U5251 (N_5251,N_3153,N_2522);
or U5252 (N_5252,N_1329,N_4871);
nand U5253 (N_5253,N_1277,N_1485);
or U5254 (N_5254,N_4044,N_1681);
nor U5255 (N_5255,N_3041,N_3234);
nor U5256 (N_5256,N_1200,N_3336);
xor U5257 (N_5257,N_2224,N_301);
nand U5258 (N_5258,N_2328,N_4481);
nor U5259 (N_5259,N_1762,N_3467);
nor U5260 (N_5260,N_3015,N_2845);
and U5261 (N_5261,N_2061,N_3311);
xnor U5262 (N_5262,N_4038,N_2603);
or U5263 (N_5263,N_525,N_1466);
nand U5264 (N_5264,N_1224,N_4929);
nor U5265 (N_5265,N_4385,N_2840);
or U5266 (N_5266,N_3968,N_584);
nor U5267 (N_5267,N_750,N_2832);
nand U5268 (N_5268,N_469,N_4252);
nor U5269 (N_5269,N_299,N_3945);
or U5270 (N_5270,N_4176,N_3431);
nand U5271 (N_5271,N_1182,N_3122);
xnor U5272 (N_5272,N_1664,N_2059);
or U5273 (N_5273,N_1572,N_4251);
or U5274 (N_5274,N_4769,N_4430);
nand U5275 (N_5275,N_2080,N_4735);
or U5276 (N_5276,N_4002,N_4400);
nand U5277 (N_5277,N_2725,N_2988);
and U5278 (N_5278,N_1078,N_4835);
xnor U5279 (N_5279,N_1464,N_2737);
and U5280 (N_5280,N_1545,N_2647);
or U5281 (N_5281,N_3568,N_2249);
or U5282 (N_5282,N_310,N_1908);
nor U5283 (N_5283,N_4463,N_3425);
nand U5284 (N_5284,N_4349,N_878);
and U5285 (N_5285,N_2192,N_698);
nand U5286 (N_5286,N_266,N_4428);
nor U5287 (N_5287,N_3213,N_744);
xor U5288 (N_5288,N_2334,N_4742);
nor U5289 (N_5289,N_3659,N_2524);
xor U5290 (N_5290,N_4080,N_1645);
xnor U5291 (N_5291,N_1902,N_3332);
or U5292 (N_5292,N_3436,N_2939);
xnor U5293 (N_5293,N_2242,N_4897);
nand U5294 (N_5294,N_664,N_3486);
xor U5295 (N_5295,N_3316,N_1344);
or U5296 (N_5296,N_4041,N_8);
or U5297 (N_5297,N_1402,N_2890);
nand U5298 (N_5298,N_4087,N_2398);
nor U5299 (N_5299,N_3092,N_3476);
and U5300 (N_5300,N_3983,N_986);
or U5301 (N_5301,N_1641,N_4977);
or U5302 (N_5302,N_42,N_2700);
or U5303 (N_5303,N_2951,N_4351);
xor U5304 (N_5304,N_247,N_979);
xor U5305 (N_5305,N_2729,N_2576);
nand U5306 (N_5306,N_3768,N_2528);
nand U5307 (N_5307,N_748,N_1918);
and U5308 (N_5308,N_4402,N_2385);
and U5309 (N_5309,N_4314,N_3334);
xor U5310 (N_5310,N_4027,N_1423);
xor U5311 (N_5311,N_3879,N_4258);
and U5312 (N_5312,N_1486,N_1130);
nand U5313 (N_5313,N_2288,N_909);
or U5314 (N_5314,N_4173,N_927);
nand U5315 (N_5315,N_3144,N_4243);
or U5316 (N_5316,N_2690,N_995);
xor U5317 (N_5317,N_183,N_3657);
xor U5318 (N_5318,N_1628,N_1113);
nor U5319 (N_5319,N_4140,N_4304);
or U5320 (N_5320,N_4571,N_676);
and U5321 (N_5321,N_2258,N_1034);
xor U5322 (N_5322,N_1333,N_1640);
nand U5323 (N_5323,N_1690,N_1808);
nand U5324 (N_5324,N_764,N_3540);
nor U5325 (N_5325,N_4979,N_298);
nor U5326 (N_5326,N_1661,N_3223);
and U5327 (N_5327,N_706,N_1272);
and U5328 (N_5328,N_1911,N_3924);
nand U5329 (N_5329,N_1982,N_2715);
nand U5330 (N_5330,N_4549,N_369);
and U5331 (N_5331,N_2677,N_970);
xor U5332 (N_5332,N_2935,N_2379);
nor U5333 (N_5333,N_1586,N_3858);
xor U5334 (N_5334,N_4846,N_3516);
nand U5335 (N_5335,N_2809,N_91);
nor U5336 (N_5336,N_2128,N_4447);
nand U5337 (N_5337,N_4319,N_387);
nor U5338 (N_5338,N_2744,N_173);
nand U5339 (N_5339,N_1774,N_874);
xnor U5340 (N_5340,N_661,N_1476);
nand U5341 (N_5341,N_3917,N_3226);
and U5342 (N_5342,N_4292,N_1446);
or U5343 (N_5343,N_3065,N_2531);
nor U5344 (N_5344,N_1102,N_2269);
nand U5345 (N_5345,N_4609,N_4516);
xnor U5346 (N_5346,N_2551,N_811);
and U5347 (N_5347,N_4224,N_4991);
or U5348 (N_5348,N_2179,N_32);
or U5349 (N_5349,N_140,N_2506);
or U5350 (N_5350,N_4000,N_19);
and U5351 (N_5351,N_862,N_109);
and U5352 (N_5352,N_3823,N_3170);
nand U5353 (N_5353,N_1706,N_3771);
or U5354 (N_5354,N_3648,N_4763);
and U5355 (N_5355,N_3358,N_2302);
nand U5356 (N_5356,N_2013,N_1995);
or U5357 (N_5357,N_3113,N_4962);
or U5358 (N_5358,N_4765,N_3202);
nand U5359 (N_5359,N_4364,N_643);
nor U5360 (N_5360,N_22,N_4788);
nor U5361 (N_5361,N_765,N_3889);
xnor U5362 (N_5362,N_438,N_550);
and U5363 (N_5363,N_2499,N_4076);
or U5364 (N_5364,N_4373,N_3072);
nor U5365 (N_5365,N_2692,N_4598);
nand U5366 (N_5366,N_1021,N_4523);
nor U5367 (N_5367,N_3446,N_4767);
xnor U5368 (N_5368,N_1760,N_3155);
or U5369 (N_5369,N_553,N_1265);
and U5370 (N_5370,N_2836,N_1132);
nand U5371 (N_5371,N_1314,N_2253);
xor U5372 (N_5372,N_2884,N_1310);
and U5373 (N_5373,N_3892,N_1962);
and U5374 (N_5374,N_4885,N_1577);
xnor U5375 (N_5375,N_2618,N_3550);
nand U5376 (N_5376,N_3724,N_804);
nand U5377 (N_5377,N_1048,N_3053);
nor U5378 (N_5378,N_945,N_1389);
xnor U5379 (N_5379,N_4611,N_2979);
nand U5380 (N_5380,N_825,N_854);
nor U5381 (N_5381,N_1120,N_1196);
and U5382 (N_5382,N_3760,N_3580);
nand U5383 (N_5383,N_1734,N_2560);
and U5384 (N_5384,N_3929,N_3662);
nand U5385 (N_5385,N_52,N_3337);
nor U5386 (N_5386,N_4404,N_3809);
nor U5387 (N_5387,N_1289,N_3719);
nand U5388 (N_5388,N_2835,N_1324);
xor U5389 (N_5389,N_842,N_4425);
nor U5390 (N_5390,N_3362,N_89);
or U5391 (N_5391,N_1956,N_1873);
or U5392 (N_5392,N_2794,N_3789);
or U5393 (N_5393,N_3498,N_2800);
or U5394 (N_5394,N_3765,N_4952);
nor U5395 (N_5395,N_4208,N_2035);
xnor U5396 (N_5396,N_3264,N_3974);
nand U5397 (N_5397,N_4408,N_1790);
nand U5398 (N_5398,N_942,N_3133);
nand U5399 (N_5399,N_2768,N_2147);
and U5400 (N_5400,N_2339,N_4993);
xnor U5401 (N_5401,N_3168,N_2760);
xnor U5402 (N_5402,N_4542,N_2811);
and U5403 (N_5403,N_1655,N_715);
or U5404 (N_5404,N_81,N_2121);
xnor U5405 (N_5405,N_4197,N_3921);
nand U5406 (N_5406,N_1444,N_4988);
xor U5407 (N_5407,N_3073,N_3637);
nand U5408 (N_5408,N_2186,N_1653);
nor U5409 (N_5409,N_1028,N_2634);
and U5410 (N_5410,N_3220,N_851);
or U5411 (N_5411,N_1240,N_365);
or U5412 (N_5412,N_2468,N_4957);
nor U5413 (N_5413,N_3174,N_386);
nand U5414 (N_5414,N_3606,N_4565);
or U5415 (N_5415,N_26,N_957);
xor U5416 (N_5416,N_1473,N_2089);
nor U5417 (N_5417,N_836,N_2863);
or U5418 (N_5418,N_2959,N_3129);
xnor U5419 (N_5419,N_2038,N_1410);
and U5420 (N_5420,N_3755,N_4473);
xor U5421 (N_5421,N_4492,N_1678);
or U5422 (N_5422,N_214,N_952);
and U5423 (N_5423,N_2578,N_2425);
xnor U5424 (N_5424,N_2291,N_2829);
nand U5425 (N_5425,N_4211,N_3070);
or U5426 (N_5426,N_3288,N_1795);
nor U5427 (N_5427,N_4768,N_291);
xnor U5428 (N_5428,N_3319,N_3578);
and U5429 (N_5429,N_4694,N_39);
or U5430 (N_5430,N_4090,N_4025);
and U5431 (N_5431,N_4535,N_1270);
xnor U5432 (N_5432,N_2070,N_2471);
nor U5433 (N_5433,N_1242,N_557);
and U5434 (N_5434,N_4440,N_3688);
and U5435 (N_5435,N_3355,N_1932);
nor U5436 (N_5436,N_2256,N_2219);
or U5437 (N_5437,N_440,N_1552);
or U5438 (N_5438,N_1296,N_2807);
xor U5439 (N_5439,N_1315,N_4799);
or U5440 (N_5440,N_4637,N_885);
or U5441 (N_5441,N_1527,N_1396);
and U5442 (N_5442,N_3512,N_2989);
or U5443 (N_5443,N_1072,N_2259);
and U5444 (N_5444,N_1362,N_2694);
xnor U5445 (N_5445,N_1506,N_1222);
or U5446 (N_5446,N_4154,N_4244);
or U5447 (N_5447,N_3204,N_2557);
nand U5448 (N_5448,N_2488,N_4948);
nor U5449 (N_5449,N_911,N_3785);
and U5450 (N_5450,N_2198,N_3877);
nor U5451 (N_5451,N_1700,N_898);
or U5452 (N_5452,N_2304,N_2981);
or U5453 (N_5453,N_3638,N_364);
or U5454 (N_5454,N_2230,N_1117);
or U5455 (N_5455,N_1388,N_13);
or U5456 (N_5456,N_4518,N_737);
or U5457 (N_5457,N_3366,N_4043);
nor U5458 (N_5458,N_2246,N_656);
nor U5459 (N_5459,N_1839,N_1696);
or U5460 (N_5460,N_1352,N_4017);
nand U5461 (N_5461,N_2273,N_4356);
nand U5462 (N_5462,N_1281,N_1778);
and U5463 (N_5463,N_1944,N_4528);
or U5464 (N_5464,N_2894,N_1276);
nor U5465 (N_5465,N_4467,N_3171);
or U5466 (N_5466,N_3782,N_511);
and U5467 (N_5467,N_103,N_1820);
nand U5468 (N_5468,N_1407,N_1161);
xor U5469 (N_5469,N_1233,N_2132);
or U5470 (N_5470,N_3882,N_1071);
nor U5471 (N_5471,N_1596,N_3032);
or U5472 (N_5472,N_416,N_1937);
and U5473 (N_5473,N_4713,N_128);
nand U5474 (N_5474,N_2999,N_2529);
nand U5475 (N_5475,N_1693,N_4547);
nor U5476 (N_5476,N_4387,N_441);
nor U5477 (N_5477,N_4235,N_860);
nand U5478 (N_5478,N_4247,N_230);
xor U5479 (N_5479,N_1342,N_4773);
xnor U5480 (N_5480,N_4355,N_3084);
nor U5481 (N_5481,N_1988,N_4118);
or U5482 (N_5482,N_1763,N_4237);
and U5483 (N_5483,N_3977,N_2303);
and U5484 (N_5484,N_1702,N_4281);
nor U5485 (N_5485,N_3893,N_509);
nand U5486 (N_5486,N_4574,N_1639);
nand U5487 (N_5487,N_3,N_810);
or U5488 (N_5488,N_3203,N_196);
xnor U5489 (N_5489,N_556,N_2448);
and U5490 (N_5490,N_4845,N_4661);
xnor U5491 (N_5491,N_2813,N_3927);
and U5492 (N_5492,N_1564,N_4226);
or U5493 (N_5493,N_1866,N_4487);
nand U5494 (N_5494,N_4188,N_989);
or U5495 (N_5495,N_92,N_2910);
xnor U5496 (N_5496,N_798,N_304);
nand U5497 (N_5497,N_3581,N_58);
nand U5498 (N_5498,N_891,N_4001);
nor U5499 (N_5499,N_195,N_3187);
xor U5500 (N_5500,N_3233,N_2200);
and U5501 (N_5501,N_604,N_2722);
xnor U5502 (N_5502,N_3059,N_2309);
nand U5503 (N_5503,N_460,N_4709);
nand U5504 (N_5504,N_3900,N_2313);
or U5505 (N_5505,N_2676,N_505);
nand U5506 (N_5506,N_3740,N_4288);
and U5507 (N_5507,N_747,N_3156);
nand U5508 (N_5508,N_778,N_815);
nor U5509 (N_5509,N_1671,N_1621);
or U5510 (N_5510,N_4310,N_3731);
xor U5511 (N_5511,N_1337,N_3717);
nand U5512 (N_5512,N_3322,N_2424);
or U5513 (N_5513,N_4564,N_2650);
xor U5514 (N_5514,N_2699,N_3367);
nand U5515 (N_5515,N_2433,N_378);
nand U5516 (N_5516,N_4671,N_2347);
xor U5517 (N_5517,N_1618,N_3697);
nor U5518 (N_5518,N_2953,N_4097);
nand U5519 (N_5519,N_1708,N_795);
nor U5520 (N_5520,N_4501,N_250);
and U5521 (N_5521,N_3031,N_3620);
nor U5522 (N_5522,N_2395,N_4433);
and U5523 (N_5523,N_4908,N_2220);
xor U5524 (N_5524,N_892,N_1946);
or U5525 (N_5525,N_966,N_4954);
or U5526 (N_5526,N_4191,N_3834);
and U5527 (N_5527,N_2308,N_2311);
xnor U5528 (N_5528,N_159,N_4588);
xor U5529 (N_5529,N_401,N_1896);
nand U5530 (N_5530,N_2438,N_502);
or U5531 (N_5531,N_4151,N_3190);
and U5532 (N_5532,N_577,N_770);
or U5533 (N_5533,N_185,N_3468);
nand U5534 (N_5534,N_1041,N_4888);
and U5535 (N_5535,N_1387,N_3718);
nand U5536 (N_5536,N_641,N_1742);
nor U5537 (N_5537,N_3542,N_4020);
or U5538 (N_5538,N_1419,N_4864);
xnor U5539 (N_5539,N_2958,N_4263);
and U5540 (N_5540,N_3042,N_2372);
nor U5541 (N_5541,N_2329,N_3449);
and U5542 (N_5542,N_2763,N_220);
nand U5543 (N_5543,N_4098,N_2180);
and U5544 (N_5544,N_3806,N_1403);
nand U5545 (N_5545,N_2422,N_3237);
xor U5546 (N_5546,N_4909,N_4214);
or U5547 (N_5547,N_4353,N_3950);
xor U5548 (N_5548,N_49,N_423);
nand U5549 (N_5549,N_3626,N_3861);
or U5550 (N_5550,N_3668,N_3807);
and U5551 (N_5551,N_4105,N_1143);
xor U5552 (N_5552,N_4383,N_1672);
nand U5553 (N_5553,N_517,N_1447);
nand U5554 (N_5554,N_124,N_779);
xnor U5555 (N_5555,N_2649,N_2238);
xnor U5556 (N_5556,N_2033,N_3193);
and U5557 (N_5557,N_616,N_4690);
nor U5558 (N_5558,N_16,N_2786);
and U5559 (N_5559,N_290,N_864);
nand U5560 (N_5560,N_4706,N_463);
or U5561 (N_5561,N_3303,N_2621);
and U5562 (N_5562,N_962,N_2980);
nand U5563 (N_5563,N_1489,N_3574);
nor U5564 (N_5564,N_2097,N_4648);
and U5565 (N_5565,N_3830,N_2095);
xnor U5566 (N_5566,N_1583,N_248);
and U5567 (N_5567,N_1569,N_2145);
nor U5568 (N_5568,N_4095,N_1753);
nor U5569 (N_5569,N_200,N_516);
xnor U5570 (N_5570,N_2757,N_1408);
or U5571 (N_5571,N_1603,N_23);
or U5572 (N_5572,N_1451,N_1526);
nand U5573 (N_5573,N_2214,N_318);
nand U5574 (N_5574,N_1391,N_2162);
or U5575 (N_5575,N_4822,N_4143);
or U5576 (N_5576,N_238,N_2969);
or U5577 (N_5577,N_2965,N_2571);
or U5578 (N_5578,N_1024,N_4298);
nand U5579 (N_5579,N_3656,N_1254);
and U5580 (N_5580,N_958,N_4532);
nand U5581 (N_5581,N_3548,N_648);
nand U5582 (N_5582,N_410,N_4485);
and U5583 (N_5583,N_2718,N_822);
nor U5584 (N_5584,N_2568,N_1717);
or U5585 (N_5585,N_3988,N_2726);
or U5586 (N_5586,N_2389,N_129);
nand U5587 (N_5587,N_3191,N_1687);
nor U5588 (N_5588,N_4166,N_2324);
nor U5589 (N_5589,N_3702,N_4334);
or U5590 (N_5590,N_2325,N_3044);
nand U5591 (N_5591,N_1079,N_1897);
nand U5592 (N_5592,N_68,N_4786);
nand U5593 (N_5593,N_1057,N_2821);
nand U5594 (N_5594,N_3937,N_4723);
nor U5595 (N_5595,N_4142,N_4283);
nor U5596 (N_5596,N_4842,N_1695);
xor U5597 (N_5597,N_3692,N_749);
xor U5598 (N_5598,N_2495,N_2799);
or U5599 (N_5599,N_1913,N_1399);
xor U5600 (N_5600,N_202,N_902);
and U5601 (N_5601,N_424,N_3689);
nand U5602 (N_5602,N_2864,N_3272);
or U5603 (N_5603,N_125,N_3241);
xnor U5604 (N_5604,N_3038,N_1784);
and U5605 (N_5605,N_3360,N_2236);
xnor U5606 (N_5606,N_3549,N_3388);
nand U5607 (N_5607,N_3235,N_2357);
or U5608 (N_5608,N_1869,N_4445);
xor U5609 (N_5609,N_2915,N_1893);
xor U5610 (N_5610,N_895,N_2312);
nor U5611 (N_5611,N_3424,N_4915);
nand U5612 (N_5612,N_787,N_4789);
or U5613 (N_5613,N_2961,N_2825);
and U5614 (N_5614,N_237,N_4578);
nand U5615 (N_5615,N_827,N_2674);
and U5616 (N_5616,N_3239,N_4393);
nand U5617 (N_5617,N_4654,N_4212);
xor U5618 (N_5618,N_834,N_4797);
nand U5619 (N_5619,N_4495,N_530);
and U5620 (N_5620,N_182,N_920);
and U5621 (N_5621,N_144,N_80);
nand U5622 (N_5622,N_1493,N_4708);
xor U5623 (N_5623,N_2742,N_4216);
and U5624 (N_5624,N_1907,N_4031);
and U5625 (N_5625,N_2232,N_948);
xnor U5626 (N_5626,N_3140,N_3862);
nor U5627 (N_5627,N_928,N_163);
xnor U5628 (N_5628,N_63,N_2814);
and U5629 (N_5629,N_1416,N_2704);
nor U5630 (N_5630,N_4730,N_2820);
or U5631 (N_5631,N_4984,N_1898);
xnor U5632 (N_5632,N_2507,N_3186);
nor U5633 (N_5633,N_411,N_1978);
nor U5634 (N_5634,N_3248,N_4600);
or U5635 (N_5635,N_4457,N_24);
nor U5636 (N_5636,N_3091,N_2923);
nand U5637 (N_5637,N_1116,N_1415);
and U5638 (N_5638,N_4617,N_4602);
nand U5639 (N_5639,N_493,N_2352);
and U5640 (N_5640,N_2613,N_2360);
nor U5641 (N_5641,N_2109,N_218);
nor U5642 (N_5642,N_1025,N_4683);
or U5643 (N_5643,N_2454,N_1312);
nand U5644 (N_5644,N_3919,N_926);
nand U5645 (N_5645,N_2957,N_1934);
or U5646 (N_5646,N_4514,N_1158);
xor U5647 (N_5647,N_3324,N_1477);
or U5648 (N_5648,N_3905,N_4615);
and U5649 (N_5649,N_3531,N_2777);
or U5650 (N_5650,N_2274,N_4410);
xor U5651 (N_5651,N_4975,N_4427);
nor U5652 (N_5652,N_4455,N_3695);
nand U5653 (N_5653,N_2680,N_1418);
xnor U5654 (N_5654,N_1865,N_4854);
nand U5655 (N_5655,N_4033,N_1255);
nor U5656 (N_5656,N_838,N_555);
nand U5657 (N_5657,N_932,N_349);
xor U5658 (N_5658,N_2869,N_4946);
and U5659 (N_5659,N_2686,N_2769);
or U5660 (N_5660,N_1765,N_1355);
xnor U5661 (N_5661,N_515,N_4660);
or U5662 (N_5662,N_2645,N_36);
or U5663 (N_5663,N_2891,N_3266);
and U5664 (N_5664,N_4577,N_3434);
or U5665 (N_5665,N_3159,N_3125);
or U5666 (N_5666,N_4696,N_4625);
nor U5667 (N_5667,N_3930,N_435);
and U5668 (N_5668,N_2449,N_2525);
or U5669 (N_5669,N_4205,N_117);
xor U5670 (N_5670,N_1522,N_2209);
nor U5671 (N_5671,N_790,N_1436);
and U5672 (N_5672,N_1633,N_313);
or U5673 (N_5673,N_4606,N_2934);
nand U5674 (N_5674,N_3518,N_1052);
nor U5675 (N_5675,N_2972,N_1591);
xor U5676 (N_5676,N_4030,N_271);
xor U5677 (N_5677,N_919,N_1985);
and U5678 (N_5678,N_1571,N_2888);
and U5679 (N_5679,N_351,N_2364);
xor U5680 (N_5680,N_2491,N_1590);
or U5681 (N_5681,N_4736,N_3976);
and U5682 (N_5682,N_4236,N_978);
and U5683 (N_5683,N_1632,N_357);
or U5684 (N_5684,N_809,N_2601);
nand U5685 (N_5685,N_784,N_2527);
xor U5686 (N_5686,N_4777,N_708);
nand U5687 (N_5687,N_400,N_3727);
xnor U5688 (N_5688,N_3295,N_767);
xor U5689 (N_5689,N_1115,N_4141);
and U5690 (N_5690,N_3847,N_1890);
and U5691 (N_5691,N_3457,N_4563);
nor U5692 (N_5692,N_3286,N_4204);
xor U5693 (N_5693,N_1334,N_3301);
or U5694 (N_5694,N_373,N_3247);
or U5695 (N_5695,N_3737,N_2388);
and U5696 (N_5696,N_1173,N_3488);
or U5697 (N_5697,N_4361,N_1916);
or U5698 (N_5698,N_1871,N_3212);
nor U5699 (N_5699,N_1666,N_2175);
and U5700 (N_5700,N_2587,N_2535);
nand U5701 (N_5701,N_1587,N_3117);
nand U5702 (N_5702,N_1559,N_41);
or U5703 (N_5703,N_2305,N_3786);
nor U5704 (N_5704,N_476,N_3653);
and U5705 (N_5705,N_587,N_1615);
xor U5706 (N_5706,N_2103,N_4358);
and U5707 (N_5707,N_4647,N_1889);
and U5708 (N_5708,N_3969,N_988);
and U5709 (N_5709,N_146,N_3006);
nand U5710 (N_5710,N_499,N_3208);
xnor U5711 (N_5711,N_339,N_4850);
and U5712 (N_5712,N_627,N_1761);
and U5713 (N_5713,N_3216,N_1566);
nand U5714 (N_5714,N_3419,N_2144);
or U5715 (N_5715,N_2077,N_2602);
and U5716 (N_5716,N_380,N_4646);
xnor U5717 (N_5717,N_1297,N_3040);
nor U5718 (N_5718,N_1731,N_3951);
and U5719 (N_5719,N_154,N_178);
xor U5720 (N_5720,N_1938,N_2974);
and U5721 (N_5721,N_4094,N_3074);
and U5722 (N_5722,N_1204,N_2191);
or U5723 (N_5723,N_987,N_896);
nand U5724 (N_5724,N_1063,N_669);
xor U5725 (N_5725,N_1300,N_1186);
or U5726 (N_5726,N_1164,N_855);
and U5727 (N_5727,N_6,N_2106);
xor U5728 (N_5728,N_3185,N_2419);
or U5729 (N_5729,N_852,N_2287);
or U5730 (N_5730,N_285,N_2463);
nand U5731 (N_5731,N_210,N_2591);
or U5732 (N_5732,N_2565,N_3126);
nor U5733 (N_5733,N_1967,N_2713);
nor U5734 (N_5734,N_276,N_4014);
and U5735 (N_5735,N_4061,N_3296);
or U5736 (N_5736,N_4520,N_31);
and U5737 (N_5737,N_3707,N_4716);
and U5738 (N_5738,N_2666,N_1727);
nor U5739 (N_5739,N_2789,N_2262);
or U5740 (N_5740,N_2377,N_1500);
xor U5741 (N_5741,N_1812,N_2194);
nand U5742 (N_5742,N_2174,N_2299);
nor U5743 (N_5743,N_2950,N_3649);
or U5744 (N_5744,N_21,N_4849);
xor U5745 (N_5745,N_2656,N_3245);
and U5746 (N_5746,N_2203,N_3320);
and U5747 (N_5747,N_635,N_412);
xnor U5748 (N_5748,N_3410,N_2310);
nand U5749 (N_5749,N_2717,N_2041);
and U5750 (N_5750,N_4558,N_923);
nand U5751 (N_5751,N_3475,N_2153);
or U5752 (N_5752,N_4376,N_4144);
and U5753 (N_5753,N_760,N_322);
and U5754 (N_5754,N_2407,N_161);
nand U5755 (N_5755,N_999,N_334);
nor U5756 (N_5756,N_2626,N_2051);
or U5757 (N_5757,N_2373,N_4505);
or U5758 (N_5758,N_3496,N_4418);
nor U5759 (N_5759,N_2090,N_3469);
or U5760 (N_5760,N_3867,N_450);
and U5761 (N_5761,N_2410,N_2582);
nor U5762 (N_5762,N_1903,N_2251);
nor U5763 (N_5763,N_1787,N_703);
or U5764 (N_5764,N_72,N_865);
or U5765 (N_5765,N_1216,N_3109);
nor U5766 (N_5766,N_3716,N_1171);
and U5767 (N_5767,N_2751,N_1612);
or U5768 (N_5768,N_3625,N_4414);
and U5769 (N_5769,N_1286,N_4969);
or U5770 (N_5770,N_3050,N_38);
and U5771 (N_5771,N_4106,N_1345);
nand U5772 (N_5772,N_2062,N_1027);
nand U5773 (N_5773,N_4354,N_3321);
and U5774 (N_5774,N_3030,N_408);
or U5775 (N_5775,N_2337,N_3918);
nor U5776 (N_5776,N_2185,N_2927);
nand U5777 (N_5777,N_670,N_3472);
nor U5778 (N_5778,N_4745,N_4475);
or U5779 (N_5779,N_292,N_3928);
and U5780 (N_5780,N_3704,N_3818);
or U5781 (N_5781,N_600,N_2);
nand U5782 (N_5782,N_2476,N_4820);
xor U5783 (N_5783,N_3832,N_1005);
or U5784 (N_5784,N_4645,N_4344);
xor U5785 (N_5785,N_497,N_2474);
xnor U5786 (N_5786,N_2903,N_1688);
nand U5787 (N_5787,N_950,N_3935);
nor U5788 (N_5788,N_2020,N_4903);
and U5789 (N_5789,N_4956,N_1458);
nand U5790 (N_5790,N_768,N_3746);
and U5791 (N_5791,N_752,N_208);
xor U5792 (N_5792,N_4689,N_1015);
nand U5793 (N_5793,N_3344,N_362);
nor U5794 (N_5794,N_1570,N_2773);
and U5795 (N_5795,N_1056,N_729);
nor U5796 (N_5796,N_3914,N_43);
or U5797 (N_5797,N_3490,N_3551);
nor U5798 (N_5798,N_1535,N_4780);
nor U5799 (N_5799,N_2189,N_1764);
nor U5800 (N_5800,N_425,N_3471);
xnor U5801 (N_5801,N_3661,N_4996);
xnor U5802 (N_5802,N_3735,N_592);
nand U5803 (N_5803,N_3543,N_3505);
or U5804 (N_5804,N_4787,N_654);
nor U5805 (N_5805,N_2375,N_1804);
and U5806 (N_5806,N_2064,N_4700);
and U5807 (N_5807,N_3705,N_4684);
and U5808 (N_5808,N_4245,N_4294);
xnor U5809 (N_5809,N_538,N_2301);
and U5810 (N_5810,N_2233,N_756);
nor U5811 (N_5811,N_2815,N_256);
or U5812 (N_5812,N_3312,N_1533);
xor U5813 (N_5813,N_2250,N_4336);
nor U5814 (N_5814,N_2216,N_4295);
xor U5815 (N_5815,N_4172,N_662);
and U5816 (N_5816,N_3837,N_289);
nand U5817 (N_5817,N_2349,N_3990);
xor U5818 (N_5818,N_2055,N_2843);
or U5819 (N_5819,N_3780,N_2486);
nand U5820 (N_5820,N_37,N_796);
nor U5821 (N_5821,N_1134,N_771);
and U5822 (N_5822,N_4497,N_843);
and U5823 (N_5823,N_308,N_802);
or U5824 (N_5824,N_2651,N_3934);
nor U5825 (N_5825,N_2105,N_2741);
and U5826 (N_5826,N_819,N_1617);
nor U5827 (N_5827,N_3641,N_1322);
xor U5828 (N_5828,N_3992,N_3576);
and U5829 (N_5829,N_1965,N_3012);
xnor U5830 (N_5830,N_465,N_3902);
nor U5831 (N_5831,N_718,N_973);
nand U5832 (N_5832,N_385,N_3843);
nand U5833 (N_5833,N_4537,N_330);
nand U5834 (N_5834,N_1592,N_1963);
and U5835 (N_5835,N_637,N_3558);
and U5836 (N_5836,N_2520,N_3949);
xor U5837 (N_5837,N_3579,N_2907);
or U5838 (N_5838,N_4267,N_4347);
nand U5839 (N_5839,N_2143,N_4703);
nand U5840 (N_5840,N_2719,N_930);
nor U5841 (N_5841,N_2655,N_1974);
or U5842 (N_5842,N_3217,N_3926);
or U5843 (N_5843,N_4711,N_3687);
or U5844 (N_5844,N_4365,N_3784);
xnor U5845 (N_5845,N_1424,N_2212);
or U5846 (N_5846,N_3957,N_4307);
xor U5847 (N_5847,N_759,N_4423);
and U5848 (N_5848,N_388,N_4053);
and U5849 (N_5849,N_4500,N_2548);
or U5850 (N_5850,N_2430,N_3121);
xor U5851 (N_5851,N_2684,N_2765);
xor U5852 (N_5852,N_1748,N_916);
and U5853 (N_5853,N_3341,N_1180);
xor U5854 (N_5854,N_2188,N_2920);
or U5855 (N_5855,N_4910,N_1877);
xor U5856 (N_5856,N_2852,N_758);
nand U5857 (N_5857,N_1971,N_3137);
xor U5858 (N_5858,N_4075,N_2662);
nor U5859 (N_5859,N_4860,N_782);
and U5860 (N_5860,N_3564,N_2343);
xnor U5861 (N_5861,N_4359,N_4562);
xor U5862 (N_5862,N_2630,N_4887);
xor U5863 (N_5863,N_2370,N_617);
nand U5864 (N_5864,N_4146,N_1654);
nand U5865 (N_5865,N_506,N_2493);
nor U5866 (N_5866,N_699,N_801);
nor U5867 (N_5867,N_565,N_3933);
nand U5868 (N_5868,N_4801,N_1112);
nor U5869 (N_5869,N_1453,N_3014);
xnor U5870 (N_5870,N_1004,N_1860);
nand U5871 (N_5871,N_1125,N_1172);
nand U5872 (N_5872,N_1230,N_755);
and U5873 (N_5873,N_720,N_2752);
or U5874 (N_5874,N_2878,N_1450);
nand U5875 (N_5875,N_3062,N_1235);
xnor U5876 (N_5876,N_4739,N_4792);
or U5877 (N_5877,N_332,N_4133);
nor U5878 (N_5878,N_481,N_392);
nor U5879 (N_5879,N_1719,N_1588);
and U5880 (N_5880,N_3289,N_1332);
nand U5881 (N_5881,N_3629,N_3001);
nand U5882 (N_5882,N_3282,N_2397);
xnor U5883 (N_5883,N_1082,N_3438);
and U5884 (N_5884,N_246,N_1409);
nor U5885 (N_5885,N_2862,N_1721);
or U5886 (N_5886,N_226,N_4100);
or U5887 (N_5887,N_3872,N_4092);
or U5888 (N_5888,N_2123,N_2496);
or U5889 (N_5889,N_1293,N_2941);
and U5890 (N_5890,N_1092,N_1437);
nor U5891 (N_5891,N_2991,N_1604);
nand U5892 (N_5892,N_1711,N_3194);
nand U5893 (N_5893,N_2093,N_3936);
xor U5894 (N_5894,N_1925,N_4275);
and U5895 (N_5895,N_625,N_610);
xor U5896 (N_5896,N_1213,N_1543);
or U5897 (N_5897,N_2558,N_3940);
or U5898 (N_5898,N_171,N_1049);
nor U5899 (N_5899,N_4056,N_1100);
xor U5900 (N_5900,N_1022,N_4838);
nand U5901 (N_5901,N_863,N_2117);
or U5902 (N_5902,N_1741,N_3331);
or U5903 (N_5903,N_2196,N_84);
xnor U5904 (N_5904,N_3593,N_1144);
nand U5905 (N_5905,N_4744,N_1178);
nand U5906 (N_5906,N_2321,N_325);
nor U5907 (N_5907,N_3064,N_594);
nand U5908 (N_5908,N_443,N_2932);
nor U5909 (N_5909,N_104,N_2428);
or U5910 (N_5910,N_3863,N_430);
nor U5911 (N_5911,N_3010,N_740);
or U5912 (N_5912,N_4232,N_3011);
xor U5913 (N_5913,N_1799,N_120);
and U5914 (N_5914,N_2279,N_181);
nand U5915 (N_5915,N_3249,N_2017);
xor U5916 (N_5916,N_3418,N_3308);
and U5917 (N_5917,N_2019,N_2633);
nor U5918 (N_5918,N_3416,N_4512);
xnor U5919 (N_5919,N_4762,N_4379);
or U5920 (N_5920,N_498,N_789);
nand U5921 (N_5921,N_2532,N_4164);
nor U5922 (N_5922,N_2183,N_442);
xor U5923 (N_5923,N_1449,N_4884);
or U5924 (N_5924,N_3880,N_2962);
nor U5925 (N_5925,N_3136,N_3157);
xnor U5926 (N_5926,N_2614,N_2550);
xnor U5927 (N_5927,N_490,N_3525);
or U5928 (N_5928,N_3757,N_3478);
xnor U5929 (N_5929,N_4007,N_100);
nand U5930 (N_5930,N_2866,N_1779);
nand U5931 (N_5931,N_1858,N_3376);
xnor U5932 (N_5932,N_300,N_4900);
and U5933 (N_5933,N_2122,N_2453);
or U5934 (N_5934,N_2348,N_1192);
and U5935 (N_5935,N_3887,N_921);
xnor U5936 (N_5936,N_965,N_2009);
and U5937 (N_5937,N_329,N_4509);
or U5938 (N_5938,N_354,N_4008);
and U5939 (N_5939,N_4942,N_4733);
and U5940 (N_5940,N_1926,N_3904);
or U5941 (N_5941,N_4348,N_2163);
or U5942 (N_5942,N_1524,N_3759);
xor U5943 (N_5943,N_4930,N_3176);
nand U5944 (N_5944,N_448,N_4179);
nand U5945 (N_5945,N_2735,N_2345);
nand U5946 (N_5946,N_1271,N_2919);
nor U5947 (N_5947,N_4758,N_3630);
nand U5948 (N_5948,N_4055,N_4734);
xnor U5949 (N_5949,N_853,N_4966);
and U5950 (N_5950,N_915,N_3980);
nand U5951 (N_5951,N_2750,N_1457);
xor U5952 (N_5952,N_612,N_571);
nand U5953 (N_5953,N_1794,N_1826);
xor U5954 (N_5954,N_2336,N_947);
and U5955 (N_5955,N_1381,N_1226);
nor U5956 (N_5956,N_1351,N_603);
xnor U5957 (N_5957,N_2609,N_1377);
xnor U5958 (N_5958,N_780,N_1363);
nand U5959 (N_5959,N_4757,N_4453);
or U5960 (N_5960,N_309,N_3314);
or U5961 (N_5961,N_994,N_4870);
or U5962 (N_5962,N_2976,N_2400);
nand U5963 (N_5963,N_4775,N_1947);
and U5964 (N_5964,N_2883,N_1199);
or U5965 (N_5965,N_4413,N_1266);
nor U5966 (N_5966,N_1058,N_3340);
nor U5967 (N_5967,N_1811,N_4624);
nand U5968 (N_5968,N_2393,N_3745);
and U5969 (N_5969,N_3885,N_1622);
nor U5970 (N_5970,N_2992,N_4806);
nor U5971 (N_5971,N_3236,N_1643);
xor U5972 (N_5972,N_4066,N_3339);
or U5973 (N_5973,N_1776,N_1151);
and U5974 (N_5974,N_3583,N_114);
and U5975 (N_5975,N_494,N_2795);
xor U5976 (N_5976,N_1750,N_791);
or U5977 (N_5977,N_532,N_1601);
nand U5978 (N_5978,N_2223,N_2802);
and U5979 (N_5979,N_1665,N_2997);
xnor U5980 (N_5980,N_1441,N_3066);
nand U5981 (N_5981,N_2776,N_2739);
xor U5982 (N_5982,N_2573,N_2975);
xnor U5983 (N_5983,N_4790,N_4938);
and U5984 (N_5984,N_3333,N_3947);
nor U5985 (N_5985,N_826,N_4559);
and U5986 (N_5986,N_4135,N_143);
nand U5987 (N_5987,N_4126,N_3506);
nor U5988 (N_5988,N_3590,N_961);
xnor U5989 (N_5989,N_3570,N_3615);
or U5990 (N_5990,N_3604,N_1573);
nand U5991 (N_5991,N_4999,N_4005);
nand U5992 (N_5992,N_4980,N_302);
or U5993 (N_5993,N_4394,N_345);
and U5994 (N_5994,N_711,N_4573);
nand U5995 (N_5995,N_3989,N_870);
and U5996 (N_5996,N_3679,N_4685);
xor U5997 (N_5997,N_2451,N_2622);
and U5998 (N_5998,N_3713,N_2575);
nor U5999 (N_5999,N_99,N_275);
xnor U6000 (N_6000,N_1040,N_946);
xor U6001 (N_6001,N_1009,N_2005);
or U6002 (N_6002,N_2319,N_444);
nor U6003 (N_6003,N_3665,N_3821);
and U6004 (N_6004,N_1827,N_4168);
xor U6005 (N_6005,N_1460,N_2142);
or U6006 (N_6006,N_4184,N_4277);
or U6007 (N_6007,N_3592,N_1652);
and U6008 (N_6008,N_4229,N_2260);
xnor U6009 (N_6009,N_3443,N_65);
nand U6010 (N_6010,N_4728,N_1728);
nand U6011 (N_6011,N_917,N_4856);
nand U6012 (N_6012,N_3997,N_3544);
or U6013 (N_6013,N_1074,N_2581);
nor U6014 (N_6014,N_2447,N_3374);
or U6015 (N_6015,N_4308,N_2046);
nor U6016 (N_6016,N_1796,N_2597);
or U6017 (N_6017,N_1481,N_1979);
or U6018 (N_6018,N_2455,N_4978);
nor U6019 (N_6019,N_1999,N_4274);
and U6020 (N_6020,N_3115,N_4526);
nor U6021 (N_6021,N_3810,N_984);
or U6022 (N_6022,N_3489,N_1755);
nand U6023 (N_6023,N_4371,N_1994);
and U6024 (N_6024,N_4115,N_2015);
nand U6025 (N_6025,N_1961,N_3146);
nor U6026 (N_6026,N_3445,N_1059);
nand U6027 (N_6027,N_2767,N_2411);
xor U6028 (N_6028,N_2758,N_638);
and U6029 (N_6029,N_2870,N_1791);
xnor U6030 (N_6030,N_4967,N_3483);
nand U6031 (N_6031,N_631,N_4839);
nand U6032 (N_6032,N_1738,N_615);
nand U6033 (N_6033,N_3738,N_652);
and U6034 (N_6034,N_2118,N_1682);
and U6035 (N_6035,N_350,N_3485);
nand U6036 (N_6036,N_429,N_4919);
nand U6037 (N_6037,N_2363,N_1899);
nor U6038 (N_6038,N_3259,N_500);
nand U6039 (N_6039,N_2738,N_1066);
xor U6040 (N_6040,N_512,N_1507);
xnor U6041 (N_6041,N_4431,N_2139);
nor U6042 (N_6042,N_2664,N_2521);
nand U6043 (N_6043,N_2104,N_4022);
or U6044 (N_6044,N_4280,N_2873);
xnor U6045 (N_6045,N_3164,N_2056);
nor U6046 (N_6046,N_204,N_3105);
nor U6047 (N_6047,N_3831,N_2537);
nand U6048 (N_6048,N_2667,N_4965);
nand U6049 (N_6049,N_287,N_3346);
xnor U6050 (N_6050,N_1759,N_249);
or U6051 (N_6051,N_3618,N_1558);
xor U6052 (N_6052,N_491,N_3849);
and U6053 (N_6053,N_3572,N_1733);
xnor U6054 (N_6054,N_3993,N_3891);
or U6055 (N_6055,N_2460,N_1917);
xor U6056 (N_6056,N_1854,N_1800);
xor U6057 (N_6057,N_57,N_1878);
nand U6058 (N_6058,N_2501,N_2906);
and U6059 (N_6059,N_4269,N_3973);
nor U6060 (N_6060,N_2712,N_622);
and U6061 (N_6061,N_2971,N_3095);
nor U6062 (N_6062,N_1221,N_3546);
or U6063 (N_6063,N_3058,N_981);
and U6064 (N_6064,N_177,N_1468);
and U6065 (N_6065,N_4862,N_3128);
or U6066 (N_6066,N_2205,N_3451);
and U6067 (N_6067,N_2365,N_2306);
or U6068 (N_6068,N_3036,N_2648);
and U6069 (N_6069,N_873,N_2678);
nand U6070 (N_6070,N_766,N_1704);
nand U6071 (N_6071,N_4881,N_3448);
or U6072 (N_6072,N_4561,N_3481);
nand U6073 (N_6073,N_3622,N_134);
nor U6074 (N_6074,N_4779,N_1855);
or U6075 (N_6075,N_823,N_3828);
nand U6076 (N_6076,N_1133,N_1176);
nand U6077 (N_6077,N_4958,N_3805);
nand U6078 (N_6078,N_1338,N_1256);
nor U6079 (N_6079,N_4253,N_2327);
xor U6080 (N_6080,N_4296,N_1542);
nand U6081 (N_6081,N_1549,N_4360);
nor U6082 (N_6082,N_3206,N_990);
nand U6083 (N_6083,N_1294,N_3955);
or U6084 (N_6084,N_4420,N_1638);
and U6085 (N_6085,N_1075,N_2006);
and U6086 (N_6086,N_1433,N_3447);
nor U6087 (N_6087,N_4955,N_2596);
and U6088 (N_6088,N_2234,N_1782);
nand U6089 (N_6089,N_1605,N_3864);
xnor U6090 (N_6090,N_3088,N_4818);
and U6091 (N_6091,N_484,N_2458);
nor U6092 (N_6092,N_608,N_2512);
xor U6093 (N_6093,N_3654,N_3348);
and U6094 (N_6094,N_3753,N_2564);
xor U6095 (N_6095,N_4719,N_2265);
or U6096 (N_6096,N_2159,N_4198);
nor U6097 (N_6097,N_3464,N_3369);
or U6098 (N_6098,N_2173,N_2671);
nand U6099 (N_6099,N_1421,N_3826);
xnor U6100 (N_6100,N_315,N_268);
nand U6101 (N_6101,N_261,N_3770);
and U6102 (N_6102,N_518,N_2711);
and U6103 (N_6103,N_3315,N_4107);
and U6104 (N_6104,N_1308,N_3846);
and U6105 (N_6105,N_4612,N_3979);
or U6106 (N_6106,N_3046,N_1939);
or U6107 (N_6107,N_167,N_138);
or U6108 (N_6108,N_1611,N_630);
nand U6109 (N_6109,N_1335,N_4058);
xor U6110 (N_6110,N_4970,N_3152);
nor U6111 (N_6111,N_2086,N_2748);
xnor U6112 (N_6112,N_1014,N_845);
and U6113 (N_6113,N_4873,N_229);
and U6114 (N_6114,N_623,N_2624);
nand U6115 (N_6115,N_879,N_4234);
xnor U6116 (N_6116,N_4717,N_1885);
nor U6117 (N_6117,N_1442,N_3200);
nand U6118 (N_6118,N_2367,N_2054);
nand U6119 (N_6119,N_374,N_1857);
xor U6120 (N_6120,N_3801,N_1928);
and U6121 (N_6121,N_533,N_1055);
nor U6122 (N_6122,N_2225,N_4907);
nand U6123 (N_6123,N_4582,N_492);
or U6124 (N_6124,N_964,N_975);
nand U6125 (N_6125,N_1901,N_4138);
nor U6126 (N_6126,N_2837,N_572);
xor U6127 (N_6127,N_3382,N_3696);
nand U6128 (N_6128,N_4285,N_844);
or U6129 (N_6129,N_644,N_4346);
xor U6130 (N_6130,N_4550,N_1285);
or U6131 (N_6131,N_2416,N_4207);
nor U6132 (N_6132,N_1887,N_405);
nor U6133 (N_6133,N_1306,N_3616);
nand U6134 (N_6134,N_258,N_3177);
nand U6135 (N_6135,N_1775,N_3000);
xnor U6136 (N_6136,N_1008,N_4368);
xor U6137 (N_6137,N_4323,N_1175);
nand U6138 (N_6138,N_2818,N_4810);
nor U6139 (N_6139,N_403,N_25);
nand U6140 (N_6140,N_828,N_4325);
xor U6141 (N_6141,N_1000,N_1519);
nor U6142 (N_6142,N_4342,N_3503);
xor U6143 (N_6143,N_4386,N_4629);
xor U6144 (N_6144,N_2473,N_1146);
nor U6145 (N_6145,N_4441,N_242);
nand U6146 (N_6146,N_3897,N_3995);
xor U6147 (N_6147,N_105,N_4155);
nand U6148 (N_6148,N_3426,N_203);
nand U6149 (N_6149,N_1707,N_1358);
or U6150 (N_6150,N_3857,N_1948);
xor U6151 (N_6151,N_4940,N_2396);
or U6152 (N_6152,N_1081,N_618);
xor U6153 (N_6153,N_613,N_126);
and U6154 (N_6154,N_4951,N_3684);
nor U6155 (N_6155,N_2160,N_2036);
or U6156 (N_6156,N_4776,N_2937);
nand U6157 (N_6157,N_4941,N_3643);
xor U6158 (N_6158,N_4153,N_3938);
xnor U6159 (N_6159,N_4201,N_3279);
and U6160 (N_6160,N_95,N_3743);
nor U6161 (N_6161,N_4515,N_1325);
nand U6162 (N_6162,N_1236,N_4720);
and U6163 (N_6163,N_1061,N_1426);
or U6164 (N_6164,N_4619,N_2264);
nand U6165 (N_6165,N_925,N_761);
or U6166 (N_6166,N_4464,N_797);
nand U6167 (N_6167,N_4626,N_130);
nor U6168 (N_6168,N_1579,N_3037);
or U6169 (N_6169,N_1973,N_3886);
or U6170 (N_6170,N_3775,N_225);
nand U6171 (N_6171,N_4282,N_4770);
nand U6172 (N_6172,N_4189,N_833);
and U6173 (N_6173,N_2285,N_561);
or U6174 (N_6174,N_2380,N_1087);
and U6175 (N_6175,N_980,N_2298);
xor U6176 (N_6176,N_2629,N_829);
nor U6177 (N_6177,N_3406,N_1536);
and U6178 (N_6178,N_4572,N_653);
xor U6179 (N_6179,N_164,N_4791);
and U6180 (N_6180,N_2135,N_4465);
nor U6181 (N_6181,N_4367,N_3987);
xor U6182 (N_6182,N_1220,N_2698);
and U6183 (N_6183,N_1386,N_1798);
or U6184 (N_6184,N_3381,N_4230);
nand U6185 (N_6185,N_3850,N_4051);
nand U6186 (N_6186,N_701,N_259);
nand U6187 (N_6187,N_595,N_4678);
nand U6188 (N_6188,N_2612,N_1958);
and U6189 (N_6189,N_1019,N_803);
xnor U6190 (N_6190,N_2227,N_1350);
xor U6191 (N_6191,N_4202,N_1709);
nand U6192 (N_6192,N_536,N_4398);
nand U6193 (N_6193,N_397,N_4868);
or U6194 (N_6194,N_2037,N_4436);
nor U6195 (N_6195,N_3184,N_1989);
and U6196 (N_6196,N_2562,N_4778);
nand U6197 (N_6197,N_1375,N_221);
xnor U6198 (N_6198,N_2076,N_1343);
nor U6199 (N_6199,N_4494,N_50);
nand U6200 (N_6200,N_554,N_348);
nor U6201 (N_6201,N_2538,N_4366);
or U6202 (N_6202,N_821,N_4309);
or U6203 (N_6203,N_2530,N_4452);
nand U6204 (N_6204,N_2759,N_2113);
and U6205 (N_6205,N_3591,N_998);
xnor U6206 (N_6206,N_3681,N_573);
or U6207 (N_6207,N_355,N_3795);
nor U6208 (N_6208,N_4037,N_3143);
and U6209 (N_6209,N_3671,N_4673);
xor U6210 (N_6210,N_4830,N_282);
and U6211 (N_6211,N_954,N_4084);
or U6212 (N_6212,N_2237,N_806);
nor U6213 (N_6213,N_1904,N_2652);
and U6214 (N_6214,N_2636,N_3326);
nand U6215 (N_6215,N_264,N_1035);
or U6216 (N_6216,N_191,N_585);
nand U6217 (N_6217,N_111,N_3594);
nand U6218 (N_6218,N_1011,N_193);
nor U6219 (N_6219,N_991,N_4293);
and U6220 (N_6220,N_813,N_4177);
and U6221 (N_6221,N_2709,N_363);
and U6222 (N_6222,N_2877,N_399);
xor U6223 (N_6223,N_2778,N_1563);
nand U6224 (N_6224,N_235,N_2351);
or U6225 (N_6225,N_3816,N_2823);
and U6226 (N_6226,N_2466,N_3792);
nand U6227 (N_6227,N_4192,N_172);
xnor U6228 (N_6228,N_1274,N_713);
xnor U6229 (N_6229,N_4451,N_1094);
nand U6230 (N_6230,N_3494,N_2444);
xor U6231 (N_6231,N_1248,N_2247);
xnor U6232 (N_6232,N_1269,N_4131);
xnor U6233 (N_6233,N_17,N_2593);
xnor U6234 (N_6234,N_2091,N_288);
and U6235 (N_6235,N_1478,N_4026);
and U6236 (N_6236,N_619,N_3963);
and U6237 (N_6237,N_835,N_1829);
and U6238 (N_6238,N_224,N_3465);
nand U6239 (N_6239,N_1624,N_15);
or U6240 (N_6240,N_4109,N_2027);
or U6241 (N_6241,N_1045,N_935);
nor U6242 (N_6242,N_2475,N_3350);
nand U6243 (N_6243,N_2154,N_3394);
xor U6244 (N_6244,N_34,N_3644);
xor U6245 (N_6245,N_1712,N_1813);
nor U6246 (N_6246,N_1121,N_281);
and U6247 (N_6247,N_4718,N_90);
xnor U6248 (N_6248,N_4892,N_1397);
xnor U6249 (N_6249,N_2749,N_1429);
xor U6250 (N_6250,N_2585,N_76);
nor U6251 (N_6251,N_4242,N_2518);
xor U6252 (N_6252,N_2987,N_668);
xnor U6253 (N_6253,N_4601,N_3869);
or U6254 (N_6254,N_3492,N_4599);
nor U6255 (N_6255,N_3736,N_4101);
nand U6256 (N_6256,N_1849,N_356);
xnor U6257 (N_6257,N_933,N_2842);
and U6258 (N_6258,N_2099,N_3252);
nor U6259 (N_6259,N_2569,N_2383);
and U6260 (N_6260,N_2912,N_3219);
or U6261 (N_6261,N_467,N_1479);
nor U6262 (N_6262,N_3229,N_4271);
nor U6263 (N_6263,N_3493,N_2456);
and U6264 (N_6264,N_745,N_2544);
xor U6265 (N_6265,N_135,N_2924);
xor U6266 (N_6266,N_4320,N_4707);
and U6267 (N_6267,N_483,N_763);
nand U6268 (N_6268,N_4918,N_263);
nor U6269 (N_6269,N_4738,N_849);
and U6270 (N_6270,N_316,N_3224);
and U6271 (N_6271,N_4931,N_1859);
nor U6272 (N_6272,N_1367,N_2579);
nand U6273 (N_6273,N_4524,N_1508);
or U6274 (N_6274,N_1840,N_3953);
xnor U6275 (N_6275,N_2450,N_2566);
or U6276 (N_6276,N_4264,N_2369);
and U6277 (N_6277,N_3378,N_4877);
or U6278 (N_6278,N_3327,N_1757);
xnor U6279 (N_6279,N_2102,N_1541);
nand U6280 (N_6280,N_3715,N_689);
nor U6281 (N_6281,N_2567,N_4687);
nor U6282 (N_6282,N_4793,N_1914);
nand U6283 (N_6283,N_4019,N_1422);
nand U6284 (N_6284,N_1821,N_2272);
or U6285 (N_6285,N_2730,N_3700);
or U6286 (N_6286,N_3412,N_4039);
xor U6287 (N_6287,N_739,N_2502);
xor U6288 (N_6288,N_11,N_522);
nor U6289 (N_6289,N_3080,N_972);
and U6290 (N_6290,N_4439,N_2048);
or U6291 (N_6291,N_236,N_1023);
nor U6292 (N_6292,N_4478,N_4751);
xnor U6293 (N_6293,N_3674,N_3874);
or U6294 (N_6294,N_3756,N_1210);
nor U6295 (N_6295,N_3397,N_4540);
nor U6296 (N_6296,N_3368,N_2785);
or U6297 (N_6297,N_534,N_4712);
nand U6298 (N_6298,N_2901,N_3357);
or U6299 (N_6299,N_4397,N_251);
xor U6300 (N_6300,N_3435,N_3764);
or U6301 (N_6301,N_905,N_2254);
nand U6302 (N_6302,N_414,N_1053);
and U6303 (N_6303,N_4395,N_3099);
nand U6304 (N_6304,N_2632,N_28);
nand U6305 (N_6305,N_2793,N_4333);
or U6306 (N_6306,N_3160,N_3134);
nor U6307 (N_6307,N_4893,N_724);
and U6308 (N_6308,N_1768,N_3287);
and U6309 (N_6309,N_4989,N_1243);
or U6310 (N_6310,N_1137,N_2503);
and U6311 (N_6311,N_1565,N_2654);
or U6312 (N_6312,N_2001,N_4362);
xnor U6313 (N_6313,N_2908,N_4496);
and U6314 (N_6314,N_478,N_3163);
nand U6315 (N_6315,N_3480,N_3387);
nand U6316 (N_6316,N_4502,N_186);
xor U6317 (N_6317,N_547,N_4449);
nor U6318 (N_6318,N_3002,N_2936);
nand U6319 (N_6319,N_141,N_4169);
nand U6320 (N_6320,N_963,N_3127);
xor U6321 (N_6321,N_4,N_1980);
nor U6322 (N_6322,N_1951,N_2834);
nor U6323 (N_6323,N_1188,N_3427);
nand U6324 (N_6324,N_4771,N_2235);
nand U6325 (N_6325,N_3270,N_4182);
nor U6326 (N_6326,N_2635,N_169);
nand U6327 (N_6327,N_1346,N_2441);
nor U6328 (N_6328,N_1491,N_1455);
or U6329 (N_6329,N_1614,N_4203);
or U6330 (N_6330,N_3539,N_3384);
or U6331 (N_6331,N_496,N_4357);
nor U6332 (N_6332,N_1975,N_1881);
xnor U6333 (N_6333,N_4904,N_2707);
nand U6334 (N_6334,N_1142,N_3710);
xor U6335 (N_6335,N_1987,N_3285);
xnor U6336 (N_6336,N_3712,N_60);
nor U6337 (N_6337,N_4419,N_1411);
or U6338 (N_6338,N_3139,N_3856);
or U6339 (N_6339,N_2482,N_3663);
and U6340 (N_6340,N_4575,N_716);
and U6341 (N_6341,N_1353,N_1789);
and U6342 (N_6342,N_4290,N_3769);
and U6343 (N_6343,N_1384,N_3680);
nor U6344 (N_6344,N_2485,N_4705);
xor U6345 (N_6345,N_3676,N_4372);
nand U6346 (N_6346,N_1568,N_4088);
nand U6347 (N_6347,N_2042,N_1924);
nor U6348 (N_6348,N_682,N_1955);
nand U6349 (N_6349,N_3460,N_1872);
or U6350 (N_6350,N_260,N_4747);
and U6351 (N_6351,N_1503,N_3361);
or U6352 (N_6352,N_4150,N_323);
nand U6353 (N_6353,N_4122,N_1844);
nor U6354 (N_6354,N_611,N_4727);
and U6355 (N_6355,N_4987,N_352);
nor U6356 (N_6356,N_1189,N_1152);
xor U6357 (N_6357,N_3043,N_1976);
xor U6358 (N_6358,N_2073,N_2331);
nor U6359 (N_6359,N_4180,N_3195);
nor U6360 (N_6360,N_2261,N_4538);
nand U6361 (N_6361,N_4426,N_1038);
nand U6362 (N_6362,N_4508,N_3952);
and U6363 (N_6363,N_910,N_1773);
and U6364 (N_6364,N_4077,N_2545);
nor U6365 (N_6365,N_2620,N_2943);
nor U6366 (N_6366,N_4639,N_588);
nor U6367 (N_6367,N_3300,N_839);
nor U6368 (N_6368,N_3975,N_199);
xnor U6369 (N_6369,N_850,N_2948);
nor U6370 (N_6370,N_1253,N_1966);
nor U6371 (N_6371,N_4448,N_1850);
or U6372 (N_6372,N_2779,N_4468);
xor U6373 (N_6373,N_2549,N_3825);
nor U6374 (N_6374,N_3998,N_3256);
or U6375 (N_6375,N_1227,N_647);
nand U6376 (N_6376,N_112,N_1817);
nand U6377 (N_6377,N_305,N_1463);
and U6378 (N_6378,N_3569,N_2157);
and U6379 (N_6379,N_655,N_2949);
nor U6380 (N_6380,N_3189,N_2341);
xor U6381 (N_6381,N_4843,N_1919);
nor U6382 (N_6382,N_461,N_3306);
nand U6383 (N_6383,N_1168,N_976);
xnor U6384 (N_6384,N_4662,N_4536);
nand U6385 (N_6385,N_3829,N_2049);
nor U6386 (N_6386,N_4886,N_3842);
or U6387 (N_6387,N_2703,N_1513);
nor U6388 (N_6388,N_228,N_3151);
or U6389 (N_6389,N_3884,N_1140);
nor U6390 (N_6390,N_4865,N_523);
or U6391 (N_6391,N_4833,N_2058);
nor U6392 (N_6392,N_2899,N_2638);
nand U6393 (N_6393,N_1459,N_3198);
nand U6394 (N_6394,N_4898,N_2595);
or U6395 (N_6395,N_3798,N_929);
xnor U6396 (N_6396,N_692,N_4255);
and U6397 (N_6397,N_949,N_1383);
nor U6398 (N_6398,N_2408,N_3214);
nand U6399 (N_6399,N_3923,N_690);
xnor U6400 (N_6400,N_314,N_3650);
and U6401 (N_6401,N_3172,N_3552);
nand U6402 (N_6402,N_3690,N_2300);
nand U6403 (N_6403,N_2916,N_394);
or U6404 (N_6404,N_132,N_1089);
or U6405 (N_6405,N_1417,N_4261);
and U6406 (N_6406,N_2072,N_3575);
nor U6407 (N_6407,N_4933,N_776);
nand U6408 (N_6408,N_4248,N_1194);
nand U6409 (N_6409,N_4469,N_867);
and U6410 (N_6410,N_4484,N_1284);
nor U6411 (N_6411,N_1252,N_4815);
nand U6412 (N_6412,N_4675,N_426);
nand U6413 (N_6413,N_1547,N_2599);
nor U6414 (N_6414,N_324,N_328);
xor U6415 (N_6415,N_2511,N_3021);
nand U6416 (N_6416,N_2657,N_2342);
or U6417 (N_6417,N_3221,N_4529);
xor U6418 (N_6418,N_3328,N_4352);
and U6419 (N_6419,N_2176,N_2025);
xnor U6420 (N_6420,N_1107,N_1983);
and U6421 (N_6421,N_2897,N_3677);
xnor U6422 (N_6422,N_3607,N_4699);
nor U6423 (N_6423,N_694,N_4217);
nand U6424 (N_6424,N_29,N_4317);
and U6425 (N_6425,N_78,N_2822);
nor U6426 (N_6426,N_2101,N_3621);
xor U6427 (N_6427,N_2847,N_743);
xor U6428 (N_6428,N_3108,N_3075);
xor U6429 (N_6429,N_3848,N_2366);
and U6430 (N_6430,N_4998,N_605);
nor U6431 (N_6431,N_4083,N_4060);
xnor U6432 (N_6432,N_3345,N_1886);
xor U6433 (N_6433,N_3225,N_4906);
nand U6434 (N_6434,N_3870,N_2688);
nand U6435 (N_6435,N_2978,N_1713);
xor U6436 (N_6436,N_1394,N_2574);
or U6437 (N_6437,N_3956,N_1258);
nor U6438 (N_6438,N_2740,N_3119);
nor U6439 (N_6439,N_1511,N_632);
and U6440 (N_6440,N_1634,N_574);
nor U6441 (N_6441,N_1674,N_3741);
nor U6442 (N_6442,N_1785,N_2721);
or U6443 (N_6443,N_1167,N_277);
or U6444 (N_6444,N_4794,N_4489);
or U6445 (N_6445,N_1556,N_1357);
nand U6446 (N_6446,N_814,N_2640);
xnor U6447 (N_6447,N_1179,N_3087);
nor U6448 (N_6448,N_3509,N_4808);
and U6449 (N_6449,N_2376,N_3675);
xor U6450 (N_6450,N_274,N_2806);
xnor U6451 (N_6451,N_331,N_1637);
or U6452 (N_6452,N_636,N_2762);
xor U6453 (N_6453,N_1801,N_1126);
or U6454 (N_6454,N_1340,N_142);
xor U6455 (N_6455,N_269,N_4844);
and U6456 (N_6456,N_1395,N_3624);
or U6457 (N_6457,N_4923,N_4676);
xnor U6458 (N_6458,N_707,N_2248);
and U6459 (N_6459,N_529,N_4396);
xor U6460 (N_6460,N_3777,N_3999);
and U6461 (N_6461,N_4315,N_4531);
nand U6462 (N_6462,N_1105,N_1909);
nor U6463 (N_6463,N_1,N_1290);
xor U6464 (N_6464,N_213,N_307);
or U6465 (N_6465,N_1663,N_4102);
xnor U6466 (N_6466,N_2149,N_2270);
and U6467 (N_6467,N_3586,N_4466);
nor U6468 (N_6468,N_428,N_1567);
nand U6469 (N_6469,N_4985,N_1321);
nand U6470 (N_6470,N_3154,N_10);
nand U6471 (N_6471,N_2069,N_734);
xor U6472 (N_6472,N_1607,N_1283);
or U6473 (N_6473,N_1943,N_3612);
and U6474 (N_6474,N_1251,N_2047);
or U6475 (N_6475,N_3169,N_3299);
or U6476 (N_6476,N_1470,N_507);
xor U6477 (N_6477,N_4082,N_4632);
or U6478 (N_6478,N_2679,N_3051);
nor U6479 (N_6479,N_996,N_1927);
xnor U6480 (N_6480,N_4220,N_1780);
xnor U6481 (N_6481,N_216,N_639);
or U6482 (N_6482,N_3747,N_1083);
and U6483 (N_6483,N_3852,N_2964);
nand U6484 (N_6484,N_1990,N_1680);
and U6485 (N_6485,N_446,N_4557);
xor U6486 (N_6486,N_2498,N_2354);
xnor U6487 (N_6487,N_2007,N_1534);
xor U6488 (N_6488,N_66,N_2222);
nand U6489 (N_6489,N_3403,N_2465);
nor U6490 (N_6490,N_691,N_2387);
xnor U6491 (N_6491,N_868,N_33);
or U6492 (N_6492,N_2057,N_3253);
nand U6493 (N_6493,N_2022,N_2689);
xnor U6494 (N_6494,N_3197,N_3330);
and U6495 (N_6495,N_578,N_1703);
nor U6496 (N_6496,N_2338,N_2141);
or U6497 (N_6497,N_2314,N_212);
or U6498 (N_6498,N_3067,N_4679);
xor U6499 (N_6499,N_4832,N_3722);
or U6500 (N_6500,N_253,N_194);
or U6501 (N_6501,N_2402,N_4876);
nand U6502 (N_6502,N_2754,N_477);
xor U6503 (N_6503,N_4521,N_3946);
nand U6504 (N_6504,N_4651,N_1802);
xnor U6505 (N_6505,N_3033,N_1726);
nand U6506 (N_6506,N_3797,N_2315);
xor U6507 (N_6507,N_1225,N_1737);
nand U6508 (N_6508,N_344,N_4674);
xor U6509 (N_6509,N_742,N_3599);
and U6510 (N_6510,N_941,N_3605);
nand U6511 (N_6511,N_1686,N_3571);
nand U6512 (N_6512,N_4190,N_396);
and U6513 (N_6513,N_3903,N_3899);
nor U6514 (N_6514,N_4161,N_3104);
nand U6515 (N_6515,N_940,N_1166);
nand U6516 (N_6516,N_418,N_4493);
nor U6517 (N_6517,N_3788,N_2152);
and U6518 (N_6518,N_922,N_805);
xnor U6519 (N_6519,N_317,N_333);
nand U6520 (N_6520,N_3158,N_1692);
xnor U6521 (N_6521,N_2484,N_4165);
or U6522 (N_6522,N_1147,N_4603);
and U6523 (N_6523,N_4241,N_2043);
xnor U6524 (N_6524,N_3477,N_1482);
or U6525 (N_6525,N_1504,N_1439);
and U6526 (N_6526,N_1287,N_4784);
or U6527 (N_6527,N_3281,N_18);
and U6528 (N_6528,N_1347,N_4587);
nand U6529 (N_6529,N_2892,N_4836);
or U6530 (N_6530,N_3284,N_4896);
or U6531 (N_6531,N_2490,N_4028);
nand U6532 (N_6532,N_1090,N_4552);
nand U6533 (N_6533,N_3868,N_2068);
xor U6534 (N_6534,N_3524,N_1317);
xor U6535 (N_6535,N_311,N_3895);
nand U6536 (N_6536,N_1792,N_1077);
or U6537 (N_6537,N_1830,N_2727);
nand U6538 (N_6538,N_2590,N_3392);
nand U6539 (N_6539,N_722,N_1039);
xnor U6540 (N_6540,N_4964,N_1017);
and U6541 (N_6541,N_527,N_2766);
xor U6542 (N_6542,N_2190,N_596);
nor U6543 (N_6543,N_2670,N_2452);
or U6544 (N_6544,N_2607,N_2096);
nor U6545 (N_6545,N_4556,N_4754);
and U6546 (N_6546,N_4185,N_3554);
and U6547 (N_6547,N_2374,N_2746);
xor U6548 (N_6548,N_1309,N_4974);
xnor U6549 (N_6549,N_4128,N_684);
nor U6550 (N_6550,N_383,N_155);
xnor U6551 (N_6551,N_4620,N_3790);
and U6552 (N_6552,N_3896,N_3526);
nand U6553 (N_6553,N_1906,N_4855);
nand U6554 (N_6554,N_1096,N_3210);
nor U6555 (N_6555,N_2148,N_650);
nand U6556 (N_6556,N_614,N_1390);
or U6557 (N_6557,N_2555,N_75);
xnor U6558 (N_6558,N_35,N_2083);
and U6559 (N_6559,N_153,N_1414);
nand U6560 (N_6560,N_2819,N_4120);
nand U6561 (N_6561,N_1512,N_1848);
or U6562 (N_6562,N_4961,N_4149);
or U6563 (N_6563,N_3761,N_280);
or U6564 (N_6564,N_2346,N_106);
xnor U6565 (N_6565,N_3750,N_3582);
or U6566 (N_6566,N_3377,N_2952);
xor U6567 (N_6567,N_735,N_3138);
nand U6568 (N_6568,N_4852,N_439);
nor U6569 (N_6569,N_3986,N_1474);
and U6570 (N_6570,N_1010,N_757);
xnor U6571 (N_6571,N_3698,N_880);
nand U6572 (N_6572,N_44,N_137);
nor U6573 (N_6573,N_3422,N_4592);
nor U6574 (N_6574,N_1510,N_846);
and U6575 (N_6575,N_4363,N_4922);
or U6576 (N_6576,N_897,N_918);
nor U6577 (N_6577,N_4905,N_2505);
nor U6578 (N_6578,N_3501,N_73);
or U6579 (N_6579,N_4193,N_4472);
and U6580 (N_6580,N_3029,N_3565);
or U6581 (N_6581,N_3102,N_3646);
nor U6582 (N_6582,N_4250,N_4103);
nand U6583 (N_6583,N_3318,N_2542);
and U6584 (N_6584,N_2350,N_2211);
nor U6585 (N_6585,N_3273,N_1589);
and U6586 (N_6586,N_2641,N_457);
nand U6587 (N_6587,N_451,N_906);
xor U6588 (N_6588,N_4667,N_1097);
and U6589 (N_6589,N_1884,N_2876);
nor U6590 (N_6590,N_688,N_3584);
nor U6591 (N_6591,N_1861,N_4814);
nand U6592 (N_6592,N_7,N_422);
xor U6593 (N_6593,N_634,N_2683);
nand U6594 (N_6594,N_3502,N_487);
and U6595 (N_6595,N_1667,N_2706);
nor U6596 (N_6596,N_4953,N_736);
or U6597 (N_6597,N_971,N_3383);
and U6598 (N_6598,N_3495,N_3199);
xnor U6599 (N_6599,N_3238,N_2263);
nor U6600 (N_6600,N_4802,N_2435);
or U6601 (N_6601,N_152,N_581);
nand U6602 (N_6602,N_3196,N_1647);
nand U6603 (N_6603,N_3553,N_1259);
nor U6604 (N_6604,N_149,N_1223);
xnor U6605 (N_6605,N_168,N_3634);
or U6606 (N_6606,N_4257,N_406);
nand U6607 (N_6607,N_1736,N_4837);
nand U6608 (N_6608,N_4339,N_2552);
nor U6609 (N_6609,N_3532,N_2079);
nor U6610 (N_6610,N_1968,N_3639);
xor U6611 (N_6611,N_3853,N_2202);
and U6612 (N_6612,N_2994,N_255);
xor U6613 (N_6613,N_1141,N_2184);
nand U6614 (N_6614,N_1685,N_4746);
nand U6615 (N_6615,N_3844,N_2841);
or U6616 (N_6616,N_2510,N_3811);
nor U6617 (N_6617,N_466,N_2774);
and U6618 (N_6618,N_2092,N_2215);
nor U6619 (N_6619,N_859,N_714);
xnor U6620 (N_6620,N_3907,N_1735);
nand U6621 (N_6621,N_2100,N_2421);
nand U6622 (N_6622,N_2856,N_4756);
or U6623 (N_6623,N_4047,N_4089);
or U6624 (N_6624,N_2598,N_4329);
xnor U6625 (N_6625,N_2026,N_4504);
and U6626 (N_6626,N_4527,N_4874);
xor U6627 (N_6627,N_1279,N_3271);
nor U6628 (N_6628,N_4488,N_4883);
nor U6629 (N_6629,N_2764,N_4401);
xnor U6630 (N_6630,N_234,N_2071);
or U6631 (N_6631,N_1537,N_2127);
nor U6632 (N_6632,N_1705,N_2504);
nor U6633 (N_6633,N_4054,N_3439);
or U6634 (N_6634,N_543,N_3640);
nand U6635 (N_6635,N_1036,N_1331);
or U6636 (N_6636,N_884,N_4755);
xor U6637 (N_6637,N_1380,N_20);
and U6638 (N_6638,N_2478,N_2330);
or U6639 (N_6639,N_1699,N_1148);
and U6640 (N_6640,N_2904,N_1319);
or U6641 (N_6641,N_3452,N_4223);
nand U6642 (N_6642,N_4530,N_3232);
nor U6643 (N_6643,N_4009,N_2399);
nor U6644 (N_6644,N_4834,N_1716);
and U6645 (N_6645,N_156,N_2848);
xor U6646 (N_6646,N_1668,N_14);
nand U6647 (N_6647,N_2151,N_3916);
and U6648 (N_6648,N_3694,N_4681);
xnor U6649 (N_6649,N_475,N_4011);
nand U6650 (N_6650,N_2515,N_3359);
nand U6651 (N_6651,N_3342,N_3165);
xor U6652 (N_6652,N_1743,N_3925);
and U6653 (N_6653,N_2572,N_326);
nor U6654 (N_6654,N_2556,N_4517);
or U6655 (N_6655,N_1443,N_542);
nor U6656 (N_6656,N_1845,N_3734);
or U6657 (N_6657,N_3721,N_4741);
or U6658 (N_6658,N_4299,N_1842);
xor U6659 (N_6659,N_1495,N_888);
nor U6660 (N_6660,N_883,N_1623);
xor U6661 (N_6661,N_4672,N_1181);
xor U6662 (N_6662,N_136,N_3430);
nand U6663 (N_6663,N_3453,N_1431);
or U6664 (N_6664,N_1234,N_1327);
nor U6665 (N_6665,N_1406,N_2120);
nor U6666 (N_6666,N_4391,N_2293);
and U6667 (N_6667,N_1546,N_3116);
nand U6668 (N_6668,N_2420,N_3635);
and U6669 (N_6669,N_3263,N_2831);
or U6670 (N_6670,N_27,N_4926);
and U6671 (N_6671,N_3534,N_3293);
nand U6672 (N_6672,N_409,N_1341);
xor U6673 (N_6673,N_869,N_3996);
xor U6674 (N_6674,N_3751,N_3742);
and U6675 (N_6675,N_1620,N_2362);
xnor U6676 (N_6676,N_4316,N_2540);
nor U6677 (N_6677,N_2137,N_1751);
nand U6678 (N_6678,N_1532,N_2440);
nor U6679 (N_6679,N_4078,N_1806);
nor U6680 (N_6680,N_4256,N_985);
xor U6681 (N_6681,N_3335,N_1149);
nand U6682 (N_6682,N_1745,N_4990);
or U6683 (N_6683,N_389,N_3778);
or U6684 (N_6684,N_3118,N_1805);
and U6685 (N_6685,N_753,N_2583);
nand U6686 (N_6686,N_1339,N_3049);
nor U6687 (N_6687,N_3802,N_3401);
nand U6688 (N_6688,N_2087,N_1307);
nand U6689 (N_6689,N_2464,N_2745);
xnor U6690 (N_6690,N_87,N_1012);
and U6691 (N_6691,N_1648,N_2094);
and U6692 (N_6692,N_2944,N_3007);
and U6693 (N_6693,N_61,N_4013);
nor U6694 (N_6694,N_1585,N_2606);
nor U6695 (N_6695,N_3714,N_1218);
or U6696 (N_6696,N_4568,N_2229);
nand U6697 (N_6697,N_677,N_914);
nand U6698 (N_6698,N_4857,N_1305);
xor U6699 (N_6699,N_102,N_1379);
nand U6700 (N_6700,N_4525,N_943);
and U6701 (N_6701,N_270,N_2391);
nand U6702 (N_6702,N_890,N_1076);
nand U6703 (N_6703,N_4302,N_645);
and U6704 (N_6704,N_1575,N_1122);
xnor U6705 (N_6705,N_4750,N_4863);
nor U6706 (N_6706,N_3954,N_4658);
xor U6707 (N_6707,N_207,N_1521);
nor U6708 (N_6708,N_1747,N_2245);
nor U6709 (N_6709,N_1268,N_3723);
or U6710 (N_6710,N_2140,N_2701);
or U6711 (N_6711,N_283,N_3772);
nand U6712 (N_6712,N_3888,N_1425);
nor U6713 (N_6713,N_4643,N_2956);
nand U6714 (N_6714,N_3536,N_772);
xnor U6715 (N_6715,N_3866,N_3589);
or U6716 (N_6716,N_3207,N_2497);
nand U6717 (N_6717,N_4976,N_4016);
or U6718 (N_6718,N_820,N_1398);
nand U6719 (N_6719,N_3603,N_4623);
nand U6720 (N_6720,N_151,N_558);
or U6721 (N_6721,N_1530,N_3519);
nor U6722 (N_6722,N_1492,N_2850);
nand U6723 (N_6723,N_2085,N_1679);
and U6724 (N_6724,N_2116,N_857);
nand U6725 (N_6725,N_1783,N_3254);
nand U6726 (N_6726,N_1843,N_2431);
xnor U6727 (N_6727,N_421,N_3283);
nor U6728 (N_6728,N_959,N_513);
nor U6729 (N_6729,N_609,N_3758);
nor U6730 (N_6730,N_3912,N_807);
xnor U6731 (N_6731,N_3601,N_3667);
nor U6732 (N_6732,N_671,N_2861);
nand U6733 (N_6733,N_404,N_1996);
xnor U6734 (N_6734,N_3754,N_4110);
xnor U6735 (N_6735,N_3078,N_1683);
nand U6736 (N_6736,N_2045,N_3875);
or U6737 (N_6737,N_1467,N_1864);
and U6738 (N_6738,N_3277,N_4692);
xor U6739 (N_6739,N_3517,N_3514);
and U6740 (N_6740,N_1070,N_3405);
and U6741 (N_6741,N_956,N_2589);
nand U6742 (N_6742,N_1659,N_2281);
nor U6743 (N_6743,N_960,N_3669);
nor U6744 (N_6744,N_4324,N_4657);
nor U6745 (N_6745,N_3725,N_4826);
and U6746 (N_6746,N_3559,N_1578);
and U6747 (N_6747,N_786,N_4388);
nor U6748 (N_6748,N_519,N_2443);
xnor U6749 (N_6749,N_3941,N_3242);
nand U6750 (N_6750,N_2546,N_2833);
or U6751 (N_6751,N_3611,N_3763);
and U6752 (N_6752,N_2138,N_2126);
nand U6753 (N_6753,N_3835,N_4313);
nor U6754 (N_6754,N_367,N_419);
xnor U6755 (N_6755,N_2382,N_4604);
nor U6756 (N_6756,N_4099,N_1326);
and U6757 (N_6757,N_3508,N_1769);
xnor U6758 (N_6758,N_2053,N_4722);
nand U6759 (N_6759,N_1895,N_2608);
xnor U6760 (N_6760,N_3347,N_3965);
and U6761 (N_6761,N_2446,N_2432);
and U6762 (N_6762,N_4622,N_3783);
or U6763 (N_6763,N_1006,N_924);
nand U6764 (N_6764,N_3045,N_559);
nand U6765 (N_6765,N_2788,N_876);
nand U6766 (N_6766,N_3482,N_4067);
and U6767 (N_6767,N_658,N_3528);
or U6768 (N_6768,N_2323,N_4259);
and U6769 (N_6769,N_4273,N_4656);
and U6770 (N_6770,N_1856,N_3008);
or U6771 (N_6771,N_3081,N_1498);
nand U6772 (N_6772,N_2536,N_3454);
xor U6773 (N_6773,N_267,N_2921);
nand U6774 (N_6774,N_794,N_672);
xnor U6775 (N_6775,N_415,N_3890);
nor U6776 (N_6776,N_3086,N_2983);
nor U6777 (N_6777,N_4454,N_1642);
or U6778 (N_6778,N_3876,N_4221);
nand U6779 (N_6779,N_1368,N_3056);
and U6780 (N_6780,N_1619,N_1208);
nor U6781 (N_6781,N_649,N_2775);
or U6782 (N_6782,N_3513,N_1232);
or U6783 (N_6783,N_4759,N_4491);
and U6784 (N_6784,N_1950,N_3244);
and U6785 (N_6785,N_2917,N_3421);
xor U6786 (N_6786,N_4343,N_3703);
xnor U6787 (N_6787,N_3479,N_2326);
and U6788 (N_6788,N_816,N_3628);
or U6789 (N_6789,N_858,N_4715);
nand U6790 (N_6790,N_1942,N_4912);
or U6791 (N_6791,N_939,N_4800);
xor U6792 (N_6792,N_1548,N_453);
or U6793 (N_6793,N_1496,N_3466);
xnor U6794 (N_6794,N_2461,N_1754);
or U6795 (N_6795,N_3566,N_3035);
xnor U6796 (N_6796,N_818,N_1646);
and U6797 (N_6797,N_2816,N_2523);
and U6798 (N_6798,N_2930,N_3838);
or U6799 (N_6799,N_1361,N_239);
nand U6800 (N_6800,N_2201,N_1718);
and U6801 (N_6801,N_586,N_360);
and U6802 (N_6802,N_4458,N_646);
and U6803 (N_6803,N_2067,N_4698);
and U6804 (N_6804,N_2697,N_3182);
nand U6805 (N_6805,N_1561,N_537);
nand U6806 (N_6806,N_2289,N_165);
or U6807 (N_6807,N_1193,N_2294);
or U6808 (N_6808,N_2702,N_101);
and U6809 (N_6809,N_2909,N_4167);
nor U6810 (N_6810,N_1065,N_82);
or U6811 (N_6811,N_871,N_3098);
or U6812 (N_6812,N_2012,N_2902);
xor U6813 (N_6813,N_3450,N_157);
nor U6814 (N_6814,N_3683,N_3380);
or U6815 (N_6815,N_2710,N_2857);
or U6816 (N_6816,N_3682,N_900);
or U6817 (N_6817,N_2880,N_1029);
nor U6818 (N_6818,N_2600,N_233);
nand U6819 (N_6819,N_113,N_4046);
and U6820 (N_6820,N_2653,N_3205);
and U6821 (N_6821,N_3942,N_4093);
and U6822 (N_6822,N_817,N_593);
nor U6823 (N_6823,N_2723,N_728);
xnor U6824 (N_6824,N_286,N_30);
and U6825 (N_6825,N_2213,N_983);
or U6826 (N_6826,N_723,N_665);
and U6827 (N_6827,N_2016,N_4901);
xnor U6828 (N_6828,N_4284,N_3175);
and U6829 (N_6829,N_4847,N_1582);
and U6830 (N_6830,N_1085,N_4318);
nand U6831 (N_6831,N_3567,N_1191);
xnor U6832 (N_6832,N_4200,N_162);
and U6833 (N_6833,N_2470,N_1264);
and U6834 (N_6834,N_4050,N_3652);
and U6835 (N_6835,N_861,N_3547);
xnor U6836 (N_6836,N_4049,N_2838);
nor U6837 (N_6837,N_2787,N_4085);
nand U6838 (N_6838,N_899,N_3260);
nor U6839 (N_6839,N_3018,N_2442);
or U6840 (N_6840,N_967,N_1207);
nor U6841 (N_6841,N_2165,N_4227);
xnor U6842 (N_6842,N_4262,N_1651);
xnor U6843 (N_6843,N_3609,N_4541);
nor U6844 (N_6844,N_1366,N_4749);
or U6845 (N_6845,N_4114,N_3623);
and U6846 (N_6846,N_563,N_3428);
or U6847 (N_6847,N_4895,N_4305);
and U6848 (N_6848,N_3749,N_1701);
nor U6849 (N_6849,N_4688,N_3373);
and U6850 (N_6850,N_53,N_2084);
nor U6851 (N_6851,N_3404,N_1020);
nor U6852 (N_6852,N_2659,N_1231);
xnor U6853 (N_6853,N_633,N_3473);
or U6854 (N_6854,N_1777,N_3145);
nor U6855 (N_6855,N_284,N_370);
nor U6856 (N_6856,N_2332,N_4045);
nand U6857 (N_6857,N_2098,N_295);
nand U6858 (N_6858,N_1484,N_1874);
nor U6859 (N_6859,N_2830,N_1456);
nand U6860 (N_6860,N_719,N_2164);
nor U6861 (N_6861,N_4416,N_2115);
and U6862 (N_6862,N_2911,N_2050);
xnor U6863 (N_6863,N_4752,N_3726);
nor U6864 (N_6864,N_4761,N_3148);
and U6865 (N_6865,N_1520,N_2577);
xor U6866 (N_6866,N_3026,N_3470);
nor U6867 (N_6867,N_1405,N_1594);
nand U6868 (N_6868,N_190,N_2207);
nand U6869 (N_6869,N_4875,N_189);
nand U6870 (N_6870,N_4579,N_3351);
or U6871 (N_6871,N_88,N_115);
nor U6872 (N_6872,N_240,N_1694);
and U6873 (N_6873,N_1299,N_524);
and U6874 (N_6874,N_4125,N_160);
xnor U6875 (N_6875,N_3617,N_1169);
and U6876 (N_6876,N_4840,N_4841);
nor U6877 (N_6877,N_872,N_1910);
or U6878 (N_6878,N_1676,N_1891);
nor U6879 (N_6879,N_2014,N_3251);
and U6880 (N_6880,N_3529,N_4415);
and U6881 (N_6881,N_4680,N_2146);
xor U6882 (N_6882,N_1452,N_252);
xor U6883 (N_6883,N_4939,N_371);
xor U6884 (N_6884,N_4798,N_831);
xnor U6885 (N_6885,N_2124,N_1249);
and U6886 (N_6886,N_4370,N_4829);
and U6887 (N_6887,N_4170,N_3082);
nor U6888 (N_6888,N_353,N_272);
or U6889 (N_6889,N_1562,N_769);
or U6890 (N_6890,N_793,N_4456);
nand U6891 (N_6891,N_3521,N_2872);
or U6892 (N_6892,N_3250,N_2368);
nor U6893 (N_6893,N_3413,N_783);
and U6894 (N_6894,N_2851,N_1862);
and U6895 (N_6895,N_1501,N_4286);
or U6896 (N_6896,N_1597,N_2695);
or U6897 (N_6897,N_3673,N_1003);
and U6898 (N_6898,N_217,N_3913);
nand U6899 (N_6899,N_1923,N_4669);
nor U6900 (N_6900,N_1206,N_4499);
and U6901 (N_6901,N_1952,N_2418);
nand U6902 (N_6902,N_1509,N_1525);
nor U6903 (N_6903,N_4548,N_2868);
xnor U6904 (N_6904,N_3068,N_2669);
nor U6905 (N_6905,N_413,N_1257);
and U6906 (N_6906,N_951,N_79);
or U6907 (N_6907,N_2125,N_2810);
and U6908 (N_6908,N_1413,N_4889);
xor U6909 (N_6909,N_4052,N_222);
xnor U6910 (N_6910,N_2002,N_4424);
xor U6911 (N_6911,N_2239,N_1302);
and U6912 (N_6912,N_4409,N_3520);
or U6913 (N_6913,N_1698,N_4522);
or U6914 (N_6914,N_1043,N_642);
and U6915 (N_6915,N_2668,N_2226);
or U6916 (N_6916,N_4156,N_1905);
nand U6917 (N_6917,N_257,N_1118);
and U6918 (N_6918,N_1894,N_540);
nor U6919 (N_6919,N_931,N_4432);
and U6920 (N_6920,N_4740,N_1616);
xor U6921 (N_6921,N_2508,N_2244);
or U6922 (N_6922,N_3354,N_4997);
xor U6923 (N_6923,N_3819,N_1867);
nand U6924 (N_6924,N_2672,N_4817);
nor U6925 (N_6925,N_3845,N_1062);
and U6926 (N_6926,N_1382,N_1823);
or U6927 (N_6927,N_2439,N_3827);
nand U6928 (N_6928,N_1673,N_3415);
nand U6929 (N_6929,N_4482,N_1018);
xnor U6930 (N_6930,N_3150,N_4147);
nor U6931 (N_6931,N_3596,N_2784);
or U6932 (N_6932,N_2412,N_1136);
nor U6933 (N_6933,N_1336,N_1846);
nand U6934 (N_6934,N_3215,N_2494);
xnor U6935 (N_6935,N_3391,N_209);
nand U6936 (N_6936,N_4381,N_666);
xor U6937 (N_6937,N_1518,N_197);
nand U6938 (N_6938,N_4266,N_3909);
or U6939 (N_6939,N_1993,N_4422);
and U6940 (N_6940,N_4890,N_432);
nor U6941 (N_6941,N_2467,N_1544);
nor U6942 (N_6942,N_721,N_1608);
or U6943 (N_6943,N_4644,N_2519);
and U6944 (N_6944,N_4971,N_508);
xor U6945 (N_6945,N_1123,N_480);
and U6946 (N_6946,N_2023,N_1150);
nand U6947 (N_6947,N_1766,N_2761);
or U6948 (N_6948,N_2995,N_4613);
nor U6949 (N_6949,N_847,N_96);
nand U6950 (N_6950,N_601,N_1214);
nor U6951 (N_6951,N_992,N_4279);
nor U6952 (N_6952,N_12,N_1064);
and U6953 (N_6953,N_1781,N_4369);
xnor U6954 (N_6954,N_4950,N_2169);
nand U6955 (N_6955,N_2855,N_3752);
and U6956 (N_6956,N_4111,N_211);
xor U6957 (N_6957,N_2889,N_4511);
nand U6958 (N_6958,N_1876,N_2828);
or U6959 (N_6959,N_1863,N_4390);
nor U6960 (N_6960,N_4137,N_841);
nand U6961 (N_6961,N_215,N_1593);
nor U6962 (N_6962,N_347,N_4480);
and U6963 (N_6963,N_4486,N_4959);
nor U6964 (N_6964,N_2895,N_1356);
nor U6965 (N_6965,N_4554,N_3132);
xnor U6966 (N_6966,N_3985,N_4196);
nand U6967 (N_6967,N_3192,N_4641);
xor U6968 (N_6968,N_730,N_3836);
and U6969 (N_6969,N_2114,N_3961);
xor U6970 (N_6970,N_1124,N_1013);
and U6971 (N_6971,N_1986,N_2181);
and U6972 (N_6972,N_2885,N_1462);
or U6973 (N_6973,N_9,N_376);
nand U6974 (N_6974,N_2133,N_1084);
or U6975 (N_6975,N_407,N_51);
nand U6976 (N_6976,N_4311,N_1033);
xnor U6977 (N_6977,N_3149,N_2206);
or U6978 (N_6978,N_4081,N_4062);
xnor U6979 (N_6979,N_4642,N_1599);
nand U6980 (N_6980,N_3135,N_1330);
xnor U6981 (N_6981,N_3538,N_4921);
nor U6982 (N_6982,N_4490,N_4803);
nor U6983 (N_6983,N_4392,N_4807);
and U6984 (N_6984,N_4994,N_974);
nor U6985 (N_6985,N_781,N_3441);
and U6986 (N_6986,N_667,N_3456);
and U6987 (N_6987,N_3276,N_712);
xnor U6988 (N_6988,N_1292,N_148);
xnor U6989 (N_6989,N_3309,N_4341);
or U6990 (N_6990,N_4992,N_1740);
or U6991 (N_6991,N_4194,N_2426);
nand U6992 (N_6992,N_531,N_2011);
or U6993 (N_6993,N_3130,N_4983);
or U6994 (N_6994,N_4072,N_420);
nand U6995 (N_6995,N_4327,N_4510);
nor U6996 (N_6996,N_679,N_3462);
xor U6997 (N_6997,N_3343,N_4332);
nand U6998 (N_6998,N_4312,N_1997);
xnor U6999 (N_6999,N_254,N_1981);
nor U7000 (N_7000,N_4816,N_2643);
xor U7001 (N_7001,N_2812,N_4949);
nor U7002 (N_7002,N_4403,N_223);
nor U7003 (N_7003,N_3739,N_3931);
nand U7004 (N_7004,N_4634,N_3672);
xor U7005 (N_7005,N_1557,N_4059);
nand U7006 (N_7006,N_231,N_504);
nand U7007 (N_7007,N_1267,N_937);
xor U7008 (N_7008,N_427,N_3278);
or U7009 (N_7009,N_1598,N_4879);
nor U7010 (N_7010,N_86,N_1814);
and U7011 (N_7011,N_4417,N_4238);
and U7012 (N_7012,N_47,N_3085);
xnor U7013 (N_7013,N_2584,N_3822);
xnor U7014 (N_7014,N_327,N_3787);
nand U7015 (N_7015,N_2296,N_1786);
nor U7016 (N_7016,N_4091,N_2197);
and U7017 (N_7017,N_1054,N_3047);
nand U7018 (N_7018,N_294,N_685);
and U7019 (N_7019,N_3393,N_2252);
or U7020 (N_7020,N_3958,N_1882);
nand U7021 (N_7021,N_4653,N_2946);
and U7022 (N_7022,N_968,N_3600);
nor U7023 (N_7023,N_3302,N_320);
nor U7024 (N_7024,N_2631,N_1461);
nor U7025 (N_7025,N_1374,N_731);
and U7026 (N_7026,N_4322,N_1953);
nand U7027 (N_7027,N_2107,N_741);
nand U7028 (N_7028,N_3800,N_4331);
nand U7029 (N_7029,N_1725,N_3915);
nor U7030 (N_7030,N_2405,N_2406);
xnor U7031 (N_7031,N_3004,N_904);
and U7032 (N_7032,N_2156,N_456);
nor U7033 (N_7033,N_2858,N_762);
or U7034 (N_7034,N_1487,N_2685);
nor U7035 (N_7035,N_3094,N_1610);
nor U7036 (N_7036,N_4035,N_1772);
or U7037 (N_7037,N_4567,N_3329);
and U7038 (N_7038,N_2967,N_570);
and U7039 (N_7039,N_4702,N_2290);
nand U7040 (N_7040,N_4301,N_2078);
and U7041 (N_7041,N_2720,N_501);
xor U7042 (N_7042,N_4174,N_1970);
xnor U7043 (N_7043,N_2963,N_3557);
nand U7044 (N_7044,N_2384,N_4869);
and U7045 (N_7045,N_3814,N_3019);
or U7046 (N_7046,N_2130,N_510);
and U7047 (N_7047,N_903,N_1434);
xnor U7048 (N_7048,N_4891,N_3023);
xor U7049 (N_7049,N_2865,N_4181);
xnor U7050 (N_7050,N_4483,N_3363);
nand U7051 (N_7051,N_4159,N_127);
or U7052 (N_7052,N_2728,N_2240);
nor U7053 (N_7053,N_1371,N_110);
xor U7054 (N_7054,N_3658,N_2217);
and U7055 (N_7055,N_1093,N_606);
and U7056 (N_7056,N_727,N_2335);
and U7057 (N_7057,N_1190,N_620);
nand U7058 (N_7058,N_856,N_629);
nor U7059 (N_7059,N_358,N_535);
nor U7060 (N_7060,N_1392,N_2492);
xnor U7061 (N_7061,N_4139,N_2984);
nor U7062 (N_7062,N_4804,N_4003);
nor U7063 (N_7063,N_4345,N_3389);
nor U7064 (N_7064,N_1135,N_907);
xor U7065 (N_7065,N_2413,N_4809);
xor U7066 (N_7066,N_2483,N_2616);
nor U7067 (N_7067,N_1935,N_2681);
nor U7068 (N_7068,N_1471,N_2266);
xnor U7069 (N_7069,N_1095,N_2926);
xor U7070 (N_7070,N_4973,N_1475);
nor U7071 (N_7071,N_4960,N_681);
and U7072 (N_7072,N_3209,N_2436);
xnor U7073 (N_7073,N_2539,N_1756);
and U7074 (N_7074,N_751,N_4872);
and U7075 (N_7075,N_2604,N_3020);
xor U7076 (N_7076,N_3563,N_297);
nor U7077 (N_7077,N_2028,N_1880);
nand U7078 (N_7078,N_3292,N_455);
and U7079 (N_7079,N_3865,N_3265);
nand U7080 (N_7080,N_695,N_3408);
and U7081 (N_7081,N_2158,N_4986);
xor U7082 (N_7082,N_3114,N_366);
and U7083 (N_7083,N_4555,N_3729);
nand U7084 (N_7084,N_705,N_2000);
nor U7085 (N_7085,N_3417,N_1250);
or U7086 (N_7086,N_1354,N_2195);
and U7087 (N_7087,N_2611,N_74);
nand U7088 (N_7088,N_3791,N_4866);
nor U7089 (N_7089,N_4437,N_4621);
or U7090 (N_7090,N_2605,N_2065);
or U7091 (N_7091,N_2403,N_2044);
xor U7092 (N_7092,N_4944,N_278);
nor U7093 (N_7093,N_2798,N_3851);
or U7094 (N_7094,N_521,N_564);
nand U7095 (N_7095,N_3720,N_3120);
or U7096 (N_7096,N_3141,N_982);
or U7097 (N_7097,N_4664,N_607);
xnor U7098 (N_7098,N_3815,N_2580);
nor U7099 (N_7099,N_2168,N_219);
or U7100 (N_7100,N_3733,N_4265);
xnor U7101 (N_7101,N_3459,N_1275);
or U7102 (N_7102,N_1262,N_180);
or U7103 (N_7103,N_4442,N_2708);
and U7104 (N_7104,N_158,N_56);
xor U7105 (N_7105,N_3499,N_1037);
nor U7106 (N_7106,N_912,N_4772);
nor U7107 (N_7107,N_4306,N_3352);
xnor U7108 (N_7108,N_340,N_2040);
and U7109 (N_7109,N_1091,N_2875);
nor U7110 (N_7110,N_1154,N_1187);
nor U7111 (N_7111,N_2356,N_1128);
nor U7112 (N_7112,N_4104,N_4697);
nand U7113 (N_7113,N_2378,N_3257);
or U7114 (N_7114,N_1658,N_3812);
or U7115 (N_7115,N_4614,N_205);
nand U7116 (N_7116,N_4569,N_3338);
and U7117 (N_7117,N_3881,N_2663);
or U7118 (N_7118,N_4399,N_3871);
nand U7119 (N_7119,N_3906,N_3054);
nor U7120 (N_7120,N_4378,N_1101);
and U7121 (N_7121,N_1960,N_866);
nand U7122 (N_7122,N_3939,N_2665);
and U7123 (N_7123,N_1103,N_576);
nor U7124 (N_7124,N_1129,N_726);
nand U7125 (N_7125,N_4411,N_4610);
and U7126 (N_7126,N_2716,N_4287);
nand U7127 (N_7127,N_1936,N_4134);
nor U7128 (N_7128,N_1841,N_4932);
and U7129 (N_7129,N_123,N_4476);
xor U7130 (N_7130,N_1318,N_2960);
nand U7131 (N_7131,N_1104,N_4828);
nand U7132 (N_7132,N_336,N_3647);
or U7133 (N_7133,N_1502,N_1497);
xor U7134 (N_7134,N_3744,N_4589);
nand U7135 (N_7135,N_1972,N_3911);
nor U7136 (N_7136,N_3142,N_3458);
or U7137 (N_7137,N_2457,N_4659);
xor U7138 (N_7138,N_3545,N_4630);
or U7139 (N_7139,N_2586,N_1606);
nor U7140 (N_7140,N_3400,N_4714);
nor U7141 (N_7141,N_1098,N_3820);
nor U7142 (N_7142,N_2973,N_717);
nand U7143 (N_7143,N_2797,N_4805);
or U7144 (N_7144,N_3728,N_2278);
and U7145 (N_7145,N_582,N_1026);
nand U7146 (N_7146,N_955,N_4584);
and U7147 (N_7147,N_3602,N_1912);
xor U7148 (N_7148,N_2913,N_2514);
xnor U7149 (N_7149,N_4677,N_2178);
or U7150 (N_7150,N_4693,N_997);
xnor U7151 (N_7151,N_1184,N_4040);
nor U7152 (N_7152,N_4209,N_877);
and U7153 (N_7153,N_449,N_3631);
or U7154 (N_7154,N_3971,N_241);
xnor U7155 (N_7155,N_4782,N_3227);
xor U7156 (N_7156,N_3409,N_4668);
and U7157 (N_7157,N_4429,N_2318);
xnor U7158 (N_7158,N_4995,N_2277);
or U7159 (N_7159,N_361,N_3920);
and U7160 (N_7160,N_1675,N_4596);
xnor U7161 (N_7161,N_1879,N_2268);
nor U7162 (N_7162,N_1514,N_4618);
and U7163 (N_7163,N_1892,N_788);
xor U7164 (N_7164,N_1788,N_1954);
and U7165 (N_7165,N_4132,N_4635);
xor U7166 (N_7166,N_4070,N_3500);
and U7167 (N_7167,N_1540,N_4407);
xor U7168 (N_7168,N_1499,N_2283);
or U7169 (N_7169,N_3395,N_4710);
and U7170 (N_7170,N_1793,N_4321);
or U7171 (N_7171,N_4732,N_1584);
xor U7172 (N_7172,N_4328,N_343);
and U7173 (N_7173,N_683,N_575);
or U7174 (N_7174,N_243,N_3841);
nor U7175 (N_7175,N_2860,N_2361);
xor U7176 (N_7176,N_3313,N_1809);
or U7177 (N_7177,N_3793,N_875);
xor U7178 (N_7178,N_4597,N_4534);
nor U7179 (N_7179,N_3860,N_1211);
or U7180 (N_7180,N_1073,N_1002);
nand U7181 (N_7181,N_1810,N_1832);
or U7182 (N_7182,N_602,N_3779);
nor U7183 (N_7183,N_116,N_3855);
and U7184 (N_7184,N_660,N_4340);
or U7185 (N_7185,N_1929,N_3701);
nand U7186 (N_7186,N_2307,N_2563);
nand U7187 (N_7187,N_2966,N_4811);
nand U7188 (N_7188,N_2060,N_2714);
nand U7189 (N_7189,N_4853,N_693);
xnor U7190 (N_7190,N_2977,N_4914);
and U7191 (N_7191,N_1260,N_2193);
and U7192 (N_7192,N_4691,N_3535);
nand U7193 (N_7193,N_4029,N_2772);
or U7194 (N_7194,N_4006,N_4506);
nor U7195 (N_7195,N_2879,N_673);
xor U7196 (N_7196,N_2687,N_2918);
nor U7197 (N_7197,N_1365,N_2705);
or U7198 (N_7198,N_2755,N_2129);
or U7199 (N_7199,N_341,N_1110);
nor U7200 (N_7200,N_1016,N_2320);
xnor U7201 (N_7201,N_2434,N_3613);
or U7202 (N_7202,N_3039,N_2390);
or U7203 (N_7203,N_321,N_1237);
and U7204 (N_7204,N_2513,N_3730);
or U7205 (N_7205,N_4553,N_2108);
nand U7206 (N_7206,N_3699,N_4152);
or U7207 (N_7207,N_1304,N_4073);
xnor U7208 (N_7208,N_589,N_3894);
xnor U7209 (N_7209,N_709,N_4936);
xor U7210 (N_7210,N_379,N_2359);
or U7211 (N_7211,N_1229,N_3491);
or U7212 (N_7212,N_3510,N_1165);
xor U7213 (N_7213,N_4063,N_4590);
or U7214 (N_7214,N_3766,N_3555);
or U7215 (N_7215,N_431,N_2371);
nor U7216 (N_7216,N_3533,N_4112);
xnor U7217 (N_7217,N_4666,N_1752);
nor U7218 (N_7218,N_567,N_2414);
nand U7219 (N_7219,N_1724,N_3433);
xnor U7220 (N_7220,N_3089,N_3402);
and U7221 (N_7221,N_886,N_1626);
nor U7222 (N_7222,N_3796,N_4068);
or U7223 (N_7223,N_1815,N_1940);
and U7224 (N_7224,N_4330,N_4858);
and U7225 (N_7225,N_293,N_1852);
and U7226 (N_7226,N_4123,N_2340);
and U7227 (N_7227,N_1749,N_368);
xor U7228 (N_7228,N_545,N_560);
xnor U7229 (N_7229,N_3123,N_549);
or U7230 (N_7230,N_1625,N_840);
nor U7231 (N_7231,N_2867,N_1241);
or U7232 (N_7232,N_2938,N_1261);
xnor U7233 (N_7233,N_1900,N_2675);
xnor U7234 (N_7234,N_3183,N_2940);
and U7235 (N_7235,N_1280,N_108);
xor U7236 (N_7236,N_1629,N_1630);
nor U7237 (N_7237,N_4278,N_3962);
nor U7238 (N_7238,N_792,N_3162);
nand U7239 (N_7239,N_372,N_4023);
and U7240 (N_7240,N_2228,N_3280);
and U7241 (N_7241,N_3034,N_4384);
or U7242 (N_7242,N_3055,N_598);
nand U7243 (N_7243,N_458,N_4636);
and U7244 (N_7244,N_3103,N_4291);
nand U7245 (N_7245,N_1219,N_433);
xnor U7246 (N_7246,N_4848,N_2547);
and U7247 (N_7247,N_3833,N_1044);
and U7248 (N_7248,N_54,N_4796);
xor U7249 (N_7249,N_4795,N_4268);
and U7250 (N_7250,N_1001,N_4831);
and U7251 (N_7251,N_4546,N_4498);
nand U7252 (N_7252,N_3527,N_2386);
xor U7253 (N_7253,N_1828,N_663);
and U7254 (N_7254,N_3541,N_503);
and U7255 (N_7255,N_1401,N_544);
xor U7256 (N_7256,N_4276,N_179);
nand U7257 (N_7257,N_4119,N_3025);
xor U7258 (N_7258,N_312,N_1369);
and U7259 (N_7259,N_1602,N_2134);
or U7260 (N_7260,N_3922,N_4187);
and U7261 (N_7261,N_2827,N_4663);
nand U7262 (N_7262,N_4593,N_3096);
and U7263 (N_7263,N_1803,N_3474);
xnor U7264 (N_7264,N_4760,N_4382);
or U7265 (N_7265,N_4375,N_2241);
nor U7266 (N_7266,N_4916,N_4270);
or U7267 (N_7267,N_3948,N_3537);
xor U7268 (N_7268,N_2243,N_3633);
and U7269 (N_7269,N_1539,N_1516);
nand U7270 (N_7270,N_1851,N_2570);
or U7271 (N_7271,N_887,N_3706);
or U7272 (N_7272,N_4460,N_2487);
nor U7273 (N_7273,N_934,N_3585);
or U7274 (N_7274,N_4461,N_3112);
xnor U7275 (N_7275,N_3619,N_2295);
xnor U7276 (N_7276,N_3052,N_3932);
nand U7277 (N_7277,N_1174,N_837);
xnor U7278 (N_7278,N_3964,N_1153);
or U7279 (N_7279,N_2724,N_384);
xor U7280 (N_7280,N_4015,N_3627);
nor U7281 (N_7281,N_2081,N_1454);
and U7282 (N_7282,N_2333,N_2770);
nand U7283 (N_7283,N_832,N_2783);
nand U7284 (N_7284,N_2553,N_359);
nand U7285 (N_7285,N_98,N_4924);
nand U7286 (N_7286,N_4218,N_3349);
and U7287 (N_7287,N_1631,N_1888);
nand U7288 (N_7288,N_1202,N_4163);
nor U7289 (N_7289,N_4594,N_1198);
and U7290 (N_7290,N_2509,N_2008);
or U7291 (N_7291,N_4670,N_3522);
nor U7292 (N_7292,N_1032,N_3632);
xnor U7293 (N_7293,N_77,N_4725);
and U7294 (N_7294,N_4925,N_3817);
nand U7295 (N_7295,N_680,N_3573);
nor U7296 (N_7296,N_2166,N_3258);
and U7297 (N_7297,N_2032,N_3274);
nand U7298 (N_7298,N_3222,N_1964);
nand U7299 (N_7299,N_1047,N_4743);
xor U7300 (N_7300,N_3290,N_133);
nor U7301 (N_7301,N_1360,N_710);
xor U7302 (N_7302,N_2781,N_640);
nor U7303 (N_7303,N_4086,N_3813);
nor U7304 (N_7304,N_3463,N_3211);
nand U7305 (N_7305,N_437,N_3686);
nor U7306 (N_7306,N_2353,N_4148);
and U7307 (N_7307,N_2480,N_1472);
nand U7308 (N_7308,N_1574,N_569);
and U7309 (N_7309,N_3269,N_3325);
or U7310 (N_7310,N_1465,N_1819);
and U7311 (N_7311,N_2317,N_3243);
and U7312 (N_7312,N_2846,N_3967);
xor U7313 (N_7313,N_3556,N_4254);
or U7314 (N_7314,N_2267,N_2824);
nand U7315 (N_7315,N_4823,N_147);
xnor U7316 (N_7316,N_2112,N_3407);
nand U7317 (N_7317,N_3003,N_4079);
nand U7318 (N_7318,N_1159,N_4585);
xnor U7319 (N_7319,N_3944,N_3079);
nand U7320 (N_7320,N_3399,N_2172);
nor U7321 (N_7321,N_1282,N_4503);
nand U7322 (N_7322,N_1677,N_4655);
nor U7323 (N_7323,N_1920,N_4215);
and U7324 (N_7324,N_3664,N_4785);
nor U7325 (N_7325,N_4783,N_2423);
nor U7326 (N_7326,N_2594,N_4627);
nor U7327 (N_7327,N_3371,N_1835);
nor U7328 (N_7328,N_977,N_3310);
or U7329 (N_7329,N_2839,N_2996);
xnor U7330 (N_7330,N_893,N_830);
nor U7331 (N_7331,N_2316,N_4477);
nand U7332 (N_7332,N_45,N_3685);
and U7333 (N_7333,N_2276,N_1373);
nor U7334 (N_7334,N_2208,N_3390);
and U7335 (N_7335,N_2642,N_1771);
or U7336 (N_7336,N_2477,N_1670);
nor U7337 (N_7337,N_702,N_4812);
xnor U7338 (N_7338,N_4551,N_3111);
xnor U7339 (N_7339,N_2736,N_4206);
xnor U7340 (N_7340,N_2358,N_4753);
or U7341 (N_7341,N_2231,N_4434);
nor U7342 (N_7342,N_85,N_4444);
nor U7343 (N_7343,N_3455,N_4074);
nand U7344 (N_7344,N_1435,N_3854);
and U7345 (N_7345,N_2639,N_4021);
and U7346 (N_7346,N_3385,N_3608);
nor U7347 (N_7347,N_1445,N_3437);
nand U7348 (N_7348,N_1273,N_2481);
or U7349 (N_7349,N_479,N_3294);
nand U7350 (N_7350,N_2627,N_1838);
nand U7351 (N_7351,N_4228,N_4474);
and U7352 (N_7352,N_894,N_3024);
nor U7353 (N_7353,N_4560,N_3124);
xnor U7354 (N_7354,N_1203,N_2990);
or U7355 (N_7355,N_732,N_4412);
nand U7356 (N_7356,N_3442,N_4160);
xor U7357 (N_7357,N_4443,N_1523);
xnor U7358 (N_7358,N_1554,N_139);
nand U7359 (N_7359,N_1636,N_1163);
xnor U7360 (N_7360,N_3991,N_1244);
xnor U7361 (N_7361,N_97,N_1870);
nor U7362 (N_7362,N_3061,N_3978);
or U7363 (N_7363,N_659,N_520);
xor U7364 (N_7364,N_597,N_2753);
xnor U7365 (N_7365,N_1393,N_3356);
nor U7366 (N_7366,N_3530,N_4928);
nand U7367 (N_7367,N_452,N_4774);
and U7368 (N_7368,N_2161,N_3230);
nor U7369 (N_7369,N_3839,N_4981);
or U7370 (N_7370,N_746,N_2415);
xnor U7371 (N_7371,N_800,N_4544);
and U7372 (N_7372,N_2063,N_4616);
xnor U7373 (N_7373,N_2030,N_2673);
xnor U7374 (N_7374,N_1185,N_1550);
nor U7375 (N_7375,N_4300,N_1921);
nor U7376 (N_7376,N_1941,N_2280);
and U7377 (N_7377,N_3507,N_2177);
xnor U7378 (N_7378,N_2322,N_4048);
or U7379 (N_7379,N_697,N_4018);
and U7380 (N_7380,N_1480,N_3693);
or U7381 (N_7381,N_1031,N_2743);
nand U7382 (N_7382,N_3022,N_4127);
or U7383 (N_7383,N_1767,N_170);
or U7384 (N_7384,N_1580,N_4034);
or U7385 (N_7385,N_306,N_1581);
and U7386 (N_7386,N_1430,N_2417);
nand U7387 (N_7387,N_4438,N_2896);
xnor U7388 (N_7388,N_3440,N_2533);
and U7389 (N_7389,N_3353,N_1162);
xnor U7390 (N_7390,N_3651,N_4130);
and U7391 (N_7391,N_4899,N_3147);
nor U7392 (N_7392,N_4825,N_3709);
nand U7393 (N_7393,N_3984,N_4374);
nand U7394 (N_7394,N_391,N_472);
and U7395 (N_7395,N_4326,N_3297);
and U7396 (N_7396,N_2929,N_2780);
nand U7397 (N_7397,N_2427,N_3364);
nor U7398 (N_7398,N_3678,N_1246);
nor U7399 (N_7399,N_3487,N_4117);
and U7400 (N_7400,N_2945,N_2933);
and U7401 (N_7401,N_2998,N_2947);
nand U7402 (N_7402,N_1114,N_1438);
and U7403 (N_7403,N_2404,N_486);
nand U7404 (N_7404,N_1370,N_1825);
nor U7405 (N_7405,N_436,N_4462);
nand U7406 (N_7406,N_3267,N_4178);
and U7407 (N_7407,N_4113,N_2394);
nor U7408 (N_7408,N_1067,N_2479);
or U7409 (N_7409,N_3097,N_514);
xnor U7410 (N_7410,N_725,N_2559);
nor U7411 (N_7411,N_1551,N_3016);
and U7412 (N_7412,N_3060,N_273);
and U7413 (N_7413,N_1108,N_4781);
xor U7414 (N_7414,N_1359,N_244);
xnor U7415 (N_7415,N_1991,N_1494);
xnor U7416 (N_7416,N_4927,N_1758);
nor U7417 (N_7417,N_262,N_4682);
nand U7418 (N_7418,N_4233,N_4583);
and U7419 (N_7419,N_4450,N_390);
nor U7420 (N_7420,N_3808,N_3181);
nor U7421 (N_7421,N_1555,N_464);
and U7422 (N_7422,N_3048,N_4595);
nor U7423 (N_7423,N_2543,N_3804);
xnor U7424 (N_7424,N_188,N_2792);
nor U7425 (N_7425,N_901,N_4421);
nand U7426 (N_7426,N_3275,N_2204);
nand U7427 (N_7427,N_1313,N_2881);
or U7428 (N_7428,N_4175,N_485);
xor U7429 (N_7429,N_3365,N_4827);
xor U7430 (N_7430,N_1238,N_4240);
or U7431 (N_7431,N_4729,N_1155);
and U7432 (N_7432,N_3017,N_1868);
and U7433 (N_7433,N_3179,N_799);
nor U7434 (N_7434,N_3093,N_2826);
nand U7435 (N_7435,N_1291,N_566);
or U7436 (N_7436,N_1412,N_2808);
xor U7437 (N_7437,N_1930,N_3901);
xnor U7438 (N_7438,N_3262,N_2732);
and U7439 (N_7439,N_1432,N_2004);
xnor U7440 (N_7440,N_3240,N_0);
or U7441 (N_7441,N_4337,N_774);
or U7442 (N_7442,N_3161,N_1042);
or U7443 (N_7443,N_459,N_1922);
xor U7444 (N_7444,N_2734,N_2804);
and U7445 (N_7445,N_882,N_2526);
xor U7446 (N_7446,N_4972,N_1157);
xnor U7447 (N_7447,N_2900,N_2970);
or U7448 (N_7448,N_2469,N_1385);
or U7449 (N_7449,N_686,N_3304);
or U7450 (N_7450,N_145,N_4882);
or U7451 (N_7451,N_4513,N_1328);
nand U7452 (N_7452,N_1949,N_591);
or U7453 (N_7453,N_624,N_1529);
nand U7454 (N_7454,N_626,N_4686);
nand U7455 (N_7455,N_2517,N_4186);
and U7456 (N_7456,N_3180,N_3420);
and U7457 (N_7457,N_3910,N_2459);
nand U7458 (N_7458,N_2893,N_1644);
and U7459 (N_7459,N_2150,N_3013);
nor U7460 (N_7460,N_3981,N_2803);
nor U7461 (N_7461,N_2731,N_4859);
nor U7462 (N_7462,N_2782,N_2849);
or U7463 (N_7463,N_187,N_1239);
or U7464 (N_7464,N_4638,N_4183);
or U7465 (N_7465,N_3878,N_3597);
and U7466 (N_7466,N_1744,N_1723);
or U7467 (N_7467,N_1797,N_4071);
and U7468 (N_7468,N_2993,N_1969);
and U7469 (N_7469,N_2437,N_3057);
xor U7470 (N_7470,N_71,N_4239);
nor U7471 (N_7471,N_3100,N_2617);
xor U7472 (N_7472,N_552,N_1303);
xnor U7473 (N_7473,N_3414,N_4650);
nand U7474 (N_7474,N_1119,N_3497);
nor U7475 (N_7475,N_539,N_4545);
and U7476 (N_7476,N_1080,N_1730);
nand U7477 (N_7477,N_46,N_3610);
nand U7478 (N_7478,N_1138,N_2119);
or U7479 (N_7479,N_2637,N_2661);
or U7480 (N_7480,N_944,N_1420);
nand U7481 (N_7481,N_3228,N_3660);
nand U7482 (N_7482,N_59,N_3218);
nor U7483 (N_7483,N_657,N_3960);
nor U7484 (N_7484,N_993,N_1691);
or U7485 (N_7485,N_4459,N_2887);
and U7486 (N_7486,N_150,N_2955);
or U7487 (N_7487,N_3178,N_4586);
xnor U7488 (N_7488,N_4851,N_4064);
and U7489 (N_7489,N_4057,N_546);
nand U7490 (N_7490,N_1088,N_1729);
nand U7491 (N_7491,N_488,N_3587);
or U7492 (N_7492,N_4640,N_1635);
xnor U7493 (N_7493,N_1807,N_2075);
xor U7494 (N_7494,N_3305,N_773);
nand U7495 (N_7495,N_1739,N_4124);
nor U7496 (N_7496,N_3005,N_279);
and U7497 (N_7497,N_1215,N_3598);
nor U7498 (N_7498,N_4519,N_4406);
and U7499 (N_7499,N_913,N_3523);
and U7500 (N_7500,N_2485,N_1593);
xnor U7501 (N_7501,N_133,N_1934);
nor U7502 (N_7502,N_3905,N_1601);
xor U7503 (N_7503,N_4336,N_4965);
nand U7504 (N_7504,N_3935,N_1512);
nand U7505 (N_7505,N_4566,N_294);
xor U7506 (N_7506,N_4734,N_1917);
nor U7507 (N_7507,N_425,N_806);
xor U7508 (N_7508,N_1758,N_4540);
nand U7509 (N_7509,N_4185,N_261);
xnor U7510 (N_7510,N_3771,N_2125);
xor U7511 (N_7511,N_3584,N_940);
and U7512 (N_7512,N_1940,N_2104);
or U7513 (N_7513,N_695,N_2342);
and U7514 (N_7514,N_4025,N_1133);
xnor U7515 (N_7515,N_2602,N_1676);
xnor U7516 (N_7516,N_2535,N_4180);
nor U7517 (N_7517,N_933,N_850);
xnor U7518 (N_7518,N_2089,N_3444);
and U7519 (N_7519,N_1103,N_3940);
nor U7520 (N_7520,N_3511,N_3889);
nand U7521 (N_7521,N_3120,N_2547);
or U7522 (N_7522,N_3078,N_846);
nand U7523 (N_7523,N_1333,N_1789);
or U7524 (N_7524,N_1879,N_3551);
xnor U7525 (N_7525,N_175,N_1879);
and U7526 (N_7526,N_2245,N_2090);
xnor U7527 (N_7527,N_2659,N_3719);
or U7528 (N_7528,N_4335,N_1293);
xnor U7529 (N_7529,N_2502,N_2351);
xnor U7530 (N_7530,N_635,N_4972);
and U7531 (N_7531,N_1838,N_2837);
nand U7532 (N_7532,N_932,N_4985);
nand U7533 (N_7533,N_4089,N_3824);
nor U7534 (N_7534,N_992,N_166);
and U7535 (N_7535,N_2545,N_995);
or U7536 (N_7536,N_1749,N_692);
and U7537 (N_7537,N_3120,N_4429);
nand U7538 (N_7538,N_1541,N_538);
and U7539 (N_7539,N_2951,N_1497);
nor U7540 (N_7540,N_4742,N_581);
nor U7541 (N_7541,N_251,N_669);
xor U7542 (N_7542,N_2308,N_138);
nor U7543 (N_7543,N_4109,N_3309);
nand U7544 (N_7544,N_1469,N_4890);
and U7545 (N_7545,N_1755,N_3821);
and U7546 (N_7546,N_970,N_1684);
nand U7547 (N_7547,N_4681,N_2464);
nor U7548 (N_7548,N_1745,N_3902);
xnor U7549 (N_7549,N_4791,N_756);
and U7550 (N_7550,N_1499,N_4933);
and U7551 (N_7551,N_2459,N_3988);
nor U7552 (N_7552,N_616,N_1946);
nand U7553 (N_7553,N_2860,N_3208);
or U7554 (N_7554,N_4553,N_1892);
xor U7555 (N_7555,N_3170,N_4006);
or U7556 (N_7556,N_4002,N_1366);
xor U7557 (N_7557,N_980,N_3082);
xnor U7558 (N_7558,N_4666,N_4147);
and U7559 (N_7559,N_4854,N_2111);
or U7560 (N_7560,N_1607,N_1545);
nor U7561 (N_7561,N_2755,N_4067);
nor U7562 (N_7562,N_2246,N_3714);
xor U7563 (N_7563,N_4984,N_3465);
or U7564 (N_7564,N_3995,N_4687);
or U7565 (N_7565,N_1235,N_2365);
nor U7566 (N_7566,N_4054,N_3519);
xor U7567 (N_7567,N_214,N_2194);
and U7568 (N_7568,N_1759,N_954);
xor U7569 (N_7569,N_3886,N_2832);
nor U7570 (N_7570,N_4186,N_4671);
nand U7571 (N_7571,N_1888,N_1122);
xnor U7572 (N_7572,N_1143,N_4902);
xor U7573 (N_7573,N_3193,N_2327);
nand U7574 (N_7574,N_1016,N_4335);
or U7575 (N_7575,N_770,N_2660);
and U7576 (N_7576,N_316,N_977);
nor U7577 (N_7577,N_3796,N_2854);
or U7578 (N_7578,N_949,N_554);
or U7579 (N_7579,N_3461,N_912);
or U7580 (N_7580,N_4597,N_1422);
xor U7581 (N_7581,N_3504,N_1141);
or U7582 (N_7582,N_415,N_3249);
or U7583 (N_7583,N_3529,N_20);
nor U7584 (N_7584,N_4866,N_1864);
xnor U7585 (N_7585,N_918,N_2718);
nand U7586 (N_7586,N_4500,N_4926);
xnor U7587 (N_7587,N_801,N_4115);
and U7588 (N_7588,N_1316,N_3343);
and U7589 (N_7589,N_629,N_872);
nand U7590 (N_7590,N_637,N_347);
nand U7591 (N_7591,N_2614,N_2245);
or U7592 (N_7592,N_1930,N_2856);
xor U7593 (N_7593,N_3025,N_2632);
nor U7594 (N_7594,N_4455,N_137);
nor U7595 (N_7595,N_135,N_3950);
xor U7596 (N_7596,N_2320,N_83);
or U7597 (N_7597,N_3526,N_3361);
xor U7598 (N_7598,N_1517,N_2910);
nor U7599 (N_7599,N_1407,N_4502);
or U7600 (N_7600,N_3382,N_4310);
xnor U7601 (N_7601,N_3427,N_1684);
xnor U7602 (N_7602,N_1209,N_346);
and U7603 (N_7603,N_3327,N_3707);
xnor U7604 (N_7604,N_4725,N_3927);
or U7605 (N_7605,N_1414,N_3533);
or U7606 (N_7606,N_2730,N_838);
xnor U7607 (N_7607,N_892,N_3059);
xor U7608 (N_7608,N_3435,N_2209);
xnor U7609 (N_7609,N_694,N_3575);
or U7610 (N_7610,N_2978,N_2733);
nor U7611 (N_7611,N_3315,N_2093);
nor U7612 (N_7612,N_3687,N_1337);
nor U7613 (N_7613,N_466,N_2272);
xor U7614 (N_7614,N_2833,N_4879);
and U7615 (N_7615,N_1351,N_3522);
and U7616 (N_7616,N_3951,N_4783);
nor U7617 (N_7617,N_1169,N_2965);
or U7618 (N_7618,N_569,N_4326);
and U7619 (N_7619,N_66,N_1655);
nor U7620 (N_7620,N_862,N_3827);
and U7621 (N_7621,N_839,N_3952);
nor U7622 (N_7622,N_2446,N_2738);
or U7623 (N_7623,N_4021,N_4929);
or U7624 (N_7624,N_287,N_4001);
nand U7625 (N_7625,N_515,N_1231);
and U7626 (N_7626,N_4664,N_1642);
and U7627 (N_7627,N_4209,N_2071);
or U7628 (N_7628,N_4603,N_2466);
nand U7629 (N_7629,N_4058,N_3392);
nor U7630 (N_7630,N_122,N_4781);
nand U7631 (N_7631,N_720,N_3476);
xor U7632 (N_7632,N_84,N_289);
nand U7633 (N_7633,N_4553,N_1278);
nor U7634 (N_7634,N_200,N_3744);
or U7635 (N_7635,N_1527,N_258);
xor U7636 (N_7636,N_1833,N_943);
or U7637 (N_7637,N_4101,N_3919);
or U7638 (N_7638,N_3035,N_3389);
nand U7639 (N_7639,N_3510,N_4904);
or U7640 (N_7640,N_391,N_496);
and U7641 (N_7641,N_1377,N_3268);
and U7642 (N_7642,N_3611,N_4963);
xnor U7643 (N_7643,N_4004,N_65);
nor U7644 (N_7644,N_3576,N_726);
and U7645 (N_7645,N_4178,N_2223);
nand U7646 (N_7646,N_1306,N_4237);
xnor U7647 (N_7647,N_3540,N_2223);
nand U7648 (N_7648,N_2218,N_1729);
or U7649 (N_7649,N_2699,N_3220);
xor U7650 (N_7650,N_1180,N_346);
and U7651 (N_7651,N_1846,N_278);
or U7652 (N_7652,N_4154,N_2249);
nor U7653 (N_7653,N_2677,N_1197);
and U7654 (N_7654,N_392,N_3404);
or U7655 (N_7655,N_4106,N_3419);
xnor U7656 (N_7656,N_3949,N_932);
or U7657 (N_7657,N_1428,N_2064);
and U7658 (N_7658,N_2527,N_3459);
nor U7659 (N_7659,N_926,N_3921);
nand U7660 (N_7660,N_4598,N_551);
nand U7661 (N_7661,N_1925,N_585);
xnor U7662 (N_7662,N_3293,N_4693);
nand U7663 (N_7663,N_1143,N_2804);
nand U7664 (N_7664,N_4903,N_4638);
or U7665 (N_7665,N_653,N_339);
and U7666 (N_7666,N_1780,N_4633);
xor U7667 (N_7667,N_1655,N_1753);
or U7668 (N_7668,N_1024,N_4779);
or U7669 (N_7669,N_73,N_4177);
or U7670 (N_7670,N_3398,N_2066);
nor U7671 (N_7671,N_2255,N_833);
and U7672 (N_7672,N_1882,N_1239);
and U7673 (N_7673,N_122,N_1239);
and U7674 (N_7674,N_832,N_1587);
xor U7675 (N_7675,N_494,N_4010);
nand U7676 (N_7676,N_626,N_1129);
nand U7677 (N_7677,N_2551,N_1573);
nand U7678 (N_7678,N_462,N_3443);
or U7679 (N_7679,N_1410,N_1943);
or U7680 (N_7680,N_3556,N_3290);
nor U7681 (N_7681,N_2468,N_1060);
or U7682 (N_7682,N_4927,N_2730);
nand U7683 (N_7683,N_2241,N_3335);
and U7684 (N_7684,N_4790,N_2667);
xnor U7685 (N_7685,N_319,N_77);
or U7686 (N_7686,N_2534,N_71);
or U7687 (N_7687,N_3254,N_3018);
xor U7688 (N_7688,N_1743,N_3607);
nand U7689 (N_7689,N_3648,N_3751);
xnor U7690 (N_7690,N_4846,N_4566);
and U7691 (N_7691,N_3074,N_4421);
nor U7692 (N_7692,N_3983,N_2860);
nand U7693 (N_7693,N_863,N_3402);
nor U7694 (N_7694,N_4032,N_1800);
nand U7695 (N_7695,N_821,N_482);
nand U7696 (N_7696,N_4266,N_30);
xnor U7697 (N_7697,N_3717,N_70);
or U7698 (N_7698,N_4548,N_1641);
or U7699 (N_7699,N_3297,N_3557);
nor U7700 (N_7700,N_2221,N_131);
nand U7701 (N_7701,N_4309,N_1000);
and U7702 (N_7702,N_3738,N_2623);
nor U7703 (N_7703,N_214,N_4865);
xnor U7704 (N_7704,N_4155,N_2823);
xnor U7705 (N_7705,N_2037,N_1436);
nand U7706 (N_7706,N_2028,N_1102);
nor U7707 (N_7707,N_883,N_476);
nand U7708 (N_7708,N_3964,N_3194);
xnor U7709 (N_7709,N_4871,N_2617);
or U7710 (N_7710,N_1023,N_915);
nor U7711 (N_7711,N_3387,N_1910);
xor U7712 (N_7712,N_3717,N_3106);
nor U7713 (N_7713,N_3198,N_2626);
nor U7714 (N_7714,N_3076,N_3016);
or U7715 (N_7715,N_324,N_3183);
nor U7716 (N_7716,N_230,N_3848);
xnor U7717 (N_7717,N_794,N_2883);
nand U7718 (N_7718,N_1868,N_3782);
and U7719 (N_7719,N_3086,N_4718);
and U7720 (N_7720,N_3377,N_1739);
xnor U7721 (N_7721,N_1539,N_4201);
xnor U7722 (N_7722,N_2055,N_1826);
nor U7723 (N_7723,N_4313,N_2208);
nand U7724 (N_7724,N_4320,N_4185);
or U7725 (N_7725,N_2779,N_2952);
or U7726 (N_7726,N_1549,N_1921);
or U7727 (N_7727,N_1935,N_3328);
xnor U7728 (N_7728,N_2314,N_1418);
or U7729 (N_7729,N_3208,N_3112);
nor U7730 (N_7730,N_4843,N_648);
xnor U7731 (N_7731,N_1912,N_1318);
and U7732 (N_7732,N_2780,N_626);
or U7733 (N_7733,N_1441,N_3596);
xor U7734 (N_7734,N_766,N_3007);
and U7735 (N_7735,N_2017,N_2144);
nand U7736 (N_7736,N_3865,N_3667);
and U7737 (N_7737,N_514,N_4490);
and U7738 (N_7738,N_670,N_4534);
or U7739 (N_7739,N_4322,N_2114);
nand U7740 (N_7740,N_1744,N_2414);
or U7741 (N_7741,N_3493,N_4246);
xor U7742 (N_7742,N_3087,N_592);
nor U7743 (N_7743,N_3864,N_3491);
or U7744 (N_7744,N_1238,N_1696);
or U7745 (N_7745,N_4744,N_679);
nand U7746 (N_7746,N_2138,N_4796);
nand U7747 (N_7747,N_2919,N_790);
and U7748 (N_7748,N_564,N_3325);
or U7749 (N_7749,N_3043,N_3064);
and U7750 (N_7750,N_281,N_1858);
nor U7751 (N_7751,N_4029,N_2643);
or U7752 (N_7752,N_1991,N_2042);
and U7753 (N_7753,N_2179,N_2538);
or U7754 (N_7754,N_677,N_3604);
and U7755 (N_7755,N_3909,N_4010);
nand U7756 (N_7756,N_4140,N_3273);
xor U7757 (N_7757,N_4169,N_4269);
nor U7758 (N_7758,N_2820,N_1633);
nor U7759 (N_7759,N_2825,N_836);
nor U7760 (N_7760,N_3207,N_535);
nor U7761 (N_7761,N_4021,N_3328);
xnor U7762 (N_7762,N_3424,N_2044);
nor U7763 (N_7763,N_1776,N_214);
and U7764 (N_7764,N_1495,N_4288);
and U7765 (N_7765,N_2472,N_4341);
xor U7766 (N_7766,N_2193,N_2991);
or U7767 (N_7767,N_4402,N_2962);
nand U7768 (N_7768,N_4763,N_1368);
or U7769 (N_7769,N_2008,N_1420);
nor U7770 (N_7770,N_1083,N_3309);
xnor U7771 (N_7771,N_280,N_1767);
and U7772 (N_7772,N_490,N_3822);
and U7773 (N_7773,N_729,N_4335);
nand U7774 (N_7774,N_4078,N_4780);
nor U7775 (N_7775,N_1393,N_130);
xnor U7776 (N_7776,N_1879,N_4764);
xnor U7777 (N_7777,N_1047,N_2583);
xnor U7778 (N_7778,N_1802,N_3936);
nor U7779 (N_7779,N_3114,N_2105);
xor U7780 (N_7780,N_1842,N_663);
or U7781 (N_7781,N_3803,N_1752);
xnor U7782 (N_7782,N_1296,N_4962);
and U7783 (N_7783,N_7,N_4479);
nand U7784 (N_7784,N_2337,N_4186);
or U7785 (N_7785,N_4054,N_3421);
nand U7786 (N_7786,N_2801,N_2209);
nand U7787 (N_7787,N_4716,N_4238);
and U7788 (N_7788,N_338,N_717);
and U7789 (N_7789,N_3406,N_899);
nor U7790 (N_7790,N_3419,N_4762);
nand U7791 (N_7791,N_3191,N_837);
nor U7792 (N_7792,N_2271,N_3364);
nand U7793 (N_7793,N_1193,N_1010);
xnor U7794 (N_7794,N_3240,N_2573);
nand U7795 (N_7795,N_3717,N_4152);
nor U7796 (N_7796,N_1970,N_3826);
and U7797 (N_7797,N_1072,N_1546);
nor U7798 (N_7798,N_3623,N_4011);
nor U7799 (N_7799,N_3563,N_2445);
or U7800 (N_7800,N_3661,N_3192);
nor U7801 (N_7801,N_1793,N_3081);
nand U7802 (N_7802,N_222,N_4625);
nor U7803 (N_7803,N_4354,N_3027);
and U7804 (N_7804,N_4714,N_2758);
or U7805 (N_7805,N_3653,N_1354);
and U7806 (N_7806,N_4575,N_3033);
and U7807 (N_7807,N_3352,N_4296);
xnor U7808 (N_7808,N_1068,N_845);
nand U7809 (N_7809,N_4854,N_4660);
nor U7810 (N_7810,N_3905,N_3818);
and U7811 (N_7811,N_1414,N_1956);
xnor U7812 (N_7812,N_607,N_807);
xnor U7813 (N_7813,N_164,N_1924);
xnor U7814 (N_7814,N_1962,N_1634);
xnor U7815 (N_7815,N_1214,N_3575);
xor U7816 (N_7816,N_4632,N_4285);
nand U7817 (N_7817,N_2018,N_294);
or U7818 (N_7818,N_2064,N_3995);
xnor U7819 (N_7819,N_1943,N_4489);
and U7820 (N_7820,N_1200,N_91);
nor U7821 (N_7821,N_4329,N_4669);
nor U7822 (N_7822,N_4771,N_4848);
nor U7823 (N_7823,N_4812,N_1715);
nand U7824 (N_7824,N_3382,N_4903);
and U7825 (N_7825,N_813,N_4294);
xnor U7826 (N_7826,N_1327,N_3229);
nand U7827 (N_7827,N_2479,N_2689);
nand U7828 (N_7828,N_4553,N_4695);
and U7829 (N_7829,N_4291,N_3165);
and U7830 (N_7830,N_2284,N_1093);
nor U7831 (N_7831,N_2948,N_868);
xnor U7832 (N_7832,N_1624,N_3410);
xor U7833 (N_7833,N_3686,N_4316);
nand U7834 (N_7834,N_4579,N_2351);
or U7835 (N_7835,N_1125,N_4870);
nor U7836 (N_7836,N_1220,N_83);
xor U7837 (N_7837,N_4613,N_795);
nand U7838 (N_7838,N_1858,N_1987);
xnor U7839 (N_7839,N_4812,N_633);
nand U7840 (N_7840,N_1193,N_1690);
nor U7841 (N_7841,N_4369,N_3827);
nor U7842 (N_7842,N_1084,N_1212);
nand U7843 (N_7843,N_1527,N_3361);
nor U7844 (N_7844,N_1964,N_4976);
or U7845 (N_7845,N_297,N_3630);
and U7846 (N_7846,N_3354,N_500);
nor U7847 (N_7847,N_3867,N_4520);
nand U7848 (N_7848,N_4893,N_4879);
or U7849 (N_7849,N_1699,N_661);
xor U7850 (N_7850,N_3232,N_3855);
xor U7851 (N_7851,N_4804,N_2402);
nor U7852 (N_7852,N_4835,N_510);
nand U7853 (N_7853,N_50,N_4594);
xor U7854 (N_7854,N_1279,N_2935);
nor U7855 (N_7855,N_36,N_3405);
nor U7856 (N_7856,N_865,N_3539);
and U7857 (N_7857,N_664,N_3171);
nor U7858 (N_7858,N_3318,N_1858);
xnor U7859 (N_7859,N_4486,N_2049);
nor U7860 (N_7860,N_4733,N_445);
xor U7861 (N_7861,N_1866,N_2437);
xor U7862 (N_7862,N_4141,N_4063);
or U7863 (N_7863,N_4310,N_1172);
or U7864 (N_7864,N_3952,N_3709);
nor U7865 (N_7865,N_4810,N_4626);
xor U7866 (N_7866,N_4213,N_1347);
nor U7867 (N_7867,N_4191,N_2052);
nor U7868 (N_7868,N_250,N_1636);
or U7869 (N_7869,N_1941,N_4652);
and U7870 (N_7870,N_3784,N_1312);
and U7871 (N_7871,N_2833,N_2646);
nor U7872 (N_7872,N_3095,N_4677);
and U7873 (N_7873,N_3438,N_3365);
and U7874 (N_7874,N_216,N_863);
nand U7875 (N_7875,N_4654,N_3844);
or U7876 (N_7876,N_3087,N_1000);
or U7877 (N_7877,N_331,N_3012);
nand U7878 (N_7878,N_4128,N_1079);
nand U7879 (N_7879,N_1102,N_1272);
nand U7880 (N_7880,N_893,N_1033);
nand U7881 (N_7881,N_4807,N_3188);
xnor U7882 (N_7882,N_4130,N_452);
nor U7883 (N_7883,N_379,N_3105);
or U7884 (N_7884,N_2631,N_3762);
nor U7885 (N_7885,N_2806,N_4327);
nand U7886 (N_7886,N_4329,N_283);
nand U7887 (N_7887,N_4054,N_3189);
or U7888 (N_7888,N_2437,N_4105);
or U7889 (N_7889,N_1539,N_4566);
or U7890 (N_7890,N_4813,N_2587);
and U7891 (N_7891,N_3485,N_846);
xor U7892 (N_7892,N_3778,N_3628);
nor U7893 (N_7893,N_1430,N_2504);
nor U7894 (N_7894,N_511,N_465);
xor U7895 (N_7895,N_2561,N_2448);
or U7896 (N_7896,N_1478,N_1512);
and U7897 (N_7897,N_4828,N_2268);
nand U7898 (N_7898,N_2418,N_4956);
nand U7899 (N_7899,N_609,N_1848);
nor U7900 (N_7900,N_1698,N_4625);
nor U7901 (N_7901,N_4249,N_728);
nor U7902 (N_7902,N_3878,N_4593);
nor U7903 (N_7903,N_4559,N_3899);
and U7904 (N_7904,N_842,N_113);
and U7905 (N_7905,N_4403,N_1988);
xor U7906 (N_7906,N_2877,N_4189);
and U7907 (N_7907,N_2315,N_3517);
or U7908 (N_7908,N_1095,N_4256);
nor U7909 (N_7909,N_1097,N_1502);
and U7910 (N_7910,N_3680,N_1149);
nor U7911 (N_7911,N_274,N_600);
nand U7912 (N_7912,N_3256,N_2546);
xnor U7913 (N_7913,N_1205,N_2288);
nor U7914 (N_7914,N_2471,N_4481);
and U7915 (N_7915,N_747,N_1619);
and U7916 (N_7916,N_4207,N_1147);
and U7917 (N_7917,N_311,N_2895);
and U7918 (N_7918,N_4957,N_3458);
nand U7919 (N_7919,N_811,N_877);
nand U7920 (N_7920,N_4707,N_3997);
or U7921 (N_7921,N_3756,N_161);
nand U7922 (N_7922,N_796,N_4490);
or U7923 (N_7923,N_3215,N_4579);
nor U7924 (N_7924,N_4436,N_3187);
nor U7925 (N_7925,N_3565,N_4453);
nor U7926 (N_7926,N_1423,N_3103);
and U7927 (N_7927,N_1783,N_3902);
and U7928 (N_7928,N_934,N_1662);
xnor U7929 (N_7929,N_1760,N_574);
and U7930 (N_7930,N_3598,N_3875);
or U7931 (N_7931,N_3462,N_3773);
or U7932 (N_7932,N_3670,N_4518);
nand U7933 (N_7933,N_4416,N_4135);
and U7934 (N_7934,N_2793,N_4513);
nor U7935 (N_7935,N_1408,N_447);
xnor U7936 (N_7936,N_876,N_1810);
or U7937 (N_7937,N_4190,N_2999);
or U7938 (N_7938,N_2389,N_2417);
nand U7939 (N_7939,N_2476,N_553);
xor U7940 (N_7940,N_2538,N_3354);
nor U7941 (N_7941,N_3638,N_2262);
xor U7942 (N_7942,N_2621,N_3936);
nand U7943 (N_7943,N_590,N_1467);
nor U7944 (N_7944,N_3607,N_3899);
xor U7945 (N_7945,N_4875,N_4694);
nor U7946 (N_7946,N_2829,N_2026);
nand U7947 (N_7947,N_4044,N_4185);
or U7948 (N_7948,N_27,N_548);
xnor U7949 (N_7949,N_1950,N_4649);
nor U7950 (N_7950,N_97,N_443);
nand U7951 (N_7951,N_3358,N_2713);
or U7952 (N_7952,N_3094,N_1862);
nor U7953 (N_7953,N_2609,N_2093);
nor U7954 (N_7954,N_1992,N_3971);
nor U7955 (N_7955,N_1586,N_1581);
or U7956 (N_7956,N_1746,N_1665);
and U7957 (N_7957,N_3100,N_4843);
or U7958 (N_7958,N_3984,N_4763);
or U7959 (N_7959,N_4825,N_2078);
or U7960 (N_7960,N_4041,N_3000);
and U7961 (N_7961,N_1563,N_2421);
xnor U7962 (N_7962,N_4877,N_4330);
or U7963 (N_7963,N_1392,N_4605);
nor U7964 (N_7964,N_4868,N_1762);
xnor U7965 (N_7965,N_3929,N_995);
and U7966 (N_7966,N_613,N_3632);
or U7967 (N_7967,N_3028,N_1188);
nand U7968 (N_7968,N_3469,N_1882);
or U7969 (N_7969,N_1938,N_488);
nor U7970 (N_7970,N_4879,N_1456);
nand U7971 (N_7971,N_248,N_4717);
nand U7972 (N_7972,N_4467,N_829);
and U7973 (N_7973,N_1882,N_1621);
nor U7974 (N_7974,N_3686,N_3075);
or U7975 (N_7975,N_14,N_2400);
xor U7976 (N_7976,N_2617,N_2101);
and U7977 (N_7977,N_3896,N_2714);
or U7978 (N_7978,N_3582,N_1709);
and U7979 (N_7979,N_4899,N_4627);
nand U7980 (N_7980,N_3324,N_3233);
nor U7981 (N_7981,N_749,N_3165);
and U7982 (N_7982,N_3844,N_3056);
nand U7983 (N_7983,N_4068,N_2858);
nor U7984 (N_7984,N_148,N_884);
or U7985 (N_7985,N_4852,N_1226);
and U7986 (N_7986,N_834,N_3545);
and U7987 (N_7987,N_829,N_4353);
nand U7988 (N_7988,N_3946,N_4780);
xor U7989 (N_7989,N_4762,N_464);
or U7990 (N_7990,N_4815,N_1986);
nor U7991 (N_7991,N_4704,N_2984);
nand U7992 (N_7992,N_4491,N_1506);
or U7993 (N_7993,N_3040,N_1230);
nand U7994 (N_7994,N_2358,N_4811);
nor U7995 (N_7995,N_48,N_4964);
and U7996 (N_7996,N_701,N_1984);
nand U7997 (N_7997,N_221,N_1654);
nand U7998 (N_7998,N_1687,N_657);
or U7999 (N_7999,N_510,N_3923);
xnor U8000 (N_8000,N_786,N_3148);
xnor U8001 (N_8001,N_3094,N_3220);
nor U8002 (N_8002,N_991,N_3977);
nor U8003 (N_8003,N_687,N_3104);
and U8004 (N_8004,N_1805,N_3555);
nor U8005 (N_8005,N_4863,N_4684);
or U8006 (N_8006,N_3129,N_491);
and U8007 (N_8007,N_3506,N_1513);
or U8008 (N_8008,N_4809,N_1405);
and U8009 (N_8009,N_2721,N_3806);
and U8010 (N_8010,N_223,N_2037);
xor U8011 (N_8011,N_2851,N_4980);
nor U8012 (N_8012,N_4763,N_2021);
nor U8013 (N_8013,N_512,N_2910);
nor U8014 (N_8014,N_1803,N_614);
xor U8015 (N_8015,N_3173,N_2784);
and U8016 (N_8016,N_3512,N_3105);
and U8017 (N_8017,N_2696,N_2612);
and U8018 (N_8018,N_3534,N_4111);
xor U8019 (N_8019,N_2186,N_4477);
nand U8020 (N_8020,N_1470,N_4588);
nor U8021 (N_8021,N_3379,N_1595);
xnor U8022 (N_8022,N_3124,N_3689);
nand U8023 (N_8023,N_4769,N_729);
nor U8024 (N_8024,N_1136,N_806);
and U8025 (N_8025,N_3764,N_3078);
xnor U8026 (N_8026,N_3829,N_2227);
xor U8027 (N_8027,N_1980,N_1373);
nand U8028 (N_8028,N_3340,N_2688);
and U8029 (N_8029,N_3029,N_4899);
or U8030 (N_8030,N_426,N_2322);
xnor U8031 (N_8031,N_4020,N_974);
and U8032 (N_8032,N_380,N_4491);
xor U8033 (N_8033,N_1068,N_4373);
nor U8034 (N_8034,N_602,N_2533);
nor U8035 (N_8035,N_243,N_3194);
or U8036 (N_8036,N_4223,N_4420);
nor U8037 (N_8037,N_756,N_3598);
nor U8038 (N_8038,N_475,N_1407);
and U8039 (N_8039,N_701,N_981);
or U8040 (N_8040,N_2098,N_1518);
or U8041 (N_8041,N_3241,N_2046);
nor U8042 (N_8042,N_1949,N_4635);
and U8043 (N_8043,N_3629,N_3025);
and U8044 (N_8044,N_907,N_3287);
xor U8045 (N_8045,N_4612,N_2318);
or U8046 (N_8046,N_3008,N_4987);
nor U8047 (N_8047,N_1372,N_4974);
nor U8048 (N_8048,N_1525,N_4135);
or U8049 (N_8049,N_3423,N_908);
and U8050 (N_8050,N_2289,N_3363);
xor U8051 (N_8051,N_1836,N_2205);
or U8052 (N_8052,N_2484,N_4373);
nand U8053 (N_8053,N_2398,N_4554);
nor U8054 (N_8054,N_557,N_4379);
xor U8055 (N_8055,N_1231,N_1919);
nand U8056 (N_8056,N_362,N_4169);
nand U8057 (N_8057,N_393,N_639);
xor U8058 (N_8058,N_3301,N_4022);
or U8059 (N_8059,N_3871,N_4453);
nor U8060 (N_8060,N_2576,N_4573);
nor U8061 (N_8061,N_1648,N_1464);
and U8062 (N_8062,N_1786,N_2828);
nand U8063 (N_8063,N_4073,N_3494);
or U8064 (N_8064,N_3519,N_2250);
xnor U8065 (N_8065,N_3711,N_3153);
or U8066 (N_8066,N_1216,N_958);
and U8067 (N_8067,N_2466,N_3479);
or U8068 (N_8068,N_1003,N_3073);
xnor U8069 (N_8069,N_4358,N_150);
and U8070 (N_8070,N_3331,N_3716);
nor U8071 (N_8071,N_3076,N_530);
xor U8072 (N_8072,N_631,N_1466);
and U8073 (N_8073,N_4284,N_2915);
or U8074 (N_8074,N_1637,N_4785);
xor U8075 (N_8075,N_1077,N_2724);
nor U8076 (N_8076,N_938,N_4045);
and U8077 (N_8077,N_990,N_2686);
xnor U8078 (N_8078,N_4020,N_2062);
or U8079 (N_8079,N_855,N_1900);
and U8080 (N_8080,N_3114,N_1380);
nor U8081 (N_8081,N_4364,N_3013);
and U8082 (N_8082,N_589,N_3020);
nand U8083 (N_8083,N_2594,N_2796);
or U8084 (N_8084,N_3134,N_4329);
nor U8085 (N_8085,N_1050,N_2594);
nor U8086 (N_8086,N_3911,N_804);
nand U8087 (N_8087,N_3133,N_3580);
nor U8088 (N_8088,N_4238,N_4594);
xnor U8089 (N_8089,N_2855,N_2167);
xnor U8090 (N_8090,N_4395,N_3206);
nor U8091 (N_8091,N_581,N_3753);
xor U8092 (N_8092,N_3263,N_1638);
nand U8093 (N_8093,N_4894,N_4049);
and U8094 (N_8094,N_1139,N_2489);
nor U8095 (N_8095,N_1054,N_1892);
xnor U8096 (N_8096,N_4985,N_2905);
or U8097 (N_8097,N_4744,N_3768);
nand U8098 (N_8098,N_836,N_3984);
or U8099 (N_8099,N_4012,N_4538);
or U8100 (N_8100,N_1233,N_3168);
nor U8101 (N_8101,N_4666,N_1847);
nor U8102 (N_8102,N_269,N_3781);
xor U8103 (N_8103,N_2672,N_208);
or U8104 (N_8104,N_1727,N_617);
nor U8105 (N_8105,N_2351,N_2908);
xnor U8106 (N_8106,N_3318,N_204);
nand U8107 (N_8107,N_394,N_16);
and U8108 (N_8108,N_826,N_3710);
and U8109 (N_8109,N_1754,N_562);
and U8110 (N_8110,N_1879,N_1938);
and U8111 (N_8111,N_2592,N_3885);
or U8112 (N_8112,N_2488,N_2974);
nor U8113 (N_8113,N_4749,N_1942);
nor U8114 (N_8114,N_2576,N_1270);
xor U8115 (N_8115,N_98,N_1918);
nand U8116 (N_8116,N_4806,N_1389);
xor U8117 (N_8117,N_4769,N_89);
xnor U8118 (N_8118,N_1360,N_3353);
nand U8119 (N_8119,N_2089,N_393);
and U8120 (N_8120,N_149,N_4627);
and U8121 (N_8121,N_2474,N_2080);
or U8122 (N_8122,N_262,N_4132);
nand U8123 (N_8123,N_4046,N_1051);
and U8124 (N_8124,N_2841,N_3028);
nor U8125 (N_8125,N_4785,N_3479);
or U8126 (N_8126,N_944,N_928);
nand U8127 (N_8127,N_2783,N_1977);
and U8128 (N_8128,N_1387,N_887);
nor U8129 (N_8129,N_1681,N_2537);
xnor U8130 (N_8130,N_1634,N_2988);
or U8131 (N_8131,N_3423,N_614);
xor U8132 (N_8132,N_4936,N_4545);
or U8133 (N_8133,N_2357,N_2386);
nor U8134 (N_8134,N_3299,N_2184);
nand U8135 (N_8135,N_1068,N_444);
and U8136 (N_8136,N_1648,N_1238);
xnor U8137 (N_8137,N_2321,N_2575);
and U8138 (N_8138,N_2622,N_701);
nand U8139 (N_8139,N_1388,N_4030);
and U8140 (N_8140,N_2747,N_4109);
xnor U8141 (N_8141,N_3443,N_4144);
and U8142 (N_8142,N_2627,N_3177);
xor U8143 (N_8143,N_4106,N_219);
nand U8144 (N_8144,N_136,N_2151);
xnor U8145 (N_8145,N_315,N_1382);
nor U8146 (N_8146,N_3455,N_4635);
nor U8147 (N_8147,N_3447,N_4189);
and U8148 (N_8148,N_3298,N_3337);
nor U8149 (N_8149,N_966,N_640);
nor U8150 (N_8150,N_3922,N_1298);
xnor U8151 (N_8151,N_1889,N_2663);
nand U8152 (N_8152,N_4681,N_2609);
or U8153 (N_8153,N_2110,N_2971);
and U8154 (N_8154,N_1829,N_4000);
or U8155 (N_8155,N_1522,N_159);
xor U8156 (N_8156,N_1130,N_2533);
or U8157 (N_8157,N_4581,N_138);
nand U8158 (N_8158,N_207,N_1300);
nand U8159 (N_8159,N_3245,N_3862);
nand U8160 (N_8160,N_4832,N_2815);
or U8161 (N_8161,N_992,N_1201);
and U8162 (N_8162,N_4527,N_4207);
or U8163 (N_8163,N_1264,N_4642);
or U8164 (N_8164,N_536,N_4142);
nor U8165 (N_8165,N_4772,N_2074);
nand U8166 (N_8166,N_4913,N_4180);
or U8167 (N_8167,N_4577,N_437);
nor U8168 (N_8168,N_1481,N_474);
nor U8169 (N_8169,N_2764,N_1306);
nand U8170 (N_8170,N_1858,N_4515);
and U8171 (N_8171,N_1934,N_4746);
nor U8172 (N_8172,N_1304,N_453);
and U8173 (N_8173,N_3895,N_2789);
nand U8174 (N_8174,N_3643,N_3939);
nor U8175 (N_8175,N_818,N_3164);
xor U8176 (N_8176,N_2818,N_3854);
or U8177 (N_8177,N_4919,N_4814);
nand U8178 (N_8178,N_1406,N_601);
or U8179 (N_8179,N_480,N_3090);
or U8180 (N_8180,N_4024,N_2949);
or U8181 (N_8181,N_3214,N_1014);
nor U8182 (N_8182,N_1593,N_1093);
nand U8183 (N_8183,N_3913,N_2679);
nor U8184 (N_8184,N_979,N_4878);
nand U8185 (N_8185,N_1107,N_1172);
nor U8186 (N_8186,N_2169,N_465);
nand U8187 (N_8187,N_4233,N_4048);
nand U8188 (N_8188,N_2176,N_3310);
xor U8189 (N_8189,N_3799,N_3825);
nand U8190 (N_8190,N_2951,N_265);
nand U8191 (N_8191,N_516,N_4421);
nor U8192 (N_8192,N_849,N_1522);
or U8193 (N_8193,N_2451,N_2057);
or U8194 (N_8194,N_4269,N_2620);
nor U8195 (N_8195,N_3938,N_2410);
xor U8196 (N_8196,N_3148,N_520);
and U8197 (N_8197,N_1193,N_355);
nor U8198 (N_8198,N_3207,N_3823);
and U8199 (N_8199,N_4739,N_3228);
nand U8200 (N_8200,N_4786,N_315);
nor U8201 (N_8201,N_1823,N_3392);
or U8202 (N_8202,N_2564,N_228);
xnor U8203 (N_8203,N_2737,N_3196);
nor U8204 (N_8204,N_1699,N_166);
and U8205 (N_8205,N_1412,N_2025);
nor U8206 (N_8206,N_125,N_2035);
and U8207 (N_8207,N_2640,N_4643);
xnor U8208 (N_8208,N_1454,N_265);
nor U8209 (N_8209,N_2713,N_631);
xnor U8210 (N_8210,N_1392,N_3220);
and U8211 (N_8211,N_933,N_4933);
or U8212 (N_8212,N_3492,N_45);
or U8213 (N_8213,N_1310,N_3708);
nor U8214 (N_8214,N_1513,N_1238);
nand U8215 (N_8215,N_4448,N_2268);
xnor U8216 (N_8216,N_996,N_4921);
xnor U8217 (N_8217,N_3369,N_105);
nor U8218 (N_8218,N_3424,N_696);
or U8219 (N_8219,N_2986,N_1355);
and U8220 (N_8220,N_2037,N_4499);
nor U8221 (N_8221,N_4302,N_4399);
nand U8222 (N_8222,N_985,N_3636);
and U8223 (N_8223,N_4391,N_3228);
nand U8224 (N_8224,N_2318,N_2344);
and U8225 (N_8225,N_4968,N_2866);
and U8226 (N_8226,N_4020,N_4337);
xnor U8227 (N_8227,N_1088,N_2711);
or U8228 (N_8228,N_1049,N_735);
or U8229 (N_8229,N_4686,N_2702);
xnor U8230 (N_8230,N_355,N_178);
or U8231 (N_8231,N_214,N_4891);
or U8232 (N_8232,N_1043,N_2932);
nand U8233 (N_8233,N_2709,N_3754);
xnor U8234 (N_8234,N_455,N_2457);
or U8235 (N_8235,N_306,N_304);
nand U8236 (N_8236,N_1664,N_3261);
nor U8237 (N_8237,N_3484,N_1512);
nor U8238 (N_8238,N_722,N_3056);
and U8239 (N_8239,N_4758,N_4059);
nand U8240 (N_8240,N_990,N_111);
nor U8241 (N_8241,N_3047,N_3321);
nand U8242 (N_8242,N_1928,N_4388);
or U8243 (N_8243,N_2575,N_499);
nand U8244 (N_8244,N_1168,N_2264);
nand U8245 (N_8245,N_2987,N_1626);
nor U8246 (N_8246,N_3010,N_224);
xnor U8247 (N_8247,N_3324,N_3294);
and U8248 (N_8248,N_602,N_2715);
nand U8249 (N_8249,N_1750,N_1676);
nand U8250 (N_8250,N_689,N_2690);
nor U8251 (N_8251,N_2903,N_405);
nand U8252 (N_8252,N_2065,N_2044);
or U8253 (N_8253,N_4005,N_1694);
or U8254 (N_8254,N_146,N_1115);
xor U8255 (N_8255,N_2699,N_4019);
and U8256 (N_8256,N_2537,N_4240);
or U8257 (N_8257,N_1142,N_733);
nor U8258 (N_8258,N_3954,N_3125);
xor U8259 (N_8259,N_1636,N_657);
nor U8260 (N_8260,N_3223,N_825);
or U8261 (N_8261,N_398,N_501);
or U8262 (N_8262,N_2911,N_250);
and U8263 (N_8263,N_2186,N_122);
or U8264 (N_8264,N_2685,N_4779);
and U8265 (N_8265,N_698,N_710);
nand U8266 (N_8266,N_4309,N_3683);
or U8267 (N_8267,N_783,N_1093);
and U8268 (N_8268,N_1463,N_2291);
and U8269 (N_8269,N_826,N_2373);
or U8270 (N_8270,N_617,N_1691);
or U8271 (N_8271,N_1537,N_3644);
nand U8272 (N_8272,N_4853,N_3506);
or U8273 (N_8273,N_4028,N_865);
nor U8274 (N_8274,N_1352,N_3276);
and U8275 (N_8275,N_4020,N_771);
or U8276 (N_8276,N_1127,N_2726);
xnor U8277 (N_8277,N_4577,N_3983);
or U8278 (N_8278,N_3734,N_4853);
xnor U8279 (N_8279,N_4108,N_3223);
or U8280 (N_8280,N_4415,N_1598);
nand U8281 (N_8281,N_1176,N_4091);
and U8282 (N_8282,N_1048,N_436);
and U8283 (N_8283,N_406,N_858);
or U8284 (N_8284,N_4480,N_4743);
or U8285 (N_8285,N_66,N_3512);
or U8286 (N_8286,N_4312,N_4120);
xor U8287 (N_8287,N_4753,N_2673);
or U8288 (N_8288,N_1118,N_1126);
xor U8289 (N_8289,N_674,N_2116);
nor U8290 (N_8290,N_418,N_2804);
nor U8291 (N_8291,N_4368,N_1920);
and U8292 (N_8292,N_477,N_1610);
nand U8293 (N_8293,N_1379,N_3866);
nand U8294 (N_8294,N_512,N_1280);
or U8295 (N_8295,N_1748,N_2936);
or U8296 (N_8296,N_1494,N_1107);
nor U8297 (N_8297,N_1949,N_2142);
or U8298 (N_8298,N_3247,N_4489);
or U8299 (N_8299,N_4381,N_2427);
and U8300 (N_8300,N_630,N_1918);
xor U8301 (N_8301,N_931,N_3784);
nand U8302 (N_8302,N_4093,N_3167);
nor U8303 (N_8303,N_1921,N_4186);
nor U8304 (N_8304,N_3674,N_974);
and U8305 (N_8305,N_1072,N_4991);
nand U8306 (N_8306,N_1772,N_1472);
or U8307 (N_8307,N_2877,N_4708);
nand U8308 (N_8308,N_1710,N_1516);
or U8309 (N_8309,N_2055,N_1405);
nand U8310 (N_8310,N_4545,N_1510);
xnor U8311 (N_8311,N_2041,N_1483);
or U8312 (N_8312,N_2766,N_1623);
nor U8313 (N_8313,N_3032,N_4908);
nor U8314 (N_8314,N_4158,N_2795);
nand U8315 (N_8315,N_3250,N_2679);
nand U8316 (N_8316,N_2206,N_4884);
nor U8317 (N_8317,N_4919,N_3919);
nand U8318 (N_8318,N_2439,N_2427);
and U8319 (N_8319,N_1443,N_4615);
and U8320 (N_8320,N_2861,N_512);
nor U8321 (N_8321,N_2790,N_1451);
and U8322 (N_8322,N_3735,N_3267);
and U8323 (N_8323,N_2626,N_409);
nor U8324 (N_8324,N_36,N_2119);
xor U8325 (N_8325,N_1387,N_4147);
and U8326 (N_8326,N_3418,N_2324);
and U8327 (N_8327,N_1715,N_2043);
or U8328 (N_8328,N_775,N_2615);
or U8329 (N_8329,N_3311,N_2148);
nand U8330 (N_8330,N_881,N_4011);
and U8331 (N_8331,N_2759,N_4892);
and U8332 (N_8332,N_931,N_1033);
nor U8333 (N_8333,N_4064,N_2653);
nand U8334 (N_8334,N_1315,N_3412);
nand U8335 (N_8335,N_3165,N_2871);
and U8336 (N_8336,N_685,N_1218);
xor U8337 (N_8337,N_2275,N_537);
nor U8338 (N_8338,N_1105,N_2395);
or U8339 (N_8339,N_0,N_3623);
xnor U8340 (N_8340,N_4887,N_3895);
nand U8341 (N_8341,N_906,N_3165);
or U8342 (N_8342,N_3275,N_4184);
or U8343 (N_8343,N_1046,N_4701);
nand U8344 (N_8344,N_1649,N_4526);
nor U8345 (N_8345,N_539,N_4252);
nand U8346 (N_8346,N_4652,N_3149);
and U8347 (N_8347,N_146,N_4243);
nand U8348 (N_8348,N_3083,N_4846);
nand U8349 (N_8349,N_1259,N_2436);
xnor U8350 (N_8350,N_3311,N_3875);
or U8351 (N_8351,N_3230,N_2418);
nand U8352 (N_8352,N_2844,N_1598);
xnor U8353 (N_8353,N_3495,N_2804);
xor U8354 (N_8354,N_1557,N_1565);
nor U8355 (N_8355,N_4229,N_3089);
nor U8356 (N_8356,N_4309,N_2243);
xor U8357 (N_8357,N_807,N_4996);
or U8358 (N_8358,N_823,N_3063);
or U8359 (N_8359,N_1698,N_591);
xor U8360 (N_8360,N_2155,N_4973);
nand U8361 (N_8361,N_2012,N_1615);
nor U8362 (N_8362,N_2692,N_4643);
nor U8363 (N_8363,N_3966,N_2078);
nand U8364 (N_8364,N_2947,N_4934);
or U8365 (N_8365,N_1352,N_186);
nor U8366 (N_8366,N_18,N_3464);
and U8367 (N_8367,N_3600,N_4886);
and U8368 (N_8368,N_3559,N_4261);
nand U8369 (N_8369,N_4438,N_586);
and U8370 (N_8370,N_2236,N_4183);
nor U8371 (N_8371,N_522,N_3307);
xnor U8372 (N_8372,N_908,N_3872);
or U8373 (N_8373,N_4712,N_4200);
xor U8374 (N_8374,N_1654,N_731);
and U8375 (N_8375,N_856,N_4751);
or U8376 (N_8376,N_1752,N_1093);
and U8377 (N_8377,N_4616,N_3277);
and U8378 (N_8378,N_3966,N_985);
or U8379 (N_8379,N_4864,N_2635);
xor U8380 (N_8380,N_3640,N_1227);
nand U8381 (N_8381,N_3301,N_3719);
nor U8382 (N_8382,N_1638,N_406);
nand U8383 (N_8383,N_210,N_4207);
xnor U8384 (N_8384,N_4457,N_1631);
or U8385 (N_8385,N_3514,N_2818);
xor U8386 (N_8386,N_1886,N_2278);
xor U8387 (N_8387,N_2514,N_2623);
or U8388 (N_8388,N_1730,N_3878);
nand U8389 (N_8389,N_1525,N_3547);
and U8390 (N_8390,N_4149,N_1714);
nor U8391 (N_8391,N_3394,N_3636);
nor U8392 (N_8392,N_4528,N_4636);
xor U8393 (N_8393,N_2888,N_401);
or U8394 (N_8394,N_2383,N_157);
nand U8395 (N_8395,N_3251,N_1468);
nor U8396 (N_8396,N_2548,N_4919);
nand U8397 (N_8397,N_1169,N_1963);
and U8398 (N_8398,N_2599,N_1359);
xnor U8399 (N_8399,N_1127,N_1815);
or U8400 (N_8400,N_3668,N_1128);
nand U8401 (N_8401,N_4077,N_4436);
xor U8402 (N_8402,N_614,N_320);
and U8403 (N_8403,N_3003,N_1255);
nand U8404 (N_8404,N_2739,N_4648);
xnor U8405 (N_8405,N_3104,N_2525);
nor U8406 (N_8406,N_3457,N_944);
and U8407 (N_8407,N_917,N_3493);
nand U8408 (N_8408,N_2720,N_1943);
nor U8409 (N_8409,N_3935,N_4341);
nor U8410 (N_8410,N_977,N_203);
nand U8411 (N_8411,N_248,N_4368);
and U8412 (N_8412,N_3494,N_272);
nor U8413 (N_8413,N_4164,N_732);
nand U8414 (N_8414,N_4774,N_3420);
nor U8415 (N_8415,N_3211,N_3210);
nor U8416 (N_8416,N_3953,N_4429);
and U8417 (N_8417,N_627,N_707);
xor U8418 (N_8418,N_4313,N_694);
nand U8419 (N_8419,N_2706,N_2713);
or U8420 (N_8420,N_3521,N_4865);
and U8421 (N_8421,N_4292,N_3833);
nor U8422 (N_8422,N_3670,N_913);
nand U8423 (N_8423,N_3925,N_4280);
nor U8424 (N_8424,N_3887,N_1079);
nand U8425 (N_8425,N_2988,N_133);
and U8426 (N_8426,N_4025,N_4228);
nor U8427 (N_8427,N_1422,N_4341);
xor U8428 (N_8428,N_4856,N_2715);
nand U8429 (N_8429,N_1109,N_3430);
xor U8430 (N_8430,N_4328,N_2729);
nand U8431 (N_8431,N_2471,N_3868);
and U8432 (N_8432,N_1628,N_3739);
or U8433 (N_8433,N_3902,N_900);
xor U8434 (N_8434,N_1354,N_3780);
nor U8435 (N_8435,N_4750,N_467);
and U8436 (N_8436,N_1686,N_2592);
or U8437 (N_8437,N_4446,N_1578);
nand U8438 (N_8438,N_3122,N_2288);
nor U8439 (N_8439,N_3315,N_245);
or U8440 (N_8440,N_2228,N_1579);
xnor U8441 (N_8441,N_4890,N_3200);
nor U8442 (N_8442,N_1798,N_11);
nand U8443 (N_8443,N_990,N_1103);
or U8444 (N_8444,N_4628,N_4366);
or U8445 (N_8445,N_4913,N_3700);
and U8446 (N_8446,N_1024,N_157);
nor U8447 (N_8447,N_735,N_4799);
nand U8448 (N_8448,N_4738,N_3409);
or U8449 (N_8449,N_1459,N_4331);
or U8450 (N_8450,N_1156,N_4847);
or U8451 (N_8451,N_1168,N_4540);
and U8452 (N_8452,N_995,N_1833);
xnor U8453 (N_8453,N_698,N_4834);
nor U8454 (N_8454,N_1627,N_3117);
and U8455 (N_8455,N_426,N_2971);
and U8456 (N_8456,N_2084,N_1039);
or U8457 (N_8457,N_2814,N_2465);
nor U8458 (N_8458,N_3533,N_2696);
and U8459 (N_8459,N_4567,N_2774);
xnor U8460 (N_8460,N_4647,N_1271);
nor U8461 (N_8461,N_166,N_4217);
xnor U8462 (N_8462,N_3270,N_2350);
nor U8463 (N_8463,N_2919,N_2904);
nor U8464 (N_8464,N_181,N_1615);
or U8465 (N_8465,N_952,N_3429);
and U8466 (N_8466,N_3280,N_4053);
nand U8467 (N_8467,N_1130,N_1533);
xnor U8468 (N_8468,N_1227,N_1842);
and U8469 (N_8469,N_1674,N_3773);
nand U8470 (N_8470,N_717,N_1096);
nand U8471 (N_8471,N_2741,N_1001);
nand U8472 (N_8472,N_3588,N_341);
nand U8473 (N_8473,N_1013,N_1393);
xor U8474 (N_8474,N_4625,N_3574);
nand U8475 (N_8475,N_3863,N_3443);
or U8476 (N_8476,N_4941,N_2107);
xor U8477 (N_8477,N_3426,N_2177);
and U8478 (N_8478,N_2274,N_1424);
and U8479 (N_8479,N_4009,N_1054);
nand U8480 (N_8480,N_4063,N_1696);
nand U8481 (N_8481,N_2557,N_2786);
or U8482 (N_8482,N_697,N_2365);
nand U8483 (N_8483,N_1374,N_3516);
nor U8484 (N_8484,N_3447,N_177);
nand U8485 (N_8485,N_3405,N_2413);
xnor U8486 (N_8486,N_4121,N_1017);
nor U8487 (N_8487,N_193,N_3938);
nand U8488 (N_8488,N_3848,N_753);
nand U8489 (N_8489,N_2575,N_4065);
and U8490 (N_8490,N_2274,N_2117);
nand U8491 (N_8491,N_1951,N_3341);
or U8492 (N_8492,N_4570,N_1382);
xor U8493 (N_8493,N_3454,N_3349);
nand U8494 (N_8494,N_468,N_1403);
nand U8495 (N_8495,N_1809,N_1365);
and U8496 (N_8496,N_1334,N_1224);
xor U8497 (N_8497,N_2654,N_2660);
nor U8498 (N_8498,N_2685,N_3648);
and U8499 (N_8499,N_3909,N_539);
or U8500 (N_8500,N_87,N_20);
or U8501 (N_8501,N_4263,N_1588);
nand U8502 (N_8502,N_2206,N_3126);
or U8503 (N_8503,N_2107,N_1882);
nand U8504 (N_8504,N_1606,N_4633);
and U8505 (N_8505,N_1655,N_4154);
xor U8506 (N_8506,N_3931,N_3768);
or U8507 (N_8507,N_635,N_100);
or U8508 (N_8508,N_1434,N_3171);
nor U8509 (N_8509,N_2381,N_3203);
xnor U8510 (N_8510,N_974,N_4447);
or U8511 (N_8511,N_4600,N_1502);
nand U8512 (N_8512,N_4265,N_1989);
or U8513 (N_8513,N_2387,N_762);
nor U8514 (N_8514,N_185,N_3531);
nor U8515 (N_8515,N_4990,N_846);
nand U8516 (N_8516,N_3193,N_2528);
nor U8517 (N_8517,N_3914,N_1747);
nor U8518 (N_8518,N_4718,N_3420);
and U8519 (N_8519,N_4091,N_1220);
xnor U8520 (N_8520,N_2114,N_2541);
or U8521 (N_8521,N_3087,N_692);
xor U8522 (N_8522,N_45,N_2244);
nor U8523 (N_8523,N_1011,N_368);
nor U8524 (N_8524,N_3837,N_4223);
xnor U8525 (N_8525,N_71,N_2324);
nor U8526 (N_8526,N_3096,N_4938);
nand U8527 (N_8527,N_4489,N_3845);
xor U8528 (N_8528,N_693,N_446);
nor U8529 (N_8529,N_1991,N_1537);
xnor U8530 (N_8530,N_3277,N_643);
nor U8531 (N_8531,N_4803,N_918);
and U8532 (N_8532,N_1135,N_3600);
or U8533 (N_8533,N_3914,N_4971);
nor U8534 (N_8534,N_2268,N_1401);
nand U8535 (N_8535,N_3854,N_629);
xor U8536 (N_8536,N_4327,N_2157);
xnor U8537 (N_8537,N_3933,N_1988);
and U8538 (N_8538,N_2232,N_1063);
or U8539 (N_8539,N_4391,N_1133);
nor U8540 (N_8540,N_1931,N_3173);
and U8541 (N_8541,N_4930,N_1846);
nand U8542 (N_8542,N_915,N_2978);
or U8543 (N_8543,N_2600,N_1867);
xor U8544 (N_8544,N_3867,N_4425);
nand U8545 (N_8545,N_947,N_124);
or U8546 (N_8546,N_2100,N_742);
and U8547 (N_8547,N_1634,N_1632);
nand U8548 (N_8548,N_1094,N_2007);
nor U8549 (N_8549,N_4116,N_1399);
nor U8550 (N_8550,N_3056,N_1140);
xnor U8551 (N_8551,N_2336,N_2735);
nor U8552 (N_8552,N_2042,N_910);
nor U8553 (N_8553,N_430,N_192);
nand U8554 (N_8554,N_4109,N_2224);
nor U8555 (N_8555,N_3916,N_3246);
and U8556 (N_8556,N_63,N_4798);
xnor U8557 (N_8557,N_1087,N_3201);
nand U8558 (N_8558,N_1771,N_2167);
or U8559 (N_8559,N_416,N_2645);
nor U8560 (N_8560,N_2596,N_3625);
and U8561 (N_8561,N_218,N_4318);
nand U8562 (N_8562,N_98,N_4347);
nor U8563 (N_8563,N_2444,N_860);
and U8564 (N_8564,N_4323,N_4523);
nand U8565 (N_8565,N_3474,N_3762);
nand U8566 (N_8566,N_4492,N_1976);
nand U8567 (N_8567,N_2913,N_479);
or U8568 (N_8568,N_4393,N_340);
xnor U8569 (N_8569,N_1130,N_2359);
and U8570 (N_8570,N_3060,N_4399);
nand U8571 (N_8571,N_586,N_1547);
nor U8572 (N_8572,N_665,N_354);
xor U8573 (N_8573,N_11,N_1007);
nor U8574 (N_8574,N_2223,N_489);
and U8575 (N_8575,N_2899,N_4985);
nor U8576 (N_8576,N_4483,N_4507);
xnor U8577 (N_8577,N_2302,N_2338);
or U8578 (N_8578,N_4918,N_2946);
nand U8579 (N_8579,N_3859,N_429);
or U8580 (N_8580,N_1849,N_2076);
and U8581 (N_8581,N_1709,N_3237);
nor U8582 (N_8582,N_853,N_3177);
nor U8583 (N_8583,N_4702,N_2815);
nor U8584 (N_8584,N_1337,N_2347);
nand U8585 (N_8585,N_3100,N_3954);
nor U8586 (N_8586,N_1863,N_720);
or U8587 (N_8587,N_4699,N_2932);
and U8588 (N_8588,N_4505,N_4786);
or U8589 (N_8589,N_1658,N_4608);
xnor U8590 (N_8590,N_4841,N_2227);
xnor U8591 (N_8591,N_2455,N_942);
nor U8592 (N_8592,N_4968,N_1404);
xnor U8593 (N_8593,N_486,N_4656);
and U8594 (N_8594,N_2111,N_870);
nor U8595 (N_8595,N_1108,N_1961);
nor U8596 (N_8596,N_197,N_243);
and U8597 (N_8597,N_4437,N_3358);
nor U8598 (N_8598,N_1650,N_3413);
nand U8599 (N_8599,N_573,N_133);
xnor U8600 (N_8600,N_2170,N_437);
and U8601 (N_8601,N_4094,N_3653);
xor U8602 (N_8602,N_2259,N_3187);
and U8603 (N_8603,N_4541,N_2917);
nor U8604 (N_8604,N_4029,N_2022);
and U8605 (N_8605,N_3644,N_4150);
or U8606 (N_8606,N_3358,N_1266);
nor U8607 (N_8607,N_3791,N_3512);
or U8608 (N_8608,N_4785,N_4086);
and U8609 (N_8609,N_186,N_2686);
or U8610 (N_8610,N_2596,N_2707);
or U8611 (N_8611,N_4452,N_1834);
nor U8612 (N_8612,N_79,N_4924);
or U8613 (N_8613,N_1163,N_2058);
nand U8614 (N_8614,N_1458,N_4596);
and U8615 (N_8615,N_1297,N_3929);
nor U8616 (N_8616,N_2060,N_2741);
nor U8617 (N_8617,N_1051,N_3791);
xor U8618 (N_8618,N_294,N_4730);
nor U8619 (N_8619,N_3336,N_4607);
nand U8620 (N_8620,N_4577,N_2565);
nand U8621 (N_8621,N_3087,N_3091);
or U8622 (N_8622,N_2044,N_3190);
and U8623 (N_8623,N_3218,N_4473);
xnor U8624 (N_8624,N_2158,N_3095);
and U8625 (N_8625,N_3941,N_3421);
nor U8626 (N_8626,N_875,N_4818);
xnor U8627 (N_8627,N_1316,N_2542);
xor U8628 (N_8628,N_1464,N_2334);
nor U8629 (N_8629,N_347,N_4316);
xor U8630 (N_8630,N_1939,N_4912);
xnor U8631 (N_8631,N_1173,N_3754);
xnor U8632 (N_8632,N_309,N_2448);
nand U8633 (N_8633,N_972,N_3125);
xor U8634 (N_8634,N_872,N_4143);
xor U8635 (N_8635,N_661,N_3648);
and U8636 (N_8636,N_108,N_3314);
and U8637 (N_8637,N_528,N_1434);
nand U8638 (N_8638,N_2231,N_4196);
nand U8639 (N_8639,N_2459,N_2738);
xor U8640 (N_8640,N_2809,N_3033);
or U8641 (N_8641,N_4218,N_2892);
nor U8642 (N_8642,N_3638,N_3950);
nand U8643 (N_8643,N_781,N_1981);
or U8644 (N_8644,N_4807,N_2720);
and U8645 (N_8645,N_171,N_273);
and U8646 (N_8646,N_2880,N_1750);
nor U8647 (N_8647,N_2626,N_363);
or U8648 (N_8648,N_2565,N_2229);
xor U8649 (N_8649,N_4103,N_3086);
nor U8650 (N_8650,N_1259,N_2705);
nor U8651 (N_8651,N_1259,N_794);
nand U8652 (N_8652,N_4000,N_3739);
and U8653 (N_8653,N_1049,N_4926);
nand U8654 (N_8654,N_3672,N_194);
and U8655 (N_8655,N_3533,N_2543);
xnor U8656 (N_8656,N_4852,N_529);
and U8657 (N_8657,N_1156,N_1789);
nor U8658 (N_8658,N_3598,N_3077);
nand U8659 (N_8659,N_434,N_3604);
nand U8660 (N_8660,N_417,N_3130);
or U8661 (N_8661,N_1425,N_959);
and U8662 (N_8662,N_1697,N_2055);
and U8663 (N_8663,N_2968,N_3932);
xor U8664 (N_8664,N_4302,N_3291);
xor U8665 (N_8665,N_2530,N_1813);
and U8666 (N_8666,N_1687,N_3737);
xnor U8667 (N_8667,N_1191,N_962);
xor U8668 (N_8668,N_2751,N_147);
xor U8669 (N_8669,N_1161,N_3084);
nor U8670 (N_8670,N_3645,N_3338);
nand U8671 (N_8671,N_3029,N_2880);
nand U8672 (N_8672,N_3566,N_1769);
nor U8673 (N_8673,N_4331,N_2839);
xor U8674 (N_8674,N_3823,N_930);
and U8675 (N_8675,N_3176,N_4959);
nor U8676 (N_8676,N_2213,N_2126);
nor U8677 (N_8677,N_2773,N_806);
or U8678 (N_8678,N_3440,N_402);
xnor U8679 (N_8679,N_2758,N_210);
and U8680 (N_8680,N_474,N_1751);
or U8681 (N_8681,N_919,N_4354);
and U8682 (N_8682,N_1914,N_669);
nand U8683 (N_8683,N_4754,N_1366);
nand U8684 (N_8684,N_4317,N_870);
or U8685 (N_8685,N_2501,N_3524);
nand U8686 (N_8686,N_4164,N_2849);
xor U8687 (N_8687,N_4075,N_1598);
or U8688 (N_8688,N_3195,N_3164);
and U8689 (N_8689,N_1869,N_4137);
xor U8690 (N_8690,N_4646,N_733);
and U8691 (N_8691,N_1256,N_3355);
nand U8692 (N_8692,N_4461,N_3388);
xor U8693 (N_8693,N_4778,N_3690);
or U8694 (N_8694,N_1993,N_2605);
nor U8695 (N_8695,N_4627,N_2206);
xor U8696 (N_8696,N_3024,N_2625);
nor U8697 (N_8697,N_4049,N_2693);
xnor U8698 (N_8698,N_2092,N_4105);
xor U8699 (N_8699,N_1801,N_3975);
and U8700 (N_8700,N_1182,N_1100);
or U8701 (N_8701,N_3543,N_1749);
and U8702 (N_8702,N_732,N_2483);
nor U8703 (N_8703,N_4255,N_293);
nor U8704 (N_8704,N_1181,N_1369);
or U8705 (N_8705,N_1742,N_3443);
or U8706 (N_8706,N_2520,N_3653);
or U8707 (N_8707,N_390,N_4832);
xnor U8708 (N_8708,N_3328,N_2738);
nand U8709 (N_8709,N_961,N_4234);
or U8710 (N_8710,N_3217,N_3962);
xor U8711 (N_8711,N_1575,N_1782);
nand U8712 (N_8712,N_996,N_3304);
xor U8713 (N_8713,N_1671,N_2867);
nand U8714 (N_8714,N_403,N_2514);
or U8715 (N_8715,N_3686,N_1822);
xor U8716 (N_8716,N_4926,N_1487);
xor U8717 (N_8717,N_2400,N_4975);
nor U8718 (N_8718,N_3653,N_1192);
xnor U8719 (N_8719,N_3131,N_1590);
nor U8720 (N_8720,N_1537,N_2205);
xnor U8721 (N_8721,N_4694,N_993);
nand U8722 (N_8722,N_4759,N_3029);
nand U8723 (N_8723,N_4916,N_4650);
and U8724 (N_8724,N_4563,N_496);
or U8725 (N_8725,N_3176,N_1043);
nor U8726 (N_8726,N_1506,N_1787);
nand U8727 (N_8727,N_630,N_1130);
or U8728 (N_8728,N_894,N_4316);
or U8729 (N_8729,N_2255,N_3522);
or U8730 (N_8730,N_3231,N_2473);
nand U8731 (N_8731,N_4255,N_1002);
xor U8732 (N_8732,N_3625,N_735);
or U8733 (N_8733,N_3133,N_3130);
and U8734 (N_8734,N_728,N_2908);
xor U8735 (N_8735,N_2209,N_940);
and U8736 (N_8736,N_4424,N_2329);
and U8737 (N_8737,N_4672,N_1588);
xor U8738 (N_8738,N_4831,N_1596);
nand U8739 (N_8739,N_668,N_4627);
or U8740 (N_8740,N_1485,N_2344);
and U8741 (N_8741,N_695,N_4356);
nor U8742 (N_8742,N_2845,N_3239);
or U8743 (N_8743,N_2170,N_3317);
nand U8744 (N_8744,N_696,N_4876);
xor U8745 (N_8745,N_2355,N_204);
nor U8746 (N_8746,N_2546,N_1223);
nor U8747 (N_8747,N_1060,N_3611);
or U8748 (N_8748,N_2738,N_2713);
nor U8749 (N_8749,N_2405,N_2090);
xor U8750 (N_8750,N_1957,N_3614);
and U8751 (N_8751,N_2563,N_802);
nor U8752 (N_8752,N_4185,N_1877);
xor U8753 (N_8753,N_33,N_2074);
nand U8754 (N_8754,N_640,N_4454);
or U8755 (N_8755,N_4822,N_224);
nand U8756 (N_8756,N_1896,N_253);
nand U8757 (N_8757,N_3290,N_1118);
or U8758 (N_8758,N_1844,N_3511);
and U8759 (N_8759,N_2519,N_2884);
xnor U8760 (N_8760,N_358,N_3175);
nand U8761 (N_8761,N_2813,N_2507);
nor U8762 (N_8762,N_2994,N_1781);
or U8763 (N_8763,N_2537,N_1089);
nor U8764 (N_8764,N_4246,N_829);
xnor U8765 (N_8765,N_2381,N_4815);
nand U8766 (N_8766,N_4941,N_4817);
nand U8767 (N_8767,N_1302,N_541);
nor U8768 (N_8768,N_1349,N_3363);
nand U8769 (N_8769,N_3855,N_4492);
nand U8770 (N_8770,N_4049,N_2519);
nand U8771 (N_8771,N_550,N_854);
xor U8772 (N_8772,N_2525,N_4094);
nor U8773 (N_8773,N_3530,N_1340);
xnor U8774 (N_8774,N_1650,N_359);
or U8775 (N_8775,N_3976,N_3324);
xor U8776 (N_8776,N_3208,N_67);
and U8777 (N_8777,N_4809,N_2076);
nor U8778 (N_8778,N_1256,N_1193);
or U8779 (N_8779,N_2630,N_1809);
xor U8780 (N_8780,N_3749,N_2484);
and U8781 (N_8781,N_1963,N_1143);
and U8782 (N_8782,N_2068,N_2029);
nand U8783 (N_8783,N_3467,N_1041);
xnor U8784 (N_8784,N_2604,N_290);
nand U8785 (N_8785,N_2863,N_672);
and U8786 (N_8786,N_3253,N_4883);
or U8787 (N_8787,N_1705,N_120);
nor U8788 (N_8788,N_386,N_2908);
and U8789 (N_8789,N_3569,N_4989);
and U8790 (N_8790,N_2993,N_4531);
xor U8791 (N_8791,N_238,N_2176);
or U8792 (N_8792,N_60,N_945);
nand U8793 (N_8793,N_4223,N_1604);
nor U8794 (N_8794,N_4444,N_4429);
and U8795 (N_8795,N_889,N_3652);
nor U8796 (N_8796,N_3205,N_891);
nand U8797 (N_8797,N_2221,N_545);
nand U8798 (N_8798,N_759,N_4181);
or U8799 (N_8799,N_4047,N_2192);
nor U8800 (N_8800,N_352,N_1798);
and U8801 (N_8801,N_1485,N_3634);
nor U8802 (N_8802,N_1541,N_178);
and U8803 (N_8803,N_4143,N_4102);
xor U8804 (N_8804,N_2656,N_565);
xor U8805 (N_8805,N_4005,N_3620);
and U8806 (N_8806,N_2226,N_4623);
nand U8807 (N_8807,N_2598,N_3263);
nor U8808 (N_8808,N_4612,N_3624);
or U8809 (N_8809,N_1199,N_4046);
nand U8810 (N_8810,N_3515,N_2469);
xnor U8811 (N_8811,N_1573,N_3078);
nand U8812 (N_8812,N_1177,N_967);
and U8813 (N_8813,N_1218,N_714);
nand U8814 (N_8814,N_2868,N_3600);
nand U8815 (N_8815,N_4024,N_1121);
nand U8816 (N_8816,N_1869,N_4925);
and U8817 (N_8817,N_579,N_4491);
nand U8818 (N_8818,N_430,N_4534);
nand U8819 (N_8819,N_1654,N_4891);
or U8820 (N_8820,N_3768,N_1968);
or U8821 (N_8821,N_707,N_3813);
nand U8822 (N_8822,N_456,N_3135);
or U8823 (N_8823,N_1594,N_4821);
nor U8824 (N_8824,N_3464,N_3170);
and U8825 (N_8825,N_1001,N_2076);
and U8826 (N_8826,N_2376,N_2681);
nand U8827 (N_8827,N_259,N_3057);
xnor U8828 (N_8828,N_752,N_682);
and U8829 (N_8829,N_2471,N_55);
xnor U8830 (N_8830,N_4042,N_2453);
or U8831 (N_8831,N_2068,N_4478);
and U8832 (N_8832,N_2547,N_2618);
nor U8833 (N_8833,N_2015,N_3531);
nor U8834 (N_8834,N_2717,N_10);
nand U8835 (N_8835,N_1514,N_1167);
nor U8836 (N_8836,N_3766,N_2503);
xnor U8837 (N_8837,N_2596,N_3921);
nor U8838 (N_8838,N_4497,N_3832);
and U8839 (N_8839,N_1422,N_2641);
nand U8840 (N_8840,N_3534,N_4366);
xnor U8841 (N_8841,N_689,N_2619);
or U8842 (N_8842,N_2420,N_4034);
xor U8843 (N_8843,N_4729,N_1316);
xnor U8844 (N_8844,N_49,N_2054);
nand U8845 (N_8845,N_1990,N_1306);
nand U8846 (N_8846,N_3563,N_2862);
xor U8847 (N_8847,N_3170,N_170);
or U8848 (N_8848,N_1193,N_1843);
or U8849 (N_8849,N_4173,N_4634);
or U8850 (N_8850,N_4447,N_3721);
nand U8851 (N_8851,N_649,N_1144);
xor U8852 (N_8852,N_3607,N_2195);
or U8853 (N_8853,N_572,N_4085);
xor U8854 (N_8854,N_4958,N_111);
xor U8855 (N_8855,N_2686,N_342);
and U8856 (N_8856,N_730,N_4254);
and U8857 (N_8857,N_2684,N_362);
and U8858 (N_8858,N_3259,N_356);
or U8859 (N_8859,N_3887,N_113);
and U8860 (N_8860,N_3336,N_296);
or U8861 (N_8861,N_3519,N_3944);
or U8862 (N_8862,N_2712,N_2297);
xor U8863 (N_8863,N_3625,N_834);
nand U8864 (N_8864,N_2432,N_257);
or U8865 (N_8865,N_3651,N_2619);
xor U8866 (N_8866,N_629,N_2063);
or U8867 (N_8867,N_2548,N_3861);
or U8868 (N_8868,N_2488,N_4563);
nand U8869 (N_8869,N_2405,N_1927);
xnor U8870 (N_8870,N_2757,N_934);
xor U8871 (N_8871,N_3849,N_3333);
xnor U8872 (N_8872,N_126,N_136);
and U8873 (N_8873,N_125,N_2159);
and U8874 (N_8874,N_1492,N_4908);
nor U8875 (N_8875,N_4521,N_1329);
nor U8876 (N_8876,N_4554,N_2734);
nor U8877 (N_8877,N_4268,N_4950);
xnor U8878 (N_8878,N_3270,N_2697);
nand U8879 (N_8879,N_684,N_872);
nor U8880 (N_8880,N_2854,N_3919);
nand U8881 (N_8881,N_1169,N_4031);
nor U8882 (N_8882,N_2117,N_2580);
nor U8883 (N_8883,N_2927,N_3616);
and U8884 (N_8884,N_2081,N_781);
xnor U8885 (N_8885,N_2811,N_3075);
xnor U8886 (N_8886,N_4271,N_2481);
nor U8887 (N_8887,N_2890,N_3021);
xor U8888 (N_8888,N_3554,N_2410);
nand U8889 (N_8889,N_163,N_1274);
nor U8890 (N_8890,N_3050,N_1213);
nand U8891 (N_8891,N_812,N_1492);
nor U8892 (N_8892,N_1729,N_3324);
nand U8893 (N_8893,N_2167,N_4849);
and U8894 (N_8894,N_2555,N_1114);
nand U8895 (N_8895,N_784,N_1174);
and U8896 (N_8896,N_2585,N_4456);
nand U8897 (N_8897,N_3252,N_1756);
nor U8898 (N_8898,N_1074,N_4918);
nor U8899 (N_8899,N_107,N_2377);
nor U8900 (N_8900,N_2669,N_135);
nor U8901 (N_8901,N_3339,N_1463);
nor U8902 (N_8902,N_3301,N_1198);
or U8903 (N_8903,N_2841,N_2923);
xor U8904 (N_8904,N_4492,N_4787);
nor U8905 (N_8905,N_4895,N_1234);
xnor U8906 (N_8906,N_3110,N_2544);
or U8907 (N_8907,N_2729,N_3779);
xnor U8908 (N_8908,N_718,N_114);
nand U8909 (N_8909,N_4618,N_2150);
xnor U8910 (N_8910,N_2156,N_2812);
nand U8911 (N_8911,N_2391,N_4834);
xor U8912 (N_8912,N_3776,N_1960);
nand U8913 (N_8913,N_391,N_4886);
nor U8914 (N_8914,N_667,N_1033);
nor U8915 (N_8915,N_3903,N_4646);
or U8916 (N_8916,N_425,N_476);
nor U8917 (N_8917,N_3440,N_4879);
xor U8918 (N_8918,N_1611,N_1932);
nor U8919 (N_8919,N_2327,N_3137);
xor U8920 (N_8920,N_2946,N_4312);
nor U8921 (N_8921,N_148,N_4882);
xnor U8922 (N_8922,N_4855,N_4933);
xnor U8923 (N_8923,N_268,N_1910);
or U8924 (N_8924,N_3616,N_1170);
or U8925 (N_8925,N_1755,N_43);
or U8926 (N_8926,N_1603,N_2233);
nor U8927 (N_8927,N_4866,N_4969);
nor U8928 (N_8928,N_3354,N_209);
or U8929 (N_8929,N_283,N_555);
xnor U8930 (N_8930,N_1171,N_1912);
and U8931 (N_8931,N_4874,N_3084);
xor U8932 (N_8932,N_1416,N_3696);
and U8933 (N_8933,N_3165,N_149);
or U8934 (N_8934,N_2506,N_258);
nand U8935 (N_8935,N_486,N_4077);
xor U8936 (N_8936,N_4062,N_214);
and U8937 (N_8937,N_1608,N_4107);
and U8938 (N_8938,N_3137,N_2802);
nand U8939 (N_8939,N_1114,N_2587);
nor U8940 (N_8940,N_2401,N_3918);
xnor U8941 (N_8941,N_3030,N_4772);
and U8942 (N_8942,N_641,N_4279);
xnor U8943 (N_8943,N_2829,N_2108);
or U8944 (N_8944,N_3462,N_3846);
xor U8945 (N_8945,N_1713,N_1190);
nor U8946 (N_8946,N_4099,N_2801);
nand U8947 (N_8947,N_1553,N_2294);
and U8948 (N_8948,N_1605,N_2720);
nor U8949 (N_8949,N_3551,N_1059);
nor U8950 (N_8950,N_3746,N_122);
or U8951 (N_8951,N_3049,N_4695);
nand U8952 (N_8952,N_392,N_2280);
and U8953 (N_8953,N_4126,N_2869);
nand U8954 (N_8954,N_1078,N_2857);
or U8955 (N_8955,N_1925,N_1748);
and U8956 (N_8956,N_643,N_1905);
or U8957 (N_8957,N_93,N_904);
or U8958 (N_8958,N_3436,N_2893);
or U8959 (N_8959,N_2909,N_4325);
and U8960 (N_8960,N_883,N_4595);
or U8961 (N_8961,N_4402,N_4048);
nand U8962 (N_8962,N_4096,N_237);
and U8963 (N_8963,N_3432,N_2243);
nor U8964 (N_8964,N_1905,N_3270);
nand U8965 (N_8965,N_1777,N_2077);
xnor U8966 (N_8966,N_1890,N_728);
nor U8967 (N_8967,N_1520,N_2096);
or U8968 (N_8968,N_370,N_3826);
and U8969 (N_8969,N_2091,N_4759);
xnor U8970 (N_8970,N_4207,N_1084);
or U8971 (N_8971,N_548,N_1737);
or U8972 (N_8972,N_4048,N_4323);
nand U8973 (N_8973,N_716,N_29);
or U8974 (N_8974,N_62,N_3588);
and U8975 (N_8975,N_2401,N_1761);
or U8976 (N_8976,N_4017,N_1655);
nor U8977 (N_8977,N_4240,N_159);
and U8978 (N_8978,N_4984,N_4077);
and U8979 (N_8979,N_3210,N_1497);
or U8980 (N_8980,N_2049,N_528);
nor U8981 (N_8981,N_2823,N_988);
nor U8982 (N_8982,N_2747,N_2400);
nand U8983 (N_8983,N_3219,N_2014);
nor U8984 (N_8984,N_3131,N_3256);
nand U8985 (N_8985,N_3728,N_281);
or U8986 (N_8986,N_2163,N_1873);
nand U8987 (N_8987,N_1677,N_4477);
nor U8988 (N_8988,N_2198,N_4846);
or U8989 (N_8989,N_3248,N_927);
and U8990 (N_8990,N_4506,N_2982);
xor U8991 (N_8991,N_4727,N_2601);
xor U8992 (N_8992,N_890,N_1094);
or U8993 (N_8993,N_119,N_4716);
and U8994 (N_8994,N_2043,N_3427);
nand U8995 (N_8995,N_3640,N_2208);
xor U8996 (N_8996,N_3583,N_551);
xnor U8997 (N_8997,N_873,N_4427);
nand U8998 (N_8998,N_949,N_439);
nand U8999 (N_8999,N_4465,N_3613);
nor U9000 (N_9000,N_684,N_2803);
xnor U9001 (N_9001,N_553,N_2460);
and U9002 (N_9002,N_3944,N_1457);
and U9003 (N_9003,N_3489,N_3118);
or U9004 (N_9004,N_1722,N_4447);
nand U9005 (N_9005,N_2071,N_1070);
nor U9006 (N_9006,N_800,N_3315);
and U9007 (N_9007,N_3582,N_3723);
nand U9008 (N_9008,N_864,N_1630);
nand U9009 (N_9009,N_1543,N_1227);
xnor U9010 (N_9010,N_1441,N_2850);
xnor U9011 (N_9011,N_1179,N_3660);
nor U9012 (N_9012,N_4474,N_4609);
or U9013 (N_9013,N_2585,N_4273);
nor U9014 (N_9014,N_4508,N_3965);
or U9015 (N_9015,N_133,N_1903);
and U9016 (N_9016,N_4350,N_1243);
nor U9017 (N_9017,N_1760,N_3138);
nor U9018 (N_9018,N_2873,N_1561);
nor U9019 (N_9019,N_99,N_1951);
and U9020 (N_9020,N_4114,N_3595);
xor U9021 (N_9021,N_745,N_2200);
and U9022 (N_9022,N_4687,N_2954);
and U9023 (N_9023,N_4923,N_4994);
and U9024 (N_9024,N_3280,N_2085);
or U9025 (N_9025,N_1689,N_741);
xnor U9026 (N_9026,N_1659,N_3785);
nor U9027 (N_9027,N_2305,N_3734);
or U9028 (N_9028,N_1975,N_4760);
and U9029 (N_9029,N_2160,N_3372);
nand U9030 (N_9030,N_67,N_1320);
nand U9031 (N_9031,N_3414,N_1684);
nand U9032 (N_9032,N_145,N_4630);
xnor U9033 (N_9033,N_1936,N_3160);
and U9034 (N_9034,N_3309,N_2847);
nor U9035 (N_9035,N_776,N_3583);
nand U9036 (N_9036,N_233,N_797);
and U9037 (N_9037,N_1140,N_3232);
or U9038 (N_9038,N_1053,N_3515);
nand U9039 (N_9039,N_1079,N_1869);
nand U9040 (N_9040,N_3095,N_2076);
or U9041 (N_9041,N_4203,N_4625);
and U9042 (N_9042,N_2291,N_498);
or U9043 (N_9043,N_4844,N_4959);
xnor U9044 (N_9044,N_4445,N_4772);
nand U9045 (N_9045,N_1458,N_2684);
and U9046 (N_9046,N_1743,N_3827);
or U9047 (N_9047,N_3337,N_3855);
nor U9048 (N_9048,N_1998,N_3746);
nand U9049 (N_9049,N_1552,N_274);
and U9050 (N_9050,N_2963,N_1673);
nor U9051 (N_9051,N_3103,N_1885);
xor U9052 (N_9052,N_2124,N_377);
nand U9053 (N_9053,N_3818,N_2593);
and U9054 (N_9054,N_3089,N_4830);
or U9055 (N_9055,N_3274,N_1330);
nand U9056 (N_9056,N_997,N_2804);
and U9057 (N_9057,N_969,N_3602);
nor U9058 (N_9058,N_3807,N_427);
and U9059 (N_9059,N_2681,N_688);
nor U9060 (N_9060,N_1112,N_4940);
xnor U9061 (N_9061,N_204,N_3638);
nand U9062 (N_9062,N_4317,N_4603);
nor U9063 (N_9063,N_440,N_846);
nand U9064 (N_9064,N_3486,N_4607);
and U9065 (N_9065,N_1855,N_456);
and U9066 (N_9066,N_1775,N_4558);
xnor U9067 (N_9067,N_4766,N_969);
xnor U9068 (N_9068,N_2133,N_1149);
nand U9069 (N_9069,N_1091,N_1631);
nand U9070 (N_9070,N_2808,N_3367);
xnor U9071 (N_9071,N_3119,N_3516);
xor U9072 (N_9072,N_4185,N_4980);
nand U9073 (N_9073,N_1345,N_304);
xor U9074 (N_9074,N_4198,N_2820);
nor U9075 (N_9075,N_3619,N_2282);
and U9076 (N_9076,N_4903,N_2287);
or U9077 (N_9077,N_4862,N_882);
nor U9078 (N_9078,N_403,N_1536);
or U9079 (N_9079,N_1216,N_2833);
and U9080 (N_9080,N_1967,N_3920);
or U9081 (N_9081,N_1,N_510);
or U9082 (N_9082,N_4972,N_4315);
and U9083 (N_9083,N_1001,N_422);
nand U9084 (N_9084,N_3172,N_3384);
and U9085 (N_9085,N_3397,N_1678);
xnor U9086 (N_9086,N_4558,N_2089);
or U9087 (N_9087,N_3382,N_3997);
and U9088 (N_9088,N_4764,N_2306);
and U9089 (N_9089,N_4392,N_1938);
and U9090 (N_9090,N_345,N_580);
and U9091 (N_9091,N_2182,N_2576);
and U9092 (N_9092,N_792,N_184);
xor U9093 (N_9093,N_4773,N_2692);
nand U9094 (N_9094,N_3926,N_818);
xor U9095 (N_9095,N_178,N_434);
xnor U9096 (N_9096,N_3388,N_3498);
xor U9097 (N_9097,N_2550,N_3786);
and U9098 (N_9098,N_4581,N_1627);
xor U9099 (N_9099,N_1595,N_2071);
nand U9100 (N_9100,N_999,N_804);
nor U9101 (N_9101,N_178,N_1868);
or U9102 (N_9102,N_1415,N_3228);
and U9103 (N_9103,N_3311,N_1856);
nand U9104 (N_9104,N_4123,N_3477);
nor U9105 (N_9105,N_1674,N_95);
xnor U9106 (N_9106,N_2292,N_4145);
nand U9107 (N_9107,N_3642,N_4209);
or U9108 (N_9108,N_4282,N_4817);
and U9109 (N_9109,N_156,N_1105);
nand U9110 (N_9110,N_3937,N_4342);
or U9111 (N_9111,N_3952,N_2188);
xor U9112 (N_9112,N_4699,N_3469);
nand U9113 (N_9113,N_2837,N_2411);
nor U9114 (N_9114,N_1913,N_3860);
or U9115 (N_9115,N_589,N_2595);
xor U9116 (N_9116,N_4868,N_4765);
nand U9117 (N_9117,N_311,N_4322);
and U9118 (N_9118,N_2002,N_4535);
and U9119 (N_9119,N_4886,N_2850);
and U9120 (N_9120,N_3174,N_4553);
and U9121 (N_9121,N_4031,N_492);
and U9122 (N_9122,N_4604,N_2774);
xnor U9123 (N_9123,N_4419,N_3463);
nand U9124 (N_9124,N_4500,N_764);
or U9125 (N_9125,N_1611,N_4373);
xnor U9126 (N_9126,N_789,N_1699);
and U9127 (N_9127,N_1951,N_1795);
xor U9128 (N_9128,N_1597,N_4939);
or U9129 (N_9129,N_4612,N_1457);
nand U9130 (N_9130,N_684,N_4430);
or U9131 (N_9131,N_1793,N_4302);
and U9132 (N_9132,N_694,N_3117);
and U9133 (N_9133,N_170,N_446);
or U9134 (N_9134,N_1544,N_2765);
and U9135 (N_9135,N_2002,N_2915);
and U9136 (N_9136,N_3453,N_4142);
and U9137 (N_9137,N_1259,N_4773);
and U9138 (N_9138,N_2555,N_4443);
and U9139 (N_9139,N_4663,N_2774);
nor U9140 (N_9140,N_1528,N_1500);
xnor U9141 (N_9141,N_3762,N_600);
nand U9142 (N_9142,N_611,N_4561);
nor U9143 (N_9143,N_2491,N_3297);
xor U9144 (N_9144,N_896,N_717);
or U9145 (N_9145,N_3626,N_3276);
or U9146 (N_9146,N_2886,N_4700);
or U9147 (N_9147,N_1450,N_2362);
nor U9148 (N_9148,N_2022,N_37);
and U9149 (N_9149,N_4844,N_3138);
nand U9150 (N_9150,N_1079,N_3023);
and U9151 (N_9151,N_208,N_1735);
nor U9152 (N_9152,N_52,N_3958);
xor U9153 (N_9153,N_4075,N_3400);
nand U9154 (N_9154,N_4407,N_4570);
and U9155 (N_9155,N_1130,N_1743);
and U9156 (N_9156,N_2723,N_1209);
nand U9157 (N_9157,N_4459,N_1444);
and U9158 (N_9158,N_63,N_4804);
nand U9159 (N_9159,N_536,N_4124);
nor U9160 (N_9160,N_2909,N_3098);
nor U9161 (N_9161,N_870,N_3569);
or U9162 (N_9162,N_3728,N_3676);
nand U9163 (N_9163,N_2767,N_2577);
or U9164 (N_9164,N_4494,N_862);
or U9165 (N_9165,N_265,N_2197);
nor U9166 (N_9166,N_2502,N_2020);
xor U9167 (N_9167,N_900,N_2427);
and U9168 (N_9168,N_1694,N_1941);
nor U9169 (N_9169,N_235,N_4751);
nand U9170 (N_9170,N_285,N_1129);
or U9171 (N_9171,N_2845,N_2372);
xor U9172 (N_9172,N_4648,N_422);
xnor U9173 (N_9173,N_1276,N_1461);
xnor U9174 (N_9174,N_4791,N_3000);
or U9175 (N_9175,N_3648,N_780);
and U9176 (N_9176,N_1553,N_4957);
and U9177 (N_9177,N_3750,N_3391);
and U9178 (N_9178,N_4827,N_2553);
and U9179 (N_9179,N_3798,N_3285);
nor U9180 (N_9180,N_624,N_3468);
nor U9181 (N_9181,N_626,N_2668);
xor U9182 (N_9182,N_1332,N_4005);
and U9183 (N_9183,N_968,N_594);
nor U9184 (N_9184,N_2464,N_762);
xor U9185 (N_9185,N_555,N_2848);
xnor U9186 (N_9186,N_4390,N_3236);
nand U9187 (N_9187,N_937,N_7);
and U9188 (N_9188,N_3957,N_4325);
nor U9189 (N_9189,N_3857,N_1443);
nand U9190 (N_9190,N_4415,N_150);
nand U9191 (N_9191,N_2925,N_3484);
and U9192 (N_9192,N_1872,N_1129);
or U9193 (N_9193,N_1301,N_3962);
and U9194 (N_9194,N_3448,N_593);
nand U9195 (N_9195,N_3558,N_758);
nor U9196 (N_9196,N_190,N_3749);
and U9197 (N_9197,N_3437,N_2789);
xnor U9198 (N_9198,N_88,N_4599);
xor U9199 (N_9199,N_2791,N_3790);
and U9200 (N_9200,N_2717,N_3745);
and U9201 (N_9201,N_4328,N_932);
xor U9202 (N_9202,N_4676,N_811);
xnor U9203 (N_9203,N_4368,N_4049);
xor U9204 (N_9204,N_616,N_3998);
or U9205 (N_9205,N_1605,N_3220);
and U9206 (N_9206,N_3754,N_1865);
and U9207 (N_9207,N_1356,N_3481);
or U9208 (N_9208,N_1112,N_1945);
nand U9209 (N_9209,N_551,N_1400);
nand U9210 (N_9210,N_1117,N_778);
nor U9211 (N_9211,N_2496,N_2205);
and U9212 (N_9212,N_4544,N_1108);
and U9213 (N_9213,N_3916,N_2421);
and U9214 (N_9214,N_1811,N_4905);
nor U9215 (N_9215,N_2657,N_3859);
nand U9216 (N_9216,N_1959,N_256);
and U9217 (N_9217,N_487,N_31);
xor U9218 (N_9218,N_504,N_1236);
and U9219 (N_9219,N_4625,N_1608);
or U9220 (N_9220,N_2140,N_1733);
and U9221 (N_9221,N_4626,N_4867);
or U9222 (N_9222,N_474,N_4267);
or U9223 (N_9223,N_884,N_1941);
nor U9224 (N_9224,N_2543,N_2593);
nand U9225 (N_9225,N_2248,N_1846);
or U9226 (N_9226,N_1160,N_3867);
nand U9227 (N_9227,N_4757,N_2545);
nor U9228 (N_9228,N_3742,N_719);
xor U9229 (N_9229,N_274,N_1660);
nand U9230 (N_9230,N_777,N_1000);
or U9231 (N_9231,N_4923,N_2223);
xor U9232 (N_9232,N_3579,N_2034);
nor U9233 (N_9233,N_1105,N_534);
or U9234 (N_9234,N_843,N_3040);
xor U9235 (N_9235,N_3269,N_3206);
and U9236 (N_9236,N_3268,N_2344);
nor U9237 (N_9237,N_4968,N_2090);
nand U9238 (N_9238,N_4548,N_4714);
nand U9239 (N_9239,N_4367,N_4950);
xor U9240 (N_9240,N_4738,N_1218);
or U9241 (N_9241,N_3750,N_3157);
nor U9242 (N_9242,N_1124,N_2632);
nor U9243 (N_9243,N_2791,N_818);
xnor U9244 (N_9244,N_48,N_2549);
xor U9245 (N_9245,N_1801,N_1163);
nor U9246 (N_9246,N_4852,N_2655);
and U9247 (N_9247,N_2455,N_1142);
and U9248 (N_9248,N_390,N_4165);
xnor U9249 (N_9249,N_707,N_839);
nand U9250 (N_9250,N_2677,N_2372);
xor U9251 (N_9251,N_2114,N_3982);
xor U9252 (N_9252,N_2420,N_1921);
nand U9253 (N_9253,N_1113,N_151);
or U9254 (N_9254,N_343,N_3786);
xnor U9255 (N_9255,N_301,N_905);
nor U9256 (N_9256,N_4530,N_1861);
and U9257 (N_9257,N_3616,N_190);
nor U9258 (N_9258,N_3161,N_3925);
xnor U9259 (N_9259,N_3267,N_1276);
nor U9260 (N_9260,N_4215,N_879);
xor U9261 (N_9261,N_15,N_3917);
nor U9262 (N_9262,N_4492,N_1735);
nand U9263 (N_9263,N_4490,N_357);
xnor U9264 (N_9264,N_1104,N_1200);
or U9265 (N_9265,N_1811,N_4098);
nor U9266 (N_9266,N_282,N_2869);
nand U9267 (N_9267,N_518,N_4188);
nor U9268 (N_9268,N_1573,N_2565);
xor U9269 (N_9269,N_2011,N_1004);
xnor U9270 (N_9270,N_4243,N_994);
nor U9271 (N_9271,N_4817,N_1893);
nand U9272 (N_9272,N_4690,N_1610);
xor U9273 (N_9273,N_2698,N_3195);
or U9274 (N_9274,N_2390,N_3904);
nand U9275 (N_9275,N_3356,N_1246);
nand U9276 (N_9276,N_3044,N_3826);
and U9277 (N_9277,N_3399,N_4094);
or U9278 (N_9278,N_1838,N_2417);
or U9279 (N_9279,N_4995,N_4762);
nor U9280 (N_9280,N_1527,N_4584);
or U9281 (N_9281,N_4006,N_2342);
and U9282 (N_9282,N_962,N_2906);
xnor U9283 (N_9283,N_2491,N_2961);
and U9284 (N_9284,N_2106,N_533);
nor U9285 (N_9285,N_3202,N_1908);
nor U9286 (N_9286,N_4716,N_2528);
and U9287 (N_9287,N_2700,N_2146);
and U9288 (N_9288,N_4329,N_1441);
nor U9289 (N_9289,N_4739,N_3629);
nand U9290 (N_9290,N_2804,N_2216);
or U9291 (N_9291,N_2097,N_2647);
or U9292 (N_9292,N_2889,N_1853);
nor U9293 (N_9293,N_1466,N_1479);
or U9294 (N_9294,N_1671,N_2610);
and U9295 (N_9295,N_4892,N_2256);
nor U9296 (N_9296,N_4971,N_1479);
xor U9297 (N_9297,N_469,N_1302);
or U9298 (N_9298,N_120,N_3721);
nand U9299 (N_9299,N_597,N_828);
or U9300 (N_9300,N_2661,N_2524);
nor U9301 (N_9301,N_1277,N_1694);
xor U9302 (N_9302,N_528,N_3365);
xor U9303 (N_9303,N_1592,N_3257);
or U9304 (N_9304,N_1790,N_3492);
nor U9305 (N_9305,N_1398,N_3336);
nand U9306 (N_9306,N_467,N_303);
or U9307 (N_9307,N_3010,N_217);
and U9308 (N_9308,N_4090,N_2200);
nand U9309 (N_9309,N_3322,N_11);
nand U9310 (N_9310,N_377,N_3587);
and U9311 (N_9311,N_4416,N_3013);
nand U9312 (N_9312,N_4770,N_2400);
or U9313 (N_9313,N_808,N_1293);
nand U9314 (N_9314,N_1253,N_3998);
or U9315 (N_9315,N_3976,N_504);
nand U9316 (N_9316,N_4646,N_4045);
or U9317 (N_9317,N_4363,N_772);
nor U9318 (N_9318,N_3898,N_3124);
or U9319 (N_9319,N_503,N_4183);
nand U9320 (N_9320,N_4201,N_824);
nor U9321 (N_9321,N_1599,N_889);
or U9322 (N_9322,N_4936,N_453);
or U9323 (N_9323,N_2758,N_1557);
xnor U9324 (N_9324,N_1314,N_4647);
and U9325 (N_9325,N_1988,N_4162);
xnor U9326 (N_9326,N_3778,N_3267);
nor U9327 (N_9327,N_1227,N_3817);
nand U9328 (N_9328,N_4222,N_1588);
nor U9329 (N_9329,N_1237,N_2642);
or U9330 (N_9330,N_831,N_1294);
xor U9331 (N_9331,N_1590,N_4913);
nor U9332 (N_9332,N_1050,N_3281);
and U9333 (N_9333,N_665,N_512);
or U9334 (N_9334,N_434,N_2716);
xnor U9335 (N_9335,N_2286,N_2219);
nor U9336 (N_9336,N_2434,N_3457);
nor U9337 (N_9337,N_853,N_3030);
xor U9338 (N_9338,N_4618,N_3427);
xnor U9339 (N_9339,N_2671,N_3309);
or U9340 (N_9340,N_272,N_446);
nand U9341 (N_9341,N_4304,N_3437);
nor U9342 (N_9342,N_2485,N_552);
and U9343 (N_9343,N_197,N_666);
or U9344 (N_9344,N_121,N_3702);
nand U9345 (N_9345,N_1405,N_516);
and U9346 (N_9346,N_68,N_3150);
and U9347 (N_9347,N_3097,N_4805);
xor U9348 (N_9348,N_4793,N_4327);
nand U9349 (N_9349,N_1238,N_4362);
nand U9350 (N_9350,N_4302,N_4741);
nor U9351 (N_9351,N_2612,N_3587);
and U9352 (N_9352,N_2682,N_1684);
nand U9353 (N_9353,N_2923,N_4514);
or U9354 (N_9354,N_1224,N_995);
nand U9355 (N_9355,N_3003,N_4212);
nand U9356 (N_9356,N_3877,N_2915);
xor U9357 (N_9357,N_1566,N_1733);
nor U9358 (N_9358,N_3897,N_2478);
xnor U9359 (N_9359,N_2821,N_759);
nor U9360 (N_9360,N_2095,N_4509);
or U9361 (N_9361,N_1063,N_3906);
or U9362 (N_9362,N_3647,N_1364);
and U9363 (N_9363,N_2019,N_3434);
and U9364 (N_9364,N_1556,N_4753);
nor U9365 (N_9365,N_282,N_4720);
nor U9366 (N_9366,N_1085,N_2997);
xnor U9367 (N_9367,N_2128,N_752);
xor U9368 (N_9368,N_95,N_1506);
nor U9369 (N_9369,N_565,N_343);
and U9370 (N_9370,N_403,N_1067);
xnor U9371 (N_9371,N_2428,N_3181);
or U9372 (N_9372,N_670,N_1789);
xnor U9373 (N_9373,N_4700,N_1669);
or U9374 (N_9374,N_4200,N_2250);
nand U9375 (N_9375,N_4417,N_4274);
nand U9376 (N_9376,N_2601,N_3853);
nor U9377 (N_9377,N_4100,N_4538);
or U9378 (N_9378,N_3406,N_3750);
and U9379 (N_9379,N_514,N_3909);
or U9380 (N_9380,N_3453,N_2065);
xnor U9381 (N_9381,N_2248,N_84);
xnor U9382 (N_9382,N_2492,N_383);
or U9383 (N_9383,N_4586,N_1633);
and U9384 (N_9384,N_696,N_2074);
or U9385 (N_9385,N_4543,N_491);
nand U9386 (N_9386,N_177,N_701);
nand U9387 (N_9387,N_2330,N_2314);
and U9388 (N_9388,N_3849,N_4400);
nor U9389 (N_9389,N_4852,N_2414);
xnor U9390 (N_9390,N_3312,N_1966);
nor U9391 (N_9391,N_238,N_2307);
or U9392 (N_9392,N_4714,N_1075);
nand U9393 (N_9393,N_741,N_2880);
and U9394 (N_9394,N_1485,N_3007);
nor U9395 (N_9395,N_2594,N_1223);
xor U9396 (N_9396,N_4716,N_3103);
or U9397 (N_9397,N_1716,N_2078);
or U9398 (N_9398,N_3853,N_1569);
nand U9399 (N_9399,N_2701,N_534);
or U9400 (N_9400,N_1977,N_1019);
xor U9401 (N_9401,N_3396,N_947);
or U9402 (N_9402,N_3673,N_1543);
xor U9403 (N_9403,N_4112,N_1016);
nand U9404 (N_9404,N_3299,N_4481);
nand U9405 (N_9405,N_2645,N_4804);
xnor U9406 (N_9406,N_873,N_552);
and U9407 (N_9407,N_4526,N_3466);
nor U9408 (N_9408,N_3225,N_953);
and U9409 (N_9409,N_2745,N_3709);
xnor U9410 (N_9410,N_3284,N_18);
nor U9411 (N_9411,N_1410,N_2086);
nor U9412 (N_9412,N_3918,N_1100);
xnor U9413 (N_9413,N_142,N_2617);
or U9414 (N_9414,N_2017,N_134);
nand U9415 (N_9415,N_149,N_1837);
and U9416 (N_9416,N_999,N_1910);
and U9417 (N_9417,N_512,N_4913);
and U9418 (N_9418,N_1195,N_644);
and U9419 (N_9419,N_4537,N_48);
nor U9420 (N_9420,N_3341,N_2810);
and U9421 (N_9421,N_763,N_1404);
xor U9422 (N_9422,N_4188,N_1896);
and U9423 (N_9423,N_1390,N_2781);
and U9424 (N_9424,N_602,N_3970);
nand U9425 (N_9425,N_1635,N_425);
nor U9426 (N_9426,N_1858,N_1968);
nor U9427 (N_9427,N_4245,N_230);
nor U9428 (N_9428,N_1377,N_1589);
or U9429 (N_9429,N_4907,N_4530);
nor U9430 (N_9430,N_1815,N_969);
xnor U9431 (N_9431,N_1148,N_2624);
xor U9432 (N_9432,N_1285,N_4901);
nor U9433 (N_9433,N_203,N_542);
nand U9434 (N_9434,N_2032,N_1190);
xnor U9435 (N_9435,N_2387,N_3415);
and U9436 (N_9436,N_729,N_1032);
nand U9437 (N_9437,N_1869,N_2816);
or U9438 (N_9438,N_4242,N_1592);
nor U9439 (N_9439,N_922,N_2241);
xnor U9440 (N_9440,N_14,N_1763);
xor U9441 (N_9441,N_4890,N_3484);
nand U9442 (N_9442,N_291,N_826);
xor U9443 (N_9443,N_3420,N_200);
and U9444 (N_9444,N_4298,N_3964);
xnor U9445 (N_9445,N_2598,N_1981);
xor U9446 (N_9446,N_3551,N_3157);
and U9447 (N_9447,N_3652,N_367);
nand U9448 (N_9448,N_1594,N_2715);
nor U9449 (N_9449,N_1948,N_347);
and U9450 (N_9450,N_2718,N_1200);
nand U9451 (N_9451,N_3891,N_59);
nor U9452 (N_9452,N_1324,N_4677);
and U9453 (N_9453,N_3940,N_970);
xor U9454 (N_9454,N_1975,N_3877);
nor U9455 (N_9455,N_579,N_907);
or U9456 (N_9456,N_1648,N_2935);
xnor U9457 (N_9457,N_2579,N_4491);
nor U9458 (N_9458,N_1431,N_1397);
nand U9459 (N_9459,N_3620,N_286);
nand U9460 (N_9460,N_4154,N_273);
nand U9461 (N_9461,N_1796,N_1142);
nand U9462 (N_9462,N_2577,N_3286);
nand U9463 (N_9463,N_3465,N_4619);
xnor U9464 (N_9464,N_679,N_241);
xor U9465 (N_9465,N_722,N_3131);
or U9466 (N_9466,N_2562,N_1417);
or U9467 (N_9467,N_803,N_2555);
nand U9468 (N_9468,N_3676,N_1361);
or U9469 (N_9469,N_3359,N_196);
and U9470 (N_9470,N_836,N_3206);
or U9471 (N_9471,N_3002,N_3871);
xor U9472 (N_9472,N_1551,N_1071);
and U9473 (N_9473,N_683,N_4323);
nor U9474 (N_9474,N_3065,N_3345);
and U9475 (N_9475,N_4509,N_378);
nand U9476 (N_9476,N_2363,N_780);
nand U9477 (N_9477,N_1855,N_4629);
nand U9478 (N_9478,N_441,N_73);
and U9479 (N_9479,N_958,N_2575);
xor U9480 (N_9480,N_1601,N_1387);
xor U9481 (N_9481,N_4449,N_4475);
and U9482 (N_9482,N_2595,N_3587);
nand U9483 (N_9483,N_2191,N_2750);
nor U9484 (N_9484,N_4991,N_484);
nand U9485 (N_9485,N_2579,N_3940);
xor U9486 (N_9486,N_1177,N_4845);
and U9487 (N_9487,N_4349,N_3665);
nand U9488 (N_9488,N_2769,N_3108);
and U9489 (N_9489,N_4175,N_3572);
or U9490 (N_9490,N_1218,N_4058);
or U9491 (N_9491,N_1667,N_1430);
xnor U9492 (N_9492,N_2997,N_3683);
xor U9493 (N_9493,N_385,N_15);
or U9494 (N_9494,N_1121,N_4647);
and U9495 (N_9495,N_326,N_270);
and U9496 (N_9496,N_2271,N_1971);
nand U9497 (N_9497,N_212,N_2434);
nand U9498 (N_9498,N_2317,N_1357);
and U9499 (N_9499,N_2344,N_942);
nand U9500 (N_9500,N_994,N_374);
nor U9501 (N_9501,N_1296,N_574);
nor U9502 (N_9502,N_3554,N_1365);
nor U9503 (N_9503,N_2760,N_333);
or U9504 (N_9504,N_842,N_4207);
nor U9505 (N_9505,N_3328,N_267);
xnor U9506 (N_9506,N_564,N_20);
xnor U9507 (N_9507,N_4077,N_3401);
or U9508 (N_9508,N_1550,N_1374);
or U9509 (N_9509,N_2874,N_268);
nand U9510 (N_9510,N_4140,N_3855);
nor U9511 (N_9511,N_1193,N_3541);
xor U9512 (N_9512,N_1042,N_4307);
nand U9513 (N_9513,N_604,N_4025);
and U9514 (N_9514,N_4949,N_2582);
nor U9515 (N_9515,N_329,N_3998);
or U9516 (N_9516,N_2637,N_1925);
nand U9517 (N_9517,N_821,N_350);
xor U9518 (N_9518,N_893,N_1244);
or U9519 (N_9519,N_3247,N_2064);
nor U9520 (N_9520,N_3094,N_3995);
or U9521 (N_9521,N_2487,N_2081);
nor U9522 (N_9522,N_4525,N_2786);
or U9523 (N_9523,N_996,N_4059);
and U9524 (N_9524,N_7,N_1081);
xnor U9525 (N_9525,N_710,N_4942);
or U9526 (N_9526,N_2430,N_864);
nor U9527 (N_9527,N_17,N_2136);
nand U9528 (N_9528,N_1619,N_2224);
xnor U9529 (N_9529,N_3009,N_3539);
nand U9530 (N_9530,N_1446,N_823);
or U9531 (N_9531,N_1897,N_1390);
nand U9532 (N_9532,N_1471,N_2552);
xor U9533 (N_9533,N_1059,N_1123);
nor U9534 (N_9534,N_2571,N_3716);
nand U9535 (N_9535,N_2426,N_3210);
or U9536 (N_9536,N_4925,N_1340);
nor U9537 (N_9537,N_665,N_692);
nand U9538 (N_9538,N_894,N_1328);
nor U9539 (N_9539,N_3532,N_1935);
nor U9540 (N_9540,N_4588,N_267);
or U9541 (N_9541,N_3487,N_3013);
nand U9542 (N_9542,N_559,N_3133);
nand U9543 (N_9543,N_634,N_1620);
nand U9544 (N_9544,N_4561,N_136);
nor U9545 (N_9545,N_4270,N_1940);
and U9546 (N_9546,N_4517,N_3034);
nor U9547 (N_9547,N_459,N_3245);
nand U9548 (N_9548,N_4138,N_2124);
nor U9549 (N_9549,N_1065,N_1264);
xnor U9550 (N_9550,N_2000,N_2859);
nor U9551 (N_9551,N_1141,N_3408);
nand U9552 (N_9552,N_2941,N_4792);
or U9553 (N_9553,N_2880,N_4058);
and U9554 (N_9554,N_3568,N_4632);
nor U9555 (N_9555,N_4792,N_2285);
or U9556 (N_9556,N_2582,N_996);
or U9557 (N_9557,N_1603,N_3253);
nor U9558 (N_9558,N_1418,N_2396);
xor U9559 (N_9559,N_17,N_1440);
or U9560 (N_9560,N_1970,N_1881);
and U9561 (N_9561,N_1934,N_2330);
nor U9562 (N_9562,N_86,N_2708);
and U9563 (N_9563,N_1606,N_3919);
nand U9564 (N_9564,N_4164,N_3359);
nand U9565 (N_9565,N_2677,N_2200);
nor U9566 (N_9566,N_3663,N_4154);
nor U9567 (N_9567,N_2236,N_3511);
or U9568 (N_9568,N_3368,N_3287);
xnor U9569 (N_9569,N_2035,N_2446);
xor U9570 (N_9570,N_533,N_3473);
or U9571 (N_9571,N_4811,N_2244);
xnor U9572 (N_9572,N_4294,N_4809);
and U9573 (N_9573,N_2050,N_489);
xor U9574 (N_9574,N_845,N_3352);
xor U9575 (N_9575,N_861,N_666);
nor U9576 (N_9576,N_2692,N_3183);
and U9577 (N_9577,N_4339,N_3569);
or U9578 (N_9578,N_2560,N_372);
nand U9579 (N_9579,N_150,N_2226);
nand U9580 (N_9580,N_974,N_297);
xnor U9581 (N_9581,N_1963,N_4056);
xor U9582 (N_9582,N_4936,N_2515);
nor U9583 (N_9583,N_653,N_4750);
nand U9584 (N_9584,N_4851,N_1943);
xor U9585 (N_9585,N_2649,N_876);
nand U9586 (N_9586,N_2242,N_4414);
nor U9587 (N_9587,N_4680,N_4037);
or U9588 (N_9588,N_1608,N_2235);
xnor U9589 (N_9589,N_1613,N_3175);
and U9590 (N_9590,N_3599,N_3934);
xor U9591 (N_9591,N_4967,N_2049);
xor U9592 (N_9592,N_2106,N_1458);
nand U9593 (N_9593,N_1903,N_3063);
or U9594 (N_9594,N_1871,N_1087);
nand U9595 (N_9595,N_1035,N_1231);
nor U9596 (N_9596,N_2315,N_3819);
and U9597 (N_9597,N_4703,N_2223);
xnor U9598 (N_9598,N_1142,N_1573);
nor U9599 (N_9599,N_930,N_1012);
nor U9600 (N_9600,N_3240,N_1331);
xnor U9601 (N_9601,N_1405,N_1277);
xor U9602 (N_9602,N_3450,N_3930);
or U9603 (N_9603,N_2521,N_4009);
nand U9604 (N_9604,N_1161,N_4509);
xor U9605 (N_9605,N_1850,N_3259);
and U9606 (N_9606,N_810,N_2598);
nand U9607 (N_9607,N_1533,N_2118);
xnor U9608 (N_9608,N_2737,N_2134);
nand U9609 (N_9609,N_890,N_3322);
or U9610 (N_9610,N_323,N_181);
nand U9611 (N_9611,N_3680,N_1200);
or U9612 (N_9612,N_638,N_4561);
xor U9613 (N_9613,N_2500,N_754);
xnor U9614 (N_9614,N_1700,N_4378);
xor U9615 (N_9615,N_2827,N_849);
and U9616 (N_9616,N_2296,N_2305);
nor U9617 (N_9617,N_4963,N_1829);
nor U9618 (N_9618,N_1460,N_113);
nor U9619 (N_9619,N_2241,N_1962);
or U9620 (N_9620,N_4507,N_3452);
nor U9621 (N_9621,N_151,N_698);
nand U9622 (N_9622,N_1696,N_4721);
or U9623 (N_9623,N_846,N_3174);
xnor U9624 (N_9624,N_654,N_2623);
nand U9625 (N_9625,N_2537,N_1472);
and U9626 (N_9626,N_2733,N_1830);
xor U9627 (N_9627,N_2280,N_25);
nor U9628 (N_9628,N_3374,N_1997);
and U9629 (N_9629,N_2831,N_4773);
nand U9630 (N_9630,N_4973,N_3342);
nor U9631 (N_9631,N_2172,N_3257);
xor U9632 (N_9632,N_2735,N_4323);
nand U9633 (N_9633,N_763,N_4284);
or U9634 (N_9634,N_4842,N_3107);
xnor U9635 (N_9635,N_2943,N_1811);
and U9636 (N_9636,N_2789,N_4105);
nor U9637 (N_9637,N_2910,N_2704);
or U9638 (N_9638,N_1858,N_987);
and U9639 (N_9639,N_4997,N_2780);
nand U9640 (N_9640,N_4577,N_392);
or U9641 (N_9641,N_2043,N_4866);
nand U9642 (N_9642,N_1448,N_998);
xnor U9643 (N_9643,N_479,N_4303);
nor U9644 (N_9644,N_2021,N_1861);
or U9645 (N_9645,N_2715,N_3962);
nor U9646 (N_9646,N_4807,N_245);
or U9647 (N_9647,N_4136,N_2981);
or U9648 (N_9648,N_2588,N_2437);
xor U9649 (N_9649,N_1916,N_3279);
or U9650 (N_9650,N_2639,N_3771);
nand U9651 (N_9651,N_1014,N_3594);
and U9652 (N_9652,N_221,N_2991);
or U9653 (N_9653,N_2583,N_1657);
nor U9654 (N_9654,N_4007,N_4123);
xnor U9655 (N_9655,N_4829,N_2486);
nand U9656 (N_9656,N_2909,N_62);
and U9657 (N_9657,N_1729,N_4085);
or U9658 (N_9658,N_234,N_2676);
nand U9659 (N_9659,N_2135,N_1361);
xnor U9660 (N_9660,N_1028,N_3628);
or U9661 (N_9661,N_1466,N_533);
xor U9662 (N_9662,N_2475,N_1700);
or U9663 (N_9663,N_651,N_3252);
and U9664 (N_9664,N_1585,N_1179);
nand U9665 (N_9665,N_3722,N_3785);
nand U9666 (N_9666,N_4912,N_4340);
nor U9667 (N_9667,N_4245,N_613);
or U9668 (N_9668,N_4328,N_963);
and U9669 (N_9669,N_1867,N_877);
and U9670 (N_9670,N_4228,N_551);
nand U9671 (N_9671,N_3670,N_3416);
or U9672 (N_9672,N_621,N_2315);
or U9673 (N_9673,N_4331,N_958);
nand U9674 (N_9674,N_1182,N_439);
or U9675 (N_9675,N_2100,N_1075);
nand U9676 (N_9676,N_1025,N_4778);
or U9677 (N_9677,N_3529,N_2726);
and U9678 (N_9678,N_1574,N_3444);
nor U9679 (N_9679,N_1010,N_3131);
xor U9680 (N_9680,N_1048,N_4235);
xnor U9681 (N_9681,N_4453,N_2334);
or U9682 (N_9682,N_3613,N_4389);
xnor U9683 (N_9683,N_4608,N_1068);
nand U9684 (N_9684,N_446,N_2684);
and U9685 (N_9685,N_3343,N_448);
nor U9686 (N_9686,N_4269,N_4635);
nor U9687 (N_9687,N_3550,N_2078);
nor U9688 (N_9688,N_1659,N_2792);
or U9689 (N_9689,N_463,N_1988);
nand U9690 (N_9690,N_905,N_4816);
nand U9691 (N_9691,N_1699,N_920);
xnor U9692 (N_9692,N_240,N_3112);
nand U9693 (N_9693,N_4944,N_2729);
nor U9694 (N_9694,N_2423,N_1130);
xnor U9695 (N_9695,N_3571,N_768);
or U9696 (N_9696,N_1789,N_3532);
and U9697 (N_9697,N_2470,N_617);
xor U9698 (N_9698,N_4406,N_1438);
or U9699 (N_9699,N_4700,N_4405);
nand U9700 (N_9700,N_225,N_1683);
or U9701 (N_9701,N_1076,N_1782);
or U9702 (N_9702,N_1004,N_1318);
xnor U9703 (N_9703,N_748,N_3270);
nor U9704 (N_9704,N_3050,N_605);
nand U9705 (N_9705,N_4794,N_2695);
nand U9706 (N_9706,N_3946,N_4080);
nand U9707 (N_9707,N_2358,N_278);
xor U9708 (N_9708,N_2640,N_936);
nor U9709 (N_9709,N_1355,N_3376);
xor U9710 (N_9710,N_4324,N_1733);
or U9711 (N_9711,N_2488,N_37);
nor U9712 (N_9712,N_3456,N_2997);
or U9713 (N_9713,N_4351,N_2686);
or U9714 (N_9714,N_2609,N_1225);
nand U9715 (N_9715,N_321,N_1736);
or U9716 (N_9716,N_4660,N_927);
or U9717 (N_9717,N_4237,N_1451);
nor U9718 (N_9718,N_935,N_4324);
or U9719 (N_9719,N_1736,N_3731);
and U9720 (N_9720,N_2732,N_3207);
or U9721 (N_9721,N_1721,N_4972);
nor U9722 (N_9722,N_795,N_1505);
or U9723 (N_9723,N_2674,N_4650);
xor U9724 (N_9724,N_4500,N_2733);
and U9725 (N_9725,N_1537,N_2236);
xor U9726 (N_9726,N_2073,N_2224);
xnor U9727 (N_9727,N_3842,N_1852);
nand U9728 (N_9728,N_4815,N_2789);
and U9729 (N_9729,N_1939,N_4441);
xnor U9730 (N_9730,N_1358,N_3746);
nand U9731 (N_9731,N_1953,N_681);
xor U9732 (N_9732,N_2513,N_460);
nor U9733 (N_9733,N_2508,N_4035);
and U9734 (N_9734,N_3169,N_2449);
nand U9735 (N_9735,N_251,N_2617);
or U9736 (N_9736,N_581,N_3768);
or U9737 (N_9737,N_2625,N_2933);
and U9738 (N_9738,N_2103,N_4608);
xnor U9739 (N_9739,N_225,N_4358);
xnor U9740 (N_9740,N_1867,N_1209);
nand U9741 (N_9741,N_3615,N_1416);
xnor U9742 (N_9742,N_1409,N_3397);
xor U9743 (N_9743,N_3245,N_2939);
or U9744 (N_9744,N_1319,N_3657);
xor U9745 (N_9745,N_3226,N_1547);
or U9746 (N_9746,N_289,N_977);
or U9747 (N_9747,N_3316,N_1395);
xor U9748 (N_9748,N_4869,N_2194);
xor U9749 (N_9749,N_2938,N_4480);
xnor U9750 (N_9750,N_918,N_3841);
or U9751 (N_9751,N_1511,N_1051);
xor U9752 (N_9752,N_979,N_1861);
and U9753 (N_9753,N_23,N_4775);
and U9754 (N_9754,N_4820,N_1027);
nand U9755 (N_9755,N_2526,N_3029);
nand U9756 (N_9756,N_3930,N_3157);
nand U9757 (N_9757,N_3382,N_522);
and U9758 (N_9758,N_245,N_873);
and U9759 (N_9759,N_4693,N_2179);
nand U9760 (N_9760,N_2345,N_2328);
xor U9761 (N_9761,N_3883,N_4426);
nand U9762 (N_9762,N_3341,N_2482);
xnor U9763 (N_9763,N_725,N_4371);
or U9764 (N_9764,N_1705,N_2967);
xnor U9765 (N_9765,N_1616,N_2134);
and U9766 (N_9766,N_981,N_4261);
or U9767 (N_9767,N_2694,N_1226);
and U9768 (N_9768,N_4947,N_3804);
or U9769 (N_9769,N_93,N_1930);
and U9770 (N_9770,N_1991,N_3354);
nand U9771 (N_9771,N_2043,N_4132);
nand U9772 (N_9772,N_1715,N_3314);
or U9773 (N_9773,N_3811,N_2753);
nand U9774 (N_9774,N_2927,N_2163);
or U9775 (N_9775,N_3926,N_281);
or U9776 (N_9776,N_3217,N_3080);
nor U9777 (N_9777,N_2631,N_2477);
xor U9778 (N_9778,N_740,N_2183);
and U9779 (N_9779,N_3196,N_2532);
xor U9780 (N_9780,N_4544,N_2867);
xnor U9781 (N_9781,N_399,N_218);
or U9782 (N_9782,N_2305,N_2570);
nor U9783 (N_9783,N_2314,N_4754);
or U9784 (N_9784,N_3855,N_321);
xor U9785 (N_9785,N_4930,N_864);
and U9786 (N_9786,N_4655,N_1459);
or U9787 (N_9787,N_562,N_277);
nor U9788 (N_9788,N_559,N_4816);
or U9789 (N_9789,N_3974,N_4470);
xor U9790 (N_9790,N_793,N_4692);
nor U9791 (N_9791,N_3325,N_4271);
xor U9792 (N_9792,N_4757,N_4107);
xnor U9793 (N_9793,N_2193,N_908);
nor U9794 (N_9794,N_1746,N_1731);
xor U9795 (N_9795,N_2130,N_2541);
and U9796 (N_9796,N_2231,N_3967);
nand U9797 (N_9797,N_1270,N_393);
xor U9798 (N_9798,N_113,N_2007);
or U9799 (N_9799,N_3443,N_572);
or U9800 (N_9800,N_2195,N_4478);
xnor U9801 (N_9801,N_4382,N_4535);
nand U9802 (N_9802,N_504,N_2083);
nor U9803 (N_9803,N_4531,N_3228);
nor U9804 (N_9804,N_2140,N_3252);
xnor U9805 (N_9805,N_2969,N_2725);
or U9806 (N_9806,N_202,N_782);
xnor U9807 (N_9807,N_3608,N_4149);
nor U9808 (N_9808,N_1384,N_4624);
xor U9809 (N_9809,N_4483,N_3823);
nand U9810 (N_9810,N_1225,N_2973);
or U9811 (N_9811,N_605,N_3661);
xor U9812 (N_9812,N_3570,N_3457);
xnor U9813 (N_9813,N_4078,N_340);
nand U9814 (N_9814,N_3141,N_4823);
nor U9815 (N_9815,N_3310,N_2938);
or U9816 (N_9816,N_399,N_826);
nor U9817 (N_9817,N_3656,N_4631);
nor U9818 (N_9818,N_4382,N_4137);
or U9819 (N_9819,N_4317,N_1578);
and U9820 (N_9820,N_2871,N_434);
xnor U9821 (N_9821,N_1256,N_3552);
nand U9822 (N_9822,N_4433,N_2846);
xor U9823 (N_9823,N_2358,N_4127);
or U9824 (N_9824,N_1043,N_1248);
or U9825 (N_9825,N_4402,N_915);
xor U9826 (N_9826,N_4667,N_2300);
xnor U9827 (N_9827,N_4275,N_2324);
xnor U9828 (N_9828,N_4235,N_1225);
nor U9829 (N_9829,N_3054,N_3854);
or U9830 (N_9830,N_4125,N_4246);
nor U9831 (N_9831,N_1527,N_611);
nand U9832 (N_9832,N_827,N_98);
and U9833 (N_9833,N_4963,N_1711);
nand U9834 (N_9834,N_4735,N_1040);
or U9835 (N_9835,N_2973,N_70);
nand U9836 (N_9836,N_933,N_4352);
or U9837 (N_9837,N_1266,N_1546);
nand U9838 (N_9838,N_1617,N_1282);
or U9839 (N_9839,N_4691,N_593);
and U9840 (N_9840,N_2550,N_115);
and U9841 (N_9841,N_3499,N_4964);
or U9842 (N_9842,N_4115,N_3425);
or U9843 (N_9843,N_3307,N_4408);
xnor U9844 (N_9844,N_2309,N_3700);
nor U9845 (N_9845,N_4260,N_4363);
xnor U9846 (N_9846,N_2809,N_2421);
nor U9847 (N_9847,N_2439,N_1942);
nor U9848 (N_9848,N_1223,N_1233);
and U9849 (N_9849,N_477,N_749);
and U9850 (N_9850,N_2489,N_2025);
xnor U9851 (N_9851,N_2318,N_2311);
nor U9852 (N_9852,N_4640,N_2224);
nand U9853 (N_9853,N_3939,N_3269);
nand U9854 (N_9854,N_120,N_4987);
nand U9855 (N_9855,N_554,N_3225);
nand U9856 (N_9856,N_4364,N_2959);
nor U9857 (N_9857,N_4923,N_3798);
nor U9858 (N_9858,N_1693,N_1466);
or U9859 (N_9859,N_4309,N_1236);
xnor U9860 (N_9860,N_4416,N_238);
nor U9861 (N_9861,N_2154,N_601);
nand U9862 (N_9862,N_1817,N_477);
nand U9863 (N_9863,N_2277,N_4556);
nor U9864 (N_9864,N_3730,N_1948);
nand U9865 (N_9865,N_2555,N_3406);
nand U9866 (N_9866,N_498,N_1665);
nand U9867 (N_9867,N_4512,N_4982);
or U9868 (N_9868,N_4161,N_2641);
xor U9869 (N_9869,N_3083,N_4362);
or U9870 (N_9870,N_458,N_2340);
xnor U9871 (N_9871,N_668,N_431);
nor U9872 (N_9872,N_4169,N_4815);
and U9873 (N_9873,N_1573,N_4329);
nand U9874 (N_9874,N_3817,N_2983);
nand U9875 (N_9875,N_2827,N_825);
xor U9876 (N_9876,N_94,N_3511);
nand U9877 (N_9877,N_4546,N_33);
or U9878 (N_9878,N_2142,N_631);
and U9879 (N_9879,N_2586,N_2116);
nor U9880 (N_9880,N_1598,N_963);
or U9881 (N_9881,N_10,N_3267);
or U9882 (N_9882,N_2919,N_1770);
or U9883 (N_9883,N_4782,N_928);
or U9884 (N_9884,N_1394,N_834);
or U9885 (N_9885,N_3692,N_2999);
nand U9886 (N_9886,N_2966,N_261);
and U9887 (N_9887,N_82,N_4177);
xnor U9888 (N_9888,N_2334,N_2779);
and U9889 (N_9889,N_2851,N_992);
nor U9890 (N_9890,N_4865,N_3931);
nor U9891 (N_9891,N_2877,N_3522);
nand U9892 (N_9892,N_4740,N_2243);
nand U9893 (N_9893,N_499,N_1117);
and U9894 (N_9894,N_1912,N_157);
nand U9895 (N_9895,N_1193,N_4312);
nor U9896 (N_9896,N_1425,N_4585);
xor U9897 (N_9897,N_27,N_566);
xnor U9898 (N_9898,N_2559,N_647);
xnor U9899 (N_9899,N_3024,N_44);
nor U9900 (N_9900,N_4895,N_1186);
and U9901 (N_9901,N_918,N_4530);
and U9902 (N_9902,N_838,N_2925);
or U9903 (N_9903,N_2643,N_549);
or U9904 (N_9904,N_2341,N_432);
or U9905 (N_9905,N_848,N_2845);
nor U9906 (N_9906,N_2845,N_4292);
and U9907 (N_9907,N_4387,N_1220);
and U9908 (N_9908,N_2547,N_1300);
and U9909 (N_9909,N_845,N_2094);
or U9910 (N_9910,N_2935,N_2586);
xnor U9911 (N_9911,N_2783,N_85);
and U9912 (N_9912,N_802,N_1200);
and U9913 (N_9913,N_1919,N_3310);
and U9914 (N_9914,N_1152,N_1822);
xor U9915 (N_9915,N_3144,N_362);
xnor U9916 (N_9916,N_3755,N_1726);
nor U9917 (N_9917,N_4248,N_685);
nor U9918 (N_9918,N_4209,N_1092);
and U9919 (N_9919,N_2886,N_4598);
nor U9920 (N_9920,N_2549,N_4529);
nor U9921 (N_9921,N_1513,N_4722);
xor U9922 (N_9922,N_4993,N_4829);
or U9923 (N_9923,N_2858,N_166);
and U9924 (N_9924,N_2769,N_57);
nand U9925 (N_9925,N_4629,N_4721);
nand U9926 (N_9926,N_344,N_3759);
nand U9927 (N_9927,N_1251,N_487);
nand U9928 (N_9928,N_2253,N_3185);
nor U9929 (N_9929,N_1393,N_2215);
nand U9930 (N_9930,N_397,N_2242);
nand U9931 (N_9931,N_2219,N_1500);
nand U9932 (N_9932,N_4665,N_1970);
and U9933 (N_9933,N_900,N_3894);
or U9934 (N_9934,N_3891,N_1442);
or U9935 (N_9935,N_4,N_2711);
nor U9936 (N_9936,N_4578,N_4070);
or U9937 (N_9937,N_1246,N_1947);
nand U9938 (N_9938,N_3914,N_4029);
nand U9939 (N_9939,N_820,N_1248);
and U9940 (N_9940,N_3995,N_2466);
nand U9941 (N_9941,N_1196,N_2936);
or U9942 (N_9942,N_96,N_3920);
nor U9943 (N_9943,N_2203,N_1678);
nor U9944 (N_9944,N_3898,N_4791);
and U9945 (N_9945,N_155,N_1331);
nor U9946 (N_9946,N_3758,N_2574);
nand U9947 (N_9947,N_2005,N_1474);
xnor U9948 (N_9948,N_115,N_446);
nor U9949 (N_9949,N_3554,N_1169);
xnor U9950 (N_9950,N_961,N_230);
xnor U9951 (N_9951,N_2808,N_1156);
or U9952 (N_9952,N_4438,N_3315);
or U9953 (N_9953,N_3580,N_2854);
xnor U9954 (N_9954,N_3291,N_2204);
nor U9955 (N_9955,N_1354,N_4712);
nand U9956 (N_9956,N_1302,N_1725);
or U9957 (N_9957,N_1678,N_4753);
nand U9958 (N_9958,N_1301,N_4016);
and U9959 (N_9959,N_964,N_2649);
or U9960 (N_9960,N_4745,N_558);
xor U9961 (N_9961,N_1072,N_552);
and U9962 (N_9962,N_2304,N_718);
nor U9963 (N_9963,N_1273,N_1055);
nor U9964 (N_9964,N_3228,N_3361);
nand U9965 (N_9965,N_196,N_3762);
and U9966 (N_9966,N_937,N_4207);
nand U9967 (N_9967,N_3194,N_1043);
nand U9968 (N_9968,N_20,N_1973);
and U9969 (N_9969,N_1940,N_3990);
or U9970 (N_9970,N_3968,N_2589);
nand U9971 (N_9971,N_1667,N_4484);
nand U9972 (N_9972,N_4861,N_806);
nand U9973 (N_9973,N_3596,N_1866);
nor U9974 (N_9974,N_1156,N_1687);
nand U9975 (N_9975,N_641,N_474);
or U9976 (N_9976,N_1088,N_4666);
xor U9977 (N_9977,N_2666,N_3534);
or U9978 (N_9978,N_2356,N_2988);
nor U9979 (N_9979,N_1999,N_1153);
nand U9980 (N_9980,N_181,N_4804);
nand U9981 (N_9981,N_689,N_4249);
xor U9982 (N_9982,N_3253,N_3351);
nand U9983 (N_9983,N_2438,N_4880);
xor U9984 (N_9984,N_1134,N_185);
nand U9985 (N_9985,N_1997,N_425);
nor U9986 (N_9986,N_688,N_4495);
nor U9987 (N_9987,N_4064,N_1993);
or U9988 (N_9988,N_3757,N_2896);
nor U9989 (N_9989,N_1687,N_1957);
and U9990 (N_9990,N_2530,N_3068);
nand U9991 (N_9991,N_2722,N_463);
xor U9992 (N_9992,N_3726,N_3992);
nand U9993 (N_9993,N_3923,N_4754);
or U9994 (N_9994,N_561,N_1058);
and U9995 (N_9995,N_2602,N_3593);
and U9996 (N_9996,N_4570,N_341);
or U9997 (N_9997,N_2656,N_1228);
nor U9998 (N_9998,N_300,N_4281);
nor U9999 (N_9999,N_3446,N_89);
and U10000 (N_10000,N_9182,N_7193);
xnor U10001 (N_10001,N_9860,N_8994);
nor U10002 (N_10002,N_6090,N_8698);
or U10003 (N_10003,N_7097,N_8093);
and U10004 (N_10004,N_7353,N_9708);
or U10005 (N_10005,N_8724,N_5030);
nor U10006 (N_10006,N_5694,N_6410);
nand U10007 (N_10007,N_9630,N_6506);
or U10008 (N_10008,N_7774,N_5750);
and U10009 (N_10009,N_5630,N_6976);
and U10010 (N_10010,N_6863,N_9219);
or U10011 (N_10011,N_7874,N_8842);
xor U10012 (N_10012,N_5318,N_7098);
nor U10013 (N_10013,N_8098,N_7535);
or U10014 (N_10014,N_7767,N_5353);
or U10015 (N_10015,N_5168,N_5032);
nand U10016 (N_10016,N_5818,N_8816);
nor U10017 (N_10017,N_5598,N_6583);
or U10018 (N_10018,N_5913,N_9933);
xnor U10019 (N_10019,N_9442,N_5171);
nor U10020 (N_10020,N_9212,N_6787);
and U10021 (N_10021,N_6276,N_6980);
nand U10022 (N_10022,N_7472,N_8573);
and U10023 (N_10023,N_8380,N_9114);
xor U10024 (N_10024,N_6711,N_8574);
nand U10025 (N_10025,N_7152,N_9908);
and U10026 (N_10026,N_7790,N_6886);
or U10027 (N_10027,N_8596,N_5926);
nor U10028 (N_10028,N_8719,N_5036);
and U10029 (N_10029,N_5385,N_8314);
nor U10030 (N_10030,N_8649,N_8772);
or U10031 (N_10031,N_7748,N_8120);
or U10032 (N_10032,N_9177,N_8915);
xnor U10033 (N_10033,N_5577,N_5535);
or U10034 (N_10034,N_7492,N_7876);
and U10035 (N_10035,N_5065,N_5956);
nor U10036 (N_10036,N_7736,N_5636);
nor U10037 (N_10037,N_5402,N_8088);
or U10038 (N_10038,N_9236,N_8959);
nor U10039 (N_10039,N_7449,N_5780);
and U10040 (N_10040,N_5056,N_5253);
xnor U10041 (N_10041,N_5165,N_6926);
xor U10042 (N_10042,N_9095,N_5914);
nand U10043 (N_10043,N_9365,N_5125);
nand U10044 (N_10044,N_6086,N_7778);
nor U10045 (N_10045,N_5071,N_7336);
and U10046 (N_10046,N_5644,N_5453);
nand U10047 (N_10047,N_7595,N_8067);
nor U10048 (N_10048,N_6057,N_9075);
xor U10049 (N_10049,N_8004,N_6284);
or U10050 (N_10050,N_8256,N_9352);
or U10051 (N_10051,N_8116,N_8722);
and U10052 (N_10052,N_7342,N_7641);
xor U10053 (N_10053,N_9698,N_7265);
nand U10054 (N_10054,N_7697,N_5786);
or U10055 (N_10055,N_7077,N_6330);
nor U10056 (N_10056,N_7993,N_7263);
nor U10057 (N_10057,N_6543,N_9466);
xnor U10058 (N_10058,N_7416,N_9658);
or U10059 (N_10059,N_5518,N_6581);
nor U10060 (N_10060,N_5995,N_7822);
nor U10061 (N_10061,N_5434,N_6887);
and U10062 (N_10062,N_6296,N_9404);
nor U10063 (N_10063,N_5428,N_9391);
or U10064 (N_10064,N_7709,N_9976);
nor U10065 (N_10065,N_5330,N_8893);
nor U10066 (N_10066,N_6142,N_5185);
or U10067 (N_10067,N_5215,N_6434);
or U10068 (N_10068,N_8730,N_7598);
nand U10069 (N_10069,N_5369,N_7232);
nor U10070 (N_10070,N_5025,N_8788);
nand U10071 (N_10071,N_9356,N_5472);
or U10072 (N_10072,N_5564,N_5234);
nor U10073 (N_10073,N_9041,N_8773);
xnor U10074 (N_10074,N_8358,N_8274);
and U10075 (N_10075,N_6352,N_6809);
nand U10076 (N_10076,N_9597,N_7500);
or U10077 (N_10077,N_9227,N_8750);
or U10078 (N_10078,N_7567,N_9646);
and U10079 (N_10079,N_8907,N_8412);
or U10080 (N_10080,N_6587,N_6006);
xnor U10081 (N_10081,N_8237,N_8250);
and U10082 (N_10082,N_9045,N_9047);
xnor U10083 (N_10083,N_9462,N_8972);
and U10084 (N_10084,N_5864,N_6510);
and U10085 (N_10085,N_5389,N_6430);
and U10086 (N_10086,N_9372,N_9131);
xor U10087 (N_10087,N_6579,N_9485);
or U10088 (N_10088,N_8987,N_6946);
and U10089 (N_10089,N_9531,N_9039);
or U10090 (N_10090,N_9617,N_5752);
nand U10091 (N_10091,N_8034,N_7180);
nor U10092 (N_10092,N_8103,N_8621);
nand U10093 (N_10093,N_9011,N_9827);
and U10094 (N_10094,N_6639,N_5695);
nor U10095 (N_10095,N_8762,N_7276);
nor U10096 (N_10096,N_8326,N_8000);
xor U10097 (N_10097,N_7387,N_9984);
and U10098 (N_10098,N_9302,N_7105);
nand U10099 (N_10099,N_9512,N_5210);
nand U10100 (N_10100,N_5593,N_7322);
and U10101 (N_10101,N_6575,N_8674);
xor U10102 (N_10102,N_7292,N_5126);
nand U10103 (N_10103,N_7929,N_9437);
or U10104 (N_10104,N_6677,N_8243);
nor U10105 (N_10105,N_5997,N_6165);
nand U10106 (N_10106,N_8595,N_7884);
or U10107 (N_10107,N_5785,N_6349);
xor U10108 (N_10108,N_9887,N_5287);
xor U10109 (N_10109,N_7286,N_9825);
nand U10110 (N_10110,N_8268,N_5885);
or U10111 (N_10111,N_9754,N_5090);
nor U10112 (N_10112,N_9395,N_9870);
and U10113 (N_10113,N_6236,N_8108);
nand U10114 (N_10114,N_7801,N_8348);
or U10115 (N_10115,N_5658,N_5713);
nand U10116 (N_10116,N_6784,N_8160);
nor U10117 (N_10117,N_5180,N_9059);
nor U10118 (N_10118,N_8017,N_8028);
nand U10119 (N_10119,N_6032,N_5849);
nand U10120 (N_10120,N_6621,N_9405);
and U10121 (N_10121,N_8578,N_9504);
nor U10122 (N_10122,N_8204,N_8803);
or U10123 (N_10123,N_6868,N_8693);
and U10124 (N_10124,N_8001,N_9916);
nor U10125 (N_10125,N_5037,N_9776);
and U10126 (N_10126,N_9930,N_6564);
nand U10127 (N_10127,N_7399,N_5294);
and U10128 (N_10128,N_8132,N_9146);
xnor U10129 (N_10129,N_6785,N_8137);
or U10130 (N_10130,N_8853,N_6951);
nand U10131 (N_10131,N_8196,N_6456);
and U10132 (N_10132,N_9601,N_5272);
nand U10133 (N_10133,N_9559,N_9299);
or U10134 (N_10134,N_5905,N_5595);
and U10135 (N_10135,N_9256,N_9621);
or U10136 (N_10136,N_7448,N_8511);
nand U10137 (N_10137,N_7502,N_9021);
xor U10138 (N_10138,N_8884,N_7957);
nor U10139 (N_10139,N_8325,N_7633);
or U10140 (N_10140,N_6999,N_6527);
nand U10141 (N_10141,N_8520,N_5875);
and U10142 (N_10142,N_8593,N_9018);
nand U10143 (N_10143,N_9517,N_6336);
and U10144 (N_10144,N_7344,N_7084);
nor U10145 (N_10145,N_8230,N_8659);
xnor U10146 (N_10146,N_9833,N_8066);
or U10147 (N_10147,N_5502,N_9838);
or U10148 (N_10148,N_6152,N_7791);
nor U10149 (N_10149,N_5328,N_9062);
nor U10150 (N_10150,N_8537,N_6808);
nand U10151 (N_10151,N_9730,N_9524);
or U10152 (N_10152,N_7427,N_9050);
and U10153 (N_10153,N_9064,N_9202);
nand U10154 (N_10154,N_7946,N_9040);
nand U10155 (N_10155,N_5553,N_5408);
nor U10156 (N_10156,N_6985,N_5541);
nor U10157 (N_10157,N_8423,N_6962);
xor U10158 (N_10158,N_8080,N_7686);
nor U10159 (N_10159,N_8565,N_6744);
xor U10160 (N_10160,N_6553,N_6550);
nand U10161 (N_10161,N_7312,N_9478);
xnor U10162 (N_10162,N_6033,N_7580);
nor U10163 (N_10163,N_9910,N_9259);
or U10164 (N_10164,N_5932,N_7751);
or U10165 (N_10165,N_6747,N_7256);
xor U10166 (N_10166,N_5202,N_8707);
xor U10167 (N_10167,N_6478,N_8272);
nand U10168 (N_10168,N_8921,N_9967);
and U10169 (N_10169,N_5580,N_8214);
or U10170 (N_10170,N_7046,N_8006);
and U10171 (N_10171,N_8126,N_9966);
nor U10172 (N_10172,N_8641,N_9412);
nor U10173 (N_10173,N_7547,N_9544);
xor U10174 (N_10174,N_7906,N_5742);
or U10175 (N_10175,N_5439,N_5018);
nor U10176 (N_10176,N_7779,N_5578);
xor U10177 (N_10177,N_7991,N_7269);
nor U10178 (N_10178,N_5591,N_8322);
nor U10179 (N_10179,N_7316,N_5679);
and U10180 (N_10180,N_6930,N_9238);
nor U10181 (N_10181,N_7786,N_5231);
or U10182 (N_10182,N_8181,N_9164);
or U10183 (N_10183,N_7446,N_7585);
xor U10184 (N_10184,N_7123,N_8530);
nand U10185 (N_10185,N_6728,N_9433);
xor U10186 (N_10186,N_5829,N_9648);
nor U10187 (N_10187,N_8435,N_8642);
xor U10188 (N_10188,N_9837,N_6634);
and U10189 (N_10189,N_7627,N_8880);
xnor U10190 (N_10190,N_8540,N_8118);
nand U10191 (N_10191,N_9266,N_5496);
or U10192 (N_10192,N_7341,N_9510);
xor U10193 (N_10193,N_6188,N_5664);
xor U10194 (N_10194,N_7985,N_5170);
xnor U10195 (N_10195,N_5371,N_9168);
and U10196 (N_10196,N_5384,N_5311);
nor U10197 (N_10197,N_9798,N_9420);
nor U10198 (N_10198,N_9906,N_9361);
nand U10199 (N_10199,N_7209,N_8763);
nor U10200 (N_10200,N_5506,N_9201);
xor U10201 (N_10201,N_5226,N_6977);
or U10202 (N_10202,N_5850,N_9226);
and U10203 (N_10203,N_9211,N_9281);
xor U10204 (N_10204,N_7015,N_6753);
xnor U10205 (N_10205,N_7293,N_6066);
or U10206 (N_10206,N_9743,N_5859);
and U10207 (N_10207,N_7240,N_6451);
xnor U10208 (N_10208,N_8896,N_5024);
and U10209 (N_10209,N_6338,N_6323);
nor U10210 (N_10210,N_8532,N_9096);
nor U10211 (N_10211,N_5620,N_6242);
nor U10212 (N_10212,N_9812,N_6221);
nor U10213 (N_10213,N_5298,N_8462);
and U10214 (N_10214,N_5604,N_5751);
nor U10215 (N_10215,N_7719,N_9272);
nor U10216 (N_10216,N_8253,N_9962);
nor U10217 (N_10217,N_7470,N_8504);
xor U10218 (N_10218,N_6866,N_9098);
or U10219 (N_10219,N_7150,N_9097);
xor U10220 (N_10220,N_5055,N_9101);
and U10221 (N_10221,N_9348,N_6992);
xnor U10222 (N_10222,N_6883,N_5728);
nand U10223 (N_10223,N_8170,N_9473);
nand U10224 (N_10224,N_9756,N_6523);
nor U10225 (N_10225,N_7082,N_6148);
nand U10226 (N_10226,N_6648,N_7587);
or U10227 (N_10227,N_7700,N_9513);
and U10228 (N_10228,N_5201,N_7408);
xnor U10229 (N_10229,N_8023,N_7808);
xnor U10230 (N_10230,N_9959,N_9858);
nand U10231 (N_10231,N_6849,N_5974);
or U10232 (N_10232,N_7760,N_6731);
xnor U10233 (N_10233,N_8197,N_8426);
xor U10234 (N_10234,N_7441,N_6365);
xnor U10235 (N_10235,N_9616,N_7166);
xor U10236 (N_10236,N_8644,N_8517);
and U10237 (N_10237,N_9100,N_8374);
xnor U10238 (N_10238,N_7029,N_9618);
xnor U10239 (N_10239,N_9042,N_6015);
nand U10240 (N_10240,N_7707,N_8536);
xnor U10241 (N_10241,N_5810,N_7729);
nand U10242 (N_10242,N_9195,N_5808);
or U10243 (N_10243,N_9083,N_6052);
or U10244 (N_10244,N_9336,N_8922);
xor U10245 (N_10245,N_8456,N_9613);
and U10246 (N_10246,N_7458,N_6439);
and U10247 (N_10247,N_6133,N_7924);
xor U10248 (N_10248,N_9492,N_6822);
nand U10249 (N_10249,N_5590,N_6697);
or U10250 (N_10250,N_9581,N_7372);
nand U10251 (N_10251,N_7157,N_9903);
nand U10252 (N_10252,N_9203,N_8252);
nor U10253 (N_10253,N_5207,N_7583);
or U10254 (N_10254,N_9566,N_9475);
or U10255 (N_10255,N_9922,N_8282);
nand U10256 (N_10256,N_7664,N_8737);
nor U10257 (N_10257,N_8012,N_8809);
nor U10258 (N_10258,N_5793,N_5080);
nor U10259 (N_10259,N_5661,N_6620);
nand U10260 (N_10260,N_9242,N_7491);
xnor U10261 (N_10261,N_5783,N_5657);
nor U10262 (N_10262,N_9969,N_9483);
nor U10263 (N_10263,N_7056,N_9895);
nand U10264 (N_10264,N_8557,N_7309);
and U10265 (N_10265,N_7167,N_9555);
xor U10266 (N_10266,N_8923,N_8223);
and U10267 (N_10267,N_7154,N_7266);
and U10268 (N_10268,N_5817,N_9243);
nor U10269 (N_10269,N_8311,N_5895);
xor U10270 (N_10270,N_6661,N_7969);
nor U10271 (N_10271,N_8710,N_9204);
and U10272 (N_10272,N_7691,N_8671);
and U10273 (N_10273,N_9993,N_7188);
and U10274 (N_10274,N_7165,N_7435);
xnor U10275 (N_10275,N_9148,N_8136);
and U10276 (N_10276,N_7572,N_7880);
or U10277 (N_10277,N_6315,N_9593);
nor U10278 (N_10278,N_6271,N_5978);
nor U10279 (N_10279,N_7813,N_8075);
and U10280 (N_10280,N_8634,N_8900);
xnor U10281 (N_10281,N_5331,N_9332);
nand U10282 (N_10282,N_8777,N_9161);
and U10283 (N_10283,N_8944,N_6720);
or U10284 (N_10284,N_7307,N_6791);
nor U10285 (N_10285,N_7130,N_5976);
nand U10286 (N_10286,N_8433,N_8432);
nand U10287 (N_10287,N_6125,N_5455);
nor U10288 (N_10288,N_6508,N_9907);
and U10289 (N_10289,N_8560,N_9255);
or U10290 (N_10290,N_6282,N_6056);
and U10291 (N_10291,N_6975,N_6937);
and U10292 (N_10292,N_8344,N_8185);
nand U10293 (N_10293,N_9803,N_8062);
nor U10294 (N_10294,N_5006,N_7800);
nor U10295 (N_10295,N_8400,N_5345);
nor U10296 (N_10296,N_6905,N_7228);
nor U10297 (N_10297,N_7501,N_7296);
nand U10298 (N_10298,N_8631,N_7932);
nand U10299 (N_10299,N_6774,N_6568);
and U10300 (N_10300,N_6150,N_8375);
nand U10301 (N_10301,N_7163,N_9821);
or U10302 (N_10302,N_9123,N_6041);
nand U10303 (N_10303,N_5368,N_8270);
xor U10304 (N_10304,N_7095,N_5592);
xnor U10305 (N_10305,N_6989,N_5915);
or U10306 (N_10306,N_7835,N_7783);
or U10307 (N_10307,N_6021,N_6162);
nor U10308 (N_10308,N_7184,N_6708);
or U10309 (N_10309,N_9024,N_6346);
nor U10310 (N_10310,N_9179,N_9487);
nand U10311 (N_10311,N_5473,N_5939);
or U10312 (N_10312,N_9126,N_8962);
and U10313 (N_10313,N_5745,N_8757);
and U10314 (N_10314,N_7814,N_6763);
and U10315 (N_10315,N_6812,N_5460);
and U10316 (N_10316,N_6299,N_6403);
nor U10317 (N_10317,N_5306,N_8904);
nor U10318 (N_10318,N_5557,N_7350);
nor U10319 (N_10319,N_8917,N_7909);
nand U10320 (N_10320,N_8011,N_9809);
xor U10321 (N_10321,N_8948,N_7087);
nor U10322 (N_10322,N_8863,N_9106);
or U10323 (N_10323,N_7635,N_8657);
nor U10324 (N_10324,N_5175,N_6357);
xor U10325 (N_10325,N_6144,N_5527);
and U10326 (N_10326,N_9304,N_6795);
and U10327 (N_10327,N_9188,N_8971);
nand U10328 (N_10328,N_8830,N_8060);
nor U10329 (N_10329,N_8209,N_5393);
or U10330 (N_10330,N_6574,N_6079);
xnor U10331 (N_10331,N_5756,N_5250);
or U10332 (N_10332,N_7857,N_6860);
nand U10333 (N_10333,N_7379,N_5585);
and U10334 (N_10334,N_6804,N_9122);
and U10335 (N_10335,N_6420,N_5089);
nand U10336 (N_10336,N_9783,N_7223);
nor U10337 (N_10337,N_8302,N_5243);
nor U10338 (N_10338,N_6504,N_5245);
xor U10339 (N_10339,N_7190,N_9217);
nand U10340 (N_10340,N_7085,N_7531);
nor U10341 (N_10341,N_7608,N_5899);
xnor U10342 (N_10342,N_5269,N_9878);
or U10343 (N_10343,N_7904,N_5217);
nand U10344 (N_10344,N_7925,N_6379);
nor U10345 (N_10345,N_7144,N_8133);
nand U10346 (N_10346,N_5836,N_7413);
nand U10347 (N_10347,N_6754,N_5383);
and U10348 (N_10348,N_6654,N_5765);
xor U10349 (N_10349,N_5327,N_5004);
nand U10350 (N_10350,N_7395,N_8129);
and U10351 (N_10351,N_7033,N_5696);
and U10352 (N_10352,N_5888,N_5156);
nand U10353 (N_10353,N_6054,N_5626);
and U10354 (N_10354,N_6279,N_5601);
nand U10355 (N_10355,N_5826,N_7812);
nor U10356 (N_10356,N_7628,N_7770);
or U10357 (N_10357,N_5929,N_7078);
nand U10358 (N_10358,N_5998,N_6442);
and U10359 (N_10359,N_6094,N_5088);
or U10360 (N_10360,N_6676,N_9841);
xnor U10361 (N_10361,N_7114,N_9789);
xnor U10362 (N_10362,N_5367,N_8381);
xnor U10363 (N_10363,N_9094,N_5319);
xor U10364 (N_10364,N_8384,N_8403);
nand U10365 (N_10365,N_9093,N_7680);
and U10366 (N_10366,N_5757,N_7565);
or U10367 (N_10367,N_9955,N_7644);
nand U10368 (N_10368,N_9897,N_6828);
and U10369 (N_10369,N_6716,N_5329);
nand U10370 (N_10370,N_9500,N_6996);
and U10371 (N_10371,N_8482,N_7047);
and U10372 (N_10372,N_9713,N_6653);
or U10373 (N_10373,N_6727,N_6803);
nor U10374 (N_10374,N_7933,N_8643);
and U10375 (N_10375,N_6684,N_6360);
and U10376 (N_10376,N_6331,N_9873);
and U10377 (N_10377,N_6907,N_9479);
nand U10378 (N_10378,N_7001,N_5407);
or U10379 (N_10379,N_5680,N_6594);
nor U10380 (N_10380,N_5183,N_5724);
xor U10381 (N_10381,N_9773,N_9808);
nor U10382 (N_10382,N_9975,N_8691);
xor U10383 (N_10383,N_8798,N_8056);
xor U10384 (N_10384,N_8989,N_8814);
xnor U10385 (N_10385,N_8254,N_6370);
or U10386 (N_10386,N_8488,N_6069);
or U10387 (N_10387,N_5164,N_7410);
and U10388 (N_10388,N_6465,N_6561);
and U10389 (N_10389,N_5641,N_5001);
or U10390 (N_10390,N_5034,N_6705);
xor U10391 (N_10391,N_9419,N_9885);
nand U10392 (N_10392,N_8609,N_8276);
xnor U10393 (N_10393,N_8501,N_9354);
nor U10394 (N_10394,N_5952,N_7558);
xnor U10395 (N_10395,N_9175,N_8470);
or U10396 (N_10396,N_7231,N_9430);
and U10397 (N_10397,N_6721,N_9797);
or U10398 (N_10398,N_8594,N_5377);
nor U10399 (N_10399,N_8387,N_9722);
nor U10400 (N_10400,N_9664,N_9516);
nand U10401 (N_10401,N_6990,N_7378);
xnor U10402 (N_10402,N_7109,N_9127);
nor U10403 (N_10403,N_5878,N_8873);
or U10404 (N_10404,N_8357,N_7230);
xnor U10405 (N_10405,N_9252,N_7026);
nor U10406 (N_10406,N_6958,N_5147);
and U10407 (N_10407,N_5683,N_8548);
xnor U10408 (N_10408,N_7170,N_6179);
and U10409 (N_10409,N_5360,N_9382);
nand U10410 (N_10410,N_6590,N_5275);
xnor U10411 (N_10411,N_6232,N_8109);
or U10412 (N_10412,N_7949,N_6986);
nor U10413 (N_10413,N_5011,N_5971);
xnor U10414 (N_10414,N_6843,N_7043);
and U10415 (N_10415,N_5127,N_5283);
nand U10416 (N_10416,N_9029,N_9518);
xor U10417 (N_10417,N_7058,N_8717);
or U10418 (N_10418,N_8284,N_7377);
and U10419 (N_10419,N_6807,N_7164);
and U10420 (N_10420,N_9163,N_6898);
nor U10421 (N_10421,N_5337,N_9857);
or U10422 (N_10422,N_8937,N_6153);
or U10423 (N_10423,N_7299,N_9685);
nor U10424 (N_10424,N_9153,N_8031);
nor U10425 (N_10425,N_6577,N_7022);
nor U10426 (N_10426,N_6901,N_9786);
xnor U10427 (N_10427,N_8319,N_7131);
nor U10428 (N_10428,N_5802,N_6806);
and U10429 (N_10429,N_9181,N_8114);
xor U10430 (N_10430,N_9245,N_7529);
and U10431 (N_10431,N_8844,N_6637);
nor U10432 (N_10432,N_6224,N_6083);
and U10433 (N_10433,N_6077,N_7673);
nor U10434 (N_10434,N_7636,N_5975);
nand U10435 (N_10435,N_5312,N_7571);
nand U10436 (N_10436,N_9089,N_5300);
xor U10437 (N_10437,N_9457,N_5159);
or U10438 (N_10438,N_5520,N_5775);
xnor U10439 (N_10439,N_6521,N_8484);
and U10440 (N_10440,N_6319,N_7390);
xnor U10441 (N_10441,N_8756,N_9687);
or U10442 (N_10442,N_6948,N_9138);
nand U10443 (N_10443,N_5840,N_5709);
nor U10444 (N_10444,N_5012,N_9541);
nor U10445 (N_10445,N_6136,N_8113);
and U10446 (N_10446,N_9896,N_8094);
nor U10447 (N_10447,N_6546,N_7310);
nor U10448 (N_10448,N_7036,N_9452);
nor U10449 (N_10449,N_9936,N_9811);
nand U10450 (N_10450,N_6961,N_7749);
or U10451 (N_10451,N_5264,N_7384);
xor U10452 (N_10452,N_5687,N_8019);
and U10453 (N_10453,N_6337,N_9189);
nor U10454 (N_10454,N_9961,N_6555);
and U10455 (N_10455,N_6857,N_7692);
nor U10456 (N_10456,N_5744,N_8350);
or U10457 (N_10457,N_5040,N_9794);
or U10458 (N_10458,N_8207,N_6757);
nor U10459 (N_10459,N_9710,N_5076);
nor U10460 (N_10460,N_5419,N_6364);
nor U10461 (N_10461,N_7337,N_8163);
and U10462 (N_10462,N_8390,N_9052);
and U10463 (N_10463,N_9494,N_8810);
nor U10464 (N_10464,N_6191,N_7126);
xnor U10465 (N_10465,N_9261,N_6115);
xnor U10466 (N_10466,N_8526,N_6818);
and U10467 (N_10467,N_9944,N_8224);
and U10468 (N_10468,N_9180,N_7096);
or U10469 (N_10469,N_8580,N_6036);
xnor U10470 (N_10470,N_8852,N_9902);
nand U10471 (N_10471,N_9271,N_6397);
xor U10472 (N_10472,N_8147,N_5440);
or U10473 (N_10473,N_8575,N_7249);
nor U10474 (N_10474,N_9805,N_5705);
nor U10475 (N_10475,N_8891,N_5602);
nor U10476 (N_10476,N_6794,N_9628);
nand U10477 (N_10477,N_5618,N_5957);
xor U10478 (N_10478,N_8257,N_8910);
or U10479 (N_10479,N_8813,N_5124);
and U10480 (N_10480,N_7329,N_5152);
or U10481 (N_10481,N_6207,N_7267);
nand U10482 (N_10482,N_9288,N_5522);
xor U10483 (N_10483,N_7903,N_6674);
and U10484 (N_10484,N_7679,N_9254);
nor U10485 (N_10485,N_9577,N_6585);
nor U10486 (N_10486,N_6802,N_5133);
or U10487 (N_10487,N_9265,N_6699);
or U10488 (N_10488,N_5853,N_9366);
nor U10489 (N_10489,N_9576,N_6245);
xnor U10490 (N_10490,N_7678,N_6969);
and U10491 (N_10491,N_8812,N_6342);
or U10492 (N_10492,N_7151,N_6702);
nor U10493 (N_10493,N_6216,N_6378);
nor U10494 (N_10494,N_8155,N_8329);
nand U10495 (N_10495,N_7260,N_6117);
nand U10496 (N_10496,N_9550,N_9362);
and U10497 (N_10497,N_5246,N_7479);
and U10498 (N_10498,N_5281,N_9057);
xnor U10499 (N_10499,N_9495,N_7672);
or U10500 (N_10500,N_6089,N_5515);
or U10501 (N_10501,N_6058,N_9842);
nand U10502 (N_10502,N_7326,N_6396);
nor U10503 (N_10503,N_5471,N_5596);
xnor U10504 (N_10504,N_9184,N_5890);
xor U10505 (N_10505,N_8571,N_8205);
and U10506 (N_10506,N_6020,N_6790);
or U10507 (N_10507,N_9739,N_9234);
nor U10508 (N_10508,N_9546,N_9166);
and U10509 (N_10509,N_9926,N_8452);
nand U10510 (N_10510,N_6260,N_6124);
or U10511 (N_10511,N_5928,N_9696);
xnor U10512 (N_10512,N_5736,N_6250);
and U10513 (N_10513,N_6797,N_8027);
nor U10514 (N_10514,N_5700,N_8766);
xnor U10515 (N_10515,N_6773,N_6931);
xor U10516 (N_10516,N_5721,N_6668);
nor U10517 (N_10517,N_5174,N_8178);
and U10518 (N_10518,N_8780,N_6895);
and U10519 (N_10519,N_9568,N_8854);
xnor U10520 (N_10520,N_7233,N_7784);
xor U10521 (N_10521,N_8799,N_8899);
nor U10522 (N_10522,N_8729,N_8183);
or U10523 (N_10523,N_5588,N_7219);
or U10524 (N_10524,N_9570,N_5042);
nand U10525 (N_10525,N_8622,N_8686);
nand U10526 (N_10526,N_7039,N_5392);
nand U10527 (N_10527,N_9898,N_9250);
xnor U10528 (N_10528,N_8601,N_5186);
nor U10529 (N_10529,N_7469,N_7609);
xor U10530 (N_10530,N_5203,N_9737);
or U10531 (N_10531,N_5852,N_8587);
or U10532 (N_10532,N_8886,N_8916);
nand U10533 (N_10533,N_8267,N_9591);
and U10534 (N_10534,N_8738,N_9493);
and U10535 (N_10535,N_9191,N_8468);
nor U10536 (N_10536,N_8555,N_8275);
nand U10537 (N_10537,N_5136,N_8656);
xnor U10538 (N_10538,N_8365,N_5413);
nand U10539 (N_10539,N_9080,N_8882);
nor U10540 (N_10540,N_5148,N_6468);
or U10541 (N_10541,N_5537,N_7334);
nor U10542 (N_10542,N_7509,N_6760);
nand U10543 (N_10543,N_8503,N_7365);
nand U10544 (N_10544,N_6729,N_6043);
and U10545 (N_10545,N_7002,N_8592);
nor U10546 (N_10546,N_7145,N_8797);
and U10547 (N_10547,N_6602,N_5454);
and U10548 (N_10548,N_9140,N_7229);
nand U10549 (N_10549,N_5629,N_9178);
xnor U10550 (N_10550,N_9197,N_5674);
and U10551 (N_10551,N_5121,N_9567);
nor U10552 (N_10552,N_6252,N_6334);
nand U10553 (N_10553,N_8032,N_7092);
or U10554 (N_10554,N_8743,N_8124);
xor U10555 (N_10555,N_9160,N_7194);
xnor U10556 (N_10556,N_6861,N_7281);
xnor U10557 (N_10557,N_6481,N_8958);
xnor U10558 (N_10558,N_7238,N_5923);
and U10559 (N_10559,N_7422,N_7147);
or U10560 (N_10560,N_9751,N_7351);
xor U10561 (N_10561,N_5397,N_8632);
xor U10562 (N_10562,N_9706,N_7206);
or U10563 (N_10563,N_7425,N_8317);
xor U10564 (N_10564,N_7507,N_9914);
or U10565 (N_10565,N_7136,N_9767);
xor U10566 (N_10566,N_8991,N_9012);
nor U10567 (N_10567,N_5375,N_9644);
or U10568 (N_10568,N_8874,N_7769);
xnor U10569 (N_10569,N_8258,N_6914);
nand U10570 (N_10570,N_5359,N_8059);
xnor U10571 (N_10571,N_7785,N_7037);
nor U10572 (N_10572,N_7703,N_8924);
xnor U10573 (N_10573,N_5204,N_9680);
and U10574 (N_10574,N_8083,N_7918);
nand U10575 (N_10575,N_8623,N_5943);
and U10576 (N_10576,N_8553,N_9322);
and U10577 (N_10577,N_6302,N_7020);
or U10578 (N_10578,N_6655,N_9919);
and U10579 (N_10579,N_5142,N_8668);
xor U10580 (N_10580,N_5466,N_6904);
or U10581 (N_10581,N_7948,N_5884);
xnor U10582 (N_10582,N_8550,N_7288);
nor U10583 (N_10583,N_8391,N_8127);
nor U10584 (N_10584,N_6925,N_7772);
nand U10585 (N_10585,N_7964,N_5342);
or U10586 (N_10586,N_9370,N_7839);
nand U10587 (N_10587,N_7573,N_9766);
nand U10588 (N_10588,N_7004,N_6464);
nor U10589 (N_10589,N_9571,N_5326);
nand U10590 (N_10590,N_7295,N_8694);
or U10591 (N_10591,N_5809,N_5449);
nor U10592 (N_10592,N_5739,N_8527);
nor U10593 (N_10593,N_5340,N_5967);
xor U10594 (N_10594,N_8008,N_6308);
xor U10595 (N_10595,N_7665,N_7423);
nand U10596 (N_10596,N_8184,N_9724);
and U10597 (N_10597,N_8747,N_6921);
or U10598 (N_10598,N_8786,N_8347);
nor U10599 (N_10599,N_7889,N_8042);
nand U10600 (N_10600,N_9393,N_5430);
and U10601 (N_10601,N_9258,N_5417);
nand U10602 (N_10602,N_6896,N_5289);
and U10603 (N_10603,N_7603,N_7073);
nor U10604 (N_10604,N_7428,N_6567);
nand U10605 (N_10605,N_8770,N_9686);
nand U10606 (N_10606,N_9744,N_5020);
and U10607 (N_10607,N_7466,N_6423);
and U10608 (N_10608,N_8529,N_7156);
nand U10609 (N_10609,N_7647,N_8140);
or U10610 (N_10610,N_9102,N_8428);
nand U10611 (N_10611,N_6301,N_6709);
and U10612 (N_10612,N_9295,N_5224);
and U10613 (N_10613,N_7622,N_6678);
or U10614 (N_10614,N_9929,N_6325);
nand U10615 (N_10615,N_6394,N_5077);
nor U10616 (N_10616,N_9283,N_9727);
and U10617 (N_10617,N_9788,N_9241);
or U10618 (N_10618,N_9409,N_6368);
nor U10619 (N_10619,N_5619,N_7420);
nand U10620 (N_10620,N_5665,N_5053);
or U10621 (N_10621,N_7526,N_7725);
and U10622 (N_10622,N_8605,N_9427);
and U10623 (N_10623,N_7090,N_5351);
nor U10624 (N_10624,N_5084,N_9912);
xor U10625 (N_10625,N_5758,N_7134);
and U10626 (N_10626,N_6872,N_7768);
nor U10627 (N_10627,N_6775,N_7186);
xnor U10628 (N_10628,N_6435,N_8281);
or U10629 (N_10629,N_6122,N_6833);
nand U10630 (N_10630,N_8486,N_7120);
nor U10631 (N_10631,N_6053,N_6457);
nand U10632 (N_10632,N_6328,N_6288);
and U10633 (N_10633,N_5867,N_9364);
or U10634 (N_10634,N_8279,N_8897);
nor U10635 (N_10635,N_9522,N_6858);
nand U10636 (N_10636,N_5902,N_6453);
nor U10637 (N_10637,N_9121,N_9679);
nand U10638 (N_10638,N_9545,N_9221);
xnor U10639 (N_10639,N_8521,N_8968);
xnor U10640 (N_10640,N_9677,N_8417);
and U10641 (N_10641,N_7205,N_6950);
xor U10642 (N_10642,N_9958,N_6826);
and U10643 (N_10643,N_9028,N_8036);
xnor U10644 (N_10644,N_7559,N_9987);
nand U10645 (N_10645,N_9306,N_7273);
nand U10646 (N_10646,N_9904,N_7275);
or U10647 (N_10647,N_6470,N_8611);
nand U10648 (N_10648,N_9355,N_7331);
or U10649 (N_10649,N_9455,N_7970);
xor U10650 (N_10650,N_5343,N_9999);
or U10651 (N_10651,N_6789,N_5333);
or U10652 (N_10652,N_8070,N_9249);
and U10653 (N_10653,N_9503,N_9726);
xor U10654 (N_10654,N_6387,N_5247);
or U10655 (N_10655,N_7747,N_6092);
nand U10656 (N_10656,N_8259,N_8202);
xnor U10657 (N_10657,N_7129,N_7108);
xor U10658 (N_10658,N_5963,N_6862);
nand U10659 (N_10659,N_8919,N_8159);
and U10660 (N_10660,N_6599,N_8078);
and U10661 (N_10661,N_8655,N_8356);
nand U10662 (N_10662,N_8260,N_7174);
nand U10663 (N_10663,N_5458,N_8176);
nand U10664 (N_10664,N_6326,N_5304);
nor U10665 (N_10665,N_7439,N_9782);
nor U10666 (N_10666,N_6672,N_6151);
and U10667 (N_10667,N_7782,N_5871);
and U10668 (N_10668,N_7728,N_5094);
and U10669 (N_10669,N_7837,N_8003);
and U10670 (N_10670,N_5816,N_8542);
nor U10671 (N_10671,N_5092,N_9596);
or U10672 (N_10672,N_9777,N_8827);
and U10673 (N_10673,N_8463,N_9632);
or U10674 (N_10674,N_5767,N_7214);
and U10675 (N_10675,N_5624,N_9051);
nand U10676 (N_10676,N_7542,N_5941);
xnor U10677 (N_10677,N_6204,N_6452);
nand U10678 (N_10678,N_7168,N_8065);
nor U10679 (N_10679,N_8878,N_5822);
nor U10680 (N_10680,N_5769,N_5819);
xnor U10681 (N_10681,N_5107,N_5373);
or U10682 (N_10682,N_9997,N_9351);
and U10683 (N_10683,N_9032,N_5847);
nor U10684 (N_10684,N_5669,N_8861);
nand U10685 (N_10685,N_5116,N_5008);
nor U10686 (N_10686,N_5480,N_6966);
or U10687 (N_10687,N_6321,N_7733);
or U10688 (N_10688,N_5937,N_8226);
nand U10689 (N_10689,N_5313,N_9893);
nand U10690 (N_10690,N_9714,N_7886);
nor U10691 (N_10691,N_7057,N_9659);
or U10692 (N_10692,N_7737,N_7667);
nor U10693 (N_10693,N_6289,N_8020);
xnor U10694 (N_10694,N_8685,N_6865);
nor U10695 (N_10695,N_6759,N_9759);
or U10696 (N_10696,N_9066,N_6130);
nor U10697 (N_10697,N_6220,N_5364);
or U10698 (N_10698,N_8338,N_9505);
xnor U10699 (N_10699,N_9931,N_8165);
and U10700 (N_10700,N_6198,N_6884);
nand U10701 (N_10701,N_7781,N_5828);
or U10702 (N_10702,N_5688,N_9871);
xnor U10703 (N_10703,N_7773,N_6519);
xor U10704 (N_10704,N_8726,N_5555);
and U10705 (N_10705,N_6813,N_9169);
xnor U10706 (N_10706,N_9915,N_6174);
and U10707 (N_10707,N_8033,N_6888);
nor U10708 (N_10708,N_7975,N_7766);
or U10709 (N_10709,N_8781,N_8359);
nor U10710 (N_10710,N_8096,N_7346);
nor U10711 (N_10711,N_7332,N_5452);
nand U10712 (N_10712,N_7640,N_8121);
or U10713 (N_10713,N_7135,N_9235);
nand U10714 (N_10714,N_5891,N_6161);
or U10715 (N_10715,N_5365,N_9087);
nand U10716 (N_10716,N_8041,N_7248);
nor U10717 (N_10717,N_5293,N_9027);
and U10718 (N_10718,N_6536,N_6345);
or U10719 (N_10719,N_8602,N_5427);
nor U10720 (N_10720,N_8832,N_8841);
nor U10721 (N_10721,N_8363,N_9538);
and U10722 (N_10722,N_8425,N_6399);
and U10723 (N_10723,N_7451,N_5192);
xnor U10724 (N_10724,N_8335,N_8287);
and U10725 (N_10725,N_6067,N_8934);
nand U10726 (N_10726,N_6262,N_6178);
or U10727 (N_10727,N_9194,N_5132);
and U10728 (N_10728,N_8796,N_8064);
or U10729 (N_10729,N_6320,N_6024);
and U10730 (N_10730,N_9519,N_9852);
and U10731 (N_10731,N_8551,N_9552);
xor U10732 (N_10732,N_7927,N_6606);
and U10733 (N_10733,N_5946,N_8975);
nand U10734 (N_10734,N_5999,N_8408);
nand U10735 (N_10735,N_7431,N_9026);
nor U10736 (N_10736,N_5307,N_9030);
or U10737 (N_10737,N_7817,N_6752);
xnor U10738 (N_10738,N_9623,N_6592);
or U10739 (N_10739,N_7621,N_9270);
and U10740 (N_10740,N_8321,N_6997);
xnor U10741 (N_10741,N_9553,N_5559);
nand U10742 (N_10742,N_9055,N_6380);
nand U10743 (N_10743,N_8157,N_7995);
and U10744 (N_10744,N_7894,N_9344);
nor U10745 (N_10745,N_8288,N_6761);
nor U10746 (N_10746,N_6736,N_6595);
xor U10747 (N_10747,N_9701,N_9770);
and U10748 (N_10748,N_9285,N_9584);
xnor U10749 (N_10749,N_8723,N_9639);
xor U10750 (N_10750,N_8889,N_6683);
or U10751 (N_10751,N_6383,N_5184);
xor U10752 (N_10752,N_5172,N_9237);
nand U10753 (N_10753,N_6428,N_9508);
or U10754 (N_10754,N_5844,N_8188);
and U10755 (N_10755,N_5980,N_5093);
nor U10756 (N_10756,N_5642,N_8353);
nand U10757 (N_10757,N_9711,N_9985);
nand U10758 (N_10758,N_7404,N_6350);
nor U10759 (N_10759,N_9982,N_5542);
xnor U10760 (N_10760,N_5163,N_8111);
and U10761 (N_10761,N_5015,N_7196);
nor U10762 (N_10762,N_5550,N_5344);
and U10763 (N_10763,N_6596,N_8149);
xor U10764 (N_10764,N_5741,N_6934);
and U10765 (N_10765,N_9565,N_8449);
nor U10766 (N_10766,N_9672,N_5917);
nor U10767 (N_10767,N_9866,N_5078);
and U10768 (N_10768,N_5607,N_7869);
nor U10769 (N_10769,N_5066,N_9154);
nand U10770 (N_10770,N_5760,N_8528);
nand U10771 (N_10771,N_7021,N_9839);
xor U10772 (N_10772,N_9823,N_6332);
or U10773 (N_10773,N_7055,N_7411);
xor U10774 (N_10774,N_7675,N_8681);
and U10775 (N_10775,N_7069,N_6016);
and U10776 (N_10776,N_9888,N_7028);
or U10777 (N_10777,N_7270,N_9015);
or U10778 (N_10778,N_9432,N_7328);
nand U10779 (N_10779,N_5706,N_6967);
xor U10780 (N_10780,N_8481,N_9590);
or U10781 (N_10781,N_8999,N_9514);
xor U10782 (N_10782,N_7107,N_6084);
or U10783 (N_10783,N_8351,N_9308);
nor U10784 (N_10784,N_6129,N_6181);
nand U10785 (N_10785,N_6261,N_8499);
xnor U10786 (N_10786,N_7272,N_7549);
or U10787 (N_10787,N_8376,N_7983);
xnor U10788 (N_10788,N_7612,N_8662);
or U10789 (N_10789,N_9377,N_5335);
or U10790 (N_10790,N_8496,N_9115);
nor U10791 (N_10791,N_6235,N_7788);
or U10792 (N_10792,N_8301,N_8245);
nor U10793 (N_10793,N_9425,N_6395);
xnor U10794 (N_10794,N_7634,N_9778);
nor U10795 (N_10795,N_5474,N_9345);
xor U10796 (N_10796,N_5697,N_5111);
and U10797 (N_10797,N_5489,N_5465);
nor U10798 (N_10798,N_9832,N_7841);
and U10799 (N_10799,N_5446,N_7916);
xor U10800 (N_10800,N_6266,N_7899);
xor U10801 (N_10801,N_8782,N_5182);
nand U10802 (N_10802,N_5823,N_8926);
and U10803 (N_10803,N_9521,N_5761);
and U10804 (N_10804,N_8952,N_9631);
or U10805 (N_10805,N_6793,N_9334);
and U10806 (N_10806,N_9269,N_5206);
xnor U10807 (N_10807,N_7794,N_5784);
or U10808 (N_10808,N_7982,N_8379);
or U10809 (N_10809,N_7605,N_6876);
and U10810 (N_10810,N_7396,N_7202);
nand U10811 (N_10811,N_8877,N_6737);
nand U10812 (N_10812,N_8984,N_7996);
or U10813 (N_10813,N_7942,N_6311);
nand U10814 (N_10814,N_5019,N_8586);
and U10815 (N_10815,N_9337,N_5612);
and U10816 (N_10816,N_8123,N_6482);
xnor U10817 (N_10817,N_8389,N_7759);
or U10818 (N_10818,N_9699,N_5112);
nand U10819 (N_10819,N_5195,N_5969);
xor U10820 (N_10820,N_6707,N_8289);
and U10821 (N_10821,N_8996,N_6576);
or U10822 (N_10822,N_5305,N_9670);
xor U10823 (N_10823,N_7177,N_8549);
nand U10824 (N_10824,N_9340,N_6267);
or U10825 (N_10825,N_6362,N_8413);
and U10826 (N_10826,N_6317,N_6758);
xnor U10827 (N_10827,N_8672,N_9035);
or U10828 (N_10828,N_6155,N_6666);
and U10829 (N_10829,N_8342,N_7075);
xnor U10830 (N_10830,N_5505,N_8687);
nor U10831 (N_10831,N_9091,N_9867);
and U10832 (N_10832,N_8930,N_5723);
or U10833 (N_10833,N_5500,N_8784);
nand U10834 (N_10834,N_7741,N_8857);
and U10835 (N_10835,N_7668,N_8945);
nand U10836 (N_10836,N_7519,N_5625);
nand U10837 (N_10837,N_8776,N_8581);
and U10838 (N_10838,N_6598,N_5350);
nand U10839 (N_10839,N_8544,N_9656);
nor U10840 (N_10840,N_8746,N_9939);
and U10841 (N_10841,N_9228,N_6257);
nand U10842 (N_10842,N_8366,N_7239);
nor U10843 (N_10843,N_7005,N_8091);
or U10844 (N_10844,N_5101,N_6283);
nand U10845 (N_10845,N_5961,N_7574);
or U10846 (N_10846,N_7913,N_5692);
and U10847 (N_10847,N_8404,N_7158);
xnor U10848 (N_10848,N_7682,N_9608);
xor U10849 (N_10849,N_7457,N_7264);
nand U10850 (N_10850,N_5114,N_6968);
nor U10851 (N_10851,N_6776,N_7990);
xnor U10852 (N_10852,N_9386,N_7080);
and U10853 (N_10853,N_5666,N_6126);
and U10854 (N_10854,N_6014,N_7943);
nor U10855 (N_10855,N_8957,N_5273);
or U10856 (N_10856,N_6646,N_6878);
xor U10857 (N_10857,N_6484,N_9574);
xnor U10858 (N_10858,N_6377,N_5778);
nand U10859 (N_10859,N_7262,N_8978);
nand U10860 (N_10860,N_5927,N_5870);
nand U10861 (N_10861,N_6128,N_5861);
and U10862 (N_10862,N_7514,N_9619);
or U10863 (N_10863,N_8558,N_8684);
xor U10864 (N_10864,N_8084,N_5958);
nand U10865 (N_10865,N_8227,N_7693);
or U10866 (N_10866,N_9880,N_7083);
and U10867 (N_10867,N_9025,N_9397);
or U10868 (N_10868,N_6042,N_6938);
nor U10869 (N_10869,N_6113,N_8879);
nand U10870 (N_10870,N_5800,N_5608);
or U10871 (N_10871,N_6663,N_5491);
nand U10872 (N_10872,N_7054,N_6525);
nand U10873 (N_10873,N_6923,N_5731);
or U10874 (N_10874,N_8221,N_8584);
xor U10875 (N_10875,N_9627,N_5945);
nand U10876 (N_10876,N_9557,N_7517);
nor U10877 (N_10877,N_6147,N_5574);
nand U10878 (N_10878,N_8361,N_8386);
nor U10879 (N_10879,N_8073,N_9031);
nand U10880 (N_10880,N_7877,N_6382);
nand U10881 (N_10881,N_5551,N_5981);
nor U10882 (N_10882,N_6013,N_5734);
nor U10883 (N_10883,N_6294,N_7945);
nor U10884 (N_10884,N_9983,N_8369);
xor U10885 (N_10885,N_7802,N_9850);
and U10886 (N_10886,N_9141,N_6643);
or U10887 (N_10887,N_8732,N_5322);
nand U10888 (N_10888,N_5645,N_8461);
xor U10889 (N_10889,N_5498,N_9527);
nand U10890 (N_10890,N_5447,N_6687);
nand U10891 (N_10891,N_9232,N_9463);
or U10892 (N_10892,N_6940,N_8533);
xor U10893 (N_10893,N_9292,N_5843);
and U10894 (N_10894,N_5951,N_7268);
nor U10895 (N_10895,N_6917,N_7620);
nand U10896 (N_10896,N_7582,N_5655);
or U10897 (N_10897,N_6891,N_7840);
or U10898 (N_10898,N_8818,N_8225);
nor U10899 (N_10899,N_7744,N_5187);
or U10900 (N_10900,N_9310,N_6704);
or U10901 (N_10901,N_9128,N_7473);
nand U10902 (N_10902,N_5442,N_6832);
or U10903 (N_10903,N_9702,N_7368);
or U10904 (N_10904,N_6935,N_6880);
or U10905 (N_10905,N_9496,N_8286);
nand U10906 (N_10906,N_5396,N_6589);
nor U10907 (N_10907,N_5561,N_8055);
xnor U10908 (N_10908,N_7118,N_5379);
or U10909 (N_10909,N_9740,N_9647);
nor U10910 (N_10910,N_9588,N_6819);
nor U10911 (N_10911,N_6398,N_9856);
and U10912 (N_10912,N_7858,N_8085);
or U10913 (N_10913,N_9429,N_9357);
xor U10914 (N_10914,N_8045,N_5668);
xor U10915 (N_10915,N_8437,N_9022);
or U10916 (N_10916,N_5737,N_5119);
xnor U10917 (N_10917,N_8395,N_7972);
or U10918 (N_10918,N_8473,N_5494);
nor U10919 (N_10919,N_8806,N_9174);
xnor U10920 (N_10920,N_9881,N_6417);
and U10921 (N_10921,N_6238,N_8169);
nand U10922 (N_10922,N_9507,N_5433);
nor U10923 (N_10923,N_8332,N_6280);
or U10924 (N_10924,N_7007,N_6569);
nand U10925 (N_10925,N_8568,N_7257);
xor U10926 (N_10926,N_9673,N_5703);
and U10927 (N_10927,N_6838,N_7074);
xnor U10928 (N_10928,N_8569,N_7541);
and U10929 (N_10929,N_7204,N_9119);
or U10930 (N_10930,N_5029,N_6075);
nor U10931 (N_10931,N_7430,N_7917);
and U10932 (N_10932,N_8507,N_6875);
xnor U10933 (N_10933,N_5267,N_7540);
xor U10934 (N_10934,N_5418,N_5883);
nand U10935 (N_10935,N_6526,N_9927);
and U10936 (N_10936,N_7732,N_7604);
and U10937 (N_10937,N_6074,N_6617);
or U10938 (N_10938,N_6081,N_9279);
xnor U10939 (N_10939,N_6303,N_5567);
nor U10940 (N_10940,N_9814,N_9276);
or U10941 (N_10941,N_5271,N_6495);
xor U10942 (N_10942,N_8443,N_8048);
and U10943 (N_10943,N_8758,N_5429);
nor U10944 (N_10944,N_5792,N_9263);
or U10945 (N_10945,N_7030,N_8434);
and U10946 (N_10946,N_8493,N_6170);
and U10947 (N_10947,N_6259,N_5423);
nand U10948 (N_10948,N_5807,N_7484);
xor U10949 (N_10949,N_5834,N_8949);
nor U10950 (N_10950,N_6406,N_7226);
nand U10951 (N_10951,N_9979,N_7968);
xor U10952 (N_10952,N_5879,N_7706);
xor U10953 (N_10953,N_8354,N_7720);
nor U10954 (N_10954,N_8362,N_6800);
or U10955 (N_10955,N_5290,N_6316);
and U10956 (N_10956,N_7203,N_9060);
nand U10957 (N_10957,N_6638,N_5067);
nand U10958 (N_10958,N_6488,N_6473);
nor U10959 (N_10959,N_6586,N_6055);
and U10960 (N_10960,N_7038,N_7116);
and U10961 (N_10961,N_5401,N_5652);
nand U10962 (N_10962,N_9248,N_8309);
nor U10963 (N_10963,N_8051,N_9378);
nand U10964 (N_10964,N_8865,N_6017);
or U10965 (N_10965,N_8914,N_5131);
nand U10966 (N_10966,N_7872,N_8410);
or U10967 (N_10967,N_8464,N_8239);
and U10968 (N_10968,N_9440,N_5572);
and U10969 (N_10969,N_5191,N_6682);
and U10970 (N_10970,N_9426,N_6771);
xor U10971 (N_10971,N_9257,N_7495);
and U10972 (N_10972,N_7433,N_8545);
nor U10973 (N_10973,N_8822,N_6624);
or U10974 (N_10974,N_7797,N_5445);
xor U10975 (N_10975,N_6856,N_8367);
or U10976 (N_10976,N_9130,N_8106);
nand U10977 (N_10977,N_8278,N_8162);
and U10978 (N_10978,N_5716,N_7753);
nand U10979 (N_10979,N_8487,N_5603);
xnor U10980 (N_10980,N_6545,N_9450);
and U10981 (N_10981,N_5930,N_5123);
xor U10982 (N_10982,N_6916,N_6409);
xnor U10983 (N_10983,N_9600,N_7881);
nor U10984 (N_10984,N_8836,N_9350);
and U10985 (N_10985,N_8764,N_5390);
nand U10986 (N_10986,N_8151,N_7081);
nand U10987 (N_10987,N_6234,N_7067);
or U10988 (N_10988,N_8817,N_6498);
nor U10989 (N_10989,N_8236,N_7690);
nand U10990 (N_10990,N_6194,N_5616);
and U10991 (N_10991,N_5513,N_7062);
and U10992 (N_10992,N_8742,N_8734);
nand U10993 (N_10993,N_7516,N_6740);
nor U10994 (N_10994,N_5530,N_8429);
and U10995 (N_10995,N_6534,N_9886);
nor U10996 (N_10996,N_7796,N_6820);
and U10997 (N_10997,N_8328,N_6879);
and U10998 (N_10998,N_7362,N_7704);
and U10999 (N_10999,N_9246,N_5575);
or U11000 (N_11000,N_6817,N_9991);
and U11001 (N_11001,N_6487,N_7467);
nor U11002 (N_11002,N_8002,N_7560);
nor U11003 (N_11003,N_9851,N_8807);
and U11004 (N_11004,N_8457,N_5403);
xnor U11005 (N_11005,N_5528,N_8599);
or U11006 (N_11006,N_6027,N_5918);
xor U11007 (N_11007,N_9477,N_6112);
and U11008 (N_11008,N_6281,N_6805);
xor U11009 (N_11009,N_6195,N_5255);
nand U11010 (N_11010,N_6448,N_7375);
xor U11011 (N_11011,N_5903,N_6418);
or U11012 (N_11012,N_6700,N_9771);
or U11013 (N_11013,N_8186,N_5581);
and U11014 (N_11014,N_8480,N_5424);
or U11015 (N_11015,N_9315,N_9467);
xor U11016 (N_11016,N_6098,N_7160);
nor U11017 (N_11017,N_8485,N_8967);
nor U11018 (N_11018,N_8406,N_5643);
and U11019 (N_11019,N_8769,N_8990);
or U11020 (N_11020,N_5812,N_7579);
xor U11021 (N_11021,N_7799,N_5623);
xnor U11022 (N_11022,N_9683,N_9207);
xor U11023 (N_11023,N_5382,N_6208);
nor U11024 (N_11024,N_8079,N_9394);
nor U11025 (N_11025,N_8713,N_7566);
nor U11026 (N_11026,N_5992,N_8217);
nand U11027 (N_11027,N_9834,N_9088);
and U11028 (N_11028,N_6531,N_7715);
and U11029 (N_11029,N_5621,N_6571);
nand U11030 (N_11030,N_9410,N_5242);
or U11031 (N_11031,N_8299,N_5820);
nor U11032 (N_11032,N_9665,N_8736);
and U11033 (N_11033,N_7227,N_8833);
and U11034 (N_11034,N_5876,N_8292);
xnor U11035 (N_11035,N_9497,N_9830);
or U11036 (N_11036,N_9210,N_6982);
or U11037 (N_11037,N_5258,N_5516);
and U11038 (N_11038,N_9657,N_9173);
xnor U11039 (N_11039,N_6358,N_7317);
nor U11040 (N_11040,N_5470,N_8613);
and U11041 (N_11041,N_9167,N_7695);
and U11042 (N_11042,N_9705,N_5411);
xnor U11043 (N_11043,N_7225,N_9653);
nor U11044 (N_11044,N_9220,N_7740);
nand U11045 (N_11045,N_5960,N_9005);
or U11046 (N_11046,N_6915,N_9074);
and U11047 (N_11047,N_7860,N_5953);
xor U11048 (N_11048,N_6258,N_9651);
or U11049 (N_11049,N_5966,N_7590);
and U11050 (N_11050,N_6924,N_5803);
xnor U11051 (N_11051,N_6449,N_5074);
nand U11052 (N_11052,N_5662,N_9940);
and U11053 (N_11053,N_9824,N_6928);
or U11054 (N_11054,N_5804,N_7426);
or U11055 (N_11055,N_9142,N_6706);
nand U11056 (N_11056,N_6698,N_7013);
nand U11057 (N_11057,N_6168,N_9883);
or U11058 (N_11058,N_9379,N_5635);
nand U11059 (N_11059,N_9671,N_6339);
and U11060 (N_11060,N_7153,N_7245);
nand U11061 (N_11061,N_6840,N_9117);
nand U11062 (N_11062,N_9109,N_9785);
or U11063 (N_11063,N_9548,N_6607);
and U11064 (N_11064,N_6189,N_5022);
nor U11065 (N_11065,N_5150,N_8887);
nor U11066 (N_11066,N_7064,N_5378);
and U11067 (N_11067,N_5865,N_5108);
nand U11068 (N_11068,N_5855,N_5188);
and U11069 (N_11069,N_5795,N_5991);
nand U11070 (N_11070,N_9693,N_9398);
xor U11071 (N_11071,N_7258,N_7259);
or U11072 (N_11072,N_5560,N_7506);
and U11073 (N_11073,N_5057,N_8134);
and U11074 (N_11074,N_9599,N_8150);
nand U11075 (N_11075,N_5763,N_6855);
and U11076 (N_11076,N_7754,N_5027);
xnor U11077 (N_11077,N_7453,N_9363);
or U11078 (N_11078,N_7807,N_6123);
nand U11079 (N_11079,N_8617,N_6913);
nand U11080 (N_11080,N_6933,N_6665);
and U11081 (N_11081,N_9481,N_7589);
nor U11082 (N_11082,N_5838,N_5232);
and U11083 (N_11083,N_6340,N_6505);
xor U11084 (N_11084,N_7597,N_7551);
nand U11085 (N_11085,N_6514,N_8745);
xor U11086 (N_11086,N_7189,N_9589);
nand U11087 (N_11087,N_8725,N_9224);
or U11088 (N_11088,N_5660,N_6823);
nand U11089 (N_11089,N_8973,N_7887);
or U11090 (N_11090,N_9534,N_8728);
and U11091 (N_11091,N_9341,N_7113);
or U11092 (N_11092,N_9300,N_9675);
and U11093 (N_11093,N_6746,N_5007);
nor U11094 (N_11094,N_5488,N_5989);
nor U11095 (N_11095,N_7830,N_6847);
and U11096 (N_11096,N_6559,N_7878);
nand U11097 (N_11097,N_9614,N_8194);
xor U11098 (N_11098,N_5988,N_6097);
nand U11099 (N_11099,N_9360,N_9585);
nand U11100 (N_11100,N_5942,N_6724);
and U11101 (N_11101,N_9399,N_6783);
nand U11102 (N_11102,N_5363,N_7133);
nand U11103 (N_11103,N_8688,N_9470);
and U11104 (N_11104,N_7816,N_8040);
xnor U11105 (N_11105,N_8232,N_7978);
or U11106 (N_11106,N_6751,N_5041);
nor U11107 (N_11107,N_8543,N_5831);
xnor U11108 (N_11108,N_6520,N_9105);
nor U11109 (N_11109,N_7122,N_6312);
or U11110 (N_11110,N_5681,N_7959);
or U11111 (N_11111,N_9994,N_7546);
nand U11112 (N_11112,N_5324,N_8508);
xnor U11113 (N_11113,N_6386,N_5811);
or U11114 (N_11114,N_6529,N_6954);
nor U11115 (N_11115,N_9333,N_7825);
nor U11116 (N_11116,N_7014,N_5987);
and U11117 (N_11117,N_5667,N_5073);
or U11118 (N_11118,N_5854,N_6834);
nand U11119 (N_11119,N_5295,N_6093);
and U11120 (N_11120,N_9697,N_7127);
nor U11121 (N_11121,N_7059,N_6018);
and U11122 (N_11122,N_6732,N_5348);
nand U11123 (N_11123,N_6610,N_9054);
nand U11124 (N_11124,N_9779,N_6341);
or U11125 (N_11125,N_6109,N_9509);
nor U11126 (N_11126,N_8385,N_7215);
nand U11127 (N_11127,N_8615,N_5198);
and U11128 (N_11128,N_6801,N_5196);
xnor U11129 (N_11129,N_8840,N_7775);
nand U11130 (N_11130,N_5050,N_7520);
and U11131 (N_11131,N_8475,N_7011);
nor U11132 (N_11132,N_8255,N_5205);
xor U11133 (N_11133,N_9303,N_8439);
nor U11134 (N_11134,N_9828,N_6146);
or U11135 (N_11135,N_8053,N_6344);
and U11136 (N_11136,N_8107,N_7302);
or U11137 (N_11137,N_8119,N_7461);
or U11138 (N_11138,N_7111,N_6483);
nor U11139 (N_11139,N_7955,N_6611);
nor U11140 (N_11140,N_9129,N_6273);
or U11141 (N_11141,N_7844,N_6566);
xor U11142 (N_11142,N_9845,N_8440);
xor U11143 (N_11143,N_5499,N_8039);
nor U11144 (N_11144,N_6503,N_6591);
xnor U11145 (N_11145,N_8597,N_6959);
and U11146 (N_11146,N_7515,N_5519);
nor U11147 (N_11147,N_8965,N_7142);
or U11148 (N_11148,N_6965,N_9311);
or U11149 (N_11149,N_7859,N_7499);
or U11150 (N_11150,N_6248,N_7552);
nand U11151 (N_11151,N_5118,N_8570);
nand U11152 (N_11152,N_6507,N_6641);
or U11153 (N_11153,N_6254,N_6247);
xor U11154 (N_11154,N_5257,N_8054);
and U11155 (N_11155,N_9603,N_7383);
nand U11156 (N_11156,N_9387,N_6333);
nor U11157 (N_11157,N_6748,N_6811);
nor U11158 (N_11158,N_9446,N_7155);
xor U11159 (N_11159,N_5230,N_7905);
and U11160 (N_11160,N_6243,N_9716);
or U11161 (N_11161,N_5239,N_6735);
nor U11162 (N_11162,N_9176,N_6159);
or U11163 (N_11163,N_8340,N_9660);
nor U11164 (N_11164,N_6291,N_9321);
nor U11165 (N_11165,N_5699,N_8345);
xnor U11166 (N_11166,N_7052,N_8198);
or U11167 (N_11167,N_7182,N_9645);
xor U11168 (N_11168,N_9569,N_6588);
nor U11169 (N_11169,N_6186,N_6446);
and U11170 (N_11170,N_9891,N_5686);
or U11171 (N_11171,N_5862,N_8808);
nand U11172 (N_11172,N_6903,N_6768);
nand U11173 (N_11173,N_6071,N_8313);
or U11174 (N_11174,N_7656,N_5994);
xnor U11175 (N_11175,N_7482,N_8946);
and U11176 (N_11176,N_9454,N_6101);
nor U11177 (N_11177,N_6467,N_9612);
nor U11178 (N_11178,N_9539,N_6060);
or U11179 (N_11179,N_6660,N_7141);
and U11180 (N_11180,N_6955,N_8566);
nand U11181 (N_11181,N_9305,N_5558);
nor U11182 (N_11182,N_8970,N_9638);
and U11183 (N_11183,N_9144,N_7803);
nand U11184 (N_11184,N_7456,N_6064);
nor U11185 (N_11185,N_5436,N_6310);
nand U11186 (N_11186,N_8834,N_8172);
xor U11187 (N_11187,N_5982,N_5211);
nor U11188 (N_11188,N_7389,N_8838);
and U11189 (N_11189,N_7750,N_5189);
or U11190 (N_11190,N_5912,N_9741);
xnor U11191 (N_11191,N_5613,N_5589);
or U11192 (N_11192,N_8679,N_9489);
and U11193 (N_11193,N_8883,N_5144);
and U11194 (N_11194,N_8651,N_7861);
nand U11195 (N_11195,N_9899,N_7490);
xnor U11196 (N_11196,N_9369,N_9268);
nor U11197 (N_11197,N_7354,N_6249);
or U11198 (N_11198,N_7843,N_8110);
nand U11199 (N_11199,N_8588,N_6359);
or U11200 (N_11200,N_5314,N_5356);
and U11201 (N_11201,N_7557,N_9058);
and U11202 (N_11202,N_9358,N_6203);
nand U11203 (N_11203,N_8427,N_9937);
nor U11204 (N_11204,N_9620,N_8956);
and U11205 (N_11205,N_8639,N_5548);
and U11206 (N_11206,N_8392,N_9718);
or U11207 (N_11207,N_9667,N_9464);
or U11208 (N_11208,N_8633,N_9872);
and U11209 (N_11209,N_7132,N_8567);
or U11210 (N_11210,N_6211,N_6255);
or U11211 (N_11211,N_7289,N_8974);
nor U11212 (N_11212,N_9835,N_8585);
nand U11213 (N_11213,N_9763,N_9950);
xnor U11214 (N_11214,N_5678,N_6600);
nand U11215 (N_11215,N_7651,N_7373);
nand U11216 (N_11216,N_9000,N_5002);
nand U11217 (N_11217,N_8148,N_5414);
xor U11218 (N_11218,N_7394,N_7654);
xnor U11219 (N_11219,N_9213,N_6530);
and U11220 (N_11220,N_5848,N_7581);
or U11221 (N_11221,N_7855,N_9652);
nand U11222 (N_11222,N_8767,N_9604);
nor U11223 (N_11223,N_9461,N_5544);
or U11224 (N_11224,N_6718,N_9655);
xor U11225 (N_11225,N_7827,N_9662);
xnor U11226 (N_11226,N_5113,N_6814);
nand U11227 (N_11227,N_5405,N_7347);
nor U11228 (N_11228,N_5095,N_9707);
nor U11229 (N_11229,N_9952,N_7117);
and U11230 (N_11230,N_5157,N_8215);
and U11231 (N_11231,N_6200,N_5719);
xor U11232 (N_11232,N_5582,N_8303);
and U11233 (N_11233,N_7973,N_8905);
nand U11234 (N_11234,N_7988,N_9415);
or U11235 (N_11235,N_7382,N_5948);
and U11236 (N_11236,N_8190,N_6212);
and U11237 (N_11237,N_7761,N_6685);
nor U11238 (N_11238,N_9225,N_9298);
and U11239 (N_11239,N_7907,N_6554);
or U11240 (N_11240,N_9564,N_6767);
xor U11241 (N_11241,N_8988,N_7243);
and U11242 (N_11242,N_9859,N_8802);
xor U11243 (N_11243,N_7137,N_9199);
and U11244 (N_11244,N_8875,N_7247);
and U11245 (N_11245,N_9934,N_9925);
or U11246 (N_11246,N_5399,N_5543);
xnor U11247 (N_11247,N_9316,N_9854);
xnor U11248 (N_11248,N_8402,N_9678);
and U11249 (N_11249,N_7805,N_9116);
xnor U11250 (N_11250,N_7977,N_5693);
nor U11251 (N_11251,N_6816,N_7532);
and U11252 (N_11252,N_7086,N_7366);
and U11253 (N_11253,N_7617,N_5650);
xor U11254 (N_11254,N_8007,N_6474);
and U11255 (N_11255,N_7333,N_8903);
and U11256 (N_11256,N_8831,N_8189);
and U11257 (N_11257,N_6141,N_6353);
xnor U11258 (N_11258,N_6623,N_5909);
nor U11259 (N_11259,N_8191,N_9147);
and U11260 (N_11260,N_7345,N_7818);
nor U11261 (N_11261,N_7297,N_5711);
nor U11262 (N_11262,N_7922,N_6253);
and U11263 (N_11263,N_7738,N_9458);
xor U11264 (N_11264,N_9381,N_6535);
nand U11265 (N_11265,N_8173,N_6681);
xor U11266 (N_11266,N_6183,N_7938);
nor U11267 (N_11267,N_6137,N_7242);
xnor U11268 (N_11268,N_6991,N_8666);
xnor U11269 (N_11269,N_5160,N_7698);
or U11270 (N_11270,N_9874,N_8071);
nand U11271 (N_11271,N_6227,N_6778);
and U11272 (N_11272,N_6265,N_9535);
nor U11273 (N_11273,N_6635,N_7099);
or U11274 (N_11274,N_5099,N_9165);
nand U11275 (N_11275,N_5787,N_6908);
xnor U11276 (N_11276,N_9323,N_9244);
xnor U11277 (N_11277,N_5422,N_9586);
nand U11278 (N_11278,N_7965,N_5754);
nor U11279 (N_11279,N_9884,N_5768);
and U11280 (N_11280,N_7320,N_9594);
nand U11281 (N_11281,N_5278,N_5511);
nor U11282 (N_11282,N_7213,N_9965);
nor U11283 (N_11283,N_8416,N_5219);
xor U11284 (N_11284,N_6372,N_5675);
or U11285 (N_11285,N_7192,N_7392);
and U11286 (N_11286,N_5199,N_6714);
and U11287 (N_11287,N_6947,N_6656);
and U11288 (N_11288,N_5571,N_9307);
nor U11289 (N_11289,N_7765,N_5799);
nand U11290 (N_11290,N_7685,N_8316);
or U11291 (N_11291,N_9449,N_6612);
nor U11292 (N_11292,N_5615,N_8383);
nor U11293 (N_11293,N_8804,N_6738);
nand U11294 (N_11294,N_9728,N_7600);
nand U11295 (N_11295,N_7044,N_7804);
xnor U11296 (N_11296,N_8336,N_8296);
nand U11297 (N_11297,N_7386,N_5996);
and U11298 (N_11298,N_5597,N_9909);
or U11299 (N_11299,N_6011,N_9044);
and U11300 (N_11300,N_9293,N_6039);
xor U11301 (N_11301,N_9864,N_9107);
and U11302 (N_11302,N_6078,N_7504);
xor U11303 (N_11303,N_6485,N_7789);
nand U11304 (N_11304,N_7568,N_5223);
and U11305 (N_11305,N_7632,N_5486);
nand U11306 (N_11306,N_7498,N_9445);
nand U11307 (N_11307,N_9070,N_6762);
or U11308 (N_11308,N_7355,N_9529);
xor U11309 (N_11309,N_5135,N_7569);
and U11310 (N_11310,N_7361,N_6769);
xor U11311 (N_11311,N_6630,N_6106);
xor U11312 (N_11312,N_5476,N_9229);
or U11313 (N_11313,N_6994,N_7115);
nor U11314 (N_11314,N_5857,N_6906);
xor U11315 (N_11315,N_6900,N_6095);
or U11316 (N_11316,N_7997,N_6573);
nand U11317 (N_11317,N_9036,N_9407);
or U11318 (N_11318,N_9963,N_9816);
nor U11319 (N_11319,N_6348,N_5292);
xnor U11320 (N_11320,N_8711,N_9951);
nand U11321 (N_11321,N_7762,N_9918);
nand U11322 (N_11322,N_9384,N_7689);
nor U11323 (N_11323,N_5362,N_5789);
nand U11324 (N_11324,N_9320,N_6400);
xnor U11325 (N_11325,N_9843,N_5733);
nand U11326 (N_11326,N_5005,N_5638);
and U11327 (N_11327,N_5238,N_8564);
nand U11328 (N_11328,N_6167,N_8995);
or U11329 (N_11329,N_5837,N_7311);
nor U11330 (N_11330,N_7708,N_7032);
or U11331 (N_11331,N_7660,N_5432);
nand U11332 (N_11332,N_8733,N_5863);
and U11333 (N_11333,N_7187,N_6401);
xor U11334 (N_11334,N_6864,N_8337);
and U11335 (N_11335,N_6411,N_8727);
and U11336 (N_11336,N_7181,N_6138);
nor U11337 (N_11337,N_9920,N_5670);
xor U11338 (N_11338,N_6347,N_5646);
nand U11339 (N_11339,N_8787,N_6725);
nor U11340 (N_11340,N_7091,N_5370);
nor U11341 (N_11341,N_5893,N_8636);
and U11342 (N_11342,N_8431,N_5079);
xnor U11343 (N_11343,N_8057,N_6477);
nand U11344 (N_11344,N_7771,N_8977);
and U11345 (N_11345,N_9996,N_9411);
and U11346 (N_11346,N_8203,N_7034);
nand U11347 (N_11347,N_6942,N_8829);
and U11348 (N_11348,N_5354,N_7162);
xor U11349 (N_11349,N_7637,N_8872);
and U11350 (N_11350,N_9134,N_6517);
or U11351 (N_11351,N_6445,N_9768);
and U11352 (N_11352,N_5497,N_8563);
nor U11353 (N_11353,N_5880,N_5782);
nor U11354 (N_11354,N_6193,N_5774);
nand U11355 (N_11355,N_9704,N_7003);
nor U11356 (N_11356,N_5478,N_6373);
and U11357 (N_11357,N_7793,N_9402);
nand U11358 (N_11358,N_5220,N_9286);
nand U11359 (N_11359,N_6848,N_7586);
nor U11360 (N_11360,N_6777,N_8648);
or U11361 (N_11361,N_8591,N_8305);
and U11362 (N_11362,N_6743,N_7851);
or U11363 (N_11363,N_7195,N_7967);
or U11364 (N_11364,N_7954,N_8775);
nand U11365 (N_11365,N_5922,N_7911);
and U11366 (N_11366,N_7533,N_7246);
xor U11367 (N_11367,N_7402,N_5701);
nand U11368 (N_11368,N_7562,N_9551);
xor U11369 (N_11369,N_5797,N_6454);
xor U11370 (N_11370,N_8925,N_5842);
nand U11371 (N_11371,N_9444,N_9013);
nand U11372 (N_11372,N_7677,N_7244);
or U11373 (N_11373,N_9367,N_8828);
and U11374 (N_11374,N_7255,N_5208);
xnor U11375 (N_11375,N_6413,N_9375);
nor U11376 (N_11376,N_8323,N_8438);
or U11377 (N_11377,N_6547,N_5082);
or U11378 (N_11378,N_9720,N_7649);
or U11379 (N_11379,N_7831,N_8709);
nor U11380 (N_11380,N_5138,N_7846);
xor U11381 (N_11381,N_5755,N_5033);
or U11382 (N_11382,N_6105,N_6010);
nor U11383 (N_11383,N_8442,N_8240);
nor U11384 (N_11384,N_5740,N_8640);
nand U11385 (N_11385,N_9643,N_5827);
xnor U11386 (N_11386,N_6798,N_9692);
nor U11387 (N_11387,N_6416,N_6197);
or U11388 (N_11388,N_5308,N_7327);
nand U11389 (N_11389,N_8200,N_5940);
or U11390 (N_11390,N_7575,N_9694);
nand U11391 (N_11391,N_9368,N_5691);
nor U11392 (N_11392,N_9736,N_6292);
nor U11393 (N_11393,N_5376,N_6671);
nor U11394 (N_11394,N_7053,N_9079);
and U11395 (N_11395,N_8906,N_5832);
or U11396 (N_11396,N_5507,N_7815);
nand U11397 (N_11397,N_6419,N_5176);
xor U11398 (N_11398,N_8213,N_8660);
nand U11399 (N_11399,N_8608,N_5702);
xor U11400 (N_11400,N_8625,N_7676);
nand U11401 (N_11401,N_7638,N_8016);
nor U11402 (N_11402,N_9296,N_7198);
and U11403 (N_11403,N_8037,N_7436);
nand U11404 (N_11404,N_6001,N_6172);
or U11405 (N_11405,N_6100,N_5512);
and U11406 (N_11406,N_8495,N_7931);
and U11407 (N_11407,N_7143,N_8607);
or U11408 (N_11408,N_9729,N_8740);
xor U11409 (N_11409,N_5708,N_6548);
or U11410 (N_11410,N_9145,N_6871);
or U11411 (N_11411,N_9869,N_7463);
nor U11412 (N_11412,N_5746,N_8409);
and U11413 (N_11413,N_6217,N_6792);
or U11414 (N_11414,N_5237,N_5689);
xor U11415 (N_11415,N_9418,N_9048);
or U11416 (N_11416,N_6026,N_8154);
and U11417 (N_11417,N_9390,N_6750);
nand U11418 (N_11418,N_9327,N_6002);
nor U11419 (N_11419,N_5510,N_8441);
xnor U11420 (N_11420,N_7745,N_7040);
nand U11421 (N_11421,N_5256,N_6515);
xor U11422 (N_11422,N_7348,N_5043);
nor U11423 (N_11423,N_6593,N_9063);
xnor U11424 (N_11424,N_5735,N_8265);
nand U11425 (N_11425,N_5685,N_8061);
nor U11426 (N_11426,N_9636,N_9506);
and U11427 (N_11427,N_6432,N_6726);
and U11428 (N_11428,N_5936,N_8676);
nor U11429 (N_11429,N_9605,N_7646);
nand U11430 (N_11430,N_9640,N_9637);
xnor U11431 (N_11431,N_9760,N_5627);
nand U11432 (N_11432,N_8370,N_5584);
or U11433 (N_11433,N_9674,N_9171);
and U11434 (N_11434,N_6327,N_6290);
or U11435 (N_11435,N_8702,N_7397);
nor U11436 (N_11436,N_7606,N_9339);
or U11437 (N_11437,N_7643,N_9436);
nand U11438 (N_11438,N_6163,N_7035);
and U11439 (N_11439,N_7464,N_9417);
nand U11440 (N_11440,N_6499,N_9826);
xnor U11441 (N_11441,N_5791,N_6755);
or U11442 (N_11442,N_8665,N_9795);
and U11443 (N_11443,N_7966,N_7944);
and U11444 (N_11444,N_5279,N_7545);
nor U11445 (N_11445,N_7722,N_9331);
nor U11446 (N_11446,N_6070,N_5482);
or U11447 (N_11447,N_7834,N_6158);
nand U11448 (N_11448,N_6354,N_9329);
nor U11449 (N_11449,N_7653,N_6645);
nor U11450 (N_11450,N_7992,N_7110);
nand U11451 (N_11451,N_7730,N_5759);
xor U11452 (N_11452,N_5676,N_9284);
and U11453 (N_11453,N_6263,N_6541);
or U11454 (N_11454,N_5395,N_6309);
xor U11455 (N_11455,N_9515,N_7313);
nor U11456 (N_11456,N_9725,N_6277);
xor U11457 (N_11457,N_7824,N_5730);
or U11458 (N_11458,N_9231,N_5044);
nand U11459 (N_11459,N_9149,N_5441);
nor U11460 (N_11460,N_7440,N_6615);
nand U11461 (N_11461,N_7161,N_7897);
nor U11462 (N_11462,N_8378,N_7371);
nand U11463 (N_11463,N_9764,N_9009);
xnor U11464 (N_11464,N_6414,N_8478);
nor U11465 (N_11465,N_5900,N_9661);
nor U11466 (N_11466,N_6770,N_8614);
nor U11467 (N_11467,N_7681,N_6494);
and U11468 (N_11468,N_6949,N_6190);
xnor U11469 (N_11469,N_8546,N_9875);
or U11470 (N_11470,N_9017,N_7027);
nand U11471 (N_11471,N_8018,N_6246);
or U11472 (N_11472,N_8531,N_6385);
or U11473 (N_11473,N_6244,N_9156);
nor U11474 (N_11474,N_7508,N_8283);
nand U11475 (N_11475,N_8705,N_6932);
nand U11476 (N_11476,N_7179,N_7994);
xnor U11477 (N_11477,N_5444,N_9239);
and U11478 (N_11478,N_6119,N_7717);
xnor U11479 (N_11479,N_7979,N_7868);
or U11480 (N_11480,N_9453,N_5717);
and U11481 (N_11481,N_8125,N_6177);
xnor U11482 (N_11482,N_8263,N_9990);
and U11483 (N_11483,N_9359,N_8739);
and U11484 (N_11484,N_7705,N_9973);
nand U11485 (N_11485,N_9946,N_7763);
nor U11486 (N_11486,N_9753,N_9267);
xor U11487 (N_11487,N_5045,N_8628);
and U11488 (N_11488,N_9490,N_8943);
or U11489 (N_11489,N_8616,N_7358);
or U11490 (N_11490,N_5539,N_9530);
xor U11491 (N_11491,N_6730,N_8415);
nand U11492 (N_11492,N_9061,N_7956);
or U11493 (N_11493,N_5450,N_9615);
or U11494 (N_11494,N_8518,N_5400);
or U11495 (N_11495,N_5718,N_6580);
nor U11496 (N_11496,N_8046,N_8821);
or U11497 (N_11497,N_7071,N_8087);
nor U11498 (N_11498,N_8131,N_9078);
nand U11499 (N_11499,N_8143,N_5394);
nor U11500 (N_11500,N_7883,N_8815);
nand U11501 (N_11501,N_9587,N_7335);
nor U11502 (N_11502,N_7369,N_6444);
and U11503 (N_11503,N_9847,N_6127);
nand U11504 (N_11504,N_8513,N_5218);
nand U11505 (N_11505,N_9330,N_5725);
nor U11506 (N_11506,N_5762,N_5896);
or U11507 (N_11507,N_5120,N_5594);
xor U11508 (N_11508,N_7121,N_5806);
xor U11509 (N_11509,N_8049,N_6391);
and U11510 (N_11510,N_9151,N_6004);
or U11511 (N_11511,N_7962,N_9681);
nand U11512 (N_11512,N_5102,N_7618);
and U11513 (N_11513,N_9921,N_7407);
xnor U11514 (N_11514,N_9297,N_7971);
xor U11515 (N_11515,N_9046,N_5063);
xnor U11516 (N_11516,N_6476,N_9396);
nor U11517 (N_11517,N_5712,N_6029);
or U11518 (N_11518,N_8793,N_6502);
and U11519 (N_11519,N_9112,N_6210);
or U11520 (N_11520,N_6171,N_7950);
and U11521 (N_11521,N_9787,N_7553);
xor U11522 (N_11522,N_5777,N_7339);
xnor U11523 (N_11523,N_7380,N_9525);
nor U11524 (N_11524,N_9319,N_5347);
nor U11525 (N_11525,N_5263,N_5285);
xor U11526 (N_11526,N_6329,N_9923);
xor U11527 (N_11527,N_6664,N_5825);
and U11528 (N_11528,N_9371,N_7974);
xor U11529 (N_11529,N_6640,N_9669);
xnor U11530 (N_11530,N_9389,N_8669);
or U11531 (N_11531,N_8145,N_8650);
nor U11532 (N_11532,N_8445,N_6228);
nor U11533 (N_11533,N_5280,N_7898);
nor U11534 (N_11534,N_8626,N_9200);
or U11535 (N_11535,N_6642,N_9001);
and U11536 (N_11536,N_9014,N_8074);
and U11537 (N_11537,N_7625,N_5868);
nand U11538 (N_11538,N_6516,N_9755);
nor U11539 (N_11539,N_9807,N_6745);
and U11540 (N_11540,N_6486,N_5690);
and U11541 (N_11541,N_6511,N_8512);
nor U11542 (N_11542,N_9010,N_9981);
or U11543 (N_11543,N_8955,N_5451);
and U11544 (N_11544,N_6114,N_6285);
nand U11545 (N_11545,N_8115,N_9749);
and U11546 (N_11546,N_6658,N_5153);
and U11547 (N_11547,N_6059,N_8122);
nand U11548 (N_11548,N_8372,N_5964);
nand U11549 (N_11549,N_7438,N_5610);
or U11550 (N_11550,N_9547,N_7234);
and U11551 (N_11551,N_9143,N_8238);
xor U11552 (N_11552,N_5216,N_7076);
nor U11553 (N_11553,N_8744,N_9894);
xor U11554 (N_11554,N_5911,N_9273);
or U11555 (N_11555,N_8771,N_6509);
or U11556 (N_11556,N_9932,N_6715);
and U11557 (N_11557,N_9865,N_8839);
and U11558 (N_11558,N_7356,N_7577);
xnor U11559 (N_11559,N_6145,N_7101);
nor U11560 (N_11560,N_8219,N_8396);
and U11561 (N_11561,N_9892,N_8976);
nand U11562 (N_11562,N_6719,N_6472);
or U11563 (N_11563,N_6558,N_6542);
nor U11564 (N_11564,N_6068,N_5933);
or U11565 (N_11565,N_7393,N_8029);
nand U11566 (N_11566,N_6945,N_9343);
and U11567 (N_11567,N_7031,N_9275);
or U11568 (N_11568,N_6230,N_7891);
xor U11569 (N_11569,N_7536,N_6723);
nor U11570 (N_11570,N_7713,N_7360);
xor U11571 (N_11571,N_6918,N_6433);
nand U11572 (N_11572,N_8448,N_8579);
or U11573 (N_11573,N_6688,N_8885);
or U11574 (N_11574,N_8026,N_6851);
or U11575 (N_11575,N_9342,N_6496);
and U11576 (N_11576,N_9004,N_9049);
nand U11577 (N_11577,N_6970,N_9019);
nor U11578 (N_11578,N_5462,N_6233);
nor U11579 (N_11579,N_6201,N_9280);
and U11580 (N_11580,N_7070,N_8618);
and U11581 (N_11581,N_9819,N_8167);
nand U11582 (N_11582,N_8939,N_8424);
xor U11583 (N_11583,N_7528,N_5355);
nand U11584 (N_11584,N_9413,N_6429);
xor U11585 (N_11585,N_5228,N_7976);
xnor U11586 (N_11586,N_6981,N_5483);
and U11587 (N_11587,N_9099,N_8422);
nor U11588 (N_11588,N_7623,N_5538);
nand U11589 (N_11589,N_8795,N_8851);
nand U11590 (N_11590,N_5833,N_8908);
and U11591 (N_11591,N_5251,N_5898);
nor U11592 (N_11592,N_7671,N_6437);
xnor U11593 (N_11593,N_7901,N_8983);
nand U11594 (N_11594,N_7870,N_6415);
and U11595 (N_11595,N_9104,N_6972);
xnor U11596 (N_11596,N_8966,N_5805);
and U11597 (N_11597,N_7735,N_7613);
or U11598 (N_11598,N_7570,N_7882);
or U11599 (N_11599,N_9085,N_7854);
and U11600 (N_11600,N_7639,N_5622);
and U11601 (N_11601,N_6085,N_7626);
nand U11602 (N_11602,N_5039,N_7920);
nand U11603 (N_11603,N_6549,N_7885);
and U11604 (N_11604,N_7659,N_5753);
or U11605 (N_11605,N_7024,N_9498);
nand U11606 (N_11606,N_6422,N_7810);
xor U11607 (N_11607,N_7611,N_7867);
nand U11608 (N_11608,N_8646,N_7836);
or U11609 (N_11609,N_7564,N_8022);
nand U11610 (N_11610,N_7935,N_6652);
nand U11611 (N_11611,N_7197,N_6000);
or U11612 (N_11612,N_6180,N_6050);
nand U11613 (N_11613,N_5072,N_6570);
or U11614 (N_11614,N_8928,N_6897);
or U11615 (N_11615,N_5628,N_5100);
and U11616 (N_11616,N_5841,N_8069);
and U11617 (N_11617,N_8894,N_5456);
or U11618 (N_11618,N_5993,N_9829);
nand U11619 (N_11619,N_5317,N_6072);
xor U11620 (N_11620,N_5779,N_6651);
and U11621 (N_11621,N_6690,N_5990);
nand U11622 (N_11622,N_6632,N_5128);
and U11623 (N_11623,N_7298,N_8936);
and U11624 (N_11624,N_7702,N_5860);
and U11625 (N_11625,N_7450,N_9215);
and U11626 (N_11626,N_6829,N_8572);
nand U11627 (N_11627,N_9264,N_7543);
nor U11628 (N_11628,N_9742,N_5732);
xnor U11629 (N_11629,N_5302,N_8689);
nand U11630 (N_11630,N_6633,N_9034);
nand U11631 (N_11631,N_9309,N_5260);
xor U11632 (N_11632,N_5639,N_8576);
and U11633 (N_11633,N_9949,N_6694);
nor U11634 (N_11634,N_9849,N_7217);
and U11635 (N_11635,N_9385,N_5962);
nand U11636 (N_11636,N_8135,N_9799);
nand U11637 (N_11637,N_7173,N_5169);
nor U11638 (N_11638,N_7363,N_7902);
or U11639 (N_11639,N_5656,N_7699);
xor U11640 (N_11640,N_5813,N_9072);
xor U11641 (N_11641,N_9033,N_7731);
xnor U11642 (N_11642,N_5325,N_6873);
nor U11643 (N_11643,N_8811,N_5122);
xnor U11644 (N_11644,N_9676,N_6139);
xor U11645 (N_11645,N_5438,N_8229);
nand U11646 (N_11646,N_7657,N_8494);
nor U11647 (N_11647,N_7303,N_8577);
or U11648 (N_11648,N_9572,N_9205);
nor U11649 (N_11649,N_6438,N_7401);
xnor U11650 (N_11650,N_8846,N_8785);
or U11651 (N_11651,N_5493,N_6425);
nor U11652 (N_11652,N_5794,N_7010);
or U11653 (N_11653,N_7119,N_5086);
and U11654 (N_11654,N_5776,N_9761);
xnor U11655 (N_11655,N_5738,N_5965);
nor U11656 (N_11656,N_8421,N_7465);
nand U11657 (N_11657,N_6956,N_6019);
xnor U11658 (N_11658,N_9748,N_6885);
nor U11659 (N_11659,N_8466,N_9314);
or U11660 (N_11660,N_6274,N_8171);
nor U11661 (N_11661,N_5233,N_6306);
nand U11662 (N_11662,N_9216,N_9401);
xor U11663 (N_11663,N_9629,N_5901);
and U11664 (N_11664,N_5252,N_8858);
nand U11665 (N_11665,N_6890,N_6978);
or U11666 (N_11666,N_5649,N_7777);
nor U11667 (N_11667,N_8339,N_5984);
xor U11668 (N_11668,N_9511,N_9198);
nor U11669 (N_11669,N_7199,N_7599);
and U11670 (N_11670,N_9003,N_8920);
nand U11671 (N_11671,N_9439,N_7222);
xnor U11672 (N_11672,N_8152,N_5130);
nand U11673 (N_11673,N_6229,N_5749);
nor U11674 (N_11674,N_8506,N_8324);
or U11675 (N_11675,N_5798,N_6766);
nor U11676 (N_11676,N_7650,N_7208);
and U11677 (N_11677,N_8604,N_8489);
xor U11678 (N_11678,N_9953,N_8753);
or U11679 (N_11679,N_5016,N_7687);
nor U11680 (N_11680,N_8177,N_6782);
and U11681 (N_11681,N_6120,N_8295);
xnor U11682 (N_11682,N_9978,N_5672);
nand U11683 (N_11683,N_7415,N_8712);
or U11684 (N_11684,N_9443,N_7254);
or U11685 (N_11685,N_9738,N_6691);
nor U11686 (N_11686,N_5573,N_5332);
nor U11687 (N_11687,N_5374,N_6995);
and U11688 (N_11688,N_5105,N_7806);
xor U11689 (N_11689,N_9943,N_8454);
xnor U11690 (N_11690,N_9733,N_9152);
and U11691 (N_11691,N_8635,N_6537);
nor U11692 (N_11692,N_6501,N_6987);
and U11693 (N_11693,N_8538,N_9945);
nand U11694 (N_11694,N_8352,N_7093);
nor U11695 (N_11695,N_9392,N_5908);
and U11696 (N_11696,N_9563,N_8128);
and U11697 (N_11697,N_9688,N_7261);
xor U11698 (N_11698,N_7795,N_8714);
and U11699 (N_11699,N_8420,N_6215);
and U11700 (N_11700,N_9957,N_9561);
and U11701 (N_11701,N_7721,N_6099);
nand U11702 (N_11702,N_6102,N_8092);
and U11703 (N_11703,N_9190,N_6087);
and U11704 (N_11704,N_6984,N_7666);
nand U11705 (N_11705,N_8180,N_7391);
nor U11706 (N_11706,N_7478,N_7106);
nand U11707 (N_11707,N_6939,N_6390);
and U11708 (N_11708,N_7629,N_9434);
or U11709 (N_11709,N_7447,N_8654);
xnor U11710 (N_11710,N_8820,N_5334);
nor U11711 (N_11711,N_9579,N_6157);
nand U11712 (N_11712,N_7417,N_9501);
nand U11713 (N_11713,N_5009,N_7584);
xnor U11714 (N_11714,N_6859,N_8869);
nor U11715 (N_11715,N_5194,N_9625);
xnor U11716 (N_11716,N_7838,N_7952);
and U11717 (N_11717,N_8701,N_7149);
or U11718 (N_11718,N_8102,N_8918);
nand U11719 (N_11719,N_8942,N_5054);
xnor U11720 (N_11720,N_9037,N_6275);
and U11721 (N_11721,N_6497,N_8931);
and U11722 (N_11722,N_6424,N_6765);
nor U11723 (N_11723,N_5291,N_6063);
xnor U11724 (N_11724,N_7139,N_7485);
or U11725 (N_11725,N_7041,N_6466);
nand U11726 (N_11726,N_8954,N_5083);
nor U11727 (N_11727,N_6143,N_8755);
and U11728 (N_11728,N_9947,N_6404);
or U11729 (N_11729,N_5222,N_5983);
and U11730 (N_11730,N_7159,N_7826);
nand U11731 (N_11731,N_9595,N_9533);
nor U11732 (N_11732,N_8320,N_5058);
and U11733 (N_11733,N_6650,N_9719);
or U11734 (N_11734,N_5437,N_8637);
and U11735 (N_11735,N_6307,N_7998);
or U11736 (N_11736,N_5023,N_6693);
or U11737 (N_11737,N_6518,N_5907);
nand U11738 (N_11738,N_5361,N_9820);
xor U11739 (N_11739,N_7175,N_5830);
and U11740 (N_11740,N_8182,N_8912);
or U11741 (N_11741,N_6209,N_6625);
nor U11742 (N_11742,N_6447,N_9124);
xor U11743 (N_11743,N_7910,N_6140);
and U11744 (N_11744,N_8300,N_7066);
and U11745 (N_11745,N_5115,N_7856);
and U11746 (N_11746,N_5484,N_7980);
xnor U11747 (N_11747,N_9421,N_6649);
or U11748 (N_11748,N_7757,N_8837);
or U11749 (N_11749,N_6713,N_8269);
nand U11750 (N_11750,N_9575,N_6971);
and U11751 (N_11751,N_8768,N_8638);
nor U11752 (N_11752,N_8678,N_5406);
and U11753 (N_11753,N_7455,N_9092);
nor U11754 (N_11754,N_7494,N_5788);
nand U11755 (N_11755,N_5209,N_9650);
and U11756 (N_11756,N_8208,N_5881);
nor U11757 (N_11757,N_5261,N_6367);
or U11758 (N_11758,N_9448,N_9081);
xnor U11759 (N_11759,N_8502,N_7863);
or U11760 (N_11760,N_9469,N_9995);
nand U11761 (N_11761,N_7477,N_6973);
or U11762 (N_11762,N_8327,N_6692);
nor U11763 (N_11763,N_8683,N_7443);
xnor U11764 (N_11764,N_8964,N_6786);
nand U11765 (N_11765,N_8343,N_6551);
nor U11766 (N_11766,N_9971,N_7525);
nand U11767 (N_11767,N_8675,N_8929);
xnor U11768 (N_11768,N_7385,N_8951);
nand U11769 (N_11769,N_5106,N_9262);
or U11770 (N_11770,N_7591,N_6287);
or U11771 (N_11771,N_6952,N_5139);
xor U11772 (N_11772,N_9642,N_8867);
nand U11773 (N_11773,N_8212,N_8741);
and U11774 (N_11774,N_9472,N_9282);
nand U11775 (N_11775,N_6226,N_5137);
or U11776 (N_11776,N_7279,N_7459);
nor U11777 (N_11777,N_8430,N_7862);
and U11778 (N_11778,N_6440,N_7537);
nor U11779 (N_11779,N_8341,N_8562);
and U11780 (N_11780,N_9474,N_8752);
xnor U11781 (N_11781,N_9905,N_9007);
and U11782 (N_11782,N_5968,N_5479);
xor U11783 (N_11783,N_7934,N_6842);
xnor U11784 (N_11784,N_7712,N_6149);
nand U11785 (N_11785,N_9196,N_8658);
or U11786 (N_11786,N_5110,N_6231);
and U11787 (N_11787,N_6910,N_8790);
xnor U11788 (N_11788,N_6609,N_8220);
or U11789 (N_11789,N_7481,N_6627);
and U11790 (N_11790,N_7284,N_8860);
xnor U11791 (N_11791,N_9781,N_8013);
nand U11792 (N_11792,N_6960,N_8297);
nand U11793 (N_11793,N_8397,N_7497);
nor U11794 (N_11794,N_5346,N_5503);
xor U11795 (N_11795,N_8419,N_8334);
or U11796 (N_11796,N_8393,N_8491);
nand U11797 (N_11797,N_6023,N_6619);
nor U11798 (N_11798,N_8144,N_5087);
and U11799 (N_11799,N_5162,N_7305);
xnor U11800 (N_11800,N_7414,N_9065);
and U11801 (N_11801,N_8467,N_6469);
or U11802 (N_11802,N_8791,N_6107);
or U11803 (N_11803,N_5748,N_9218);
nand U11804 (N_11804,N_6936,N_7511);
nand U11805 (N_11805,N_9414,N_6852);
or U11806 (N_11806,N_5904,N_5605);
and U11807 (N_11807,N_6402,N_6268);
xor U11808 (N_11808,N_7518,N_8015);
and U11809 (N_11809,N_5977,N_7374);
nor U11810 (N_11810,N_8695,N_6108);
nand U11811 (N_11811,N_7176,N_8539);
xor U11812 (N_11812,N_9800,N_6524);
nand U11813 (N_11813,N_7148,N_9125);
and U11814 (N_11814,N_6185,N_9598);
or U11815 (N_11815,N_5495,N_6213);
nor U11816 (N_11816,N_7006,N_8377);
xnor U11817 (N_11817,N_8556,N_9067);
and U11818 (N_11818,N_5726,N_5244);
xor U11819 (N_11819,N_7530,N_8703);
xnor U11820 (N_11820,N_5443,N_8097);
xor U11821 (N_11821,N_5161,N_5897);
nand U11822 (N_11822,N_5038,N_9388);
xor U11823 (N_11823,N_5193,N_8716);
xor U11824 (N_11824,N_6657,N_5614);
or U11825 (N_11825,N_5146,N_9313);
xor U11826 (N_11826,N_5003,N_5772);
nor U11827 (N_11827,N_5583,N_7009);
or U11828 (N_11828,N_5047,N_8765);
and U11829 (N_11829,N_9073,N_9818);
or U11830 (N_11830,N_6557,N_5545);
or U11831 (N_11831,N_7442,N_9682);
or U11832 (N_11832,N_7112,N_9373);
xnor U11833 (N_11833,N_9641,N_6286);
and U11834 (N_11834,N_7315,N_9935);
and U11835 (N_11835,N_7088,N_7908);
and U11836 (N_11836,N_8310,N_5770);
or U11837 (N_11837,N_5270,N_6869);
nor U11838 (N_11838,N_8534,N_8794);
and U11839 (N_11839,N_6920,N_8706);
and U11840 (N_11840,N_8469,N_8835);
xor U11841 (N_11841,N_8472,N_9502);
or U11842 (N_11842,N_7102,N_8663);
and U11843 (N_11843,N_6717,N_5919);
or U11844 (N_11844,N_7323,N_9848);
and U11845 (N_11845,N_6028,N_9876);
and U11846 (N_11846,N_9277,N_8043);
or U11847 (N_11847,N_8285,N_8876);
nand U11848 (N_11848,N_5475,N_8847);
and U11849 (N_11849,N_7940,N_6647);
xor U11850 (N_11850,N_8010,N_5068);
and U11851 (N_11851,N_6269,N_8349);
nand U11852 (N_11852,N_7424,N_8241);
nor U11853 (N_11853,N_8523,N_5366);
and U11854 (N_11854,N_9717,N_8801);
nor U11855 (N_11855,N_5421,N_6629);
or U11856 (N_11856,N_9734,N_7674);
nand U11857 (N_11857,N_5051,N_9038);
nand U11858 (N_11858,N_6489,N_6412);
and U11859 (N_11859,N_6988,N_9416);
xor U11860 (N_11860,N_6458,N_8479);
nor U11861 (N_11861,N_9170,N_9403);
or U11862 (N_11862,N_6408,N_7343);
xor U11863 (N_11863,N_5892,N_8856);
nor U11864 (N_11864,N_7340,N_6815);
or U11865 (N_11865,N_9775,N_9582);
nor U11866 (N_11866,N_8248,N_5925);
xor U11867 (N_11867,N_8960,N_7201);
xor U11868 (N_11868,N_6492,N_9523);
or U11869 (N_11869,N_6893,N_6206);
xor U11870 (N_11870,N_9374,N_7561);
xnor U11871 (N_11871,N_7241,N_7642);
nand U11872 (N_11872,N_5098,N_8824);
nor U11873 (N_11873,N_7527,N_5075);
nand U11874 (N_11874,N_6667,N_8009);
nor U11875 (N_11875,N_8673,N_9484);
or U11876 (N_11876,N_5521,N_5526);
nor U11877 (N_11877,N_8864,N_8700);
xor U11878 (N_11878,N_6421,N_7601);
nor U11879 (N_11879,N_5177,N_5064);
xor U11880 (N_11880,N_5722,N_9633);
nor U11881 (N_11881,N_5179,N_9654);
or U11882 (N_11882,N_9353,N_6218);
and U11883 (N_11883,N_7523,N_9964);
nand U11884 (N_11884,N_9185,N_6927);
nor U11885 (N_11885,N_9020,N_7873);
and U11886 (N_11886,N_5611,N_8950);
and U11887 (N_11887,N_7847,N_6532);
or U11888 (N_11888,N_8112,N_8677);
nand U11889 (N_11889,N_9294,N_5469);
and U11890 (N_11890,N_8630,N_9108);
and U11891 (N_11891,N_9844,N_5288);
and U11892 (N_11892,N_7483,N_7212);
nand U11893 (N_11893,N_9855,N_7505);
or U11894 (N_11894,N_7809,N_7216);
or U11895 (N_11895,N_5565,N_8682);
or U11896 (N_11896,N_6825,N_5972);
or U11897 (N_11897,N_8911,N_7089);
nor U11898 (N_11898,N_6835,N_8081);
or U11899 (N_11899,N_6047,N_8138);
nor U11900 (N_11900,N_7914,N_8940);
xor U11901 (N_11901,N_8465,N_6827);
and U11902 (N_11902,N_7607,N_7842);
nor U11903 (N_11903,N_6626,N_9023);
nor U11904 (N_11904,N_6824,N_7489);
nand U11905 (N_11905,N_6902,N_7124);
and U11906 (N_11906,N_6562,N_8453);
nor U11907 (N_11907,N_7025,N_5684);
xor U11908 (N_11908,N_9206,N_9578);
xnor U11909 (N_11909,N_7953,N_6963);
nand U11910 (N_11910,N_5894,N_9924);
nand U11911 (N_11911,N_6733,N_6799);
nor U11912 (N_11912,N_9573,N_9609);
xnor U11913 (N_11913,N_7060,N_7688);
and U11914 (N_11914,N_5415,N_7282);
nor U11915 (N_11915,N_9762,N_8266);
or U11916 (N_11916,N_6845,N_7510);
xor U11917 (N_11917,N_5869,N_8888);
or U11918 (N_11918,N_8715,N_8076);
or U11919 (N_11919,N_6441,N_5214);
nor U11920 (N_11920,N_8800,N_9972);
and U11921 (N_11921,N_8222,N_8981);
and U11922 (N_11922,N_5525,N_7923);
nor U11923 (N_11923,N_5081,N_7522);
xor U11924 (N_11924,N_9721,N_5570);
xnor U11925 (N_11925,N_7352,N_6810);
xor U11926 (N_11926,N_6614,N_9172);
and U11927 (N_11927,N_8231,N_7274);
nor U11928 (N_11928,N_9428,N_8843);
nor U11929 (N_11929,N_7103,N_8318);
nand U11930 (N_11930,N_8789,N_9691);
xor U11931 (N_11931,N_6764,N_5349);
and U11932 (N_11932,N_6622,N_7756);
xor U11933 (N_11933,N_6490,N_9383);
and U11934 (N_11934,N_5190,N_6187);
nand U11935 (N_11935,N_6156,N_9622);
xor U11936 (N_11936,N_7330,N_6749);
or U11937 (N_11937,N_5021,N_7845);
nand U11938 (N_11938,N_9158,N_9135);
and U11939 (N_11939,N_8590,N_9086);
xor U11940 (N_11940,N_5013,N_7325);
nor U11941 (N_11941,N_7318,N_8371);
xnor U11942 (N_11942,N_6779,N_7475);
nand U11943 (N_11943,N_7220,N_8941);
nand U11944 (N_11944,N_7051,N_9223);
nand U11945 (N_11945,N_7961,N_9791);
xor U11946 (N_11946,N_6556,N_8104);
xnor U11947 (N_11947,N_5715,N_5487);
or U11948 (N_11948,N_8235,N_8982);
nor U11949 (N_11949,N_7250,N_6005);
nand U11950 (N_11950,N_5284,N_8497);
and U11951 (N_11951,N_5921,N_7398);
and U11952 (N_11952,N_8398,N_7792);
xor U11953 (N_11953,N_7171,N_7588);
and U11954 (N_11954,N_9772,N_6998);
nor U11955 (N_11955,N_8866,N_5637);
or U11956 (N_11956,N_6008,N_8312);
or U11957 (N_11957,N_7125,N_7357);
nor U11958 (N_11958,N_9471,N_7850);
or U11959 (N_11959,N_9536,N_9214);
and U11960 (N_11960,N_9960,N_8418);
nor U11961 (N_11961,N_7701,N_9139);
and U11962 (N_11962,N_6475,N_9890);
and U11963 (N_11963,N_5651,N_5935);
or U11964 (N_11964,N_7454,N_5944);
nor U11965 (N_11965,N_5872,N_5017);
or U11966 (N_11966,N_5906,N_7277);
and U11967 (N_11967,N_6772,N_5035);
or U11968 (N_11968,N_9491,N_5790);
nor U11969 (N_11969,N_5532,N_5950);
nor U11970 (N_11970,N_8935,N_8044);
nor U11971 (N_11971,N_5028,N_8690);
nor U11972 (N_11972,N_7936,N_7734);
nand U11973 (N_11973,N_6405,N_6830);
and U11974 (N_11974,N_5682,N_8047);
nand U11975 (N_11975,N_7364,N_8095);
or U11976 (N_11976,N_8035,N_5398);
nor U11977 (N_11977,N_9954,N_6552);
nor U11978 (N_11978,N_8490,N_7294);
and U11979 (N_11979,N_6241,N_5536);
nor U11980 (N_11980,N_7017,N_8436);
nand U11981 (N_11981,N_9917,N_9602);
xnor U11982 (N_11982,N_6459,N_7787);
nor U11983 (N_11983,N_7476,N_5154);
or U11984 (N_11984,N_8206,N_6821);
nor U11985 (N_11985,N_5970,N_7833);
and U11986 (N_11986,N_5556,N_5221);
nor U11987 (N_11987,N_5866,N_6278);
or U11988 (N_11988,N_8474,N_8168);
xor U11989 (N_11989,N_9110,N_7183);
nand U11990 (N_11990,N_6601,N_9438);
nor U11991 (N_11991,N_9251,N_5600);
xor U11992 (N_11992,N_5634,N_6909);
nand U11993 (N_11993,N_9941,N_9810);
or U11994 (N_11994,N_8515,N_9861);
nand U11995 (N_11995,N_8195,N_6613);
nand U11996 (N_11996,N_6297,N_6616);
or U11997 (N_11997,N_7434,N_9460);
nor U11998 (N_11998,N_6695,N_5720);
nor U11999 (N_11999,N_9889,N_6313);
or U12000 (N_12000,N_8735,N_5947);
and U12001 (N_12001,N_5409,N_5096);
or U12002 (N_12002,N_5856,N_9301);
or U12003 (N_12003,N_7893,N_9695);
and U12004 (N_12004,N_8871,N_5410);
or U12005 (N_12005,N_9666,N_5358);
and U12006 (N_12006,N_7921,N_7338);
nand U12007 (N_12007,N_8246,N_8612);
xnor U12008 (N_12008,N_8247,N_5714);
nand U12009 (N_12009,N_5886,N_8458);
nand U12010 (N_12010,N_7513,N_5979);
nor U12011 (N_12011,N_5097,N_7624);
nor U12012 (N_12012,N_5846,N_5877);
nand U12013 (N_12013,N_7544,N_5134);
xor U12014 (N_12014,N_7548,N_6371);
or U12015 (N_12015,N_7324,N_8961);
nor U12016 (N_12016,N_6854,N_6455);
or U12017 (N_12017,N_5773,N_9526);
nand U12018 (N_12018,N_7661,N_6788);
and U12019 (N_12019,N_9318,N_5858);
xnor U12020 (N_12020,N_8038,N_5704);
or U12021 (N_12021,N_9836,N_7207);
nand U12022 (N_12022,N_9408,N_9347);
or U12023 (N_12023,N_9757,N_7896);
nor U12024 (N_12024,N_5059,N_9376);
nand U12025 (N_12025,N_6160,N_5149);
nor U12026 (N_12026,N_7251,N_8680);
nor U12027 (N_12027,N_5653,N_7742);
nand U12028 (N_12028,N_5814,N_9780);
xnor U12029 (N_12029,N_9431,N_8234);
and U12030 (N_12030,N_7875,N_5299);
and U12031 (N_12031,N_9877,N_7556);
and U12032 (N_12032,N_5524,N_8749);
xor U12033 (N_12033,N_9634,N_9002);
and U12034 (N_12034,N_6493,N_6264);
and U12035 (N_12035,N_9520,N_7185);
or U12036 (N_12036,N_6831,N_8401);
nand U12037 (N_12037,N_7718,N_7723);
xnor U12038 (N_12038,N_6544,N_8997);
xor U12039 (N_12039,N_5633,N_9016);
nor U12040 (N_12040,N_5529,N_5576);
nand U12041 (N_12041,N_9862,N_7429);
nand U12042 (N_12042,N_6324,N_6030);
and U12043 (N_12043,N_6844,N_8451);
and U12044 (N_12044,N_7042,N_6436);
nand U12045 (N_12045,N_9948,N_9900);
xor U12046 (N_12046,N_7068,N_8933);
nor U12047 (N_12047,N_6565,N_8561);
and U12048 (N_12048,N_6035,N_7023);
nand U12049 (N_12049,N_9626,N_9053);
xnor U12050 (N_12050,N_8100,N_5710);
or U12051 (N_12051,N_5352,N_7474);
xnor U12052 (N_12052,N_8218,N_9103);
xor U12053 (N_12053,N_9499,N_9136);
and U12054 (N_12054,N_9380,N_5282);
or U12055 (N_12055,N_5517,N_9325);
nor U12056 (N_12056,N_7710,N_5648);
nor U12057 (N_12057,N_8895,N_8331);
xor U12058 (N_12058,N_8819,N_5241);
and U12059 (N_12059,N_5617,N_7403);
nor U12060 (N_12060,N_5381,N_8450);
or U12061 (N_12061,N_6710,N_9974);
nand U12062 (N_12062,N_8174,N_7432);
xnor U12063 (N_12063,N_8619,N_8606);
nor U12064 (N_12064,N_6322,N_9076);
nor U12065 (N_12065,N_8082,N_8101);
or U12066 (N_12066,N_6450,N_7820);
nand U12067 (N_12067,N_6110,N_6214);
nand U12068 (N_12068,N_7290,N_6491);
and U12069 (N_12069,N_9846,N_8627);
nand U12070 (N_12070,N_5062,N_7534);
nand U12071 (N_12071,N_5568,N_5155);
nor U12072 (N_12072,N_8510,N_5143);
nand U12073 (N_12073,N_8661,N_9746);
xor U12074 (N_12074,N_6922,N_8077);
nor U12075 (N_12075,N_9287,N_6091);
or U12076 (N_12076,N_6009,N_5296);
nand U12077 (N_12077,N_6680,N_5145);
and U12078 (N_12078,N_7683,N_6512);
or U12079 (N_12079,N_8514,N_7460);
xor U12080 (N_12080,N_6082,N_6712);
nor U12081 (N_12081,N_7253,N_8086);
nand U12082 (N_12082,N_7419,N_9668);
xor U12083 (N_12083,N_5091,N_6427);
xnor U12084 (N_12084,N_6076,N_6270);
xnor U12085 (N_12085,N_8388,N_5014);
xnor U12086 (N_12086,N_7871,N_9988);
xor U12087 (N_12087,N_9802,N_6983);
nor U12088 (N_12088,N_8792,N_5954);
and U12089 (N_12089,N_8552,N_8444);
xnor U12090 (N_12090,N_8519,N_8696);
xnor U12091 (N_12091,N_8647,N_5481);
nor U12092 (N_12092,N_8368,N_5955);
and U12093 (N_12093,N_7367,N_6363);
xnor U12094 (N_12094,N_7852,N_5457);
nand U12095 (N_12095,N_6219,N_6892);
xnor U12096 (N_12096,N_5103,N_5647);
nor U12097 (N_12097,N_8072,N_9423);
or U12098 (N_12098,N_8855,N_5873);
or U12099 (N_12099,N_7669,N_7079);
xor U12100 (N_12100,N_5461,N_7578);
nor U12101 (N_12101,N_6533,N_8692);
nand U12102 (N_12102,N_5151,N_8913);
and U12103 (N_12103,N_9790,N_7237);
and U12104 (N_12104,N_5341,N_7670);
nor U12105 (N_12105,N_6846,N_6540);
and U12106 (N_12106,N_6096,N_7828);
xor U12107 (N_12107,N_6882,N_9700);
or U12108 (N_12108,N_6239,N_6582);
xor U12109 (N_12109,N_8089,N_9942);
and U12110 (N_12110,N_5387,N_8653);
nor U12111 (N_12111,N_7989,N_7319);
and U12112 (N_12112,N_6374,N_7811);
nor U12113 (N_12113,N_5249,N_5301);
nor U12114 (N_12114,N_5026,N_9868);
nand U12115 (N_12115,N_7406,N_5339);
and U12116 (N_12116,N_8870,N_5212);
or U12117 (N_12117,N_9317,N_9157);
xnor U12118 (N_12118,N_7444,N_7049);
xnor U12119 (N_12119,N_8141,N_6237);
or U12120 (N_12120,N_7468,N_6500);
nand U12121 (N_12121,N_6407,N_5632);
xnor U12122 (N_12122,N_9554,N_6604);
nor U12123 (N_12123,N_9290,N_6173);
and U12124 (N_12124,N_6361,N_5959);
and U12125 (N_12125,N_8525,N_8476);
xnor U12126 (N_12126,N_6080,N_6355);
and U12127 (N_12127,N_8583,N_8927);
nor U12128 (N_12128,N_5031,N_6603);
and U12129 (N_12129,N_5606,N_9183);
and U12130 (N_12130,N_5000,N_7409);
or U12131 (N_12131,N_5764,N_9465);
or U12132 (N_12132,N_8211,N_5599);
and U12133 (N_12133,N_7776,N_5178);
or U12134 (N_12134,N_8998,N_7879);
nor U12135 (N_12135,N_8902,N_7555);
or U12136 (N_12136,N_7658,N_8130);
or U12137 (N_12137,N_8210,N_7376);
or U12138 (N_12138,N_6046,N_7892);
xor U12139 (N_12139,N_6943,N_5566);
and U12140 (N_12140,N_8505,N_9752);
nand U12141 (N_12141,N_7823,N_7412);
or U12142 (N_12142,N_6049,N_6741);
nand U12143 (N_12143,N_8748,N_7930);
xor U12144 (N_12144,N_6479,N_5821);
nand U12145 (N_12145,N_7050,N_7008);
or U12146 (N_12146,N_9745,N_7947);
and U12147 (N_12147,N_8993,N_8355);
xnor U12148 (N_12148,N_7218,N_8589);
nand U12149 (N_12149,N_7063,N_5464);
xnor U12150 (N_12150,N_6132,N_9338);
nand U12151 (N_12151,N_5747,N_6560);
or U12152 (N_12152,N_5049,N_6919);
xnor U12153 (N_12153,N_7308,N_5085);
nand U12154 (N_12154,N_9712,N_9611);
and U12155 (N_12155,N_7593,N_5276);
or U12156 (N_12156,N_8783,N_8242);
or U12157 (N_12157,N_9607,N_6012);
or U12158 (N_12158,N_7000,N_8447);
nand U12159 (N_12159,N_7349,N_8014);
nand U12160 (N_12160,N_8315,N_7138);
nand U12161 (N_12161,N_6662,N_8021);
and U12162 (N_12162,N_6037,N_6912);
nor U12163 (N_12163,N_7235,N_8667);
and U12164 (N_12164,N_6184,N_6443);
xnor U12165 (N_12165,N_7524,N_8761);
or U12166 (N_12166,N_8105,N_7694);
nor U12167 (N_12167,N_5309,N_9133);
nor U12168 (N_12168,N_7912,N_7172);
or U12169 (N_12169,N_7798,N_7521);
xnor U12170 (N_12170,N_7480,N_8261);
and U12171 (N_12171,N_8848,N_9913);
nor U12172 (N_12172,N_9468,N_7619);
xor U12173 (N_12173,N_7758,N_7726);
and U12174 (N_12174,N_6431,N_7016);
nand U12175 (N_12175,N_7714,N_8850);
or U12176 (N_12176,N_5227,N_9137);
and U12177 (N_12177,N_5372,N_5640);
xor U12178 (N_12178,N_5534,N_6048);
and U12179 (N_12179,N_5259,N_8280);
xnor U12180 (N_12180,N_5274,N_6993);
or U12181 (N_12181,N_6343,N_6061);
or U12182 (N_12182,N_8859,N_8938);
nor U12183 (N_12183,N_5851,N_5060);
nand U12184 (N_12184,N_6300,N_9709);
xor U12185 (N_12185,N_7941,N_5416);
nor U12186 (N_12186,N_6889,N_9758);
nand U12187 (N_12187,N_6460,N_7981);
and U12188 (N_12188,N_7864,N_9247);
and U12189 (N_12189,N_5459,N_9043);
and U12190 (N_12190,N_5552,N_6941);
or U12191 (N_12191,N_5531,N_5236);
nor U12192 (N_12192,N_8455,N_9732);
xnor U12193 (N_12193,N_9289,N_9424);
nor U12194 (N_12194,N_9649,N_7012);
and U12195 (N_12195,N_6366,N_9911);
nand U12196 (N_12196,N_9111,N_6644);
nor U12197 (N_12197,N_5916,N_7018);
nor U12198 (N_12198,N_7554,N_5562);
and U12199 (N_12199,N_6867,N_9451);
nor U12200 (N_12200,N_6131,N_9583);
nand U12201 (N_12201,N_5727,N_5492);
nand U12202 (N_12202,N_7853,N_9537);
nor U12203 (N_12203,N_8953,N_5338);
nor U12204 (N_12204,N_5315,N_5569);
xnor U12205 (N_12205,N_7128,N_5815);
and U12206 (N_12206,N_9480,N_6192);
xnor U12207 (N_12207,N_8161,N_6088);
or U12208 (N_12208,N_7819,N_7596);
nor U12209 (N_12209,N_7486,N_7958);
and U12210 (N_12210,N_7610,N_6031);
nor U12211 (N_12211,N_7780,N_7739);
or U12212 (N_12212,N_9233,N_5048);
xor U12213 (N_12213,N_7200,N_9349);
nand U12214 (N_12214,N_6135,N_5501);
and U12215 (N_12215,N_9542,N_5986);
nand U12216 (N_12216,N_7576,N_7211);
xor U12217 (N_12217,N_6223,N_8187);
nor U12218 (N_12218,N_9970,N_9476);
nand U12219 (N_12219,N_6877,N_6964);
and U12220 (N_12220,N_8898,N_7984);
nand U12221 (N_12221,N_6351,N_7663);
nand U12222 (N_12222,N_5141,N_6957);
or U12223 (N_12223,N_9312,N_8652);
and U12224 (N_12224,N_6701,N_6742);
nand U12225 (N_12225,N_5540,N_9435);
and U12226 (N_12226,N_7437,N_9222);
xor U12227 (N_12227,N_6689,N_5839);
or U12228 (N_12228,N_5426,N_8156);
nand U12229 (N_12229,N_7100,N_9560);
or U12230 (N_12230,N_8193,N_7301);
or U12231 (N_12231,N_9840,N_6974);
nor U12232 (N_12232,N_6318,N_7381);
and U12233 (N_12233,N_9817,N_6176);
nand U12234 (N_12234,N_8890,N_6305);
or U12235 (N_12235,N_6572,N_6304);
xnor U12236 (N_12236,N_6461,N_6205);
and U12237 (N_12237,N_5659,N_5240);
nand U12238 (N_12238,N_9624,N_8620);
nand U12239 (N_12239,N_9879,N_8364);
nor U12240 (N_12240,N_6240,N_9690);
and U12241 (N_12241,N_6335,N_6899);
or U12242 (N_12242,N_9291,N_7939);
xor U12243 (N_12243,N_8582,N_7191);
nand U12244 (N_12244,N_6381,N_5129);
nand U12245 (N_12245,N_8699,N_8477);
nand U12246 (N_12246,N_5698,N_6480);
nor U12247 (N_12247,N_9747,N_5677);
nor U12248 (N_12248,N_6295,N_5262);
nor U12249 (N_12249,N_8823,N_7488);
or U12250 (N_12250,N_9689,N_8201);
xnor U12251 (N_12251,N_9008,N_8373);
or U12252 (N_12252,N_7538,N_7746);
nor U12253 (N_12253,N_8233,N_5514);
or U12254 (N_12254,N_9882,N_5167);
or U12255 (N_12255,N_6388,N_7550);
and U12256 (N_12256,N_9774,N_8868);
nand U12257 (N_12257,N_6522,N_8664);
nor U12258 (N_12258,N_8030,N_5225);
xor U12259 (N_12259,N_6696,N_6166);
nand U12260 (N_12260,N_7400,N_6045);
xor U12261 (N_12261,N_6874,N_7743);
or U12262 (N_12262,N_8277,N_9831);
or U12263 (N_12263,N_6881,N_6111);
nand U12264 (N_12264,N_9703,N_7563);
xor U12265 (N_12265,N_8718,N_7866);
and U12266 (N_12266,N_7684,N_8932);
nor U12267 (N_12267,N_8731,N_8307);
nand U12268 (N_12268,N_5310,N_7221);
nand U12269 (N_12269,N_7496,N_8670);
or U12270 (N_12270,N_9077,N_8471);
and U12271 (N_12271,N_8460,N_8881);
xor U12272 (N_12272,N_6384,N_7662);
xnor U12273 (N_12273,N_5563,N_9230);
and U12274 (N_12274,N_7140,N_6734);
nor U12275 (N_12275,N_7045,N_8980);
xor U12276 (N_12276,N_8909,N_8849);
and U12277 (N_12277,N_9992,N_8199);
nor U12278 (N_12278,N_8298,N_7919);
xor U12279 (N_12279,N_7724,N_6202);
nand U12280 (N_12280,N_8600,N_6850);
or U12281 (N_12281,N_8139,N_5425);
nand U12282 (N_12282,N_6182,N_6298);
xor U12283 (N_12283,N_7252,N_8760);
xor U12284 (N_12284,N_9956,N_9723);
or U12285 (N_12285,N_8405,N_9193);
or U12286 (N_12286,N_7614,N_7849);
or U12287 (N_12287,N_5796,N_6314);
or U12288 (N_12288,N_9765,N_5104);
nor U12289 (N_12289,N_7888,N_6022);
and U12290 (N_12290,N_8697,N_7471);
or U12291 (N_12291,N_9400,N_5579);
nand U12292 (N_12292,N_9253,N_9346);
and U12293 (N_12293,N_7602,N_5303);
nand U12294 (N_12294,N_7445,N_6272);
nand U12295 (N_12295,N_9813,N_9977);
or U12296 (N_12296,N_7986,N_8304);
and U12297 (N_12297,N_5173,N_5316);
nand U12298 (N_12298,N_9863,N_7462);
or U12299 (N_12299,N_5297,N_8947);
nor U12300 (N_12300,N_9806,N_9528);
nor U12301 (N_12301,N_9482,N_5158);
nand U12302 (N_12302,N_8986,N_6841);
xnor U12303 (N_12303,N_7648,N_8273);
nand U12304 (N_12304,N_5357,N_7630);
xnor U12305 (N_12305,N_8411,N_6222);
xor U12306 (N_12306,N_8228,N_8216);
nand U12307 (N_12307,N_7832,N_7716);
nand U12308 (N_12308,N_6044,N_7711);
or U12309 (N_12309,N_9610,N_6870);
nor U12310 (N_12310,N_7271,N_8992);
nand U12311 (N_12311,N_8541,N_8629);
xor U12312 (N_12312,N_5463,N_8166);
nor U12313 (N_12313,N_8751,N_9486);
xor U12314 (N_12314,N_8142,N_6979);
or U12315 (N_12315,N_5117,N_6796);
or U12316 (N_12316,N_6062,N_8407);
or U12317 (N_12317,N_9580,N_8330);
or U12318 (N_12318,N_9328,N_5254);
nand U12319 (N_12319,N_5766,N_9901);
xnor U12320 (N_12320,N_8498,N_9488);
nor U12321 (N_12321,N_5931,N_9562);
nor U12322 (N_12322,N_7304,N_9155);
nor U12323 (N_12323,N_6389,N_9540);
or U12324 (N_12324,N_7421,N_8963);
or U12325 (N_12325,N_7951,N_6034);
nand U12326 (N_12326,N_9069,N_6722);
nand U12327 (N_12327,N_8063,N_6169);
nor U12328 (N_12328,N_7146,N_7306);
xnor U12329 (N_12329,N_8754,N_7829);
xnor U12330 (N_12330,N_8271,N_5468);
nand U12331 (N_12331,N_8117,N_7314);
nand U12332 (N_12332,N_6103,N_5546);
nor U12333 (N_12333,N_9132,N_7224);
xnor U12334 (N_12334,N_9750,N_6154);
or U12335 (N_12335,N_5934,N_5587);
xor U12336 (N_12336,N_5654,N_5523);
nand U12337 (N_12337,N_7280,N_6853);
nand U12338 (N_12338,N_7418,N_8985);
xnor U12339 (N_12339,N_9928,N_8708);
or U12340 (N_12340,N_9796,N_9592);
nor U12341 (N_12341,N_5533,N_8346);
or U12342 (N_12342,N_9456,N_6376);
xnor U12343 (N_12343,N_6539,N_9793);
or U12344 (N_12344,N_9209,N_5835);
and U12345 (N_12345,N_7652,N_6426);
nand U12346 (N_12346,N_9120,N_5920);
and U12347 (N_12347,N_8759,N_9150);
and U12348 (N_12348,N_5586,N_9815);
or U12349 (N_12349,N_9784,N_6756);
or U12350 (N_12350,N_5235,N_6134);
nand U12351 (N_12351,N_5061,N_7291);
nor U12352 (N_12352,N_5609,N_6392);
xor U12353 (N_12353,N_9663,N_8249);
xnor U12354 (N_12354,N_5052,N_5771);
xnor U12355 (N_12355,N_5781,N_6836);
nand U12356 (N_12356,N_5286,N_7655);
nor U12357 (N_12357,N_6251,N_8524);
and U12358 (N_12358,N_7926,N_7764);
and U12359 (N_12359,N_8778,N_6703);
and U12360 (N_12360,N_6686,N_7487);
nand U12361 (N_12361,N_7072,N_9459);
or U12362 (N_12362,N_8610,N_7615);
nor U12363 (N_12363,N_5321,N_6025);
nand U12364 (N_12364,N_9422,N_6199);
nand U12365 (N_12365,N_7755,N_5949);
and U12366 (N_12366,N_9853,N_6911);
xor U12367 (N_12367,N_9068,N_6471);
xor U12368 (N_12368,N_8459,N_6393);
or U12369 (N_12369,N_6196,N_6040);
nand U12370 (N_12370,N_7937,N_5181);
or U12371 (N_12371,N_5248,N_7388);
or U12372 (N_12372,N_5467,N_8805);
nand U12373 (N_12373,N_7594,N_8024);
xor U12374 (N_12374,N_9543,N_5671);
xnor U12375 (N_12375,N_5887,N_6118);
nand U12376 (N_12376,N_6116,N_5824);
or U12377 (N_12377,N_9192,N_6739);
and U12378 (N_12378,N_8294,N_8603);
or U12379 (N_12379,N_5412,N_5477);
nand U12380 (N_12380,N_9090,N_8969);
nor U12381 (N_12381,N_6837,N_5631);
xor U12382 (N_12382,N_6513,N_7848);
xor U12383 (N_12383,N_8862,N_5435);
xor U12384 (N_12384,N_6636,N_9335);
and U12385 (N_12385,N_7539,N_7210);
nor U12386 (N_12386,N_5448,N_6605);
xor U12387 (N_12387,N_6673,N_7048);
xor U12388 (N_12388,N_8645,N_5320);
and U12389 (N_12389,N_8892,N_6631);
xor U12390 (N_12390,N_8547,N_6293);
nand U12391 (N_12391,N_5547,N_6528);
and U12392 (N_12392,N_6659,N_7865);
nand U12393 (N_12393,N_7821,N_9801);
xnor U12394 (N_12394,N_6839,N_8264);
nand U12395 (N_12395,N_7752,N_7283);
nand U12396 (N_12396,N_5388,N_7094);
nor U12397 (N_12397,N_5845,N_7890);
and U12398 (N_12398,N_9532,N_5490);
and U12399 (N_12399,N_7900,N_5663);
xor U12400 (N_12400,N_9324,N_8721);
nor U12401 (N_12401,N_8399,N_7631);
nand U12402 (N_12402,N_8979,N_8825);
nor U12403 (N_12403,N_8262,N_8308);
nand U12404 (N_12404,N_5889,N_9274);
and U12405 (N_12405,N_8559,N_9118);
xor U12406 (N_12406,N_9406,N_7452);
and U12407 (N_12407,N_9208,N_7503);
or U12408 (N_12408,N_9735,N_7915);
xor U12409 (N_12409,N_7370,N_7019);
or U12410 (N_12410,N_6356,N_9006);
and U12411 (N_12411,N_9556,N_6375);
or U12412 (N_12412,N_6781,N_5910);
and U12413 (N_12413,N_8025,N_8779);
xnor U12414 (N_12414,N_9998,N_7928);
nand U12415 (N_12415,N_8394,N_9186);
and U12416 (N_12416,N_7321,N_8774);
or U12417 (N_12417,N_6225,N_8516);
xor U12418 (N_12418,N_8414,N_8624);
or U12419 (N_12419,N_8050,N_6104);
or U12420 (N_12420,N_8704,N_5985);
and U12421 (N_12421,N_6953,N_7512);
xnor U12422 (N_12422,N_9071,N_7285);
or U12423 (N_12423,N_6462,N_8598);
and U12424 (N_12424,N_9822,N_6618);
nor U12425 (N_12425,N_5707,N_7999);
nand U12426 (N_12426,N_8500,N_7616);
xor U12427 (N_12427,N_6538,N_8333);
or U12428 (N_12428,N_5266,N_9980);
nand U12429 (N_12429,N_9968,N_5166);
or U12430 (N_12430,N_8306,N_5673);
and U12431 (N_12431,N_6675,N_9989);
nand U12432 (N_12432,N_5213,N_6584);
and U12433 (N_12433,N_8522,N_5549);
nand U12434 (N_12434,N_7895,N_6679);
xnor U12435 (N_12435,N_7592,N_5069);
or U12436 (N_12436,N_8164,N_7169);
nor U12437 (N_12437,N_8052,N_8090);
or U12438 (N_12438,N_5109,N_5070);
and U12439 (N_12439,N_5386,N_5938);
nand U12440 (N_12440,N_8293,N_9056);
nor U12441 (N_12441,N_7960,N_6669);
nand U12442 (N_12442,N_8058,N_9447);
nor U12443 (N_12443,N_5336,N_6369);
nor U12444 (N_12444,N_6256,N_9159);
xnor U12445 (N_12445,N_9635,N_8153);
nand U12446 (N_12446,N_6038,N_7987);
xnor U12447 (N_12447,N_8446,N_6578);
or U12448 (N_12448,N_9441,N_7287);
nor U12449 (N_12449,N_6608,N_6670);
and U12450 (N_12450,N_8068,N_5882);
nor U12451 (N_12451,N_6007,N_8554);
nor U12452 (N_12452,N_6121,N_5729);
nor U12453 (N_12453,N_5268,N_9769);
and U12454 (N_12454,N_9549,N_5197);
and U12455 (N_12455,N_5046,N_9684);
nand U12456 (N_12456,N_9187,N_8099);
xor U12457 (N_12457,N_5801,N_8845);
xor U12458 (N_12458,N_5504,N_5229);
nor U12459 (N_12459,N_5874,N_8492);
xnor U12460 (N_12460,N_5265,N_7104);
xor U12461 (N_12461,N_7493,N_7405);
and U12462 (N_12462,N_8146,N_6175);
nand U12463 (N_12463,N_8720,N_6929);
and U12464 (N_12464,N_8901,N_6164);
xnor U12465 (N_12465,N_8179,N_8535);
or U12466 (N_12466,N_9278,N_8382);
nand U12467 (N_12467,N_7061,N_5485);
or U12468 (N_12468,N_9260,N_7300);
xor U12469 (N_12469,N_7278,N_5200);
and U12470 (N_12470,N_6463,N_5380);
nor U12471 (N_12471,N_8360,N_7236);
xnor U12472 (N_12472,N_5420,N_9792);
or U12473 (N_12473,N_8291,N_5431);
xnor U12474 (N_12474,N_6065,N_6780);
nand U12475 (N_12475,N_8158,N_6563);
xor U12476 (N_12476,N_9731,N_6894);
nand U12477 (N_12477,N_7065,N_9606);
xor U12478 (N_12478,N_8175,N_8244);
or U12479 (N_12479,N_8005,N_8483);
xnor U12480 (N_12480,N_6944,N_9113);
nor U12481 (N_12481,N_7359,N_5010);
xor U12482 (N_12482,N_5140,N_6628);
xor U12483 (N_12483,N_5924,N_9715);
nor U12484 (N_12484,N_9162,N_8826);
or U12485 (N_12485,N_8251,N_5743);
nand U12486 (N_12486,N_6073,N_5323);
and U12487 (N_12487,N_7178,N_9084);
nor U12488 (N_12488,N_5508,N_8509);
nand U12489 (N_12489,N_9082,N_5404);
or U12490 (N_12490,N_6003,N_9986);
or U12491 (N_12491,N_9804,N_5554);
nand U12492 (N_12492,N_5509,N_8192);
xor U12493 (N_12493,N_6051,N_9558);
or U12494 (N_12494,N_6597,N_7963);
nor U12495 (N_12495,N_5391,N_7727);
and U12496 (N_12496,N_7645,N_9240);
or U12497 (N_12497,N_9326,N_7696);
nor U12498 (N_12498,N_8290,N_5277);
or U12499 (N_12499,N_9938,N_5973);
nor U12500 (N_12500,N_7895,N_6896);
xnor U12501 (N_12501,N_6236,N_8268);
nand U12502 (N_12502,N_6542,N_9783);
xor U12503 (N_12503,N_7842,N_7743);
or U12504 (N_12504,N_6226,N_6099);
nor U12505 (N_12505,N_5507,N_5155);
nand U12506 (N_12506,N_6727,N_9327);
or U12507 (N_12507,N_6155,N_9386);
nand U12508 (N_12508,N_5520,N_9766);
nor U12509 (N_12509,N_6262,N_8491);
or U12510 (N_12510,N_9813,N_7974);
nand U12511 (N_12511,N_7801,N_7423);
xnor U12512 (N_12512,N_9911,N_8323);
and U12513 (N_12513,N_8359,N_8377);
xor U12514 (N_12514,N_7711,N_5432);
and U12515 (N_12515,N_5027,N_7102);
nand U12516 (N_12516,N_7184,N_9375);
xnor U12517 (N_12517,N_6612,N_5090);
nor U12518 (N_12518,N_5919,N_5512);
nand U12519 (N_12519,N_9703,N_7609);
and U12520 (N_12520,N_7809,N_7456);
nand U12521 (N_12521,N_9008,N_9774);
and U12522 (N_12522,N_8777,N_6487);
or U12523 (N_12523,N_7236,N_6501);
xnor U12524 (N_12524,N_7421,N_9676);
and U12525 (N_12525,N_6198,N_6092);
or U12526 (N_12526,N_9825,N_9424);
nor U12527 (N_12527,N_8270,N_9299);
or U12528 (N_12528,N_5296,N_6606);
and U12529 (N_12529,N_5519,N_5318);
or U12530 (N_12530,N_9648,N_7118);
nand U12531 (N_12531,N_5947,N_9050);
and U12532 (N_12532,N_7280,N_5604);
nor U12533 (N_12533,N_6813,N_5930);
or U12534 (N_12534,N_9355,N_8484);
or U12535 (N_12535,N_5235,N_8357);
and U12536 (N_12536,N_5114,N_7888);
or U12537 (N_12537,N_7379,N_5698);
or U12538 (N_12538,N_9033,N_9064);
or U12539 (N_12539,N_7403,N_8940);
and U12540 (N_12540,N_6594,N_9112);
nand U12541 (N_12541,N_8917,N_7553);
xor U12542 (N_12542,N_7097,N_9779);
and U12543 (N_12543,N_5717,N_7875);
or U12544 (N_12544,N_6604,N_5553);
nor U12545 (N_12545,N_8063,N_5148);
nor U12546 (N_12546,N_7764,N_6633);
or U12547 (N_12547,N_9887,N_7423);
and U12548 (N_12548,N_9078,N_7581);
nor U12549 (N_12549,N_6284,N_9171);
xnor U12550 (N_12550,N_9307,N_5130);
nand U12551 (N_12551,N_5446,N_6508);
and U12552 (N_12552,N_7054,N_9161);
or U12553 (N_12553,N_6884,N_5513);
nor U12554 (N_12554,N_7415,N_6372);
and U12555 (N_12555,N_5086,N_7713);
and U12556 (N_12556,N_9795,N_7884);
nand U12557 (N_12557,N_9175,N_9833);
nand U12558 (N_12558,N_9796,N_5106);
or U12559 (N_12559,N_6019,N_9249);
xnor U12560 (N_12560,N_7774,N_9237);
and U12561 (N_12561,N_8189,N_6819);
xnor U12562 (N_12562,N_6595,N_8385);
nor U12563 (N_12563,N_7193,N_6425);
nand U12564 (N_12564,N_8562,N_8790);
and U12565 (N_12565,N_8647,N_6611);
nand U12566 (N_12566,N_7772,N_9578);
xor U12567 (N_12567,N_6944,N_7993);
nand U12568 (N_12568,N_9861,N_8618);
and U12569 (N_12569,N_7867,N_5997);
and U12570 (N_12570,N_5762,N_6985);
xnor U12571 (N_12571,N_6128,N_8461);
and U12572 (N_12572,N_6934,N_6796);
or U12573 (N_12573,N_9198,N_8008);
and U12574 (N_12574,N_8499,N_7036);
xor U12575 (N_12575,N_8836,N_8278);
xor U12576 (N_12576,N_7284,N_6737);
nand U12577 (N_12577,N_5820,N_7935);
nand U12578 (N_12578,N_7185,N_7113);
and U12579 (N_12579,N_7978,N_7019);
nand U12580 (N_12580,N_6411,N_7900);
or U12581 (N_12581,N_9193,N_7424);
nor U12582 (N_12582,N_5307,N_6861);
and U12583 (N_12583,N_8720,N_7473);
nand U12584 (N_12584,N_7772,N_5475);
nor U12585 (N_12585,N_7768,N_9726);
nor U12586 (N_12586,N_9103,N_7674);
nand U12587 (N_12587,N_7366,N_9810);
or U12588 (N_12588,N_5766,N_8202);
nor U12589 (N_12589,N_8511,N_5420);
and U12590 (N_12590,N_8538,N_9704);
nor U12591 (N_12591,N_6130,N_8806);
and U12592 (N_12592,N_6798,N_5228);
nor U12593 (N_12593,N_7155,N_7167);
nor U12594 (N_12594,N_6001,N_9042);
and U12595 (N_12595,N_6389,N_8028);
and U12596 (N_12596,N_8506,N_9766);
or U12597 (N_12597,N_7691,N_6204);
and U12598 (N_12598,N_8268,N_9295);
nand U12599 (N_12599,N_9176,N_5411);
nand U12600 (N_12600,N_8638,N_7795);
or U12601 (N_12601,N_9896,N_7324);
xnor U12602 (N_12602,N_5162,N_9124);
or U12603 (N_12603,N_7233,N_8418);
nand U12604 (N_12604,N_7026,N_9185);
nand U12605 (N_12605,N_7934,N_8308);
or U12606 (N_12606,N_8756,N_6971);
nor U12607 (N_12607,N_8087,N_5861);
nor U12608 (N_12608,N_9259,N_8262);
xnor U12609 (N_12609,N_7710,N_8701);
nor U12610 (N_12610,N_8143,N_9739);
xor U12611 (N_12611,N_6076,N_5925);
and U12612 (N_12612,N_5480,N_5058);
xor U12613 (N_12613,N_6275,N_9160);
nor U12614 (N_12614,N_5829,N_8677);
nor U12615 (N_12615,N_8100,N_8040);
nand U12616 (N_12616,N_6864,N_7817);
and U12617 (N_12617,N_5245,N_6015);
nor U12618 (N_12618,N_7889,N_6044);
or U12619 (N_12619,N_5698,N_5031);
or U12620 (N_12620,N_8203,N_5280);
and U12621 (N_12621,N_5856,N_5360);
nor U12622 (N_12622,N_9996,N_5553);
and U12623 (N_12623,N_6036,N_7841);
or U12624 (N_12624,N_7656,N_7983);
nand U12625 (N_12625,N_6809,N_9908);
or U12626 (N_12626,N_7093,N_6415);
nand U12627 (N_12627,N_9282,N_9406);
or U12628 (N_12628,N_9164,N_8354);
and U12629 (N_12629,N_5376,N_7692);
or U12630 (N_12630,N_8114,N_7196);
nor U12631 (N_12631,N_5592,N_9887);
xnor U12632 (N_12632,N_6625,N_7258);
nor U12633 (N_12633,N_6299,N_7564);
or U12634 (N_12634,N_5023,N_7370);
or U12635 (N_12635,N_8444,N_8517);
and U12636 (N_12636,N_8498,N_6459);
nand U12637 (N_12637,N_7938,N_6910);
nor U12638 (N_12638,N_6615,N_6794);
xnor U12639 (N_12639,N_8302,N_5268);
or U12640 (N_12640,N_9067,N_5658);
or U12641 (N_12641,N_8587,N_6653);
xnor U12642 (N_12642,N_5454,N_8713);
nand U12643 (N_12643,N_5490,N_8714);
nand U12644 (N_12644,N_9155,N_6961);
nor U12645 (N_12645,N_5866,N_8412);
nand U12646 (N_12646,N_9139,N_8507);
nand U12647 (N_12647,N_5028,N_7946);
xor U12648 (N_12648,N_5129,N_6984);
or U12649 (N_12649,N_5270,N_9295);
nand U12650 (N_12650,N_5950,N_6653);
nand U12651 (N_12651,N_5546,N_6343);
or U12652 (N_12652,N_7435,N_8188);
xnor U12653 (N_12653,N_7511,N_5679);
xor U12654 (N_12654,N_8864,N_9525);
nor U12655 (N_12655,N_8790,N_8254);
or U12656 (N_12656,N_6476,N_6083);
nor U12657 (N_12657,N_9139,N_7748);
nand U12658 (N_12658,N_5982,N_8497);
nor U12659 (N_12659,N_7266,N_6855);
xor U12660 (N_12660,N_5741,N_6209);
nor U12661 (N_12661,N_5131,N_7740);
xnor U12662 (N_12662,N_6315,N_9190);
nand U12663 (N_12663,N_8332,N_6528);
xor U12664 (N_12664,N_7342,N_8211);
nor U12665 (N_12665,N_6454,N_9734);
nand U12666 (N_12666,N_5059,N_5767);
xnor U12667 (N_12667,N_5462,N_6440);
nand U12668 (N_12668,N_5272,N_9214);
nor U12669 (N_12669,N_8402,N_9597);
and U12670 (N_12670,N_6650,N_5443);
or U12671 (N_12671,N_9702,N_8730);
nand U12672 (N_12672,N_6791,N_7992);
and U12673 (N_12673,N_5560,N_9826);
and U12674 (N_12674,N_8409,N_8830);
xnor U12675 (N_12675,N_6576,N_9923);
and U12676 (N_12676,N_8352,N_7156);
and U12677 (N_12677,N_7037,N_6028);
nor U12678 (N_12678,N_8716,N_6887);
nor U12679 (N_12679,N_8155,N_6968);
and U12680 (N_12680,N_5043,N_5530);
or U12681 (N_12681,N_6987,N_8781);
nand U12682 (N_12682,N_7454,N_5473);
or U12683 (N_12683,N_9116,N_5367);
nand U12684 (N_12684,N_6819,N_8562);
nor U12685 (N_12685,N_6469,N_5240);
nand U12686 (N_12686,N_8309,N_7168);
nand U12687 (N_12687,N_6538,N_5129);
nor U12688 (N_12688,N_5848,N_9037);
xnor U12689 (N_12689,N_9915,N_6256);
nor U12690 (N_12690,N_5550,N_8740);
xor U12691 (N_12691,N_5223,N_9010);
and U12692 (N_12692,N_8435,N_7741);
and U12693 (N_12693,N_5471,N_5290);
nand U12694 (N_12694,N_6002,N_8532);
or U12695 (N_12695,N_5586,N_9215);
or U12696 (N_12696,N_6085,N_6763);
or U12697 (N_12697,N_7242,N_8722);
nand U12698 (N_12698,N_5128,N_6246);
nor U12699 (N_12699,N_9351,N_9912);
nor U12700 (N_12700,N_8821,N_5311);
nor U12701 (N_12701,N_7395,N_8452);
and U12702 (N_12702,N_5455,N_7064);
or U12703 (N_12703,N_5269,N_9969);
or U12704 (N_12704,N_5554,N_6235);
nand U12705 (N_12705,N_9802,N_7273);
nand U12706 (N_12706,N_9145,N_8478);
and U12707 (N_12707,N_7752,N_8405);
nor U12708 (N_12708,N_9937,N_7246);
and U12709 (N_12709,N_6500,N_5040);
xor U12710 (N_12710,N_9358,N_7251);
xnor U12711 (N_12711,N_9374,N_7770);
or U12712 (N_12712,N_9714,N_7851);
xnor U12713 (N_12713,N_6491,N_9564);
and U12714 (N_12714,N_8273,N_9195);
nor U12715 (N_12715,N_8911,N_7619);
and U12716 (N_12716,N_5660,N_5733);
nor U12717 (N_12717,N_6146,N_7200);
xor U12718 (N_12718,N_7196,N_7479);
or U12719 (N_12719,N_7012,N_5419);
xnor U12720 (N_12720,N_8973,N_6889);
nor U12721 (N_12721,N_8301,N_7125);
and U12722 (N_12722,N_5482,N_7437);
and U12723 (N_12723,N_8261,N_9175);
or U12724 (N_12724,N_5560,N_7220);
and U12725 (N_12725,N_6153,N_6220);
nor U12726 (N_12726,N_9306,N_5105);
xnor U12727 (N_12727,N_7496,N_6738);
xor U12728 (N_12728,N_8673,N_6074);
xnor U12729 (N_12729,N_6103,N_9402);
and U12730 (N_12730,N_5920,N_8354);
xor U12731 (N_12731,N_9863,N_6554);
and U12732 (N_12732,N_7978,N_5035);
nand U12733 (N_12733,N_9725,N_6767);
nor U12734 (N_12734,N_8011,N_6796);
xnor U12735 (N_12735,N_9994,N_7964);
xnor U12736 (N_12736,N_8809,N_5208);
nand U12737 (N_12737,N_7503,N_7316);
and U12738 (N_12738,N_6390,N_5065);
nor U12739 (N_12739,N_5832,N_7620);
nand U12740 (N_12740,N_5172,N_8747);
xor U12741 (N_12741,N_5221,N_7922);
nor U12742 (N_12742,N_6913,N_7319);
nor U12743 (N_12743,N_5599,N_8771);
and U12744 (N_12744,N_8037,N_6823);
or U12745 (N_12745,N_9926,N_9002);
nand U12746 (N_12746,N_9764,N_9190);
nor U12747 (N_12747,N_8819,N_7070);
nand U12748 (N_12748,N_8246,N_6539);
xor U12749 (N_12749,N_5261,N_9335);
and U12750 (N_12750,N_9814,N_9279);
and U12751 (N_12751,N_9039,N_8974);
nor U12752 (N_12752,N_9127,N_5995);
or U12753 (N_12753,N_5973,N_6022);
nor U12754 (N_12754,N_8183,N_6785);
or U12755 (N_12755,N_9799,N_5662);
nor U12756 (N_12756,N_7130,N_7434);
nor U12757 (N_12757,N_9656,N_7080);
and U12758 (N_12758,N_5642,N_8543);
nor U12759 (N_12759,N_7789,N_6701);
nor U12760 (N_12760,N_6460,N_8826);
or U12761 (N_12761,N_5496,N_5924);
nand U12762 (N_12762,N_7736,N_7595);
xnor U12763 (N_12763,N_6040,N_8534);
or U12764 (N_12764,N_5957,N_8246);
and U12765 (N_12765,N_7413,N_5723);
xnor U12766 (N_12766,N_8084,N_6896);
nand U12767 (N_12767,N_8535,N_8109);
and U12768 (N_12768,N_6331,N_8310);
and U12769 (N_12769,N_6398,N_8574);
nand U12770 (N_12770,N_5204,N_8922);
xnor U12771 (N_12771,N_5821,N_9749);
xor U12772 (N_12772,N_9927,N_9672);
nor U12773 (N_12773,N_7034,N_5037);
xor U12774 (N_12774,N_8781,N_7499);
nor U12775 (N_12775,N_6656,N_5372);
xnor U12776 (N_12776,N_9357,N_5515);
nand U12777 (N_12777,N_7976,N_8016);
xor U12778 (N_12778,N_9540,N_9389);
or U12779 (N_12779,N_7712,N_8114);
or U12780 (N_12780,N_7979,N_8033);
nand U12781 (N_12781,N_8511,N_6783);
nand U12782 (N_12782,N_9635,N_5156);
nand U12783 (N_12783,N_7856,N_6061);
nand U12784 (N_12784,N_8829,N_8344);
and U12785 (N_12785,N_9881,N_5542);
nand U12786 (N_12786,N_8779,N_7569);
or U12787 (N_12787,N_6235,N_5176);
and U12788 (N_12788,N_5938,N_5213);
nand U12789 (N_12789,N_5443,N_6037);
and U12790 (N_12790,N_9300,N_9562);
nand U12791 (N_12791,N_8684,N_5637);
nand U12792 (N_12792,N_8761,N_7362);
xnor U12793 (N_12793,N_9944,N_5159);
nand U12794 (N_12794,N_8998,N_5472);
nand U12795 (N_12795,N_6360,N_9126);
xnor U12796 (N_12796,N_6191,N_5406);
nand U12797 (N_12797,N_9729,N_5935);
nand U12798 (N_12798,N_9354,N_8551);
and U12799 (N_12799,N_8520,N_8156);
and U12800 (N_12800,N_8797,N_6867);
nor U12801 (N_12801,N_5807,N_7259);
nand U12802 (N_12802,N_8325,N_6511);
nor U12803 (N_12803,N_7634,N_9111);
and U12804 (N_12804,N_5328,N_8072);
nor U12805 (N_12805,N_9137,N_8038);
or U12806 (N_12806,N_8325,N_9843);
xor U12807 (N_12807,N_9171,N_9046);
or U12808 (N_12808,N_7640,N_8442);
and U12809 (N_12809,N_6189,N_9898);
or U12810 (N_12810,N_7484,N_8118);
nand U12811 (N_12811,N_7629,N_6599);
and U12812 (N_12812,N_5261,N_7430);
xor U12813 (N_12813,N_9491,N_5699);
xnor U12814 (N_12814,N_7965,N_6172);
or U12815 (N_12815,N_8604,N_7051);
and U12816 (N_12816,N_5820,N_6826);
and U12817 (N_12817,N_9910,N_7738);
xnor U12818 (N_12818,N_9691,N_6077);
or U12819 (N_12819,N_5351,N_8601);
and U12820 (N_12820,N_6494,N_6997);
nor U12821 (N_12821,N_9399,N_9055);
xnor U12822 (N_12822,N_7926,N_8144);
and U12823 (N_12823,N_6478,N_8898);
or U12824 (N_12824,N_7343,N_5963);
nor U12825 (N_12825,N_5556,N_9214);
and U12826 (N_12826,N_7164,N_5095);
nand U12827 (N_12827,N_6230,N_5407);
nor U12828 (N_12828,N_8875,N_6887);
xor U12829 (N_12829,N_6326,N_6830);
and U12830 (N_12830,N_9023,N_6305);
xor U12831 (N_12831,N_7480,N_8744);
and U12832 (N_12832,N_5522,N_8216);
nor U12833 (N_12833,N_9285,N_8877);
or U12834 (N_12834,N_5917,N_6586);
nand U12835 (N_12835,N_6885,N_8515);
and U12836 (N_12836,N_6947,N_9384);
nor U12837 (N_12837,N_8289,N_9127);
nor U12838 (N_12838,N_6239,N_7010);
nand U12839 (N_12839,N_6739,N_5473);
nor U12840 (N_12840,N_9285,N_5629);
and U12841 (N_12841,N_9341,N_7105);
or U12842 (N_12842,N_9227,N_9841);
and U12843 (N_12843,N_7268,N_8037);
nor U12844 (N_12844,N_7520,N_5198);
or U12845 (N_12845,N_6929,N_5920);
and U12846 (N_12846,N_9238,N_5218);
or U12847 (N_12847,N_5137,N_9675);
or U12848 (N_12848,N_9169,N_6013);
or U12849 (N_12849,N_8339,N_9961);
xor U12850 (N_12850,N_6822,N_6278);
or U12851 (N_12851,N_9685,N_6715);
and U12852 (N_12852,N_6663,N_7877);
xnor U12853 (N_12853,N_7664,N_8209);
xnor U12854 (N_12854,N_7399,N_5947);
or U12855 (N_12855,N_5821,N_8350);
nor U12856 (N_12856,N_9530,N_5041);
or U12857 (N_12857,N_8409,N_5358);
or U12858 (N_12858,N_7143,N_8519);
nor U12859 (N_12859,N_7618,N_6916);
nand U12860 (N_12860,N_5983,N_6266);
xnor U12861 (N_12861,N_9540,N_5874);
nand U12862 (N_12862,N_9826,N_9315);
and U12863 (N_12863,N_5900,N_9034);
nand U12864 (N_12864,N_7561,N_9304);
xnor U12865 (N_12865,N_9677,N_6749);
or U12866 (N_12866,N_6078,N_8644);
or U12867 (N_12867,N_8346,N_6702);
xor U12868 (N_12868,N_9428,N_8801);
or U12869 (N_12869,N_5477,N_8791);
xor U12870 (N_12870,N_8224,N_8376);
nand U12871 (N_12871,N_9038,N_5559);
or U12872 (N_12872,N_9010,N_7655);
nor U12873 (N_12873,N_8352,N_5225);
nor U12874 (N_12874,N_7467,N_5636);
nor U12875 (N_12875,N_8429,N_9145);
nor U12876 (N_12876,N_5973,N_8509);
or U12877 (N_12877,N_9722,N_7484);
and U12878 (N_12878,N_6980,N_6737);
nand U12879 (N_12879,N_7725,N_6675);
and U12880 (N_12880,N_5811,N_9767);
or U12881 (N_12881,N_9474,N_9682);
xnor U12882 (N_12882,N_9402,N_9595);
or U12883 (N_12883,N_6820,N_9011);
xnor U12884 (N_12884,N_5025,N_7280);
nand U12885 (N_12885,N_7984,N_9648);
and U12886 (N_12886,N_5417,N_7859);
xnor U12887 (N_12887,N_8819,N_9740);
xnor U12888 (N_12888,N_5097,N_6543);
nand U12889 (N_12889,N_6670,N_8461);
and U12890 (N_12890,N_7601,N_5800);
nor U12891 (N_12891,N_6280,N_7143);
and U12892 (N_12892,N_9484,N_7366);
xnor U12893 (N_12893,N_8268,N_9799);
nand U12894 (N_12894,N_5344,N_5240);
nand U12895 (N_12895,N_8089,N_6534);
xor U12896 (N_12896,N_6927,N_6548);
nand U12897 (N_12897,N_8715,N_6203);
nor U12898 (N_12898,N_6239,N_5928);
xnor U12899 (N_12899,N_8593,N_8710);
or U12900 (N_12900,N_6799,N_5190);
or U12901 (N_12901,N_9207,N_7188);
nor U12902 (N_12902,N_9818,N_8204);
xnor U12903 (N_12903,N_7977,N_9301);
nand U12904 (N_12904,N_6367,N_9601);
or U12905 (N_12905,N_8870,N_6809);
and U12906 (N_12906,N_7170,N_5561);
and U12907 (N_12907,N_8720,N_5592);
or U12908 (N_12908,N_7904,N_8147);
nor U12909 (N_12909,N_7065,N_7696);
or U12910 (N_12910,N_8039,N_8635);
and U12911 (N_12911,N_9904,N_8961);
and U12912 (N_12912,N_8459,N_9544);
nand U12913 (N_12913,N_8798,N_5583);
or U12914 (N_12914,N_9796,N_7919);
or U12915 (N_12915,N_8106,N_5518);
xor U12916 (N_12916,N_8139,N_9987);
xor U12917 (N_12917,N_5079,N_7115);
and U12918 (N_12918,N_9073,N_8516);
and U12919 (N_12919,N_8997,N_6341);
nand U12920 (N_12920,N_8634,N_9160);
or U12921 (N_12921,N_8151,N_6056);
nand U12922 (N_12922,N_5166,N_7701);
and U12923 (N_12923,N_6786,N_5274);
nor U12924 (N_12924,N_7779,N_9363);
or U12925 (N_12925,N_8997,N_7133);
and U12926 (N_12926,N_7367,N_5993);
and U12927 (N_12927,N_7653,N_9105);
nor U12928 (N_12928,N_9567,N_6383);
xor U12929 (N_12929,N_6316,N_9541);
nand U12930 (N_12930,N_5172,N_5940);
and U12931 (N_12931,N_9240,N_9092);
xor U12932 (N_12932,N_8678,N_9660);
nand U12933 (N_12933,N_5845,N_5201);
xnor U12934 (N_12934,N_7069,N_5666);
nor U12935 (N_12935,N_9769,N_8144);
nor U12936 (N_12936,N_5385,N_5922);
xnor U12937 (N_12937,N_7078,N_7151);
xnor U12938 (N_12938,N_7583,N_6197);
and U12939 (N_12939,N_9014,N_5566);
nand U12940 (N_12940,N_8996,N_6360);
nand U12941 (N_12941,N_7204,N_9583);
nor U12942 (N_12942,N_7675,N_7224);
xnor U12943 (N_12943,N_8764,N_6252);
or U12944 (N_12944,N_8684,N_5972);
and U12945 (N_12945,N_9621,N_9747);
nor U12946 (N_12946,N_6417,N_7964);
nand U12947 (N_12947,N_9470,N_9010);
nor U12948 (N_12948,N_8041,N_9591);
nand U12949 (N_12949,N_5692,N_5991);
or U12950 (N_12950,N_6237,N_5862);
xnor U12951 (N_12951,N_7445,N_6204);
nand U12952 (N_12952,N_9575,N_7604);
or U12953 (N_12953,N_9194,N_7503);
nand U12954 (N_12954,N_5307,N_5537);
nor U12955 (N_12955,N_6115,N_8309);
and U12956 (N_12956,N_8174,N_9467);
nor U12957 (N_12957,N_7897,N_6312);
nor U12958 (N_12958,N_9429,N_7103);
and U12959 (N_12959,N_7137,N_7374);
nand U12960 (N_12960,N_7368,N_5183);
xor U12961 (N_12961,N_9278,N_7273);
nor U12962 (N_12962,N_9736,N_9969);
and U12963 (N_12963,N_8048,N_7977);
nor U12964 (N_12964,N_5667,N_6294);
xnor U12965 (N_12965,N_8198,N_8966);
or U12966 (N_12966,N_8026,N_5900);
or U12967 (N_12967,N_8960,N_5397);
nand U12968 (N_12968,N_5801,N_9206);
nor U12969 (N_12969,N_9849,N_8893);
xor U12970 (N_12970,N_8087,N_7160);
nand U12971 (N_12971,N_9612,N_5952);
and U12972 (N_12972,N_8991,N_6653);
nand U12973 (N_12973,N_7447,N_6964);
or U12974 (N_12974,N_6810,N_6612);
or U12975 (N_12975,N_5096,N_5012);
and U12976 (N_12976,N_9268,N_8885);
xor U12977 (N_12977,N_7064,N_9689);
xnor U12978 (N_12978,N_6704,N_8269);
or U12979 (N_12979,N_6856,N_7663);
and U12980 (N_12980,N_9538,N_6237);
nand U12981 (N_12981,N_5941,N_5544);
and U12982 (N_12982,N_9550,N_7227);
nand U12983 (N_12983,N_9592,N_7824);
or U12984 (N_12984,N_9481,N_6535);
nor U12985 (N_12985,N_9768,N_8863);
nand U12986 (N_12986,N_7270,N_5886);
or U12987 (N_12987,N_6867,N_7939);
nand U12988 (N_12988,N_8486,N_9451);
xnor U12989 (N_12989,N_6036,N_8217);
or U12990 (N_12990,N_9027,N_7829);
nor U12991 (N_12991,N_8232,N_8451);
nor U12992 (N_12992,N_9744,N_6905);
and U12993 (N_12993,N_9331,N_7679);
xor U12994 (N_12994,N_7301,N_5359);
xor U12995 (N_12995,N_7805,N_7875);
or U12996 (N_12996,N_6960,N_9760);
nand U12997 (N_12997,N_7619,N_6611);
nand U12998 (N_12998,N_9617,N_8029);
nand U12999 (N_12999,N_9044,N_9197);
nor U13000 (N_13000,N_7460,N_7280);
xnor U13001 (N_13001,N_8493,N_5586);
nor U13002 (N_13002,N_9297,N_8389);
nor U13003 (N_13003,N_6212,N_9017);
and U13004 (N_13004,N_8876,N_7514);
or U13005 (N_13005,N_7739,N_8853);
or U13006 (N_13006,N_6220,N_5603);
xnor U13007 (N_13007,N_8551,N_9268);
nor U13008 (N_13008,N_6853,N_7898);
nand U13009 (N_13009,N_9234,N_7316);
nand U13010 (N_13010,N_8232,N_6811);
nor U13011 (N_13011,N_5769,N_7661);
and U13012 (N_13012,N_7880,N_7853);
nor U13013 (N_13013,N_9623,N_6660);
and U13014 (N_13014,N_7867,N_9233);
xor U13015 (N_13015,N_8857,N_7846);
and U13016 (N_13016,N_5239,N_7669);
xor U13017 (N_13017,N_9854,N_5453);
xor U13018 (N_13018,N_6956,N_9779);
and U13019 (N_13019,N_7257,N_5207);
or U13020 (N_13020,N_7666,N_7582);
nor U13021 (N_13021,N_8303,N_8466);
nand U13022 (N_13022,N_5239,N_8374);
and U13023 (N_13023,N_8735,N_6752);
and U13024 (N_13024,N_5785,N_5108);
nand U13025 (N_13025,N_8912,N_8334);
nand U13026 (N_13026,N_8994,N_8399);
xor U13027 (N_13027,N_7506,N_6147);
and U13028 (N_13028,N_6815,N_7141);
xor U13029 (N_13029,N_5219,N_5970);
and U13030 (N_13030,N_5700,N_9178);
xnor U13031 (N_13031,N_7807,N_5469);
xnor U13032 (N_13032,N_9742,N_5181);
or U13033 (N_13033,N_9923,N_8522);
nor U13034 (N_13034,N_6933,N_6936);
nor U13035 (N_13035,N_7207,N_6338);
nor U13036 (N_13036,N_7285,N_7872);
nand U13037 (N_13037,N_9433,N_8974);
and U13038 (N_13038,N_6700,N_6893);
nand U13039 (N_13039,N_8179,N_8809);
nor U13040 (N_13040,N_8651,N_7400);
nand U13041 (N_13041,N_5968,N_8110);
or U13042 (N_13042,N_8459,N_9579);
or U13043 (N_13043,N_6401,N_6183);
or U13044 (N_13044,N_6412,N_5021);
xnor U13045 (N_13045,N_7703,N_7968);
and U13046 (N_13046,N_8332,N_8547);
nor U13047 (N_13047,N_8583,N_7046);
and U13048 (N_13048,N_6393,N_7832);
or U13049 (N_13049,N_5424,N_6561);
nor U13050 (N_13050,N_8460,N_7606);
or U13051 (N_13051,N_9628,N_8782);
nor U13052 (N_13052,N_7354,N_8132);
or U13053 (N_13053,N_6737,N_5846);
and U13054 (N_13054,N_7810,N_5441);
xnor U13055 (N_13055,N_5712,N_6897);
nor U13056 (N_13056,N_5635,N_9208);
and U13057 (N_13057,N_9449,N_6151);
nand U13058 (N_13058,N_7399,N_8757);
and U13059 (N_13059,N_6164,N_7398);
nand U13060 (N_13060,N_7859,N_9338);
nand U13061 (N_13061,N_5826,N_9945);
xor U13062 (N_13062,N_9033,N_7820);
nand U13063 (N_13063,N_9279,N_6851);
xor U13064 (N_13064,N_8581,N_7343);
nor U13065 (N_13065,N_9851,N_8632);
nand U13066 (N_13066,N_5779,N_8975);
nor U13067 (N_13067,N_6461,N_5537);
nand U13068 (N_13068,N_9247,N_8564);
nand U13069 (N_13069,N_8424,N_5832);
and U13070 (N_13070,N_8745,N_7712);
or U13071 (N_13071,N_6458,N_5924);
and U13072 (N_13072,N_5067,N_6314);
or U13073 (N_13073,N_8125,N_5805);
xnor U13074 (N_13074,N_7396,N_8771);
or U13075 (N_13075,N_8086,N_9648);
and U13076 (N_13076,N_6633,N_5040);
or U13077 (N_13077,N_8353,N_7970);
or U13078 (N_13078,N_5930,N_6404);
or U13079 (N_13079,N_5979,N_5506);
xor U13080 (N_13080,N_8899,N_5313);
nand U13081 (N_13081,N_5864,N_9153);
and U13082 (N_13082,N_7824,N_6893);
and U13083 (N_13083,N_6233,N_9190);
nand U13084 (N_13084,N_8429,N_5980);
nor U13085 (N_13085,N_5395,N_7322);
and U13086 (N_13086,N_5124,N_6654);
and U13087 (N_13087,N_5968,N_8866);
or U13088 (N_13088,N_5084,N_5522);
xnor U13089 (N_13089,N_5186,N_7223);
nor U13090 (N_13090,N_8420,N_6978);
or U13091 (N_13091,N_9743,N_5855);
and U13092 (N_13092,N_6464,N_5301);
or U13093 (N_13093,N_6317,N_6585);
and U13094 (N_13094,N_5062,N_6938);
nor U13095 (N_13095,N_5380,N_6709);
and U13096 (N_13096,N_9671,N_8746);
xor U13097 (N_13097,N_7573,N_8282);
xnor U13098 (N_13098,N_7827,N_6396);
and U13099 (N_13099,N_9738,N_9315);
nor U13100 (N_13100,N_9111,N_5094);
nand U13101 (N_13101,N_7106,N_9919);
nand U13102 (N_13102,N_8893,N_7103);
xnor U13103 (N_13103,N_6528,N_7362);
or U13104 (N_13104,N_6739,N_5903);
xor U13105 (N_13105,N_9639,N_6642);
nand U13106 (N_13106,N_5775,N_7443);
xor U13107 (N_13107,N_6587,N_8736);
nand U13108 (N_13108,N_5522,N_8169);
nand U13109 (N_13109,N_9343,N_8344);
nor U13110 (N_13110,N_9019,N_9756);
and U13111 (N_13111,N_5964,N_6375);
xnor U13112 (N_13112,N_8668,N_8938);
and U13113 (N_13113,N_7416,N_8734);
xor U13114 (N_13114,N_8225,N_5968);
nor U13115 (N_13115,N_6882,N_5805);
nor U13116 (N_13116,N_7090,N_6961);
nor U13117 (N_13117,N_5401,N_9350);
xnor U13118 (N_13118,N_6992,N_7640);
and U13119 (N_13119,N_8352,N_7623);
and U13120 (N_13120,N_5345,N_8744);
nor U13121 (N_13121,N_7946,N_9486);
nand U13122 (N_13122,N_7202,N_6931);
nand U13123 (N_13123,N_7572,N_5714);
nand U13124 (N_13124,N_9562,N_6926);
nand U13125 (N_13125,N_7074,N_8782);
nand U13126 (N_13126,N_5445,N_6177);
xor U13127 (N_13127,N_5745,N_8068);
and U13128 (N_13128,N_5306,N_5365);
nor U13129 (N_13129,N_7575,N_5636);
and U13130 (N_13130,N_8932,N_5683);
or U13131 (N_13131,N_8403,N_5321);
xor U13132 (N_13132,N_7831,N_6216);
and U13133 (N_13133,N_8194,N_5793);
nand U13134 (N_13134,N_5620,N_9023);
and U13135 (N_13135,N_5541,N_5916);
xor U13136 (N_13136,N_6184,N_8040);
nor U13137 (N_13137,N_9187,N_7642);
and U13138 (N_13138,N_7426,N_6015);
xor U13139 (N_13139,N_9558,N_8719);
and U13140 (N_13140,N_6008,N_8127);
or U13141 (N_13141,N_6444,N_5186);
nor U13142 (N_13142,N_7236,N_7029);
and U13143 (N_13143,N_5388,N_7892);
and U13144 (N_13144,N_7040,N_7501);
xor U13145 (N_13145,N_8276,N_5770);
nand U13146 (N_13146,N_8087,N_9523);
and U13147 (N_13147,N_8821,N_5041);
xor U13148 (N_13148,N_9608,N_7078);
or U13149 (N_13149,N_8304,N_7561);
nand U13150 (N_13150,N_7197,N_9944);
xnor U13151 (N_13151,N_6925,N_5796);
nand U13152 (N_13152,N_7729,N_9688);
or U13153 (N_13153,N_9420,N_5501);
and U13154 (N_13154,N_5693,N_5836);
or U13155 (N_13155,N_5195,N_8693);
nand U13156 (N_13156,N_7666,N_6522);
xnor U13157 (N_13157,N_9655,N_9377);
nor U13158 (N_13158,N_5243,N_8365);
and U13159 (N_13159,N_6205,N_8202);
nor U13160 (N_13160,N_6853,N_6419);
xor U13161 (N_13161,N_6840,N_6127);
and U13162 (N_13162,N_9700,N_5083);
xor U13163 (N_13163,N_6977,N_5524);
and U13164 (N_13164,N_6071,N_9836);
nor U13165 (N_13165,N_8519,N_9211);
nor U13166 (N_13166,N_5114,N_6174);
and U13167 (N_13167,N_8334,N_8154);
and U13168 (N_13168,N_5124,N_7791);
and U13169 (N_13169,N_8258,N_6919);
and U13170 (N_13170,N_9306,N_8673);
or U13171 (N_13171,N_9591,N_8028);
or U13172 (N_13172,N_7024,N_7819);
nor U13173 (N_13173,N_8214,N_5564);
and U13174 (N_13174,N_6704,N_9207);
xnor U13175 (N_13175,N_9879,N_5713);
nor U13176 (N_13176,N_9527,N_8743);
and U13177 (N_13177,N_7198,N_8944);
xor U13178 (N_13178,N_7479,N_5644);
or U13179 (N_13179,N_6067,N_8109);
xnor U13180 (N_13180,N_5343,N_8129);
nand U13181 (N_13181,N_8760,N_6097);
xnor U13182 (N_13182,N_5471,N_8717);
nor U13183 (N_13183,N_8973,N_8877);
nand U13184 (N_13184,N_6148,N_8944);
nand U13185 (N_13185,N_8059,N_5593);
nand U13186 (N_13186,N_5414,N_6491);
nand U13187 (N_13187,N_9772,N_9086);
nand U13188 (N_13188,N_7727,N_7212);
xor U13189 (N_13189,N_6790,N_6754);
nand U13190 (N_13190,N_9895,N_9807);
and U13191 (N_13191,N_5329,N_5679);
and U13192 (N_13192,N_8049,N_6937);
and U13193 (N_13193,N_9211,N_8297);
nor U13194 (N_13194,N_9620,N_8925);
xor U13195 (N_13195,N_6487,N_6608);
nand U13196 (N_13196,N_8566,N_6413);
nor U13197 (N_13197,N_8225,N_6052);
nand U13198 (N_13198,N_8419,N_6124);
xor U13199 (N_13199,N_9610,N_5034);
or U13200 (N_13200,N_6697,N_9336);
or U13201 (N_13201,N_6048,N_6411);
nand U13202 (N_13202,N_8870,N_9572);
nor U13203 (N_13203,N_7086,N_9084);
or U13204 (N_13204,N_9131,N_6390);
and U13205 (N_13205,N_5312,N_7496);
xor U13206 (N_13206,N_5862,N_8312);
nor U13207 (N_13207,N_8417,N_6727);
nand U13208 (N_13208,N_5120,N_7950);
xnor U13209 (N_13209,N_6209,N_7375);
xor U13210 (N_13210,N_8538,N_8808);
and U13211 (N_13211,N_5940,N_7938);
nand U13212 (N_13212,N_6906,N_9739);
nand U13213 (N_13213,N_7356,N_8516);
or U13214 (N_13214,N_7894,N_5000);
nor U13215 (N_13215,N_5930,N_9238);
xnor U13216 (N_13216,N_9045,N_7097);
or U13217 (N_13217,N_7702,N_5068);
nand U13218 (N_13218,N_7428,N_6400);
and U13219 (N_13219,N_8022,N_9463);
or U13220 (N_13220,N_6751,N_7970);
xor U13221 (N_13221,N_6650,N_9335);
nand U13222 (N_13222,N_5097,N_5145);
xor U13223 (N_13223,N_9540,N_5571);
nand U13224 (N_13224,N_6213,N_9830);
xor U13225 (N_13225,N_8882,N_8650);
nand U13226 (N_13226,N_7491,N_5530);
or U13227 (N_13227,N_7395,N_9845);
and U13228 (N_13228,N_7309,N_9905);
or U13229 (N_13229,N_8368,N_7366);
xor U13230 (N_13230,N_9090,N_5559);
xor U13231 (N_13231,N_5968,N_5459);
nand U13232 (N_13232,N_9970,N_5284);
nand U13233 (N_13233,N_8218,N_5856);
nand U13234 (N_13234,N_6897,N_5901);
nor U13235 (N_13235,N_6969,N_8748);
and U13236 (N_13236,N_5014,N_8102);
nor U13237 (N_13237,N_7385,N_6619);
and U13238 (N_13238,N_5144,N_5060);
or U13239 (N_13239,N_8139,N_6877);
and U13240 (N_13240,N_5432,N_8155);
or U13241 (N_13241,N_8980,N_7307);
and U13242 (N_13242,N_6495,N_5931);
xnor U13243 (N_13243,N_6410,N_8503);
and U13244 (N_13244,N_9265,N_9021);
and U13245 (N_13245,N_6811,N_5738);
nand U13246 (N_13246,N_9078,N_6243);
nand U13247 (N_13247,N_5285,N_6730);
xnor U13248 (N_13248,N_6638,N_6542);
and U13249 (N_13249,N_6715,N_6268);
nor U13250 (N_13250,N_9871,N_9626);
and U13251 (N_13251,N_6281,N_7252);
nor U13252 (N_13252,N_6476,N_9678);
nand U13253 (N_13253,N_6864,N_8929);
nand U13254 (N_13254,N_6570,N_5472);
nand U13255 (N_13255,N_6570,N_6984);
nor U13256 (N_13256,N_6783,N_6746);
or U13257 (N_13257,N_5888,N_8910);
xnor U13258 (N_13258,N_5318,N_9131);
nor U13259 (N_13259,N_8914,N_5480);
or U13260 (N_13260,N_8899,N_8672);
nor U13261 (N_13261,N_5740,N_5164);
nor U13262 (N_13262,N_9788,N_7207);
xnor U13263 (N_13263,N_6187,N_8359);
or U13264 (N_13264,N_6748,N_5023);
and U13265 (N_13265,N_8864,N_7434);
xnor U13266 (N_13266,N_8447,N_9533);
xnor U13267 (N_13267,N_7012,N_8917);
nand U13268 (N_13268,N_6614,N_6702);
or U13269 (N_13269,N_9687,N_8702);
nand U13270 (N_13270,N_7325,N_7107);
or U13271 (N_13271,N_9466,N_8509);
nor U13272 (N_13272,N_7056,N_7166);
xor U13273 (N_13273,N_5609,N_6705);
nor U13274 (N_13274,N_5489,N_6295);
or U13275 (N_13275,N_9068,N_7595);
xor U13276 (N_13276,N_5659,N_7042);
or U13277 (N_13277,N_9114,N_8522);
nand U13278 (N_13278,N_5964,N_8190);
nand U13279 (N_13279,N_5000,N_5029);
nand U13280 (N_13280,N_6463,N_9648);
xnor U13281 (N_13281,N_7406,N_8296);
and U13282 (N_13282,N_5916,N_9383);
xor U13283 (N_13283,N_6991,N_6134);
nand U13284 (N_13284,N_5642,N_5596);
or U13285 (N_13285,N_7684,N_6823);
nand U13286 (N_13286,N_9488,N_6989);
nor U13287 (N_13287,N_5956,N_6166);
or U13288 (N_13288,N_7897,N_9691);
nand U13289 (N_13289,N_9240,N_9421);
or U13290 (N_13290,N_6294,N_7767);
or U13291 (N_13291,N_5430,N_5708);
nor U13292 (N_13292,N_9207,N_8726);
nand U13293 (N_13293,N_7436,N_9808);
nor U13294 (N_13294,N_6587,N_9088);
and U13295 (N_13295,N_7627,N_5286);
nand U13296 (N_13296,N_7014,N_5007);
or U13297 (N_13297,N_9996,N_7322);
nand U13298 (N_13298,N_7451,N_9646);
nor U13299 (N_13299,N_9864,N_7796);
nor U13300 (N_13300,N_5722,N_7229);
nor U13301 (N_13301,N_9700,N_9181);
nor U13302 (N_13302,N_5352,N_5190);
nand U13303 (N_13303,N_7609,N_7278);
and U13304 (N_13304,N_6218,N_9283);
nand U13305 (N_13305,N_7121,N_7539);
nor U13306 (N_13306,N_8883,N_9171);
xor U13307 (N_13307,N_6370,N_8999);
xnor U13308 (N_13308,N_9673,N_9016);
nor U13309 (N_13309,N_9260,N_5053);
xor U13310 (N_13310,N_5857,N_6587);
nand U13311 (N_13311,N_5501,N_9513);
nor U13312 (N_13312,N_5966,N_7282);
nand U13313 (N_13313,N_9374,N_7067);
and U13314 (N_13314,N_5863,N_5257);
nor U13315 (N_13315,N_6620,N_6979);
xor U13316 (N_13316,N_5736,N_7177);
xor U13317 (N_13317,N_6337,N_7664);
nor U13318 (N_13318,N_7460,N_6855);
nand U13319 (N_13319,N_7210,N_5276);
nand U13320 (N_13320,N_5284,N_7881);
nand U13321 (N_13321,N_8561,N_6630);
and U13322 (N_13322,N_9753,N_7057);
xnor U13323 (N_13323,N_5352,N_6684);
nand U13324 (N_13324,N_9456,N_8094);
nor U13325 (N_13325,N_8964,N_5889);
nor U13326 (N_13326,N_7617,N_9573);
nand U13327 (N_13327,N_6294,N_6487);
nor U13328 (N_13328,N_9785,N_5684);
nand U13329 (N_13329,N_7218,N_7105);
nor U13330 (N_13330,N_8085,N_8315);
or U13331 (N_13331,N_9660,N_7024);
xnor U13332 (N_13332,N_6989,N_9016);
xor U13333 (N_13333,N_5491,N_5229);
nand U13334 (N_13334,N_8907,N_9743);
xor U13335 (N_13335,N_9190,N_5943);
xor U13336 (N_13336,N_6521,N_9505);
or U13337 (N_13337,N_6114,N_9867);
and U13338 (N_13338,N_7612,N_9116);
nor U13339 (N_13339,N_5573,N_7917);
nor U13340 (N_13340,N_7610,N_7965);
nor U13341 (N_13341,N_5413,N_5333);
xnor U13342 (N_13342,N_9980,N_5157);
or U13343 (N_13343,N_9467,N_9587);
nand U13344 (N_13344,N_5321,N_9545);
and U13345 (N_13345,N_9143,N_8524);
or U13346 (N_13346,N_7081,N_9621);
or U13347 (N_13347,N_5119,N_7763);
nor U13348 (N_13348,N_5240,N_7220);
or U13349 (N_13349,N_9073,N_5384);
xnor U13350 (N_13350,N_6172,N_9366);
or U13351 (N_13351,N_9347,N_7356);
and U13352 (N_13352,N_7497,N_5387);
nand U13353 (N_13353,N_6877,N_6204);
xnor U13354 (N_13354,N_5963,N_7643);
nor U13355 (N_13355,N_8868,N_8189);
and U13356 (N_13356,N_9228,N_7644);
nand U13357 (N_13357,N_7366,N_8572);
nor U13358 (N_13358,N_8705,N_6726);
nand U13359 (N_13359,N_9661,N_5345);
nor U13360 (N_13360,N_5690,N_6247);
and U13361 (N_13361,N_9535,N_6672);
nor U13362 (N_13362,N_7346,N_9611);
nand U13363 (N_13363,N_9245,N_8708);
and U13364 (N_13364,N_9386,N_8670);
or U13365 (N_13365,N_7202,N_6868);
nand U13366 (N_13366,N_8284,N_7733);
nor U13367 (N_13367,N_7247,N_7025);
or U13368 (N_13368,N_9723,N_6344);
xnor U13369 (N_13369,N_7060,N_5568);
and U13370 (N_13370,N_8026,N_8210);
and U13371 (N_13371,N_8397,N_7877);
xor U13372 (N_13372,N_8199,N_6522);
xnor U13373 (N_13373,N_7589,N_7072);
xor U13374 (N_13374,N_5503,N_6423);
nand U13375 (N_13375,N_8238,N_8603);
and U13376 (N_13376,N_5200,N_6171);
and U13377 (N_13377,N_7770,N_8516);
xor U13378 (N_13378,N_6731,N_5261);
and U13379 (N_13379,N_5015,N_5093);
nand U13380 (N_13380,N_9797,N_9648);
nand U13381 (N_13381,N_5985,N_5952);
nor U13382 (N_13382,N_7032,N_9812);
nor U13383 (N_13383,N_5176,N_8377);
nand U13384 (N_13384,N_9940,N_8887);
nor U13385 (N_13385,N_7973,N_9960);
and U13386 (N_13386,N_7452,N_7077);
nand U13387 (N_13387,N_9660,N_9342);
nor U13388 (N_13388,N_8745,N_9229);
or U13389 (N_13389,N_6325,N_7073);
nor U13390 (N_13390,N_5807,N_7519);
or U13391 (N_13391,N_6197,N_6105);
or U13392 (N_13392,N_8037,N_7185);
and U13393 (N_13393,N_7951,N_5939);
nor U13394 (N_13394,N_8894,N_9271);
nor U13395 (N_13395,N_8352,N_6925);
nor U13396 (N_13396,N_5780,N_7478);
nor U13397 (N_13397,N_6598,N_6003);
nand U13398 (N_13398,N_8136,N_7378);
and U13399 (N_13399,N_6050,N_6446);
and U13400 (N_13400,N_7567,N_5995);
and U13401 (N_13401,N_6169,N_7099);
nor U13402 (N_13402,N_8373,N_8174);
and U13403 (N_13403,N_7648,N_8169);
or U13404 (N_13404,N_6485,N_6207);
nor U13405 (N_13405,N_7506,N_9450);
xnor U13406 (N_13406,N_7637,N_7492);
and U13407 (N_13407,N_6709,N_5983);
nand U13408 (N_13408,N_9138,N_9062);
and U13409 (N_13409,N_7339,N_6871);
xnor U13410 (N_13410,N_8578,N_5685);
and U13411 (N_13411,N_9438,N_7508);
xnor U13412 (N_13412,N_8015,N_7074);
or U13413 (N_13413,N_7759,N_9322);
nor U13414 (N_13414,N_6674,N_7295);
or U13415 (N_13415,N_9722,N_5738);
nor U13416 (N_13416,N_6205,N_5349);
or U13417 (N_13417,N_5031,N_6709);
nand U13418 (N_13418,N_8034,N_8172);
nor U13419 (N_13419,N_9703,N_6829);
nand U13420 (N_13420,N_8094,N_8621);
or U13421 (N_13421,N_9432,N_5460);
or U13422 (N_13422,N_8213,N_8911);
nand U13423 (N_13423,N_5597,N_7086);
xnor U13424 (N_13424,N_9603,N_6809);
nor U13425 (N_13425,N_7984,N_6882);
xnor U13426 (N_13426,N_6697,N_6778);
or U13427 (N_13427,N_6983,N_6196);
xor U13428 (N_13428,N_8476,N_7747);
or U13429 (N_13429,N_6657,N_9787);
or U13430 (N_13430,N_7539,N_7207);
or U13431 (N_13431,N_5256,N_6245);
or U13432 (N_13432,N_9095,N_9584);
or U13433 (N_13433,N_8931,N_8924);
or U13434 (N_13434,N_6506,N_5123);
nor U13435 (N_13435,N_8790,N_8992);
nor U13436 (N_13436,N_7114,N_9851);
and U13437 (N_13437,N_9740,N_7982);
xnor U13438 (N_13438,N_8481,N_8624);
nand U13439 (N_13439,N_6981,N_9569);
nand U13440 (N_13440,N_7358,N_7940);
and U13441 (N_13441,N_9916,N_6767);
and U13442 (N_13442,N_6908,N_7879);
nor U13443 (N_13443,N_8313,N_5957);
xor U13444 (N_13444,N_5851,N_8288);
or U13445 (N_13445,N_9332,N_9154);
xor U13446 (N_13446,N_8233,N_7038);
nand U13447 (N_13447,N_7821,N_7455);
or U13448 (N_13448,N_6998,N_6217);
xor U13449 (N_13449,N_5801,N_6068);
nor U13450 (N_13450,N_7800,N_7720);
or U13451 (N_13451,N_6443,N_5928);
and U13452 (N_13452,N_9423,N_7820);
nand U13453 (N_13453,N_7860,N_5319);
nand U13454 (N_13454,N_8480,N_6153);
nor U13455 (N_13455,N_7974,N_5165);
xnor U13456 (N_13456,N_5470,N_7024);
xor U13457 (N_13457,N_5849,N_7596);
xnor U13458 (N_13458,N_6795,N_7932);
and U13459 (N_13459,N_8950,N_6586);
or U13460 (N_13460,N_8476,N_8281);
nand U13461 (N_13461,N_5148,N_7832);
nor U13462 (N_13462,N_8455,N_9887);
xor U13463 (N_13463,N_5602,N_5128);
nand U13464 (N_13464,N_8129,N_6971);
xnor U13465 (N_13465,N_9934,N_8992);
and U13466 (N_13466,N_9119,N_6561);
xor U13467 (N_13467,N_9906,N_8420);
nor U13468 (N_13468,N_6586,N_8944);
xor U13469 (N_13469,N_9839,N_5386);
or U13470 (N_13470,N_8558,N_8683);
and U13471 (N_13471,N_8948,N_7822);
nand U13472 (N_13472,N_7853,N_8266);
and U13473 (N_13473,N_7344,N_8986);
xor U13474 (N_13474,N_6747,N_7425);
nand U13475 (N_13475,N_8405,N_9334);
xnor U13476 (N_13476,N_9011,N_8014);
nor U13477 (N_13477,N_6316,N_5152);
nor U13478 (N_13478,N_7492,N_7163);
and U13479 (N_13479,N_5508,N_6125);
and U13480 (N_13480,N_5372,N_6486);
xnor U13481 (N_13481,N_6973,N_5395);
nand U13482 (N_13482,N_7869,N_9588);
and U13483 (N_13483,N_9182,N_9026);
or U13484 (N_13484,N_9244,N_9316);
or U13485 (N_13485,N_8788,N_9240);
xor U13486 (N_13486,N_7179,N_6014);
and U13487 (N_13487,N_5986,N_7411);
nor U13488 (N_13488,N_5290,N_5030);
xor U13489 (N_13489,N_5237,N_8509);
nor U13490 (N_13490,N_6630,N_9742);
and U13491 (N_13491,N_5049,N_8943);
or U13492 (N_13492,N_7612,N_7795);
nor U13493 (N_13493,N_6748,N_9843);
nand U13494 (N_13494,N_6255,N_5530);
nand U13495 (N_13495,N_9401,N_5704);
nor U13496 (N_13496,N_8087,N_9514);
and U13497 (N_13497,N_6231,N_6099);
xnor U13498 (N_13498,N_8339,N_9137);
nand U13499 (N_13499,N_5511,N_5566);
nand U13500 (N_13500,N_6976,N_6736);
xnor U13501 (N_13501,N_8570,N_8484);
nand U13502 (N_13502,N_7871,N_9784);
xnor U13503 (N_13503,N_5029,N_6738);
nand U13504 (N_13504,N_5999,N_5881);
or U13505 (N_13505,N_7313,N_7347);
and U13506 (N_13506,N_6821,N_8612);
or U13507 (N_13507,N_9314,N_7490);
nor U13508 (N_13508,N_5006,N_5361);
nor U13509 (N_13509,N_9150,N_8605);
xor U13510 (N_13510,N_6868,N_9848);
and U13511 (N_13511,N_8872,N_7692);
nand U13512 (N_13512,N_5525,N_6865);
nor U13513 (N_13513,N_7829,N_9331);
or U13514 (N_13514,N_9788,N_7295);
or U13515 (N_13515,N_7425,N_8538);
nand U13516 (N_13516,N_6706,N_7382);
nor U13517 (N_13517,N_6443,N_8551);
xnor U13518 (N_13518,N_7536,N_5595);
or U13519 (N_13519,N_7798,N_7229);
xor U13520 (N_13520,N_6832,N_9258);
nor U13521 (N_13521,N_7174,N_9548);
or U13522 (N_13522,N_6013,N_6152);
or U13523 (N_13523,N_9770,N_9958);
nand U13524 (N_13524,N_6839,N_7056);
nor U13525 (N_13525,N_7387,N_8655);
xnor U13526 (N_13526,N_9797,N_8796);
and U13527 (N_13527,N_6617,N_5261);
or U13528 (N_13528,N_8783,N_8269);
nor U13529 (N_13529,N_7472,N_5496);
or U13530 (N_13530,N_9409,N_9178);
and U13531 (N_13531,N_7201,N_6080);
nand U13532 (N_13532,N_6665,N_7211);
or U13533 (N_13533,N_8813,N_5727);
nor U13534 (N_13534,N_7169,N_7138);
and U13535 (N_13535,N_8711,N_8291);
nor U13536 (N_13536,N_6713,N_5674);
and U13537 (N_13537,N_8590,N_6608);
nand U13538 (N_13538,N_9508,N_8271);
xor U13539 (N_13539,N_9052,N_7388);
and U13540 (N_13540,N_7043,N_8324);
and U13541 (N_13541,N_9264,N_9826);
xor U13542 (N_13542,N_5639,N_5701);
and U13543 (N_13543,N_5825,N_6359);
or U13544 (N_13544,N_9259,N_6752);
nand U13545 (N_13545,N_5076,N_5026);
or U13546 (N_13546,N_7286,N_8687);
xor U13547 (N_13547,N_8438,N_5933);
xor U13548 (N_13548,N_8650,N_7514);
xnor U13549 (N_13549,N_5554,N_8542);
nand U13550 (N_13550,N_5181,N_6912);
nand U13551 (N_13551,N_8120,N_9400);
or U13552 (N_13552,N_7195,N_5596);
or U13553 (N_13553,N_7669,N_9120);
and U13554 (N_13554,N_6106,N_5506);
and U13555 (N_13555,N_6529,N_5905);
and U13556 (N_13556,N_6100,N_9013);
xnor U13557 (N_13557,N_7152,N_8124);
nor U13558 (N_13558,N_9618,N_8074);
nor U13559 (N_13559,N_9278,N_7383);
and U13560 (N_13560,N_5299,N_9337);
or U13561 (N_13561,N_7145,N_8903);
or U13562 (N_13562,N_5229,N_8788);
nor U13563 (N_13563,N_8220,N_9762);
nand U13564 (N_13564,N_9495,N_5734);
nor U13565 (N_13565,N_8480,N_5641);
xnor U13566 (N_13566,N_6242,N_7173);
nor U13567 (N_13567,N_9645,N_7686);
or U13568 (N_13568,N_8399,N_9311);
xnor U13569 (N_13569,N_5846,N_9695);
or U13570 (N_13570,N_5063,N_7720);
nor U13571 (N_13571,N_9309,N_9233);
and U13572 (N_13572,N_8825,N_7181);
nor U13573 (N_13573,N_8241,N_8023);
xor U13574 (N_13574,N_5960,N_7942);
xnor U13575 (N_13575,N_8156,N_7624);
nand U13576 (N_13576,N_5003,N_9082);
or U13577 (N_13577,N_6131,N_6805);
nand U13578 (N_13578,N_8986,N_7285);
nor U13579 (N_13579,N_6185,N_5380);
or U13580 (N_13580,N_9797,N_8353);
nor U13581 (N_13581,N_7505,N_5642);
and U13582 (N_13582,N_7550,N_8342);
or U13583 (N_13583,N_7727,N_8457);
xnor U13584 (N_13584,N_8251,N_5401);
and U13585 (N_13585,N_8957,N_6485);
nand U13586 (N_13586,N_5959,N_5261);
nand U13587 (N_13587,N_6861,N_6264);
nor U13588 (N_13588,N_8348,N_9326);
xor U13589 (N_13589,N_6879,N_6318);
and U13590 (N_13590,N_5135,N_5497);
or U13591 (N_13591,N_9871,N_7598);
and U13592 (N_13592,N_7770,N_6769);
and U13593 (N_13593,N_6476,N_7735);
xnor U13594 (N_13594,N_8811,N_5200);
xor U13595 (N_13595,N_9162,N_8854);
nand U13596 (N_13596,N_6458,N_8242);
xnor U13597 (N_13597,N_6368,N_6810);
nor U13598 (N_13598,N_6009,N_6720);
or U13599 (N_13599,N_7166,N_8443);
nor U13600 (N_13600,N_9682,N_5741);
and U13601 (N_13601,N_6814,N_8557);
xor U13602 (N_13602,N_8846,N_8790);
or U13603 (N_13603,N_6698,N_7301);
xor U13604 (N_13604,N_7847,N_5176);
and U13605 (N_13605,N_7353,N_7099);
nand U13606 (N_13606,N_8369,N_5140);
nand U13607 (N_13607,N_7112,N_5234);
xnor U13608 (N_13608,N_5166,N_6520);
and U13609 (N_13609,N_5351,N_7171);
nand U13610 (N_13610,N_5876,N_8154);
xor U13611 (N_13611,N_8724,N_7732);
nand U13612 (N_13612,N_7796,N_7078);
or U13613 (N_13613,N_7637,N_5279);
xor U13614 (N_13614,N_7228,N_7608);
nand U13615 (N_13615,N_6957,N_9760);
nor U13616 (N_13616,N_9809,N_7974);
or U13617 (N_13617,N_9042,N_7748);
nor U13618 (N_13618,N_8040,N_8008);
xnor U13619 (N_13619,N_7000,N_7064);
nand U13620 (N_13620,N_7529,N_7633);
nand U13621 (N_13621,N_7683,N_5863);
xor U13622 (N_13622,N_9994,N_9725);
xor U13623 (N_13623,N_7706,N_9634);
nor U13624 (N_13624,N_5663,N_7398);
nand U13625 (N_13625,N_6396,N_6442);
xor U13626 (N_13626,N_6270,N_8470);
and U13627 (N_13627,N_8157,N_5754);
nor U13628 (N_13628,N_8234,N_6519);
nand U13629 (N_13629,N_5842,N_6770);
nor U13630 (N_13630,N_7456,N_8041);
nand U13631 (N_13631,N_9482,N_9457);
xnor U13632 (N_13632,N_5303,N_5437);
xor U13633 (N_13633,N_8676,N_5191);
or U13634 (N_13634,N_6820,N_5522);
and U13635 (N_13635,N_5825,N_9039);
and U13636 (N_13636,N_5781,N_8540);
and U13637 (N_13637,N_9711,N_8410);
or U13638 (N_13638,N_6115,N_5098);
nor U13639 (N_13639,N_8653,N_9353);
nor U13640 (N_13640,N_6584,N_7626);
nand U13641 (N_13641,N_8507,N_6930);
and U13642 (N_13642,N_8593,N_5395);
nor U13643 (N_13643,N_8242,N_9258);
or U13644 (N_13644,N_5957,N_8361);
nand U13645 (N_13645,N_6011,N_7632);
nand U13646 (N_13646,N_7389,N_7767);
and U13647 (N_13647,N_7461,N_6643);
xnor U13648 (N_13648,N_9256,N_9763);
nand U13649 (N_13649,N_7115,N_6717);
nand U13650 (N_13650,N_8264,N_9464);
xnor U13651 (N_13651,N_7082,N_6482);
nand U13652 (N_13652,N_7673,N_5230);
and U13653 (N_13653,N_6083,N_8842);
nand U13654 (N_13654,N_9256,N_6247);
xor U13655 (N_13655,N_9043,N_8888);
nor U13656 (N_13656,N_7114,N_6122);
xnor U13657 (N_13657,N_9502,N_9716);
and U13658 (N_13658,N_7061,N_5478);
or U13659 (N_13659,N_6889,N_7963);
nor U13660 (N_13660,N_6662,N_5258);
xor U13661 (N_13661,N_7098,N_7050);
and U13662 (N_13662,N_5166,N_7485);
and U13663 (N_13663,N_9380,N_7494);
nor U13664 (N_13664,N_8347,N_8262);
xor U13665 (N_13665,N_6836,N_8965);
nor U13666 (N_13666,N_9592,N_8960);
and U13667 (N_13667,N_7019,N_5673);
nand U13668 (N_13668,N_9700,N_5676);
xor U13669 (N_13669,N_9421,N_8987);
nor U13670 (N_13670,N_6421,N_9276);
nor U13671 (N_13671,N_7505,N_8129);
xnor U13672 (N_13672,N_8845,N_8112);
xnor U13673 (N_13673,N_9980,N_8470);
or U13674 (N_13674,N_5371,N_5246);
nor U13675 (N_13675,N_5219,N_6493);
and U13676 (N_13676,N_5788,N_5432);
xor U13677 (N_13677,N_9898,N_6571);
or U13678 (N_13678,N_8096,N_7893);
xnor U13679 (N_13679,N_7402,N_5400);
nor U13680 (N_13680,N_7934,N_8284);
or U13681 (N_13681,N_7658,N_9932);
and U13682 (N_13682,N_6701,N_6895);
nor U13683 (N_13683,N_7886,N_6571);
and U13684 (N_13684,N_8648,N_7221);
nor U13685 (N_13685,N_7575,N_7672);
xor U13686 (N_13686,N_8835,N_6055);
and U13687 (N_13687,N_7310,N_9783);
or U13688 (N_13688,N_8943,N_6514);
or U13689 (N_13689,N_5514,N_6868);
xnor U13690 (N_13690,N_9001,N_9662);
nand U13691 (N_13691,N_5924,N_9285);
or U13692 (N_13692,N_8526,N_5708);
or U13693 (N_13693,N_9482,N_7495);
nand U13694 (N_13694,N_5628,N_8174);
nor U13695 (N_13695,N_8624,N_9417);
nor U13696 (N_13696,N_7203,N_8643);
nand U13697 (N_13697,N_9871,N_5307);
nand U13698 (N_13698,N_6461,N_7922);
and U13699 (N_13699,N_7873,N_9170);
or U13700 (N_13700,N_5606,N_6343);
and U13701 (N_13701,N_7952,N_9191);
and U13702 (N_13702,N_6884,N_7655);
xor U13703 (N_13703,N_6851,N_5909);
or U13704 (N_13704,N_8281,N_7628);
nand U13705 (N_13705,N_8463,N_8481);
xnor U13706 (N_13706,N_8750,N_8330);
and U13707 (N_13707,N_7284,N_8304);
or U13708 (N_13708,N_6139,N_8305);
or U13709 (N_13709,N_9717,N_6609);
nor U13710 (N_13710,N_9252,N_6110);
xor U13711 (N_13711,N_6705,N_5884);
xor U13712 (N_13712,N_5699,N_8617);
xor U13713 (N_13713,N_5739,N_7190);
nand U13714 (N_13714,N_9301,N_7410);
nand U13715 (N_13715,N_9704,N_7256);
nor U13716 (N_13716,N_7397,N_5138);
nor U13717 (N_13717,N_9225,N_6530);
nand U13718 (N_13718,N_6301,N_6692);
and U13719 (N_13719,N_8061,N_6835);
and U13720 (N_13720,N_8330,N_8937);
nand U13721 (N_13721,N_5927,N_7990);
nor U13722 (N_13722,N_5188,N_6204);
and U13723 (N_13723,N_6858,N_5025);
nand U13724 (N_13724,N_8332,N_5833);
and U13725 (N_13725,N_5299,N_7581);
or U13726 (N_13726,N_9863,N_9733);
or U13727 (N_13727,N_7563,N_9773);
and U13728 (N_13728,N_8361,N_9166);
and U13729 (N_13729,N_7435,N_5522);
xor U13730 (N_13730,N_9509,N_7114);
or U13731 (N_13731,N_6612,N_6317);
nor U13732 (N_13732,N_7736,N_8776);
nor U13733 (N_13733,N_7241,N_8411);
nand U13734 (N_13734,N_5392,N_8311);
nand U13735 (N_13735,N_6662,N_8261);
and U13736 (N_13736,N_8834,N_7112);
nor U13737 (N_13737,N_6417,N_8141);
nand U13738 (N_13738,N_7957,N_6453);
nor U13739 (N_13739,N_5069,N_9102);
xnor U13740 (N_13740,N_9457,N_6259);
or U13741 (N_13741,N_8807,N_5549);
or U13742 (N_13742,N_7719,N_6980);
xor U13743 (N_13743,N_6430,N_9178);
nand U13744 (N_13744,N_7359,N_9457);
and U13745 (N_13745,N_7774,N_7926);
xor U13746 (N_13746,N_7794,N_9193);
xnor U13747 (N_13747,N_6851,N_5336);
and U13748 (N_13748,N_9493,N_5545);
and U13749 (N_13749,N_5084,N_8927);
nand U13750 (N_13750,N_9754,N_9903);
and U13751 (N_13751,N_5043,N_9080);
nand U13752 (N_13752,N_8373,N_8475);
and U13753 (N_13753,N_6175,N_8009);
nand U13754 (N_13754,N_6915,N_9861);
or U13755 (N_13755,N_9574,N_5939);
xnor U13756 (N_13756,N_8149,N_5122);
and U13757 (N_13757,N_9610,N_5591);
and U13758 (N_13758,N_8434,N_6622);
and U13759 (N_13759,N_7986,N_6423);
and U13760 (N_13760,N_7094,N_5553);
xnor U13761 (N_13761,N_6371,N_6203);
or U13762 (N_13762,N_7492,N_7867);
xor U13763 (N_13763,N_9670,N_8177);
nor U13764 (N_13764,N_6979,N_5990);
and U13765 (N_13765,N_7129,N_5470);
nor U13766 (N_13766,N_8267,N_9782);
xor U13767 (N_13767,N_7899,N_9054);
or U13768 (N_13768,N_6097,N_6025);
and U13769 (N_13769,N_9516,N_7121);
or U13770 (N_13770,N_6159,N_7266);
nand U13771 (N_13771,N_7041,N_9520);
nand U13772 (N_13772,N_6194,N_7984);
xor U13773 (N_13773,N_7912,N_5631);
or U13774 (N_13774,N_5373,N_6578);
nor U13775 (N_13775,N_8717,N_9702);
nor U13776 (N_13776,N_8521,N_5338);
nor U13777 (N_13777,N_7169,N_8432);
nand U13778 (N_13778,N_6523,N_5434);
xnor U13779 (N_13779,N_9184,N_9784);
and U13780 (N_13780,N_6204,N_6719);
nand U13781 (N_13781,N_7410,N_7383);
nand U13782 (N_13782,N_9243,N_7975);
or U13783 (N_13783,N_8244,N_8677);
or U13784 (N_13784,N_6131,N_5109);
and U13785 (N_13785,N_8480,N_9185);
nor U13786 (N_13786,N_9551,N_5442);
xnor U13787 (N_13787,N_6515,N_7106);
or U13788 (N_13788,N_5190,N_7284);
xnor U13789 (N_13789,N_6107,N_8013);
xor U13790 (N_13790,N_5623,N_9253);
nand U13791 (N_13791,N_7686,N_5336);
nor U13792 (N_13792,N_6473,N_7282);
nand U13793 (N_13793,N_8602,N_7178);
nand U13794 (N_13794,N_9686,N_8521);
and U13795 (N_13795,N_9036,N_9998);
xnor U13796 (N_13796,N_6386,N_5502);
and U13797 (N_13797,N_9825,N_7657);
or U13798 (N_13798,N_7377,N_6177);
xnor U13799 (N_13799,N_8103,N_5750);
xor U13800 (N_13800,N_9487,N_7726);
and U13801 (N_13801,N_6413,N_9633);
or U13802 (N_13802,N_9140,N_9350);
or U13803 (N_13803,N_9002,N_7169);
xor U13804 (N_13804,N_9820,N_8001);
xnor U13805 (N_13805,N_7901,N_9501);
nand U13806 (N_13806,N_9065,N_7260);
nor U13807 (N_13807,N_8479,N_6319);
xor U13808 (N_13808,N_6308,N_8969);
xor U13809 (N_13809,N_6526,N_5437);
nand U13810 (N_13810,N_5360,N_9304);
or U13811 (N_13811,N_5942,N_6288);
nand U13812 (N_13812,N_8483,N_7214);
xnor U13813 (N_13813,N_7426,N_5576);
xnor U13814 (N_13814,N_7201,N_7952);
nand U13815 (N_13815,N_8711,N_8305);
nand U13816 (N_13816,N_6381,N_9674);
or U13817 (N_13817,N_8932,N_7671);
nand U13818 (N_13818,N_9535,N_8997);
or U13819 (N_13819,N_6501,N_5425);
or U13820 (N_13820,N_6567,N_9809);
xor U13821 (N_13821,N_9041,N_9362);
and U13822 (N_13822,N_7218,N_9074);
nand U13823 (N_13823,N_7517,N_9612);
nor U13824 (N_13824,N_7689,N_9088);
xnor U13825 (N_13825,N_5181,N_6673);
or U13826 (N_13826,N_5019,N_8157);
nand U13827 (N_13827,N_6430,N_7721);
or U13828 (N_13828,N_6268,N_8722);
xnor U13829 (N_13829,N_9997,N_7429);
or U13830 (N_13830,N_9149,N_8767);
or U13831 (N_13831,N_9990,N_8942);
and U13832 (N_13832,N_7098,N_5766);
and U13833 (N_13833,N_9344,N_7325);
xor U13834 (N_13834,N_7493,N_9431);
nor U13835 (N_13835,N_7382,N_9691);
nand U13836 (N_13836,N_7305,N_7610);
and U13837 (N_13837,N_5235,N_7322);
nand U13838 (N_13838,N_7773,N_7928);
xor U13839 (N_13839,N_6968,N_5295);
xor U13840 (N_13840,N_5798,N_7604);
and U13841 (N_13841,N_7627,N_9816);
or U13842 (N_13842,N_5505,N_7210);
nand U13843 (N_13843,N_6737,N_8255);
nand U13844 (N_13844,N_5819,N_9662);
nand U13845 (N_13845,N_8531,N_8175);
xnor U13846 (N_13846,N_6176,N_9666);
xnor U13847 (N_13847,N_8825,N_8643);
or U13848 (N_13848,N_5005,N_7665);
nor U13849 (N_13849,N_5109,N_9122);
and U13850 (N_13850,N_6871,N_5519);
xor U13851 (N_13851,N_6321,N_8490);
xnor U13852 (N_13852,N_9727,N_5968);
or U13853 (N_13853,N_8507,N_9943);
and U13854 (N_13854,N_5161,N_9755);
nor U13855 (N_13855,N_8055,N_6427);
nand U13856 (N_13856,N_9400,N_6257);
nor U13857 (N_13857,N_9125,N_7492);
xnor U13858 (N_13858,N_5839,N_8140);
and U13859 (N_13859,N_5877,N_7346);
nand U13860 (N_13860,N_7234,N_5271);
nor U13861 (N_13861,N_6755,N_9765);
nand U13862 (N_13862,N_8788,N_6731);
nand U13863 (N_13863,N_6387,N_7261);
nand U13864 (N_13864,N_5570,N_7097);
xor U13865 (N_13865,N_7102,N_9710);
or U13866 (N_13866,N_7658,N_8172);
or U13867 (N_13867,N_7972,N_8820);
nor U13868 (N_13868,N_5798,N_5423);
and U13869 (N_13869,N_9436,N_7742);
nor U13870 (N_13870,N_8471,N_8909);
and U13871 (N_13871,N_5837,N_6246);
nor U13872 (N_13872,N_6895,N_7944);
or U13873 (N_13873,N_8485,N_8093);
nand U13874 (N_13874,N_5548,N_9490);
xor U13875 (N_13875,N_9445,N_5274);
and U13876 (N_13876,N_9476,N_9543);
or U13877 (N_13877,N_5981,N_8491);
or U13878 (N_13878,N_6801,N_8034);
and U13879 (N_13879,N_9894,N_5009);
or U13880 (N_13880,N_8371,N_9776);
nor U13881 (N_13881,N_5443,N_6501);
or U13882 (N_13882,N_8814,N_7846);
nor U13883 (N_13883,N_7968,N_9288);
and U13884 (N_13884,N_7376,N_8027);
nand U13885 (N_13885,N_7347,N_7234);
nor U13886 (N_13886,N_5024,N_7782);
nor U13887 (N_13887,N_6221,N_5983);
nand U13888 (N_13888,N_5617,N_9971);
or U13889 (N_13889,N_5864,N_8380);
and U13890 (N_13890,N_8486,N_9953);
and U13891 (N_13891,N_6435,N_7621);
and U13892 (N_13892,N_5116,N_5602);
and U13893 (N_13893,N_9865,N_5468);
nand U13894 (N_13894,N_5657,N_8791);
or U13895 (N_13895,N_9339,N_5568);
nor U13896 (N_13896,N_5177,N_9128);
xor U13897 (N_13897,N_9384,N_8902);
or U13898 (N_13898,N_9208,N_6547);
xnor U13899 (N_13899,N_8021,N_7964);
xnor U13900 (N_13900,N_6411,N_5133);
or U13901 (N_13901,N_7188,N_5066);
xor U13902 (N_13902,N_8586,N_9229);
xnor U13903 (N_13903,N_6765,N_8861);
xor U13904 (N_13904,N_5084,N_7780);
nor U13905 (N_13905,N_6533,N_9210);
nand U13906 (N_13906,N_5133,N_6218);
or U13907 (N_13907,N_9566,N_6174);
nand U13908 (N_13908,N_7621,N_5023);
nor U13909 (N_13909,N_5468,N_5174);
or U13910 (N_13910,N_8227,N_9892);
nor U13911 (N_13911,N_9902,N_5931);
nor U13912 (N_13912,N_7674,N_7604);
or U13913 (N_13913,N_7739,N_5376);
or U13914 (N_13914,N_7364,N_5454);
xor U13915 (N_13915,N_8300,N_8376);
nand U13916 (N_13916,N_7883,N_7709);
and U13917 (N_13917,N_6590,N_9708);
nor U13918 (N_13918,N_8732,N_8524);
nand U13919 (N_13919,N_7838,N_7770);
xnor U13920 (N_13920,N_7290,N_6297);
xor U13921 (N_13921,N_5407,N_9994);
or U13922 (N_13922,N_9338,N_8114);
xor U13923 (N_13923,N_5132,N_6969);
nand U13924 (N_13924,N_5430,N_9628);
xnor U13925 (N_13925,N_7045,N_9535);
nor U13926 (N_13926,N_5521,N_7811);
or U13927 (N_13927,N_5062,N_7602);
xnor U13928 (N_13928,N_5999,N_5428);
or U13929 (N_13929,N_7797,N_5151);
nand U13930 (N_13930,N_9700,N_5316);
nand U13931 (N_13931,N_8353,N_5108);
and U13932 (N_13932,N_9887,N_6911);
or U13933 (N_13933,N_7599,N_9527);
nor U13934 (N_13934,N_7249,N_6526);
and U13935 (N_13935,N_7873,N_5541);
nand U13936 (N_13936,N_6796,N_5388);
and U13937 (N_13937,N_9842,N_5142);
nand U13938 (N_13938,N_9891,N_9473);
nand U13939 (N_13939,N_8682,N_9805);
and U13940 (N_13940,N_7827,N_7898);
or U13941 (N_13941,N_7673,N_9123);
or U13942 (N_13942,N_6722,N_8889);
and U13943 (N_13943,N_9641,N_7250);
nand U13944 (N_13944,N_6357,N_9948);
xnor U13945 (N_13945,N_9557,N_6119);
nor U13946 (N_13946,N_5490,N_5754);
and U13947 (N_13947,N_8964,N_6767);
xnor U13948 (N_13948,N_7070,N_7812);
nand U13949 (N_13949,N_5713,N_6792);
xnor U13950 (N_13950,N_5379,N_8740);
and U13951 (N_13951,N_7246,N_6610);
nor U13952 (N_13952,N_6500,N_8987);
or U13953 (N_13953,N_9656,N_7447);
nor U13954 (N_13954,N_8042,N_7587);
xor U13955 (N_13955,N_6536,N_6967);
and U13956 (N_13956,N_5114,N_7013);
nor U13957 (N_13957,N_6294,N_7066);
nor U13958 (N_13958,N_9106,N_5928);
xor U13959 (N_13959,N_6032,N_8949);
or U13960 (N_13960,N_9165,N_9103);
nand U13961 (N_13961,N_6693,N_5968);
xnor U13962 (N_13962,N_6721,N_6783);
nor U13963 (N_13963,N_5641,N_6712);
nand U13964 (N_13964,N_9886,N_9588);
xor U13965 (N_13965,N_8650,N_6072);
xnor U13966 (N_13966,N_5110,N_9875);
or U13967 (N_13967,N_6616,N_6320);
nand U13968 (N_13968,N_9487,N_7719);
xor U13969 (N_13969,N_9437,N_6211);
nor U13970 (N_13970,N_5447,N_6198);
and U13971 (N_13971,N_9755,N_7116);
xor U13972 (N_13972,N_6267,N_7585);
or U13973 (N_13973,N_6365,N_8835);
nor U13974 (N_13974,N_5657,N_8461);
and U13975 (N_13975,N_9601,N_5394);
nand U13976 (N_13976,N_7618,N_8139);
nand U13977 (N_13977,N_8560,N_8825);
or U13978 (N_13978,N_7378,N_6805);
nand U13979 (N_13979,N_9390,N_9106);
or U13980 (N_13980,N_6517,N_8814);
nor U13981 (N_13981,N_5012,N_5212);
or U13982 (N_13982,N_8541,N_8290);
and U13983 (N_13983,N_8447,N_5437);
or U13984 (N_13984,N_5099,N_5404);
and U13985 (N_13985,N_9716,N_7680);
or U13986 (N_13986,N_5605,N_6290);
or U13987 (N_13987,N_6556,N_6093);
nor U13988 (N_13988,N_7345,N_5311);
nand U13989 (N_13989,N_6771,N_6664);
or U13990 (N_13990,N_6782,N_6659);
or U13991 (N_13991,N_8275,N_9029);
nor U13992 (N_13992,N_7207,N_7469);
nand U13993 (N_13993,N_7446,N_8588);
xnor U13994 (N_13994,N_6153,N_9625);
nand U13995 (N_13995,N_6037,N_8568);
nor U13996 (N_13996,N_5128,N_5123);
and U13997 (N_13997,N_8322,N_6425);
or U13998 (N_13998,N_5716,N_8818);
nor U13999 (N_13999,N_6193,N_5009);
and U14000 (N_14000,N_9435,N_9704);
xor U14001 (N_14001,N_9406,N_9639);
or U14002 (N_14002,N_9569,N_7048);
or U14003 (N_14003,N_9882,N_5019);
nor U14004 (N_14004,N_5032,N_5953);
and U14005 (N_14005,N_8101,N_9851);
or U14006 (N_14006,N_9049,N_6411);
or U14007 (N_14007,N_5356,N_8326);
nand U14008 (N_14008,N_6445,N_8725);
nand U14009 (N_14009,N_9620,N_7502);
and U14010 (N_14010,N_9192,N_8456);
xnor U14011 (N_14011,N_6608,N_6554);
nor U14012 (N_14012,N_9928,N_8158);
nor U14013 (N_14013,N_5990,N_5800);
nand U14014 (N_14014,N_5021,N_5883);
nand U14015 (N_14015,N_8686,N_9655);
and U14016 (N_14016,N_7878,N_8263);
nand U14017 (N_14017,N_9538,N_6890);
xnor U14018 (N_14018,N_9744,N_8292);
xnor U14019 (N_14019,N_5846,N_9855);
nor U14020 (N_14020,N_6355,N_5143);
and U14021 (N_14021,N_5081,N_5385);
xor U14022 (N_14022,N_6763,N_6605);
and U14023 (N_14023,N_5367,N_6222);
xnor U14024 (N_14024,N_7944,N_7317);
or U14025 (N_14025,N_7239,N_7883);
nor U14026 (N_14026,N_5251,N_9831);
and U14027 (N_14027,N_5731,N_8528);
or U14028 (N_14028,N_8366,N_8102);
xnor U14029 (N_14029,N_5408,N_7524);
or U14030 (N_14030,N_7933,N_6363);
nor U14031 (N_14031,N_5844,N_5284);
and U14032 (N_14032,N_7014,N_5572);
nand U14033 (N_14033,N_5424,N_7618);
or U14034 (N_14034,N_9235,N_7765);
nand U14035 (N_14035,N_9331,N_8302);
nor U14036 (N_14036,N_6286,N_7814);
xor U14037 (N_14037,N_9021,N_9681);
and U14038 (N_14038,N_6206,N_7481);
xor U14039 (N_14039,N_8400,N_6165);
and U14040 (N_14040,N_5516,N_8251);
nand U14041 (N_14041,N_7728,N_9281);
or U14042 (N_14042,N_7827,N_8877);
and U14043 (N_14043,N_6308,N_6406);
nand U14044 (N_14044,N_9103,N_5141);
nor U14045 (N_14045,N_7760,N_7562);
or U14046 (N_14046,N_5266,N_5628);
nor U14047 (N_14047,N_5704,N_9831);
nor U14048 (N_14048,N_7901,N_7504);
xor U14049 (N_14049,N_9621,N_5820);
xnor U14050 (N_14050,N_8878,N_7379);
and U14051 (N_14051,N_5113,N_5867);
or U14052 (N_14052,N_5743,N_6031);
nor U14053 (N_14053,N_5092,N_7515);
xor U14054 (N_14054,N_7148,N_5445);
nor U14055 (N_14055,N_5508,N_8204);
xnor U14056 (N_14056,N_5825,N_9662);
nor U14057 (N_14057,N_9133,N_5371);
or U14058 (N_14058,N_5000,N_8790);
or U14059 (N_14059,N_8579,N_8880);
and U14060 (N_14060,N_9446,N_9793);
nand U14061 (N_14061,N_7829,N_6257);
or U14062 (N_14062,N_9733,N_8367);
xnor U14063 (N_14063,N_6671,N_6369);
or U14064 (N_14064,N_9745,N_5556);
nand U14065 (N_14065,N_7997,N_9013);
and U14066 (N_14066,N_5090,N_9918);
xor U14067 (N_14067,N_7733,N_7590);
nand U14068 (N_14068,N_5899,N_9554);
or U14069 (N_14069,N_9438,N_6201);
or U14070 (N_14070,N_8626,N_8969);
and U14071 (N_14071,N_6703,N_5288);
nand U14072 (N_14072,N_5874,N_5077);
and U14073 (N_14073,N_9278,N_9647);
nor U14074 (N_14074,N_5598,N_8961);
and U14075 (N_14075,N_6177,N_9342);
nor U14076 (N_14076,N_5847,N_7049);
nor U14077 (N_14077,N_5383,N_8531);
nor U14078 (N_14078,N_7145,N_7046);
xnor U14079 (N_14079,N_9400,N_6898);
and U14080 (N_14080,N_6858,N_5131);
nor U14081 (N_14081,N_6346,N_5432);
xnor U14082 (N_14082,N_8969,N_6777);
and U14083 (N_14083,N_5083,N_5624);
nand U14084 (N_14084,N_8880,N_7799);
nand U14085 (N_14085,N_9594,N_9499);
or U14086 (N_14086,N_6863,N_8623);
and U14087 (N_14087,N_8349,N_5224);
nor U14088 (N_14088,N_5650,N_9892);
and U14089 (N_14089,N_6576,N_9960);
or U14090 (N_14090,N_7767,N_8124);
nor U14091 (N_14091,N_5950,N_8120);
nor U14092 (N_14092,N_7348,N_5504);
nor U14093 (N_14093,N_7251,N_8861);
nand U14094 (N_14094,N_5014,N_9188);
or U14095 (N_14095,N_7789,N_8074);
nor U14096 (N_14096,N_9030,N_7026);
xor U14097 (N_14097,N_5205,N_9907);
xnor U14098 (N_14098,N_6320,N_6944);
xor U14099 (N_14099,N_8416,N_5460);
nand U14100 (N_14100,N_6489,N_6244);
xnor U14101 (N_14101,N_9261,N_9203);
or U14102 (N_14102,N_9173,N_8289);
or U14103 (N_14103,N_9359,N_6017);
or U14104 (N_14104,N_8590,N_6700);
nor U14105 (N_14105,N_9250,N_9200);
and U14106 (N_14106,N_8519,N_7136);
and U14107 (N_14107,N_9570,N_8793);
nor U14108 (N_14108,N_9033,N_7777);
nor U14109 (N_14109,N_9141,N_9052);
nor U14110 (N_14110,N_5849,N_5753);
and U14111 (N_14111,N_5051,N_9152);
nor U14112 (N_14112,N_9044,N_7054);
nor U14113 (N_14113,N_7279,N_9873);
xor U14114 (N_14114,N_5993,N_6726);
nor U14115 (N_14115,N_9528,N_9681);
nor U14116 (N_14116,N_7910,N_8879);
or U14117 (N_14117,N_6981,N_8468);
nand U14118 (N_14118,N_6961,N_9533);
and U14119 (N_14119,N_9068,N_8279);
xor U14120 (N_14120,N_5736,N_6077);
nor U14121 (N_14121,N_6347,N_5577);
nor U14122 (N_14122,N_6611,N_5754);
xor U14123 (N_14123,N_7458,N_6974);
and U14124 (N_14124,N_6873,N_8293);
nor U14125 (N_14125,N_6786,N_7555);
and U14126 (N_14126,N_9460,N_7053);
nand U14127 (N_14127,N_6269,N_5920);
and U14128 (N_14128,N_6661,N_8311);
xnor U14129 (N_14129,N_8494,N_5509);
nand U14130 (N_14130,N_7146,N_7554);
nor U14131 (N_14131,N_6066,N_8103);
nand U14132 (N_14132,N_9707,N_9021);
xor U14133 (N_14133,N_7360,N_8324);
nand U14134 (N_14134,N_8181,N_7165);
nor U14135 (N_14135,N_9654,N_5860);
nand U14136 (N_14136,N_6409,N_5859);
and U14137 (N_14137,N_6140,N_6549);
or U14138 (N_14138,N_5938,N_6774);
xnor U14139 (N_14139,N_8120,N_9044);
and U14140 (N_14140,N_5635,N_7509);
xor U14141 (N_14141,N_8554,N_9181);
or U14142 (N_14142,N_5164,N_9593);
xor U14143 (N_14143,N_7515,N_8520);
xnor U14144 (N_14144,N_5206,N_7064);
nor U14145 (N_14145,N_9487,N_8662);
nor U14146 (N_14146,N_9842,N_7536);
nor U14147 (N_14147,N_5883,N_5012);
or U14148 (N_14148,N_5318,N_6120);
xor U14149 (N_14149,N_8850,N_7396);
or U14150 (N_14150,N_9351,N_6612);
or U14151 (N_14151,N_9129,N_7026);
xor U14152 (N_14152,N_7642,N_7394);
nand U14153 (N_14153,N_8887,N_6394);
nor U14154 (N_14154,N_7115,N_7756);
and U14155 (N_14155,N_7194,N_6512);
and U14156 (N_14156,N_8588,N_8908);
xor U14157 (N_14157,N_6561,N_6068);
and U14158 (N_14158,N_8172,N_5905);
and U14159 (N_14159,N_9837,N_9692);
xnor U14160 (N_14160,N_5136,N_7832);
and U14161 (N_14161,N_5382,N_6349);
and U14162 (N_14162,N_7202,N_8190);
nor U14163 (N_14163,N_9894,N_9063);
or U14164 (N_14164,N_5245,N_7341);
and U14165 (N_14165,N_6791,N_6343);
xnor U14166 (N_14166,N_9082,N_5376);
and U14167 (N_14167,N_9249,N_7805);
nor U14168 (N_14168,N_8665,N_6129);
nand U14169 (N_14169,N_8144,N_6459);
or U14170 (N_14170,N_6397,N_8404);
and U14171 (N_14171,N_6079,N_6808);
xnor U14172 (N_14172,N_7060,N_9877);
and U14173 (N_14173,N_7450,N_6773);
xnor U14174 (N_14174,N_5426,N_8021);
nor U14175 (N_14175,N_7280,N_7093);
nor U14176 (N_14176,N_9488,N_7995);
nand U14177 (N_14177,N_7009,N_5264);
nor U14178 (N_14178,N_6113,N_6268);
nand U14179 (N_14179,N_5184,N_7951);
nand U14180 (N_14180,N_9994,N_7571);
xnor U14181 (N_14181,N_6001,N_5901);
or U14182 (N_14182,N_9814,N_7131);
nor U14183 (N_14183,N_9577,N_5401);
nor U14184 (N_14184,N_6607,N_9887);
nor U14185 (N_14185,N_5408,N_9077);
nor U14186 (N_14186,N_6308,N_5810);
xor U14187 (N_14187,N_5968,N_9781);
xor U14188 (N_14188,N_5741,N_5620);
nand U14189 (N_14189,N_7719,N_9098);
and U14190 (N_14190,N_8047,N_9486);
or U14191 (N_14191,N_5091,N_6623);
xnor U14192 (N_14192,N_6017,N_8956);
or U14193 (N_14193,N_6167,N_5537);
nor U14194 (N_14194,N_7896,N_7765);
nor U14195 (N_14195,N_7716,N_7482);
nor U14196 (N_14196,N_7098,N_8243);
nand U14197 (N_14197,N_6070,N_8598);
nand U14198 (N_14198,N_5360,N_7259);
nand U14199 (N_14199,N_5270,N_5534);
xor U14200 (N_14200,N_9300,N_8279);
nand U14201 (N_14201,N_7276,N_6406);
nor U14202 (N_14202,N_6597,N_7028);
xnor U14203 (N_14203,N_7966,N_9173);
and U14204 (N_14204,N_5622,N_7139);
or U14205 (N_14205,N_9806,N_8058);
nor U14206 (N_14206,N_9804,N_6417);
and U14207 (N_14207,N_9011,N_5273);
xor U14208 (N_14208,N_6287,N_8907);
and U14209 (N_14209,N_5923,N_5449);
nand U14210 (N_14210,N_6015,N_6007);
and U14211 (N_14211,N_8504,N_7221);
and U14212 (N_14212,N_5262,N_6308);
xor U14213 (N_14213,N_5288,N_6841);
and U14214 (N_14214,N_5975,N_7241);
nand U14215 (N_14215,N_5634,N_5426);
nand U14216 (N_14216,N_9299,N_9214);
or U14217 (N_14217,N_6158,N_9724);
or U14218 (N_14218,N_5808,N_6701);
or U14219 (N_14219,N_9913,N_7595);
or U14220 (N_14220,N_6908,N_6230);
or U14221 (N_14221,N_9543,N_8279);
or U14222 (N_14222,N_9350,N_8946);
xnor U14223 (N_14223,N_7487,N_6815);
or U14224 (N_14224,N_5036,N_9918);
or U14225 (N_14225,N_5946,N_8623);
xor U14226 (N_14226,N_5048,N_5103);
nor U14227 (N_14227,N_9948,N_6692);
nand U14228 (N_14228,N_6193,N_6413);
nor U14229 (N_14229,N_8992,N_5602);
xnor U14230 (N_14230,N_7951,N_9733);
nor U14231 (N_14231,N_5561,N_8132);
and U14232 (N_14232,N_6244,N_7574);
or U14233 (N_14233,N_7782,N_9541);
xor U14234 (N_14234,N_7931,N_7552);
or U14235 (N_14235,N_9451,N_8888);
xor U14236 (N_14236,N_5461,N_9067);
and U14237 (N_14237,N_8219,N_5296);
or U14238 (N_14238,N_9286,N_9866);
nor U14239 (N_14239,N_7094,N_7647);
xor U14240 (N_14240,N_7470,N_9104);
xnor U14241 (N_14241,N_6504,N_5321);
xor U14242 (N_14242,N_5265,N_8398);
xnor U14243 (N_14243,N_9757,N_5227);
or U14244 (N_14244,N_7054,N_7999);
and U14245 (N_14245,N_6913,N_5049);
nor U14246 (N_14246,N_7090,N_8661);
nor U14247 (N_14247,N_5115,N_9617);
or U14248 (N_14248,N_8371,N_7297);
nand U14249 (N_14249,N_7007,N_8842);
nand U14250 (N_14250,N_9869,N_6059);
nand U14251 (N_14251,N_9649,N_8227);
or U14252 (N_14252,N_9655,N_5424);
and U14253 (N_14253,N_8317,N_6039);
xnor U14254 (N_14254,N_6425,N_5907);
nor U14255 (N_14255,N_7271,N_9076);
xnor U14256 (N_14256,N_5250,N_7534);
nor U14257 (N_14257,N_8090,N_8385);
xor U14258 (N_14258,N_7982,N_6343);
nand U14259 (N_14259,N_6351,N_9124);
nor U14260 (N_14260,N_9128,N_8101);
nand U14261 (N_14261,N_8330,N_6364);
or U14262 (N_14262,N_6216,N_8159);
nand U14263 (N_14263,N_6793,N_8777);
or U14264 (N_14264,N_7789,N_5456);
nand U14265 (N_14265,N_5673,N_7677);
or U14266 (N_14266,N_6253,N_9852);
or U14267 (N_14267,N_5550,N_7019);
or U14268 (N_14268,N_8772,N_5028);
nor U14269 (N_14269,N_6429,N_6033);
xnor U14270 (N_14270,N_9906,N_5732);
nor U14271 (N_14271,N_9922,N_7503);
and U14272 (N_14272,N_6870,N_9626);
xnor U14273 (N_14273,N_7037,N_8929);
and U14274 (N_14274,N_5279,N_7702);
xor U14275 (N_14275,N_9271,N_5898);
or U14276 (N_14276,N_6658,N_5379);
nor U14277 (N_14277,N_5897,N_5627);
and U14278 (N_14278,N_7092,N_8796);
nor U14279 (N_14279,N_7946,N_5636);
xor U14280 (N_14280,N_8202,N_8073);
nand U14281 (N_14281,N_5265,N_7936);
xor U14282 (N_14282,N_7330,N_6704);
and U14283 (N_14283,N_5527,N_8542);
nor U14284 (N_14284,N_5178,N_9749);
and U14285 (N_14285,N_6104,N_5036);
or U14286 (N_14286,N_8312,N_6941);
and U14287 (N_14287,N_9671,N_5543);
or U14288 (N_14288,N_6266,N_7677);
xnor U14289 (N_14289,N_5401,N_9694);
xor U14290 (N_14290,N_5298,N_6562);
nand U14291 (N_14291,N_5992,N_7945);
nor U14292 (N_14292,N_9799,N_9372);
or U14293 (N_14293,N_5178,N_8001);
and U14294 (N_14294,N_9562,N_8311);
and U14295 (N_14295,N_7220,N_5672);
nor U14296 (N_14296,N_8971,N_7536);
nor U14297 (N_14297,N_6188,N_5611);
or U14298 (N_14298,N_7520,N_7851);
xor U14299 (N_14299,N_8862,N_5877);
and U14300 (N_14300,N_6449,N_7574);
nor U14301 (N_14301,N_5778,N_8785);
nand U14302 (N_14302,N_5247,N_9964);
and U14303 (N_14303,N_9842,N_6442);
and U14304 (N_14304,N_8181,N_5305);
xor U14305 (N_14305,N_6533,N_5211);
and U14306 (N_14306,N_7180,N_8104);
xor U14307 (N_14307,N_8297,N_5318);
or U14308 (N_14308,N_6120,N_6247);
and U14309 (N_14309,N_6119,N_5130);
or U14310 (N_14310,N_6115,N_5448);
or U14311 (N_14311,N_6782,N_5395);
xor U14312 (N_14312,N_8230,N_9127);
or U14313 (N_14313,N_5613,N_9917);
nor U14314 (N_14314,N_6698,N_9753);
xor U14315 (N_14315,N_7713,N_9500);
or U14316 (N_14316,N_7342,N_7236);
xnor U14317 (N_14317,N_8070,N_5747);
nand U14318 (N_14318,N_9168,N_6015);
and U14319 (N_14319,N_7656,N_7067);
nor U14320 (N_14320,N_7143,N_5752);
and U14321 (N_14321,N_5545,N_9909);
or U14322 (N_14322,N_9846,N_9774);
and U14323 (N_14323,N_8635,N_8866);
nor U14324 (N_14324,N_5713,N_5021);
nand U14325 (N_14325,N_5673,N_5039);
and U14326 (N_14326,N_8218,N_8279);
nand U14327 (N_14327,N_8373,N_6874);
nor U14328 (N_14328,N_5281,N_5130);
and U14329 (N_14329,N_6737,N_9392);
nand U14330 (N_14330,N_6219,N_6405);
nand U14331 (N_14331,N_9469,N_5499);
xnor U14332 (N_14332,N_7493,N_7755);
nor U14333 (N_14333,N_8347,N_8827);
xnor U14334 (N_14334,N_6082,N_9793);
xor U14335 (N_14335,N_5613,N_9214);
and U14336 (N_14336,N_8067,N_8333);
xor U14337 (N_14337,N_5814,N_6541);
and U14338 (N_14338,N_8793,N_5197);
xnor U14339 (N_14339,N_5592,N_9975);
and U14340 (N_14340,N_7376,N_8928);
xor U14341 (N_14341,N_5238,N_5942);
nor U14342 (N_14342,N_6404,N_7660);
nand U14343 (N_14343,N_8077,N_5525);
xor U14344 (N_14344,N_5586,N_9041);
nand U14345 (N_14345,N_9240,N_5177);
nand U14346 (N_14346,N_6259,N_5659);
xor U14347 (N_14347,N_8661,N_9072);
nor U14348 (N_14348,N_8623,N_8511);
or U14349 (N_14349,N_9719,N_9702);
nand U14350 (N_14350,N_8197,N_7290);
nor U14351 (N_14351,N_8452,N_9808);
xor U14352 (N_14352,N_6069,N_9716);
xnor U14353 (N_14353,N_9037,N_6376);
or U14354 (N_14354,N_5173,N_9627);
xnor U14355 (N_14355,N_7168,N_6980);
and U14356 (N_14356,N_5095,N_6746);
nand U14357 (N_14357,N_9481,N_7037);
or U14358 (N_14358,N_7010,N_9545);
nand U14359 (N_14359,N_7972,N_9046);
and U14360 (N_14360,N_7630,N_5527);
xnor U14361 (N_14361,N_8838,N_9979);
and U14362 (N_14362,N_5469,N_5609);
xor U14363 (N_14363,N_7293,N_6054);
nand U14364 (N_14364,N_9511,N_9034);
nor U14365 (N_14365,N_9992,N_9692);
nor U14366 (N_14366,N_7284,N_8532);
nand U14367 (N_14367,N_8734,N_9797);
or U14368 (N_14368,N_5603,N_8115);
or U14369 (N_14369,N_9038,N_9243);
or U14370 (N_14370,N_9390,N_8803);
and U14371 (N_14371,N_5058,N_6947);
xor U14372 (N_14372,N_7396,N_8601);
nor U14373 (N_14373,N_6579,N_5998);
or U14374 (N_14374,N_7140,N_9936);
and U14375 (N_14375,N_7661,N_6134);
xor U14376 (N_14376,N_7954,N_6668);
nor U14377 (N_14377,N_6945,N_5351);
or U14378 (N_14378,N_5745,N_8893);
nand U14379 (N_14379,N_6176,N_8371);
nand U14380 (N_14380,N_7752,N_7302);
nand U14381 (N_14381,N_9433,N_8326);
and U14382 (N_14382,N_7026,N_7059);
nand U14383 (N_14383,N_5501,N_9151);
and U14384 (N_14384,N_5883,N_5288);
and U14385 (N_14385,N_6502,N_8684);
nor U14386 (N_14386,N_5853,N_6970);
nor U14387 (N_14387,N_5471,N_8050);
nand U14388 (N_14388,N_5350,N_5681);
or U14389 (N_14389,N_8879,N_7550);
and U14390 (N_14390,N_5237,N_6221);
and U14391 (N_14391,N_8190,N_5772);
or U14392 (N_14392,N_6988,N_6835);
nor U14393 (N_14393,N_5169,N_6888);
or U14394 (N_14394,N_9889,N_8968);
nand U14395 (N_14395,N_9715,N_6470);
nor U14396 (N_14396,N_7859,N_7134);
nand U14397 (N_14397,N_9717,N_8987);
xnor U14398 (N_14398,N_8915,N_7079);
nand U14399 (N_14399,N_9735,N_7999);
or U14400 (N_14400,N_6848,N_9811);
and U14401 (N_14401,N_7611,N_5831);
xor U14402 (N_14402,N_5792,N_8733);
xor U14403 (N_14403,N_9638,N_6892);
and U14404 (N_14404,N_7687,N_8809);
xnor U14405 (N_14405,N_6727,N_9506);
and U14406 (N_14406,N_7009,N_8189);
nor U14407 (N_14407,N_8992,N_7445);
xnor U14408 (N_14408,N_8736,N_7492);
or U14409 (N_14409,N_5920,N_5888);
and U14410 (N_14410,N_7579,N_6694);
and U14411 (N_14411,N_9088,N_9906);
nand U14412 (N_14412,N_7057,N_5506);
nand U14413 (N_14413,N_8177,N_6621);
or U14414 (N_14414,N_7295,N_7124);
nor U14415 (N_14415,N_8169,N_9911);
or U14416 (N_14416,N_8138,N_9805);
xnor U14417 (N_14417,N_9051,N_6218);
nand U14418 (N_14418,N_7392,N_9175);
xor U14419 (N_14419,N_5975,N_6283);
or U14420 (N_14420,N_5514,N_5727);
xnor U14421 (N_14421,N_8866,N_9088);
xnor U14422 (N_14422,N_9655,N_5845);
or U14423 (N_14423,N_8929,N_8978);
xor U14424 (N_14424,N_7494,N_8221);
or U14425 (N_14425,N_8533,N_7230);
and U14426 (N_14426,N_5232,N_7748);
xnor U14427 (N_14427,N_9725,N_7587);
nand U14428 (N_14428,N_5450,N_8954);
nor U14429 (N_14429,N_8588,N_7103);
nand U14430 (N_14430,N_7669,N_5157);
xnor U14431 (N_14431,N_8135,N_8942);
nor U14432 (N_14432,N_7120,N_7974);
xor U14433 (N_14433,N_8760,N_5837);
nand U14434 (N_14434,N_6511,N_8172);
nor U14435 (N_14435,N_7907,N_8590);
and U14436 (N_14436,N_6921,N_5834);
and U14437 (N_14437,N_7525,N_8234);
or U14438 (N_14438,N_7862,N_7550);
xor U14439 (N_14439,N_5944,N_5162);
nand U14440 (N_14440,N_5528,N_6182);
and U14441 (N_14441,N_5757,N_8211);
or U14442 (N_14442,N_6582,N_6721);
xor U14443 (N_14443,N_5364,N_7049);
and U14444 (N_14444,N_7574,N_5422);
nor U14445 (N_14445,N_8884,N_7930);
and U14446 (N_14446,N_7078,N_6488);
nor U14447 (N_14447,N_8277,N_6224);
xor U14448 (N_14448,N_9696,N_8152);
nor U14449 (N_14449,N_7753,N_5022);
xor U14450 (N_14450,N_7761,N_7539);
nand U14451 (N_14451,N_5008,N_7489);
nand U14452 (N_14452,N_9274,N_7001);
nand U14453 (N_14453,N_5289,N_5097);
nor U14454 (N_14454,N_7169,N_5667);
nor U14455 (N_14455,N_5233,N_9821);
nand U14456 (N_14456,N_9694,N_6858);
xor U14457 (N_14457,N_9272,N_7426);
or U14458 (N_14458,N_5213,N_5658);
or U14459 (N_14459,N_8510,N_9084);
xor U14460 (N_14460,N_6151,N_8162);
and U14461 (N_14461,N_7349,N_9893);
or U14462 (N_14462,N_8393,N_8232);
or U14463 (N_14463,N_6851,N_6896);
nand U14464 (N_14464,N_7036,N_6239);
nor U14465 (N_14465,N_7635,N_8476);
nor U14466 (N_14466,N_9769,N_6152);
or U14467 (N_14467,N_6152,N_9627);
nor U14468 (N_14468,N_7417,N_6325);
nand U14469 (N_14469,N_6318,N_9560);
or U14470 (N_14470,N_8957,N_9763);
or U14471 (N_14471,N_5421,N_6024);
xor U14472 (N_14472,N_8574,N_9337);
and U14473 (N_14473,N_9016,N_5869);
and U14474 (N_14474,N_7234,N_6807);
nand U14475 (N_14475,N_9972,N_9830);
and U14476 (N_14476,N_8268,N_8766);
nor U14477 (N_14477,N_5911,N_8303);
nand U14478 (N_14478,N_8770,N_7455);
xnor U14479 (N_14479,N_7737,N_5328);
nand U14480 (N_14480,N_5274,N_8795);
nand U14481 (N_14481,N_7628,N_8873);
nand U14482 (N_14482,N_8548,N_8944);
xnor U14483 (N_14483,N_6471,N_8156);
and U14484 (N_14484,N_7578,N_7592);
nor U14485 (N_14485,N_5636,N_5942);
nand U14486 (N_14486,N_9321,N_9956);
nand U14487 (N_14487,N_8658,N_8488);
xor U14488 (N_14488,N_7081,N_7994);
xor U14489 (N_14489,N_7579,N_9391);
and U14490 (N_14490,N_5049,N_5165);
nor U14491 (N_14491,N_5471,N_7509);
or U14492 (N_14492,N_8176,N_5854);
or U14493 (N_14493,N_7843,N_5831);
nand U14494 (N_14494,N_8317,N_9633);
or U14495 (N_14495,N_6695,N_5004);
and U14496 (N_14496,N_5643,N_5142);
xor U14497 (N_14497,N_9236,N_8411);
or U14498 (N_14498,N_7610,N_7977);
and U14499 (N_14499,N_9928,N_9648);
nor U14500 (N_14500,N_9812,N_5145);
nor U14501 (N_14501,N_8885,N_5751);
xnor U14502 (N_14502,N_5613,N_8983);
nand U14503 (N_14503,N_5845,N_6410);
or U14504 (N_14504,N_8914,N_5517);
nor U14505 (N_14505,N_9950,N_6922);
xor U14506 (N_14506,N_8159,N_9617);
and U14507 (N_14507,N_9478,N_9391);
nor U14508 (N_14508,N_5343,N_7065);
nor U14509 (N_14509,N_7278,N_8203);
nor U14510 (N_14510,N_9817,N_6183);
nand U14511 (N_14511,N_5076,N_6485);
or U14512 (N_14512,N_6598,N_5975);
and U14513 (N_14513,N_6646,N_5771);
nor U14514 (N_14514,N_5662,N_8325);
xnor U14515 (N_14515,N_5685,N_5944);
xnor U14516 (N_14516,N_8882,N_6602);
nand U14517 (N_14517,N_7966,N_7845);
or U14518 (N_14518,N_5167,N_6193);
nor U14519 (N_14519,N_6322,N_9683);
xnor U14520 (N_14520,N_9705,N_9345);
and U14521 (N_14521,N_6338,N_8523);
or U14522 (N_14522,N_6651,N_9906);
or U14523 (N_14523,N_9681,N_7821);
nor U14524 (N_14524,N_8052,N_8236);
and U14525 (N_14525,N_5140,N_6991);
xor U14526 (N_14526,N_5668,N_6817);
or U14527 (N_14527,N_7561,N_7704);
nand U14528 (N_14528,N_8338,N_8057);
xnor U14529 (N_14529,N_8193,N_8371);
nor U14530 (N_14530,N_5654,N_5697);
and U14531 (N_14531,N_5245,N_7955);
xnor U14532 (N_14532,N_8073,N_9124);
and U14533 (N_14533,N_7905,N_7234);
nand U14534 (N_14534,N_7728,N_6156);
or U14535 (N_14535,N_9376,N_5211);
nand U14536 (N_14536,N_5981,N_7779);
nor U14537 (N_14537,N_7218,N_7392);
or U14538 (N_14538,N_6257,N_5282);
xnor U14539 (N_14539,N_6960,N_7862);
or U14540 (N_14540,N_7532,N_8920);
or U14541 (N_14541,N_8330,N_9305);
nor U14542 (N_14542,N_5837,N_8295);
xnor U14543 (N_14543,N_8755,N_5846);
nor U14544 (N_14544,N_8767,N_7518);
or U14545 (N_14545,N_5946,N_9957);
and U14546 (N_14546,N_6511,N_8554);
or U14547 (N_14547,N_8878,N_9016);
or U14548 (N_14548,N_8612,N_8519);
nor U14549 (N_14549,N_7950,N_7251);
and U14550 (N_14550,N_6790,N_8024);
nand U14551 (N_14551,N_5331,N_6740);
or U14552 (N_14552,N_9481,N_6096);
and U14553 (N_14553,N_5417,N_6347);
and U14554 (N_14554,N_7822,N_5719);
and U14555 (N_14555,N_6885,N_7373);
nor U14556 (N_14556,N_6315,N_7038);
nand U14557 (N_14557,N_8831,N_8754);
nand U14558 (N_14558,N_6149,N_9901);
or U14559 (N_14559,N_5515,N_9982);
or U14560 (N_14560,N_7782,N_6765);
and U14561 (N_14561,N_8139,N_5764);
and U14562 (N_14562,N_5791,N_8512);
and U14563 (N_14563,N_9900,N_5253);
nor U14564 (N_14564,N_7084,N_7535);
nand U14565 (N_14565,N_8756,N_9652);
nor U14566 (N_14566,N_7101,N_8507);
nor U14567 (N_14567,N_8844,N_5543);
nor U14568 (N_14568,N_6001,N_7311);
or U14569 (N_14569,N_6051,N_9559);
and U14570 (N_14570,N_9248,N_7699);
nand U14571 (N_14571,N_5725,N_5225);
and U14572 (N_14572,N_7807,N_8916);
and U14573 (N_14573,N_6829,N_6452);
nand U14574 (N_14574,N_7161,N_9567);
and U14575 (N_14575,N_6366,N_9845);
nand U14576 (N_14576,N_7903,N_8740);
nand U14577 (N_14577,N_8318,N_7688);
xnor U14578 (N_14578,N_6005,N_9058);
and U14579 (N_14579,N_7002,N_7501);
or U14580 (N_14580,N_7548,N_6524);
nor U14581 (N_14581,N_5384,N_5413);
or U14582 (N_14582,N_7121,N_6503);
and U14583 (N_14583,N_9037,N_7042);
nand U14584 (N_14584,N_8051,N_6347);
xor U14585 (N_14585,N_7316,N_6314);
nand U14586 (N_14586,N_6996,N_9779);
and U14587 (N_14587,N_7138,N_9996);
or U14588 (N_14588,N_6529,N_8481);
nor U14589 (N_14589,N_9957,N_8392);
nand U14590 (N_14590,N_9358,N_8551);
nor U14591 (N_14591,N_8919,N_6315);
or U14592 (N_14592,N_5162,N_9511);
and U14593 (N_14593,N_7458,N_5487);
xor U14594 (N_14594,N_5246,N_6645);
or U14595 (N_14595,N_9190,N_7258);
nor U14596 (N_14596,N_6834,N_8978);
xnor U14597 (N_14597,N_5784,N_8522);
and U14598 (N_14598,N_5102,N_9562);
xor U14599 (N_14599,N_8008,N_8360);
and U14600 (N_14600,N_9066,N_6166);
or U14601 (N_14601,N_7319,N_9681);
or U14602 (N_14602,N_5661,N_5566);
nor U14603 (N_14603,N_6551,N_8569);
nand U14604 (N_14604,N_6284,N_5491);
nand U14605 (N_14605,N_8779,N_5716);
nor U14606 (N_14606,N_9670,N_5115);
xor U14607 (N_14607,N_9250,N_5375);
nand U14608 (N_14608,N_8259,N_5672);
nand U14609 (N_14609,N_8703,N_7402);
nor U14610 (N_14610,N_7850,N_8613);
or U14611 (N_14611,N_7073,N_9237);
nand U14612 (N_14612,N_8925,N_8842);
or U14613 (N_14613,N_5415,N_6518);
or U14614 (N_14614,N_5223,N_5342);
or U14615 (N_14615,N_7628,N_6643);
nand U14616 (N_14616,N_5324,N_7003);
nand U14617 (N_14617,N_5302,N_6493);
nor U14618 (N_14618,N_9432,N_7720);
or U14619 (N_14619,N_5070,N_5990);
and U14620 (N_14620,N_7867,N_7068);
or U14621 (N_14621,N_6256,N_8065);
or U14622 (N_14622,N_9826,N_8245);
nor U14623 (N_14623,N_5197,N_9450);
nor U14624 (N_14624,N_9698,N_5839);
xor U14625 (N_14625,N_6164,N_7993);
nand U14626 (N_14626,N_7361,N_7296);
or U14627 (N_14627,N_9311,N_8905);
or U14628 (N_14628,N_6117,N_7616);
nand U14629 (N_14629,N_5213,N_8095);
and U14630 (N_14630,N_8382,N_6793);
or U14631 (N_14631,N_8126,N_7400);
nand U14632 (N_14632,N_6913,N_5298);
or U14633 (N_14633,N_7927,N_8398);
nor U14634 (N_14634,N_6300,N_6150);
nor U14635 (N_14635,N_5299,N_5407);
or U14636 (N_14636,N_5932,N_5234);
nand U14637 (N_14637,N_8359,N_5461);
xor U14638 (N_14638,N_7049,N_7107);
and U14639 (N_14639,N_6807,N_7673);
nor U14640 (N_14640,N_7202,N_9588);
nand U14641 (N_14641,N_6627,N_9325);
nand U14642 (N_14642,N_8918,N_5980);
xor U14643 (N_14643,N_5225,N_9385);
or U14644 (N_14644,N_6932,N_9625);
nand U14645 (N_14645,N_6571,N_6842);
and U14646 (N_14646,N_7221,N_5714);
nor U14647 (N_14647,N_7677,N_6328);
nand U14648 (N_14648,N_9267,N_7970);
and U14649 (N_14649,N_5260,N_6213);
or U14650 (N_14650,N_6013,N_6649);
nand U14651 (N_14651,N_8258,N_6946);
or U14652 (N_14652,N_5044,N_9592);
xor U14653 (N_14653,N_8559,N_6544);
nand U14654 (N_14654,N_5189,N_8355);
nor U14655 (N_14655,N_9411,N_7269);
or U14656 (N_14656,N_8948,N_5312);
and U14657 (N_14657,N_9899,N_8477);
nor U14658 (N_14658,N_7920,N_5025);
nand U14659 (N_14659,N_9675,N_6362);
xor U14660 (N_14660,N_9143,N_5834);
or U14661 (N_14661,N_9421,N_8943);
nor U14662 (N_14662,N_7041,N_7215);
or U14663 (N_14663,N_6845,N_8856);
and U14664 (N_14664,N_9597,N_7439);
and U14665 (N_14665,N_9717,N_7032);
nor U14666 (N_14666,N_6754,N_8326);
or U14667 (N_14667,N_7886,N_7186);
nand U14668 (N_14668,N_9319,N_9525);
nand U14669 (N_14669,N_7668,N_5548);
or U14670 (N_14670,N_6045,N_8434);
and U14671 (N_14671,N_7307,N_7535);
xnor U14672 (N_14672,N_8496,N_9389);
and U14673 (N_14673,N_7547,N_5555);
and U14674 (N_14674,N_5826,N_5578);
and U14675 (N_14675,N_9478,N_6239);
nand U14676 (N_14676,N_8344,N_9032);
xnor U14677 (N_14677,N_9944,N_9360);
nor U14678 (N_14678,N_6370,N_8555);
nand U14679 (N_14679,N_6679,N_9586);
and U14680 (N_14680,N_5321,N_7465);
nand U14681 (N_14681,N_7700,N_5926);
or U14682 (N_14682,N_6080,N_8518);
and U14683 (N_14683,N_7244,N_8279);
nand U14684 (N_14684,N_9636,N_7576);
and U14685 (N_14685,N_5492,N_5841);
xnor U14686 (N_14686,N_8266,N_5569);
nor U14687 (N_14687,N_8118,N_9283);
or U14688 (N_14688,N_5649,N_9001);
or U14689 (N_14689,N_6978,N_7531);
or U14690 (N_14690,N_5158,N_7763);
and U14691 (N_14691,N_6345,N_6688);
or U14692 (N_14692,N_6667,N_7284);
and U14693 (N_14693,N_7886,N_9870);
nor U14694 (N_14694,N_5609,N_5292);
or U14695 (N_14695,N_7296,N_8498);
or U14696 (N_14696,N_7940,N_7588);
or U14697 (N_14697,N_7034,N_6097);
xnor U14698 (N_14698,N_5290,N_9919);
nand U14699 (N_14699,N_9537,N_6376);
nor U14700 (N_14700,N_9509,N_8211);
xnor U14701 (N_14701,N_9502,N_7555);
nand U14702 (N_14702,N_9126,N_7383);
and U14703 (N_14703,N_6239,N_5827);
nand U14704 (N_14704,N_7518,N_8522);
and U14705 (N_14705,N_8765,N_6345);
nand U14706 (N_14706,N_8052,N_8458);
nand U14707 (N_14707,N_5039,N_9801);
nor U14708 (N_14708,N_7834,N_9041);
xnor U14709 (N_14709,N_9177,N_6700);
nand U14710 (N_14710,N_7096,N_8692);
or U14711 (N_14711,N_6955,N_7268);
nand U14712 (N_14712,N_8525,N_7127);
or U14713 (N_14713,N_8140,N_5875);
xor U14714 (N_14714,N_6064,N_6684);
nand U14715 (N_14715,N_5825,N_8231);
nand U14716 (N_14716,N_9887,N_9890);
or U14717 (N_14717,N_6389,N_5114);
nor U14718 (N_14718,N_7045,N_9346);
xor U14719 (N_14719,N_6211,N_5324);
or U14720 (N_14720,N_7928,N_7930);
nand U14721 (N_14721,N_6699,N_9972);
nand U14722 (N_14722,N_7394,N_6921);
or U14723 (N_14723,N_6926,N_5999);
xnor U14724 (N_14724,N_6400,N_7150);
nand U14725 (N_14725,N_7089,N_9004);
and U14726 (N_14726,N_5783,N_6512);
and U14727 (N_14727,N_5228,N_9459);
and U14728 (N_14728,N_6270,N_7296);
or U14729 (N_14729,N_8306,N_7286);
xor U14730 (N_14730,N_7800,N_7518);
and U14731 (N_14731,N_6122,N_6685);
nand U14732 (N_14732,N_5013,N_7060);
and U14733 (N_14733,N_5274,N_8509);
nand U14734 (N_14734,N_9519,N_9218);
and U14735 (N_14735,N_5649,N_9401);
nand U14736 (N_14736,N_7323,N_6743);
xnor U14737 (N_14737,N_7603,N_9483);
nand U14738 (N_14738,N_5458,N_8939);
or U14739 (N_14739,N_8921,N_8524);
nor U14740 (N_14740,N_7037,N_8426);
nand U14741 (N_14741,N_7192,N_7988);
nand U14742 (N_14742,N_6688,N_9355);
or U14743 (N_14743,N_6176,N_6173);
xor U14744 (N_14744,N_9301,N_7108);
or U14745 (N_14745,N_6877,N_9396);
or U14746 (N_14746,N_7414,N_6596);
nand U14747 (N_14747,N_9062,N_8969);
or U14748 (N_14748,N_6971,N_7149);
nor U14749 (N_14749,N_5974,N_8390);
and U14750 (N_14750,N_9611,N_7354);
or U14751 (N_14751,N_8608,N_9579);
nand U14752 (N_14752,N_7490,N_7271);
xor U14753 (N_14753,N_8605,N_9778);
xor U14754 (N_14754,N_7777,N_5884);
xor U14755 (N_14755,N_9789,N_9580);
xor U14756 (N_14756,N_7327,N_8177);
xnor U14757 (N_14757,N_9235,N_9138);
xor U14758 (N_14758,N_5810,N_9090);
nand U14759 (N_14759,N_5739,N_6226);
nand U14760 (N_14760,N_8094,N_5950);
nand U14761 (N_14761,N_7932,N_8282);
xor U14762 (N_14762,N_6183,N_7952);
or U14763 (N_14763,N_8086,N_7943);
nor U14764 (N_14764,N_5251,N_5133);
nand U14765 (N_14765,N_6653,N_5387);
and U14766 (N_14766,N_9712,N_5247);
nand U14767 (N_14767,N_9616,N_8413);
nor U14768 (N_14768,N_8588,N_5436);
xnor U14769 (N_14769,N_6978,N_9593);
and U14770 (N_14770,N_7867,N_7556);
and U14771 (N_14771,N_5344,N_7907);
xnor U14772 (N_14772,N_9757,N_6025);
nor U14773 (N_14773,N_5570,N_9663);
nand U14774 (N_14774,N_6208,N_5472);
nand U14775 (N_14775,N_6135,N_8438);
xnor U14776 (N_14776,N_6210,N_5564);
and U14777 (N_14777,N_9958,N_9587);
nand U14778 (N_14778,N_8806,N_6274);
and U14779 (N_14779,N_5747,N_9467);
nand U14780 (N_14780,N_5918,N_9517);
nor U14781 (N_14781,N_7548,N_9531);
and U14782 (N_14782,N_5924,N_5742);
or U14783 (N_14783,N_8677,N_9892);
nand U14784 (N_14784,N_7108,N_9018);
xor U14785 (N_14785,N_5650,N_5378);
or U14786 (N_14786,N_7087,N_8904);
nor U14787 (N_14787,N_5510,N_7426);
nand U14788 (N_14788,N_7485,N_5233);
nand U14789 (N_14789,N_6721,N_9356);
nor U14790 (N_14790,N_5293,N_9439);
xnor U14791 (N_14791,N_6499,N_9020);
nor U14792 (N_14792,N_8767,N_6923);
xnor U14793 (N_14793,N_6301,N_9049);
nand U14794 (N_14794,N_7744,N_6312);
nor U14795 (N_14795,N_9916,N_7034);
xnor U14796 (N_14796,N_8645,N_6839);
xnor U14797 (N_14797,N_9268,N_6218);
and U14798 (N_14798,N_6078,N_5012);
and U14799 (N_14799,N_5399,N_9312);
nand U14800 (N_14800,N_6130,N_6807);
nor U14801 (N_14801,N_5211,N_5345);
xor U14802 (N_14802,N_6389,N_6547);
or U14803 (N_14803,N_6637,N_7412);
nand U14804 (N_14804,N_5486,N_5681);
and U14805 (N_14805,N_9741,N_7542);
xnor U14806 (N_14806,N_6038,N_7232);
and U14807 (N_14807,N_7642,N_5392);
nand U14808 (N_14808,N_5527,N_5226);
nor U14809 (N_14809,N_6115,N_8814);
and U14810 (N_14810,N_6095,N_7677);
nand U14811 (N_14811,N_8323,N_5224);
or U14812 (N_14812,N_5471,N_9984);
and U14813 (N_14813,N_8400,N_7106);
nor U14814 (N_14814,N_9441,N_8696);
and U14815 (N_14815,N_9058,N_7957);
and U14816 (N_14816,N_9859,N_8305);
or U14817 (N_14817,N_5259,N_5688);
nor U14818 (N_14818,N_8695,N_7456);
or U14819 (N_14819,N_6003,N_6252);
nand U14820 (N_14820,N_7680,N_9711);
or U14821 (N_14821,N_9636,N_9253);
xor U14822 (N_14822,N_9497,N_9314);
nor U14823 (N_14823,N_8636,N_5848);
nor U14824 (N_14824,N_5806,N_5798);
or U14825 (N_14825,N_5825,N_5430);
xor U14826 (N_14826,N_5602,N_5256);
nand U14827 (N_14827,N_6497,N_5080);
nand U14828 (N_14828,N_7117,N_9369);
or U14829 (N_14829,N_6073,N_7481);
xor U14830 (N_14830,N_8632,N_6038);
or U14831 (N_14831,N_5125,N_5486);
or U14832 (N_14832,N_6539,N_9595);
nand U14833 (N_14833,N_6147,N_5983);
and U14834 (N_14834,N_7498,N_8926);
or U14835 (N_14835,N_6722,N_5165);
xnor U14836 (N_14836,N_5122,N_7210);
or U14837 (N_14837,N_9420,N_7290);
xnor U14838 (N_14838,N_8450,N_8267);
xor U14839 (N_14839,N_9442,N_6967);
nor U14840 (N_14840,N_7218,N_9262);
xnor U14841 (N_14841,N_5165,N_5807);
xor U14842 (N_14842,N_6001,N_7569);
and U14843 (N_14843,N_5365,N_5058);
or U14844 (N_14844,N_8938,N_7557);
or U14845 (N_14845,N_5999,N_8447);
nor U14846 (N_14846,N_9660,N_6527);
xor U14847 (N_14847,N_7102,N_9689);
nand U14848 (N_14848,N_5936,N_9628);
nand U14849 (N_14849,N_9316,N_8699);
or U14850 (N_14850,N_7628,N_9776);
nor U14851 (N_14851,N_5555,N_6571);
xor U14852 (N_14852,N_8083,N_7160);
nand U14853 (N_14853,N_6046,N_7527);
or U14854 (N_14854,N_8191,N_6723);
xnor U14855 (N_14855,N_7697,N_7931);
xnor U14856 (N_14856,N_8404,N_6264);
and U14857 (N_14857,N_7461,N_7600);
and U14858 (N_14858,N_5077,N_6781);
nor U14859 (N_14859,N_5631,N_6356);
and U14860 (N_14860,N_5530,N_8907);
nor U14861 (N_14861,N_8492,N_6324);
xor U14862 (N_14862,N_8989,N_7714);
nor U14863 (N_14863,N_5384,N_8487);
or U14864 (N_14864,N_8972,N_5809);
and U14865 (N_14865,N_9426,N_8370);
nand U14866 (N_14866,N_8083,N_9501);
and U14867 (N_14867,N_8205,N_7229);
nor U14868 (N_14868,N_9562,N_6858);
nand U14869 (N_14869,N_7703,N_7597);
nand U14870 (N_14870,N_5653,N_7642);
xnor U14871 (N_14871,N_5271,N_6488);
and U14872 (N_14872,N_9542,N_9083);
nor U14873 (N_14873,N_8911,N_6147);
xor U14874 (N_14874,N_6468,N_8193);
or U14875 (N_14875,N_9094,N_6659);
xor U14876 (N_14876,N_7559,N_9396);
nor U14877 (N_14877,N_5116,N_7646);
nand U14878 (N_14878,N_8636,N_5839);
xnor U14879 (N_14879,N_5281,N_5057);
xor U14880 (N_14880,N_7714,N_5897);
or U14881 (N_14881,N_9933,N_9433);
nand U14882 (N_14882,N_9464,N_7257);
and U14883 (N_14883,N_6603,N_9891);
nor U14884 (N_14884,N_9287,N_6122);
and U14885 (N_14885,N_8701,N_5943);
xnor U14886 (N_14886,N_7263,N_8020);
xnor U14887 (N_14887,N_6575,N_5183);
and U14888 (N_14888,N_8214,N_9246);
nand U14889 (N_14889,N_5625,N_7358);
or U14890 (N_14890,N_6637,N_5681);
and U14891 (N_14891,N_7951,N_5693);
xnor U14892 (N_14892,N_7596,N_8821);
nand U14893 (N_14893,N_8691,N_7308);
or U14894 (N_14894,N_5555,N_7092);
and U14895 (N_14895,N_8536,N_5114);
nand U14896 (N_14896,N_7893,N_6557);
nor U14897 (N_14897,N_9631,N_8404);
and U14898 (N_14898,N_7110,N_8244);
and U14899 (N_14899,N_8196,N_9651);
and U14900 (N_14900,N_9341,N_5912);
xor U14901 (N_14901,N_5852,N_6574);
nor U14902 (N_14902,N_6039,N_6208);
nor U14903 (N_14903,N_7594,N_8050);
or U14904 (N_14904,N_6704,N_7634);
nand U14905 (N_14905,N_6235,N_8910);
and U14906 (N_14906,N_7826,N_9792);
nand U14907 (N_14907,N_7471,N_7734);
or U14908 (N_14908,N_5182,N_6223);
nand U14909 (N_14909,N_5994,N_9680);
nand U14910 (N_14910,N_7327,N_8703);
nor U14911 (N_14911,N_7123,N_5483);
nor U14912 (N_14912,N_5829,N_7235);
nand U14913 (N_14913,N_6992,N_9870);
and U14914 (N_14914,N_5256,N_7174);
nand U14915 (N_14915,N_7129,N_9424);
or U14916 (N_14916,N_6375,N_5544);
nand U14917 (N_14917,N_7534,N_5480);
xor U14918 (N_14918,N_7755,N_8022);
nor U14919 (N_14919,N_7672,N_5775);
or U14920 (N_14920,N_6408,N_8999);
nor U14921 (N_14921,N_9417,N_6678);
and U14922 (N_14922,N_5808,N_5618);
and U14923 (N_14923,N_9907,N_6001);
or U14924 (N_14924,N_7199,N_5852);
or U14925 (N_14925,N_8087,N_8983);
xor U14926 (N_14926,N_6287,N_9620);
xor U14927 (N_14927,N_9220,N_9038);
nor U14928 (N_14928,N_5334,N_9475);
nand U14929 (N_14929,N_5085,N_7330);
nor U14930 (N_14930,N_7904,N_8537);
or U14931 (N_14931,N_6031,N_7667);
or U14932 (N_14932,N_6408,N_6977);
nand U14933 (N_14933,N_5972,N_8799);
nor U14934 (N_14934,N_6074,N_5234);
or U14935 (N_14935,N_6922,N_6115);
nor U14936 (N_14936,N_9223,N_8060);
nor U14937 (N_14937,N_8208,N_8558);
xor U14938 (N_14938,N_5383,N_5417);
nand U14939 (N_14939,N_8837,N_9283);
and U14940 (N_14940,N_8982,N_9040);
xor U14941 (N_14941,N_7866,N_8225);
or U14942 (N_14942,N_5313,N_8483);
xor U14943 (N_14943,N_9710,N_5662);
and U14944 (N_14944,N_9872,N_5140);
and U14945 (N_14945,N_5624,N_6636);
or U14946 (N_14946,N_6131,N_6024);
xnor U14947 (N_14947,N_6369,N_9159);
nor U14948 (N_14948,N_9419,N_6620);
nand U14949 (N_14949,N_9661,N_6722);
xnor U14950 (N_14950,N_9082,N_9676);
or U14951 (N_14951,N_7707,N_6986);
and U14952 (N_14952,N_5623,N_6718);
nor U14953 (N_14953,N_9172,N_8377);
or U14954 (N_14954,N_9801,N_6923);
nor U14955 (N_14955,N_8356,N_7321);
nor U14956 (N_14956,N_5798,N_6313);
nand U14957 (N_14957,N_9004,N_7616);
or U14958 (N_14958,N_5809,N_7152);
nor U14959 (N_14959,N_9402,N_6632);
and U14960 (N_14960,N_5090,N_8470);
nand U14961 (N_14961,N_8711,N_6571);
nor U14962 (N_14962,N_7120,N_5232);
nor U14963 (N_14963,N_5368,N_5633);
nor U14964 (N_14964,N_8825,N_7255);
and U14965 (N_14965,N_5830,N_7087);
nand U14966 (N_14966,N_7151,N_5444);
and U14967 (N_14967,N_6124,N_9279);
nand U14968 (N_14968,N_8370,N_6372);
nand U14969 (N_14969,N_5870,N_7200);
xor U14970 (N_14970,N_7637,N_6391);
or U14971 (N_14971,N_8527,N_6542);
or U14972 (N_14972,N_7974,N_5204);
nand U14973 (N_14973,N_6888,N_6435);
nand U14974 (N_14974,N_8543,N_6516);
and U14975 (N_14975,N_7581,N_9607);
nor U14976 (N_14976,N_9252,N_9602);
xnor U14977 (N_14977,N_6760,N_8402);
or U14978 (N_14978,N_9515,N_9745);
nor U14979 (N_14979,N_8724,N_9506);
or U14980 (N_14980,N_6625,N_9312);
or U14981 (N_14981,N_5723,N_6764);
and U14982 (N_14982,N_9572,N_7546);
nand U14983 (N_14983,N_9796,N_6967);
or U14984 (N_14984,N_7544,N_8613);
nor U14985 (N_14985,N_5824,N_5057);
nor U14986 (N_14986,N_8268,N_9542);
nand U14987 (N_14987,N_9814,N_6425);
and U14988 (N_14988,N_6809,N_6296);
nor U14989 (N_14989,N_9860,N_5276);
or U14990 (N_14990,N_5430,N_5515);
and U14991 (N_14991,N_9713,N_8665);
nand U14992 (N_14992,N_6258,N_7747);
and U14993 (N_14993,N_6468,N_6661);
or U14994 (N_14994,N_5916,N_9235);
nand U14995 (N_14995,N_5355,N_9840);
xnor U14996 (N_14996,N_9942,N_6067);
xor U14997 (N_14997,N_9020,N_6970);
xnor U14998 (N_14998,N_5669,N_5673);
xnor U14999 (N_14999,N_5820,N_8226);
xor U15000 (N_15000,N_12850,N_11571);
or U15001 (N_15001,N_14488,N_12916);
and U15002 (N_15002,N_11092,N_13829);
nand U15003 (N_15003,N_14427,N_13366);
and U15004 (N_15004,N_12600,N_12782);
xor U15005 (N_15005,N_12460,N_10758);
nor U15006 (N_15006,N_10257,N_10963);
nor U15007 (N_15007,N_13276,N_14922);
nand U15008 (N_15008,N_12308,N_13541);
nand U15009 (N_15009,N_13217,N_14813);
xor U15010 (N_15010,N_12266,N_14859);
xor U15011 (N_15011,N_12406,N_10958);
nor U15012 (N_15012,N_11300,N_14617);
nor U15013 (N_15013,N_12310,N_12121);
nand U15014 (N_15014,N_13216,N_10846);
and U15015 (N_15015,N_14993,N_14847);
nor U15016 (N_15016,N_13860,N_12980);
nand U15017 (N_15017,N_14274,N_11792);
and U15018 (N_15018,N_13979,N_13658);
nand U15019 (N_15019,N_12612,N_11918);
and U15020 (N_15020,N_10155,N_13258);
nand U15021 (N_15021,N_12968,N_10240);
xnor U15022 (N_15022,N_11278,N_12190);
and U15023 (N_15023,N_13213,N_10157);
xor U15024 (N_15024,N_11117,N_10483);
nor U15025 (N_15025,N_10364,N_11177);
xor U15026 (N_15026,N_14067,N_11132);
xnor U15027 (N_15027,N_12154,N_13299);
and U15028 (N_15028,N_12469,N_11405);
xnor U15029 (N_15029,N_11106,N_14374);
nand U15030 (N_15030,N_14304,N_12162);
or U15031 (N_15031,N_12885,N_12050);
nor U15032 (N_15032,N_13794,N_11983);
nand U15033 (N_15033,N_10278,N_10225);
xor U15034 (N_15034,N_12854,N_14283);
or U15035 (N_15035,N_13898,N_12407);
and U15036 (N_15036,N_13520,N_14347);
and U15037 (N_15037,N_11305,N_10287);
xnor U15038 (N_15038,N_14610,N_13825);
xor U15039 (N_15039,N_13219,N_14723);
nor U15040 (N_15040,N_12151,N_14215);
or U15041 (N_15041,N_12393,N_10368);
and U15042 (N_15042,N_11167,N_14756);
nor U15043 (N_15043,N_10588,N_12258);
nor U15044 (N_15044,N_13273,N_12982);
and U15045 (N_15045,N_12205,N_14360);
and U15046 (N_15046,N_13716,N_13082);
nand U15047 (N_15047,N_12478,N_11265);
nand U15048 (N_15048,N_12092,N_11270);
and U15049 (N_15049,N_11394,N_14064);
nor U15050 (N_15050,N_11052,N_13813);
xor U15051 (N_15051,N_11023,N_14117);
and U15052 (N_15052,N_14528,N_13667);
xnor U15053 (N_15053,N_11842,N_12536);
and U15054 (N_15054,N_12135,N_10150);
nor U15055 (N_15055,N_10297,N_12865);
xnor U15056 (N_15056,N_10980,N_13095);
nor U15057 (N_15057,N_14025,N_11252);
or U15058 (N_15058,N_10977,N_14870);
xnor U15059 (N_15059,N_13048,N_14997);
xnor U15060 (N_15060,N_12119,N_14907);
and U15061 (N_15061,N_14709,N_11097);
nand U15062 (N_15062,N_11328,N_11745);
and U15063 (N_15063,N_12966,N_12963);
or U15064 (N_15064,N_14371,N_13274);
or U15065 (N_15065,N_13339,N_10581);
or U15066 (N_15066,N_10123,N_10578);
nand U15067 (N_15067,N_12847,N_12664);
nand U15068 (N_15068,N_11743,N_14494);
and U15069 (N_15069,N_12087,N_10487);
nand U15070 (N_15070,N_12260,N_12335);
nor U15071 (N_15071,N_14110,N_12957);
or U15072 (N_15072,N_10622,N_12570);
nand U15073 (N_15073,N_14896,N_14812);
nand U15074 (N_15074,N_11088,N_10815);
xor U15075 (N_15075,N_11863,N_14683);
or U15076 (N_15076,N_12530,N_14231);
nand U15077 (N_15077,N_12811,N_12663);
nand U15078 (N_15078,N_12036,N_14157);
xor U15079 (N_15079,N_12419,N_11469);
nor U15080 (N_15080,N_11815,N_12784);
xor U15081 (N_15081,N_14111,N_13348);
or U15082 (N_15082,N_14971,N_13915);
xnor U15083 (N_15083,N_10825,N_12483);
nand U15084 (N_15084,N_11374,N_11478);
xor U15085 (N_15085,N_11967,N_10139);
nor U15086 (N_15086,N_10677,N_14841);
or U15087 (N_15087,N_12384,N_12629);
and U15088 (N_15088,N_14006,N_10989);
and U15089 (N_15089,N_13368,N_10300);
nand U15090 (N_15090,N_10058,N_12449);
nor U15091 (N_15091,N_14832,N_10057);
nand U15092 (N_15092,N_12007,N_11690);
nor U15093 (N_15093,N_10724,N_10370);
and U15094 (N_15094,N_11181,N_10356);
xnor U15095 (N_15095,N_14702,N_11636);
xor U15096 (N_15096,N_12696,N_12858);
or U15097 (N_15097,N_10496,N_10263);
xor U15098 (N_15098,N_12262,N_11003);
nand U15099 (N_15099,N_14513,N_10988);
or U15100 (N_15100,N_11507,N_10735);
and U15101 (N_15101,N_12311,N_13247);
nor U15102 (N_15102,N_12741,N_13579);
nor U15103 (N_15103,N_14718,N_13812);
and U15104 (N_15104,N_10498,N_13014);
nand U15105 (N_15105,N_13557,N_12021);
xor U15106 (N_15106,N_11018,N_13294);
xor U15107 (N_15107,N_11190,N_13266);
xor U15108 (N_15108,N_14563,N_14018);
nand U15109 (N_15109,N_11198,N_13789);
or U15110 (N_15110,N_12585,N_10961);
nand U15111 (N_15111,N_10252,N_14102);
and U15112 (N_15112,N_13868,N_12099);
xnor U15113 (N_15113,N_13469,N_14155);
and U15114 (N_15114,N_13859,N_13310);
nor U15115 (N_15115,N_10184,N_10290);
nor U15116 (N_15116,N_12548,N_13561);
xnor U15117 (N_15117,N_14092,N_14272);
or U15118 (N_15118,N_14009,N_12947);
nand U15119 (N_15119,N_11620,N_11799);
nor U15120 (N_15120,N_12773,N_12690);
xor U15121 (N_15121,N_10407,N_11931);
or U15122 (N_15122,N_11233,N_11896);
or U15123 (N_15123,N_13050,N_14378);
or U15124 (N_15124,N_14176,N_14988);
nand U15125 (N_15125,N_13827,N_14763);
nor U15126 (N_15126,N_10933,N_11050);
xor U15127 (N_15127,N_10379,N_13526);
xor U15128 (N_15128,N_14869,N_12654);
xor U15129 (N_15129,N_10066,N_11515);
and U15130 (N_15130,N_10227,N_10213);
nand U15131 (N_15131,N_12497,N_13023);
or U15132 (N_15132,N_11149,N_13575);
nand U15133 (N_15133,N_11325,N_12286);
or U15134 (N_15134,N_14071,N_14467);
and U15135 (N_15135,N_11686,N_13865);
and U15136 (N_15136,N_12875,N_13096);
or U15137 (N_15137,N_12775,N_10171);
and U15138 (N_15138,N_11638,N_14086);
and U15139 (N_15139,N_11361,N_11975);
xnor U15140 (N_15140,N_13834,N_10342);
xor U15141 (N_15141,N_12821,N_11037);
nand U15142 (N_15142,N_13307,N_10995);
xor U15143 (N_15143,N_13650,N_11007);
and U15144 (N_15144,N_10306,N_12757);
and U15145 (N_15145,N_10937,N_11164);
and U15146 (N_15146,N_11669,N_11200);
xnor U15147 (N_15147,N_10755,N_13199);
or U15148 (N_15148,N_11929,N_13434);
nand U15149 (N_15149,N_12026,N_10733);
and U15150 (N_15150,N_10160,N_14320);
nand U15151 (N_15151,N_13830,N_12785);
or U15152 (N_15152,N_10595,N_11191);
xnor U15153 (N_15153,N_13560,N_12411);
xnor U15154 (N_15154,N_14555,N_12048);
nand U15155 (N_15155,N_14539,N_13828);
nor U15156 (N_15156,N_11939,N_13704);
nand U15157 (N_15157,N_10305,N_12823);
nand U15158 (N_15158,N_14823,N_11676);
xor U15159 (N_15159,N_14357,N_12013);
nand U15160 (N_15160,N_11295,N_12900);
xnor U15161 (N_15161,N_14962,N_11528);
nand U15162 (N_15162,N_12032,N_10628);
and U15163 (N_15163,N_13964,N_10143);
or U15164 (N_15164,N_10585,N_10999);
nor U15165 (N_15165,N_10475,N_12242);
nand U15166 (N_15166,N_13137,N_13395);
nor U15167 (N_15167,N_10237,N_10249);
and U15168 (N_15168,N_12978,N_11470);
nor U15169 (N_15169,N_13823,N_12630);
xnor U15170 (N_15170,N_12115,N_14692);
nand U15171 (N_15171,N_14126,N_14259);
nand U15172 (N_15172,N_11214,N_14850);
nor U15173 (N_15173,N_13479,N_11483);
and U15174 (N_15174,N_14490,N_14878);
and U15175 (N_15175,N_11958,N_12710);
and U15176 (N_15176,N_12147,N_13343);
nand U15177 (N_15177,N_13694,N_14161);
or U15178 (N_15178,N_13383,N_11310);
or U15179 (N_15179,N_14738,N_11093);
xnor U15180 (N_15180,N_11701,N_13935);
nand U15181 (N_15181,N_10486,N_11986);
xnor U15182 (N_15182,N_14815,N_11402);
nand U15183 (N_15183,N_13091,N_12694);
xor U15184 (N_15184,N_12088,N_10369);
xor U15185 (N_15185,N_11979,N_12257);
nor U15186 (N_15186,N_13897,N_11488);
or U15187 (N_15187,N_12314,N_11642);
or U15188 (N_15188,N_10871,N_11059);
xor U15189 (N_15189,N_10930,N_13452);
nor U15190 (N_15190,N_11869,N_13300);
nand U15191 (N_15191,N_10216,N_11185);
nor U15192 (N_15192,N_12336,N_10389);
nor U15193 (N_15193,N_10120,N_11639);
or U15194 (N_15194,N_10304,N_12891);
nand U15195 (N_15195,N_13461,N_12467);
nor U15196 (N_15196,N_10783,N_13278);
xnor U15197 (N_15197,N_14674,N_11268);
or U15198 (N_15198,N_13249,N_13421);
xnor U15199 (N_15199,N_11928,N_14710);
xor U15200 (N_15200,N_10878,N_11158);
nor U15201 (N_15201,N_12108,N_13358);
nor U15202 (N_15202,N_11276,N_12474);
xnor U15203 (N_15203,N_12707,N_13167);
nor U15204 (N_15204,N_10981,N_14687);
and U15205 (N_15205,N_10466,N_13530);
nor U15206 (N_15206,N_12194,N_13745);
nor U15207 (N_15207,N_12501,N_14915);
nand U15208 (N_15208,N_13040,N_13934);
nand U15209 (N_15209,N_10042,N_13907);
nor U15210 (N_15210,N_10763,N_13811);
or U15211 (N_15211,N_14821,N_14376);
xor U15212 (N_15212,N_11242,N_11903);
or U15213 (N_15213,N_11299,N_12913);
and U15214 (N_15214,N_12876,N_13911);
or U15215 (N_15215,N_11830,N_14422);
nand U15216 (N_15216,N_14305,N_13995);
or U15217 (N_15217,N_11419,N_12320);
and U15218 (N_15218,N_13439,N_12528);
or U15219 (N_15219,N_13548,N_10422);
xor U15220 (N_15220,N_13544,N_13196);
or U15221 (N_15221,N_14974,N_14854);
nand U15222 (N_15222,N_12835,N_10797);
or U15223 (N_15223,N_13097,N_12187);
and U15224 (N_15224,N_12104,N_12722);
nor U15225 (N_15225,N_14392,N_10310);
or U15226 (N_15226,N_10746,N_12273);
nor U15227 (N_15227,N_11897,N_12296);
nand U15228 (N_15228,N_14062,N_10457);
nand U15229 (N_15229,N_12074,N_14146);
nor U15230 (N_15230,N_10365,N_14010);
nand U15231 (N_15231,N_13718,N_10997);
nand U15232 (N_15232,N_11645,N_13563);
nand U15233 (N_15233,N_13426,N_14496);
or U15234 (N_15234,N_13886,N_10134);
or U15235 (N_15235,N_13737,N_13677);
xnor U15236 (N_15236,N_14606,N_10720);
and U15237 (N_15237,N_13204,N_11540);
nor U15238 (N_15238,N_12290,N_12085);
and U15239 (N_15239,N_10118,N_14678);
nor U15240 (N_15240,N_13736,N_10083);
and U15241 (N_15241,N_11518,N_11513);
nand U15242 (N_15242,N_12921,N_14000);
xnor U15243 (N_15243,N_14767,N_13618);
and U15244 (N_15244,N_13275,N_11882);
and U15245 (N_15245,N_14943,N_10072);
xnor U15246 (N_15246,N_10488,N_13078);
or U15247 (N_15247,N_12987,N_10831);
or U15248 (N_15248,N_14391,N_14120);
nand U15249 (N_15249,N_11788,N_12889);
xor U15250 (N_15250,N_12636,N_13448);
xor U15251 (N_15251,N_10653,N_12948);
and U15252 (N_15252,N_11294,N_11022);
nand U15253 (N_15253,N_11562,N_14151);
nand U15254 (N_15254,N_14397,N_12562);
nand U15255 (N_15255,N_14039,N_11921);
xor U15256 (N_15256,N_11121,N_12477);
or U15257 (N_15257,N_14594,N_10807);
and U15258 (N_15258,N_13245,N_12874);
and U15259 (N_15259,N_10111,N_10392);
xor U15260 (N_15260,N_14226,N_11077);
nor U15261 (N_15261,N_11737,N_14044);
nor U15262 (N_15262,N_14852,N_11703);
xor U15263 (N_15263,N_13500,N_11110);
and U15264 (N_15264,N_13387,N_14957);
xor U15265 (N_15265,N_11395,N_11641);
or U15266 (N_15266,N_10556,N_13115);
or U15267 (N_15267,N_11692,N_10378);
nand U15268 (N_15268,N_11917,N_10561);
nand U15269 (N_15269,N_11687,N_14354);
or U15270 (N_15270,N_11100,N_14860);
nand U15271 (N_15271,N_10013,N_12575);
xor U15272 (N_15272,N_10241,N_12880);
xor U15273 (N_15273,N_12898,N_12372);
nand U15274 (N_15274,N_14779,N_14370);
and U15275 (N_15275,N_13382,N_13547);
and U15276 (N_15276,N_14216,N_10312);
nand U15277 (N_15277,N_11234,N_14441);
xor U15278 (N_15278,N_11187,N_11152);
or U15279 (N_15279,N_14826,N_13011);
or U15280 (N_15280,N_10405,N_13003);
and U15281 (N_15281,N_10253,N_14855);
xor U15282 (N_15282,N_13021,N_10991);
and U15283 (N_15283,N_14797,N_12596);
and U15284 (N_15284,N_14138,N_13151);
and U15285 (N_15285,N_10008,N_13488);
nand U15286 (N_15286,N_11752,N_12264);
or U15287 (N_15287,N_13427,N_13616);
xnor U15288 (N_15288,N_10520,N_14569);
or U15289 (N_15289,N_14578,N_10149);
xor U15290 (N_15290,N_13960,N_12339);
nor U15291 (N_15291,N_11162,N_11914);
and U15292 (N_15292,N_10215,N_11750);
and U15293 (N_15293,N_10102,N_12992);
and U15294 (N_15294,N_12798,N_13337);
nand U15295 (N_15295,N_12186,N_14352);
and U15296 (N_15296,N_10456,N_14950);
xnor U15297 (N_15297,N_13729,N_10440);
nor U15298 (N_15298,N_10446,N_11410);
nor U15299 (N_15299,N_10404,N_14275);
nand U15300 (N_15300,N_12917,N_13946);
or U15301 (N_15301,N_10881,N_12441);
xnor U15302 (N_15302,N_12044,N_10395);
nor U15303 (N_15303,N_10776,N_11220);
xor U15304 (N_15304,N_13218,N_13491);
or U15305 (N_15305,N_12576,N_13558);
xor U15306 (N_15306,N_11377,N_12328);
xnor U15307 (N_15307,N_11780,N_12253);
nand U15308 (N_15308,N_10564,N_10490);
nor U15309 (N_15309,N_12578,N_13397);
nor U15310 (N_15310,N_10450,N_10135);
nor U15311 (N_15311,N_14287,N_11664);
nor U15312 (N_15312,N_14103,N_13759);
nand U15313 (N_15313,N_10203,N_13471);
nor U15314 (N_15314,N_13068,N_14681);
or U15315 (N_15315,N_10941,N_14114);
or U15316 (N_15316,N_10484,N_13663);
nor U15317 (N_15317,N_10584,N_13872);
xnor U15318 (N_15318,N_12373,N_14492);
nor U15319 (N_15319,N_12025,N_11487);
nand U15320 (N_15320,N_10522,N_12881);
nor U15321 (N_15321,N_12998,N_14335);
or U15322 (N_15322,N_14686,N_12820);
or U15323 (N_15323,N_13788,N_13973);
or U15324 (N_15324,N_10965,N_11738);
nand U15325 (N_15325,N_12790,N_10175);
nor U15326 (N_15326,N_14060,N_12571);
xor U15327 (N_15327,N_12816,N_12472);
nand U15328 (N_15328,N_10718,N_11679);
or U15329 (N_15329,N_13485,N_13892);
nand U15330 (N_15330,N_10550,N_10799);
nand U15331 (N_15331,N_14144,N_10231);
nor U15332 (N_15332,N_12270,N_11546);
xnor U15333 (N_15333,N_14368,N_13494);
nor U15334 (N_15334,N_12506,N_10590);
or U15335 (N_15335,N_12397,N_14790);
or U15336 (N_15336,N_13783,N_12959);
xnor U15337 (N_15337,N_13063,N_13401);
nor U15338 (N_15338,N_14145,N_11708);
or U15339 (N_15339,N_14373,N_13436);
and U15340 (N_15340,N_11083,N_13220);
nand U15341 (N_15341,N_14433,N_11659);
xnor U15342 (N_15342,N_14295,N_12346);
or U15343 (N_15343,N_11485,N_14525);
xor U15344 (N_15344,N_14551,N_11084);
and U15345 (N_15345,N_10992,N_12806);
or U15346 (N_15346,N_10750,N_10499);
or U15347 (N_15347,N_11026,N_10303);
xor U15348 (N_15348,N_10146,N_12323);
or U15349 (N_15349,N_12860,N_12042);
and U15350 (N_15350,N_10476,N_14658);
and U15351 (N_15351,N_14769,N_11250);
xor U15352 (N_15352,N_12637,N_11962);
and U15353 (N_15353,N_10766,N_14432);
or U15354 (N_15354,N_12701,N_13422);
nor U15355 (N_15355,N_11391,N_13227);
nor U15356 (N_15356,N_14233,N_11934);
xor U15357 (N_15357,N_10728,N_12661);
xor U15358 (N_15358,N_14503,N_13851);
and U15359 (N_15359,N_11860,N_13020);
nand U15360 (N_15360,N_10412,N_10398);
nand U15361 (N_15361,N_11120,N_10829);
xor U15362 (N_15362,N_14675,N_10798);
and U15363 (N_15363,N_14362,N_11396);
nor U15364 (N_15364,N_10903,N_14534);
and U15365 (N_15365,N_12867,N_10599);
xnor U15366 (N_15366,N_14065,N_12890);
nor U15367 (N_15367,N_12772,N_12139);
nor U15368 (N_15368,N_10245,N_11206);
or U15369 (N_15369,N_14237,N_11304);
nand U15370 (N_15370,N_14839,N_13836);
or U15371 (N_15371,N_10915,N_14153);
or U15372 (N_15372,N_11383,N_10777);
or U15373 (N_15373,N_10283,N_14833);
xor U15374 (N_15374,N_14246,N_10038);
nor U15375 (N_15375,N_10824,N_10608);
nor U15376 (N_15376,N_12969,N_10383);
and U15377 (N_15377,N_12148,N_11494);
xnor U15378 (N_15378,N_12836,N_14123);
or U15379 (N_15379,N_10060,N_11027);
xor U15380 (N_15380,N_14053,N_14508);
nor U15381 (N_15381,N_10692,N_14905);
or U15382 (N_15382,N_12069,N_10610);
xnor U15383 (N_15383,N_13320,N_11925);
nor U15384 (N_15384,N_11197,N_11864);
and U15385 (N_15385,N_10969,N_14256);
nor U15386 (N_15386,N_14003,N_14080);
or U15387 (N_15387,N_14139,N_10293);
xnor U15388 (N_15388,N_10337,N_14849);
xnor U15389 (N_15389,N_11854,N_13645);
and U15390 (N_15390,N_11791,N_14191);
nand U15391 (N_15391,N_11434,N_12468);
nor U15392 (N_15392,N_11603,N_12648);
xnor U15393 (N_15393,N_11086,N_12364);
nor U15394 (N_15394,N_14845,N_13521);
xor U15395 (N_15395,N_14482,N_14935);
nor U15396 (N_15396,N_13770,N_12613);
or U15397 (N_15397,N_14061,N_14520);
nor U15398 (N_15398,N_13141,N_13473);
and U15399 (N_15399,N_11408,N_13019);
nor U15400 (N_15400,N_11421,N_11898);
xnor U15401 (N_15401,N_14109,N_12776);
xor U15402 (N_15402,N_10021,N_11732);
nand U15403 (N_15403,N_14066,N_11323);
or U15404 (N_15404,N_10512,N_12639);
or U15405 (N_15405,N_12250,N_11036);
xnor U15406 (N_15406,N_10302,N_11244);
nand U15407 (N_15407,N_12893,N_12717);
nor U15408 (N_15408,N_10932,N_11298);
or U15409 (N_15409,N_10563,N_11427);
nand U15410 (N_15410,N_12408,N_13732);
and U15411 (N_15411,N_13033,N_11754);
nand U15412 (N_15412,N_11216,N_10199);
nand U15413 (N_15413,N_13027,N_10286);
nand U15414 (N_15414,N_14603,N_12944);
xor U15415 (N_15415,N_14472,N_10817);
or U15416 (N_15416,N_14616,N_10130);
xor U15417 (N_15417,N_13835,N_10922);
xnor U15418 (N_15418,N_14476,N_10918);
nand U15419 (N_15419,N_10684,N_10966);
xnor U15420 (N_15420,N_12208,N_14955);
xor U15421 (N_15421,N_11041,N_11624);
nor U15422 (N_15422,N_11071,N_12324);
or U15423 (N_15423,N_14181,N_10234);
nor U15424 (N_15424,N_10784,N_12796);
or U15425 (N_15425,N_12750,N_14761);
and U15426 (N_15426,N_13334,N_14387);
or U15427 (N_15427,N_13818,N_11834);
nand U15428 (N_15428,N_13372,N_11356);
nor U15429 (N_15429,N_11175,N_13280);
nor U15430 (N_15430,N_13924,N_13309);
xor U15431 (N_15431,N_14609,N_12923);
xnor U15432 (N_15432,N_14717,N_10624);
nor U15433 (N_15433,N_14011,N_13990);
nor U15434 (N_15434,N_12444,N_11286);
xor U15435 (N_15435,N_10055,N_13215);
and U15436 (N_15436,N_11592,N_10311);
nor U15437 (N_15437,N_11784,N_14499);
nor U15438 (N_15438,N_14167,N_11608);
or U15439 (N_15439,N_13302,N_12215);
nand U15440 (N_15440,N_12020,N_10949);
xnor U15441 (N_15441,N_11218,N_14280);
nor U15442 (N_15442,N_14697,N_12691);
nand U15443 (N_15443,N_11626,N_11201);
and U15444 (N_15444,N_12157,N_11390);
nor U15445 (N_15445,N_12224,N_10979);
or U15446 (N_15446,N_10793,N_10332);
or U15447 (N_15447,N_10740,N_11814);
nand U15448 (N_15448,N_12965,N_13373);
or U15449 (N_15449,N_13049,N_14873);
xnor U15450 (N_15450,N_13425,N_13997);
and U15451 (N_15451,N_13015,N_11116);
nor U15452 (N_15452,N_10339,N_12265);
xor U15453 (N_15453,N_13856,N_10164);
or U15454 (N_15454,N_13207,N_11284);
xor U15455 (N_15455,N_10468,N_10767);
or U15456 (N_15456,N_10106,N_10165);
nor U15457 (N_15457,N_10221,N_11688);
nor U15458 (N_15458,N_13511,N_13961);
and U15459 (N_15459,N_13843,N_13281);
nor U15460 (N_15460,N_12405,N_13611);
nand U15461 (N_15461,N_10528,N_11172);
and U15462 (N_15462,N_13906,N_11563);
nor U15463 (N_15463,N_11096,N_13804);
nand U15464 (N_15464,N_13628,N_13642);
nand U15465 (N_15465,N_12174,N_11632);
or U15466 (N_15466,N_10459,N_10469);
or U15467 (N_15467,N_13543,N_10591);
and U15468 (N_15468,N_14196,N_12901);
or U15469 (N_15469,N_14838,N_14661);
nand U15470 (N_15470,N_12004,N_12337);
nor U15471 (N_15471,N_13208,N_11803);
nor U15472 (N_15472,N_11911,N_12277);
nand U15473 (N_15473,N_13666,N_10887);
and U15474 (N_15474,N_14743,N_14803);
nor U15475 (N_15475,N_11699,N_13414);
or U15476 (N_15476,N_13447,N_12057);
nand U15477 (N_15477,N_10788,N_10820);
or U15478 (N_15478,N_10294,N_13714);
and U15479 (N_15479,N_11721,N_13950);
nand U15480 (N_15480,N_14049,N_13263);
nand U15481 (N_15481,N_11881,N_11057);
nand U15482 (N_15482,N_12201,N_11880);
or U15483 (N_15483,N_11612,N_12845);
nand U15484 (N_15484,N_12945,N_14512);
and U15485 (N_15485,N_14967,N_14132);
nor U15486 (N_15486,N_14208,N_13062);
nor U15487 (N_15487,N_12284,N_13507);
and U15488 (N_15488,N_12018,N_10474);
nand U15489 (N_15489,N_10865,N_10441);
or U15490 (N_15490,N_10121,N_13234);
or U15491 (N_15491,N_11030,N_14301);
xor U15492 (N_15492,N_11875,N_10521);
or U15493 (N_15493,N_10532,N_11496);
xnor U15494 (N_15494,N_12758,N_10280);
or U15495 (N_15495,N_14825,N_10435);
xor U15496 (N_15496,N_14886,N_12318);
and U15497 (N_15497,N_10905,N_14188);
xnor U15498 (N_15498,N_10539,N_10112);
or U15499 (N_15499,N_10291,N_11606);
and U15500 (N_15500,N_14953,N_11397);
nor U15501 (N_15501,N_14445,N_10658);
xnor U15502 (N_15502,N_13852,N_14269);
xnor U15503 (N_15503,N_10950,N_11399);
nor U15504 (N_15504,N_10957,N_10619);
or U15505 (N_15505,N_10009,N_12504);
and U15506 (N_15506,N_13250,N_14309);
and U15507 (N_15507,N_10886,N_13133);
and U15508 (N_15508,N_13124,N_13649);
or U15509 (N_15509,N_10179,N_14336);
nor U15510 (N_15510,N_13288,N_12852);
and U15511 (N_15511,N_12392,N_10838);
or U15512 (N_15512,N_12605,N_13882);
nand U15513 (N_15513,N_12362,N_12906);
and U15514 (N_15514,N_14254,N_11957);
nand U15515 (N_15515,N_14446,N_10244);
or U15516 (N_15516,N_11301,N_10549);
or U15517 (N_15517,N_12492,N_11163);
or U15518 (N_15518,N_10834,N_11103);
xor U15519 (N_15519,N_14438,N_12259);
or U15520 (N_15520,N_14572,N_12329);
and U15521 (N_15521,N_14273,N_10352);
nand U15522 (N_15522,N_13962,N_14349);
nor U15523 (N_15523,N_12428,N_11382);
xnor U15524 (N_15524,N_14232,N_13708);
and U15525 (N_15525,N_10258,N_11835);
and U15526 (N_15526,N_12476,N_14379);
nor U15527 (N_15527,N_11128,N_14588);
xor U15528 (N_15528,N_12256,N_14189);
nor U15529 (N_15529,N_10270,N_11165);
or U15530 (N_15530,N_14602,N_14586);
xor U15531 (N_15531,N_13508,N_13738);
xor U15532 (N_15532,N_13571,N_11544);
nand U15533 (N_15533,N_12236,N_14436);
or U15534 (N_15534,N_11663,N_10093);
nor U15535 (N_15535,N_11224,N_10248);
xnor U15536 (N_15536,N_11066,N_14415);
nor U15537 (N_15537,N_12742,N_13185);
and U15538 (N_15538,N_10073,N_11493);
nor U15539 (N_15539,N_13164,N_10453);
xor U15540 (N_15540,N_10934,N_10861);
nor U15541 (N_15541,N_13670,N_14317);
and U15542 (N_15542,N_12123,N_11153);
or U15543 (N_15543,N_12096,N_13355);
xnor U15544 (N_15544,N_13740,N_12607);
or U15545 (N_15545,N_10704,N_14649);
nor U15546 (N_15546,N_14466,N_11111);
xnor U15547 (N_15547,N_12203,N_13717);
or U15548 (N_15548,N_10367,N_13675);
nor U15549 (N_15549,N_13996,N_12306);
or U15550 (N_15550,N_13779,N_11923);
or U15551 (N_15551,N_14587,N_10069);
or U15552 (N_15552,N_10242,N_11695);
xor U15553 (N_15553,N_11763,N_10129);
xnor U15554 (N_15554,N_12176,N_14666);
xor U15555 (N_15555,N_12910,N_10562);
xnor U15556 (N_15556,N_10020,N_11677);
xor U15557 (N_15557,N_11598,N_13706);
nor U15558 (N_15558,N_14995,N_14540);
and U15559 (N_15559,N_13908,N_12396);
nand U15560 (N_15560,N_14604,N_11368);
nand U15561 (N_15561,N_13131,N_10462);
nand U15562 (N_15562,N_13766,N_13237);
nand U15563 (N_15563,N_10741,N_14814);
xnor U15564 (N_15564,N_10716,N_13166);
nand U15565 (N_15565,N_13065,N_10012);
and U15566 (N_15566,N_12354,N_12620);
nor U15567 (N_15567,N_12685,N_14529);
nand U15568 (N_15568,N_12864,N_11188);
nand U15569 (N_15569,N_10779,N_13863);
xnor U15570 (N_15570,N_14734,N_12739);
and U15571 (N_15571,N_14026,N_11558);
xnor U15572 (N_15572,N_14827,N_13370);
or U15573 (N_15573,N_14008,N_11974);
or U15574 (N_15574,N_10185,N_12665);
nand U15575 (N_15575,N_12765,N_14933);
xor U15576 (N_15576,N_11450,N_10876);
and U15577 (N_15577,N_14012,N_13956);
nor U15578 (N_15578,N_10978,N_12163);
or U15579 (N_15579,N_12495,N_11680);
nor U15580 (N_15580,N_10272,N_10541);
xnor U15581 (N_15581,N_13176,N_11051);
nor U15582 (N_15582,N_14927,N_10895);
or U15583 (N_15583,N_10202,N_11363);
xor U15584 (N_15584,N_11010,N_12252);
xor U15585 (N_15585,N_10668,N_14258);
and U15586 (N_15586,N_12967,N_13454);
nand U15587 (N_15587,N_12317,N_10371);
and U15588 (N_15588,N_13743,N_13084);
xor U15589 (N_15589,N_13008,N_13160);
and U15590 (N_15590,N_13582,N_10839);
nor U15591 (N_15591,N_13539,N_12385);
and U15592 (N_15592,N_10553,N_12699);
xor U15593 (N_15593,N_10054,N_13246);
nand U15594 (N_15594,N_13318,N_13025);
xnor U15595 (N_15595,N_12133,N_12887);
nor U15596 (N_15596,N_12184,N_14329);
or U15597 (N_15597,N_11228,N_12443);
or U15598 (N_15598,N_12167,N_14545);
or U15599 (N_15599,N_11108,N_14455);
or U15600 (N_15600,N_10122,N_12897);
xor U15601 (N_15601,N_10552,N_12994);
or U15602 (N_15602,N_14627,N_14938);
xor U15603 (N_15603,N_13171,N_14648);
nor U15604 (N_15604,N_10515,N_13653);
nor U15605 (N_15605,N_12659,N_10529);
and U15606 (N_15606,N_12173,N_12903);
or U15607 (N_15607,N_11336,N_14882);
xor U15608 (N_15608,N_13605,N_14510);
or U15609 (N_15609,N_11888,N_10324);
or U15610 (N_15610,N_13969,N_11809);
nor U15611 (N_15611,N_11662,N_11359);
xnor U15612 (N_15612,N_14521,N_13226);
or U15613 (N_15613,N_14936,N_14224);
and U15614 (N_15614,N_11465,N_11559);
nor U15615 (N_15615,N_13800,N_12538);
xnor U15616 (N_15616,N_11209,N_14978);
nor U15617 (N_15617,N_12307,N_12532);
or U15618 (N_15618,N_10211,N_10419);
xnor U15619 (N_15619,N_14543,N_12078);
xnor U15620 (N_15620,N_11087,N_10902);
nand U15621 (N_15621,N_14327,N_14024);
and U15622 (N_15622,N_11886,N_13895);
nand U15623 (N_15623,N_11966,N_10341);
nand U15624 (N_15624,N_12779,N_12660);
or U15625 (N_15625,N_13705,N_14402);
or U15626 (N_15626,N_12349,N_11433);
and U15627 (N_15627,N_12183,N_11130);
nor U15628 (N_15628,N_12682,N_14906);
nor U15629 (N_15629,N_11647,N_12643);
nor U15630 (N_15630,N_12060,N_13513);
or U15631 (N_15631,N_14430,N_10660);
or U15632 (N_15632,N_12598,N_11442);
xnor U15633 (N_15633,N_13437,N_11144);
or U15634 (N_15634,N_11366,N_14597);
xnor U15635 (N_15635,N_11203,N_13384);
xnor U15636 (N_15636,N_11594,N_13607);
nor U15637 (N_15637,N_13194,N_14424);
xor U15638 (N_15638,N_10265,N_11836);
or U15639 (N_15639,N_14590,N_13415);
nor U15640 (N_15640,N_12453,N_12412);
nand U15641 (N_15641,N_12015,N_14720);
nand U15642 (N_15642,N_11065,N_11819);
xor U15643 (N_15643,N_11885,N_10914);
and U15644 (N_15644,N_13944,N_13591);
or U15645 (N_15645,N_14834,N_12438);
nor U15646 (N_15646,N_12720,N_12204);
and U15647 (N_15647,N_14689,N_12436);
nor U15648 (N_15648,N_13057,N_11098);
and U15649 (N_15649,N_11416,N_13058);
nand U15650 (N_15650,N_12863,N_14589);
or U15651 (N_15651,N_13985,N_14735);
nor U15652 (N_15652,N_10645,N_14530);
nor U15653 (N_15653,N_10928,N_12767);
or U15654 (N_15654,N_14879,N_12950);
or U15655 (N_15655,N_11035,N_13926);
or U15656 (N_15656,N_12313,N_12431);
nand U15657 (N_15657,N_12671,N_10299);
xnor U15658 (N_15658,N_12274,N_10189);
nand U15659 (N_15659,N_12615,N_11134);
and U15660 (N_15660,N_12955,N_14787);
nor U15661 (N_15661,N_14493,N_14050);
and U15662 (N_15662,N_11385,N_12788);
xnor U15663 (N_15663,N_12631,N_12278);
or U15664 (N_15664,N_14070,N_13752);
or U15665 (N_15665,N_14579,N_12037);
or U15666 (N_15666,N_13991,N_14079);
and U15667 (N_15667,N_11147,N_10434);
or U15668 (N_15668,N_13839,N_12712);
nand U15669 (N_15669,N_12159,N_11704);
xor U15670 (N_15670,N_11346,N_13816);
nor U15671 (N_15671,N_12496,N_14727);
nand U15672 (N_15672,N_12341,N_12912);
and U15673 (N_15673,N_10614,N_13411);
xor U15674 (N_15674,N_14497,N_10086);
and U15675 (N_15675,N_12563,N_10274);
nand U15676 (N_15676,N_13482,N_12409);
nor U15677 (N_15677,N_14015,N_13702);
nor U15678 (N_15678,N_10676,N_14737);
nand U15679 (N_15679,N_10033,N_14225);
and U15680 (N_15680,N_11313,N_12452);
nand U15681 (N_15681,N_11079,N_10702);
and U15682 (N_15682,N_13165,N_14107);
xnor U15683 (N_15683,N_13862,N_12973);
and U15684 (N_15684,N_13428,N_14483);
nand U15685 (N_15685,N_10822,N_13826);
or U15686 (N_15686,N_12031,N_14523);
and U15687 (N_15687,N_10000,N_13945);
nand U15688 (N_15688,N_13925,N_10413);
nand U15689 (N_15689,N_13413,N_11335);
nor U15690 (N_15690,N_11800,N_13114);
nor U15691 (N_15691,N_10489,N_10647);
xor U15692 (N_15692,N_11537,N_12870);
and U15693 (N_15693,N_13193,N_13331);
xnor U15694 (N_15694,N_13076,N_11635);
xnor U15695 (N_15695,N_12904,N_14328);
nor U15696 (N_15696,N_10220,N_10942);
nand U15697 (N_15697,N_10212,N_14811);
and U15698 (N_15698,N_12519,N_14983);
and U15699 (N_15699,N_12479,N_14348);
or U15700 (N_15700,N_13988,N_12566);
nor U15701 (N_15701,N_10835,N_11683);
and U15702 (N_15702,N_12841,N_13287);
or U15703 (N_15703,N_10975,N_14491);
or U15704 (N_15704,N_13104,N_13903);
or U15705 (N_15705,N_13067,N_11749);
xor U15706 (N_15706,N_10001,N_11682);
nand U15707 (N_15707,N_11131,N_14238);
xnor U15708 (N_15708,N_12740,N_12746);
xor U15709 (N_15709,N_11970,N_11817);
nor U15710 (N_15710,N_13905,N_11816);
xnor U15711 (N_15711,N_11107,N_11150);
and U15712 (N_15712,N_11257,N_13874);
and U15713 (N_15713,N_13755,N_12344);
nand U15714 (N_15714,N_12729,N_11145);
and U15715 (N_15715,N_10525,N_10695);
nand U15716 (N_15716,N_14612,N_12809);
xnor U15717 (N_15717,N_14299,N_14266);
xor U15718 (N_15718,N_11342,N_14142);
nor U15719 (N_15719,N_13117,N_14419);
nand U15720 (N_15720,N_11560,N_10217);
or U15721 (N_15721,N_14417,N_12737);
xnor U15722 (N_15722,N_12866,N_11871);
xnor U15723 (N_15723,N_11500,N_10105);
and U15724 (N_15724,N_14966,N_11756);
and U15725 (N_15725,N_10207,N_11467);
xnor U15726 (N_15726,N_11309,N_12033);
xnor U15727 (N_15727,N_10016,N_10295);
or U15728 (N_15728,N_10169,N_14639);
nand U15729 (N_15729,N_12970,N_10752);
xor U15730 (N_15730,N_10142,N_12199);
nand U15731 (N_15731,N_11766,N_12633);
or U15732 (N_15732,N_11008,N_13778);
or U15733 (N_15733,N_13072,N_10626);
and U15734 (N_15734,N_12961,N_10601);
nor U15735 (N_15735,N_14165,N_13073);
xor U15736 (N_15736,N_14240,N_10723);
xnor U15737 (N_15737,N_14635,N_11833);
nand U15738 (N_15738,N_12652,N_13711);
nand U15739 (N_15739,N_12733,N_14212);
or U15740 (N_15740,N_10340,N_10629);
or U15741 (N_15741,N_10731,N_13744);
nand U15742 (N_15742,N_14888,N_10671);
nand U15743 (N_15743,N_14353,N_13968);
nand U15744 (N_15744,N_14650,N_12579);
xor U15745 (N_15745,N_13754,N_11696);
or U15746 (N_15746,N_13529,N_13034);
or U15747 (N_15747,N_11407,N_11354);
and U15748 (N_15748,N_13120,N_10375);
nand U15749 (N_15749,N_11601,N_10823);
nor U15750 (N_15750,N_14986,N_13306);
nor U15751 (N_15751,N_13931,N_12288);
and U15752 (N_15752,N_12800,N_14754);
nor U15753 (N_15753,N_11401,N_14550);
and U15754 (N_15754,N_10560,N_13198);
nand U15755 (N_15755,N_14069,N_13763);
and U15756 (N_15756,N_12943,N_13138);
nor U15757 (N_15757,N_10162,N_12540);
nand U15758 (N_15758,N_11038,N_13803);
nor U15759 (N_15759,N_14960,N_11525);
nand U15760 (N_15760,N_13292,N_10141);
nor U15761 (N_15761,N_11312,N_10206);
and U15762 (N_15762,N_10090,N_13881);
nor U15763 (N_15763,N_10663,N_14113);
xnor U15764 (N_15764,N_10699,N_12043);
or U15765 (N_15765,N_14788,N_13186);
nand U15766 (N_15766,N_10765,N_11348);
xor U15767 (N_15767,N_11707,N_12567);
and U15768 (N_15768,N_14714,N_14096);
and U15769 (N_15769,N_10868,N_12531);
and U15770 (N_15770,N_10344,N_11306);
nor U15771 (N_15771,N_11730,N_11887);
nor U15772 (N_15772,N_13636,N_11542);
or U15773 (N_15773,N_13904,N_10583);
xor U15774 (N_15774,N_14711,N_12728);
and U15775 (N_15775,N_12179,N_12815);
nor U15776 (N_15776,N_11577,N_13071);
nor U15777 (N_15777,N_13930,N_10193);
or U15778 (N_15778,N_10648,N_10463);
nand U15779 (N_15779,N_10706,N_12730);
xnor U15780 (N_15780,N_14152,N_12330);
and U15781 (N_15781,N_12082,N_11085);
or U15782 (N_15782,N_10630,N_12473);
xnor U15783 (N_15783,N_10837,N_13797);
and U15784 (N_15784,N_10425,N_14637);
and U15785 (N_15785,N_14853,N_10497);
nor U15786 (N_15786,N_10690,N_13896);
nor U15787 (N_15787,N_14704,N_13444);
nor U15788 (N_15788,N_13593,N_14668);
xor U15789 (N_15789,N_12516,N_10916);
nand U15790 (N_15790,N_11579,N_14889);
or U15791 (N_15791,N_11105,N_14747);
xor U15792 (N_15792,N_14998,N_14041);
xor U15793 (N_15793,N_14946,N_13695);
xor U15794 (N_15794,N_13232,N_13174);
and U15795 (N_15795,N_12704,N_13316);
nand U15796 (N_15796,N_11735,N_10517);
nor U15797 (N_15797,N_10172,N_13821);
xnor U15798 (N_15798,N_11316,N_14996);
xor U15799 (N_15799,N_13774,N_11940);
nor U15800 (N_15800,N_13390,N_10657);
nor U15801 (N_15801,N_12962,N_11829);
nor U15802 (N_15802,N_12997,N_14361);
or U15803 (N_15803,N_14095,N_13833);
nand U15804 (N_15804,N_11069,N_14346);
and U15805 (N_15805,N_12918,N_12144);
xnor U15806 (N_15806,N_10018,N_13807);
or U15807 (N_15807,N_11481,N_11796);
xor U15808 (N_15808,N_13179,N_12507);
and U15809 (N_15809,N_12680,N_13693);
nor U15810 (N_15810,N_10813,N_12753);
xor U15811 (N_15811,N_11256,N_12249);
xor U15812 (N_15812,N_10768,N_11223);
and U15813 (N_15813,N_10314,N_11728);
or U15814 (N_15814,N_11455,N_14830);
or U15815 (N_15815,N_12039,N_14192);
and U15816 (N_15816,N_11801,N_13772);
or U15817 (N_15817,N_10501,N_10226);
nor U15818 (N_15818,N_12369,N_11238);
and U15819 (N_15819,N_14229,N_10451);
or U15820 (N_15820,N_12077,N_10191);
nand U15821 (N_15821,N_14081,N_12180);
xnor U15822 (N_15822,N_14899,N_14031);
nand U15823 (N_15823,N_12991,N_12045);
nand U15824 (N_15824,N_11196,N_11443);
and U15825 (N_15825,N_11920,N_12494);
xnor U15826 (N_15826,N_11969,N_10970);
and U15827 (N_15827,N_11992,N_14897);
and U15828 (N_15828,N_13613,N_13967);
and U15829 (N_15829,N_12522,N_13489);
or U15830 (N_15830,N_14204,N_11585);
nand U15831 (N_15831,N_13603,N_12676);
or U15832 (N_15832,N_10260,N_11852);
nor U15833 (N_15833,N_14984,N_10470);
nand U15834 (N_15834,N_12667,N_14796);
nand U15835 (N_15835,N_10857,N_13412);
xnor U15836 (N_15836,N_13562,N_12831);
and U15837 (N_15837,N_10418,N_12394);
xnor U15838 (N_15838,N_14028,N_11661);
nand U15839 (N_15839,N_14992,N_12061);
nor U15840 (N_15840,N_11693,N_13786);
and U15841 (N_15841,N_10103,N_11122);
xor U15842 (N_15842,N_12481,N_11420);
and U15843 (N_15843,N_13269,N_14516);
or U15844 (N_15844,N_14934,N_11774);
and U15845 (N_15845,N_11883,N_13552);
nand U15846 (N_15846,N_14741,N_13966);
or U15847 (N_15847,N_12086,N_10110);
nor U15848 (N_15848,N_11668,N_13584);
nor U15849 (N_15849,N_10972,N_12543);
nor U15850 (N_15850,N_13692,N_14640);
or U15851 (N_15851,N_13070,N_13802);
and U15852 (N_15852,N_14680,N_12122);
xor U15853 (N_15853,N_11275,N_14817);
xor U15854 (N_15854,N_11597,N_10064);
nand U15855 (N_15855,N_14760,N_14458);
or U15856 (N_15856,N_12824,N_10656);
or U15857 (N_15857,N_11611,N_12138);
nand U15858 (N_15858,N_13938,N_12340);
or U15859 (N_15859,N_14007,N_14591);
xnor U15860 (N_15860,N_10634,N_11825);
nand U15861 (N_15861,N_10200,N_14963);
and U15862 (N_15862,N_12708,N_10049);
and U15863 (N_15863,N_11991,N_10430);
and U15864 (N_15864,N_12861,N_14592);
and U15865 (N_15865,N_12748,N_10003);
nand U15866 (N_15866,N_12792,N_11700);
and U15867 (N_15867,N_12533,N_11717);
and U15868 (N_15868,N_11670,N_14844);
or U15869 (N_15869,N_10557,N_12925);
nand U15870 (N_15870,N_10852,N_13286);
and U15871 (N_15871,N_12433,N_12989);
nor U15872 (N_15872,N_12672,N_10396);
nor U15873 (N_15873,N_11757,N_10326);
nand U15874 (N_15874,N_12673,N_12843);
nand U15875 (N_15875,N_10190,N_13855);
nor U15876 (N_15876,N_11798,N_10449);
xor U15877 (N_15877,N_14865,N_14338);
nand U15878 (N_15878,N_14511,N_12622);
nand U15879 (N_15879,N_12094,N_10649);
or U15880 (N_15880,N_11532,N_11906);
and U15881 (N_15881,N_10445,N_11805);
nor U15882 (N_15882,N_10170,N_10426);
xor U15883 (N_15883,N_14739,N_10114);
nand U15884 (N_15884,N_10354,N_12402);
nand U15885 (N_15885,N_14605,N_10947);
xnor U15886 (N_15886,N_10760,N_13497);
nor U15887 (N_15887,N_12465,N_14956);
and U15888 (N_15888,N_14805,N_12888);
xor U15889 (N_15889,N_12217,N_13376);
and U15890 (N_15890,N_12602,N_10124);
xor U15891 (N_15891,N_13781,N_13074);
and U15892 (N_15892,N_10713,N_11810);
nand U15893 (N_15893,N_11570,N_10044);
and U15894 (N_15894,N_14987,N_13661);
or U15895 (N_15895,N_13357,N_11126);
nor U15896 (N_15896,N_10565,N_14891);
nor U15897 (N_15897,N_12279,N_13272);
or U15898 (N_15898,N_14206,N_11091);
nor U15899 (N_15899,N_14135,N_12883);
nand U15900 (N_15900,N_14615,N_12561);
xnor U15901 (N_15901,N_12706,N_12185);
and U15902 (N_15902,N_14461,N_10719);
xor U15903 (N_15903,N_12145,N_14611);
xor U15904 (N_15904,N_14343,N_14375);
nor U15905 (N_15905,N_10749,N_13371);
xor U15906 (N_15906,N_13615,N_13920);
nor U15907 (N_15907,N_12705,N_13959);
nor U15908 (N_15908,N_10397,N_10080);
nor U15909 (N_15909,N_12059,N_11180);
and U15910 (N_15910,N_11673,N_13883);
or U15911 (N_15911,N_10888,N_14642);
or U15912 (N_15912,N_12221,N_13617);
or U15913 (N_15913,N_12230,N_14673);
nand U15914 (N_15914,N_12829,N_13244);
xnor U15915 (N_15915,N_11726,N_13606);
and U15916 (N_15916,N_11794,N_12038);
nand U15917 (N_15917,N_11615,N_11742);
and U15918 (N_15918,N_10901,N_10996);
nor U15919 (N_15919,N_11600,N_12657);
or U15920 (N_15920,N_12830,N_10391);
xor U15921 (N_15921,N_11021,N_10939);
or U15922 (N_15922,N_14369,N_13867);
and U15923 (N_15923,N_14451,N_14408);
nor U15924 (N_15924,N_14148,N_10534);
and U15925 (N_15925,N_14502,N_11297);
or U15926 (N_15926,N_11812,N_10844);
nor U15927 (N_15927,N_14084,N_13710);
xnor U15928 (N_15928,N_13085,N_13265);
nand U15929 (N_15929,N_14706,N_10465);
nor U15930 (N_15930,N_11048,N_14122);
nor U15931 (N_15931,N_10485,N_12651);
and U15932 (N_15932,N_12161,N_11955);
nor U15933 (N_15933,N_11890,N_14223);
xnor U15934 (N_15934,N_10858,N_10335);
xnor U15935 (N_15935,N_12803,N_14383);
xnor U15936 (N_15936,N_13891,N_13301);
nand U15937 (N_15937,N_14626,N_12647);
nand U15938 (N_15938,N_10447,N_12587);
nand U15939 (N_15939,N_12931,N_11081);
nor U15940 (N_15940,N_14087,N_13688);
or U15941 (N_15941,N_13523,N_14746);
nor U15942 (N_15942,N_13241,N_10219);
nand U15943 (N_15943,N_12348,N_13271);
xnor U15944 (N_15944,N_11802,N_10566);
or U15945 (N_15945,N_14013,N_11170);
xor U15946 (N_15946,N_14326,N_14194);
nand U15947 (N_15947,N_13847,N_10516);
nor U15948 (N_15948,N_13815,N_11996);
or U15949 (N_15949,N_10428,N_11511);
nor U15950 (N_15950,N_12679,N_13505);
nand U15951 (N_15951,N_12041,N_11317);
nor U15952 (N_15952,N_12872,N_13805);
xor U15953 (N_15953,N_14676,N_10537);
nand U15954 (N_15954,N_10984,N_11530);
xor U15955 (N_15955,N_12714,N_12545);
xnor U15956 (N_15956,N_10827,N_14952);
and U15957 (N_15957,N_10748,N_10675);
or U15958 (N_15958,N_13381,N_12102);
nor U15959 (N_15959,N_12426,N_13153);
or U15960 (N_15960,N_14398,N_11573);
nor U15961 (N_15961,N_12695,N_11848);
or U15962 (N_15962,N_14029,N_13742);
or U15963 (N_15963,N_10288,N_12332);
xnor U15964 (N_15964,N_12303,N_12361);
nor U15965 (N_15965,N_12292,N_12417);
and U15966 (N_15966,N_12924,N_12952);
nor U15967 (N_15967,N_13554,N_13753);
nor U15968 (N_15968,N_10604,N_13223);
or U15969 (N_15969,N_13977,N_14104);
nand U15970 (N_15970,N_14517,N_10805);
nand U15971 (N_15971,N_13949,N_14389);
nand U15972 (N_15972,N_10321,N_12556);
nor U15973 (N_15973,N_11009,N_14533);
xnor U15974 (N_15974,N_11535,N_11777);
nand U15975 (N_15975,N_10424,N_13005);
xor U15976 (N_15976,N_12034,N_12808);
nor U15977 (N_15977,N_12125,N_14620);
nand U15978 (N_15978,N_12016,N_12470);
and U15979 (N_15979,N_10953,N_12687);
xor U15980 (N_15980,N_11436,N_12911);
and U15981 (N_15981,N_11516,N_11094);
xor U15982 (N_15982,N_14440,N_12413);
or U15983 (N_15983,N_10313,N_12554);
nor U15984 (N_15984,N_13201,N_12856);
or U15985 (N_15985,N_12136,N_10007);
nand U15986 (N_15986,N_14093,N_14279);
nand U15987 (N_15987,N_14020,N_11891);
or U15988 (N_15988,N_14667,N_12616);
and U15989 (N_15989,N_11947,N_10945);
and U15990 (N_15990,N_10075,N_12107);
xnor U15991 (N_15991,N_13974,N_10973);
nor U15992 (N_15992,N_14249,N_13170);
xnor U15993 (N_15993,N_11953,N_13590);
or U15994 (N_15994,N_12589,N_10109);
or U15995 (N_15995,N_14372,N_14363);
xor U15996 (N_15996,N_14022,N_11517);
nand U15997 (N_15997,N_11415,N_10188);
nand U15998 (N_15998,N_14289,N_10736);
and U15999 (N_15999,N_14671,N_12951);
and U16000 (N_16000,N_14793,N_14920);
or U16001 (N_16001,N_14469,N_10034);
or U16002 (N_16002,N_14303,N_14048);
or U16003 (N_16003,N_12053,N_10153);
and U16004 (N_16004,N_14473,N_11378);
or U16005 (N_16005,N_13980,N_14037);
nor U16006 (N_16006,N_11943,N_10889);
nor U16007 (N_16007,N_14758,N_12603);
nor U16008 (N_16008,N_10882,N_13472);
nor U16009 (N_16009,N_12621,N_14241);
nand U16010 (N_16010,N_12555,N_10883);
nand U16011 (N_16011,N_11174,N_12071);
or U16012 (N_16012,N_14541,N_12999);
or U16013 (N_16013,N_10840,N_13715);
and U16014 (N_16014,N_11851,N_10853);
and U16015 (N_16015,N_11240,N_13354);
nand U16016 (N_16016,N_10133,N_12546);
or U16017 (N_16017,N_11133,N_14345);
and U16018 (N_16018,N_11054,N_13252);
or U16019 (N_16019,N_12169,N_11509);
nand U16020 (N_16020,N_12534,N_11184);
and U16021 (N_16021,N_14457,N_14792);
nand U16022 (N_16022,N_11557,N_12946);
xnor U16023 (N_16023,N_14990,N_13470);
nand U16024 (N_16024,N_13317,N_14701);
nand U16025 (N_16025,N_14774,N_11937);
nand U16026 (N_16026,N_14140,N_14752);
xnor U16027 (N_16027,N_13641,N_12851);
xor U16028 (N_16028,N_11364,N_14912);
xnor U16029 (N_16029,N_12238,N_14252);
xor U16030 (N_16030,N_10983,N_10362);
nand U16031 (N_16031,N_12770,N_12244);
and U16032 (N_16032,N_10107,N_12356);
nor U16033 (N_16033,N_14596,N_12756);
nand U16034 (N_16034,N_12698,N_13189);
and U16035 (N_16035,N_10990,N_14134);
or U16036 (N_16036,N_10854,N_13509);
nand U16037 (N_16037,N_12783,N_10929);
nand U16038 (N_16038,N_14623,N_14672);
nor U16039 (N_16039,N_13432,N_11029);
nand U16040 (N_16040,N_11905,N_12291);
nand U16041 (N_16041,N_12905,N_10307);
nand U16042 (N_16042,N_12211,N_10859);
nor U16043 (N_16043,N_14218,N_10912);
nand U16044 (N_16044,N_12360,N_13841);
xnor U16045 (N_16045,N_10366,N_10641);
nor U16046 (N_16046,N_12403,N_11020);
or U16047 (N_16047,N_12958,N_12134);
and U16048 (N_16048,N_11529,N_13565);
nor U16049 (N_16049,N_13467,N_14866);
xnor U16050 (N_16050,N_12029,N_10333);
nand U16051 (N_16051,N_12012,N_13947);
or U16052 (N_16052,N_13916,N_13225);
xnor U16053 (N_16053,N_13018,N_13499);
and U16054 (N_16054,N_13498,N_14643);
xnor U16055 (N_16055,N_11959,N_14452);
or U16056 (N_16056,N_12855,N_11578);
or U16057 (N_16057,N_14914,N_13101);
nand U16058 (N_16058,N_14214,N_10891);
and U16059 (N_16059,N_11720,N_11406);
xor U16060 (N_16060,N_13304,N_10631);
and U16061 (N_16061,N_12153,N_14634);
and U16062 (N_16062,N_11519,N_14396);
and U16063 (N_16063,N_10828,N_13257);
nand U16064 (N_16064,N_13296,N_13031);
xor U16065 (N_16065,N_12158,N_13588);
nor U16066 (N_16066,N_11747,N_12456);
or U16067 (N_16067,N_11212,N_10712);
or U16068 (N_16068,N_11909,N_11202);
and U16069 (N_16069,N_14562,N_13942);
or U16070 (N_16070,N_10729,N_10233);
nor U16071 (N_16071,N_10772,N_14470);
xor U16072 (N_16072,N_14726,N_10568);
nor U16073 (N_16073,N_12381,N_10567);
and U16074 (N_16074,N_10360,N_14928);
nor U16075 (N_16075,N_10301,N_10778);
or U16076 (N_16076,N_11933,N_13631);
or U16077 (N_16077,N_11572,N_14757);
and U16078 (N_16078,N_11213,N_14150);
and U16079 (N_16079,N_12231,N_12116);
nor U16080 (N_16080,N_13984,N_14768);
nor U16081 (N_16081,N_14448,N_10709);
xor U16082 (N_16082,N_12975,N_11741);
nor U16083 (N_16083,N_11208,N_14765);
nor U16084 (N_16084,N_13546,N_12606);
nor U16085 (N_16085,N_13900,N_12222);
or U16086 (N_16086,N_13791,N_14106);
nor U16087 (N_16087,N_12583,N_12725);
and U16088 (N_16088,N_11908,N_13352);
and U16089 (N_16089,N_11583,N_11355);
nand U16090 (N_16090,N_11640,N_14202);
and U16091 (N_16091,N_10059,N_14409);
xnor U16092 (N_16092,N_13623,N_13761);
nor U16093 (N_16093,N_10187,N_10275);
and U16094 (N_16094,N_12771,N_10431);
nand U16095 (N_16095,N_12304,N_12137);
or U16096 (N_16096,N_10505,N_14270);
nand U16097 (N_16097,N_13894,N_12073);
nand U16098 (N_16098,N_10707,N_12160);
and U16099 (N_16099,N_10328,N_11941);
xor U16100 (N_16100,N_10255,N_13989);
or U16101 (N_16101,N_12058,N_14924);
nand U16102 (N_16102,N_10773,N_13527);
nand U16103 (N_16103,N_13919,N_14456);
nand U16104 (N_16104,N_12715,N_12827);
nor U16105 (N_16105,N_12254,N_12482);
and U16106 (N_16106,N_11723,N_12234);
nand U16107 (N_16107,N_12377,N_13212);
nor U16108 (N_16108,N_14698,N_14072);
and U16109 (N_16109,N_13180,N_11985);
xor U16110 (N_16110,N_13893,N_14979);
nand U16111 (N_16111,N_13573,N_14484);
xor U16112 (N_16112,N_13045,N_10586);
nand U16113 (N_16113,N_11628,N_12941);
xnor U16114 (N_16114,N_10605,N_11922);
nand U16115 (N_16115,N_11643,N_10068);
xnor U16116 (N_16116,N_10192,N_10414);
nor U16117 (N_16117,N_12755,N_10238);
nor U16118 (N_16118,N_10382,N_10892);
xnor U16119 (N_16119,N_10151,N_11319);
or U16120 (N_16120,N_13169,N_14972);
nand U16121 (N_16121,N_11733,N_14863);
nor U16122 (N_16122,N_11565,N_14331);
nand U16123 (N_16123,N_14187,N_11987);
nand U16124 (N_16124,N_10471,N_13751);
xor U16125 (N_16125,N_11381,N_12593);
or U16126 (N_16126,N_14308,N_10951);
and U16127 (N_16127,N_11248,N_10993);
nand U16128 (N_16128,N_13392,N_12716);
and U16129 (N_16129,N_10180,N_14652);
or U16130 (N_16130,N_13363,N_11644);
and U16131 (N_16131,N_10536,N_12223);
or U16132 (N_16132,N_13664,N_11773);
nor U16133 (N_16133,N_10705,N_11089);
and U16134 (N_16134,N_13952,N_13293);
xnor U16135 (N_16135,N_14585,N_14871);
nand U16136 (N_16136,N_10296,N_14664);
or U16137 (N_16137,N_10787,N_12688);
nor U16138 (N_16138,N_11033,N_10454);
or U16139 (N_16139,N_12508,N_14789);
or U16140 (N_16140,N_13093,N_11412);
nor U16141 (N_16141,N_10683,N_13674);
nor U16142 (N_16142,N_12801,N_11582);
and U16143 (N_16143,N_13405,N_14964);
or U16144 (N_16144,N_13890,N_14236);
or U16145 (N_16145,N_10897,N_13943);
nand U16146 (N_16146,N_11064,N_14339);
nand U16147 (N_16147,N_10573,N_11899);
or U16148 (N_16148,N_13873,N_14219);
nand U16149 (N_16149,N_14820,N_10821);
nand U16150 (N_16150,N_14166,N_10239);
and U16151 (N_16151,N_13420,N_10284);
nor U16152 (N_16152,N_12182,N_14234);
and U16153 (N_16153,N_11124,N_14519);
xnor U16154 (N_16154,N_12458,N_13116);
or U16155 (N_16155,N_12030,N_11821);
xnor U16156 (N_16156,N_14420,N_10243);
nor U16157 (N_16157,N_13261,N_11192);
and U16158 (N_16158,N_11499,N_10514);
xor U16159 (N_16159,N_14250,N_11605);
xor U16160 (N_16160,N_12207,N_14261);
nand U16161 (N_16161,N_12627,N_12066);
and U16162 (N_16162,N_13351,N_11337);
xor U16163 (N_16163,N_12868,N_12255);
xnor U16164 (N_16164,N_14636,N_14442);
xor U16165 (N_16165,N_13039,N_13367);
or U16166 (N_16166,N_14468,N_13877);
xnor U16167 (N_16167,N_12293,N_14862);
and U16168 (N_16168,N_11758,N_13303);
and U16169 (N_16169,N_11195,N_14276);
xor U16170 (N_16170,N_13407,N_12240);
xnor U16171 (N_16171,N_12814,N_10028);
and U16172 (N_16172,N_13776,N_12512);
nand U16173 (N_16173,N_14977,N_13681);
nor U16174 (N_16174,N_12499,N_11945);
nor U16175 (N_16175,N_10971,N_11468);
nand U16176 (N_16176,N_11157,N_11490);
nand U16177 (N_16177,N_14382,N_14217);
or U16178 (N_16178,N_14581,N_13537);
nor U16179 (N_16179,N_14646,N_14314);
xor U16180 (N_16180,N_13402,N_12505);
nor U16181 (N_16181,N_10334,N_12150);
xnor U16182 (N_16182,N_11541,N_12586);
nand U16183 (N_16183,N_14647,N_13240);
nor U16184 (N_16184,N_12423,N_14804);
nand U16185 (N_16185,N_14471,N_13568);
nor U16186 (N_16186,N_10140,N_13992);
nand U16187 (N_16187,N_10350,N_13994);
and U16188 (N_16188,N_13330,N_14108);
nand U16189 (N_16189,N_11619,N_11032);
nand U16190 (N_16190,N_13460,N_14333);
nand U16191 (N_16191,N_11561,N_14858);
nand U16192 (N_16192,N_13538,N_10218);
and U16193 (N_16193,N_14271,N_12398);
xnor U16194 (N_16194,N_14776,N_10096);
or U16195 (N_16195,N_13122,N_14981);
or U16196 (N_16196,N_14265,N_11595);
nand U16197 (N_16197,N_10620,N_10943);
xnor U16198 (N_16198,N_13660,N_12067);
and U16199 (N_16199,N_12218,N_10491);
and U16200 (N_16200,N_11609,N_14088);
and U16201 (N_16201,N_11148,N_10315);
xor U16202 (N_16202,N_14559,N_14783);
or U16203 (N_16203,N_10654,N_12986);
and U16204 (N_16204,N_10251,N_13602);
and U16205 (N_16205,N_12700,N_14669);
nand U16206 (N_16206,N_11279,N_12109);
and U16207 (N_16207,N_10467,N_12674);
nand U16208 (N_16208,N_13449,N_14245);
nand U16209 (N_16209,N_14163,N_13090);
or U16210 (N_16210,N_13364,N_10316);
nand U16211 (N_16211,N_11281,N_12164);
or U16212 (N_16212,N_10935,N_11502);
xor U16213 (N_16213,N_14624,N_11075);
and U16214 (N_16214,N_12996,N_10544);
nand U16215 (N_16215,N_10098,N_13685);
xnor U16216 (N_16216,N_10385,N_11333);
or U16217 (N_16217,N_11351,N_13639);
nor U16218 (N_16218,N_10197,N_11179);
nor U16219 (N_16219,N_12267,N_12848);
xnor U16220 (N_16220,N_12956,N_13134);
xor U16221 (N_16221,N_11614,N_13909);
and U16222 (N_16222,N_10019,N_11311);
nor U16223 (N_16223,N_13326,N_10866);
and U16224 (N_16224,N_10438,N_12577);
nand U16225 (N_16225,N_14582,N_12781);
xor U16226 (N_16226,N_12379,N_10594);
nand U16227 (N_16227,N_13599,N_12487);
xnor U16228 (N_16228,N_10849,N_14532);
nand U16229 (N_16229,N_14733,N_10167);
or U16230 (N_16230,N_11604,N_12799);
xnor U16231 (N_16231,N_14824,N_12594);
and U16232 (N_16232,N_14098,N_13365);
nand U16233 (N_16233,N_12697,N_12493);
and U16234 (N_16234,N_12650,N_10535);
or U16235 (N_16235,N_10511,N_12213);
or U16236 (N_16236,N_12764,N_14574);
and U16237 (N_16237,N_13098,N_14780);
nand U16238 (N_16238,N_13495,N_11387);
nand U16239 (N_16239,N_13587,N_11705);
or U16240 (N_16240,N_10769,N_10910);
and U16241 (N_16241,N_10691,N_11534);
xor U16242 (N_16242,N_12421,N_12595);
nor U16243 (N_16243,N_11621,N_14083);
or U16244 (N_16244,N_11078,N_12592);
nor U16245 (N_16245,N_13092,N_10285);
xor U16246 (N_16246,N_10811,N_10633);
nor U16247 (N_16247,N_10955,N_11822);
or U16248 (N_16248,N_10359,N_10095);
or U16249 (N_16249,N_13130,N_12285);
nand U16250 (N_16250,N_12131,N_10890);
nand U16251 (N_16251,N_11843,N_10644);
nor U16252 (N_16252,N_13002,N_10609);
xnor U16253 (N_16253,N_11326,N_10480);
xor U16254 (N_16254,N_10010,N_10176);
nand U16255 (N_16255,N_13409,N_13673);
and U16256 (N_16256,N_11315,N_12415);
xor U16257 (N_16257,N_14478,N_11734);
and U16258 (N_16258,N_12609,N_10327);
nand U16259 (N_16259,N_14976,N_13551);
nand U16260 (N_16260,N_14872,N_12498);
nor U16261 (N_16261,N_11109,N_12188);
nand U16262 (N_16262,N_12500,N_11138);
or U16263 (N_16263,N_10987,N_11331);
xnor U16264 (N_16264,N_14486,N_11115);
nor U16265 (N_16265,N_11751,N_10099);
xnor U16266 (N_16266,N_10444,N_11769);
nor U16267 (N_16267,N_12206,N_12761);
or U16268 (N_16268,N_13087,N_14707);
and U16269 (N_16269,N_12549,N_10235);
xnor U16270 (N_16270,N_10014,N_12907);
nor U16271 (N_16271,N_10782,N_11840);
nor U16272 (N_16272,N_11341,N_12001);
xor U16273 (N_16273,N_11625,N_13941);
nand U16274 (N_16274,N_13430,N_12559);
nor U16275 (N_16275,N_12713,N_13125);
and U16276 (N_16276,N_10029,N_11893);
nor U16277 (N_16277,N_14538,N_13283);
xnor U16278 (N_16278,N_14560,N_11574);
and U16279 (N_16279,N_13456,N_14716);
xnor U16280 (N_16280,N_14951,N_14034);
or U16281 (N_16281,N_14094,N_14892);
nor U16282 (N_16282,N_12209,N_11956);
xnor U16283 (N_16283,N_13679,N_14890);
and U16284 (N_16284,N_10800,N_13668);
or U16285 (N_16285,N_13545,N_14330);
or U16286 (N_16286,N_11543,N_14629);
or U16287 (N_16287,N_14745,N_13784);
and U16288 (N_16288,N_11430,N_11946);
and U16289 (N_16289,N_11280,N_10145);
and U16290 (N_16290,N_14641,N_13379);
nand U16291 (N_16291,N_12539,N_10092);
and U16292 (N_16292,N_13214,N_12442);
or U16293 (N_16293,N_10409,N_12214);
xnor U16294 (N_16294,N_12445,N_14127);
xnor U16295 (N_16295,N_13037,N_11308);
nand U16296 (N_16296,N_11884,N_12511);
nor U16297 (N_16297,N_10152,N_12321);
and U16298 (N_16298,N_14965,N_11845);
and U16299 (N_16299,N_12853,N_13727);
or U16300 (N_16300,N_12995,N_12055);
nand U16301 (N_16301,N_13291,N_14099);
nand U16302 (N_16302,N_14290,N_11844);
and U16303 (N_16303,N_14843,N_12378);
or U16304 (N_16304,N_14178,N_14561);
xor U16305 (N_16305,N_14802,N_12810);
xor U16306 (N_16306,N_11846,N_13549);
nand U16307 (N_16307,N_14243,N_11678);
or U16308 (N_16308,N_13764,N_13589);
nor U16309 (N_16309,N_14137,N_12429);
nand U16310 (N_16310,N_12670,N_12237);
and U16311 (N_16311,N_14659,N_11667);
nor U16312 (N_16312,N_13570,N_14404);
or U16313 (N_16313,N_11569,N_13957);
nor U16314 (N_16314,N_13777,N_12484);
nor U16315 (N_16315,N_10710,N_11797);
and U16316 (N_16316,N_10841,N_12934);
or U16317 (N_16317,N_10613,N_14553);
and U16318 (N_16318,N_14184,N_12656);
nand U16319 (N_16319,N_11706,N_14601);
xnor U16320 (N_16320,N_13408,N_14524);
xnor U16321 (N_16321,N_13720,N_10796);
and U16322 (N_16322,N_12152,N_12269);
xor U16323 (N_16323,N_12719,N_12280);
xnor U16324 (N_16324,N_10781,N_13842);
nand U16325 (N_16325,N_10867,N_11781);
or U16326 (N_16326,N_10032,N_10833);
nand U16327 (N_16327,N_13046,N_14785);
or U16328 (N_16328,N_14463,N_10545);
nor U16329 (N_16329,N_12915,N_14055);
or U16330 (N_16330,N_12170,N_14546);
nand U16331 (N_16331,N_10554,N_14781);
nor U16332 (N_16332,N_14394,N_11486);
nor U16333 (N_16333,N_10406,N_13787);
nor U16334 (N_16334,N_10524,N_13400);
nor U16335 (N_16335,N_14846,N_11653);
and U16336 (N_16336,N_13480,N_12786);
xor U16337 (N_16337,N_10666,N_10982);
nor U16338 (N_16338,N_14881,N_11447);
nand U16339 (N_16339,N_11849,N_10579);
and U16340 (N_16340,N_14923,N_13321);
xor U16341 (N_16341,N_12601,N_12990);
or U16342 (N_16342,N_13578,N_11160);
nand U16343 (N_16343,N_13620,N_13362);
or U16344 (N_16344,N_12322,N_14932);
nand U16345 (N_16345,N_14557,N_13423);
or U16346 (N_16346,N_11253,N_12063);
xnor U16347 (N_16347,N_13596,N_12416);
nand U16348 (N_16348,N_14670,N_14688);
nand U16349 (N_16349,N_11258,N_10094);
nor U16350 (N_16350,N_11477,N_14173);
xor U16351 (N_16351,N_14959,N_12380);
nor U16352 (N_16352,N_13598,N_10361);
nand U16353 (N_16353,N_10623,N_13183);
and U16354 (N_16354,N_10011,N_14175);
nor U16355 (N_16355,N_14393,N_14439);
and U16356 (N_16356,N_11549,N_13404);
and U16357 (N_16357,N_11652,N_11739);
and U16358 (N_16358,N_14799,N_11393);
nor U16359 (N_16359,N_11053,N_11215);
or U16360 (N_16360,N_14917,N_14075);
nand U16361 (N_16361,N_12040,N_12940);
nor U16362 (N_16362,N_11587,N_13254);
or U16363 (N_16363,N_14182,N_13152);
nand U16364 (N_16364,N_10318,N_13353);
nand U16365 (N_16365,N_11547,N_12793);
nand U16366 (N_16366,N_13553,N_13910);
nand U16367 (N_16367,N_14864,N_12514);
or U16368 (N_16368,N_11101,N_14251);
and U16369 (N_16369,N_12374,N_11675);
xor U16370 (N_16370,N_14197,N_14255);
and U16371 (N_16371,N_14816,N_11685);
nor U16372 (N_16372,N_14450,N_14875);
and U16373 (N_16373,N_13773,N_13723);
and U16374 (N_16374,N_13690,N_13635);
xnor U16375 (N_16375,N_10289,N_10035);
or U16376 (N_16376,N_13879,N_12625);
or U16377 (N_16377,N_12289,N_13983);
nand U16378 (N_16378,N_10276,N_12846);
nor U16379 (N_16379,N_11264,N_10348);
and U16380 (N_16380,N_10685,N_10331);
nor U16381 (N_16381,N_12884,N_13260);
nor U16382 (N_16382,N_13954,N_11235);
xor U16383 (N_16383,N_12143,N_14125);
and U16384 (N_16384,N_13648,N_14341);
nand U16385 (N_16385,N_10688,N_14742);
nand U16386 (N_16386,N_10547,N_10598);
nand U16387 (N_16387,N_12448,N_14489);
xnor U16388 (N_16388,N_11205,N_12011);
nand U16389 (N_16389,N_10518,N_13933);
nand U16390 (N_16390,N_13089,N_11334);
and U16391 (N_16391,N_14323,N_10615);
and U16392 (N_16392,N_14459,N_13394);
and U16393 (N_16393,N_11999,N_13669);
nor U16394 (N_16394,N_12804,N_11813);
and U16395 (N_16395,N_14220,N_11274);
nor U16396 (N_16396,N_13209,N_12794);
and U16397 (N_16397,N_13463,N_11330);
or U16398 (N_16398,N_14351,N_14210);
xnor U16399 (N_16399,N_12624,N_13610);
xnor U16400 (N_16400,N_13013,N_10061);
or U16401 (N_16401,N_12895,N_11251);
nand U16402 (N_16402,N_11266,N_13270);
and U16403 (N_16403,N_12491,N_10229);
or U16404 (N_16404,N_11666,N_11753);
nand U16405 (N_16405,N_13975,N_10636);
xnor U16406 (N_16406,N_10161,N_13350);
nor U16407 (N_16407,N_12520,N_13443);
nand U16408 (N_16408,N_10603,N_11552);
and U16409 (N_16409,N_11432,N_10273);
nor U16410 (N_16410,N_11161,N_12896);
or U16411 (N_16411,N_11017,N_10974);
nand U16412 (N_16412,N_12692,N_11135);
xnor U16413 (N_16413,N_14713,N_14856);
and U16414 (N_16414,N_11689,N_14786);
nor U16415 (N_16415,N_10743,N_12192);
xnor U16416 (N_16416,N_11090,N_11127);
nor U16417 (N_16417,N_12014,N_10673);
nand U16418 (N_16418,N_12171,N_10804);
and U16419 (N_16419,N_11588,N_14203);
nor U16420 (N_16420,N_12455,N_13656);
nor U16421 (N_16421,N_12635,N_14613);
or U16422 (N_16422,N_13178,N_11674);
nor U16423 (N_16423,N_14778,N_12604);
nor U16424 (N_16424,N_11862,N_13793);
xor U16425 (N_16425,N_10144,N_13233);
nor U16426 (N_16426,N_13730,N_12485);
nor U16427 (N_16427,N_11411,N_13850);
nand U16428 (N_16428,N_12365,N_13698);
nand U16429 (N_16429,N_13406,N_10759);
xor U16430 (N_16430,N_11169,N_11140);
and U16431 (N_16431,N_10687,N_10125);
nor U16432 (N_16432,N_13248,N_12461);
or U16433 (N_16433,N_13728,N_12513);
xnor U16434 (N_16434,N_13709,N_13123);
nand U16435 (N_16435,N_10138,N_13510);
xor U16436 (N_16436,N_10101,N_13030);
nor U16437 (N_16437,N_10325,N_11948);
nand U16438 (N_16438,N_12686,N_12083);
xor U16439 (N_16439,N_14322,N_13739);
xnor U16440 (N_16440,N_10040,N_14719);
xnor U16441 (N_16441,N_11993,N_12232);
and U16442 (N_16442,N_12938,N_14840);
and U16443 (N_16443,N_14791,N_13746);
or U16444 (N_16444,N_13689,N_10127);
nand U16445 (N_16445,N_11113,N_10574);
and U16446 (N_16446,N_14656,N_13567);
and U16447 (N_16447,N_14449,N_13493);
xor U16448 (N_16448,N_14281,N_14762);
nand U16449 (N_16449,N_11159,N_13377);
or U16450 (N_16450,N_10855,N_11589);
nand U16451 (N_16451,N_10559,N_13963);
or U16452 (N_16452,N_12510,N_10079);
nor U16453 (N_16453,N_13154,N_10323);
and U16454 (N_16454,N_13410,N_12049);
and U16455 (N_16455,N_10998,N_14051);
nand U16456 (N_16456,N_11239,N_13518);
and U16457 (N_16457,N_14131,N_13799);
nor U16458 (N_16458,N_13884,N_12282);
xor U16459 (N_16459,N_13103,N_14097);
or U16460 (N_16460,N_10309,N_13147);
and U16461 (N_16461,N_14207,N_14522);
nand U16462 (N_16462,N_14444,N_11186);
and U16463 (N_16463,N_14819,N_14421);
nor U16464 (N_16464,N_12840,N_14515);
xnor U16465 (N_16465,N_12301,N_12248);
and U16466 (N_16466,N_11853,N_14740);
or U16467 (N_16467,N_10116,N_11681);
nor U16468 (N_16468,N_11425,N_11936);
nor U16469 (N_16469,N_11867,N_11927);
nand U16470 (N_16470,N_13760,N_11080);
or U16471 (N_16471,N_12299,N_13458);
or U16472 (N_16472,N_14227,N_12370);
nor U16473 (N_16473,N_12272,N_12420);
and U16474 (N_16474,N_10659,N_10349);
xnor U16475 (N_16475,N_13424,N_14200);
nand U16476 (N_16476,N_14715,N_11654);
xor U16477 (N_16477,N_12196,N_13010);
nor U16478 (N_16478,N_12046,N_11329);
xnor U16479 (N_16479,N_10259,N_11178);
xor U16480 (N_16480,N_11288,N_13256);
and U16481 (N_16481,N_14918,N_14158);
xor U16482 (N_16482,N_12395,N_12653);
nand U16483 (N_16483,N_13595,N_12780);
and U16484 (N_16484,N_13634,N_13533);
nor U16485 (N_16485,N_12919,N_12927);
and U16486 (N_16486,N_13840,N_10308);
nor U16487 (N_16487,N_11474,N_14027);
xnor U16488 (N_16488,N_11011,N_10228);
xor U16489 (N_16489,N_13581,N_11716);
or U16490 (N_16490,N_10472,N_10790);
or U16491 (N_16491,N_13442,N_12197);
and U16492 (N_16492,N_14296,N_11973);
nand U16493 (N_16493,N_13899,N_13555);
nor U16494 (N_16494,N_11764,N_12118);
xnor U16495 (N_16495,N_11327,N_13464);
xor U16496 (N_16496,N_13880,N_11527);
and U16497 (N_16497,N_14949,N_12177);
xor U16498 (N_16498,N_13697,N_11318);
xnor U16499 (N_16499,N_11067,N_11472);
or U16500 (N_16500,N_10158,N_11759);
xor U16501 (N_16501,N_13024,N_12080);
nor U16502 (N_16502,N_14475,N_11004);
and U16503 (N_16503,N_11232,N_11379);
xnor U16504 (N_16504,N_11613,N_13319);
nand U16505 (N_16505,N_10616,N_14209);
and U16506 (N_16506,N_13345,N_10832);
nor U16507 (N_16507,N_11633,N_13322);
nor U16508 (N_16508,N_12352,N_10482);
xor U16509 (N_16509,N_12111,N_13148);
nor U16510 (N_16510,N_13928,N_13678);
or U16511 (N_16511,N_13846,N_11272);
and U16512 (N_16512,N_10870,N_11772);
and U16513 (N_16513,N_10948,N_11977);
nor U16514 (N_16514,N_13094,N_12382);
or U16515 (N_16515,N_10920,N_14332);
xnor U16516 (N_16516,N_13756,N_14662);
nand U16517 (N_16517,N_13385,N_13235);
and U16518 (N_16518,N_11650,N_10420);
nor U16519 (N_16519,N_10732,N_13451);
and U16520 (N_16520,N_10031,N_13940);
nand U16521 (N_16521,N_11070,N_14948);
xnor U16522 (N_16522,N_13080,N_13888);
and U16523 (N_16523,N_10810,N_11901);
nor U16524 (N_16524,N_12106,N_13917);
and U16525 (N_16525,N_14518,N_10071);
and U16526 (N_16526,N_14377,N_14818);
nor U16527 (N_16527,N_12949,N_13032);
nor U16528 (N_16528,N_10163,N_12386);
or U16529 (N_16529,N_12747,N_11458);
and U16530 (N_16530,N_12838,N_11480);
xor U16531 (N_16531,N_13981,N_12404);
nand U16532 (N_16532,N_11219,N_13313);
xor U16533 (N_16533,N_10408,N_11894);
nand U16534 (N_16534,N_10411,N_10909);
nand U16535 (N_16535,N_13817,N_10400);
or U16536 (N_16536,N_12439,N_11475);
and U16537 (N_16537,N_12275,N_10555);
nand U16538 (N_16538,N_14910,N_11930);
nand U16539 (N_16539,N_11826,N_14929);
or U16540 (N_16540,N_13136,N_12626);
or U16541 (N_16541,N_10558,N_10714);
nor U16542 (N_16542,N_13128,N_13142);
and U16543 (N_16543,N_13583,N_13026);
or U16544 (N_16544,N_14277,N_12591);
xnor U16545 (N_16545,N_13986,N_12573);
or U16546 (N_16546,N_14407,N_10642);
nand U16547 (N_16547,N_14288,N_11123);
and U16548 (N_16548,N_14437,N_13501);
nand U16549 (N_16549,N_13765,N_10246);
nor U16550 (N_16550,N_10739,N_14618);
and U16551 (N_16551,N_11915,N_10177);
and U16552 (N_16552,N_10432,N_10005);
or U16553 (N_16553,N_11055,N_14480);
nor U16554 (N_16554,N_14782,N_10651);
and U16555 (N_16555,N_11482,N_13017);
or U16556 (N_16556,N_12617,N_12225);
xnor U16557 (N_16557,N_14447,N_10664);
nand U16558 (N_16558,N_12899,N_11568);
or U16559 (N_16559,N_10874,N_13939);
or U16560 (N_16560,N_10674,N_13845);
or U16561 (N_16561,N_13782,N_13243);
nor U16562 (N_16562,N_14947,N_12857);
nand U16563 (N_16563,N_11837,N_14660);
and U16564 (N_16564,N_11118,N_10247);
and U16565 (N_16565,N_12105,N_14764);
and U16566 (N_16566,N_11984,N_14423);
nor U16567 (N_16567,N_13206,N_13267);
nor U16568 (N_16568,N_12229,N_12216);
and U16569 (N_16569,N_13921,N_14425);
and U16570 (N_16570,N_13659,N_12649);
and U16571 (N_16571,N_12097,N_14101);
nand U16572 (N_16572,N_14074,N_13126);
nand U16573 (N_16573,N_14429,N_10775);
nand U16574 (N_16574,N_10320,N_14136);
xor U16575 (N_16575,N_13630,N_11462);
xnor U16576 (N_16576,N_11622,N_14677);
or U16577 (N_16577,N_13713,N_14300);
xor U16578 (N_16578,N_14566,N_13492);
xor U16579 (N_16579,N_11423,N_12984);
nand U16580 (N_16580,N_11445,N_14366);
or U16581 (N_16581,N_14119,N_14867);
and U16582 (N_16582,N_10597,N_11786);
nand U16583 (N_16583,N_13042,N_13188);
nor U16584 (N_16584,N_10493,N_13577);
and U16585 (N_16585,N_12774,N_13999);
or U16586 (N_16586,N_13236,N_14149);
and U16587 (N_16587,N_13725,N_13418);
or U16588 (N_16588,N_13044,N_11249);
nor U16589 (N_16589,N_14982,N_14576);
nor U16590 (N_16590,N_12971,N_14903);
nor U16591 (N_16591,N_13970,N_12070);
and U16592 (N_16592,N_10128,N_12523);
nand U16593 (N_16593,N_14989,N_14040);
nand U16594 (N_16594,N_14091,N_10923);
nand U16595 (N_16595,N_14900,N_12425);
or U16596 (N_16596,N_10880,N_11637);
nand U16597 (N_16597,N_10662,N_11119);
nand U16598 (N_16598,N_10771,N_11429);
xor U16599 (N_16599,N_11376,N_10232);
nor U16600 (N_16600,N_12247,N_14179);
nor U16601 (N_16601,N_13686,N_14358);
nand U16602 (N_16602,N_10026,N_12736);
nand U16603 (N_16603,N_10669,N_10495);
and U16604 (N_16604,N_11623,N_14381);
and U16605 (N_16605,N_13446,N_10358);
and U16606 (N_16606,N_10954,N_10262);
xor U16607 (N_16607,N_11980,N_12718);
nor U16608 (N_16608,N_10572,N_11646);
nand U16609 (N_16609,N_13614,N_12638);
nor U16610 (N_16610,N_13901,N_10830);
or U16611 (N_16611,N_12375,N_14784);
nor U16612 (N_16612,N_13780,N_11371);
or U16613 (N_16613,N_10646,N_11808);
nand U16614 (N_16614,N_10607,N_12009);
nor U16615 (N_16615,N_14465,N_11424);
nand U16616 (N_16616,N_12005,N_12922);
nand U16617 (N_16617,N_11892,N_11545);
nand U16618 (N_16618,N_12802,N_12435);
or U16619 (N_16619,N_14848,N_11386);
or U16620 (N_16620,N_10801,N_12475);
xor U16621 (N_16621,N_13734,N_11658);
xnor U16622 (N_16622,N_10506,N_11932);
nor U16623 (N_16623,N_11649,N_13478);
nand U16624 (N_16624,N_12623,N_14077);
or U16625 (N_16625,N_12464,N_11584);
and U16626 (N_16626,N_14685,N_14413);
nand U16627 (N_16627,N_13627,N_10986);
nor U16628 (N_16628,N_14159,N_12294);
nand U16629 (N_16629,N_10678,N_14595);
nand U16630 (N_16630,N_14991,N_10442);
or U16631 (N_16631,N_13749,N_14930);
nor U16632 (N_16632,N_11338,N_14356);
nand U16633 (N_16633,N_10178,N_12319);
nand U16634 (N_16634,N_13624,N_13028);
nor U16635 (N_16635,N_10701,N_11013);
nand U16636 (N_16636,N_14133,N_13569);
and U16637 (N_16637,N_12220,N_11506);
and U16638 (N_16638,N_14535,N_13672);
nor U16639 (N_16639,N_12634,N_14190);
nor U16640 (N_16640,N_14453,N_14315);
or U16641 (N_16641,N_14334,N_13181);
nand U16642 (N_16642,N_12791,N_13159);
and U16643 (N_16643,N_12051,N_11618);
or U16644 (N_16644,N_10004,N_10039);
nand U16645 (N_16645,N_10754,N_14968);
nand U16646 (N_16646,N_13086,N_14732);
and U16647 (N_16647,N_12930,N_14958);
or U16648 (N_16648,N_10551,N_11441);
nor U16649 (N_16649,N_10082,N_14495);
xor U16650 (N_16650,N_12437,N_14056);
or U16651 (N_16651,N_13205,N_14829);
and U16652 (N_16652,N_13887,N_10637);
and U16653 (N_16653,N_11724,N_12552);
nand U16654 (N_16654,N_14045,N_14749);
xnor U16655 (N_16655,N_12681,N_14177);
nor U16656 (N_16656,N_10104,N_12689);
or U16657 (N_16657,N_13585,N_13586);
and U16658 (N_16658,N_11142,N_11183);
or U16659 (N_16659,N_13341,N_13077);
nand U16660 (N_16660,N_10410,N_12126);
xor U16661 (N_16661,N_14129,N_12569);
and U16662 (N_16662,N_12463,N_10569);
or U16663 (N_16663,N_11804,N_13993);
and U16664 (N_16664,N_12345,N_11785);
nand U16665 (N_16665,N_14725,N_10390);
nand U16666 (N_16666,N_13360,N_11072);
xnor U16667 (N_16667,N_11972,N_10355);
xor U16668 (N_16668,N_12391,N_10403);
nor U16669 (N_16669,N_10448,N_11263);
nand U16670 (N_16670,N_14558,N_14318);
nor U16671 (N_16671,N_12389,N_10037);
or U16672 (N_16672,N_14059,N_11260);
nor U16673 (N_16673,N_13655,N_11095);
and U16674 (N_16674,N_11982,N_13806);
xnor U16675 (N_16675,N_13224,N_13481);
nor U16676 (N_16676,N_11498,N_13506);
xor U16677 (N_16677,N_12127,N_13722);
and U16678 (N_16678,N_12113,N_12909);
or U16679 (N_16679,N_12168,N_12155);
xnor U16680 (N_16680,N_10478,N_13059);
or U16681 (N_16681,N_12754,N_11765);
and U16682 (N_16682,N_12873,N_13222);
and U16683 (N_16683,N_11332,N_11762);
and U16684 (N_16684,N_13060,N_12914);
xor U16685 (N_16685,N_12777,N_14221);
and U16686 (N_16686,N_12002,N_12489);
nand U16687 (N_16687,N_11580,N_13132);
and U16688 (N_16688,N_13987,N_13998);
or U16689 (N_16689,N_13680,N_11012);
xnor U16690 (N_16690,N_14775,N_11479);
or U16691 (N_16691,N_11403,N_10508);
xor U16692 (N_16692,N_13009,N_10851);
xor U16693 (N_16693,N_10894,N_11314);
or U16694 (N_16694,N_10198,N_12432);
nand U16695 (N_16695,N_10738,N_10727);
nand U16696 (N_16696,N_11702,N_14868);
nand U16697 (N_16697,N_13221,N_13088);
or U16698 (N_16698,N_10067,N_10208);
and U16699 (N_16699,N_10734,N_14282);
and U16700 (N_16700,N_11151,N_12019);
nand U16701 (N_16701,N_10097,N_13289);
xnor U16702 (N_16702,N_13878,N_14350);
and U16703 (N_16703,N_13646,N_10070);
xor U16704 (N_16704,N_11392,N_12678);
and U16705 (N_16705,N_10896,N_11063);
nor U16706 (N_16706,N_12355,N_14975);
and U16707 (N_16707,N_12471,N_12735);
nand U16708 (N_16708,N_12387,N_11740);
nand U16709 (N_16709,N_12486,N_10696);
xnor U16710 (N_16710,N_10698,N_10336);
nand U16711 (N_16711,N_14319,N_12833);
or U16712 (N_16712,N_11456,N_12191);
or U16713 (N_16713,N_14168,N_11296);
nand U16714 (N_16714,N_13006,N_10639);
nand U16715 (N_16715,N_10686,N_11776);
or U16716 (N_16716,N_14435,N_11451);
and U16717 (N_16717,N_14406,N_13665);
or U16718 (N_16718,N_12302,N_11736);
nor U16719 (N_16719,N_12056,N_13683);
xor U16720 (N_16720,N_14567,N_11501);
xnor U16721 (N_16721,N_10737,N_13268);
xor U16722 (N_16722,N_10956,N_14230);
nor U16723 (N_16723,N_11710,N_13038);
or U16724 (N_16724,N_13305,N_10147);
nor U16725 (N_16725,N_13724,N_14729);
nand U16726 (N_16726,N_10617,N_12521);
or U16727 (N_16727,N_13055,N_12068);
or U16728 (N_16728,N_13747,N_14426);
nand U16729 (N_16729,N_10204,N_10088);
xor U16730 (N_16730,N_10436,N_10250);
and U16731 (N_16731,N_13767,N_13022);
and U16732 (N_16732,N_12632,N_13792);
xor U16733 (N_16733,N_13455,N_14973);
nand U16734 (N_16734,N_13810,N_12350);
and U16735 (N_16735,N_10926,N_13192);
and U16736 (N_16736,N_12544,N_10994);
nor U16737 (N_16737,N_13308,N_10387);
nor U16738 (N_16738,N_11916,N_12239);
or U16739 (N_16739,N_14477,N_11576);
nand U16740 (N_16740,N_10047,N_12977);
nand U16741 (N_16741,N_10089,N_14268);
nor U16742 (N_16742,N_12342,N_13601);
xnor U16743 (N_16743,N_12353,N_10267);
or U16744 (N_16744,N_14621,N_12062);
and U16745 (N_16745,N_13182,N_11727);
or U16746 (N_16746,N_10911,N_10464);
nand U16747 (N_16747,N_11156,N_10056);
or U16748 (N_16748,N_11000,N_12200);
xor U16749 (N_16749,N_12834,N_10873);
xnor U16750 (N_16750,N_14694,N_10747);
or U16751 (N_16751,N_12515,N_10527);
and U16752 (N_16752,N_12668,N_14033);
or U16753 (N_16753,N_13871,N_14999);
and U16754 (N_16754,N_13161,N_12089);
or U16755 (N_16755,N_10621,N_11352);
nand U16756 (N_16756,N_11061,N_11273);
or U16757 (N_16757,N_10940,N_13150);
xor U16758 (N_16758,N_10186,N_14264);
nor U16759 (N_16759,N_14898,N_13081);
nand U16760 (N_16760,N_13580,N_13748);
or U16761 (N_16761,N_12075,N_13453);
or U16762 (N_16762,N_13918,N_11627);
nand U16763 (N_16763,N_12763,N_10751);
and U16764 (N_16764,N_10181,N_14531);
nor U16765 (N_16765,N_14063,N_12309);
nor U16766 (N_16766,N_10661,N_13440);
or U16767 (N_16767,N_11422,N_13036);
nor U16768 (N_16768,N_10667,N_10596);
xnor U16769 (N_16769,N_10346,N_12886);
or U16770 (N_16770,N_11768,N_10842);
xor U16771 (N_16771,N_14337,N_10717);
and U16772 (N_16772,N_13129,N_13542);
or U16773 (N_16773,N_14505,N_12928);
or U16774 (N_16774,N_14038,N_11795);
nand U16775 (N_16775,N_12141,N_13099);
nor U16776 (N_16776,N_13861,N_14170);
xnor U16777 (N_16777,N_11783,N_14302);
xor U16778 (N_16778,N_14548,N_12117);
nand U16779 (N_16779,N_14902,N_11389);
nor U16780 (N_16780,N_13914,N_14705);
and U16781 (N_16781,N_12976,N_11444);
and U16782 (N_16782,N_13468,N_11452);
xnor U16783 (N_16783,N_11775,N_12590);
xor U16784 (N_16784,N_10108,N_10030);
nand U16785 (N_16785,N_14355,N_13707);
and U16786 (N_16786,N_13771,N_13652);
and U16787 (N_16787,N_14380,N_14724);
nor U16788 (N_16788,N_12325,N_10785);
or U16789 (N_16789,N_14285,N_14877);
or U16790 (N_16790,N_13168,N_10137);
nor U16791 (N_16791,N_14428,N_12787);
and U16792 (N_16792,N_13971,N_10510);
and U16793 (N_16793,N_13633,N_12894);
or U16794 (N_16794,N_13393,N_14042);
xnor U16795 (N_16795,N_14498,N_14401);
xor U16796 (N_16796,N_10115,N_10570);
nor U16797 (N_16797,N_12640,N_10254);
nand U16798 (N_16798,N_14798,N_11039);
or U16799 (N_16799,N_12684,N_10703);
nand U16800 (N_16800,N_14464,N_12954);
nor U16801 (N_16801,N_10439,N_12112);
xnor U16802 (N_16802,N_12743,N_10726);
nand U16803 (N_16803,N_11466,N_12359);
xor U16804 (N_16804,N_10022,N_10100);
and U16805 (N_16805,N_11868,N_13875);
nor U16806 (N_16806,N_12662,N_14944);
nor U16807 (N_16807,N_13671,N_10329);
and U16808 (N_16808,N_13041,N_13608);
and U16809 (N_16809,N_11952,N_12219);
and U16810 (N_16810,N_11237,N_14810);
or U16811 (N_16811,N_13450,N_13490);
nand U16812 (N_16812,N_12542,N_13328);
xor U16813 (N_16813,N_13638,N_11989);
nand U16814 (N_16814,N_11104,N_14058);
nand U16815 (N_16815,N_11971,N_12526);
nand U16816 (N_16816,N_14945,N_12129);
or U16817 (N_16817,N_14100,N_14030);
nand U16818 (N_16818,N_14580,N_13531);
and U16819 (N_16819,N_11409,N_11461);
nor U16820 (N_16820,N_13955,N_10722);
nor U16821 (N_16821,N_12812,N_13029);
nand U16822 (N_16822,N_10640,N_11729);
nor U16823 (N_16823,N_10919,N_11504);
or U16824 (N_16824,N_11575,N_13597);
nand U16825 (N_16825,N_10600,N_12312);
nor U16826 (N_16826,N_13264,N_12817);
and U16827 (N_16827,N_11715,N_12611);
and U16828 (N_16828,N_13312,N_14808);
nand U16829 (N_16829,N_12981,N_11536);
and U16830 (N_16830,N_14021,N_11292);
nand U16831 (N_16831,N_11254,N_14090);
nand U16832 (N_16832,N_10612,N_13768);
nor U16833 (N_16833,N_11995,N_10927);
xor U16834 (N_16834,N_14600,N_13476);
or U16835 (N_16835,N_13069,N_10053);
and U16836 (N_16836,N_10721,N_14755);
or U16837 (N_16837,N_12095,N_14014);
or U16838 (N_16838,N_14047,N_11199);
xor U16839 (N_16839,N_13912,N_11538);
and U16840 (N_16840,N_11154,N_11997);
nor U16841 (N_16841,N_11655,N_14994);
or U16842 (N_16842,N_10533,N_11823);
xor U16843 (N_16843,N_12572,N_11719);
or U16844 (N_16844,N_11790,N_14831);
and U16845 (N_16845,N_10507,N_10319);
and U16846 (N_16846,N_13403,N_12877);
or U16847 (N_16847,N_14851,N_11491);
and U16848 (N_16848,N_12202,N_11146);
or U16849 (N_16849,N_12723,N_13075);
and U16850 (N_16850,N_10770,N_13657);
or U16851 (N_16851,N_10205,N_12766);
nor U16852 (N_16852,N_14386,N_11722);
nor U16853 (N_16853,N_13844,N_13342);
nand U16854 (N_16854,N_13687,N_14985);
nand U16855 (N_16855,N_13762,N_13798);
xnor U16856 (N_16856,N_14260,N_10803);
nand U16857 (N_16857,N_11789,N_10546);
and U16858 (N_16858,N_14460,N_14638);
nor U16859 (N_16859,N_11787,N_12666);
nor U16860 (N_16860,N_14154,N_12724);
and U16861 (N_16861,N_13047,N_12933);
xnor U16862 (N_16862,N_14751,N_10672);
or U16863 (N_16863,N_11231,N_13061);
nand U16864 (N_16864,N_13329,N_14941);
or U16865 (N_16865,N_14141,N_10814);
xnor U16866 (N_16866,N_10809,N_13066);
xor U16867 (N_16867,N_11049,N_11879);
and U16868 (N_16868,N_12287,N_11365);
nor U16869 (N_16869,N_10904,N_13644);
and U16870 (N_16870,N_11388,N_12246);
or U16871 (N_16871,N_13284,N_13391);
nand U16872 (N_16872,N_12351,N_10548);
or U16873 (N_16873,N_11554,N_12993);
and U16874 (N_16874,N_11599,N_12557);
nand U16875 (N_16875,N_14162,N_12727);
nor U16876 (N_16876,N_14939,N_11463);
xnor U16877 (N_16877,N_10885,N_12347);
and U16878 (N_16878,N_12778,N_12064);
nand U16879 (N_16879,N_14278,N_13866);
or U16880 (N_16880,N_12547,N_12584);
xnor U16881 (N_16881,N_10582,N_13864);
nand U16882 (N_16882,N_12466,N_13109);
or U16883 (N_16883,N_14462,N_14942);
nor U16884 (N_16884,N_12529,N_14573);
xnor U16885 (N_16885,N_11526,N_13504);
or U16886 (N_16886,N_11417,N_13378);
nor U16887 (N_16887,N_12081,N_14509);
or U16888 (N_16888,N_11831,N_13550);
or U16889 (N_16889,N_12022,N_11289);
or U16890 (N_16890,N_12953,N_11990);
nand U16891 (N_16891,N_13229,N_13314);
or U16892 (N_16892,N_13298,N_14913);
or U16893 (N_16893,N_13190,N_13475);
or U16894 (N_16894,N_13556,N_14699);
xnor U16895 (N_16895,N_12535,N_12010);
nor U16896 (N_16896,N_10681,N_10416);
and U16897 (N_16897,N_10540,N_10744);
xor U16898 (N_16898,N_12172,N_13600);
or U16899 (N_16899,N_14925,N_13522);
nor U16900 (N_16900,N_14118,N_13202);
and U16901 (N_16901,N_13282,N_14443);
nor U16902 (N_16902,N_11454,N_14908);
or U16903 (N_16903,N_14753,N_13948);
nor U16904 (N_16904,N_12842,N_12146);
xor U16905 (N_16905,N_12488,N_10376);
and U16906 (N_16906,N_14124,N_11437);
nand U16907 (N_16907,N_13712,N_13079);
xor U16908 (N_16908,N_10680,N_12527);
and U16909 (N_16909,N_14665,N_10166);
or U16910 (N_16910,N_13359,N_10602);
xnor U16911 (N_16911,N_10017,N_14384);
and U16912 (N_16912,N_11230,N_12315);
nor U16913 (N_16913,N_12027,N_13958);
xnor U16914 (N_16914,N_10078,N_13929);
or U16915 (N_16915,N_11616,N_14185);
xor U16916 (N_16916,N_11339,N_12983);
xor U16917 (N_16917,N_10236,N_10580);
nor U16918 (N_16918,N_14213,N_12964);
or U16919 (N_16919,N_11861,N_11566);
nand U16920 (N_16920,N_11060,N_11373);
nor U16921 (N_16921,N_11031,N_13592);
xnor U16922 (N_16922,N_14645,N_14199);
nor U16923 (N_16923,N_11942,N_12245);
xor U16924 (N_16924,N_10789,N_11340);
and U16925 (N_16925,N_13902,N_12702);
nor U16926 (N_16926,N_11426,N_11521);
nand U16927 (N_16927,N_14728,N_11910);
or U16928 (N_16928,N_13651,N_11824);
and U16929 (N_16929,N_12446,N_12711);
and U16930 (N_16930,N_14712,N_12818);
nor U16931 (N_16931,N_14772,N_13796);
and U16932 (N_16932,N_12006,N_12558);
nor U16933 (N_16933,N_14500,N_10944);
xnor U16934 (N_16934,N_12114,N_11375);
nand U16935 (N_16935,N_13625,N_13158);
xnor U16936 (N_16936,N_11591,N_14400);
xnor U16937 (N_16937,N_14970,N_14068);
or U16938 (N_16938,N_11492,N_10050);
xor U16939 (N_16939,N_14883,N_10794);
nand U16940 (N_16940,N_14874,N_11617);
xor U16941 (N_16941,N_10655,N_14895);
nand U16942 (N_16942,N_13417,N_13102);
nor U16943 (N_16943,N_10384,N_13149);
and U16944 (N_16944,N_12744,N_12072);
nand U16945 (N_16945,N_11283,N_11287);
or U16946 (N_16946,N_10182,N_14235);
xor U16947 (N_16947,N_13536,N_10742);
xnor U16948 (N_16948,N_10906,N_10774);
or U16949 (N_16949,N_14822,N_14644);
and U16950 (N_16950,N_12430,N_11418);
nor U16951 (N_16951,N_14771,N_10816);
nand U16952 (N_16952,N_12271,N_10051);
nand U16953 (N_16953,N_12658,N_11044);
and U16954 (N_16954,N_13398,N_13007);
nor U16955 (N_16955,N_12156,N_11353);
xnor U16956 (N_16956,N_14017,N_10697);
xor U16957 (N_16957,N_11453,N_11820);
nand U16958 (N_16958,N_14263,N_10455);
or U16959 (N_16959,N_11691,N_10643);
xnor U16960 (N_16960,N_14291,N_10917);
and U16961 (N_16961,N_11320,N_12101);
or U16962 (N_16962,N_14593,N_14837);
nand U16963 (N_16963,N_13978,N_13937);
nor U16964 (N_16964,N_12447,N_13832);
nor U16965 (N_16965,N_14730,N_14228);
or U16966 (N_16966,N_14321,N_10863);
nor U16967 (N_16967,N_14487,N_11954);
or U16968 (N_16968,N_10898,N_13052);
or U16969 (N_16969,N_14583,N_11358);
nand U16970 (N_16970,N_11282,N_14663);
xnor U16971 (N_16971,N_14313,N_13106);
nand U16972 (N_16972,N_13775,N_11056);
or U16973 (N_16973,N_14607,N_11222);
nor U16974 (N_16974,N_13332,N_12376);
nand U16975 (N_16975,N_11988,N_12960);
xnor U16976 (N_16976,N_12762,N_13333);
or U16977 (N_16977,N_11303,N_11360);
nand U16978 (N_16978,N_10650,N_14800);
nand U16979 (N_16979,N_13356,N_10271);
nand U16980 (N_16980,N_10879,N_12826);
or U16981 (N_16981,N_14506,N_11755);
or U16982 (N_16982,N_11553,N_12942);
or U16983 (N_16983,N_11074,N_13927);
nand U16984 (N_16984,N_12920,N_11350);
and U16985 (N_16985,N_14239,N_13279);
or U16986 (N_16986,N_10745,N_10374);
nor U16987 (N_16987,N_12100,N_14893);
xor U16988 (N_16988,N_11839,N_11047);
and U16989 (N_16989,N_14684,N_14174);
nand U16990 (N_16990,N_11168,N_12837);
nor U16991 (N_16991,N_13054,N_10526);
and U16992 (N_16992,N_11895,N_12677);
or U16993 (N_16993,N_12582,N_12985);
nand U16994 (N_16994,N_13643,N_10967);
and U16995 (N_16995,N_11413,N_10437);
xor U16996 (N_16996,N_10877,N_14632);
and U16997 (N_16997,N_11471,N_14036);
nand U16998 (N_16998,N_12642,N_14940);
xor U16999 (N_16999,N_13622,N_11564);
nand U17000 (N_17000,N_13431,N_12709);
and U17001 (N_17001,N_12902,N_11718);
xor U17002 (N_17002,N_13483,N_10757);
nand U17003 (N_17003,N_14835,N_12434);
xor U17004 (N_17004,N_12451,N_13684);
xor U17005 (N_17005,N_10962,N_13144);
or U17006 (N_17006,N_13172,N_13853);
and U17007 (N_17007,N_10523,N_10347);
nand U17008 (N_17008,N_10786,N_13719);
xnor U17009 (N_17009,N_10461,N_11651);
nand U17010 (N_17010,N_12401,N_14481);
and U17011 (N_17011,N_10756,N_13349);
xnor U17012 (N_17012,N_12932,N_12103);
xnor U17013 (N_17013,N_13162,N_10618);
xnor U17014 (N_17014,N_10393,N_12849);
nand U17015 (N_17015,N_11226,N_13127);
or U17016 (N_17016,N_14054,N_12819);
nand U17017 (N_17017,N_10968,N_14744);
xnor U17018 (N_17018,N_12454,N_11062);
and U17019 (N_17019,N_12338,N_10908);
xor U17020 (N_17020,N_14919,N_14564);
and U17021 (N_17021,N_11114,N_10043);
nand U17022 (N_17022,N_14773,N_13438);
nor U17023 (N_17023,N_10708,N_13824);
nor U17024 (N_17024,N_13340,N_11771);
and U17025 (N_17025,N_14365,N_14434);
or U17026 (N_17026,N_13790,N_12789);
nand U17027 (N_17027,N_10531,N_11435);
or U17028 (N_17028,N_13230,N_12008);
nand U17029 (N_17029,N_10946,N_13121);
or U17030 (N_17030,N_13200,N_10477);
xnor U17031 (N_17031,N_13474,N_13735);
or U17032 (N_17032,N_14700,N_10931);
or U17033 (N_17033,N_10592,N_10159);
nand U17034 (N_17034,N_11694,N_14293);
xor U17035 (N_17035,N_13239,N_12462);
xnor U17036 (N_17036,N_10850,N_11866);
xnor U17037 (N_17037,N_10576,N_10575);
and U17038 (N_17038,N_12091,N_12574);
xor U17039 (N_17039,N_14032,N_13386);
and U17040 (N_17040,N_12140,N_13187);
nand U17041 (N_17041,N_10132,N_11964);
nand U17042 (N_17042,N_10317,N_14501);
xor U17043 (N_17043,N_12646,N_13211);
nand U17044 (N_17044,N_14608,N_13466);
and U17045 (N_17045,N_13441,N_10377);
or U17046 (N_17046,N_14631,N_12363);
nand U17047 (N_17047,N_13564,N_11744);
nor U17048 (N_17048,N_12988,N_10045);
xor U17049 (N_17049,N_10401,N_10062);
nor U17050 (N_17050,N_11938,N_11497);
nor U17051 (N_17051,N_14807,N_11631);
or U17052 (N_17052,N_12655,N_12399);
and U17053 (N_17053,N_10415,N_13184);
xnor U17054 (N_17054,N_11900,N_10960);
nand U17055 (N_17055,N_14577,N_13346);
or U17056 (N_17056,N_11508,N_10298);
and U17057 (N_17057,N_14340,N_10353);
nor U17058 (N_17058,N_13173,N_12132);
xor U17059 (N_17059,N_11459,N_12331);
nand U17060 (N_17060,N_10041,N_12683);
or U17061 (N_17061,N_13118,N_13662);
nor U17062 (N_17062,N_12879,N_11807);
and U17063 (N_17063,N_10084,N_11221);
nor U17064 (N_17064,N_10131,N_11978);
or U17065 (N_17065,N_11045,N_11112);
and U17066 (N_17066,N_11531,N_12276);
and U17067 (N_17067,N_11189,N_12641);
or U17068 (N_17068,N_13632,N_14310);
or U17069 (N_17069,N_14169,N_10730);
nand U17070 (N_17070,N_14554,N_14568);
and U17071 (N_17071,N_11019,N_13157);
xor U17072 (N_17072,N_13388,N_12305);
or U17073 (N_17073,N_10048,N_12614);
nand U17074 (N_17074,N_13528,N_10509);
nor U17075 (N_17075,N_12175,N_10864);
or U17076 (N_17076,N_11761,N_11856);
and U17077 (N_17077,N_12588,N_12871);
and U17078 (N_17078,N_12502,N_14599);
nand U17079 (N_17079,N_14297,N_12189);
xnor U17080 (N_17080,N_11068,N_13951);
nor U17081 (N_17081,N_13001,N_10791);
xor U17082 (N_17082,N_10985,N_14073);
nand U17083 (N_17083,N_14023,N_11850);
and U17084 (N_17084,N_14547,N_14172);
nand U17085 (N_17085,N_12805,N_13626);
nor U17086 (N_17086,N_13375,N_14193);
and U17087 (N_17087,N_13512,N_13757);
nand U17088 (N_17088,N_12525,N_14880);
nand U17089 (N_17089,N_13242,N_14721);
xnor U17090 (N_17090,N_12243,N_14410);
or U17091 (N_17091,N_12166,N_10281);
xor U17092 (N_17092,N_13228,N_12368);
or U17093 (N_17093,N_12333,N_11919);
and U17094 (N_17094,N_13913,N_11778);
and U17095 (N_17095,N_14298,N_11267);
and U17096 (N_17096,N_10015,N_10530);
or U17097 (N_17097,N_10913,N_12822);
nand U17098 (N_17098,N_14431,N_14284);
nor U17099 (N_17099,N_11040,N_12000);
and U17100 (N_17100,N_14052,N_14537);
xnor U17101 (N_17101,N_10113,N_11034);
xor U17102 (N_17102,N_11246,N_10795);
xor U17103 (N_17103,N_11610,N_10136);
xnor U17104 (N_17104,N_11590,N_14679);
or U17105 (N_17105,N_14399,N_12878);
nand U17106 (N_17106,N_14116,N_13502);
xor U17107 (N_17107,N_14342,N_13534);
nand U17108 (N_17108,N_11505,N_13396);
and U17109 (N_17109,N_11660,N_13143);
nor U17110 (N_17110,N_10587,N_14657);
xnor U17111 (N_17111,N_11524,N_12422);
nand U17112 (N_17112,N_12120,N_12517);
and U17113 (N_17113,N_10452,N_14901);
xnor U17114 (N_17114,N_13809,N_11713);
nor U17115 (N_17115,N_10223,N_13629);
nand U17116 (N_17116,N_12693,N_14089);
nand U17117 (N_17117,N_14485,N_12581);
nor U17118 (N_17118,N_10427,N_11005);
nand U17119 (N_17119,N_11503,N_11322);
and U17120 (N_17120,N_12731,N_11229);
or U17121 (N_17121,N_13654,N_13255);
nor U17122 (N_17122,N_10504,N_14542);
or U17123 (N_17123,N_11058,N_11291);
or U17124 (N_17124,N_11510,N_14655);
xor U17125 (N_17125,N_10700,N_13965);
and U17126 (N_17126,N_12142,N_10322);
nand U17127 (N_17127,N_13769,N_12326);
nand U17128 (N_17128,N_13477,N_14364);
nor U17129 (N_17129,N_12813,N_14403);
xor U17130 (N_17130,N_11859,N_10764);
nor U17131 (N_17131,N_10884,N_11414);
or U17132 (N_17132,N_13277,N_11976);
and U17133 (N_17133,N_11102,N_12457);
or U17134 (N_17134,N_10388,N_12235);
or U17135 (N_17135,N_12503,N_13696);
or U17136 (N_17136,N_10421,N_13112);
and U17137 (N_17137,N_10399,N_12228);
nor U17138 (N_17138,N_11357,N_10845);
and U17139 (N_17139,N_12024,N_13135);
nand U17140 (N_17140,N_11998,N_12093);
and U17141 (N_17141,N_14619,N_13604);
or U17142 (N_17142,N_14894,N_12726);
nand U17143 (N_17143,N_14628,N_14414);
nand U17144 (N_17144,N_11865,N_11963);
and U17145 (N_17145,N_10577,N_12936);
xor U17146 (N_17146,N_10423,N_11697);
xnor U17147 (N_17147,N_14367,N_13139);
or U17148 (N_17148,N_12178,N_11136);
and U17149 (N_17149,N_13156,N_13519);
or U17150 (N_17150,N_13726,N_14205);
nand U17151 (N_17151,N_12390,N_12518);
xnor U17152 (N_17152,N_11155,N_14242);
xnor U17153 (N_17153,N_10168,N_13885);
nor U17154 (N_17154,N_11372,N_11858);
xor U17155 (N_17155,N_14183,N_12003);
nand U17156 (N_17156,N_11725,N_14885);
or U17157 (N_17157,N_10819,N_12084);
xor U17158 (N_17158,N_13465,N_11255);
nor U17159 (N_17159,N_10277,N_10063);
or U17160 (N_17160,N_13253,N_13297);
and U17161 (N_17161,N_11449,N_10126);
nand U17162 (N_17162,N_10826,N_12297);
nand U17163 (N_17163,N_13251,N_14552);
nor U17164 (N_17164,N_14536,N_13814);
nor U17165 (N_17165,N_13163,N_11550);
or U17166 (N_17166,N_12251,N_13295);
or U17167 (N_17167,N_11656,N_12261);
nor U17168 (N_17168,N_14411,N_14921);
or U17169 (N_17169,N_11847,N_11367);
or U17170 (N_17170,N_10174,N_11855);
nand U17171 (N_17171,N_11889,N_10363);
or U17172 (N_17172,N_12564,N_14770);
nor U17173 (N_17173,N_14794,N_14625);
or U17174 (N_17174,N_12418,N_10196);
nor U17175 (N_17175,N_14211,N_14046);
xor U17176 (N_17176,N_14622,N_10023);
nand U17177 (N_17177,N_10679,N_10338);
xnor U17178 (N_17178,N_11439,N_11261);
and U17179 (N_17179,N_11949,N_10224);
xnor U17180 (N_17180,N_11994,N_14262);
nor U17181 (N_17181,N_11818,N_13285);
or U17182 (N_17182,N_10052,N_13035);
nor U17183 (N_17183,N_11137,N_11811);
xor U17184 (N_17184,N_11193,N_11857);
nor U17185 (N_17185,N_10402,N_11522);
and U17186 (N_17186,N_13107,N_12052);
or U17187 (N_17187,N_13785,N_14130);
or U17188 (N_17188,N_10952,N_14695);
xnor U17189 (N_17189,N_13619,N_12745);
xor U17190 (N_17190,N_13210,N_11271);
or U17191 (N_17191,N_10860,N_13315);
xnor U17192 (N_17192,N_10394,N_11139);
nor U17193 (N_17193,N_12551,N_11290);
nor U17194 (N_17194,N_13083,N_13503);
or U17195 (N_17195,N_11657,N_11182);
nor U17196 (N_17196,N_10148,N_10959);
or U17197 (N_17197,N_12882,N_14076);
nor U17198 (N_17198,N_14105,N_12732);
nand U17199 (N_17199,N_14198,N_14344);
or U17200 (N_17200,N_11016,N_13459);
nand U17201 (N_17201,N_12628,N_10076);
nand U17202 (N_17202,N_10503,N_10670);
or U17203 (N_17203,N_11711,N_11166);
nor U17204 (N_17204,N_12316,N_13462);
and U17205 (N_17205,N_12079,N_14526);
nor U17206 (N_17206,N_12440,N_13532);
nand U17207 (N_17207,N_10024,N_11384);
or U17208 (N_17208,N_11523,N_11380);
or U17209 (N_17209,N_10077,N_11344);
and U17210 (N_17210,N_10119,N_13517);
xnor U17211 (N_17211,N_11965,N_11698);
xnor U17212 (N_17212,N_10818,N_14085);
and U17213 (N_17213,N_10027,N_13838);
or U17214 (N_17214,N_12295,N_14916);
nor U17215 (N_17215,N_11269,N_14078);
and U17216 (N_17216,N_11960,N_14565);
nor U17217 (N_17217,N_14954,N_11262);
nor U17218 (N_17218,N_10900,N_14876);
or U17219 (N_17219,N_11841,N_13854);
nand U17220 (N_17220,N_12090,N_12028);
xor U17221 (N_17221,N_10762,N_12839);
xnor U17222 (N_17222,N_12768,N_13262);
and U17223 (N_17223,N_11926,N_10625);
and U17224 (N_17224,N_10330,N_14307);
nand U17225 (N_17225,N_11828,N_11567);
or U17226 (N_17226,N_11793,N_12065);
xor U17227 (N_17227,N_10209,N_11129);
and U17228 (N_17228,N_13487,N_13457);
nand U17229 (N_17229,N_14186,N_10836);
nor U17230 (N_17230,N_13808,N_14115);
and U17231 (N_17231,N_13238,N_10292);
or U17232 (N_17232,N_10417,N_14112);
xnor U17233 (N_17233,N_13231,N_14418);
nor U17234 (N_17234,N_12597,N_13831);
nand U17235 (N_17235,N_12198,N_13323);
nand U17236 (N_17236,N_11520,N_11400);
or U17237 (N_17237,N_12414,N_11874);
and U17238 (N_17238,N_14926,N_11634);
nand U17239 (N_17239,N_12807,N_12149);
or U17240 (N_17240,N_11714,N_11770);
nand U17241 (N_17241,N_10195,N_11944);
or U17242 (N_17242,N_13559,N_13064);
nor U17243 (N_17243,N_13146,N_13347);
and U17244 (N_17244,N_14016,N_13982);
nor U17245 (N_17245,N_11343,N_14160);
nand U17246 (N_17246,N_10711,N_10611);
xor U17247 (N_17247,N_10543,N_12825);
xnor U17248 (N_17248,N_11073,N_13609);
nand U17249 (N_17249,N_12343,N_13111);
and U17250 (N_17250,N_13335,N_13496);
xor U17251 (N_17251,N_14164,N_14633);
xnor U17252 (N_17252,N_13795,N_10869);
xnor U17253 (N_17253,N_10589,N_12181);
or U17254 (N_17254,N_12357,N_14514);
and U17255 (N_17255,N_13721,N_14171);
nor U17256 (N_17256,N_11760,N_10036);
nor U17257 (N_17257,N_12300,N_12869);
xor U17258 (N_17258,N_14043,N_11473);
or U17259 (N_17259,N_12130,N_10571);
and U17260 (N_17260,N_12565,N_11748);
and U17261 (N_17261,N_11935,N_10201);
xor U17262 (N_17262,N_11581,N_12832);
nand U17263 (N_17263,N_14244,N_14201);
nor U17264 (N_17264,N_11548,N_11767);
nand U17265 (N_17265,N_14961,N_11514);
and U17266 (N_17266,N_14931,N_13535);
or U17267 (N_17267,N_11907,N_12233);
xor U17268 (N_17268,N_10848,N_14306);
nor U17269 (N_17269,N_14180,N_10343);
nor U17270 (N_17270,N_10173,N_13750);
nand U17271 (N_17271,N_14253,N_12327);
nand U17272 (N_17272,N_13004,N_13016);
xor U17273 (N_17273,N_10222,N_13936);
xnor U17274 (N_17274,N_10230,N_14128);
or U17275 (N_17275,N_12560,N_12076);
nand U17276 (N_17276,N_11345,N_12023);
or U17277 (N_17277,N_13703,N_13612);
nor U17278 (N_17278,N_12568,N_13869);
nor U17279 (N_17279,N_12400,N_14795);
xor U17280 (N_17280,N_14980,N_11099);
or U17281 (N_17281,N_12553,N_12537);
nor U17282 (N_17282,N_11025,N_13290);
xor U17283 (N_17283,N_11665,N_13976);
and U17284 (N_17284,N_13259,N_11002);
and U17285 (N_17285,N_11247,N_11630);
or U17286 (N_17286,N_12524,N_10117);
nor U17287 (N_17287,N_10693,N_11227);
or U17288 (N_17288,N_12738,N_10725);
and U17289 (N_17289,N_10593,N_13113);
nand U17290 (N_17290,N_13682,N_12599);
xor U17291 (N_17291,N_10606,N_11006);
nor U17292 (N_17292,N_14316,N_13574);
nand U17293 (N_17293,N_12892,N_11285);
xnor U17294 (N_17294,N_12541,N_14696);
xnor U17295 (N_17295,N_10261,N_11245);
nor U17296 (N_17296,N_12675,N_11533);
nand U17297 (N_17297,N_11082,N_13857);
nor U17298 (N_17298,N_14828,N_10856);
nor U17299 (N_17299,N_14556,N_10458);
nand U17300 (N_17300,N_12703,N_12383);
nor U17301 (N_17301,N_11556,N_13486);
nor U17302 (N_17302,N_10183,N_11210);
and U17303 (N_17303,N_12645,N_11171);
or U17304 (N_17304,N_13516,N_12281);
xor U17305 (N_17305,N_11593,N_14809);
nand U17306 (N_17306,N_11176,N_11870);
nor U17307 (N_17307,N_13012,N_14388);
xor U17308 (N_17308,N_13051,N_14257);
or U17309 (N_17309,N_13576,N_11241);
nand U17310 (N_17310,N_13445,N_11207);
and U17311 (N_17311,N_12759,N_11779);
xnor U17312 (N_17312,N_14766,N_11981);
nand U17313 (N_17313,N_12193,N_12268);
or U17314 (N_17314,N_10872,N_13056);
or U17315 (N_17315,N_12388,N_12844);
or U17316 (N_17316,N_11125,N_14325);
nand U17317 (N_17317,N_10652,N_14311);
xor U17318 (N_17318,N_11243,N_13594);
and U17319 (N_17319,N_12165,N_13923);
xor U17320 (N_17320,N_13572,N_14247);
nand U17321 (N_17321,N_11806,N_13699);
xnor U17322 (N_17322,N_11438,N_11307);
nor U17323 (N_17323,N_10632,N_10538);
nand U17324 (N_17324,N_14019,N_12721);
nand U17325 (N_17325,N_10802,N_10753);
nor U17326 (N_17326,N_11827,N_11457);
or U17327 (N_17327,N_12509,N_11838);
nor U17328 (N_17328,N_11629,N_10380);
nor U17329 (N_17329,N_11484,N_12371);
nand U17330 (N_17330,N_12195,N_10268);
nor U17331 (N_17331,N_11648,N_10921);
and U17332 (N_17332,N_11876,N_10381);
nor U17333 (N_17333,N_13053,N_13540);
or U17334 (N_17334,N_10264,N_10046);
nor U17335 (N_17335,N_10473,N_10081);
and U17336 (N_17336,N_11968,N_11028);
nand U17337 (N_17337,N_14731,N_10429);
and U17338 (N_17338,N_11448,N_12760);
or U17339 (N_17339,N_11173,N_13515);
nand U17340 (N_17340,N_13858,N_11370);
nor U17341 (N_17341,N_13870,N_13822);
nand U17342 (N_17342,N_10638,N_10976);
xnor U17343 (N_17343,N_11489,N_14156);
and U17344 (N_17344,N_13311,N_11302);
nor U17345 (N_17345,N_12210,N_11024);
or U17346 (N_17346,N_14474,N_12226);
or U17347 (N_17347,N_14969,N_12972);
and U17348 (N_17348,N_13361,N_10085);
or U17349 (N_17349,N_14842,N_13000);
or U17350 (N_17350,N_11076,N_10542);
nand U17351 (N_17351,N_11001,N_13145);
or U17352 (N_17352,N_12619,N_14653);
xnor U17353 (N_17353,N_10875,N_13389);
and U17354 (N_17354,N_12241,N_13119);
or U17355 (N_17355,N_14286,N_12795);
or U17356 (N_17356,N_11362,N_13819);
xnor U17357 (N_17357,N_10899,N_11671);
nor U17358 (N_17358,N_14884,N_10156);
nor U17359 (N_17359,N_14722,N_12797);
nor U17360 (N_17360,N_11446,N_11015);
nand U17361 (N_17361,N_12410,N_13637);
or U17362 (N_17362,N_11014,N_14748);
nand U17363 (N_17363,N_14584,N_10862);
xor U17364 (N_17364,N_12974,N_12929);
xor U17365 (N_17365,N_13514,N_11731);
or U17366 (N_17366,N_10282,N_14598);
nor U17367 (N_17367,N_11607,N_13758);
and U17368 (N_17368,N_12939,N_10694);
and U17369 (N_17369,N_10924,N_11586);
or U17370 (N_17370,N_10210,N_10279);
xnor U17371 (N_17371,N_13105,N_14294);
xnor U17372 (N_17372,N_14504,N_12459);
and U17373 (N_17373,N_10682,N_10806);
and U17374 (N_17374,N_12734,N_14861);
or U17375 (N_17375,N_11709,N_12334);
or U17376 (N_17376,N_11398,N_12480);
nor U17377 (N_17377,N_12227,N_14571);
and U17378 (N_17378,N_12358,N_10513);
xor U17379 (N_17379,N_14806,N_11602);
or U17380 (N_17380,N_12550,N_13429);
nand U17381 (N_17381,N_12298,N_14395);
nand U17382 (N_17382,N_14121,N_12828);
nand U17383 (N_17383,N_12751,N_11672);
xnor U17384 (N_17384,N_11431,N_14385);
nand U17385 (N_17385,N_14312,N_12618);
and U17386 (N_17386,N_10006,N_13953);
or U17387 (N_17387,N_13177,N_13419);
and U17388 (N_17388,N_10519,N_14544);
and U17389 (N_17389,N_13733,N_11782);
nand U17390 (N_17390,N_14359,N_12610);
nor U17391 (N_17391,N_11347,N_11217);
or U17392 (N_17392,N_14002,N_11551);
nor U17393 (N_17393,N_11684,N_14887);
xnor U17394 (N_17394,N_10443,N_13197);
or U17395 (N_17395,N_10925,N_13110);
or U17396 (N_17396,N_10357,N_12054);
nand U17397 (N_17397,N_13191,N_11495);
nor U17398 (N_17398,N_14195,N_14708);
xor U17399 (N_17399,N_11878,N_11832);
xor U17400 (N_17400,N_11924,N_14750);
nor U17401 (N_17401,N_14412,N_13524);
xnor U17402 (N_17402,N_12128,N_11225);
or U17403 (N_17403,N_13889,N_10893);
and U17404 (N_17404,N_11951,N_13876);
or U17405 (N_17405,N_10907,N_10481);
xnor U17406 (N_17406,N_14691,N_13195);
xnor U17407 (N_17407,N_12366,N_14801);
xor U17408 (N_17408,N_12110,N_12424);
nand U17409 (N_17409,N_11404,N_14005);
nor U17410 (N_17410,N_10761,N_12644);
and U17411 (N_17411,N_14222,N_14651);
nor U17412 (N_17412,N_14690,N_10269);
xnor U17413 (N_17413,N_13525,N_12124);
and U17414 (N_17414,N_13435,N_13140);
xnor U17415 (N_17415,N_10635,N_13700);
or U17416 (N_17416,N_10345,N_11324);
nor U17417 (N_17417,N_10780,N_10964);
xnor U17418 (N_17418,N_13922,N_11912);
xor U17419 (N_17419,N_14454,N_11512);
or U17420 (N_17420,N_13374,N_10479);
nand U17421 (N_17421,N_10002,N_10500);
or U17422 (N_17422,N_14292,N_10091);
and U17423 (N_17423,N_13399,N_14082);
nand U17424 (N_17424,N_13741,N_14324);
nor U17425 (N_17425,N_14654,N_11046);
and U17426 (N_17426,N_13701,N_10502);
nand U17427 (N_17427,N_14479,N_13801);
nand U17428 (N_17428,N_14836,N_13100);
nor U17429 (N_17429,N_11194,N_10792);
nor U17430 (N_17430,N_13640,N_11293);
and U17431 (N_17431,N_10194,N_10214);
or U17432 (N_17432,N_14527,N_13108);
nor U17433 (N_17433,N_11950,N_14147);
nor U17434 (N_17434,N_13338,N_14759);
nor U17435 (N_17435,N_14777,N_13336);
nand U17436 (N_17436,N_10266,N_12212);
nor U17437 (N_17437,N_10938,N_12427);
xnor U17438 (N_17438,N_12935,N_14143);
or U17439 (N_17439,N_10386,N_10433);
nand U17440 (N_17440,N_10373,N_11143);
nor U17441 (N_17441,N_11141,N_14703);
nor U17442 (N_17442,N_14267,N_11460);
and U17443 (N_17443,N_10372,N_12752);
xor U17444 (N_17444,N_11211,N_11712);
or U17445 (N_17445,N_12749,N_14507);
nor U17446 (N_17446,N_10689,N_14405);
xor U17447 (N_17447,N_11464,N_11596);
or U17448 (N_17448,N_13484,N_12908);
and U17449 (N_17449,N_11904,N_13344);
or U17450 (N_17450,N_13932,N_11440);
xnor U17451 (N_17451,N_14857,N_12098);
nand U17452 (N_17452,N_11428,N_14911);
and U17453 (N_17453,N_13175,N_10351);
or U17454 (N_17454,N_13416,N_12862);
nand U17455 (N_17455,N_11259,N_13203);
or U17456 (N_17456,N_11877,N_11204);
or U17457 (N_17457,N_13380,N_14248);
and U17458 (N_17458,N_12017,N_14057);
or U17459 (N_17459,N_13324,N_10065);
and U17460 (N_17460,N_13731,N_10025);
nor U17461 (N_17461,N_13676,N_14682);
nand U17462 (N_17462,N_10460,N_12283);
nor U17463 (N_17463,N_11043,N_12263);
or U17464 (N_17464,N_14736,N_13820);
nand U17465 (N_17465,N_10843,N_12450);
nand U17466 (N_17466,N_11746,N_10154);
xnor U17467 (N_17467,N_10256,N_13043);
xor U17468 (N_17468,N_13647,N_12859);
nor U17469 (N_17469,N_13155,N_13848);
nor U17470 (N_17470,N_10808,N_10847);
and U17471 (N_17471,N_13691,N_11902);
or U17472 (N_17472,N_11369,N_11539);
nand U17473 (N_17473,N_12580,N_12035);
nand U17474 (N_17474,N_14614,N_13325);
nor U17475 (N_17475,N_14416,N_10715);
xor U17476 (N_17476,N_11349,N_14570);
and U17477 (N_17477,N_11236,N_14630);
and U17478 (N_17478,N_13837,N_10494);
xnor U17479 (N_17479,N_14575,N_10492);
or U17480 (N_17480,N_13369,N_14549);
xnor U17481 (N_17481,N_10074,N_11321);
nand U17482 (N_17482,N_10087,N_11277);
nand U17483 (N_17483,N_11961,N_13433);
or U17484 (N_17484,N_11872,N_12937);
nand U17485 (N_17485,N_14693,N_12367);
or U17486 (N_17486,N_14937,N_12608);
xor U17487 (N_17487,N_12047,N_14904);
and U17488 (N_17488,N_14001,N_13621);
nor U17489 (N_17489,N_14035,N_10627);
nor U17490 (N_17490,N_11873,N_12490);
nor U17491 (N_17491,N_14004,N_12979);
and U17492 (N_17492,N_11555,N_10665);
or U17493 (N_17493,N_13566,N_10812);
nand U17494 (N_17494,N_12769,N_11042);
nand U17495 (N_17495,N_13972,N_14909);
nand U17496 (N_17496,N_10936,N_12669);
nor U17497 (N_17497,N_13327,N_11913);
and U17498 (N_17498,N_13849,N_12926);
nor U17499 (N_17499,N_14390,N_11476);
and U17500 (N_17500,N_14975,N_10418);
nor U17501 (N_17501,N_11104,N_11467);
nand U17502 (N_17502,N_11985,N_12412);
or U17503 (N_17503,N_14400,N_10421);
nand U17504 (N_17504,N_10498,N_11790);
nor U17505 (N_17505,N_10138,N_12871);
xnor U17506 (N_17506,N_10136,N_14681);
xor U17507 (N_17507,N_14857,N_10964);
nor U17508 (N_17508,N_12272,N_12990);
nor U17509 (N_17509,N_11214,N_14213);
or U17510 (N_17510,N_10601,N_12882);
nor U17511 (N_17511,N_13252,N_10819);
nor U17512 (N_17512,N_13415,N_14835);
nand U17513 (N_17513,N_13307,N_13821);
xor U17514 (N_17514,N_12272,N_12740);
or U17515 (N_17515,N_13092,N_11755);
or U17516 (N_17516,N_10497,N_13844);
nor U17517 (N_17517,N_10683,N_14239);
or U17518 (N_17518,N_13804,N_11054);
and U17519 (N_17519,N_10451,N_12259);
or U17520 (N_17520,N_11497,N_10838);
nand U17521 (N_17521,N_14247,N_14593);
or U17522 (N_17522,N_10442,N_14837);
nor U17523 (N_17523,N_13859,N_11729);
nor U17524 (N_17524,N_14980,N_10596);
xor U17525 (N_17525,N_14020,N_14392);
and U17526 (N_17526,N_13312,N_11405);
and U17527 (N_17527,N_12811,N_11550);
xor U17528 (N_17528,N_10487,N_13729);
nand U17529 (N_17529,N_12830,N_12927);
nand U17530 (N_17530,N_14559,N_12725);
nand U17531 (N_17531,N_13237,N_13725);
xor U17532 (N_17532,N_14499,N_13959);
xor U17533 (N_17533,N_12580,N_11492);
or U17534 (N_17534,N_12682,N_11725);
or U17535 (N_17535,N_13995,N_14248);
nand U17536 (N_17536,N_13145,N_12053);
and U17537 (N_17537,N_14010,N_13212);
xor U17538 (N_17538,N_12231,N_14942);
nor U17539 (N_17539,N_13518,N_11226);
nor U17540 (N_17540,N_10147,N_13248);
nor U17541 (N_17541,N_11712,N_14569);
nor U17542 (N_17542,N_14321,N_12370);
or U17543 (N_17543,N_13024,N_12502);
nand U17544 (N_17544,N_10855,N_12609);
nor U17545 (N_17545,N_11349,N_13171);
and U17546 (N_17546,N_10105,N_14629);
or U17547 (N_17547,N_11939,N_10104);
xnor U17548 (N_17548,N_13694,N_10141);
xor U17549 (N_17549,N_12353,N_12989);
nand U17550 (N_17550,N_14635,N_10505);
and U17551 (N_17551,N_10475,N_14313);
nand U17552 (N_17552,N_14448,N_10811);
and U17553 (N_17553,N_10014,N_12569);
or U17554 (N_17554,N_12898,N_14262);
xnor U17555 (N_17555,N_12460,N_11000);
or U17556 (N_17556,N_13401,N_10646);
xnor U17557 (N_17557,N_11770,N_14628);
or U17558 (N_17558,N_13259,N_12074);
and U17559 (N_17559,N_12282,N_12527);
nand U17560 (N_17560,N_14034,N_10960);
nor U17561 (N_17561,N_10286,N_12450);
xor U17562 (N_17562,N_11982,N_11948);
xnor U17563 (N_17563,N_11380,N_12113);
or U17564 (N_17564,N_11029,N_13292);
nor U17565 (N_17565,N_13295,N_11471);
and U17566 (N_17566,N_12200,N_14613);
xor U17567 (N_17567,N_12655,N_13388);
or U17568 (N_17568,N_12194,N_13075);
or U17569 (N_17569,N_10528,N_10601);
nand U17570 (N_17570,N_11373,N_12781);
and U17571 (N_17571,N_13315,N_11442);
nor U17572 (N_17572,N_13239,N_14852);
nor U17573 (N_17573,N_10350,N_10902);
and U17574 (N_17574,N_10574,N_12866);
and U17575 (N_17575,N_14657,N_14812);
nor U17576 (N_17576,N_14473,N_13493);
and U17577 (N_17577,N_12351,N_10071);
and U17578 (N_17578,N_14897,N_12662);
or U17579 (N_17579,N_14811,N_14329);
or U17580 (N_17580,N_13446,N_13706);
nand U17581 (N_17581,N_13382,N_13453);
and U17582 (N_17582,N_10773,N_12307);
nor U17583 (N_17583,N_14573,N_14928);
and U17584 (N_17584,N_10722,N_13687);
xor U17585 (N_17585,N_14989,N_12385);
or U17586 (N_17586,N_14035,N_13931);
nor U17587 (N_17587,N_10538,N_12595);
or U17588 (N_17588,N_13585,N_10866);
xnor U17589 (N_17589,N_11374,N_14372);
xor U17590 (N_17590,N_10255,N_13306);
xnor U17591 (N_17591,N_10185,N_13347);
nor U17592 (N_17592,N_12436,N_12491);
nor U17593 (N_17593,N_11223,N_13517);
nand U17594 (N_17594,N_14813,N_11844);
nand U17595 (N_17595,N_12218,N_10142);
xor U17596 (N_17596,N_13324,N_12920);
and U17597 (N_17597,N_12151,N_13550);
or U17598 (N_17598,N_13690,N_12736);
and U17599 (N_17599,N_12648,N_13467);
or U17600 (N_17600,N_11701,N_14460);
and U17601 (N_17601,N_14193,N_10910);
xnor U17602 (N_17602,N_10175,N_14036);
nand U17603 (N_17603,N_11184,N_13826);
nor U17604 (N_17604,N_12178,N_14553);
and U17605 (N_17605,N_11488,N_10042);
and U17606 (N_17606,N_13985,N_12460);
nand U17607 (N_17607,N_14163,N_10440);
and U17608 (N_17608,N_11013,N_13175);
xnor U17609 (N_17609,N_12849,N_14153);
or U17610 (N_17610,N_13443,N_11895);
nor U17611 (N_17611,N_14801,N_14222);
or U17612 (N_17612,N_12479,N_10863);
nor U17613 (N_17613,N_11788,N_14079);
nand U17614 (N_17614,N_14583,N_10282);
and U17615 (N_17615,N_10902,N_14602);
xnor U17616 (N_17616,N_10189,N_14821);
nand U17617 (N_17617,N_13719,N_12337);
or U17618 (N_17618,N_10515,N_12868);
nor U17619 (N_17619,N_11499,N_10550);
xnor U17620 (N_17620,N_10587,N_13249);
and U17621 (N_17621,N_10685,N_13745);
xor U17622 (N_17622,N_10202,N_11553);
nand U17623 (N_17623,N_11033,N_12328);
and U17624 (N_17624,N_14981,N_12652);
nand U17625 (N_17625,N_14673,N_13774);
nand U17626 (N_17626,N_10374,N_14292);
xnor U17627 (N_17627,N_14558,N_10751);
nor U17628 (N_17628,N_11097,N_10894);
nand U17629 (N_17629,N_10560,N_14851);
nand U17630 (N_17630,N_14096,N_11257);
or U17631 (N_17631,N_13882,N_11956);
and U17632 (N_17632,N_11859,N_14169);
nor U17633 (N_17633,N_14841,N_11323);
nor U17634 (N_17634,N_14078,N_13213);
nor U17635 (N_17635,N_14172,N_11460);
nand U17636 (N_17636,N_10234,N_13105);
xor U17637 (N_17637,N_12939,N_12322);
nor U17638 (N_17638,N_12151,N_14738);
xor U17639 (N_17639,N_12885,N_14622);
nand U17640 (N_17640,N_14749,N_11417);
nand U17641 (N_17641,N_10848,N_11198);
nor U17642 (N_17642,N_12785,N_10950);
and U17643 (N_17643,N_11817,N_14817);
nor U17644 (N_17644,N_13765,N_11829);
or U17645 (N_17645,N_12812,N_13626);
nor U17646 (N_17646,N_11574,N_13278);
or U17647 (N_17647,N_10075,N_11182);
or U17648 (N_17648,N_14258,N_11339);
nor U17649 (N_17649,N_12354,N_13998);
or U17650 (N_17650,N_12936,N_10608);
nor U17651 (N_17651,N_10492,N_10029);
xnor U17652 (N_17652,N_14638,N_12416);
nor U17653 (N_17653,N_11820,N_10536);
xnor U17654 (N_17654,N_11714,N_14936);
xor U17655 (N_17655,N_12917,N_13311);
or U17656 (N_17656,N_11892,N_12291);
xnor U17657 (N_17657,N_13586,N_13108);
or U17658 (N_17658,N_10108,N_13485);
nor U17659 (N_17659,N_14346,N_10163);
nand U17660 (N_17660,N_12010,N_12239);
and U17661 (N_17661,N_10169,N_14143);
nand U17662 (N_17662,N_12628,N_11842);
xor U17663 (N_17663,N_13606,N_11321);
and U17664 (N_17664,N_14459,N_10329);
and U17665 (N_17665,N_12210,N_14687);
and U17666 (N_17666,N_13925,N_10214);
xor U17667 (N_17667,N_10913,N_12769);
nand U17668 (N_17668,N_10247,N_14756);
and U17669 (N_17669,N_12597,N_13892);
or U17670 (N_17670,N_14651,N_11470);
and U17671 (N_17671,N_12701,N_12684);
xor U17672 (N_17672,N_10034,N_10060);
nor U17673 (N_17673,N_14467,N_12298);
nand U17674 (N_17674,N_12875,N_13398);
xnor U17675 (N_17675,N_13553,N_10826);
nand U17676 (N_17676,N_10005,N_14893);
or U17677 (N_17677,N_13999,N_13154);
and U17678 (N_17678,N_12229,N_14029);
and U17679 (N_17679,N_12092,N_12686);
xnor U17680 (N_17680,N_14154,N_14928);
and U17681 (N_17681,N_11294,N_10299);
or U17682 (N_17682,N_11044,N_11132);
nand U17683 (N_17683,N_14590,N_11240);
nor U17684 (N_17684,N_11893,N_12766);
nor U17685 (N_17685,N_13026,N_12125);
xor U17686 (N_17686,N_14049,N_11819);
xnor U17687 (N_17687,N_13045,N_12700);
xor U17688 (N_17688,N_14258,N_10100);
nor U17689 (N_17689,N_13593,N_13135);
and U17690 (N_17690,N_13506,N_10262);
or U17691 (N_17691,N_14494,N_11857);
xor U17692 (N_17692,N_10653,N_13544);
or U17693 (N_17693,N_14536,N_13955);
nor U17694 (N_17694,N_12268,N_11984);
xor U17695 (N_17695,N_12133,N_10946);
nor U17696 (N_17696,N_13607,N_10921);
xnor U17697 (N_17697,N_14565,N_10636);
xnor U17698 (N_17698,N_12072,N_14937);
xor U17699 (N_17699,N_10815,N_13566);
nand U17700 (N_17700,N_13010,N_13483);
and U17701 (N_17701,N_10726,N_12506);
nand U17702 (N_17702,N_12593,N_12427);
nand U17703 (N_17703,N_10007,N_14212);
or U17704 (N_17704,N_10120,N_11145);
xnor U17705 (N_17705,N_14798,N_13581);
nor U17706 (N_17706,N_14597,N_11461);
xnor U17707 (N_17707,N_14652,N_11248);
nor U17708 (N_17708,N_14234,N_13866);
and U17709 (N_17709,N_13172,N_13109);
or U17710 (N_17710,N_13770,N_14031);
or U17711 (N_17711,N_11880,N_14291);
or U17712 (N_17712,N_12364,N_14632);
or U17713 (N_17713,N_13654,N_11067);
or U17714 (N_17714,N_14065,N_13434);
or U17715 (N_17715,N_12048,N_10436);
xnor U17716 (N_17716,N_10231,N_11990);
nor U17717 (N_17717,N_10849,N_10548);
nor U17718 (N_17718,N_13117,N_10593);
and U17719 (N_17719,N_11591,N_11496);
or U17720 (N_17720,N_13209,N_13642);
xnor U17721 (N_17721,N_14233,N_14764);
or U17722 (N_17722,N_12096,N_13723);
or U17723 (N_17723,N_12777,N_10838);
and U17724 (N_17724,N_14530,N_10049);
and U17725 (N_17725,N_14814,N_10953);
or U17726 (N_17726,N_12207,N_14281);
and U17727 (N_17727,N_12660,N_10047);
nor U17728 (N_17728,N_11262,N_11675);
and U17729 (N_17729,N_10102,N_11483);
nor U17730 (N_17730,N_12057,N_14583);
xor U17731 (N_17731,N_12393,N_10723);
nor U17732 (N_17732,N_14412,N_12659);
nor U17733 (N_17733,N_11819,N_10135);
nand U17734 (N_17734,N_13407,N_11514);
or U17735 (N_17735,N_12495,N_12030);
nor U17736 (N_17736,N_14634,N_11337);
xor U17737 (N_17737,N_11883,N_11851);
and U17738 (N_17738,N_10351,N_11223);
and U17739 (N_17739,N_12020,N_11848);
nand U17740 (N_17740,N_10595,N_13201);
nand U17741 (N_17741,N_13885,N_10807);
xnor U17742 (N_17742,N_12536,N_12478);
or U17743 (N_17743,N_13877,N_12382);
or U17744 (N_17744,N_12493,N_12014);
or U17745 (N_17745,N_14414,N_12077);
or U17746 (N_17746,N_11092,N_14898);
nor U17747 (N_17747,N_13244,N_13342);
xor U17748 (N_17748,N_11933,N_10755);
or U17749 (N_17749,N_10880,N_11992);
nor U17750 (N_17750,N_14825,N_10483);
nand U17751 (N_17751,N_14003,N_14698);
or U17752 (N_17752,N_14263,N_12453);
xnor U17753 (N_17753,N_11023,N_10253);
nand U17754 (N_17754,N_12102,N_14547);
or U17755 (N_17755,N_13758,N_12093);
and U17756 (N_17756,N_13083,N_10459);
and U17757 (N_17757,N_13774,N_12013);
nor U17758 (N_17758,N_13101,N_14594);
nor U17759 (N_17759,N_10805,N_12103);
xnor U17760 (N_17760,N_13992,N_12008);
xnor U17761 (N_17761,N_10861,N_14883);
and U17762 (N_17762,N_10620,N_12320);
xor U17763 (N_17763,N_11771,N_14907);
nor U17764 (N_17764,N_13019,N_10112);
or U17765 (N_17765,N_14290,N_13349);
nand U17766 (N_17766,N_10539,N_11768);
and U17767 (N_17767,N_10334,N_11879);
xor U17768 (N_17768,N_13546,N_10038);
nand U17769 (N_17769,N_10041,N_11836);
and U17770 (N_17770,N_12742,N_11450);
or U17771 (N_17771,N_13828,N_13832);
nand U17772 (N_17772,N_13322,N_14444);
nor U17773 (N_17773,N_11407,N_14449);
or U17774 (N_17774,N_11626,N_11177);
nand U17775 (N_17775,N_11383,N_11856);
nor U17776 (N_17776,N_13869,N_13604);
or U17777 (N_17777,N_11731,N_12638);
nand U17778 (N_17778,N_10432,N_11326);
nor U17779 (N_17779,N_14814,N_11794);
xnor U17780 (N_17780,N_10310,N_13313);
xnor U17781 (N_17781,N_13948,N_12806);
nand U17782 (N_17782,N_11995,N_14719);
nand U17783 (N_17783,N_13887,N_11131);
and U17784 (N_17784,N_14248,N_11616);
nand U17785 (N_17785,N_10324,N_14825);
or U17786 (N_17786,N_11674,N_11593);
and U17787 (N_17787,N_11713,N_12234);
nor U17788 (N_17788,N_13364,N_10045);
nand U17789 (N_17789,N_12810,N_14710);
and U17790 (N_17790,N_13244,N_14910);
xnor U17791 (N_17791,N_12962,N_11964);
nor U17792 (N_17792,N_13412,N_11079);
nand U17793 (N_17793,N_12633,N_13855);
nand U17794 (N_17794,N_11477,N_11030);
and U17795 (N_17795,N_13863,N_13199);
or U17796 (N_17796,N_10455,N_10541);
nand U17797 (N_17797,N_13642,N_13315);
nor U17798 (N_17798,N_14514,N_10663);
and U17799 (N_17799,N_11609,N_12806);
nand U17800 (N_17800,N_14590,N_11288);
nand U17801 (N_17801,N_13637,N_12903);
nand U17802 (N_17802,N_13718,N_13585);
nand U17803 (N_17803,N_13098,N_12441);
xor U17804 (N_17804,N_14464,N_14129);
and U17805 (N_17805,N_11361,N_11513);
nor U17806 (N_17806,N_10953,N_11681);
nor U17807 (N_17807,N_13358,N_10346);
nor U17808 (N_17808,N_13713,N_12962);
or U17809 (N_17809,N_11161,N_13126);
nor U17810 (N_17810,N_12659,N_10232);
nand U17811 (N_17811,N_14244,N_14538);
xnor U17812 (N_17812,N_12195,N_13879);
nand U17813 (N_17813,N_14416,N_10903);
or U17814 (N_17814,N_10432,N_11041);
nor U17815 (N_17815,N_10404,N_13271);
and U17816 (N_17816,N_13020,N_13161);
nand U17817 (N_17817,N_14591,N_14753);
nor U17818 (N_17818,N_11350,N_12979);
or U17819 (N_17819,N_11836,N_11424);
and U17820 (N_17820,N_12277,N_12634);
or U17821 (N_17821,N_12974,N_13478);
nand U17822 (N_17822,N_13005,N_11431);
nor U17823 (N_17823,N_12979,N_11266);
or U17824 (N_17824,N_12677,N_14951);
or U17825 (N_17825,N_12911,N_11863);
xor U17826 (N_17826,N_14463,N_10181);
and U17827 (N_17827,N_12903,N_13901);
and U17828 (N_17828,N_14869,N_13310);
and U17829 (N_17829,N_14161,N_11602);
nor U17830 (N_17830,N_10084,N_14861);
and U17831 (N_17831,N_14576,N_12386);
xor U17832 (N_17832,N_10617,N_14883);
or U17833 (N_17833,N_13356,N_10622);
nand U17834 (N_17834,N_11056,N_14961);
nand U17835 (N_17835,N_14562,N_12732);
and U17836 (N_17836,N_11612,N_11826);
nor U17837 (N_17837,N_13400,N_11562);
xnor U17838 (N_17838,N_14660,N_13248);
xor U17839 (N_17839,N_12301,N_12898);
nand U17840 (N_17840,N_11606,N_10417);
nand U17841 (N_17841,N_11220,N_12655);
and U17842 (N_17842,N_10073,N_12715);
nor U17843 (N_17843,N_14236,N_12503);
nor U17844 (N_17844,N_14253,N_10748);
and U17845 (N_17845,N_14925,N_14160);
or U17846 (N_17846,N_11482,N_11913);
and U17847 (N_17847,N_13825,N_14026);
and U17848 (N_17848,N_13855,N_11298);
xnor U17849 (N_17849,N_14027,N_13890);
and U17850 (N_17850,N_12992,N_13656);
xnor U17851 (N_17851,N_10959,N_12307);
xnor U17852 (N_17852,N_12253,N_12325);
nor U17853 (N_17853,N_10267,N_12226);
nor U17854 (N_17854,N_12771,N_12973);
xnor U17855 (N_17855,N_14721,N_13657);
xnor U17856 (N_17856,N_13805,N_14126);
nand U17857 (N_17857,N_11507,N_13367);
and U17858 (N_17858,N_11177,N_14050);
and U17859 (N_17859,N_13699,N_11233);
nand U17860 (N_17860,N_10307,N_14564);
nand U17861 (N_17861,N_13275,N_14072);
or U17862 (N_17862,N_12772,N_10650);
or U17863 (N_17863,N_13358,N_11963);
nor U17864 (N_17864,N_11878,N_14805);
nor U17865 (N_17865,N_11208,N_14045);
and U17866 (N_17866,N_14020,N_11868);
or U17867 (N_17867,N_14358,N_14230);
or U17868 (N_17868,N_14499,N_12189);
xnor U17869 (N_17869,N_12231,N_13117);
nor U17870 (N_17870,N_14944,N_14216);
nor U17871 (N_17871,N_11691,N_14551);
nand U17872 (N_17872,N_14491,N_12061);
xor U17873 (N_17873,N_10807,N_11494);
nor U17874 (N_17874,N_11258,N_11058);
xnor U17875 (N_17875,N_12421,N_14623);
xnor U17876 (N_17876,N_14967,N_10158);
nand U17877 (N_17877,N_11883,N_13266);
or U17878 (N_17878,N_11419,N_10097);
nand U17879 (N_17879,N_11114,N_14970);
nand U17880 (N_17880,N_13171,N_10015);
or U17881 (N_17881,N_12633,N_12597);
and U17882 (N_17882,N_12963,N_11047);
nand U17883 (N_17883,N_12105,N_10686);
or U17884 (N_17884,N_13157,N_13111);
nand U17885 (N_17885,N_13837,N_12079);
and U17886 (N_17886,N_12532,N_13397);
or U17887 (N_17887,N_11259,N_13020);
nor U17888 (N_17888,N_12277,N_12256);
or U17889 (N_17889,N_14631,N_14065);
xor U17890 (N_17890,N_10566,N_10158);
xor U17891 (N_17891,N_10186,N_14585);
xor U17892 (N_17892,N_13403,N_13580);
and U17893 (N_17893,N_14494,N_10869);
xor U17894 (N_17894,N_13951,N_13596);
nor U17895 (N_17895,N_11424,N_14051);
nand U17896 (N_17896,N_12597,N_13071);
nand U17897 (N_17897,N_13748,N_10005);
or U17898 (N_17898,N_10690,N_13826);
nand U17899 (N_17899,N_12340,N_11966);
xor U17900 (N_17900,N_13989,N_13992);
and U17901 (N_17901,N_11319,N_12088);
xnor U17902 (N_17902,N_10866,N_12861);
and U17903 (N_17903,N_13445,N_11110);
or U17904 (N_17904,N_12458,N_14277);
xnor U17905 (N_17905,N_13842,N_14554);
xor U17906 (N_17906,N_11142,N_11975);
xnor U17907 (N_17907,N_10788,N_10883);
nand U17908 (N_17908,N_11765,N_13114);
xor U17909 (N_17909,N_12075,N_12077);
xnor U17910 (N_17910,N_12802,N_11988);
or U17911 (N_17911,N_14695,N_13809);
nand U17912 (N_17912,N_12660,N_13744);
and U17913 (N_17913,N_10796,N_14408);
nand U17914 (N_17914,N_10896,N_10939);
xnor U17915 (N_17915,N_12822,N_11617);
nand U17916 (N_17916,N_10469,N_14556);
xor U17917 (N_17917,N_14828,N_13823);
and U17918 (N_17918,N_13787,N_12252);
and U17919 (N_17919,N_12685,N_13172);
xor U17920 (N_17920,N_13351,N_11825);
nand U17921 (N_17921,N_14792,N_10717);
xor U17922 (N_17922,N_13386,N_13691);
or U17923 (N_17923,N_12276,N_10386);
xnor U17924 (N_17924,N_11244,N_11902);
or U17925 (N_17925,N_10983,N_11236);
nor U17926 (N_17926,N_11511,N_12893);
nor U17927 (N_17927,N_10897,N_13322);
and U17928 (N_17928,N_13618,N_10290);
nor U17929 (N_17929,N_12552,N_12191);
and U17930 (N_17930,N_14585,N_13669);
or U17931 (N_17931,N_10051,N_10894);
nor U17932 (N_17932,N_14157,N_11144);
nand U17933 (N_17933,N_13327,N_10477);
nor U17934 (N_17934,N_13400,N_11638);
or U17935 (N_17935,N_12122,N_14994);
nor U17936 (N_17936,N_12999,N_14475);
or U17937 (N_17937,N_13265,N_13604);
nand U17938 (N_17938,N_12308,N_13299);
nand U17939 (N_17939,N_14557,N_10190);
nor U17940 (N_17940,N_11766,N_11666);
nor U17941 (N_17941,N_10493,N_10447);
xnor U17942 (N_17942,N_13151,N_10798);
xnor U17943 (N_17943,N_10636,N_11184);
or U17944 (N_17944,N_11913,N_12187);
or U17945 (N_17945,N_12731,N_12047);
xor U17946 (N_17946,N_12544,N_12244);
nand U17947 (N_17947,N_11704,N_11368);
or U17948 (N_17948,N_12700,N_13598);
xnor U17949 (N_17949,N_12517,N_11933);
and U17950 (N_17950,N_11190,N_12631);
nand U17951 (N_17951,N_14804,N_11949);
and U17952 (N_17952,N_11073,N_10570);
xnor U17953 (N_17953,N_14258,N_10402);
and U17954 (N_17954,N_10661,N_10527);
nand U17955 (N_17955,N_14657,N_12184);
or U17956 (N_17956,N_10416,N_12344);
or U17957 (N_17957,N_14751,N_12231);
or U17958 (N_17958,N_12714,N_11203);
or U17959 (N_17959,N_10489,N_10382);
and U17960 (N_17960,N_11839,N_13905);
and U17961 (N_17961,N_14004,N_13779);
or U17962 (N_17962,N_13420,N_14793);
xor U17963 (N_17963,N_10166,N_13820);
and U17964 (N_17964,N_13948,N_11966);
xor U17965 (N_17965,N_14237,N_14679);
and U17966 (N_17966,N_13591,N_10840);
and U17967 (N_17967,N_12318,N_11382);
or U17968 (N_17968,N_10866,N_14344);
nand U17969 (N_17969,N_12315,N_12727);
xor U17970 (N_17970,N_12459,N_13950);
and U17971 (N_17971,N_14215,N_11028);
or U17972 (N_17972,N_13174,N_11867);
or U17973 (N_17973,N_13423,N_14136);
nor U17974 (N_17974,N_12074,N_10568);
and U17975 (N_17975,N_13956,N_11969);
nor U17976 (N_17976,N_12927,N_10542);
and U17977 (N_17977,N_13311,N_12073);
and U17978 (N_17978,N_12379,N_13102);
nor U17979 (N_17979,N_12358,N_13119);
nand U17980 (N_17980,N_14271,N_14282);
nand U17981 (N_17981,N_11330,N_13584);
xor U17982 (N_17982,N_12305,N_13687);
and U17983 (N_17983,N_12884,N_10131);
xnor U17984 (N_17984,N_13407,N_10735);
nand U17985 (N_17985,N_10742,N_13074);
or U17986 (N_17986,N_14453,N_14491);
or U17987 (N_17987,N_12083,N_10864);
nor U17988 (N_17988,N_13529,N_11451);
and U17989 (N_17989,N_12265,N_12213);
nor U17990 (N_17990,N_14676,N_14272);
xor U17991 (N_17991,N_11218,N_14314);
nor U17992 (N_17992,N_10895,N_11543);
nand U17993 (N_17993,N_10234,N_13798);
xnor U17994 (N_17994,N_10636,N_12393);
nand U17995 (N_17995,N_14172,N_12966);
or U17996 (N_17996,N_14196,N_10084);
xnor U17997 (N_17997,N_11279,N_13147);
or U17998 (N_17998,N_10105,N_13533);
nand U17999 (N_17999,N_13820,N_12937);
nor U18000 (N_18000,N_11795,N_12077);
nor U18001 (N_18001,N_13235,N_14301);
xnor U18002 (N_18002,N_11599,N_13067);
and U18003 (N_18003,N_14977,N_12616);
nand U18004 (N_18004,N_13967,N_14859);
xor U18005 (N_18005,N_10176,N_11087);
or U18006 (N_18006,N_14762,N_14436);
nor U18007 (N_18007,N_11415,N_13768);
or U18008 (N_18008,N_13786,N_14078);
xnor U18009 (N_18009,N_13961,N_13302);
nand U18010 (N_18010,N_12314,N_13051);
or U18011 (N_18011,N_14236,N_11666);
xnor U18012 (N_18012,N_13391,N_10393);
xor U18013 (N_18013,N_12537,N_14453);
and U18014 (N_18014,N_12130,N_13673);
nor U18015 (N_18015,N_10579,N_10386);
and U18016 (N_18016,N_13220,N_10211);
or U18017 (N_18017,N_13313,N_10249);
nor U18018 (N_18018,N_11555,N_10835);
and U18019 (N_18019,N_10451,N_10686);
xnor U18020 (N_18020,N_12266,N_13830);
nand U18021 (N_18021,N_14598,N_14992);
nand U18022 (N_18022,N_11331,N_11421);
and U18023 (N_18023,N_12377,N_14708);
nand U18024 (N_18024,N_11012,N_11291);
xor U18025 (N_18025,N_10008,N_13402);
or U18026 (N_18026,N_10843,N_12527);
xnor U18027 (N_18027,N_12146,N_11138);
xor U18028 (N_18028,N_14729,N_13425);
nand U18029 (N_18029,N_10333,N_14023);
xnor U18030 (N_18030,N_14069,N_11858);
nand U18031 (N_18031,N_10122,N_12201);
or U18032 (N_18032,N_11899,N_12869);
xor U18033 (N_18033,N_11728,N_10387);
and U18034 (N_18034,N_10639,N_13121);
nand U18035 (N_18035,N_13142,N_10358);
xor U18036 (N_18036,N_12325,N_14140);
xor U18037 (N_18037,N_10641,N_11137);
xor U18038 (N_18038,N_10843,N_11745);
nor U18039 (N_18039,N_14757,N_14645);
nor U18040 (N_18040,N_11764,N_10350);
nand U18041 (N_18041,N_14235,N_14953);
and U18042 (N_18042,N_12630,N_11250);
xor U18043 (N_18043,N_13760,N_14121);
nand U18044 (N_18044,N_13250,N_12200);
nand U18045 (N_18045,N_10195,N_10192);
nand U18046 (N_18046,N_10769,N_11802);
and U18047 (N_18047,N_12446,N_12614);
nand U18048 (N_18048,N_11176,N_14697);
nor U18049 (N_18049,N_12721,N_11645);
xor U18050 (N_18050,N_13007,N_11100);
or U18051 (N_18051,N_13622,N_13347);
or U18052 (N_18052,N_13300,N_10842);
or U18053 (N_18053,N_12462,N_11491);
and U18054 (N_18054,N_13117,N_10591);
and U18055 (N_18055,N_10916,N_13602);
xor U18056 (N_18056,N_11510,N_13203);
or U18057 (N_18057,N_11250,N_14489);
xnor U18058 (N_18058,N_10983,N_14181);
and U18059 (N_18059,N_13544,N_10410);
and U18060 (N_18060,N_11593,N_13814);
and U18061 (N_18061,N_12757,N_10450);
and U18062 (N_18062,N_10938,N_12973);
nor U18063 (N_18063,N_10942,N_14463);
nand U18064 (N_18064,N_11529,N_14896);
or U18065 (N_18065,N_11858,N_14462);
nor U18066 (N_18066,N_11390,N_12470);
nor U18067 (N_18067,N_14245,N_12602);
xor U18068 (N_18068,N_12744,N_13024);
or U18069 (N_18069,N_12400,N_12581);
nor U18070 (N_18070,N_14912,N_10746);
nor U18071 (N_18071,N_11331,N_14902);
nand U18072 (N_18072,N_13788,N_12550);
nand U18073 (N_18073,N_11857,N_13614);
xor U18074 (N_18074,N_13567,N_12011);
nor U18075 (N_18075,N_10191,N_11401);
and U18076 (N_18076,N_11980,N_11193);
xor U18077 (N_18077,N_14003,N_10184);
nor U18078 (N_18078,N_12931,N_13004);
and U18079 (N_18079,N_10998,N_10358);
nand U18080 (N_18080,N_10903,N_10936);
or U18081 (N_18081,N_11709,N_10965);
nor U18082 (N_18082,N_14678,N_14763);
and U18083 (N_18083,N_11118,N_12094);
xor U18084 (N_18084,N_14362,N_11545);
and U18085 (N_18085,N_10743,N_13270);
xor U18086 (N_18086,N_10881,N_12511);
nor U18087 (N_18087,N_12573,N_10691);
or U18088 (N_18088,N_11763,N_13451);
and U18089 (N_18089,N_10843,N_13181);
and U18090 (N_18090,N_12790,N_12418);
nand U18091 (N_18091,N_12948,N_12994);
xor U18092 (N_18092,N_13618,N_14258);
nand U18093 (N_18093,N_12506,N_11081);
nand U18094 (N_18094,N_10921,N_10488);
xnor U18095 (N_18095,N_10586,N_11637);
nand U18096 (N_18096,N_14949,N_14638);
and U18097 (N_18097,N_13032,N_12191);
or U18098 (N_18098,N_12460,N_12256);
nor U18099 (N_18099,N_12507,N_13529);
nand U18100 (N_18100,N_11925,N_10405);
or U18101 (N_18101,N_13020,N_12155);
nand U18102 (N_18102,N_10530,N_11359);
or U18103 (N_18103,N_13964,N_10221);
xnor U18104 (N_18104,N_13778,N_11395);
and U18105 (N_18105,N_13771,N_13929);
nor U18106 (N_18106,N_13530,N_14207);
nor U18107 (N_18107,N_12772,N_11583);
and U18108 (N_18108,N_13755,N_12776);
nand U18109 (N_18109,N_14823,N_12121);
nor U18110 (N_18110,N_10577,N_13086);
or U18111 (N_18111,N_13777,N_14602);
nor U18112 (N_18112,N_13572,N_10788);
xor U18113 (N_18113,N_13632,N_13383);
nor U18114 (N_18114,N_13180,N_10563);
or U18115 (N_18115,N_11345,N_14603);
nor U18116 (N_18116,N_13625,N_11242);
xor U18117 (N_18117,N_11310,N_11813);
and U18118 (N_18118,N_13595,N_10819);
nand U18119 (N_18119,N_12152,N_14739);
nand U18120 (N_18120,N_12982,N_10690);
or U18121 (N_18121,N_12537,N_12815);
xor U18122 (N_18122,N_11976,N_10757);
and U18123 (N_18123,N_10242,N_11932);
nand U18124 (N_18124,N_13509,N_13973);
or U18125 (N_18125,N_12697,N_11593);
xnor U18126 (N_18126,N_14346,N_14249);
nand U18127 (N_18127,N_14742,N_10320);
nor U18128 (N_18128,N_12054,N_13187);
and U18129 (N_18129,N_13185,N_11917);
nor U18130 (N_18130,N_12231,N_13911);
nor U18131 (N_18131,N_12750,N_12939);
or U18132 (N_18132,N_11853,N_14027);
and U18133 (N_18133,N_12834,N_11325);
nand U18134 (N_18134,N_11512,N_11223);
xnor U18135 (N_18135,N_11895,N_14136);
nor U18136 (N_18136,N_12792,N_12111);
or U18137 (N_18137,N_14469,N_11503);
nand U18138 (N_18138,N_12552,N_11598);
and U18139 (N_18139,N_14184,N_13109);
and U18140 (N_18140,N_13446,N_14691);
and U18141 (N_18141,N_11608,N_13442);
nor U18142 (N_18142,N_14892,N_12679);
xnor U18143 (N_18143,N_13545,N_12265);
or U18144 (N_18144,N_11464,N_14774);
and U18145 (N_18145,N_11143,N_10203);
xnor U18146 (N_18146,N_11509,N_12175);
nand U18147 (N_18147,N_12269,N_11698);
nor U18148 (N_18148,N_13463,N_10954);
nand U18149 (N_18149,N_12824,N_12418);
or U18150 (N_18150,N_14763,N_13587);
nand U18151 (N_18151,N_12318,N_10369);
xor U18152 (N_18152,N_12996,N_12382);
or U18153 (N_18153,N_14608,N_14997);
xnor U18154 (N_18154,N_13831,N_10671);
or U18155 (N_18155,N_12934,N_14404);
nand U18156 (N_18156,N_11913,N_12117);
or U18157 (N_18157,N_11926,N_14830);
nand U18158 (N_18158,N_14273,N_11953);
nand U18159 (N_18159,N_13503,N_14458);
and U18160 (N_18160,N_13859,N_11765);
xnor U18161 (N_18161,N_14818,N_11115);
nand U18162 (N_18162,N_12086,N_12745);
nand U18163 (N_18163,N_14767,N_11619);
or U18164 (N_18164,N_13357,N_14112);
and U18165 (N_18165,N_11740,N_14222);
or U18166 (N_18166,N_10561,N_10700);
or U18167 (N_18167,N_13673,N_13406);
xor U18168 (N_18168,N_14132,N_10063);
or U18169 (N_18169,N_14659,N_14505);
nor U18170 (N_18170,N_11850,N_12631);
or U18171 (N_18171,N_12688,N_13953);
and U18172 (N_18172,N_12261,N_11001);
nand U18173 (N_18173,N_13810,N_14309);
nor U18174 (N_18174,N_12972,N_13340);
or U18175 (N_18175,N_13096,N_11502);
nor U18176 (N_18176,N_11263,N_12667);
nor U18177 (N_18177,N_12114,N_11205);
nand U18178 (N_18178,N_11265,N_13217);
nand U18179 (N_18179,N_11439,N_12687);
and U18180 (N_18180,N_10190,N_13458);
or U18181 (N_18181,N_10208,N_12449);
xnor U18182 (N_18182,N_13742,N_13475);
and U18183 (N_18183,N_10433,N_13160);
and U18184 (N_18184,N_14729,N_11351);
nand U18185 (N_18185,N_13936,N_13273);
nand U18186 (N_18186,N_10841,N_11261);
or U18187 (N_18187,N_10422,N_10798);
nor U18188 (N_18188,N_13645,N_13891);
or U18189 (N_18189,N_11405,N_14392);
and U18190 (N_18190,N_12048,N_14760);
or U18191 (N_18191,N_14306,N_13681);
nand U18192 (N_18192,N_13673,N_13190);
nand U18193 (N_18193,N_10473,N_12657);
and U18194 (N_18194,N_10098,N_11557);
and U18195 (N_18195,N_11443,N_11469);
nor U18196 (N_18196,N_11442,N_14408);
xnor U18197 (N_18197,N_11664,N_12637);
nand U18198 (N_18198,N_11966,N_12003);
or U18199 (N_18199,N_10824,N_11457);
nand U18200 (N_18200,N_12517,N_12371);
and U18201 (N_18201,N_13031,N_12471);
or U18202 (N_18202,N_13594,N_14215);
and U18203 (N_18203,N_13876,N_12547);
nand U18204 (N_18204,N_12870,N_10324);
nor U18205 (N_18205,N_10673,N_11866);
nor U18206 (N_18206,N_14996,N_11694);
nor U18207 (N_18207,N_11690,N_10014);
xnor U18208 (N_18208,N_14079,N_14052);
and U18209 (N_18209,N_12314,N_12515);
xor U18210 (N_18210,N_13993,N_12277);
and U18211 (N_18211,N_11824,N_11643);
nand U18212 (N_18212,N_11018,N_14955);
or U18213 (N_18213,N_12434,N_11356);
xnor U18214 (N_18214,N_14126,N_12307);
or U18215 (N_18215,N_10033,N_14068);
nor U18216 (N_18216,N_13038,N_12945);
and U18217 (N_18217,N_14521,N_10177);
xor U18218 (N_18218,N_12135,N_11377);
nand U18219 (N_18219,N_14627,N_12585);
and U18220 (N_18220,N_10047,N_12176);
nor U18221 (N_18221,N_10811,N_13927);
and U18222 (N_18222,N_12556,N_13636);
and U18223 (N_18223,N_10638,N_13720);
xnor U18224 (N_18224,N_11771,N_12488);
nor U18225 (N_18225,N_14928,N_13633);
or U18226 (N_18226,N_11481,N_12389);
xor U18227 (N_18227,N_11393,N_13301);
nor U18228 (N_18228,N_13704,N_11613);
nand U18229 (N_18229,N_14777,N_10931);
xor U18230 (N_18230,N_12756,N_12124);
nor U18231 (N_18231,N_10532,N_11957);
or U18232 (N_18232,N_12026,N_10215);
nor U18233 (N_18233,N_10910,N_10195);
or U18234 (N_18234,N_10593,N_13004);
nor U18235 (N_18235,N_11597,N_12839);
or U18236 (N_18236,N_14189,N_14080);
xor U18237 (N_18237,N_12500,N_12782);
nand U18238 (N_18238,N_14519,N_13396);
nor U18239 (N_18239,N_11897,N_12278);
xnor U18240 (N_18240,N_12591,N_10361);
nor U18241 (N_18241,N_14704,N_13122);
nor U18242 (N_18242,N_13091,N_10183);
nor U18243 (N_18243,N_14450,N_11370);
and U18244 (N_18244,N_12502,N_12789);
or U18245 (N_18245,N_13304,N_13582);
nor U18246 (N_18246,N_13934,N_12147);
nand U18247 (N_18247,N_13849,N_10599);
or U18248 (N_18248,N_12683,N_10860);
or U18249 (N_18249,N_12026,N_11054);
or U18250 (N_18250,N_14053,N_12792);
xnor U18251 (N_18251,N_14150,N_14453);
and U18252 (N_18252,N_12535,N_12959);
nor U18253 (N_18253,N_11744,N_11572);
and U18254 (N_18254,N_14640,N_14040);
nor U18255 (N_18255,N_10102,N_12171);
nor U18256 (N_18256,N_10345,N_10307);
or U18257 (N_18257,N_12477,N_12947);
nor U18258 (N_18258,N_11535,N_13025);
nand U18259 (N_18259,N_14956,N_10603);
xor U18260 (N_18260,N_14430,N_14532);
or U18261 (N_18261,N_13365,N_12989);
nand U18262 (N_18262,N_11451,N_14848);
nand U18263 (N_18263,N_11920,N_12298);
nand U18264 (N_18264,N_13521,N_14437);
xnor U18265 (N_18265,N_10120,N_12916);
nand U18266 (N_18266,N_13395,N_10411);
nand U18267 (N_18267,N_13249,N_14079);
or U18268 (N_18268,N_11911,N_12587);
nor U18269 (N_18269,N_12197,N_11160);
xor U18270 (N_18270,N_13376,N_11159);
or U18271 (N_18271,N_11750,N_13984);
and U18272 (N_18272,N_14252,N_13472);
nor U18273 (N_18273,N_13868,N_11801);
xnor U18274 (N_18274,N_13041,N_11746);
nand U18275 (N_18275,N_13237,N_11752);
nand U18276 (N_18276,N_11946,N_10879);
and U18277 (N_18277,N_14307,N_14056);
or U18278 (N_18278,N_10450,N_12034);
and U18279 (N_18279,N_13290,N_14331);
or U18280 (N_18280,N_13849,N_11587);
and U18281 (N_18281,N_13101,N_10482);
and U18282 (N_18282,N_14985,N_14792);
nand U18283 (N_18283,N_11200,N_12785);
nor U18284 (N_18284,N_14792,N_14080);
and U18285 (N_18285,N_12296,N_11253);
nor U18286 (N_18286,N_10423,N_14614);
nand U18287 (N_18287,N_14107,N_14691);
or U18288 (N_18288,N_11063,N_13317);
nand U18289 (N_18289,N_10714,N_10029);
nor U18290 (N_18290,N_13014,N_11290);
xor U18291 (N_18291,N_10297,N_14707);
xnor U18292 (N_18292,N_12613,N_14065);
and U18293 (N_18293,N_12107,N_14304);
nand U18294 (N_18294,N_10054,N_10540);
xnor U18295 (N_18295,N_12396,N_10583);
nand U18296 (N_18296,N_11517,N_10011);
nor U18297 (N_18297,N_13421,N_13832);
xor U18298 (N_18298,N_10609,N_11609);
or U18299 (N_18299,N_10532,N_11065);
xnor U18300 (N_18300,N_10269,N_14248);
nor U18301 (N_18301,N_13438,N_12067);
nand U18302 (N_18302,N_11619,N_11743);
and U18303 (N_18303,N_12266,N_13681);
and U18304 (N_18304,N_14362,N_14166);
nor U18305 (N_18305,N_13494,N_12369);
nor U18306 (N_18306,N_13305,N_11073);
nand U18307 (N_18307,N_10646,N_13259);
xnor U18308 (N_18308,N_10565,N_12739);
nor U18309 (N_18309,N_12592,N_10647);
nand U18310 (N_18310,N_14759,N_10072);
nand U18311 (N_18311,N_13176,N_13538);
and U18312 (N_18312,N_11432,N_12153);
nand U18313 (N_18313,N_12282,N_12574);
xnor U18314 (N_18314,N_13583,N_12698);
and U18315 (N_18315,N_14169,N_12323);
nor U18316 (N_18316,N_14722,N_13030);
nor U18317 (N_18317,N_10123,N_14278);
xor U18318 (N_18318,N_14646,N_10687);
xor U18319 (N_18319,N_14101,N_14404);
nor U18320 (N_18320,N_13664,N_10276);
nand U18321 (N_18321,N_14501,N_14430);
xnor U18322 (N_18322,N_12352,N_13602);
and U18323 (N_18323,N_10600,N_11046);
and U18324 (N_18324,N_13679,N_10148);
nor U18325 (N_18325,N_13757,N_12087);
nand U18326 (N_18326,N_12631,N_12235);
xnor U18327 (N_18327,N_12552,N_14292);
nor U18328 (N_18328,N_10936,N_12585);
xnor U18329 (N_18329,N_12820,N_13349);
nand U18330 (N_18330,N_13931,N_12763);
or U18331 (N_18331,N_13719,N_14893);
and U18332 (N_18332,N_12602,N_12589);
nand U18333 (N_18333,N_12358,N_11569);
and U18334 (N_18334,N_14176,N_10419);
nor U18335 (N_18335,N_12442,N_14440);
or U18336 (N_18336,N_13392,N_13671);
or U18337 (N_18337,N_14658,N_12939);
and U18338 (N_18338,N_11642,N_14299);
and U18339 (N_18339,N_13587,N_11335);
nand U18340 (N_18340,N_11931,N_13216);
xor U18341 (N_18341,N_11499,N_13439);
xor U18342 (N_18342,N_14491,N_12821);
and U18343 (N_18343,N_12298,N_11776);
or U18344 (N_18344,N_10958,N_14133);
nand U18345 (N_18345,N_14100,N_11949);
nor U18346 (N_18346,N_14445,N_10186);
and U18347 (N_18347,N_13731,N_12363);
and U18348 (N_18348,N_14205,N_13776);
and U18349 (N_18349,N_11061,N_13545);
nor U18350 (N_18350,N_14151,N_10591);
xnor U18351 (N_18351,N_11906,N_13855);
or U18352 (N_18352,N_10648,N_12029);
and U18353 (N_18353,N_13689,N_14610);
or U18354 (N_18354,N_14188,N_10361);
xnor U18355 (N_18355,N_14936,N_14433);
or U18356 (N_18356,N_13350,N_10051);
nor U18357 (N_18357,N_13059,N_13849);
nor U18358 (N_18358,N_14387,N_13657);
nor U18359 (N_18359,N_12859,N_13153);
nand U18360 (N_18360,N_11470,N_11008);
and U18361 (N_18361,N_14061,N_14691);
and U18362 (N_18362,N_10152,N_14925);
xnor U18363 (N_18363,N_12963,N_12603);
and U18364 (N_18364,N_12289,N_10743);
xnor U18365 (N_18365,N_11288,N_12250);
and U18366 (N_18366,N_13361,N_10212);
and U18367 (N_18367,N_13928,N_14499);
nand U18368 (N_18368,N_14973,N_14991);
nand U18369 (N_18369,N_11260,N_14239);
or U18370 (N_18370,N_10477,N_13675);
nand U18371 (N_18371,N_10955,N_14390);
nor U18372 (N_18372,N_10533,N_11121);
nand U18373 (N_18373,N_13773,N_11867);
or U18374 (N_18374,N_12875,N_11581);
xor U18375 (N_18375,N_12519,N_14236);
nor U18376 (N_18376,N_10850,N_12958);
nand U18377 (N_18377,N_10790,N_12130);
or U18378 (N_18378,N_13554,N_10689);
and U18379 (N_18379,N_11961,N_14907);
and U18380 (N_18380,N_13920,N_11798);
and U18381 (N_18381,N_13121,N_12029);
and U18382 (N_18382,N_14369,N_13169);
and U18383 (N_18383,N_10447,N_10553);
nor U18384 (N_18384,N_14315,N_13226);
and U18385 (N_18385,N_13326,N_13699);
nand U18386 (N_18386,N_12565,N_10829);
xnor U18387 (N_18387,N_14897,N_12578);
and U18388 (N_18388,N_10851,N_13559);
xnor U18389 (N_18389,N_12099,N_10203);
xor U18390 (N_18390,N_14568,N_12773);
xnor U18391 (N_18391,N_11513,N_14305);
nand U18392 (N_18392,N_12016,N_13691);
nand U18393 (N_18393,N_12315,N_14768);
nor U18394 (N_18394,N_12288,N_10032);
and U18395 (N_18395,N_10016,N_12048);
or U18396 (N_18396,N_13250,N_14365);
xor U18397 (N_18397,N_11980,N_12764);
or U18398 (N_18398,N_13722,N_11672);
and U18399 (N_18399,N_13051,N_14792);
nand U18400 (N_18400,N_10589,N_11849);
nand U18401 (N_18401,N_13411,N_10370);
xor U18402 (N_18402,N_12637,N_14687);
and U18403 (N_18403,N_10010,N_10921);
or U18404 (N_18404,N_12587,N_10936);
and U18405 (N_18405,N_14661,N_13044);
nand U18406 (N_18406,N_14156,N_12528);
or U18407 (N_18407,N_14762,N_14897);
and U18408 (N_18408,N_11057,N_11261);
xnor U18409 (N_18409,N_10937,N_14086);
nor U18410 (N_18410,N_10085,N_13544);
or U18411 (N_18411,N_13252,N_11516);
and U18412 (N_18412,N_13681,N_10122);
nor U18413 (N_18413,N_13765,N_11630);
or U18414 (N_18414,N_12490,N_12273);
nor U18415 (N_18415,N_11212,N_10327);
xnor U18416 (N_18416,N_12567,N_10267);
nor U18417 (N_18417,N_12641,N_13457);
nand U18418 (N_18418,N_11134,N_14845);
nand U18419 (N_18419,N_14649,N_12401);
xnor U18420 (N_18420,N_13221,N_14444);
nand U18421 (N_18421,N_11889,N_12506);
nor U18422 (N_18422,N_10871,N_10166);
nor U18423 (N_18423,N_11622,N_12237);
nand U18424 (N_18424,N_11951,N_13918);
or U18425 (N_18425,N_12314,N_12740);
nor U18426 (N_18426,N_11339,N_10978);
or U18427 (N_18427,N_12173,N_12946);
and U18428 (N_18428,N_12989,N_10327);
and U18429 (N_18429,N_12788,N_14905);
and U18430 (N_18430,N_12203,N_14671);
nor U18431 (N_18431,N_14638,N_13992);
xor U18432 (N_18432,N_10713,N_12419);
xor U18433 (N_18433,N_12276,N_10330);
nor U18434 (N_18434,N_10709,N_14021);
nor U18435 (N_18435,N_11253,N_10065);
nor U18436 (N_18436,N_10006,N_10687);
or U18437 (N_18437,N_11664,N_12574);
xor U18438 (N_18438,N_14430,N_13238);
xor U18439 (N_18439,N_11940,N_10989);
nor U18440 (N_18440,N_10774,N_14976);
and U18441 (N_18441,N_12684,N_12530);
and U18442 (N_18442,N_10078,N_12794);
or U18443 (N_18443,N_14256,N_12110);
nor U18444 (N_18444,N_12723,N_13282);
and U18445 (N_18445,N_12993,N_14223);
and U18446 (N_18446,N_11550,N_12541);
nand U18447 (N_18447,N_12851,N_10958);
nand U18448 (N_18448,N_14746,N_12756);
and U18449 (N_18449,N_11426,N_13080);
nor U18450 (N_18450,N_13034,N_10881);
nor U18451 (N_18451,N_12584,N_10294);
nand U18452 (N_18452,N_14266,N_11080);
or U18453 (N_18453,N_11378,N_11929);
nand U18454 (N_18454,N_14693,N_13850);
or U18455 (N_18455,N_13427,N_11691);
and U18456 (N_18456,N_12509,N_11217);
or U18457 (N_18457,N_13607,N_13604);
xor U18458 (N_18458,N_12667,N_11471);
nor U18459 (N_18459,N_12695,N_14674);
and U18460 (N_18460,N_12846,N_13871);
and U18461 (N_18461,N_10273,N_11551);
xnor U18462 (N_18462,N_12813,N_11685);
and U18463 (N_18463,N_12089,N_14070);
nand U18464 (N_18464,N_14781,N_10005);
and U18465 (N_18465,N_12332,N_14474);
xor U18466 (N_18466,N_12347,N_11652);
nand U18467 (N_18467,N_12941,N_14388);
nor U18468 (N_18468,N_11258,N_14639);
or U18469 (N_18469,N_13141,N_10151);
xor U18470 (N_18470,N_10480,N_12145);
xnor U18471 (N_18471,N_11202,N_10451);
nor U18472 (N_18472,N_12178,N_13386);
nand U18473 (N_18473,N_13247,N_14271);
nor U18474 (N_18474,N_11295,N_11907);
or U18475 (N_18475,N_13176,N_11039);
xnor U18476 (N_18476,N_13605,N_10770);
nand U18477 (N_18477,N_13792,N_13996);
and U18478 (N_18478,N_14384,N_12411);
nand U18479 (N_18479,N_11358,N_13221);
nor U18480 (N_18480,N_11472,N_11971);
nor U18481 (N_18481,N_13406,N_11593);
xor U18482 (N_18482,N_10384,N_11724);
or U18483 (N_18483,N_13087,N_10162);
and U18484 (N_18484,N_11404,N_11803);
xnor U18485 (N_18485,N_14635,N_10324);
xor U18486 (N_18486,N_13537,N_13069);
nor U18487 (N_18487,N_13794,N_10552);
nand U18488 (N_18488,N_11770,N_10875);
nand U18489 (N_18489,N_13899,N_12299);
nor U18490 (N_18490,N_11732,N_12354);
nor U18491 (N_18491,N_10487,N_14192);
nand U18492 (N_18492,N_10804,N_10225);
or U18493 (N_18493,N_11886,N_11867);
or U18494 (N_18494,N_14892,N_13792);
xor U18495 (N_18495,N_11595,N_12203);
xnor U18496 (N_18496,N_14829,N_13619);
nand U18497 (N_18497,N_13458,N_11583);
nand U18498 (N_18498,N_14599,N_12755);
and U18499 (N_18499,N_14763,N_14805);
and U18500 (N_18500,N_13427,N_13316);
nor U18501 (N_18501,N_10898,N_12607);
xor U18502 (N_18502,N_11259,N_13973);
xor U18503 (N_18503,N_14897,N_14579);
or U18504 (N_18504,N_11066,N_13443);
or U18505 (N_18505,N_14042,N_14704);
nor U18506 (N_18506,N_11733,N_12389);
and U18507 (N_18507,N_11013,N_13185);
nand U18508 (N_18508,N_14664,N_14489);
nand U18509 (N_18509,N_11157,N_13081);
nand U18510 (N_18510,N_10142,N_10185);
nand U18511 (N_18511,N_10740,N_10757);
and U18512 (N_18512,N_12992,N_13425);
xor U18513 (N_18513,N_13990,N_14084);
and U18514 (N_18514,N_14093,N_14098);
nor U18515 (N_18515,N_11462,N_14865);
nor U18516 (N_18516,N_11636,N_12060);
nor U18517 (N_18517,N_12346,N_10095);
xor U18518 (N_18518,N_13058,N_12661);
nor U18519 (N_18519,N_14632,N_12795);
nor U18520 (N_18520,N_12868,N_14857);
or U18521 (N_18521,N_12144,N_12832);
nand U18522 (N_18522,N_10399,N_10548);
or U18523 (N_18523,N_14990,N_10930);
xnor U18524 (N_18524,N_13065,N_13529);
nand U18525 (N_18525,N_13698,N_12012);
xor U18526 (N_18526,N_10472,N_14195);
and U18527 (N_18527,N_12425,N_13483);
or U18528 (N_18528,N_14434,N_14600);
or U18529 (N_18529,N_11488,N_13269);
nand U18530 (N_18530,N_12600,N_14652);
and U18531 (N_18531,N_12165,N_10912);
nor U18532 (N_18532,N_11573,N_11707);
or U18533 (N_18533,N_10529,N_10915);
or U18534 (N_18534,N_13999,N_11936);
or U18535 (N_18535,N_10044,N_10516);
nor U18536 (N_18536,N_13727,N_14642);
and U18537 (N_18537,N_11255,N_14367);
nand U18538 (N_18538,N_12639,N_12710);
xnor U18539 (N_18539,N_10627,N_10334);
and U18540 (N_18540,N_13134,N_12128);
nor U18541 (N_18541,N_10150,N_10496);
xor U18542 (N_18542,N_13026,N_13425);
or U18543 (N_18543,N_13543,N_11659);
xnor U18544 (N_18544,N_13503,N_12111);
nor U18545 (N_18545,N_10968,N_12148);
nand U18546 (N_18546,N_13769,N_12139);
and U18547 (N_18547,N_11849,N_14010);
nor U18548 (N_18548,N_14559,N_11210);
or U18549 (N_18549,N_12518,N_13624);
and U18550 (N_18550,N_14587,N_12067);
nand U18551 (N_18551,N_14237,N_13553);
and U18552 (N_18552,N_12946,N_11634);
or U18553 (N_18553,N_10633,N_14910);
and U18554 (N_18554,N_10446,N_10985);
or U18555 (N_18555,N_12516,N_14837);
and U18556 (N_18556,N_13070,N_14853);
and U18557 (N_18557,N_14758,N_11979);
and U18558 (N_18558,N_14279,N_11860);
or U18559 (N_18559,N_14378,N_13659);
xnor U18560 (N_18560,N_14071,N_12963);
nand U18561 (N_18561,N_10789,N_10802);
xor U18562 (N_18562,N_11379,N_14241);
xnor U18563 (N_18563,N_11932,N_13947);
nand U18564 (N_18564,N_13192,N_10486);
and U18565 (N_18565,N_11300,N_10410);
nand U18566 (N_18566,N_10007,N_10900);
xor U18567 (N_18567,N_14622,N_13133);
and U18568 (N_18568,N_13434,N_14196);
or U18569 (N_18569,N_11640,N_13449);
or U18570 (N_18570,N_11053,N_11303);
or U18571 (N_18571,N_11965,N_13810);
nand U18572 (N_18572,N_10545,N_11368);
or U18573 (N_18573,N_11399,N_14585);
nor U18574 (N_18574,N_10505,N_12713);
nand U18575 (N_18575,N_11767,N_11406);
or U18576 (N_18576,N_13272,N_13455);
and U18577 (N_18577,N_13302,N_11092);
nor U18578 (N_18578,N_14003,N_10134);
nor U18579 (N_18579,N_11344,N_11892);
xor U18580 (N_18580,N_10638,N_12474);
nor U18581 (N_18581,N_10318,N_14040);
or U18582 (N_18582,N_14476,N_11340);
nor U18583 (N_18583,N_12820,N_11900);
or U18584 (N_18584,N_12088,N_12362);
nand U18585 (N_18585,N_11456,N_10353);
nor U18586 (N_18586,N_11841,N_11448);
xnor U18587 (N_18587,N_12615,N_12416);
and U18588 (N_18588,N_12109,N_11424);
or U18589 (N_18589,N_12656,N_14175);
nor U18590 (N_18590,N_14218,N_10478);
xnor U18591 (N_18591,N_10739,N_14818);
nand U18592 (N_18592,N_12632,N_13201);
xor U18593 (N_18593,N_10979,N_12170);
or U18594 (N_18594,N_12417,N_13479);
nor U18595 (N_18595,N_13905,N_12942);
xnor U18596 (N_18596,N_13988,N_14270);
xnor U18597 (N_18597,N_11564,N_10882);
nor U18598 (N_18598,N_12826,N_14877);
nand U18599 (N_18599,N_13044,N_10051);
or U18600 (N_18600,N_12944,N_13996);
and U18601 (N_18601,N_10506,N_13108);
xnor U18602 (N_18602,N_10497,N_14448);
xnor U18603 (N_18603,N_14343,N_13385);
and U18604 (N_18604,N_10347,N_13800);
nand U18605 (N_18605,N_14375,N_10190);
and U18606 (N_18606,N_13169,N_11958);
nor U18607 (N_18607,N_14476,N_13204);
and U18608 (N_18608,N_14842,N_11151);
xor U18609 (N_18609,N_13299,N_13600);
and U18610 (N_18610,N_13557,N_14326);
or U18611 (N_18611,N_14620,N_10157);
xor U18612 (N_18612,N_14581,N_14055);
nor U18613 (N_18613,N_14998,N_10735);
nor U18614 (N_18614,N_12360,N_10081);
nor U18615 (N_18615,N_12765,N_14324);
nand U18616 (N_18616,N_13143,N_13332);
and U18617 (N_18617,N_13630,N_11160);
or U18618 (N_18618,N_10975,N_10133);
xnor U18619 (N_18619,N_11741,N_11360);
and U18620 (N_18620,N_14262,N_12387);
nand U18621 (N_18621,N_12834,N_10523);
nand U18622 (N_18622,N_10633,N_10662);
or U18623 (N_18623,N_13285,N_11929);
and U18624 (N_18624,N_14672,N_11794);
xnor U18625 (N_18625,N_14063,N_14443);
nand U18626 (N_18626,N_13799,N_10867);
nand U18627 (N_18627,N_14742,N_12355);
nand U18628 (N_18628,N_11448,N_13451);
xnor U18629 (N_18629,N_11121,N_13495);
or U18630 (N_18630,N_14037,N_14726);
xnor U18631 (N_18631,N_11174,N_11923);
or U18632 (N_18632,N_13005,N_14708);
xnor U18633 (N_18633,N_14726,N_14143);
or U18634 (N_18634,N_11413,N_11783);
xnor U18635 (N_18635,N_13181,N_11181);
and U18636 (N_18636,N_13400,N_14398);
or U18637 (N_18637,N_14325,N_14604);
xnor U18638 (N_18638,N_10328,N_13930);
nand U18639 (N_18639,N_13189,N_10224);
nand U18640 (N_18640,N_11323,N_12909);
nand U18641 (N_18641,N_11965,N_11602);
xnor U18642 (N_18642,N_12248,N_11312);
xnor U18643 (N_18643,N_10390,N_12612);
nand U18644 (N_18644,N_12171,N_10324);
or U18645 (N_18645,N_12337,N_14973);
and U18646 (N_18646,N_10696,N_14531);
nand U18647 (N_18647,N_10991,N_11338);
nor U18648 (N_18648,N_13229,N_11027);
and U18649 (N_18649,N_14215,N_13729);
nor U18650 (N_18650,N_13790,N_14802);
and U18651 (N_18651,N_12324,N_14858);
or U18652 (N_18652,N_14119,N_13210);
nand U18653 (N_18653,N_11081,N_14145);
nor U18654 (N_18654,N_11766,N_14548);
nor U18655 (N_18655,N_12229,N_12509);
or U18656 (N_18656,N_10966,N_13128);
xnor U18657 (N_18657,N_14133,N_11995);
nand U18658 (N_18658,N_12642,N_11689);
or U18659 (N_18659,N_14466,N_14346);
xor U18660 (N_18660,N_13722,N_12735);
or U18661 (N_18661,N_13903,N_13626);
or U18662 (N_18662,N_10461,N_10360);
nor U18663 (N_18663,N_13382,N_13946);
nor U18664 (N_18664,N_12247,N_12755);
xor U18665 (N_18665,N_11476,N_12528);
or U18666 (N_18666,N_14768,N_10920);
and U18667 (N_18667,N_11060,N_10708);
nor U18668 (N_18668,N_12810,N_14633);
or U18669 (N_18669,N_12987,N_11433);
and U18670 (N_18670,N_10452,N_11530);
xor U18671 (N_18671,N_12348,N_11975);
nor U18672 (N_18672,N_11816,N_14532);
and U18673 (N_18673,N_10984,N_10419);
xor U18674 (N_18674,N_12291,N_10130);
nor U18675 (N_18675,N_10347,N_10969);
or U18676 (N_18676,N_10277,N_10259);
and U18677 (N_18677,N_12900,N_11774);
nand U18678 (N_18678,N_14522,N_14559);
or U18679 (N_18679,N_12635,N_12587);
xnor U18680 (N_18680,N_13923,N_12643);
xor U18681 (N_18681,N_10045,N_13727);
nand U18682 (N_18682,N_11163,N_12635);
or U18683 (N_18683,N_12855,N_13416);
and U18684 (N_18684,N_10980,N_10378);
and U18685 (N_18685,N_12963,N_12063);
and U18686 (N_18686,N_14318,N_10844);
and U18687 (N_18687,N_10123,N_11197);
nor U18688 (N_18688,N_11802,N_14970);
and U18689 (N_18689,N_12339,N_10984);
and U18690 (N_18690,N_11762,N_11938);
xor U18691 (N_18691,N_13153,N_13114);
and U18692 (N_18692,N_12820,N_12208);
xnor U18693 (N_18693,N_12550,N_14481);
or U18694 (N_18694,N_10756,N_12051);
xnor U18695 (N_18695,N_11834,N_13747);
or U18696 (N_18696,N_12539,N_12010);
and U18697 (N_18697,N_14119,N_13907);
or U18698 (N_18698,N_14628,N_11283);
or U18699 (N_18699,N_13291,N_11622);
nand U18700 (N_18700,N_12038,N_10877);
nand U18701 (N_18701,N_12171,N_12330);
xnor U18702 (N_18702,N_13996,N_12589);
and U18703 (N_18703,N_13774,N_12537);
or U18704 (N_18704,N_14894,N_14676);
or U18705 (N_18705,N_12907,N_12318);
xnor U18706 (N_18706,N_10023,N_12775);
xor U18707 (N_18707,N_10100,N_10667);
xnor U18708 (N_18708,N_10248,N_13850);
and U18709 (N_18709,N_10987,N_13757);
xnor U18710 (N_18710,N_11324,N_10336);
nor U18711 (N_18711,N_12478,N_12262);
xor U18712 (N_18712,N_13615,N_13320);
and U18713 (N_18713,N_10486,N_13885);
and U18714 (N_18714,N_12009,N_12752);
nand U18715 (N_18715,N_14611,N_12424);
nor U18716 (N_18716,N_12734,N_11977);
and U18717 (N_18717,N_11035,N_10230);
or U18718 (N_18718,N_12395,N_13902);
or U18719 (N_18719,N_13814,N_12191);
and U18720 (N_18720,N_10639,N_13886);
nand U18721 (N_18721,N_10082,N_12839);
xnor U18722 (N_18722,N_10639,N_12930);
xor U18723 (N_18723,N_12583,N_10179);
nand U18724 (N_18724,N_10738,N_11680);
and U18725 (N_18725,N_14263,N_14799);
and U18726 (N_18726,N_12174,N_14682);
xnor U18727 (N_18727,N_14876,N_13203);
nor U18728 (N_18728,N_13180,N_12019);
nor U18729 (N_18729,N_11161,N_12495);
and U18730 (N_18730,N_14043,N_12596);
or U18731 (N_18731,N_11625,N_14810);
xor U18732 (N_18732,N_14677,N_12568);
nor U18733 (N_18733,N_14333,N_11610);
and U18734 (N_18734,N_11065,N_13557);
xnor U18735 (N_18735,N_13318,N_14298);
xnor U18736 (N_18736,N_13595,N_11460);
or U18737 (N_18737,N_14657,N_12190);
and U18738 (N_18738,N_14227,N_14050);
xor U18739 (N_18739,N_11502,N_14252);
or U18740 (N_18740,N_12102,N_14035);
nand U18741 (N_18741,N_11081,N_11788);
or U18742 (N_18742,N_12359,N_10718);
xnor U18743 (N_18743,N_14306,N_12042);
nor U18744 (N_18744,N_14067,N_12285);
nor U18745 (N_18745,N_12431,N_11995);
or U18746 (N_18746,N_10506,N_13888);
nand U18747 (N_18747,N_12190,N_11090);
nand U18748 (N_18748,N_11583,N_13532);
nor U18749 (N_18749,N_12790,N_10884);
and U18750 (N_18750,N_10570,N_13697);
or U18751 (N_18751,N_10041,N_11509);
nor U18752 (N_18752,N_12772,N_12207);
and U18753 (N_18753,N_14724,N_13018);
and U18754 (N_18754,N_10756,N_14690);
or U18755 (N_18755,N_10014,N_13718);
xnor U18756 (N_18756,N_13225,N_13601);
or U18757 (N_18757,N_13675,N_10625);
nor U18758 (N_18758,N_11605,N_13760);
and U18759 (N_18759,N_14682,N_13618);
nand U18760 (N_18760,N_12159,N_14133);
nor U18761 (N_18761,N_11132,N_13997);
nand U18762 (N_18762,N_13695,N_11099);
nand U18763 (N_18763,N_11198,N_14073);
and U18764 (N_18764,N_14877,N_10199);
or U18765 (N_18765,N_12729,N_10743);
or U18766 (N_18766,N_12949,N_12092);
xor U18767 (N_18767,N_13210,N_13044);
or U18768 (N_18768,N_12784,N_12444);
and U18769 (N_18769,N_10137,N_10978);
and U18770 (N_18770,N_11248,N_10493);
or U18771 (N_18771,N_14682,N_13762);
nor U18772 (N_18772,N_14467,N_11738);
nand U18773 (N_18773,N_12678,N_10605);
and U18774 (N_18774,N_13407,N_11695);
xor U18775 (N_18775,N_12511,N_11962);
or U18776 (N_18776,N_11747,N_14454);
or U18777 (N_18777,N_12098,N_11934);
or U18778 (N_18778,N_10424,N_14284);
and U18779 (N_18779,N_11426,N_13567);
or U18780 (N_18780,N_12142,N_11893);
nor U18781 (N_18781,N_11981,N_13878);
nor U18782 (N_18782,N_10017,N_12676);
nand U18783 (N_18783,N_12316,N_13405);
nor U18784 (N_18784,N_11206,N_10889);
nor U18785 (N_18785,N_11195,N_11673);
nand U18786 (N_18786,N_11259,N_10997);
nand U18787 (N_18787,N_10900,N_13509);
nand U18788 (N_18788,N_12519,N_13440);
xnor U18789 (N_18789,N_13793,N_12511);
xnor U18790 (N_18790,N_12143,N_14585);
nor U18791 (N_18791,N_14212,N_11563);
or U18792 (N_18792,N_14401,N_13581);
nor U18793 (N_18793,N_14506,N_10220);
or U18794 (N_18794,N_10825,N_10143);
or U18795 (N_18795,N_11168,N_13095);
and U18796 (N_18796,N_11842,N_14057);
or U18797 (N_18797,N_13256,N_12176);
xnor U18798 (N_18798,N_12168,N_14898);
xor U18799 (N_18799,N_14050,N_12961);
and U18800 (N_18800,N_13057,N_14639);
and U18801 (N_18801,N_13324,N_12276);
xor U18802 (N_18802,N_12827,N_10916);
or U18803 (N_18803,N_10567,N_13499);
nor U18804 (N_18804,N_10290,N_13224);
or U18805 (N_18805,N_12559,N_13588);
nand U18806 (N_18806,N_10906,N_14050);
nand U18807 (N_18807,N_10659,N_11709);
nand U18808 (N_18808,N_11224,N_13285);
or U18809 (N_18809,N_12823,N_14752);
nand U18810 (N_18810,N_12427,N_12678);
and U18811 (N_18811,N_10688,N_13572);
nor U18812 (N_18812,N_11973,N_14722);
nand U18813 (N_18813,N_14875,N_10565);
xor U18814 (N_18814,N_14993,N_14997);
and U18815 (N_18815,N_11073,N_10647);
or U18816 (N_18816,N_14390,N_13287);
and U18817 (N_18817,N_13088,N_14702);
or U18818 (N_18818,N_13733,N_13668);
nand U18819 (N_18819,N_14351,N_11917);
xor U18820 (N_18820,N_10104,N_13576);
xnor U18821 (N_18821,N_12188,N_10034);
nand U18822 (N_18822,N_14509,N_10089);
xnor U18823 (N_18823,N_11309,N_14494);
nand U18824 (N_18824,N_13167,N_14181);
nor U18825 (N_18825,N_11066,N_11023);
nor U18826 (N_18826,N_11613,N_12058);
and U18827 (N_18827,N_14365,N_10167);
xor U18828 (N_18828,N_13835,N_12151);
nand U18829 (N_18829,N_11897,N_10584);
or U18830 (N_18830,N_12836,N_11131);
or U18831 (N_18831,N_12082,N_10372);
nor U18832 (N_18832,N_14056,N_10748);
and U18833 (N_18833,N_11137,N_13196);
nand U18834 (N_18834,N_10183,N_11864);
nor U18835 (N_18835,N_14282,N_11070);
nand U18836 (N_18836,N_13943,N_10794);
and U18837 (N_18837,N_11902,N_11283);
nand U18838 (N_18838,N_10318,N_12565);
or U18839 (N_18839,N_11793,N_14643);
xnor U18840 (N_18840,N_10898,N_12657);
or U18841 (N_18841,N_12208,N_10835);
and U18842 (N_18842,N_11335,N_11571);
or U18843 (N_18843,N_13659,N_13585);
xnor U18844 (N_18844,N_10368,N_14910);
xnor U18845 (N_18845,N_12361,N_10102);
nor U18846 (N_18846,N_12766,N_11844);
or U18847 (N_18847,N_13847,N_13842);
xor U18848 (N_18848,N_12963,N_13766);
nor U18849 (N_18849,N_11687,N_12966);
nor U18850 (N_18850,N_10166,N_14866);
nor U18851 (N_18851,N_14366,N_13511);
xnor U18852 (N_18852,N_14989,N_12005);
nor U18853 (N_18853,N_13200,N_14292);
nand U18854 (N_18854,N_13655,N_14687);
nor U18855 (N_18855,N_12165,N_14971);
xnor U18856 (N_18856,N_13226,N_10531);
and U18857 (N_18857,N_11567,N_13338);
or U18858 (N_18858,N_12993,N_10498);
nor U18859 (N_18859,N_14577,N_10740);
xor U18860 (N_18860,N_13119,N_13712);
and U18861 (N_18861,N_13879,N_10791);
nor U18862 (N_18862,N_10584,N_10060);
and U18863 (N_18863,N_11343,N_13680);
or U18864 (N_18864,N_10434,N_13739);
or U18865 (N_18865,N_11636,N_14990);
and U18866 (N_18866,N_12175,N_10800);
xor U18867 (N_18867,N_13039,N_13246);
nor U18868 (N_18868,N_12630,N_11806);
nand U18869 (N_18869,N_11130,N_11809);
or U18870 (N_18870,N_11642,N_10439);
nor U18871 (N_18871,N_11264,N_10126);
and U18872 (N_18872,N_14476,N_11896);
or U18873 (N_18873,N_10871,N_12498);
or U18874 (N_18874,N_10342,N_14081);
or U18875 (N_18875,N_14908,N_12974);
and U18876 (N_18876,N_11824,N_13882);
nand U18877 (N_18877,N_12000,N_10661);
and U18878 (N_18878,N_11218,N_14265);
nor U18879 (N_18879,N_12259,N_11848);
or U18880 (N_18880,N_10610,N_14710);
or U18881 (N_18881,N_13690,N_11538);
xnor U18882 (N_18882,N_14447,N_10544);
or U18883 (N_18883,N_10217,N_11505);
and U18884 (N_18884,N_10992,N_11454);
nor U18885 (N_18885,N_13805,N_13649);
nand U18886 (N_18886,N_13604,N_12800);
or U18887 (N_18887,N_12883,N_11782);
nand U18888 (N_18888,N_10574,N_12718);
and U18889 (N_18889,N_11077,N_13026);
or U18890 (N_18890,N_10724,N_10595);
nor U18891 (N_18891,N_10598,N_14875);
xnor U18892 (N_18892,N_10324,N_14058);
xor U18893 (N_18893,N_14559,N_10830);
and U18894 (N_18894,N_13045,N_14974);
nor U18895 (N_18895,N_13095,N_12355);
and U18896 (N_18896,N_11700,N_12880);
nor U18897 (N_18897,N_11711,N_14932);
or U18898 (N_18898,N_14774,N_14877);
and U18899 (N_18899,N_14226,N_12868);
and U18900 (N_18900,N_11315,N_14327);
and U18901 (N_18901,N_12747,N_10763);
nand U18902 (N_18902,N_13009,N_12984);
nand U18903 (N_18903,N_13426,N_10131);
nand U18904 (N_18904,N_13592,N_11551);
nor U18905 (N_18905,N_14165,N_11955);
nand U18906 (N_18906,N_10285,N_11812);
or U18907 (N_18907,N_12061,N_11829);
nor U18908 (N_18908,N_14098,N_10287);
xnor U18909 (N_18909,N_12633,N_12622);
xor U18910 (N_18910,N_14030,N_11031);
xnor U18911 (N_18911,N_10183,N_10202);
and U18912 (N_18912,N_13625,N_14828);
nand U18913 (N_18913,N_12586,N_14238);
nand U18914 (N_18914,N_12530,N_12120);
xor U18915 (N_18915,N_10197,N_12521);
nor U18916 (N_18916,N_14933,N_10988);
xnor U18917 (N_18917,N_13588,N_11484);
xor U18918 (N_18918,N_14516,N_11507);
or U18919 (N_18919,N_11862,N_12165);
nor U18920 (N_18920,N_12000,N_13926);
or U18921 (N_18921,N_14250,N_11383);
or U18922 (N_18922,N_12084,N_12666);
nand U18923 (N_18923,N_12742,N_11011);
nor U18924 (N_18924,N_12402,N_12260);
and U18925 (N_18925,N_11731,N_14368);
nand U18926 (N_18926,N_11842,N_10919);
nor U18927 (N_18927,N_14281,N_11249);
nand U18928 (N_18928,N_11776,N_13719);
nor U18929 (N_18929,N_13492,N_13583);
xnor U18930 (N_18930,N_13964,N_14673);
xnor U18931 (N_18931,N_11493,N_11463);
nand U18932 (N_18932,N_13050,N_14272);
or U18933 (N_18933,N_12271,N_11345);
nand U18934 (N_18934,N_11613,N_14678);
nor U18935 (N_18935,N_13890,N_11839);
and U18936 (N_18936,N_10439,N_14446);
and U18937 (N_18937,N_14674,N_10565);
nor U18938 (N_18938,N_12050,N_10900);
or U18939 (N_18939,N_13861,N_11888);
xor U18940 (N_18940,N_12423,N_11242);
nor U18941 (N_18941,N_11937,N_13264);
nand U18942 (N_18942,N_12450,N_12791);
or U18943 (N_18943,N_14559,N_14927);
xor U18944 (N_18944,N_12947,N_14691);
nand U18945 (N_18945,N_11147,N_13257);
nor U18946 (N_18946,N_14111,N_12598);
nor U18947 (N_18947,N_10592,N_12089);
or U18948 (N_18948,N_11741,N_14029);
nand U18949 (N_18949,N_12620,N_10918);
nand U18950 (N_18950,N_11487,N_13067);
and U18951 (N_18951,N_11061,N_14507);
or U18952 (N_18952,N_10232,N_14617);
nor U18953 (N_18953,N_12015,N_14787);
nor U18954 (N_18954,N_11999,N_11291);
or U18955 (N_18955,N_11762,N_12042);
xnor U18956 (N_18956,N_14515,N_11376);
nand U18957 (N_18957,N_14948,N_10079);
nor U18958 (N_18958,N_11118,N_14845);
or U18959 (N_18959,N_14515,N_11796);
or U18960 (N_18960,N_14152,N_10350);
xnor U18961 (N_18961,N_10509,N_10092);
nor U18962 (N_18962,N_12285,N_12626);
and U18963 (N_18963,N_13451,N_13827);
nor U18964 (N_18964,N_14731,N_14017);
or U18965 (N_18965,N_10474,N_12360);
nor U18966 (N_18966,N_11097,N_12976);
and U18967 (N_18967,N_12693,N_11498);
nor U18968 (N_18968,N_10944,N_14950);
xor U18969 (N_18969,N_13198,N_12165);
or U18970 (N_18970,N_11129,N_12914);
and U18971 (N_18971,N_13139,N_12733);
and U18972 (N_18972,N_10918,N_10735);
or U18973 (N_18973,N_12823,N_13338);
xnor U18974 (N_18974,N_13043,N_10925);
and U18975 (N_18975,N_11588,N_11831);
xor U18976 (N_18976,N_12737,N_14017);
nand U18977 (N_18977,N_11652,N_10725);
and U18978 (N_18978,N_14045,N_10673);
xor U18979 (N_18979,N_11362,N_10274);
nor U18980 (N_18980,N_11495,N_14355);
xnor U18981 (N_18981,N_10276,N_12158);
xor U18982 (N_18982,N_11143,N_13597);
and U18983 (N_18983,N_14847,N_10744);
and U18984 (N_18984,N_10899,N_14072);
nand U18985 (N_18985,N_10026,N_14181);
nor U18986 (N_18986,N_11071,N_11747);
or U18987 (N_18987,N_12862,N_13144);
nand U18988 (N_18988,N_11686,N_10341);
nand U18989 (N_18989,N_13117,N_11188);
xnor U18990 (N_18990,N_12368,N_11749);
nor U18991 (N_18991,N_14586,N_10921);
xor U18992 (N_18992,N_12333,N_11794);
nand U18993 (N_18993,N_13267,N_11130);
nand U18994 (N_18994,N_13471,N_14035);
nand U18995 (N_18995,N_12276,N_11193);
nor U18996 (N_18996,N_11668,N_10126);
or U18997 (N_18997,N_11251,N_10137);
and U18998 (N_18998,N_12628,N_13211);
nor U18999 (N_18999,N_14278,N_10549);
and U19000 (N_19000,N_13574,N_12538);
or U19001 (N_19001,N_10049,N_10504);
nand U19002 (N_19002,N_13994,N_10606);
xnor U19003 (N_19003,N_12942,N_13541);
nor U19004 (N_19004,N_14459,N_13377);
and U19005 (N_19005,N_10227,N_10635);
xor U19006 (N_19006,N_12660,N_10618);
xnor U19007 (N_19007,N_13572,N_10686);
and U19008 (N_19008,N_13178,N_10856);
and U19009 (N_19009,N_12676,N_12592);
and U19010 (N_19010,N_11998,N_11807);
or U19011 (N_19011,N_12631,N_14483);
or U19012 (N_19012,N_10434,N_11909);
or U19013 (N_19013,N_10845,N_14944);
xnor U19014 (N_19014,N_13407,N_13520);
nand U19015 (N_19015,N_11406,N_14856);
or U19016 (N_19016,N_10116,N_13303);
xnor U19017 (N_19017,N_10569,N_10905);
nor U19018 (N_19018,N_14415,N_12677);
and U19019 (N_19019,N_13236,N_14672);
and U19020 (N_19020,N_11729,N_13705);
xnor U19021 (N_19021,N_13599,N_14016);
and U19022 (N_19022,N_11717,N_11786);
nand U19023 (N_19023,N_13902,N_12322);
nand U19024 (N_19024,N_11665,N_14981);
nand U19025 (N_19025,N_12061,N_12350);
xnor U19026 (N_19026,N_11080,N_13566);
nand U19027 (N_19027,N_11268,N_14702);
and U19028 (N_19028,N_12696,N_10197);
or U19029 (N_19029,N_14826,N_10102);
nand U19030 (N_19030,N_11302,N_10897);
or U19031 (N_19031,N_12836,N_14221);
nand U19032 (N_19032,N_12028,N_12083);
nor U19033 (N_19033,N_13450,N_11766);
or U19034 (N_19034,N_11081,N_10024);
and U19035 (N_19035,N_10963,N_14738);
nor U19036 (N_19036,N_10190,N_13161);
nand U19037 (N_19037,N_12102,N_13664);
xor U19038 (N_19038,N_12520,N_14907);
xnor U19039 (N_19039,N_14848,N_12585);
nand U19040 (N_19040,N_12323,N_14086);
and U19041 (N_19041,N_13607,N_12623);
nand U19042 (N_19042,N_10119,N_11257);
nor U19043 (N_19043,N_12722,N_12998);
nand U19044 (N_19044,N_11283,N_12927);
xor U19045 (N_19045,N_11187,N_13167);
nor U19046 (N_19046,N_10424,N_14916);
xnor U19047 (N_19047,N_13174,N_11481);
xnor U19048 (N_19048,N_11927,N_10783);
nor U19049 (N_19049,N_13518,N_12744);
or U19050 (N_19050,N_14407,N_10340);
and U19051 (N_19051,N_14720,N_13893);
nor U19052 (N_19052,N_10444,N_10311);
xnor U19053 (N_19053,N_13464,N_14757);
and U19054 (N_19054,N_11649,N_11385);
or U19055 (N_19055,N_12349,N_13686);
xor U19056 (N_19056,N_10245,N_11170);
or U19057 (N_19057,N_10607,N_14604);
xor U19058 (N_19058,N_14670,N_14560);
nor U19059 (N_19059,N_10026,N_14644);
or U19060 (N_19060,N_12625,N_13645);
or U19061 (N_19061,N_14922,N_13881);
or U19062 (N_19062,N_13264,N_13102);
or U19063 (N_19063,N_14677,N_14234);
and U19064 (N_19064,N_10356,N_13139);
nor U19065 (N_19065,N_13899,N_13560);
or U19066 (N_19066,N_11937,N_11944);
or U19067 (N_19067,N_12902,N_10150);
nor U19068 (N_19068,N_14741,N_13622);
nand U19069 (N_19069,N_13902,N_10091);
nor U19070 (N_19070,N_10399,N_11916);
nand U19071 (N_19071,N_12453,N_10791);
and U19072 (N_19072,N_12500,N_14871);
xnor U19073 (N_19073,N_14337,N_13110);
nor U19074 (N_19074,N_12667,N_14680);
nand U19075 (N_19075,N_10145,N_10918);
nor U19076 (N_19076,N_10606,N_12669);
nand U19077 (N_19077,N_14017,N_11599);
nor U19078 (N_19078,N_10158,N_10925);
nor U19079 (N_19079,N_11092,N_12977);
and U19080 (N_19080,N_14411,N_13037);
xnor U19081 (N_19081,N_13963,N_10822);
or U19082 (N_19082,N_13764,N_11066);
nand U19083 (N_19083,N_14270,N_14694);
nor U19084 (N_19084,N_13863,N_13440);
or U19085 (N_19085,N_12989,N_12952);
and U19086 (N_19086,N_14746,N_11595);
nand U19087 (N_19087,N_13593,N_14989);
or U19088 (N_19088,N_13038,N_11495);
and U19089 (N_19089,N_14489,N_12488);
nand U19090 (N_19090,N_14559,N_10639);
xnor U19091 (N_19091,N_13628,N_13760);
and U19092 (N_19092,N_14012,N_12229);
xor U19093 (N_19093,N_13556,N_10276);
xor U19094 (N_19094,N_12250,N_13949);
nand U19095 (N_19095,N_10640,N_14853);
nor U19096 (N_19096,N_12007,N_12830);
xnor U19097 (N_19097,N_14236,N_14335);
and U19098 (N_19098,N_11925,N_11631);
xnor U19099 (N_19099,N_14259,N_11071);
nor U19100 (N_19100,N_11949,N_12818);
nand U19101 (N_19101,N_10457,N_14121);
nand U19102 (N_19102,N_14544,N_13974);
xor U19103 (N_19103,N_14808,N_11394);
xnor U19104 (N_19104,N_10755,N_12437);
or U19105 (N_19105,N_13529,N_11180);
nor U19106 (N_19106,N_13016,N_14157);
nand U19107 (N_19107,N_11793,N_12283);
and U19108 (N_19108,N_13219,N_14657);
nand U19109 (N_19109,N_14282,N_14416);
xnor U19110 (N_19110,N_13414,N_10605);
and U19111 (N_19111,N_12133,N_13357);
nor U19112 (N_19112,N_14727,N_11754);
nand U19113 (N_19113,N_14266,N_13373);
or U19114 (N_19114,N_10904,N_11747);
and U19115 (N_19115,N_11456,N_12826);
xnor U19116 (N_19116,N_10993,N_11060);
or U19117 (N_19117,N_13257,N_11029);
and U19118 (N_19118,N_12773,N_13445);
nand U19119 (N_19119,N_11291,N_12031);
nand U19120 (N_19120,N_14074,N_13124);
or U19121 (N_19121,N_14433,N_13700);
nor U19122 (N_19122,N_11530,N_10304);
xor U19123 (N_19123,N_12455,N_14492);
nor U19124 (N_19124,N_11534,N_14994);
nor U19125 (N_19125,N_14200,N_11616);
or U19126 (N_19126,N_11553,N_14138);
nand U19127 (N_19127,N_13319,N_11800);
nand U19128 (N_19128,N_13729,N_14856);
or U19129 (N_19129,N_11220,N_12822);
xnor U19130 (N_19130,N_10498,N_12180);
or U19131 (N_19131,N_12914,N_14695);
or U19132 (N_19132,N_12001,N_10267);
nor U19133 (N_19133,N_12007,N_10502);
or U19134 (N_19134,N_10666,N_13384);
nor U19135 (N_19135,N_12985,N_13143);
nand U19136 (N_19136,N_10328,N_10979);
nor U19137 (N_19137,N_13655,N_13365);
xor U19138 (N_19138,N_13990,N_12061);
nand U19139 (N_19139,N_13530,N_13414);
or U19140 (N_19140,N_10732,N_14272);
nand U19141 (N_19141,N_14529,N_14413);
or U19142 (N_19142,N_10194,N_14751);
nand U19143 (N_19143,N_11204,N_14346);
or U19144 (N_19144,N_11526,N_14642);
nor U19145 (N_19145,N_10970,N_11345);
nand U19146 (N_19146,N_13228,N_10349);
xnor U19147 (N_19147,N_12271,N_10386);
xnor U19148 (N_19148,N_12088,N_11690);
or U19149 (N_19149,N_13989,N_14508);
nor U19150 (N_19150,N_11330,N_11295);
nand U19151 (N_19151,N_11258,N_14043);
or U19152 (N_19152,N_10524,N_12579);
and U19153 (N_19153,N_11222,N_13743);
and U19154 (N_19154,N_12186,N_11488);
xor U19155 (N_19155,N_13883,N_12946);
or U19156 (N_19156,N_13077,N_12618);
or U19157 (N_19157,N_11503,N_13362);
nand U19158 (N_19158,N_13757,N_13849);
and U19159 (N_19159,N_14271,N_10539);
nor U19160 (N_19160,N_13872,N_13092);
and U19161 (N_19161,N_11062,N_10738);
nand U19162 (N_19162,N_11228,N_12619);
nand U19163 (N_19163,N_10745,N_12170);
nor U19164 (N_19164,N_13532,N_10651);
or U19165 (N_19165,N_14467,N_12518);
or U19166 (N_19166,N_10173,N_12729);
nor U19167 (N_19167,N_10471,N_10915);
and U19168 (N_19168,N_14188,N_14172);
nor U19169 (N_19169,N_13975,N_11995);
or U19170 (N_19170,N_13509,N_12292);
nor U19171 (N_19171,N_11573,N_12702);
nor U19172 (N_19172,N_14184,N_10075);
nand U19173 (N_19173,N_14330,N_14558);
nor U19174 (N_19174,N_11595,N_12318);
and U19175 (N_19175,N_13427,N_10882);
nand U19176 (N_19176,N_10533,N_10050);
or U19177 (N_19177,N_10881,N_10331);
or U19178 (N_19178,N_11760,N_14817);
nor U19179 (N_19179,N_12824,N_13632);
xor U19180 (N_19180,N_13795,N_11954);
nand U19181 (N_19181,N_11453,N_11008);
xor U19182 (N_19182,N_13412,N_10961);
and U19183 (N_19183,N_11419,N_11119);
nor U19184 (N_19184,N_10447,N_13333);
nor U19185 (N_19185,N_13208,N_11545);
nand U19186 (N_19186,N_13618,N_14949);
xnor U19187 (N_19187,N_11565,N_14664);
nor U19188 (N_19188,N_10726,N_12070);
xnor U19189 (N_19189,N_12273,N_10192);
nor U19190 (N_19190,N_10011,N_14873);
or U19191 (N_19191,N_13079,N_13496);
and U19192 (N_19192,N_14036,N_11293);
nor U19193 (N_19193,N_11170,N_13042);
nand U19194 (N_19194,N_13881,N_12153);
xnor U19195 (N_19195,N_11745,N_10985);
and U19196 (N_19196,N_13349,N_11251);
and U19197 (N_19197,N_10284,N_13172);
and U19198 (N_19198,N_10054,N_13494);
and U19199 (N_19199,N_14591,N_11090);
and U19200 (N_19200,N_10023,N_13437);
xnor U19201 (N_19201,N_11411,N_14856);
xnor U19202 (N_19202,N_13719,N_10197);
nor U19203 (N_19203,N_14620,N_14857);
nor U19204 (N_19204,N_11146,N_14473);
and U19205 (N_19205,N_10533,N_11365);
xor U19206 (N_19206,N_12466,N_11721);
and U19207 (N_19207,N_11928,N_11271);
xor U19208 (N_19208,N_12718,N_11420);
or U19209 (N_19209,N_10621,N_14694);
xor U19210 (N_19210,N_14183,N_12650);
nor U19211 (N_19211,N_10861,N_13987);
xor U19212 (N_19212,N_11292,N_13841);
and U19213 (N_19213,N_14342,N_11560);
nand U19214 (N_19214,N_11599,N_13136);
nor U19215 (N_19215,N_10229,N_12068);
xnor U19216 (N_19216,N_14995,N_14121);
nand U19217 (N_19217,N_13549,N_14372);
nand U19218 (N_19218,N_13433,N_10422);
nand U19219 (N_19219,N_11018,N_11626);
or U19220 (N_19220,N_10300,N_12342);
xnor U19221 (N_19221,N_12879,N_14790);
nor U19222 (N_19222,N_13435,N_11487);
nand U19223 (N_19223,N_13154,N_13594);
or U19224 (N_19224,N_12261,N_10851);
nor U19225 (N_19225,N_14055,N_14871);
xor U19226 (N_19226,N_12070,N_11885);
nor U19227 (N_19227,N_13356,N_13291);
and U19228 (N_19228,N_10626,N_12928);
nor U19229 (N_19229,N_10586,N_14047);
nand U19230 (N_19230,N_13984,N_12088);
xor U19231 (N_19231,N_10129,N_11570);
or U19232 (N_19232,N_14185,N_11028);
nor U19233 (N_19233,N_12821,N_13051);
xnor U19234 (N_19234,N_13169,N_14462);
nor U19235 (N_19235,N_10463,N_14947);
xor U19236 (N_19236,N_12900,N_13918);
nand U19237 (N_19237,N_10162,N_10674);
nand U19238 (N_19238,N_13716,N_13309);
xnor U19239 (N_19239,N_13175,N_14112);
and U19240 (N_19240,N_12856,N_11799);
nor U19241 (N_19241,N_11729,N_12962);
nand U19242 (N_19242,N_10398,N_14603);
nand U19243 (N_19243,N_12569,N_13028);
nor U19244 (N_19244,N_14002,N_13247);
and U19245 (N_19245,N_11053,N_10118);
and U19246 (N_19246,N_12904,N_10673);
or U19247 (N_19247,N_13365,N_13560);
and U19248 (N_19248,N_11624,N_10296);
or U19249 (N_19249,N_12607,N_13829);
and U19250 (N_19250,N_14703,N_13084);
nor U19251 (N_19251,N_14248,N_14351);
and U19252 (N_19252,N_12733,N_14821);
nor U19253 (N_19253,N_13951,N_11233);
nor U19254 (N_19254,N_10374,N_11015);
and U19255 (N_19255,N_13629,N_13741);
nor U19256 (N_19256,N_13873,N_12369);
xnor U19257 (N_19257,N_13177,N_12729);
nand U19258 (N_19258,N_12522,N_11270);
and U19259 (N_19259,N_13725,N_13784);
or U19260 (N_19260,N_14771,N_14698);
nor U19261 (N_19261,N_11360,N_12187);
and U19262 (N_19262,N_13230,N_14247);
nand U19263 (N_19263,N_14857,N_10849);
nor U19264 (N_19264,N_13964,N_13827);
xnor U19265 (N_19265,N_14936,N_13588);
nor U19266 (N_19266,N_12146,N_11141);
nor U19267 (N_19267,N_14834,N_13339);
nor U19268 (N_19268,N_14247,N_11192);
or U19269 (N_19269,N_11755,N_10433);
xor U19270 (N_19270,N_11105,N_13270);
nor U19271 (N_19271,N_10101,N_10640);
and U19272 (N_19272,N_11940,N_14114);
and U19273 (N_19273,N_12083,N_12208);
xor U19274 (N_19274,N_14039,N_10438);
or U19275 (N_19275,N_13466,N_11077);
xnor U19276 (N_19276,N_12995,N_13870);
and U19277 (N_19277,N_11527,N_12353);
nand U19278 (N_19278,N_11959,N_11401);
nand U19279 (N_19279,N_12821,N_12609);
nor U19280 (N_19280,N_11209,N_11094);
and U19281 (N_19281,N_14396,N_11540);
nand U19282 (N_19282,N_10406,N_10914);
and U19283 (N_19283,N_13290,N_13431);
nand U19284 (N_19284,N_11032,N_12112);
or U19285 (N_19285,N_12162,N_12208);
nor U19286 (N_19286,N_13121,N_13022);
nor U19287 (N_19287,N_13359,N_12008);
nand U19288 (N_19288,N_13532,N_12925);
nand U19289 (N_19289,N_13093,N_11346);
or U19290 (N_19290,N_13242,N_13225);
or U19291 (N_19291,N_14815,N_14820);
nand U19292 (N_19292,N_10851,N_12204);
nor U19293 (N_19293,N_14496,N_13454);
nor U19294 (N_19294,N_12790,N_14316);
nand U19295 (N_19295,N_11101,N_12693);
and U19296 (N_19296,N_12151,N_10956);
or U19297 (N_19297,N_12055,N_12133);
nand U19298 (N_19298,N_12691,N_11249);
or U19299 (N_19299,N_11266,N_14747);
xnor U19300 (N_19300,N_10789,N_11377);
and U19301 (N_19301,N_13296,N_12701);
nand U19302 (N_19302,N_13262,N_10370);
nand U19303 (N_19303,N_14968,N_11500);
and U19304 (N_19304,N_12547,N_13614);
nor U19305 (N_19305,N_13834,N_12332);
nor U19306 (N_19306,N_12834,N_13291);
xor U19307 (N_19307,N_14097,N_12813);
or U19308 (N_19308,N_11017,N_11542);
or U19309 (N_19309,N_10673,N_10593);
nor U19310 (N_19310,N_14037,N_13415);
and U19311 (N_19311,N_12190,N_13735);
nor U19312 (N_19312,N_14506,N_12108);
or U19313 (N_19313,N_13245,N_14861);
and U19314 (N_19314,N_10034,N_12842);
nor U19315 (N_19315,N_12861,N_14399);
or U19316 (N_19316,N_12193,N_14073);
or U19317 (N_19317,N_14689,N_14230);
nor U19318 (N_19318,N_11508,N_11579);
nand U19319 (N_19319,N_12988,N_13135);
nor U19320 (N_19320,N_10706,N_10940);
nand U19321 (N_19321,N_14604,N_10729);
or U19322 (N_19322,N_12615,N_10580);
nand U19323 (N_19323,N_10297,N_10001);
and U19324 (N_19324,N_13917,N_10500);
xnor U19325 (N_19325,N_14621,N_11096);
and U19326 (N_19326,N_12122,N_12701);
xnor U19327 (N_19327,N_11217,N_14584);
nor U19328 (N_19328,N_12175,N_13997);
nand U19329 (N_19329,N_11131,N_14761);
xnor U19330 (N_19330,N_10081,N_14487);
and U19331 (N_19331,N_10236,N_13908);
nand U19332 (N_19332,N_10724,N_14766);
xor U19333 (N_19333,N_10625,N_12870);
and U19334 (N_19334,N_14713,N_10376);
nand U19335 (N_19335,N_10268,N_12485);
or U19336 (N_19336,N_13007,N_12623);
xnor U19337 (N_19337,N_14753,N_12324);
xor U19338 (N_19338,N_12529,N_14782);
nor U19339 (N_19339,N_11034,N_10651);
nand U19340 (N_19340,N_14434,N_13033);
nand U19341 (N_19341,N_13686,N_12966);
nand U19342 (N_19342,N_11934,N_13430);
and U19343 (N_19343,N_13261,N_13316);
nand U19344 (N_19344,N_10410,N_11751);
xnor U19345 (N_19345,N_13920,N_14251);
and U19346 (N_19346,N_10524,N_12519);
and U19347 (N_19347,N_13306,N_14743);
or U19348 (N_19348,N_10967,N_12501);
nor U19349 (N_19349,N_14480,N_11331);
or U19350 (N_19350,N_13454,N_10193);
or U19351 (N_19351,N_12273,N_11007);
xnor U19352 (N_19352,N_13114,N_13130);
xnor U19353 (N_19353,N_11403,N_11005);
or U19354 (N_19354,N_12962,N_12992);
or U19355 (N_19355,N_11120,N_12381);
xor U19356 (N_19356,N_10991,N_14492);
xor U19357 (N_19357,N_12319,N_10438);
and U19358 (N_19358,N_11283,N_14733);
xor U19359 (N_19359,N_12136,N_11084);
and U19360 (N_19360,N_11876,N_14922);
and U19361 (N_19361,N_12597,N_12514);
nand U19362 (N_19362,N_13482,N_13407);
xnor U19363 (N_19363,N_12853,N_11548);
nand U19364 (N_19364,N_13466,N_13179);
nor U19365 (N_19365,N_12450,N_12067);
xnor U19366 (N_19366,N_13699,N_13148);
or U19367 (N_19367,N_12485,N_13265);
xnor U19368 (N_19368,N_10900,N_12827);
or U19369 (N_19369,N_11794,N_10851);
nor U19370 (N_19370,N_10606,N_11832);
xnor U19371 (N_19371,N_13462,N_10170);
xor U19372 (N_19372,N_11506,N_10143);
or U19373 (N_19373,N_10602,N_10099);
xnor U19374 (N_19374,N_13757,N_13488);
nand U19375 (N_19375,N_13152,N_11748);
or U19376 (N_19376,N_11317,N_10814);
xor U19377 (N_19377,N_12728,N_13248);
xnor U19378 (N_19378,N_11892,N_10437);
nor U19379 (N_19379,N_13037,N_14719);
or U19380 (N_19380,N_13266,N_10501);
nor U19381 (N_19381,N_14291,N_11774);
nor U19382 (N_19382,N_13219,N_11320);
xor U19383 (N_19383,N_12408,N_11399);
or U19384 (N_19384,N_13781,N_12476);
xnor U19385 (N_19385,N_12583,N_11736);
and U19386 (N_19386,N_13035,N_14825);
and U19387 (N_19387,N_11672,N_13397);
nand U19388 (N_19388,N_11504,N_11722);
nand U19389 (N_19389,N_13147,N_14325);
xor U19390 (N_19390,N_12422,N_11937);
xnor U19391 (N_19391,N_10391,N_11973);
xor U19392 (N_19392,N_11199,N_13689);
xnor U19393 (N_19393,N_11826,N_13638);
xnor U19394 (N_19394,N_13816,N_11091);
nor U19395 (N_19395,N_14802,N_11027);
or U19396 (N_19396,N_10038,N_10578);
xnor U19397 (N_19397,N_14870,N_12151);
and U19398 (N_19398,N_11595,N_11349);
nor U19399 (N_19399,N_14865,N_10960);
or U19400 (N_19400,N_14293,N_10110);
xor U19401 (N_19401,N_13259,N_12856);
or U19402 (N_19402,N_10748,N_13250);
xor U19403 (N_19403,N_14563,N_10976);
or U19404 (N_19404,N_14117,N_11804);
and U19405 (N_19405,N_10353,N_10668);
or U19406 (N_19406,N_11337,N_14480);
nor U19407 (N_19407,N_13401,N_13317);
nor U19408 (N_19408,N_10042,N_11905);
nand U19409 (N_19409,N_14678,N_11045);
xnor U19410 (N_19410,N_11068,N_13848);
xor U19411 (N_19411,N_11131,N_10357);
and U19412 (N_19412,N_13812,N_12712);
nor U19413 (N_19413,N_14290,N_12835);
nand U19414 (N_19414,N_11077,N_10904);
and U19415 (N_19415,N_13753,N_13195);
nor U19416 (N_19416,N_10340,N_12012);
nand U19417 (N_19417,N_11905,N_13088);
xor U19418 (N_19418,N_11153,N_11718);
or U19419 (N_19419,N_13766,N_14291);
and U19420 (N_19420,N_12234,N_12815);
and U19421 (N_19421,N_12639,N_11390);
nor U19422 (N_19422,N_12797,N_10673);
xor U19423 (N_19423,N_11875,N_10866);
or U19424 (N_19424,N_13774,N_12099);
or U19425 (N_19425,N_10737,N_14034);
or U19426 (N_19426,N_13135,N_10589);
or U19427 (N_19427,N_14156,N_13209);
nor U19428 (N_19428,N_10053,N_13358);
xnor U19429 (N_19429,N_13763,N_13453);
xnor U19430 (N_19430,N_10268,N_12407);
nand U19431 (N_19431,N_13345,N_13019);
and U19432 (N_19432,N_13256,N_14662);
or U19433 (N_19433,N_12650,N_11990);
and U19434 (N_19434,N_14268,N_14158);
nor U19435 (N_19435,N_13647,N_11399);
or U19436 (N_19436,N_12798,N_14515);
nand U19437 (N_19437,N_12028,N_11662);
and U19438 (N_19438,N_12984,N_14283);
xnor U19439 (N_19439,N_10406,N_12050);
and U19440 (N_19440,N_14292,N_11322);
nor U19441 (N_19441,N_13393,N_13414);
or U19442 (N_19442,N_11787,N_13164);
or U19443 (N_19443,N_14769,N_13045);
nor U19444 (N_19444,N_14553,N_11834);
and U19445 (N_19445,N_10118,N_12465);
nand U19446 (N_19446,N_14909,N_14493);
xor U19447 (N_19447,N_13209,N_11378);
nor U19448 (N_19448,N_13999,N_12781);
nor U19449 (N_19449,N_12094,N_13465);
or U19450 (N_19450,N_12226,N_13127);
or U19451 (N_19451,N_13053,N_13257);
or U19452 (N_19452,N_14728,N_13886);
nor U19453 (N_19453,N_14119,N_14526);
nand U19454 (N_19454,N_13807,N_10875);
or U19455 (N_19455,N_12427,N_14815);
and U19456 (N_19456,N_12138,N_10459);
xor U19457 (N_19457,N_11058,N_14407);
nand U19458 (N_19458,N_14420,N_12565);
nand U19459 (N_19459,N_14218,N_12277);
nand U19460 (N_19460,N_12440,N_11740);
xnor U19461 (N_19461,N_12405,N_10309);
or U19462 (N_19462,N_13974,N_12287);
and U19463 (N_19463,N_13071,N_10397);
nor U19464 (N_19464,N_10870,N_13921);
and U19465 (N_19465,N_12483,N_13408);
nor U19466 (N_19466,N_13852,N_14420);
nor U19467 (N_19467,N_10256,N_12429);
xnor U19468 (N_19468,N_12209,N_14243);
nand U19469 (N_19469,N_12022,N_12598);
nand U19470 (N_19470,N_11746,N_13746);
nor U19471 (N_19471,N_11211,N_14321);
nand U19472 (N_19472,N_10313,N_10628);
or U19473 (N_19473,N_11420,N_12844);
and U19474 (N_19474,N_10099,N_14755);
and U19475 (N_19475,N_14736,N_12629);
xor U19476 (N_19476,N_13352,N_11951);
or U19477 (N_19477,N_11521,N_13466);
and U19478 (N_19478,N_10534,N_10635);
or U19479 (N_19479,N_12719,N_14493);
xor U19480 (N_19480,N_13024,N_14134);
nand U19481 (N_19481,N_12208,N_10276);
or U19482 (N_19482,N_13225,N_12625);
xnor U19483 (N_19483,N_13671,N_12013);
nand U19484 (N_19484,N_14879,N_12641);
and U19485 (N_19485,N_13163,N_11512);
nand U19486 (N_19486,N_10439,N_11104);
and U19487 (N_19487,N_13421,N_14928);
xnor U19488 (N_19488,N_11556,N_13990);
nor U19489 (N_19489,N_12559,N_10780);
xnor U19490 (N_19490,N_14484,N_10557);
and U19491 (N_19491,N_11392,N_11779);
nand U19492 (N_19492,N_10503,N_11150);
nand U19493 (N_19493,N_12453,N_11860);
nor U19494 (N_19494,N_11715,N_14472);
nor U19495 (N_19495,N_14184,N_11165);
nand U19496 (N_19496,N_14677,N_11194);
or U19497 (N_19497,N_13414,N_13515);
nand U19498 (N_19498,N_11469,N_12779);
or U19499 (N_19499,N_10568,N_10226);
xor U19500 (N_19500,N_12912,N_11952);
nand U19501 (N_19501,N_11195,N_11088);
nand U19502 (N_19502,N_11756,N_10678);
nand U19503 (N_19503,N_10579,N_11719);
and U19504 (N_19504,N_10303,N_13394);
or U19505 (N_19505,N_14197,N_13783);
or U19506 (N_19506,N_13663,N_10798);
or U19507 (N_19507,N_13066,N_11295);
nand U19508 (N_19508,N_10300,N_12973);
nor U19509 (N_19509,N_14918,N_12274);
nor U19510 (N_19510,N_14479,N_10019);
xnor U19511 (N_19511,N_11129,N_14639);
xnor U19512 (N_19512,N_10529,N_13216);
xnor U19513 (N_19513,N_12747,N_12733);
xor U19514 (N_19514,N_10779,N_13474);
or U19515 (N_19515,N_11738,N_12748);
xnor U19516 (N_19516,N_11691,N_12132);
nor U19517 (N_19517,N_10730,N_12491);
and U19518 (N_19518,N_12574,N_14170);
and U19519 (N_19519,N_12643,N_12850);
nand U19520 (N_19520,N_13787,N_10130);
nand U19521 (N_19521,N_12115,N_12192);
and U19522 (N_19522,N_10183,N_10251);
nand U19523 (N_19523,N_11144,N_11134);
and U19524 (N_19524,N_13631,N_14061);
and U19525 (N_19525,N_10517,N_10371);
nand U19526 (N_19526,N_12057,N_12027);
nand U19527 (N_19527,N_10760,N_10091);
nor U19528 (N_19528,N_13274,N_13404);
xor U19529 (N_19529,N_11828,N_12120);
xor U19530 (N_19530,N_10117,N_10653);
and U19531 (N_19531,N_11119,N_10266);
or U19532 (N_19532,N_11990,N_10084);
or U19533 (N_19533,N_14466,N_11639);
or U19534 (N_19534,N_12000,N_10726);
and U19535 (N_19535,N_13785,N_12589);
nand U19536 (N_19536,N_12688,N_13852);
nand U19537 (N_19537,N_14228,N_13769);
and U19538 (N_19538,N_10222,N_10496);
nand U19539 (N_19539,N_10612,N_10456);
nand U19540 (N_19540,N_12184,N_10317);
nand U19541 (N_19541,N_14566,N_10038);
nor U19542 (N_19542,N_12379,N_14831);
or U19543 (N_19543,N_10196,N_10845);
nor U19544 (N_19544,N_14294,N_14244);
nor U19545 (N_19545,N_13624,N_12633);
and U19546 (N_19546,N_11519,N_12963);
nand U19547 (N_19547,N_13159,N_10122);
nand U19548 (N_19548,N_12084,N_13190);
nor U19549 (N_19549,N_10062,N_11807);
or U19550 (N_19550,N_12802,N_11142);
nand U19551 (N_19551,N_12992,N_12594);
xnor U19552 (N_19552,N_13136,N_12914);
xnor U19553 (N_19553,N_14758,N_12483);
and U19554 (N_19554,N_13801,N_14104);
nand U19555 (N_19555,N_12934,N_10930);
nor U19556 (N_19556,N_13325,N_12411);
xnor U19557 (N_19557,N_11511,N_10446);
or U19558 (N_19558,N_10645,N_10829);
nor U19559 (N_19559,N_12437,N_12005);
nand U19560 (N_19560,N_14690,N_13796);
and U19561 (N_19561,N_10298,N_10090);
nor U19562 (N_19562,N_14784,N_14596);
nor U19563 (N_19563,N_13484,N_10452);
or U19564 (N_19564,N_13698,N_10073);
xnor U19565 (N_19565,N_11440,N_14637);
and U19566 (N_19566,N_12643,N_11728);
or U19567 (N_19567,N_11672,N_14592);
nor U19568 (N_19568,N_12981,N_13853);
and U19569 (N_19569,N_11749,N_12901);
and U19570 (N_19570,N_12520,N_14698);
nor U19571 (N_19571,N_10592,N_12987);
and U19572 (N_19572,N_14754,N_10206);
nand U19573 (N_19573,N_10905,N_13325);
or U19574 (N_19574,N_11843,N_10917);
xor U19575 (N_19575,N_11652,N_13024);
nor U19576 (N_19576,N_10378,N_13587);
and U19577 (N_19577,N_10323,N_12324);
xor U19578 (N_19578,N_11402,N_10900);
nor U19579 (N_19579,N_11318,N_14926);
xnor U19580 (N_19580,N_10149,N_10496);
and U19581 (N_19581,N_13519,N_14985);
and U19582 (N_19582,N_10971,N_10593);
nand U19583 (N_19583,N_11681,N_14904);
xnor U19584 (N_19584,N_14242,N_10992);
nand U19585 (N_19585,N_10892,N_14749);
and U19586 (N_19586,N_10258,N_12571);
xnor U19587 (N_19587,N_14673,N_14361);
xor U19588 (N_19588,N_10610,N_11535);
and U19589 (N_19589,N_11214,N_14561);
nand U19590 (N_19590,N_14202,N_14122);
or U19591 (N_19591,N_11873,N_12073);
and U19592 (N_19592,N_12146,N_12093);
and U19593 (N_19593,N_10055,N_12100);
or U19594 (N_19594,N_14644,N_10368);
xor U19595 (N_19595,N_12230,N_12324);
nor U19596 (N_19596,N_13205,N_10727);
or U19597 (N_19597,N_11110,N_14475);
and U19598 (N_19598,N_10919,N_13160);
or U19599 (N_19599,N_14419,N_11580);
and U19600 (N_19600,N_10366,N_14450);
nor U19601 (N_19601,N_13063,N_12660);
and U19602 (N_19602,N_11374,N_12911);
and U19603 (N_19603,N_14399,N_14667);
nor U19604 (N_19604,N_11945,N_13432);
and U19605 (N_19605,N_13494,N_12385);
or U19606 (N_19606,N_11002,N_14758);
and U19607 (N_19607,N_10947,N_11422);
nor U19608 (N_19608,N_14328,N_14338);
and U19609 (N_19609,N_11524,N_10318);
and U19610 (N_19610,N_14790,N_11867);
xnor U19611 (N_19611,N_10496,N_11460);
nor U19612 (N_19612,N_12155,N_14058);
and U19613 (N_19613,N_11968,N_11922);
nor U19614 (N_19614,N_13802,N_12281);
xor U19615 (N_19615,N_11719,N_10698);
and U19616 (N_19616,N_12576,N_12762);
and U19617 (N_19617,N_11130,N_10806);
or U19618 (N_19618,N_13055,N_14097);
nor U19619 (N_19619,N_14096,N_11706);
xnor U19620 (N_19620,N_12656,N_14663);
and U19621 (N_19621,N_13676,N_13616);
and U19622 (N_19622,N_14230,N_10124);
or U19623 (N_19623,N_13195,N_13053);
nor U19624 (N_19624,N_13540,N_13037);
nand U19625 (N_19625,N_14315,N_14747);
nand U19626 (N_19626,N_11532,N_13578);
or U19627 (N_19627,N_10437,N_12080);
nand U19628 (N_19628,N_11010,N_13338);
nand U19629 (N_19629,N_13740,N_12745);
nand U19630 (N_19630,N_10230,N_13993);
nor U19631 (N_19631,N_13519,N_13687);
nor U19632 (N_19632,N_13173,N_11323);
nand U19633 (N_19633,N_11103,N_11117);
xnor U19634 (N_19634,N_10448,N_10146);
or U19635 (N_19635,N_11313,N_11873);
or U19636 (N_19636,N_11325,N_12085);
nand U19637 (N_19637,N_10299,N_11620);
nand U19638 (N_19638,N_14596,N_13987);
and U19639 (N_19639,N_11111,N_14488);
xor U19640 (N_19640,N_13707,N_12844);
and U19641 (N_19641,N_12445,N_13998);
nand U19642 (N_19642,N_12443,N_14644);
and U19643 (N_19643,N_10786,N_11710);
or U19644 (N_19644,N_11221,N_12249);
nand U19645 (N_19645,N_14619,N_12279);
nand U19646 (N_19646,N_12296,N_10358);
and U19647 (N_19647,N_14371,N_10614);
nor U19648 (N_19648,N_13280,N_11040);
nor U19649 (N_19649,N_12113,N_14009);
nand U19650 (N_19650,N_14221,N_13507);
nand U19651 (N_19651,N_11220,N_11302);
or U19652 (N_19652,N_11184,N_13163);
nand U19653 (N_19653,N_11711,N_14091);
xnor U19654 (N_19654,N_14179,N_11082);
or U19655 (N_19655,N_12503,N_10197);
or U19656 (N_19656,N_11960,N_13891);
nand U19657 (N_19657,N_14084,N_13125);
nor U19658 (N_19658,N_10053,N_10448);
nor U19659 (N_19659,N_12193,N_10027);
nand U19660 (N_19660,N_10016,N_10120);
nor U19661 (N_19661,N_12719,N_14074);
xnor U19662 (N_19662,N_12784,N_12404);
and U19663 (N_19663,N_12577,N_13728);
nand U19664 (N_19664,N_10016,N_14480);
xnor U19665 (N_19665,N_13002,N_11269);
nand U19666 (N_19666,N_11536,N_12021);
or U19667 (N_19667,N_14803,N_14499);
or U19668 (N_19668,N_11778,N_12702);
xor U19669 (N_19669,N_12829,N_10513);
nand U19670 (N_19670,N_11342,N_11861);
and U19671 (N_19671,N_10179,N_13989);
xnor U19672 (N_19672,N_14018,N_14893);
or U19673 (N_19673,N_14438,N_14186);
nand U19674 (N_19674,N_14249,N_14842);
and U19675 (N_19675,N_12614,N_10747);
or U19676 (N_19676,N_12014,N_12634);
and U19677 (N_19677,N_11431,N_12747);
or U19678 (N_19678,N_10176,N_10820);
nor U19679 (N_19679,N_14448,N_14657);
and U19680 (N_19680,N_10939,N_13284);
and U19681 (N_19681,N_13941,N_13751);
nand U19682 (N_19682,N_14849,N_14033);
and U19683 (N_19683,N_11158,N_10710);
nand U19684 (N_19684,N_14199,N_13130);
and U19685 (N_19685,N_13376,N_11906);
or U19686 (N_19686,N_11016,N_12474);
nor U19687 (N_19687,N_12299,N_10658);
and U19688 (N_19688,N_13743,N_14144);
nor U19689 (N_19689,N_14321,N_11293);
nor U19690 (N_19690,N_12335,N_12425);
xor U19691 (N_19691,N_14457,N_14073);
and U19692 (N_19692,N_10410,N_12055);
xnor U19693 (N_19693,N_12453,N_14573);
nand U19694 (N_19694,N_14875,N_10282);
or U19695 (N_19695,N_10153,N_14009);
and U19696 (N_19696,N_10422,N_10697);
or U19697 (N_19697,N_14472,N_10585);
and U19698 (N_19698,N_11494,N_14980);
or U19699 (N_19699,N_12687,N_11036);
or U19700 (N_19700,N_14805,N_10628);
or U19701 (N_19701,N_10680,N_11429);
and U19702 (N_19702,N_14528,N_13965);
or U19703 (N_19703,N_11111,N_10753);
and U19704 (N_19704,N_12821,N_10176);
xnor U19705 (N_19705,N_12172,N_14316);
and U19706 (N_19706,N_14956,N_13489);
or U19707 (N_19707,N_12743,N_13389);
nor U19708 (N_19708,N_14590,N_10339);
nor U19709 (N_19709,N_10453,N_13769);
xnor U19710 (N_19710,N_13426,N_10501);
and U19711 (N_19711,N_14101,N_12775);
or U19712 (N_19712,N_10952,N_13845);
nor U19713 (N_19713,N_13335,N_14880);
nor U19714 (N_19714,N_10530,N_12269);
xor U19715 (N_19715,N_13551,N_13222);
nand U19716 (N_19716,N_11136,N_10639);
xnor U19717 (N_19717,N_12381,N_14621);
or U19718 (N_19718,N_11599,N_10275);
nand U19719 (N_19719,N_11355,N_10658);
and U19720 (N_19720,N_12552,N_10338);
or U19721 (N_19721,N_12225,N_14172);
or U19722 (N_19722,N_12785,N_11034);
nor U19723 (N_19723,N_13080,N_11508);
or U19724 (N_19724,N_12133,N_10183);
nor U19725 (N_19725,N_12097,N_10050);
and U19726 (N_19726,N_14510,N_13627);
or U19727 (N_19727,N_13523,N_11950);
and U19728 (N_19728,N_10459,N_14858);
or U19729 (N_19729,N_11015,N_11902);
or U19730 (N_19730,N_11130,N_14860);
and U19731 (N_19731,N_10803,N_12458);
nand U19732 (N_19732,N_10416,N_10370);
nand U19733 (N_19733,N_11647,N_13754);
nor U19734 (N_19734,N_12094,N_10477);
nor U19735 (N_19735,N_11956,N_11188);
and U19736 (N_19736,N_12617,N_10111);
xor U19737 (N_19737,N_12945,N_12592);
or U19738 (N_19738,N_12628,N_10590);
or U19739 (N_19739,N_10377,N_13865);
and U19740 (N_19740,N_12479,N_12024);
or U19741 (N_19741,N_10185,N_14066);
nor U19742 (N_19742,N_10821,N_13587);
or U19743 (N_19743,N_14401,N_10885);
nand U19744 (N_19744,N_10808,N_14838);
xnor U19745 (N_19745,N_11151,N_10709);
and U19746 (N_19746,N_10216,N_11519);
nand U19747 (N_19747,N_14047,N_11772);
and U19748 (N_19748,N_10590,N_13599);
or U19749 (N_19749,N_12616,N_14955);
and U19750 (N_19750,N_13957,N_13880);
xor U19751 (N_19751,N_10826,N_11473);
nand U19752 (N_19752,N_12337,N_11701);
nand U19753 (N_19753,N_12508,N_12277);
nand U19754 (N_19754,N_12110,N_12703);
and U19755 (N_19755,N_14824,N_10004);
nor U19756 (N_19756,N_13015,N_12060);
and U19757 (N_19757,N_14850,N_14082);
and U19758 (N_19758,N_12536,N_11112);
xnor U19759 (N_19759,N_14152,N_11974);
nand U19760 (N_19760,N_14086,N_14382);
nor U19761 (N_19761,N_13586,N_11032);
or U19762 (N_19762,N_11741,N_13519);
and U19763 (N_19763,N_10020,N_10752);
and U19764 (N_19764,N_10530,N_10597);
xor U19765 (N_19765,N_11647,N_13113);
or U19766 (N_19766,N_12903,N_11210);
xnor U19767 (N_19767,N_12964,N_12800);
and U19768 (N_19768,N_11786,N_11324);
or U19769 (N_19769,N_12456,N_13635);
nand U19770 (N_19770,N_14159,N_12888);
or U19771 (N_19771,N_10130,N_14818);
and U19772 (N_19772,N_11972,N_11981);
nand U19773 (N_19773,N_14209,N_14450);
or U19774 (N_19774,N_14983,N_11350);
nand U19775 (N_19775,N_12821,N_10104);
nand U19776 (N_19776,N_10509,N_11187);
xor U19777 (N_19777,N_14111,N_12803);
nor U19778 (N_19778,N_11884,N_10684);
and U19779 (N_19779,N_12345,N_13341);
and U19780 (N_19780,N_10578,N_10725);
or U19781 (N_19781,N_10532,N_12378);
xnor U19782 (N_19782,N_12433,N_13235);
nand U19783 (N_19783,N_12644,N_12473);
or U19784 (N_19784,N_13859,N_11057);
nand U19785 (N_19785,N_10821,N_13970);
xor U19786 (N_19786,N_14192,N_13938);
nand U19787 (N_19787,N_12368,N_10548);
xnor U19788 (N_19788,N_10000,N_12617);
nand U19789 (N_19789,N_12016,N_12664);
and U19790 (N_19790,N_10320,N_14508);
and U19791 (N_19791,N_12866,N_11718);
or U19792 (N_19792,N_10602,N_11210);
nand U19793 (N_19793,N_13981,N_10866);
nor U19794 (N_19794,N_11366,N_13518);
xor U19795 (N_19795,N_10967,N_14135);
or U19796 (N_19796,N_13115,N_12248);
nand U19797 (N_19797,N_13922,N_12010);
xnor U19798 (N_19798,N_10009,N_14654);
or U19799 (N_19799,N_11194,N_13904);
or U19800 (N_19800,N_13006,N_11667);
or U19801 (N_19801,N_14552,N_12925);
and U19802 (N_19802,N_14740,N_10668);
nor U19803 (N_19803,N_12626,N_10047);
nand U19804 (N_19804,N_12276,N_14028);
and U19805 (N_19805,N_10060,N_11493);
and U19806 (N_19806,N_14998,N_13658);
or U19807 (N_19807,N_13068,N_10221);
nor U19808 (N_19808,N_11388,N_14323);
nor U19809 (N_19809,N_14185,N_10304);
xor U19810 (N_19810,N_12373,N_11071);
and U19811 (N_19811,N_10841,N_12231);
or U19812 (N_19812,N_10559,N_12900);
and U19813 (N_19813,N_11680,N_13242);
nand U19814 (N_19814,N_12773,N_13032);
nand U19815 (N_19815,N_14559,N_11233);
or U19816 (N_19816,N_11793,N_10439);
xnor U19817 (N_19817,N_11406,N_11691);
or U19818 (N_19818,N_14008,N_11304);
nand U19819 (N_19819,N_10478,N_14530);
xor U19820 (N_19820,N_14579,N_13088);
and U19821 (N_19821,N_11052,N_10452);
and U19822 (N_19822,N_12938,N_12603);
or U19823 (N_19823,N_13261,N_13938);
nor U19824 (N_19824,N_11592,N_11605);
nor U19825 (N_19825,N_11289,N_12819);
nor U19826 (N_19826,N_11109,N_11574);
nor U19827 (N_19827,N_14923,N_10673);
or U19828 (N_19828,N_10981,N_11495);
nor U19829 (N_19829,N_11375,N_14452);
nand U19830 (N_19830,N_13717,N_11108);
xnor U19831 (N_19831,N_12763,N_14511);
or U19832 (N_19832,N_14690,N_10855);
or U19833 (N_19833,N_11907,N_13441);
xnor U19834 (N_19834,N_13611,N_11011);
or U19835 (N_19835,N_14018,N_10830);
xnor U19836 (N_19836,N_13988,N_13770);
or U19837 (N_19837,N_12099,N_14763);
nor U19838 (N_19838,N_14962,N_14397);
or U19839 (N_19839,N_11605,N_14856);
and U19840 (N_19840,N_11519,N_10679);
nor U19841 (N_19841,N_12812,N_11641);
nand U19842 (N_19842,N_10038,N_13573);
nand U19843 (N_19843,N_12670,N_11950);
xor U19844 (N_19844,N_13422,N_11527);
or U19845 (N_19845,N_10449,N_10786);
nor U19846 (N_19846,N_10034,N_14608);
xor U19847 (N_19847,N_13224,N_13279);
or U19848 (N_19848,N_13877,N_13746);
or U19849 (N_19849,N_13417,N_10526);
nand U19850 (N_19850,N_12397,N_11592);
and U19851 (N_19851,N_11529,N_10907);
and U19852 (N_19852,N_14880,N_13070);
xor U19853 (N_19853,N_14347,N_10380);
and U19854 (N_19854,N_12258,N_12009);
and U19855 (N_19855,N_14240,N_13987);
xnor U19856 (N_19856,N_14856,N_11358);
nand U19857 (N_19857,N_11490,N_13640);
nand U19858 (N_19858,N_12158,N_13349);
nor U19859 (N_19859,N_11819,N_10721);
nand U19860 (N_19860,N_13006,N_13257);
nand U19861 (N_19861,N_11664,N_14758);
and U19862 (N_19862,N_14702,N_11285);
nand U19863 (N_19863,N_12588,N_12477);
nand U19864 (N_19864,N_13150,N_11111);
and U19865 (N_19865,N_14430,N_13740);
and U19866 (N_19866,N_13644,N_14921);
xor U19867 (N_19867,N_12605,N_10706);
xnor U19868 (N_19868,N_13460,N_10851);
xor U19869 (N_19869,N_12233,N_12370);
xnor U19870 (N_19870,N_10583,N_13133);
nand U19871 (N_19871,N_10588,N_13116);
or U19872 (N_19872,N_11280,N_12710);
or U19873 (N_19873,N_10948,N_10383);
or U19874 (N_19874,N_13102,N_14068);
and U19875 (N_19875,N_13777,N_12261);
nand U19876 (N_19876,N_14665,N_12804);
xnor U19877 (N_19877,N_13648,N_13254);
nand U19878 (N_19878,N_10967,N_13570);
and U19879 (N_19879,N_12989,N_13341);
nor U19880 (N_19880,N_11833,N_13708);
or U19881 (N_19881,N_11356,N_12965);
nor U19882 (N_19882,N_12619,N_13764);
and U19883 (N_19883,N_13758,N_12179);
nor U19884 (N_19884,N_10101,N_12556);
or U19885 (N_19885,N_11118,N_14659);
or U19886 (N_19886,N_13277,N_10177);
nor U19887 (N_19887,N_14014,N_10402);
and U19888 (N_19888,N_12048,N_13982);
or U19889 (N_19889,N_13724,N_11003);
nor U19890 (N_19890,N_11989,N_10401);
and U19891 (N_19891,N_12067,N_14129);
and U19892 (N_19892,N_14495,N_10134);
nand U19893 (N_19893,N_11021,N_14340);
and U19894 (N_19894,N_10159,N_14808);
or U19895 (N_19895,N_12564,N_13028);
xnor U19896 (N_19896,N_10399,N_10704);
nand U19897 (N_19897,N_11274,N_13022);
or U19898 (N_19898,N_11883,N_14800);
nand U19899 (N_19899,N_11336,N_11535);
or U19900 (N_19900,N_14821,N_13177);
or U19901 (N_19901,N_11996,N_13884);
nor U19902 (N_19902,N_10972,N_14528);
nand U19903 (N_19903,N_13259,N_13768);
nor U19904 (N_19904,N_10258,N_10744);
and U19905 (N_19905,N_12158,N_14946);
and U19906 (N_19906,N_12250,N_11315);
nor U19907 (N_19907,N_14654,N_11735);
nor U19908 (N_19908,N_10493,N_13064);
xor U19909 (N_19909,N_13492,N_10200);
xor U19910 (N_19910,N_10919,N_13052);
and U19911 (N_19911,N_14780,N_14351);
nor U19912 (N_19912,N_10450,N_10336);
nand U19913 (N_19913,N_13580,N_10768);
and U19914 (N_19914,N_13401,N_14383);
xor U19915 (N_19915,N_11245,N_14344);
and U19916 (N_19916,N_11218,N_12854);
and U19917 (N_19917,N_10805,N_14180);
xor U19918 (N_19918,N_10569,N_12605);
or U19919 (N_19919,N_10000,N_11209);
nor U19920 (N_19920,N_11717,N_12355);
nor U19921 (N_19921,N_11754,N_11095);
or U19922 (N_19922,N_11114,N_10711);
or U19923 (N_19923,N_13290,N_10250);
and U19924 (N_19924,N_11097,N_10338);
nor U19925 (N_19925,N_13061,N_14403);
nand U19926 (N_19926,N_13331,N_12485);
nand U19927 (N_19927,N_11745,N_13948);
and U19928 (N_19928,N_13888,N_14256);
and U19929 (N_19929,N_13111,N_12786);
and U19930 (N_19930,N_12819,N_12670);
nor U19931 (N_19931,N_13553,N_13901);
or U19932 (N_19932,N_14627,N_11634);
or U19933 (N_19933,N_11885,N_13161);
and U19934 (N_19934,N_14183,N_11284);
xnor U19935 (N_19935,N_12269,N_13744);
nand U19936 (N_19936,N_11808,N_12661);
and U19937 (N_19937,N_13688,N_11735);
nand U19938 (N_19938,N_13041,N_11818);
xor U19939 (N_19939,N_14847,N_12196);
xor U19940 (N_19940,N_12187,N_11879);
xor U19941 (N_19941,N_11868,N_12261);
nor U19942 (N_19942,N_13622,N_11817);
and U19943 (N_19943,N_12382,N_11890);
or U19944 (N_19944,N_10600,N_13680);
nand U19945 (N_19945,N_11290,N_11934);
or U19946 (N_19946,N_13759,N_13632);
or U19947 (N_19947,N_14941,N_10581);
nand U19948 (N_19948,N_12895,N_12865);
nand U19949 (N_19949,N_14300,N_10593);
or U19950 (N_19950,N_12514,N_14592);
nor U19951 (N_19951,N_14190,N_10121);
nor U19952 (N_19952,N_10044,N_13121);
and U19953 (N_19953,N_14883,N_12155);
nor U19954 (N_19954,N_13037,N_11645);
or U19955 (N_19955,N_13859,N_14901);
and U19956 (N_19956,N_11311,N_10750);
nor U19957 (N_19957,N_14486,N_10479);
nor U19958 (N_19958,N_10666,N_13511);
nor U19959 (N_19959,N_10826,N_12189);
xnor U19960 (N_19960,N_10202,N_10388);
xnor U19961 (N_19961,N_13028,N_11727);
nand U19962 (N_19962,N_11553,N_14006);
nand U19963 (N_19963,N_12768,N_13058);
nor U19964 (N_19964,N_11211,N_11243);
nand U19965 (N_19965,N_12229,N_11577);
and U19966 (N_19966,N_10373,N_14647);
and U19967 (N_19967,N_10523,N_11567);
or U19968 (N_19968,N_11842,N_12685);
or U19969 (N_19969,N_13514,N_13027);
nand U19970 (N_19970,N_14529,N_13640);
or U19971 (N_19971,N_10899,N_13512);
and U19972 (N_19972,N_13148,N_13482);
xnor U19973 (N_19973,N_12929,N_10728);
and U19974 (N_19974,N_13748,N_10638);
nor U19975 (N_19975,N_11375,N_10952);
nor U19976 (N_19976,N_10349,N_13584);
xor U19977 (N_19977,N_14128,N_12859);
xor U19978 (N_19978,N_12309,N_14451);
and U19979 (N_19979,N_14136,N_13327);
nand U19980 (N_19980,N_10307,N_10635);
and U19981 (N_19981,N_11503,N_11742);
or U19982 (N_19982,N_11833,N_14227);
or U19983 (N_19983,N_12396,N_12644);
xor U19984 (N_19984,N_11144,N_12559);
or U19985 (N_19985,N_11639,N_13295);
nor U19986 (N_19986,N_14763,N_13138);
xnor U19987 (N_19987,N_12231,N_11214);
and U19988 (N_19988,N_14330,N_10518);
nand U19989 (N_19989,N_13265,N_13363);
or U19990 (N_19990,N_10911,N_13993);
nor U19991 (N_19991,N_12646,N_11042);
xor U19992 (N_19992,N_14398,N_11936);
and U19993 (N_19993,N_13373,N_14250);
nor U19994 (N_19994,N_13438,N_12017);
nand U19995 (N_19995,N_11689,N_13157);
and U19996 (N_19996,N_12393,N_12878);
nor U19997 (N_19997,N_10355,N_10972);
or U19998 (N_19998,N_10227,N_12852);
xnor U19999 (N_19999,N_10368,N_13458);
nor U20000 (N_20000,N_18539,N_18470);
nor U20001 (N_20001,N_16385,N_19955);
and U20002 (N_20002,N_19470,N_16065);
xnor U20003 (N_20003,N_18045,N_15968);
or U20004 (N_20004,N_19813,N_18839);
or U20005 (N_20005,N_17013,N_15216);
nor U20006 (N_20006,N_18869,N_15997);
nand U20007 (N_20007,N_17989,N_15599);
xnor U20008 (N_20008,N_17628,N_16992);
xnor U20009 (N_20009,N_16444,N_19035);
nor U20010 (N_20010,N_15585,N_15377);
nand U20011 (N_20011,N_18873,N_18416);
nor U20012 (N_20012,N_19287,N_17696);
nand U20013 (N_20013,N_19480,N_16538);
xnor U20014 (N_20014,N_16999,N_15623);
and U20015 (N_20015,N_17676,N_19407);
nor U20016 (N_20016,N_15539,N_15615);
or U20017 (N_20017,N_17450,N_15584);
xor U20018 (N_20018,N_16910,N_15261);
nor U20019 (N_20019,N_15163,N_15248);
nor U20020 (N_20020,N_18841,N_15858);
xor U20021 (N_20021,N_15045,N_17811);
xnor U20022 (N_20022,N_16152,N_17318);
xor U20023 (N_20023,N_19171,N_15378);
xnor U20024 (N_20024,N_16080,N_19368);
and U20025 (N_20025,N_16033,N_18546);
or U20026 (N_20026,N_17147,N_16455);
and U20027 (N_20027,N_19796,N_17497);
xnor U20028 (N_20028,N_17342,N_19334);
and U20029 (N_20029,N_18831,N_19843);
nand U20030 (N_20030,N_16762,N_15079);
nor U20031 (N_20031,N_15144,N_18312);
nor U20032 (N_20032,N_17003,N_16774);
nor U20033 (N_20033,N_15200,N_18924);
nand U20034 (N_20034,N_15527,N_16951);
nand U20035 (N_20035,N_17443,N_19645);
xor U20036 (N_20036,N_16682,N_17016);
or U20037 (N_20037,N_16305,N_19747);
nand U20038 (N_20038,N_15767,N_17071);
or U20039 (N_20039,N_19414,N_18610);
and U20040 (N_20040,N_17329,N_15290);
xor U20041 (N_20041,N_17861,N_17365);
nor U20042 (N_20042,N_18528,N_16454);
or U20043 (N_20043,N_16536,N_19246);
or U20044 (N_20044,N_18215,N_15949);
nor U20045 (N_20045,N_19411,N_19807);
xor U20046 (N_20046,N_18932,N_15917);
nor U20047 (N_20047,N_16038,N_15155);
nor U20048 (N_20048,N_15707,N_19136);
and U20049 (N_20049,N_19114,N_15703);
and U20050 (N_20050,N_19526,N_17137);
or U20051 (N_20051,N_16157,N_19100);
nand U20052 (N_20052,N_15728,N_17040);
or U20053 (N_20053,N_16580,N_15920);
and U20054 (N_20054,N_16758,N_19612);
and U20055 (N_20055,N_19544,N_19491);
nor U20056 (N_20056,N_17014,N_16860);
nor U20057 (N_20057,N_19503,N_18378);
nand U20058 (N_20058,N_19628,N_15669);
and U20059 (N_20059,N_17336,N_15908);
xor U20060 (N_20060,N_17974,N_16576);
and U20061 (N_20061,N_15971,N_17713);
and U20062 (N_20062,N_17991,N_18082);
nor U20063 (N_20063,N_16203,N_16153);
xor U20064 (N_20064,N_19932,N_15137);
nand U20065 (N_20065,N_16623,N_18972);
nand U20066 (N_20066,N_16957,N_19513);
or U20067 (N_20067,N_19238,N_19868);
nor U20068 (N_20068,N_16976,N_15025);
xor U20069 (N_20069,N_16832,N_19305);
and U20070 (N_20070,N_17305,N_16589);
nor U20071 (N_20071,N_19964,N_19685);
and U20072 (N_20072,N_17485,N_19935);
nor U20073 (N_20073,N_17021,N_17897);
or U20074 (N_20074,N_16629,N_19773);
nand U20075 (N_20075,N_17019,N_15138);
nand U20076 (N_20076,N_16506,N_17763);
nand U20077 (N_20077,N_17894,N_19852);
or U20078 (N_20078,N_19917,N_17002);
nand U20079 (N_20079,N_17669,N_19610);
and U20080 (N_20080,N_19657,N_16280);
or U20081 (N_20081,N_18171,N_16620);
or U20082 (N_20082,N_19438,N_16074);
or U20083 (N_20083,N_19582,N_15656);
xor U20084 (N_20084,N_19164,N_15307);
nor U20085 (N_20085,N_18785,N_17899);
xor U20086 (N_20086,N_16063,N_17623);
or U20087 (N_20087,N_19719,N_19756);
nor U20088 (N_20088,N_16324,N_18916);
nor U20089 (N_20089,N_17568,N_18217);
nor U20090 (N_20090,N_18468,N_17372);
and U20091 (N_20091,N_19995,N_18783);
and U20092 (N_20092,N_16011,N_17024);
nor U20093 (N_20093,N_19631,N_19370);
xnor U20094 (N_20094,N_19584,N_15999);
nor U20095 (N_20095,N_15485,N_17397);
or U20096 (N_20096,N_18136,N_18524);
or U20097 (N_20097,N_16140,N_18068);
nor U20098 (N_20098,N_18584,N_15477);
and U20099 (N_20099,N_19936,N_19488);
xor U20100 (N_20100,N_19863,N_15816);
and U20101 (N_20101,N_19761,N_15071);
and U20102 (N_20102,N_17709,N_15028);
and U20103 (N_20103,N_17730,N_16487);
xnor U20104 (N_20104,N_15513,N_15122);
nand U20105 (N_20105,N_15186,N_16368);
and U20106 (N_20106,N_17109,N_15791);
xnor U20107 (N_20107,N_19318,N_15826);
or U20108 (N_20108,N_17154,N_16448);
xor U20109 (N_20109,N_18501,N_17398);
or U20110 (N_20110,N_19101,N_15654);
and U20111 (N_20111,N_17087,N_19524);
xor U20112 (N_20112,N_19064,N_18994);
or U20113 (N_20113,N_15713,N_16334);
and U20114 (N_20114,N_16685,N_16907);
xor U20115 (N_20115,N_15630,N_15434);
and U20116 (N_20116,N_15531,N_17630);
and U20117 (N_20117,N_15969,N_15590);
nand U20118 (N_20118,N_17875,N_15575);
nor U20119 (N_20119,N_19426,N_15723);
nor U20120 (N_20120,N_18120,N_16472);
nor U20121 (N_20121,N_16362,N_15745);
and U20122 (N_20122,N_16799,N_17658);
nand U20123 (N_20123,N_18747,N_18991);
xor U20124 (N_20124,N_19730,N_19724);
nor U20125 (N_20125,N_18806,N_18542);
nor U20126 (N_20126,N_15680,N_19835);
nand U20127 (N_20127,N_15677,N_16803);
or U20128 (N_20128,N_15283,N_15674);
nand U20129 (N_20129,N_16676,N_17057);
and U20130 (N_20130,N_15990,N_16414);
nand U20131 (N_20131,N_16081,N_19206);
nand U20132 (N_20132,N_19460,N_19925);
or U20133 (N_20133,N_16888,N_15407);
or U20134 (N_20134,N_18922,N_18687);
and U20135 (N_20135,N_15027,N_17395);
nand U20136 (N_20136,N_15882,N_18335);
or U20137 (N_20137,N_18087,N_19071);
and U20138 (N_20138,N_15646,N_19181);
nand U20139 (N_20139,N_16467,N_18414);
nor U20140 (N_20140,N_19716,N_19344);
nor U20141 (N_20141,N_17490,N_18311);
or U20142 (N_20142,N_18022,N_16619);
nand U20143 (N_20143,N_19261,N_16727);
nor U20144 (N_20144,N_16958,N_15056);
nand U20145 (N_20145,N_19777,N_16489);
and U20146 (N_20146,N_17200,N_18187);
or U20147 (N_20147,N_16230,N_15614);
xor U20148 (N_20148,N_17680,N_16018);
nor U20149 (N_20149,N_15555,N_15102);
and U20150 (N_20150,N_19303,N_19536);
or U20151 (N_20151,N_16687,N_15945);
xor U20152 (N_20152,N_17505,N_15236);
or U20153 (N_20153,N_17053,N_15313);
xnor U20154 (N_20154,N_15251,N_15239);
and U20155 (N_20155,N_16663,N_16630);
nand U20156 (N_20156,N_17994,N_19593);
xor U20157 (N_20157,N_19384,N_17536);
or U20158 (N_20158,N_18974,N_16402);
and U20159 (N_20159,N_17161,N_18132);
nor U20160 (N_20160,N_17741,N_17525);
nand U20161 (N_20161,N_18700,N_19403);
nand U20162 (N_20162,N_17463,N_16292);
xnor U20163 (N_20163,N_16656,N_19622);
nor U20164 (N_20164,N_19643,N_15347);
nand U20165 (N_20165,N_19754,N_15503);
and U20166 (N_20166,N_18119,N_18802);
nand U20167 (N_20167,N_15124,N_18837);
xnor U20168 (N_20168,N_16673,N_16932);
xor U20169 (N_20169,N_19882,N_18977);
and U20170 (N_20170,N_18336,N_17093);
or U20171 (N_20171,N_15299,N_17364);
xnor U20172 (N_20172,N_18562,N_19375);
and U20173 (N_20173,N_15288,N_16131);
xor U20174 (N_20174,N_16555,N_15602);
nand U20175 (N_20175,N_18233,N_17130);
nand U20176 (N_20176,N_19120,N_15325);
xnor U20177 (N_20177,N_16405,N_18784);
nand U20178 (N_20178,N_18611,N_16597);
or U20179 (N_20179,N_19721,N_19710);
nor U20180 (N_20180,N_16343,N_19940);
xnor U20181 (N_20181,N_19523,N_15571);
or U20182 (N_20182,N_18526,N_18163);
nand U20183 (N_20183,N_19011,N_17564);
and U20184 (N_20184,N_15569,N_18790);
xnor U20185 (N_20185,N_17357,N_19758);
nand U20186 (N_20186,N_19728,N_19680);
and U20187 (N_20187,N_15900,N_16376);
xor U20188 (N_20188,N_19097,N_18895);
xor U20189 (N_20189,N_17784,N_17675);
or U20190 (N_20190,N_17958,N_15712);
xnor U20191 (N_20191,N_15100,N_18091);
nand U20192 (N_20192,N_17070,N_19629);
or U20193 (N_20193,N_15755,N_18502);
or U20194 (N_20194,N_17690,N_18951);
or U20195 (N_20195,N_16779,N_18061);
nand U20196 (N_20196,N_18670,N_19881);
and U20197 (N_20197,N_16425,N_17338);
nor U20198 (N_20198,N_17399,N_19175);
xor U20199 (N_20199,N_19787,N_18992);
or U20200 (N_20200,N_17387,N_19354);
and U20201 (N_20201,N_16077,N_18813);
and U20202 (N_20202,N_17551,N_18999);
xnor U20203 (N_20203,N_19128,N_17725);
or U20204 (N_20204,N_17777,N_19086);
and U20205 (N_20205,N_16450,N_17805);
and U20206 (N_20206,N_18430,N_16916);
nor U20207 (N_20207,N_15074,N_16996);
nand U20208 (N_20208,N_15692,N_16792);
nor U20209 (N_20209,N_19567,N_18791);
or U20210 (N_20210,N_16883,N_19782);
xnor U20211 (N_20211,N_19732,N_16549);
nand U20212 (N_20212,N_17442,N_17686);
and U20213 (N_20213,N_19008,N_18173);
or U20214 (N_20214,N_16045,N_19684);
or U20215 (N_20215,N_15478,N_16980);
or U20216 (N_20216,N_16151,N_16849);
or U20217 (N_20217,N_16309,N_15683);
xor U20218 (N_20218,N_17931,N_17256);
and U20219 (N_20219,N_17662,N_15603);
nor U20220 (N_20220,N_18967,N_16606);
nand U20221 (N_20221,N_18570,N_16784);
nand U20222 (N_20222,N_19545,N_16584);
xor U20223 (N_20223,N_15551,N_17473);
or U20224 (N_20224,N_19751,N_17144);
or U20225 (N_20225,N_16610,N_15068);
xor U20226 (N_20226,N_17755,N_15145);
nor U20227 (N_20227,N_18385,N_16732);
and U20228 (N_20228,N_17884,N_15730);
or U20229 (N_20229,N_19030,N_16514);
xnor U20230 (N_20230,N_15229,N_18266);
nand U20231 (N_20231,N_15412,N_19691);
or U20232 (N_20232,N_17007,N_16987);
nor U20233 (N_20233,N_19801,N_19866);
nand U20234 (N_20234,N_16880,N_19976);
or U20235 (N_20235,N_19639,N_19337);
xor U20236 (N_20236,N_16332,N_19946);
nor U20237 (N_20237,N_16276,N_17795);
or U20238 (N_20238,N_15387,N_17332);
xor U20239 (N_20239,N_15212,N_16299);
nand U20240 (N_20240,N_16041,N_16679);
or U20241 (N_20241,N_17539,N_19439);
xnor U20242 (N_20242,N_19648,N_18966);
and U20243 (N_20243,N_19587,N_15168);
nor U20244 (N_20244,N_18681,N_16139);
nor U20245 (N_20245,N_15470,N_16884);
and U20246 (N_20246,N_17436,N_17376);
xor U20247 (N_20247,N_19376,N_16782);
xnor U20248 (N_20248,N_18505,N_19799);
and U20249 (N_20249,N_15314,N_19937);
and U20250 (N_20250,N_17842,N_17594);
or U20251 (N_20251,N_15413,N_15780);
nor U20252 (N_20252,N_15764,N_19229);
and U20253 (N_20253,N_17191,N_16190);
or U20254 (N_20254,N_17258,N_17150);
or U20255 (N_20255,N_17638,N_18619);
xnor U20256 (N_20256,N_17892,N_18483);
xnor U20257 (N_20257,N_16858,N_16434);
and U20258 (N_20258,N_16941,N_19283);
nor U20259 (N_20259,N_16703,N_15397);
or U20260 (N_20260,N_19196,N_19722);
nand U20261 (N_20261,N_17544,N_17723);
nand U20262 (N_20262,N_16517,N_15828);
nand U20263 (N_20263,N_17674,N_17791);
or U20264 (N_20264,N_15833,N_19059);
or U20265 (N_20265,N_16210,N_18674);
nor U20266 (N_20266,N_15037,N_17997);
and U20267 (N_20267,N_19474,N_18073);
nor U20268 (N_20268,N_19633,N_15177);
nand U20269 (N_20269,N_18693,N_17523);
nand U20270 (N_20270,N_15847,N_16834);
or U20271 (N_20271,N_19615,N_19386);
xor U20272 (N_20272,N_18487,N_17467);
xor U20273 (N_20273,N_16918,N_17996);
nand U20274 (N_20274,N_18117,N_15912);
xnor U20275 (N_20275,N_17211,N_18309);
nor U20276 (N_20276,N_16613,N_15560);
nand U20277 (N_20277,N_18124,N_15794);
and U20278 (N_20278,N_16924,N_16962);
nand U20279 (N_20279,N_15936,N_17289);
nor U20280 (N_20280,N_18050,N_18686);
and U20281 (N_20281,N_17684,N_19806);
nor U20282 (N_20282,N_17390,N_18495);
and U20283 (N_20283,N_16241,N_16618);
nand U20284 (N_20284,N_17330,N_18098);
nor U20285 (N_20285,N_16218,N_16412);
nand U20286 (N_20286,N_17835,N_19489);
nand U20287 (N_20287,N_15052,N_16684);
or U20288 (N_20288,N_17728,N_17660);
xor U20289 (N_20289,N_19451,N_15367);
nand U20290 (N_20290,N_15655,N_19583);
xnor U20291 (N_20291,N_18758,N_18834);
nand U20292 (N_20292,N_17817,N_19404);
xnor U20293 (N_20293,N_15771,N_17361);
and U20294 (N_20294,N_16671,N_19281);
xnor U20295 (N_20295,N_15662,N_15320);
xor U20296 (N_20296,N_17718,N_19152);
nand U20297 (N_20297,N_19034,N_19585);
or U20298 (N_20298,N_15208,N_18439);
nand U20299 (N_20299,N_16361,N_15979);
or U20300 (N_20300,N_16718,N_19016);
xor U20301 (N_20301,N_15597,N_16668);
xnor U20302 (N_20302,N_19186,N_15734);
or U20303 (N_20303,N_19767,N_15849);
or U20304 (N_20304,N_19714,N_16905);
and U20305 (N_20305,N_19840,N_17032);
nor U20306 (N_20306,N_16625,N_16097);
and U20307 (N_20307,N_17550,N_17136);
or U20308 (N_20308,N_18053,N_18923);
nor U20309 (N_20309,N_17752,N_16300);
xor U20310 (N_20310,N_17993,N_15241);
nand U20311 (N_20311,N_19592,N_17980);
nand U20312 (N_20312,N_19613,N_16944);
nand U20313 (N_20313,N_15386,N_19626);
nor U20314 (N_20314,N_18874,N_18765);
xor U20315 (N_20315,N_18718,N_16936);
nor U20316 (N_20316,N_15902,N_18452);
and U20317 (N_20317,N_15639,N_17122);
and U20318 (N_20318,N_17115,N_19820);
or U20319 (N_20319,N_16662,N_17942);
xor U20320 (N_20320,N_19233,N_16461);
xnor U20321 (N_20321,N_16633,N_15157);
nor U20322 (N_20322,N_16103,N_18382);
nand U20323 (N_20323,N_15850,N_17542);
or U20324 (N_20324,N_18126,N_16469);
and U20325 (N_20325,N_15810,N_15040);
nand U20326 (N_20326,N_17411,N_16008);
nor U20327 (N_20327,N_19462,N_16503);
xnor U20328 (N_20328,N_16837,N_17691);
and U20329 (N_20329,N_15974,N_15043);
and U20330 (N_20330,N_18981,N_15537);
or U20331 (N_20331,N_18504,N_16123);
xnor U20332 (N_20332,N_15237,N_17646);
nor U20333 (N_20333,N_19464,N_15983);
xor U20334 (N_20334,N_18310,N_16548);
nand U20335 (N_20335,N_17149,N_19923);
nor U20336 (N_20336,N_19506,N_16573);
xnor U20337 (N_20337,N_18847,N_19704);
xor U20338 (N_20338,N_19252,N_19830);
or U20339 (N_20339,N_19699,N_17017);
nand U20340 (N_20340,N_19191,N_16430);
nand U20341 (N_20341,N_15581,N_15250);
nor U20342 (N_20342,N_17471,N_19504);
nand U20343 (N_20343,N_18804,N_18095);
and U20344 (N_20344,N_17821,N_19423);
nand U20345 (N_20345,N_18664,N_19793);
nand U20346 (N_20346,N_19039,N_15532);
xor U20347 (N_20347,N_19216,N_15587);
or U20348 (N_20348,N_17693,N_15107);
and U20349 (N_20349,N_16410,N_18386);
and U20350 (N_20350,N_19380,N_17293);
nand U20351 (N_20351,N_16350,N_15789);
xor U20352 (N_20352,N_17502,N_17706);
or U20353 (N_20353,N_15890,N_15670);
xnor U20354 (N_20354,N_16759,N_15883);
xnor U20355 (N_20355,N_15973,N_17212);
xnor U20356 (N_20356,N_17801,N_17670);
nand U20357 (N_20357,N_15061,N_19597);
and U20358 (N_20358,N_19262,N_19212);
and U20359 (N_20359,N_19372,N_19397);
xor U20360 (N_20360,N_18011,N_19405);
nor U20361 (N_20361,N_16114,N_18551);
xnor U20362 (N_20362,N_17378,N_15848);
nand U20363 (N_20363,N_18734,N_19307);
xnor U20364 (N_20364,N_15775,N_15516);
xnor U20365 (N_20365,N_17027,N_16771);
and U20366 (N_20366,N_17533,N_18942);
nor U20367 (N_20367,N_17822,N_15731);
nor U20368 (N_20368,N_15295,N_15473);
nand U20369 (N_20369,N_16565,N_18778);
nor U20370 (N_20370,N_15171,N_16886);
nand U20371 (N_20371,N_16856,N_19176);
nor U20372 (N_20372,N_17046,N_18421);
and U20373 (N_20373,N_15484,N_19831);
xnor U20374 (N_20374,N_16796,N_15547);
xnor U20375 (N_20375,N_15091,N_17699);
or U20376 (N_20376,N_16498,N_16829);
nor U20377 (N_20377,N_18541,N_17766);
and U20378 (N_20378,N_16465,N_18531);
nor U20379 (N_20379,N_18808,N_18027);
nor U20380 (N_20380,N_16721,N_18287);
xnor U20381 (N_20381,N_19910,N_18958);
or U20382 (N_20382,N_16559,N_18580);
or U20383 (N_20383,N_18746,N_17422);
and U20384 (N_20384,N_19740,N_18592);
nand U20385 (N_20385,N_19668,N_19260);
nand U20386 (N_20386,N_19056,N_18017);
or U20387 (N_20387,N_15181,N_17298);
nor U20388 (N_20388,N_18314,N_15266);
xnor U20389 (N_20389,N_17162,N_19124);
nand U20390 (N_20390,N_15032,N_18853);
nand U20391 (N_20391,N_15020,N_15586);
nor U20392 (N_20392,N_15658,N_15489);
xnor U20393 (N_20393,N_19891,N_18169);
or U20394 (N_20394,N_19990,N_16372);
or U20395 (N_20395,N_16272,N_17034);
nor U20396 (N_20396,N_17010,N_16838);
xnor U20397 (N_20397,N_17559,N_18275);
nand U20398 (N_20398,N_16326,N_16695);
nor U20399 (N_20399,N_19416,N_18366);
nor U20400 (N_20400,N_19485,N_16240);
xor U20401 (N_20401,N_15273,N_17300);
xnor U20402 (N_20402,N_15928,N_19836);
xor U20403 (N_20403,N_18222,N_17850);
and U20404 (N_20404,N_19515,N_17327);
nand U20405 (N_20405,N_16313,N_19422);
xor U20406 (N_20406,N_15886,N_18845);
xor U20407 (N_20407,N_18571,N_17023);
xnor U20408 (N_20408,N_19708,N_16669);
nand U20409 (N_20409,N_16228,N_18021);
or U20410 (N_20410,N_18690,N_17851);
and U20411 (N_20411,N_16383,N_18517);
xor U20412 (N_20412,N_18202,N_17350);
and U20413 (N_20413,N_18697,N_15258);
and U20414 (N_20414,N_19824,N_17654);
and U20415 (N_20415,N_17114,N_19289);
nand U20416 (N_20416,N_15776,N_15704);
nand U20417 (N_20417,N_18710,N_18934);
xor U20418 (N_20418,N_15952,N_17223);
xor U20419 (N_20419,N_17841,N_18106);
xor U20420 (N_20420,N_15829,N_15519);
or U20421 (N_20421,N_19096,N_19429);
nor U20422 (N_20422,N_18211,N_16814);
or U20423 (N_20423,N_19872,N_16302);
or U20424 (N_20424,N_16652,N_16076);
nor U20425 (N_20425,N_17274,N_16010);
nor U20426 (N_20426,N_19977,N_18828);
or U20427 (N_20427,N_16509,N_16855);
nor U20428 (N_20428,N_17260,N_18015);
or U20429 (N_20429,N_17006,N_16972);
and U20430 (N_20430,N_16994,N_17165);
nand U20431 (N_20431,N_17516,N_15717);
or U20432 (N_20432,N_16919,N_18434);
nand U20433 (N_20433,N_18070,N_16527);
and U20434 (N_20434,N_15189,N_16053);
xor U20435 (N_20435,N_17175,N_18812);
nor U20436 (N_20436,N_15401,N_16601);
nand U20437 (N_20437,N_19173,N_18466);
or U20438 (N_20438,N_17396,N_18985);
and U20439 (N_20439,N_17343,N_17059);
or U20440 (N_20440,N_17952,N_15588);
or U20441 (N_20441,N_19142,N_17880);
or U20442 (N_20442,N_16128,N_15946);
or U20443 (N_20443,N_15598,N_17197);
and U20444 (N_20444,N_15763,N_19285);
nor U20445 (N_20445,N_19017,N_17311);
nor U20446 (N_20446,N_18346,N_17173);
or U20447 (N_20447,N_17220,N_16520);
nor U20448 (N_20448,N_19562,N_18658);
and U20449 (N_20449,N_15203,N_18491);
and U20450 (N_20450,N_16483,N_18372);
xor U20451 (N_20451,N_18267,N_18576);
nor U20452 (N_20452,N_17814,N_19107);
nand U20453 (N_20453,N_17417,N_17043);
and U20454 (N_20454,N_18425,N_15404);
or U20455 (N_20455,N_16524,N_18716);
nor U20456 (N_20456,N_15440,N_18970);
xnor U20457 (N_20457,N_19550,N_17116);
nor U20458 (N_20458,N_18055,N_19218);
or U20459 (N_20459,N_18135,N_15350);
nand U20460 (N_20460,N_16438,N_16104);
nand U20461 (N_20461,N_15305,N_15753);
or U20462 (N_20462,N_16009,N_19131);
or U20463 (N_20463,N_18067,N_18506);
and U20464 (N_20464,N_15123,N_17836);
or U20465 (N_20465,N_17748,N_17827);
nand U20466 (N_20466,N_15741,N_19486);
nor U20467 (N_20467,N_16585,N_16188);
nand U20468 (N_20468,N_16870,N_18455);
xnor U20469 (N_20469,N_15962,N_18997);
nor U20470 (N_20470,N_15933,N_16787);
nand U20471 (N_20471,N_18076,N_19087);
nand U20472 (N_20472,N_19805,N_15989);
xor U20473 (N_20473,N_18249,N_15301);
or U20474 (N_20474,N_17058,N_17425);
and U20475 (N_20475,N_15904,N_17346);
xor U20476 (N_20476,N_17248,N_17129);
nand U20477 (N_20477,N_18442,N_18162);
xor U20478 (N_20478,N_18210,N_17983);
and U20479 (N_20479,N_15214,N_18380);
nand U20480 (N_20480,N_15994,N_19395);
and U20481 (N_20481,N_15732,N_15866);
and U20482 (N_20482,N_18890,N_19869);
nand U20483 (N_20483,N_18298,N_16712);
and U20484 (N_20484,N_17595,N_19983);
or U20485 (N_20485,N_19032,N_18000);
xor U20486 (N_20486,N_18767,N_17054);
or U20487 (N_20487,N_18292,N_18678);
and U20488 (N_20488,N_19814,N_15672);
and U20489 (N_20489,N_16205,N_18855);
and U20490 (N_20490,N_19897,N_17769);
and U20491 (N_20491,N_17100,N_15084);
xnor U20492 (N_20492,N_16437,N_19809);
and U20493 (N_20493,N_16426,N_19599);
xnor U20494 (N_20494,N_15106,N_16797);
nor U20495 (N_20495,N_15249,N_16657);
xnor U20496 (N_20496,N_17048,N_19076);
nor U20497 (N_20497,N_18766,N_18278);
or U20498 (N_20498,N_19466,N_17353);
xor U20499 (N_20499,N_18586,N_15768);
xnor U20500 (N_20500,N_17571,N_19343);
xnor U20501 (N_20501,N_19505,N_18982);
and U20502 (N_20502,N_19884,N_19788);
and U20503 (N_20503,N_19664,N_19853);
nor U20504 (N_20504,N_18259,N_17873);
nor U20505 (N_20505,N_16260,N_19092);
or U20506 (N_20506,N_19590,N_16885);
nor U20507 (N_20507,N_15524,N_19447);
or U20508 (N_20508,N_17039,N_16126);
nor U20509 (N_20509,N_17352,N_15365);
or U20510 (N_20510,N_17830,N_18519);
and U20511 (N_20511,N_17751,N_15869);
nand U20512 (N_20512,N_19484,N_17905);
nand U20513 (N_20513,N_19851,N_15951);
xnor U20514 (N_20514,N_15133,N_18446);
nand U20515 (N_20515,N_15443,N_15363);
xnor U20516 (N_20516,N_18324,N_17874);
or U20517 (N_20517,N_18428,N_16215);
nand U20518 (N_20518,N_18028,N_19356);
nor U20519 (N_20519,N_18500,N_19298);
nor U20520 (N_20520,N_15538,N_17299);
xnor U20521 (N_20521,N_15051,N_15835);
xor U20522 (N_20522,N_15998,N_15319);
nand U20523 (N_20523,N_17694,N_17080);
and U20524 (N_20524,N_19887,N_19069);
or U20525 (N_20525,N_16716,N_18926);
xnor U20526 (N_20526,N_15259,N_17733);
nor U20527 (N_20527,N_15981,N_18364);
xnor U20528 (N_20528,N_19725,N_18656);
or U20529 (N_20529,N_19689,N_17518);
nor U20530 (N_20530,N_16529,N_17714);
nand U20531 (N_20531,N_17852,N_19538);
and U20532 (N_20532,N_16544,N_19510);
nand U20533 (N_20533,N_18387,N_16692);
and U20534 (N_20534,N_15129,N_17253);
and U20535 (N_20535,N_16165,N_15182);
nor U20536 (N_20536,N_18702,N_15023);
xor U20537 (N_20537,N_19205,N_15867);
and U20538 (N_20538,N_15269,N_15684);
nor U20539 (N_20539,N_15198,N_19771);
and U20540 (N_20540,N_19312,N_15552);
nand U20541 (N_20541,N_15408,N_19197);
xnor U20542 (N_20542,N_16281,N_16058);
nand U20543 (N_20543,N_17572,N_19810);
or U20544 (N_20544,N_18108,N_15879);
and U20545 (N_20545,N_19862,N_15240);
nor U20546 (N_20546,N_17409,N_16666);
xnor U20547 (N_20547,N_17610,N_18559);
nor U20548 (N_20548,N_18764,N_17849);
xnor U20549 (N_20549,N_16678,N_18859);
nor U20550 (N_20550,N_17224,N_16826);
nand U20551 (N_20551,N_15148,N_15380);
xnor U20552 (N_20552,N_16765,N_17885);
or U20553 (N_20553,N_15798,N_16558);
or U20554 (N_20554,N_16744,N_15687);
nand U20555 (N_20555,N_18722,N_19314);
nand U20556 (N_20556,N_18730,N_16468);
and U20557 (N_20557,N_16198,N_15545);
or U20558 (N_20558,N_18071,N_17038);
and U20559 (N_20559,N_16966,N_16757);
nand U20560 (N_20560,N_18821,N_17470);
or U20561 (N_20561,N_15757,N_15366);
or U20562 (N_20562,N_17992,N_18188);
nand U20563 (N_20563,N_18078,N_19280);
xnor U20564 (N_20564,N_17567,N_15151);
nor U20565 (N_20565,N_15409,N_16377);
and U20566 (N_20566,N_19687,N_19251);
xor U20567 (N_20567,N_16382,N_18713);
xnor U20568 (N_20568,N_18373,N_17217);
xor U20569 (N_20569,N_17612,N_18776);
nand U20570 (N_20570,N_15842,N_19569);
nand U20571 (N_20571,N_16533,N_18342);
and U20572 (N_20572,N_16381,N_17112);
or U20573 (N_20573,N_15101,N_19046);
xor U20574 (N_20574,N_18822,N_16902);
nor U20575 (N_20575,N_17934,N_15851);
and U20576 (N_20576,N_17587,N_18737);
xor U20577 (N_20577,N_19037,N_15751);
or U20578 (N_20578,N_19768,N_15153);
or U20579 (N_20579,N_19053,N_17643);
and U20580 (N_20580,N_16583,N_17131);
nand U20581 (N_20581,N_15834,N_17500);
or U20582 (N_20582,N_16869,N_16031);
nand U20583 (N_20583,N_18885,N_19007);
or U20584 (N_20584,N_15131,N_16396);
and U20585 (N_20585,N_19507,N_16602);
nor U20586 (N_20586,N_15113,N_18411);
or U20587 (N_20587,N_16802,N_15651);
and U20588 (N_20588,N_15690,N_19928);
or U20589 (N_20589,N_19079,N_15726);
nand U20590 (N_20590,N_17616,N_17349);
and U20591 (N_20591,N_19461,N_15536);
nor U20592 (N_20592,N_19641,N_17186);
and U20593 (N_20593,N_18300,N_18864);
nand U20594 (N_20594,N_18789,N_18626);
nor U20595 (N_20595,N_18695,N_16518);
nand U20596 (N_20596,N_17192,N_19988);
xnor U20597 (N_20597,N_19457,N_16605);
nand U20598 (N_20598,N_17291,N_19847);
xnor U20599 (N_20599,N_15311,N_15224);
nand U20600 (N_20600,N_18630,N_16255);
and U20601 (N_20601,N_17132,N_17066);
and U20602 (N_20602,N_17799,N_18995);
nand U20603 (N_20603,N_16794,N_18523);
nor U20604 (N_20604,N_16761,N_17432);
or U20605 (N_20605,N_16160,N_16864);
nor U20606 (N_20606,N_16421,N_17069);
xnor U20607 (N_20607,N_16286,N_17273);
and U20608 (N_20608,N_16661,N_18435);
nand U20609 (N_20609,N_15761,N_18892);
xnor U20610 (N_20610,N_19103,N_18181);
xnor U20611 (N_20611,N_18388,N_19004);
and U20612 (N_20612,N_15736,N_15119);
xnor U20613 (N_20613,N_17499,N_17966);
or U20614 (N_20614,N_18303,N_18963);
xnor U20615 (N_20615,N_18616,N_16315);
nor U20616 (N_20616,N_15553,N_18679);
nor U20617 (N_20617,N_18887,N_17240);
nor U20618 (N_20618,N_16609,N_18140);
and U20619 (N_20619,N_18602,N_15659);
nor U20620 (N_20620,N_15395,N_15169);
and U20621 (N_20621,N_17284,N_15083);
xnor U20622 (N_20622,N_15749,N_16889);
nor U20623 (N_20623,N_18420,N_19123);
or U20624 (N_20624,N_15450,N_18396);
xnor U20625 (N_20625,N_17474,N_15081);
nor U20626 (N_20626,N_17356,N_19134);
xor U20627 (N_20627,N_19126,N_19834);
and U20628 (N_20628,N_19903,N_18127);
nor U20629 (N_20629,N_19640,N_17201);
nand U20630 (N_20630,N_17648,N_17534);
nand U20631 (N_20631,N_17645,N_17995);
xor U20632 (N_20632,N_19496,N_15748);
nand U20633 (N_20633,N_15573,N_18075);
or U20634 (N_20634,N_18458,N_18949);
or U20635 (N_20635,N_17742,N_17492);
nor U20636 (N_20636,N_17872,N_18406);
and U20637 (N_20637,N_18605,N_17444);
nand U20638 (N_20638,N_16392,N_15661);
and U20639 (N_20639,N_17011,N_18796);
and U20640 (N_20640,N_17985,N_17925);
nor U20641 (N_20641,N_15293,N_19268);
and U20642 (N_20642,N_16277,N_17092);
nand U20643 (N_20643,N_18521,N_19325);
or U20644 (N_20644,N_16102,N_18877);
and U20645 (N_20645,N_15410,N_15419);
nand U20646 (N_20646,N_17782,N_15760);
nand U20647 (N_20647,N_17018,N_17780);
and U20648 (N_20648,N_18212,N_18613);
and U20649 (N_20649,N_19189,N_18260);
nand U20650 (N_20650,N_18564,N_17581);
and U20651 (N_20651,N_15967,N_18587);
nand U20652 (N_20652,N_17824,N_16419);
nor U20653 (N_20653,N_18805,N_16263);
xnor U20654 (N_20654,N_15925,N_16923);
and U20655 (N_20655,N_18072,N_16232);
and U20656 (N_20656,N_18080,N_15063);
nor U20657 (N_20657,N_19045,N_19763);
or U20658 (N_20658,N_18047,N_19815);
nor U20659 (N_20659,N_16824,N_15953);
xor U20660 (N_20660,N_15217,N_19437);
or U20661 (N_20661,N_19345,N_17839);
nor U20662 (N_20662,N_19812,N_16681);
nand U20663 (N_20663,N_15353,N_16775);
nand U20664 (N_20664,N_15505,N_16470);
nand U20665 (N_20665,N_19455,N_16737);
or U20666 (N_20666,N_18284,N_15230);
xor U20667 (N_20667,N_16526,N_17609);
and U20668 (N_20668,N_18069,N_19705);
nand U20669 (N_20669,N_15304,N_17319);
and U20670 (N_20670,N_15285,N_15055);
xnor U20671 (N_20671,N_17077,N_16516);
nor U20672 (N_20672,N_16931,N_18285);
nand U20673 (N_20673,N_15392,N_17237);
nor U20674 (N_20674,N_16603,N_16129);
and U20675 (N_20675,N_15490,N_19446);
xnor U20676 (N_20676,N_16863,N_16604);
nand U20677 (N_20677,N_15558,N_17933);
and U20678 (N_20678,N_18755,N_18394);
and U20679 (N_20679,N_17056,N_15093);
or U20680 (N_20680,N_15574,N_16819);
nand U20681 (N_20681,N_18280,N_18946);
nand U20682 (N_20682,N_16801,N_17367);
xor U20683 (N_20683,N_18800,N_17494);
nor U20684 (N_20684,N_15117,N_19912);
or U20685 (N_20685,N_17895,N_17047);
and U20686 (N_20686,N_18301,N_15825);
xor U20687 (N_20687,N_15164,N_17401);
nand U20688 (N_20688,N_19434,N_15624);
or U20689 (N_20689,N_17668,N_16116);
nor U20690 (N_20690,N_18883,N_16812);
and U20691 (N_20691,N_15156,N_18354);
nor U20692 (N_20692,N_16688,N_17927);
or U20693 (N_20693,N_17959,N_19533);
nor U20694 (N_20694,N_17914,N_17796);
xor U20695 (N_20695,N_16346,N_16659);
nor U20696 (N_20696,N_19141,N_19794);
or U20697 (N_20697,N_17265,N_18793);
or U20698 (N_20698,N_15872,N_17266);
nand U20699 (N_20699,N_15103,N_15406);
or U20700 (N_20700,N_16279,N_19770);
nor U20701 (N_20701,N_18832,N_19207);
xnor U20702 (N_20702,N_17855,N_19358);
nand U20703 (N_20703,N_16357,N_15195);
nand U20704 (N_20704,N_16773,N_18925);
or U20705 (N_20705,N_15725,N_16841);
xnor U20706 (N_20706,N_15664,N_17252);
xor U20707 (N_20707,N_19537,N_17570);
nand U20708 (N_20708,N_16294,N_16347);
xnor U20709 (N_20709,N_19062,N_17174);
or U20710 (N_20710,N_18735,N_19558);
xnor U20711 (N_20711,N_19232,N_19182);
and U20712 (N_20712,N_19540,N_15213);
and U20713 (N_20713,N_15403,N_15557);
and U20714 (N_20714,N_17177,N_19019);
and U20715 (N_20715,N_16393,N_15604);
nand U20716 (N_20716,N_15220,N_18178);
nand U20717 (N_20717,N_17560,N_18990);
or U20718 (N_20718,N_18773,N_18961);
nand U20719 (N_20719,N_16482,N_19832);
nand U20720 (N_20720,N_19146,N_16127);
or U20721 (N_20721,N_18228,N_16048);
nor U20722 (N_20722,N_19906,N_19731);
nor U20723 (N_20723,N_17717,N_17012);
xnor U20724 (N_20724,N_19105,N_17281);
or U20725 (N_20725,N_16865,N_19255);
and U20726 (N_20726,N_18692,N_17182);
xor U20727 (N_20727,N_19642,N_19225);
xor U20728 (N_20728,N_17477,N_18928);
nand U20729 (N_20729,N_19137,N_19154);
nand U20730 (N_20730,N_19893,N_15263);
or U20731 (N_20731,N_18572,N_18084);
xor U20732 (N_20732,N_17898,N_15328);
or U20733 (N_20733,N_17277,N_15095);
or U20734 (N_20734,N_16575,N_16861);
xor U20735 (N_20735,N_19185,N_19674);
xor U20736 (N_20736,N_16823,N_15041);
or U20737 (N_20737,N_16406,N_17125);
nor U20738 (N_20738,N_16082,N_15002);
xnor U20739 (N_20739,N_16106,N_15278);
and U20740 (N_20740,N_19493,N_17716);
and U20741 (N_20741,N_19651,N_16254);
xnor U20742 (N_20742,N_15058,N_15750);
or U20743 (N_20743,N_15509,N_18851);
nor U20744 (N_20744,N_16531,N_16990);
or U20745 (N_20745,N_16701,N_18540);
and U20746 (N_20746,N_18365,N_17119);
xor U20747 (N_20747,N_19905,N_16170);
nor U20748 (N_20748,N_18440,N_18332);
nor U20749 (N_20749,N_18279,N_19098);
xnor U20750 (N_20750,N_17403,N_17437);
and U20751 (N_20751,N_16278,N_17910);
xor U20752 (N_20752,N_15905,N_19821);
and U20753 (N_20753,N_19023,N_15451);
or U20754 (N_20754,N_16284,N_17635);
xnor U20755 (N_20755,N_15801,N_16267);
and U20756 (N_20756,N_16237,N_17591);
nor U20757 (N_20757,N_16754,N_19571);
or U20758 (N_20758,N_18915,N_16379);
or U20759 (N_20759,N_16147,N_18558);
or U20760 (N_20760,N_19965,N_17649);
xnor U20761 (N_20761,N_15329,N_15582);
and U20762 (N_20762,N_18936,N_15746);
or U20763 (N_20763,N_16562,N_18633);
or U20764 (N_20764,N_18971,N_15863);
and U20765 (N_20765,N_16177,N_16341);
nand U20766 (N_20766,N_15836,N_16474);
nand U20767 (N_20767,N_17615,N_15517);
xnor U20768 (N_20768,N_15567,N_16789);
xnor U20769 (N_20769,N_15903,N_15689);
or U20770 (N_20770,N_17810,N_17903);
or U20771 (N_20771,N_19290,N_16769);
nor U20772 (N_20772,N_17164,N_18062);
or U20773 (N_20773,N_19351,N_17541);
or U20774 (N_20774,N_18103,N_16952);
nand U20775 (N_20775,N_19187,N_18515);
nor U20776 (N_20776,N_15035,N_16499);
or U20777 (N_20777,N_18927,N_15650);
nand U20778 (N_20778,N_18221,N_18433);
nor U20779 (N_20779,N_16920,N_19644);
xnor U20780 (N_20780,N_18473,N_17720);
nor U20781 (N_20781,N_17657,N_17341);
or U20782 (N_20782,N_19286,N_18732);
or U20783 (N_20783,N_15108,N_19837);
and U20784 (N_20784,N_15772,N_17377);
and U20785 (N_20785,N_17445,N_18561);
nor U20786 (N_20786,N_16098,N_17360);
xnor U20787 (N_20787,N_17563,N_15402);
nand U20788 (N_20788,N_18123,N_18413);
nor U20789 (N_20789,N_15488,N_17067);
nand U20790 (N_20790,N_17960,N_18968);
xnor U20791 (N_20791,N_17844,N_18223);
and U20792 (N_20792,N_16117,N_18389);
or U20793 (N_20793,N_16927,N_16930);
or U20794 (N_20794,N_17086,N_15711);
nand U20795 (N_20795,N_18195,N_19774);
xor U20796 (N_20796,N_15727,N_16012);
and U20797 (N_20797,N_17176,N_19919);
nor U20798 (N_20798,N_18201,N_15673);
and U20799 (N_20799,N_16390,N_17384);
and U20800 (N_20800,N_17636,N_18533);
nand U20801 (N_20801,N_19174,N_18137);
nand U20802 (N_20802,N_18448,N_17205);
and U20803 (N_20803,N_17964,N_18291);
nand U20804 (N_20804,N_16323,N_18144);
and U20805 (N_20805,N_18835,N_16013);
nand U20806 (N_20806,N_18355,N_19234);
xor U20807 (N_20807,N_19616,N_19655);
or U20808 (N_20808,N_16778,N_18122);
xnor U20809 (N_20809,N_15279,N_19121);
nand U20810 (N_20810,N_19627,N_15740);
nor U20811 (N_20811,N_15937,N_18628);
nand U20812 (N_20812,N_18004,N_17599);
xnor U20813 (N_20813,N_16500,N_18268);
xor U20814 (N_20814,N_17731,N_18530);
nand U20815 (N_20815,N_15638,N_17975);
nor U20816 (N_20816,N_16333,N_15135);
or U20817 (N_20817,N_15592,N_18729);
xor U20818 (N_20818,N_16030,N_19517);
or U20819 (N_20819,N_17882,N_16319);
xor U20820 (N_20820,N_19967,N_17199);
and U20821 (N_20821,N_16182,N_18612);
xnor U20822 (N_20822,N_17108,N_17483);
xor U20823 (N_20823,N_17999,N_17794);
nand U20824 (N_20824,N_16283,N_16632);
and U20825 (N_20825,N_15379,N_18608);
nor U20826 (N_20826,N_16100,N_19511);
and U20827 (N_20827,N_19904,N_15323);
and U20828 (N_20828,N_15192,N_17573);
xnor U20829 (N_20829,N_15528,N_18721);
or U20830 (N_20830,N_19576,N_17548);
or U20831 (N_20831,N_16653,N_18322);
xor U20832 (N_20832,N_19757,N_15919);
or U20833 (N_20833,N_15232,N_18417);
nand U20834 (N_20834,N_15207,N_15364);
xor U20835 (N_20835,N_15060,N_18891);
nor U20836 (N_20836,N_18274,N_19243);
or U20837 (N_20837,N_19803,N_19520);
xor U20838 (N_20838,N_18715,N_19335);
and U20839 (N_20839,N_18003,N_19363);
nor U20840 (N_20840,N_17806,N_15943);
or U20841 (N_20841,N_16105,N_18615);
or U20842 (N_20842,N_15959,N_15512);
or U20843 (N_20843,N_16291,N_17704);
nor U20844 (N_20844,N_19696,N_16552);
nor U20845 (N_20845,N_15455,N_17858);
nand U20846 (N_20846,N_15822,N_18214);
or U20847 (N_20847,N_17049,N_19009);
and U20848 (N_20848,N_17511,N_16977);
xor U20849 (N_20849,N_16891,N_15322);
nand U20850 (N_20850,N_18947,N_15272);
nand U20851 (N_20851,N_18983,N_17187);
and U20852 (N_20852,N_15030,N_15110);
nand U20853 (N_20853,N_17457,N_17000);
or U20854 (N_20854,N_18762,N_19132);
nand U20855 (N_20855,N_15228,N_16079);
nor U20856 (N_20856,N_18645,N_17719);
xnor U20857 (N_20857,N_15161,N_17947);
xnor U20858 (N_20858,N_19886,N_19845);
nand U20859 (N_20859,N_19822,N_16193);
xor U20860 (N_20860,N_18472,N_19734);
xnor U20861 (N_20861,N_17379,N_15565);
nand U20862 (N_20862,N_18358,N_15267);
or U20863 (N_20863,N_17621,N_18040);
or U20864 (N_20864,N_15215,N_17565);
nor U20865 (N_20865,N_15576,N_15221);
xor U20866 (N_20866,N_15481,N_17439);
nand U20867 (N_20867,N_17578,N_17637);
nand U20868 (N_20868,N_18709,N_17848);
nand U20869 (N_20869,N_19828,N_15665);
nor U20870 (N_20870,N_17083,N_19431);
nor U20871 (N_20871,N_17385,N_18344);
nor U20872 (N_20872,N_19927,N_17600);
or U20873 (N_20873,N_19360,N_15302);
nand U20874 (N_20874,N_15648,N_15921);
nand U20875 (N_20875,N_16986,N_16726);
nand U20876 (N_20876,N_15805,N_15773);
and U20877 (N_20877,N_18025,N_18089);
xnor U20878 (N_20878,N_19706,N_18115);
and U20879 (N_20879,N_16101,N_15336);
and U20880 (N_20880,N_19874,N_16015);
and U20881 (N_20881,N_17900,N_15702);
or U20882 (N_20882,N_18603,N_17813);
xnor U20883 (N_20883,N_16654,N_18818);
nand U20884 (N_20884,N_19055,N_19697);
nor U20885 (N_20885,N_16365,N_18330);
nand U20886 (N_20886,N_16644,N_19180);
and U20887 (N_20887,N_16507,N_18316);
nor U20888 (N_20888,N_16906,N_15452);
nor U20889 (N_20889,N_15694,N_17896);
nor U20890 (N_20890,N_18090,N_16848);
nor U20891 (N_20891,N_16307,N_19658);
or U20892 (N_20892,N_15686,N_15996);
or U20893 (N_20893,N_15143,N_16655);
or U20894 (N_20894,N_15383,N_16825);
or U20895 (N_20895,N_18733,N_16052);
nor U20896 (N_20896,N_16085,N_17503);
nor U20897 (N_20897,N_16935,N_15277);
nor U20898 (N_20898,N_17656,N_17761);
or U20899 (N_20899,N_19288,N_17362);
or U20900 (N_20900,N_16142,N_17886);
nor U20901 (N_20901,N_15985,N_16984);
or U20902 (N_20902,N_15464,N_17962);
nor U20903 (N_20903,N_17303,N_16462);
nor U20904 (N_20904,N_19795,N_16566);
nand U20905 (N_20905,N_17582,N_15369);
nand U20906 (N_20906,N_15445,N_17050);
nor U20907 (N_20907,N_15142,N_15790);
nand U20908 (N_20908,N_18488,N_15891);
and U20909 (N_20909,N_18669,N_19278);
and U20910 (N_20910,N_17735,N_19319);
nand U20911 (N_20911,N_15666,N_16133);
or U20912 (N_20912,N_18652,N_16233);
or U20913 (N_20913,N_15238,N_19952);
nand U20914 (N_20914,N_18810,N_19209);
or U20915 (N_20915,N_15210,N_16525);
nand U20916 (N_20916,N_16327,N_18329);
nor U20917 (N_20917,N_17103,N_19950);
xnor U20918 (N_20918,N_19454,N_19889);
nand U20919 (N_20919,N_15938,N_15641);
and U20920 (N_20920,N_18649,N_16743);
nor U20921 (N_20921,N_17745,N_19760);
nor U20922 (N_20922,N_19966,N_17681);
nor U20923 (N_20923,N_18492,N_18871);
xor U20924 (N_20924,N_17243,N_17692);
nand U20925 (N_20925,N_19839,N_19825);
nor U20926 (N_20926,N_17603,N_19392);
nand U20927 (N_20927,N_15840,N_15892);
xor U20928 (N_20928,N_19200,N_17296);
and U20929 (N_20929,N_17831,N_18093);
nor U20930 (N_20930,N_18128,N_16508);
and U20931 (N_20931,N_19534,N_17096);
nand U20932 (N_20932,N_16428,N_17845);
and U20933 (N_20933,N_19294,N_19315);
nand U20934 (N_20934,N_17420,N_17613);
xor U20935 (N_20935,N_18348,N_19638);
nor U20936 (N_20936,N_15932,N_19531);
nor U20937 (N_20937,N_18377,N_15331);
nor U20938 (N_20938,N_19797,N_15332);
and U20939 (N_20939,N_16330,N_18186);
or U20940 (N_20940,N_17700,N_17867);
and U20941 (N_20941,N_16073,N_19139);
nor U20942 (N_20942,N_15233,N_15354);
nand U20943 (N_20943,N_19202,N_17650);
or U20944 (N_20944,N_16592,N_15556);
xnor U20945 (N_20945,N_16708,N_17089);
nor U20946 (N_20946,N_15716,N_19790);
xnor U20947 (N_20947,N_16496,N_18018);
and U20948 (N_20948,N_15671,N_15426);
xor U20949 (N_20949,N_15991,N_17909);
nor U20950 (N_20950,N_16431,N_15837);
nand U20951 (N_20951,N_18565,N_16934);
nand U20952 (N_20952,N_19789,N_16367);
xnor U20953 (N_20953,N_17961,N_15196);
xnor U20954 (N_20954,N_15078,N_16217);
xor U20955 (N_20955,N_15970,N_15309);
nand U20956 (N_20956,N_15783,N_18811);
or U20957 (N_20957,N_17972,N_16892);
nor U20958 (N_20958,N_18471,N_19073);
xor U20959 (N_20959,N_18399,N_19293);
or U20960 (N_20960,N_19522,N_17005);
or U20961 (N_20961,N_17907,N_18809);
or U20962 (N_20962,N_17705,N_15578);
xnor U20963 (N_20963,N_18667,N_15341);
or U20964 (N_20964,N_19695,N_15104);
and U20965 (N_20965,N_15944,N_19435);
and U20966 (N_20966,N_18060,N_16306);
nand U20967 (N_20967,N_18066,N_18356);
or U20968 (N_20968,N_19408,N_19078);
or U20969 (N_20969,N_17504,N_17159);
xnor U20970 (N_20970,N_15026,N_18375);
nor U20971 (N_20971,N_16222,N_15911);
xor U20972 (N_20972,N_16486,N_17870);
and U20973 (N_20973,N_19339,N_18296);
nand U20974 (N_20974,N_15514,N_17798);
xnor U20975 (N_20975,N_16408,N_16873);
xnor U20976 (N_20976,N_16024,N_15067);
nand U20977 (N_20977,N_17340,N_15235);
nand U20978 (N_20978,N_17203,N_17321);
or U20979 (N_20979,N_17098,N_17226);
nand U20980 (N_20980,N_18759,N_18787);
or U20981 (N_20981,N_17757,N_19978);
or U20982 (N_20982,N_17370,N_15152);
and U20983 (N_20983,N_19266,N_15411);
xnor U20984 (N_20984,N_19111,N_16588);
or U20985 (N_20985,N_19878,N_15463);
and U20986 (N_20986,N_17627,N_19971);
and U20987 (N_20987,N_19579,N_17702);
nor U20988 (N_20988,N_18005,N_19472);
and U20989 (N_20989,N_17569,N_17371);
and U20990 (N_20990,N_15275,N_19210);
nand U20991 (N_20991,N_16704,N_19482);
xnor U20992 (N_20992,N_17929,N_19720);
or U20993 (N_20993,N_17279,N_16964);
and U20994 (N_20994,N_18086,N_17904);
nor U20995 (N_20995,N_19021,N_15972);
and U20996 (N_20996,N_15930,N_17926);
nor U20997 (N_20997,N_16752,N_18281);
xnor U20998 (N_20998,N_15338,N_19468);
xor U20999 (N_20999,N_16709,N_19391);
xnor U21000 (N_21000,N_17082,N_16409);
or U21001 (N_21001,N_19580,N_15087);
xor U21002 (N_21002,N_17060,N_19321);
or U21003 (N_21003,N_18582,N_17451);
nand U21004 (N_21004,N_18032,N_18057);
nand U21005 (N_21005,N_19811,N_15435);
or U21006 (N_21006,N_16014,N_19800);
or U21007 (N_21007,N_17758,N_16608);
nor U21008 (N_21008,N_15444,N_18930);
nand U21009 (N_21009,N_19082,N_15324);
or U21010 (N_21010,N_18289,N_16236);
or U21011 (N_21011,N_19224,N_19780);
nor U21012 (N_21012,N_15521,N_16191);
and U21013 (N_21013,N_19483,N_18450);
nor U21014 (N_21014,N_16095,N_19144);
or U21015 (N_21015,N_17493,N_18213);
or U21016 (N_21016,N_16975,N_17097);
nand U21017 (N_21017,N_19647,N_18896);
nor U21018 (N_21018,N_19006,N_18113);
nor U21019 (N_21019,N_18326,N_19880);
nor U21020 (N_21020,N_17188,N_15618);
or U21021 (N_21021,N_16593,N_18774);
nand U21022 (N_21022,N_18493,N_19296);
nand U21023 (N_21023,N_15306,N_18621);
xnor U21024 (N_21024,N_16598,N_19709);
nand U21025 (N_21025,N_17128,N_16763);
or U21026 (N_21026,N_19993,N_16821);
xnor U21027 (N_21027,N_19254,N_17807);
nor U21028 (N_21028,N_19038,N_19341);
and U21029 (N_21029,N_19700,N_19741);
nand U21030 (N_21030,N_17317,N_16607);
and U21031 (N_21031,N_18760,N_16169);
or U21032 (N_21032,N_16418,N_18352);
nor U21033 (N_21033,N_16197,N_16634);
nand U21034 (N_21034,N_17328,N_18462);
nor U21035 (N_21035,N_17037,N_19959);
or U21036 (N_21036,N_18880,N_15162);
and U21037 (N_21037,N_15899,N_17210);
nor U21038 (N_21038,N_16591,N_17911);
and U21039 (N_21039,N_17756,N_16226);
xnor U21040 (N_21040,N_16071,N_16231);
or U21041 (N_21041,N_17369,N_16348);
or U21042 (N_21042,N_19028,N_19861);
nand U21043 (N_21043,N_15415,N_19833);
and U21044 (N_21044,N_17519,N_17932);
xor U21045 (N_21045,N_17074,N_19541);
nor U21046 (N_21046,N_16815,N_17085);
nand U21047 (N_21047,N_18445,N_19449);
xor U21048 (N_21048,N_18254,N_19275);
nor U21049 (N_21049,N_17618,N_15926);
or U21050 (N_21050,N_18522,N_17712);
xor U21051 (N_21051,N_17482,N_16370);
nand U21052 (N_21052,N_19473,N_17633);
nor U21053 (N_21053,N_18065,N_15436);
or U21054 (N_21054,N_16582,N_17301);
and U21055 (N_21055,N_19340,N_18919);
and U21056 (N_21056,N_19479,N_18685);
xor U21057 (N_21057,N_17625,N_18912);
nand U21058 (N_21058,N_18568,N_15172);
xor U21059 (N_21059,N_15640,N_19941);
xnor U21060 (N_21060,N_16539,N_17275);
xnor U21061 (N_21061,N_19478,N_19495);
and U21062 (N_21062,N_15975,N_18402);
xnor U21063 (N_21063,N_18683,N_15351);
nand U21064 (N_21064,N_19560,N_16993);
xnor U21065 (N_21065,N_16022,N_18043);
nand U21066 (N_21066,N_15049,N_16363);
nor U21067 (N_21067,N_18393,N_17271);
or U21068 (N_21068,N_19726,N_16871);
nor U21069 (N_21069,N_18996,N_15094);
and U21070 (N_21070,N_17261,N_19514);
nor U21071 (N_21071,N_18817,N_16144);
xnor U21072 (N_21072,N_17076,N_19603);
xor U21073 (N_21073,N_15134,N_16164);
nand U21074 (N_21074,N_15958,N_16699);
nor U21075 (N_21075,N_16808,N_15737);
and U21076 (N_21076,N_18911,N_15631);
nand U21077 (N_21077,N_18295,N_17355);
and U21078 (N_21078,N_15159,N_19054);
and U21079 (N_21079,N_18875,N_16354);
and U21080 (N_21080,N_15802,N_17138);
nand U21081 (N_21081,N_16002,N_18192);
and U21082 (N_21082,N_19140,N_19913);
and U21083 (N_21083,N_17251,N_15873);
nor U21084 (N_21084,N_15475,N_16282);
and U21085 (N_21085,N_16730,N_19441);
xor U21086 (N_21086,N_15072,N_17979);
and U21087 (N_21087,N_15044,N_18190);
and U21088 (N_21088,N_15308,N_16945);
or U21089 (N_21089,N_15605,N_19328);
or U21090 (N_21090,N_18620,N_16092);
nor U21091 (N_21091,N_15881,N_19013);
nor U21092 (N_21092,N_16083,N_19867);
or U21093 (N_21093,N_17405,N_16969);
and U21094 (N_21094,N_16059,N_19929);
and U21095 (N_21095,N_18230,N_19349);
xor U21096 (N_21096,N_18909,N_15685);
nor U21097 (N_21097,N_16025,N_16246);
or U21098 (N_21098,N_17954,N_18944);
nor U21099 (N_21099,N_15453,N_15073);
nor U21100 (N_21100,N_18325,N_16387);
nor U21101 (N_21101,N_16805,N_18705);
xnor U21102 (N_21102,N_17513,N_18150);
nor U21103 (N_21103,N_19501,N_15812);
or U21104 (N_21104,N_17015,N_17392);
and U21105 (N_21105,N_17351,N_19099);
nor U21106 (N_21106,N_16836,N_18772);
nand U21107 (N_21107,N_19963,N_15682);
nor U21108 (N_21108,N_18838,N_19130);
nor U21109 (N_21109,N_17428,N_17295);
nor U21110 (N_21110,N_17105,N_19858);
xnor U21111 (N_21111,N_19138,N_15610);
or U21112 (N_21112,N_18815,N_16274);
or U21113 (N_21113,N_16075,N_16650);
and U21114 (N_21114,N_19487,N_17802);
or U21115 (N_21115,N_16057,N_18676);
xnor U21116 (N_21116,N_19547,N_15870);
or U21117 (N_21117,N_15733,N_16206);
nor U21118 (N_21118,N_15289,N_15533);
or U21119 (N_21119,N_15096,N_15595);
nor U21120 (N_21120,N_19944,N_15199);
nor U21121 (N_21121,N_18196,N_18339);
xnor U21122 (N_21122,N_16150,N_19333);
and U21123 (N_21123,N_16766,N_15297);
and U21124 (N_21124,N_16724,N_15187);
nand U21125 (N_21125,N_17843,N_15140);
xor U21126 (N_21126,N_19118,N_18509);
or U21127 (N_21127,N_19413,N_19755);
nor U21128 (N_21128,N_16545,N_16478);
nor U21129 (N_21129,N_19779,N_17736);
xnor U21130 (N_21130,N_16859,N_16449);
nand U21131 (N_21131,N_18130,N_17953);
nor U21132 (N_21132,N_18553,N_19424);
nand U21133 (N_21133,N_16374,N_18496);
and U21134 (N_21134,N_17965,N_16881);
and U21135 (N_21135,N_16189,N_16953);
nand U21136 (N_21136,N_16697,N_17619);
nand U21137 (N_21137,N_17133,N_18146);
or U21138 (N_21138,N_19049,N_18595);
or U21139 (N_21139,N_16235,N_18110);
nor U21140 (N_21140,N_19075,N_18644);
or U21141 (N_21141,N_19272,N_19896);
xnor U21142 (N_21142,N_17950,N_15437);
and U21143 (N_21143,N_19738,N_18037);
nor U21144 (N_21144,N_16876,N_17084);
xnor U21145 (N_21145,N_16249,N_17901);
nor U21146 (N_21146,N_16479,N_19195);
xor U21147 (N_21147,N_16921,N_18134);
nand U21148 (N_21148,N_15344,N_18889);
and U21149 (N_21149,N_18349,N_16212);
or U21150 (N_21150,N_17368,N_16475);
or U21151 (N_21151,N_18185,N_18512);
nand U21152 (N_21152,N_16268,N_18398);
nand U21153 (N_21153,N_15579,N_18390);
nor U21154 (N_21154,N_15265,N_16690);
nand U21155 (N_21155,N_15209,N_15530);
and U21156 (N_21156,N_16091,N_19083);
nand U21157 (N_21157,N_15625,N_15977);
and U21158 (N_21158,N_17206,N_18218);
xnor U21159 (N_21159,N_15420,N_15956);
or U21160 (N_21160,N_15019,N_16253);
nand U21161 (N_21161,N_15399,N_19844);
nand U21162 (N_21162,N_17033,N_19553);
and U21163 (N_21163,N_16735,N_17521);
xnor U21164 (N_21164,N_18978,N_19265);
xor U21165 (N_21165,N_16388,N_18557);
or U21166 (N_21166,N_16981,N_19306);
nand U21167 (N_21167,N_16497,N_17469);
xor U21168 (N_21168,N_19841,N_16207);
xnor U21169 (N_21169,N_16965,N_15021);
nor U21170 (N_21170,N_16943,N_18051);
nand U21171 (N_21171,N_18444,N_19970);
and U21172 (N_21172,N_19338,N_17099);
or U21173 (N_21173,N_18753,N_17647);
nor U21174 (N_21174,N_18437,N_16168);
nand U21175 (N_21175,N_19902,N_16227);
nand U21176 (N_21176,N_17928,N_16096);
nor U21177 (N_21177,N_18578,N_15754);
xnor U21178 (N_21178,N_17853,N_15818);
nor U21179 (N_21179,N_15128,N_15898);
nor U21180 (N_21180,N_17501,N_18039);
or U21181 (N_21181,N_16528,N_15281);
and U21182 (N_21182,N_15498,N_15054);
nor U21183 (N_21183,N_19532,N_15980);
xor U21184 (N_21184,N_15120,N_16060);
and U21185 (N_21185,N_16570,N_19399);
and U21186 (N_21186,N_15857,N_19996);
and U21187 (N_21187,N_15425,N_15076);
nor U21188 (N_21188,N_17078,N_15358);
or U21189 (N_21189,N_19492,N_19117);
nor U21190 (N_21190,N_16890,N_19050);
nor U21191 (N_21191,N_17246,N_18383);
nand U21192 (N_21192,N_16587,N_17793);
nor U21193 (N_21193,N_18668,N_17812);
nor U21194 (N_21194,N_19476,N_15007);
and U21195 (N_21195,N_19348,N_18353);
nand U21196 (N_21196,N_19213,N_16257);
or U21197 (N_21197,N_16173,N_17956);
xor U21198 (N_21198,N_17707,N_16070);
xor U21199 (N_21199,N_19352,N_16122);
nor U21200 (N_21200,N_15992,N_19915);
and U21201 (N_21201,N_17393,N_15724);
or U21202 (N_21202,N_18263,N_15088);
or U21203 (N_21203,N_15715,N_18412);
nand U21204 (N_21204,N_18943,N_16719);
nor U21205 (N_21205,N_19247,N_17738);
nor U21206 (N_21206,N_15468,N_15877);
nor U21207 (N_21207,N_15616,N_16039);
and U21208 (N_21208,N_15184,N_18054);
and U21209 (N_21209,N_19388,N_16463);
xor U21210 (N_21210,N_18846,N_18016);
nand U21211 (N_21211,N_17753,N_16398);
xnor U21212 (N_21212,N_16982,N_16813);
xnor U21213 (N_21213,N_18345,N_18662);
xor U21214 (N_21214,N_19783,N_18973);
xor U21215 (N_21215,N_18704,N_16167);
and U21216 (N_21216,N_15747,N_18052);
or U21217 (N_21217,N_19443,N_19942);
nor U21218 (N_21218,N_16335,N_15720);
xor U21219 (N_21219,N_17878,N_16027);
nand U21220 (N_21220,N_18499,N_15139);
or U21221 (N_21221,N_17859,N_17790);
nor U21222 (N_21222,N_15166,N_18575);
nand U21223 (N_21223,N_16464,N_19781);
nor U21224 (N_21224,N_16651,N_17386);
or U21225 (N_21225,N_15786,N_16851);
nor U21226 (N_21226,N_16162,N_18429);
and U21227 (N_21227,N_16896,N_15334);
nor U21228 (N_21228,N_18654,N_17143);
xor U21229 (N_21229,N_17322,N_16351);
nand U21230 (N_21230,N_16258,N_18133);
or U21231 (N_21231,N_18290,N_18719);
nor U21232 (N_21232,N_15889,N_17140);
xor U21233 (N_21233,N_19653,N_19292);
xor U21234 (N_21234,N_17249,N_18555);
nand U21235 (N_21235,N_19323,N_18507);
or U21236 (N_21236,N_17876,N_16738);
nor U21237 (N_21237,N_18484,N_17498);
nor U21238 (N_21238,N_18302,N_15125);
or U21239 (N_21239,N_17431,N_17309);
nand U21240 (N_21240,N_17288,N_18750);
nand U21241 (N_21241,N_18197,N_18964);
xnor U21242 (N_21242,N_15518,N_17447);
nand U21243 (N_21243,N_19273,N_16554);
nor U21244 (N_21244,N_17803,N_17156);
nand U21245 (N_21245,N_15253,N_17759);
or U21246 (N_21246,N_16956,N_16028);
or U21247 (N_21247,N_15225,N_18646);
nand U21248 (N_21248,N_19849,N_15337);
nand U21249 (N_21249,N_19330,N_19951);
nor U21250 (N_21250,N_15474,N_15950);
and U21251 (N_21251,N_17552,N_19632);
nor U21252 (N_21252,N_18698,N_15286);
and U21253 (N_21253,N_19031,N_18350);
xor U21254 (N_21254,N_18131,N_19621);
xor U21255 (N_21255,N_15257,N_17196);
or U21256 (N_21256,N_18591,N_16238);
nand U21257 (N_21257,N_16029,N_15884);
xor U21258 (N_21258,N_15064,N_16016);
or U21259 (N_21259,N_18929,N_19926);
and U21260 (N_21260,N_18632,N_17598);
and U21261 (N_21261,N_16356,N_15859);
nand U21262 (N_21262,N_17601,N_19156);
nor U21263 (N_21263,N_16502,N_16541);
xor U21264 (N_21264,N_18849,N_15008);
or U21265 (N_21265,N_15191,N_16991);
xor U21266 (N_21266,N_16795,N_19119);
xnor U21267 (N_21267,N_17489,N_17465);
nor U21268 (N_21268,N_17622,N_19529);
nand U21269 (N_21269,N_17913,N_18511);
nor U21270 (N_21270,N_17495,N_18042);
nand U21271 (N_21271,N_15915,N_16929);
xor U21272 (N_21272,N_17651,N_16035);
nor U21273 (N_21273,N_15077,N_18905);
xnor U21274 (N_21274,N_15432,N_17179);
nand U21275 (N_21275,N_15832,N_19452);
nor U21276 (N_21276,N_18307,N_19712);
xor U21277 (N_21277,N_18498,N_15206);
nand U21278 (N_21278,N_15245,N_15954);
nand U21279 (N_21279,N_15841,N_18898);
and U21280 (N_21280,N_15097,N_19361);
or U21281 (N_21281,N_18258,N_16143);
and U21282 (N_21282,N_16265,N_16435);
or U21283 (N_21283,N_16510,N_17276);
nand U21284 (N_21284,N_17374,N_15276);
and U21285 (N_21285,N_15449,N_15085);
and U21286 (N_21286,N_19477,N_16252);
or U21287 (N_21287,N_16639,N_19471);
or U21288 (N_21288,N_18744,N_18833);
or U21289 (N_21289,N_17157,N_15370);
nor U21290 (N_21290,N_19394,N_16887);
xnor U21291 (N_21291,N_15781,N_16121);
or U21292 (N_21292,N_17857,N_16846);
nor U21293 (N_21293,N_16751,N_15861);
or U21294 (N_21294,N_18463,N_17828);
and U21295 (N_21295,N_18921,N_18456);
and U21296 (N_21296,N_17526,N_16899);
or U21297 (N_21297,N_16534,N_19998);
nand U21298 (N_21298,N_18294,N_19465);
xnor U21299 (N_21299,N_16311,N_19450);
or U21300 (N_21300,N_18594,N_15722);
nor U21301 (N_21301,N_18246,N_17333);
xor U21302 (N_21302,N_17770,N_19248);
or U21303 (N_21303,N_18337,N_17977);
nand U21304 (N_21304,N_16854,N_15862);
nor U21305 (N_21305,N_17970,N_18761);
nor U21306 (N_21306,N_18798,N_15821);
nand U21307 (N_21307,N_15466,N_16897);
nor U21308 (N_21308,N_15782,N_16643);
nor U21309 (N_21309,N_16443,N_16713);
and U21310 (N_21310,N_18478,N_15016);
xor U21311 (N_21311,N_16777,N_15596);
and U21312 (N_21312,N_19235,N_19065);
or U21313 (N_21313,N_16145,N_18600);
nor U21314 (N_21314,N_15803,N_19723);
nor U21315 (N_21315,N_19609,N_18400);
and U21316 (N_21316,N_17715,N_18161);
or U21317 (N_21317,N_17661,N_18320);
nand U21318 (N_21318,N_19240,N_15183);
xor U21319 (N_21319,N_19525,N_16546);
xnor U21320 (N_21320,N_18660,N_19214);
nand U21321 (N_21321,N_18121,N_16089);
nand U21322 (N_21322,N_18629,N_17123);
or U21323 (N_21323,N_17971,N_19549);
nor U21324 (N_21324,N_16290,N_15202);
nor U21325 (N_21325,N_18908,N_19922);
and U21326 (N_21326,N_17869,N_15126);
nor U21327 (N_21327,N_18786,N_16453);
or U21328 (N_21328,N_17739,N_16728);
xnor U21329 (N_21329,N_18641,N_17866);
xnor U21330 (N_21330,N_17460,N_19994);
nand U21331 (N_21331,N_17440,N_18807);
and U21332 (N_21332,N_19972,N_17781);
nand U21333 (N_21333,N_17421,N_15190);
and U21334 (N_21334,N_15127,N_18624);
xnor U21335 (N_21335,N_18675,N_18031);
nor U21336 (N_21336,N_15197,N_18155);
nor U21337 (N_21337,N_18369,N_15393);
xor U21338 (N_21338,N_18248,N_17388);
nand U21339 (N_21339,N_19221,N_16901);
nor U21340 (N_21340,N_16733,N_17063);
nand U21341 (N_21341,N_19675,N_15619);
nor U21342 (N_21342,N_19670,N_16852);
xor U21343 (N_21343,N_19085,N_15544);
or U21344 (N_21344,N_19667,N_17124);
nand U21345 (N_21345,N_19320,N_17227);
nand U21346 (N_21346,N_15480,N_19497);
xnor U21347 (N_21347,N_18598,N_16560);
nor U21348 (N_21348,N_16384,N_17415);
and U21349 (N_21349,N_17347,N_19875);
nand U21350 (N_21350,N_17547,N_19916);
nor U21351 (N_21351,N_17418,N_17711);
or U21352 (N_21352,N_17543,N_18782);
nand U21353 (N_21353,N_19665,N_19241);
nand U21354 (N_21354,N_16099,N_19591);
xor U21355 (N_21355,N_17354,N_16471);
or U21356 (N_21356,N_15346,N_17075);
nor U21357 (N_21357,N_16616,N_19453);
and U21358 (N_21358,N_17434,N_16973);
nor U21359 (N_21359,N_18827,N_18092);
nand U21360 (N_21360,N_15814,N_15964);
and U21361 (N_21361,N_16337,N_19649);
or U21362 (N_21362,N_16155,N_15462);
xnor U21363 (N_21363,N_19469,N_16287);
nand U21364 (N_21364,N_18682,N_17400);
and U21365 (N_21365,N_18481,N_16216);
nor U21366 (N_21366,N_17545,N_15918);
or U21367 (N_21367,N_18893,N_18701);
nor U21368 (N_21368,N_16985,N_19542);
xor U21369 (N_21369,N_15778,N_18360);
or U21370 (N_21370,N_15405,N_16577);
nand U21371 (N_21371,N_18858,N_17446);
xor U21372 (N_21372,N_19744,N_15963);
nand U21373 (N_21373,N_19636,N_15806);
xnor U21374 (N_21374,N_18738,N_16898);
and U21375 (N_21375,N_17652,N_15038);
nand U21376 (N_21376,N_18199,N_18234);
or U21377 (N_21377,N_19661,N_18152);
or U21378 (N_21378,N_16314,N_17754);
xnor U21379 (N_21379,N_15676,N_17195);
or U21380 (N_21380,N_18236,N_18741);
xnor U21381 (N_21381,N_19090,N_17776);
nand U21382 (N_21382,N_18340,N_16196);
xnor U21383 (N_21383,N_16269,N_17877);
xor U21384 (N_21384,N_16456,N_17029);
xnor U21385 (N_21385,N_16369,N_16084);
and U21386 (N_21386,N_15390,N_15300);
or U21387 (N_21387,N_18950,N_18264);
nand U21388 (N_21388,N_19365,N_18665);
xor U21389 (N_21389,N_15075,N_17938);
nand U21390 (N_21390,N_19025,N_16331);
xnor U21391 (N_21391,N_16853,N_16297);
nor U21392 (N_21392,N_15391,N_15456);
nor U21393 (N_21393,N_17945,N_16244);
or U21394 (N_21394,N_15326,N_16494);
nand U21395 (N_21395,N_16521,N_15321);
and U21396 (N_21396,N_17051,N_19057);
or U21397 (N_21397,N_15114,N_18317);
nand U21398 (N_21398,N_19250,N_15880);
xor U21399 (N_21399,N_19681,N_19151);
or U21400 (N_21400,N_15845,N_19945);
and U21401 (N_21401,N_15149,N_17602);
and U21402 (N_21402,N_16894,N_17779);
or U21403 (N_21403,N_19619,N_17818);
and U21404 (N_21404,N_16441,N_16124);
nor U21405 (N_21405,N_17221,N_17285);
or U21406 (N_21406,N_16967,N_18554);
xnor U21407 (N_21407,N_19311,N_16066);
xnor U21408 (N_21408,N_16790,N_15700);
and U21409 (N_21409,N_18823,N_15705);
nand U21410 (N_21410,N_18205,N_16050);
nor U21411 (N_21411,N_15714,N_19377);
xor U21412 (N_21412,N_17747,N_15287);
or U21413 (N_21413,N_16937,N_16200);
and U21414 (N_21414,N_15398,N_17484);
nand U21415 (N_21415,N_15146,N_16702);
or U21416 (N_21416,N_17287,N_15792);
and U21417 (N_21417,N_18856,N_16325);
xnor U21418 (N_21418,N_19949,N_16638);
or U21419 (N_21419,N_15948,N_15342);
nor U21420 (N_21420,N_17113,N_16842);
and U21421 (N_21421,N_18879,N_17944);
and U21422 (N_21422,N_16138,N_19607);
or U21423 (N_21423,N_17575,N_17786);
and U21424 (N_21424,N_16649,N_17540);
nand U21425 (N_21425,N_16380,N_16706);
xnor U21426 (N_21426,N_15352,N_15601);
or U21427 (N_21427,N_18224,N_17576);
or U21428 (N_21428,N_18904,N_16017);
nor U21429 (N_21429,N_19624,N_18520);
nor U21430 (N_21430,N_19001,N_17762);
and U21431 (N_21431,N_17270,N_18293);
nand U21432 (N_21432,N_19227,N_16749);
and U21433 (N_21433,N_19559,N_15718);
nor U21434 (N_21434,N_18756,N_17267);
and U21435 (N_21435,N_15593,N_15795);
nor U21436 (N_21436,N_17816,N_18728);
and U21437 (N_21437,N_18969,N_18910);
or U21438 (N_21438,N_18604,N_16641);
nand U21439 (N_21439,N_17135,N_18227);
and U21440 (N_21440,N_19157,N_15039);
nor U21441 (N_21441,N_19276,N_18273);
and U21442 (N_21442,N_17035,N_17585);
or U21443 (N_21443,N_15368,N_16705);
nor U21444 (N_21444,N_15005,N_18648);
and U21445 (N_21445,N_18338,N_18657);
xnor U21446 (N_21446,N_16974,N_18547);
nand U21447 (N_21447,N_15796,N_19299);
or U21448 (N_21448,N_16353,N_18723);
and U21449 (N_21449,N_19125,N_18397);
or U21450 (N_21450,N_15895,N_16617);
and U21451 (N_21451,N_17228,N_17538);
xor U21452 (N_21452,N_16439,N_19637);
and U21453 (N_21453,N_19165,N_19147);
or U21454 (N_21454,N_19791,N_18145);
nor U21455 (N_21455,N_17491,N_15549);
or U21456 (N_21456,N_17940,N_17290);
nand U21457 (N_21457,N_19921,N_19163);
or U21458 (N_21458,N_19058,N_16535);
xor U21459 (N_21459,N_16933,N_16423);
and U21460 (N_21460,N_16195,N_18038);
nor U21461 (N_21461,N_16843,N_15150);
nand U21462 (N_21462,N_18371,N_17452);
xnor U21463 (N_21463,N_15371,N_19892);
xnor U21464 (N_21464,N_19650,N_17373);
nor U21465 (N_21465,N_16322,N_15000);
or U21466 (N_21466,N_18432,N_16505);
nor U21467 (N_21467,N_16519,N_18252);
nand U21468 (N_21468,N_17337,N_15433);
nor U21469 (N_21469,N_19694,N_19857);
or U21470 (N_21470,N_19702,N_15374);
xor U21471 (N_21471,N_15099,N_16672);
nand U21472 (N_21472,N_19122,N_16882);
xnor U21473 (N_21473,N_17743,N_15491);
nor U21474 (N_21474,N_15660,N_17435);
or U21475 (N_21475,N_15688,N_19003);
nand U21476 (N_21476,N_18427,N_18105);
or U21477 (N_21477,N_19063,N_16120);
or U21478 (N_21478,N_19387,N_19829);
nand U21479 (N_21479,N_18034,N_15330);
xnor U21480 (N_21480,N_19322,N_18001);
nor U21481 (N_21481,N_16557,N_18825);
nor U21482 (N_21482,N_18319,N_16289);
and U21483 (N_21483,N_16247,N_16399);
xor U21484 (N_21484,N_18170,N_16872);
or U21485 (N_21485,N_17031,N_19381);
nand U21486 (N_21486,N_16459,N_18866);
nor U21487 (N_21487,N_15600,N_18175);
nor U21488 (N_21488,N_19148,N_18590);
xor U21489 (N_21489,N_16310,N_17214);
and U21490 (N_21490,N_18107,N_16731);
xnor U21491 (N_21491,N_16698,N_15247);
nand U21492 (N_21492,N_15219,N_15649);
nand U21493 (N_21493,N_18165,N_16115);
nor U21494 (N_21494,N_17815,N_17315);
or U21495 (N_21495,N_18241,N_15606);
and U21496 (N_21496,N_16312,N_15109);
and U21497 (N_21497,N_19502,N_17984);
xnor U21498 (N_21498,N_18453,N_17348);
and U21499 (N_21499,N_16635,N_17225);
and U21500 (N_21500,N_17732,N_16046);
nand U21501 (N_21501,N_18370,N_18219);
xor U21502 (N_21502,N_18711,N_18631);
and U21503 (N_21503,N_16753,N_15271);
nand U21504 (N_21504,N_19604,N_15817);
and U21505 (N_21505,N_18826,N_18063);
nor U21506 (N_21506,N_17286,N_19194);
nor U21507 (N_21507,N_18583,N_15698);
xor U21508 (N_21508,N_15871,N_16154);
or U21509 (N_21509,N_19508,N_18475);
xor U21510 (N_21510,N_15622,N_17168);
or U21511 (N_21511,N_15335,N_18854);
nand U21512 (N_21512,N_18959,N_19984);
nand U21513 (N_21513,N_15916,N_18182);
or U21514 (N_21514,N_18688,N_17506);
or U21515 (N_21515,N_17101,N_17840);
or U21516 (N_21516,N_17860,N_17461);
or U21517 (N_21517,N_18229,N_17126);
or U21518 (N_21518,N_19530,N_16301);
xor U21519 (N_21519,N_16266,N_15529);
nor U21520 (N_21520,N_17414,N_16764);
and U21521 (N_21521,N_19129,N_15362);
or U21522 (N_21522,N_19625,N_17302);
or U21523 (N_21523,N_17294,N_16445);
nor U21524 (N_21524,N_18673,N_18588);
nand U21525 (N_21525,N_16447,N_17532);
nand U21526 (N_21526,N_16251,N_16850);
and U21527 (N_21527,N_16175,N_19018);
nand U21528 (N_21528,N_18138,N_15270);
nor U21529 (N_21529,N_17312,N_19331);
or U21530 (N_21530,N_18064,N_17924);
nor U21531 (N_21531,N_17219,N_17486);
and U21532 (N_21532,N_18757,N_19188);
nor U21533 (N_21533,N_17988,N_17772);
and U21534 (N_21534,N_15667,N_16578);
or U21535 (N_21535,N_19883,N_15564);
and U21536 (N_21536,N_18240,N_19109);
xor U21537 (N_21537,N_16248,N_18902);
nand U21538 (N_21538,N_17879,N_15627);
or U21539 (N_21539,N_16375,N_18627);
nand U21540 (N_21540,N_16998,N_15066);
xor U21541 (N_21541,N_15629,N_16395);
or U21542 (N_21542,N_15541,N_18957);
nand U21543 (N_21543,N_19080,N_18100);
or U21544 (N_21544,N_18116,N_19986);
or U21545 (N_21545,N_16078,N_19785);
xor U21546 (N_21546,N_19410,N_16954);
nor U21547 (N_21547,N_17535,N_18742);
nand U21548 (N_21548,N_17427,N_18724);
xnor U21549 (N_21549,N_16225,N_16342);
and U21550 (N_21550,N_15065,N_17255);
or U21551 (N_21551,N_17967,N_19552);
xor U21552 (N_21552,N_19490,N_18041);
xor U21553 (N_21553,N_17596,N_19982);
nand U21554 (N_21554,N_18907,N_17334);
xor U21555 (N_21555,N_15793,N_15652);
and U21556 (N_21556,N_18077,N_15476);
nand U21557 (N_21557,N_18056,N_19957);
xnor U21558 (N_21558,N_19239,N_17244);
or U21559 (N_21559,N_17441,N_15296);
and U21560 (N_21560,N_18984,N_16674);
nand U21561 (N_21561,N_19672,N_18308);
nor U21562 (N_21562,N_16250,N_15423);
or U21563 (N_21563,N_18443,N_15628);
xnor U21564 (N_21564,N_16466,N_19521);
and U21565 (N_21565,N_19765,N_17579);
and U21566 (N_21566,N_18381,N_19412);
or U21567 (N_21567,N_15626,N_18671);
and U21568 (N_21568,N_15116,N_17883);
nor U21569 (N_21569,N_16664,N_17800);
xnor U21570 (N_21570,N_15759,N_19870);
and U21571 (N_21571,N_15486,N_19992);
nand U21572 (N_21572,N_19402,N_17724);
xor U21573 (N_21573,N_19010,N_16049);
or U21574 (N_21574,N_18191,N_17462);
nand U21575 (N_21575,N_16088,N_19150);
xor U21576 (N_21576,N_15421,N_15885);
nand U21577 (N_21577,N_16862,N_17881);
nor U21578 (N_21578,N_17783,N_15785);
and U21579 (N_21579,N_18242,N_15966);
xnor U21580 (N_21580,N_16344,N_19284);
nand U21581 (N_21581,N_19300,N_19635);
nor U21582 (N_21582,N_17750,N_18906);
nor U21583 (N_21583,N_15082,N_18209);
nand U21584 (N_21584,N_19093,N_16411);
and U21585 (N_21585,N_16914,N_15838);
and U21586 (N_21586,N_16926,N_19070);
or U21587 (N_21587,N_15752,N_18058);
nand U21588 (N_21588,N_16807,N_17574);
or U21589 (N_21589,N_15105,N_19698);
xnor U21590 (N_21590,N_19516,N_18026);
nand U21591 (N_21591,N_19911,N_15846);
and U21592 (N_21592,N_17531,N_19160);
and U21593 (N_21593,N_16835,N_16922);
xor U21594 (N_21594,N_15416,N_18362);
or U21595 (N_21595,N_18262,N_15526);
xnor U21596 (N_21596,N_15010,N_15193);
and U21597 (N_21597,N_18059,N_16401);
xor U21598 (N_21598,N_17245,N_16109);
xnor U21599 (N_21599,N_19373,N_19895);
and U21600 (N_21600,N_19671,N_16912);
nand U21601 (N_21601,N_17326,N_18379);
or U21602 (N_21602,N_18661,N_16561);
or U21603 (N_21603,N_15550,N_16007);
or U21604 (N_21604,N_16113,N_19178);
or U21605 (N_21605,N_19127,N_16054);
xnor U21606 (N_21606,N_18792,N_17025);
and U21607 (N_21607,N_18257,N_15396);
or U21608 (N_21608,N_15118,N_17721);
nor U21609 (N_21609,N_18176,N_19499);
nor U21610 (N_21610,N_15360,N_15004);
and U21611 (N_21611,N_19396,N_18663);
or U21612 (N_21612,N_16371,N_18118);
nor U21613 (N_21613,N_18410,N_15372);
xor U21614 (N_21614,N_19572,N_19172);
and U21615 (N_21615,N_15735,N_17073);
or U21616 (N_21616,N_18099,N_15256);
or U21617 (N_21617,N_18872,N_17642);
or U21618 (N_21618,N_17407,N_17232);
xor U21619 (N_21619,N_18931,N_16458);
nand U21620 (N_21620,N_17081,N_17703);
xor U21621 (N_21621,N_16689,N_18010);
xnor U21622 (N_21622,N_17383,N_19282);
nand U21623 (N_21623,N_15496,N_19838);
nand U21624 (N_21624,N_16318,N_15141);
nand U21625 (N_21625,N_17141,N_18255);
xnor U21626 (N_21626,N_15343,N_17737);
or U21627 (N_21627,N_16574,N_15710);
or U21628 (N_21628,N_17153,N_15742);
nand U21629 (N_21629,N_17282,N_17204);
and U21630 (N_21630,N_18357,N_18097);
nor U21631 (N_21631,N_15154,N_17862);
nor U21632 (N_21632,N_16820,N_19934);
nand U21633 (N_21633,N_17172,N_19565);
and U21634 (N_21634,N_19953,N_19199);
or U21635 (N_21635,N_16723,N_16213);
xnor U21636 (N_21636,N_18036,N_18518);
nand U21637 (N_21637,N_15252,N_17036);
or U21638 (N_21638,N_16979,N_17710);
and U21639 (N_21639,N_17020,N_17617);
and U21640 (N_21640,N_16818,N_17955);
and U21641 (N_21641,N_17509,N_19817);
or U21642 (N_21642,N_16568,N_18870);
or U21643 (N_21643,N_17304,N_18556);
or U21644 (N_21644,N_18537,N_18745);
nor U21645 (N_21645,N_15262,N_17644);
nor U21646 (N_21646,N_17655,N_15807);
nor U21647 (N_21647,N_19848,N_16298);
or U21648 (N_21648,N_15080,N_16810);
nor U21649 (N_21649,N_17028,N_16693);
nor U21650 (N_21650,N_15218,N_18867);
or U21651 (N_21651,N_19379,N_19177);
nand U21652 (N_21652,N_18780,N_16586);
nor U21653 (N_21653,N_18876,N_16433);
and U21654 (N_21654,N_16711,N_18094);
and U21655 (N_21655,N_19539,N_17607);
nand U21656 (N_21656,N_19029,N_18850);
or U21657 (N_21657,N_19746,N_18666);
nor U21658 (N_21658,N_15523,N_18801);
and U21659 (N_21659,N_15268,N_17088);
xnor U21660 (N_21660,N_17771,N_16440);
nor U21661 (N_21661,N_18640,N_18327);
nand U21662 (N_21662,N_18727,N_16404);
and U21663 (N_21663,N_18775,N_19350);
nor U21664 (N_21664,N_19390,N_17890);
and U21665 (N_21665,N_17951,N_18962);
xor U21666 (N_21666,N_17558,N_16645);
or U21667 (N_21667,N_18232,N_15031);
nand U21668 (N_21668,N_15896,N_15438);
and U21669 (N_21669,N_18477,N_19589);
nand U21670 (N_21670,N_18634,N_17915);
nor U21671 (N_21671,N_17215,N_18842);
and U21672 (N_21672,N_16798,N_17969);
and U21673 (N_21673,N_16420,N_18083);
and U21674 (N_21674,N_18900,N_15417);
or U21675 (N_21675,N_15637,N_18532);
xor U21676 (N_21676,N_16530,N_16600);
nor U21677 (N_21677,N_17423,N_19267);
and U21678 (N_21678,N_18938,N_19954);
or U21679 (N_21679,N_17382,N_15515);
or U21680 (N_21680,N_15535,N_19618);
nand U21681 (N_21681,N_16594,N_16770);
and U21682 (N_21682,N_18606,N_19778);
nand U21683 (N_21683,N_17561,N_15211);
xor U21684 (N_21684,N_15906,N_15130);
xor U21685 (N_21685,N_18566,N_17554);
xnor U21686 (N_21686,N_17358,N_15282);
and U21687 (N_21687,N_15246,N_17167);
nor U21688 (N_21688,N_19938,N_15988);
or U21689 (N_21689,N_18049,N_17864);
nand U21690 (N_21690,N_17562,N_19027);
xor U21691 (N_21691,N_16199,N_17665);
nor U21692 (N_21692,N_19745,N_15888);
nand U21693 (N_21693,N_19894,N_16512);
nor U21694 (N_21694,N_18024,N_18593);
nand U21695 (N_21695,N_18581,N_18941);
nand U21696 (N_21696,N_15178,N_19301);
and U21697 (N_21697,N_18044,N_18636);
nand U21698 (N_21698,N_18109,N_19258);
nor U21699 (N_21699,N_17022,N_15046);
or U21700 (N_21700,N_17789,N_16895);
nor U21701 (N_21701,N_18956,N_15765);
and U21702 (N_21702,N_17163,N_18881);
nor U21703 (N_21703,N_15024,N_17090);
or U21704 (N_21704,N_17111,N_15635);
nand U21705 (N_21705,N_18225,N_19161);
and U21706 (N_21706,N_16181,N_15914);
nor U21707 (N_21707,N_17788,N_16961);
nand U21708 (N_21708,N_18035,N_17239);
nor U21709 (N_21709,N_15506,N_15566);
and U21710 (N_21710,N_18265,N_19382);
nor U21711 (N_21711,N_19162,N_18474);
nor U21712 (N_21712,N_17170,N_18989);
nor U21713 (N_21713,N_17229,N_18166);
nand U21714 (N_21714,N_16811,N_19326);
and U21715 (N_21715,N_17529,N_15929);
xor U21716 (N_21716,N_16828,N_17923);
and U21717 (N_21717,N_18677,N_15062);
nor U21718 (N_21718,N_15510,N_15643);
nand U21719 (N_21719,N_16093,N_18490);
and U21720 (N_21720,N_17404,N_18743);
nor U21721 (N_21721,N_15384,N_15375);
or U21722 (N_21722,N_18007,N_18359);
nor U21723 (N_21723,N_19688,N_18085);
or U21724 (N_21724,N_16822,N_18736);
nor U21725 (N_21725,N_19242,N_16847);
xnor U21726 (N_21726,N_16736,N_15492);
xnor U21727 (N_21727,N_18315,N_17672);
or U21728 (N_21728,N_18048,N_15381);
nor U21729 (N_21729,N_16352,N_19383);
nor U21730 (N_21730,N_15548,N_19061);
and U21731 (N_21731,N_19877,N_19776);
nor U21732 (N_21732,N_16064,N_19143);
and U21733 (N_21733,N_19961,N_19864);
or U21734 (N_21734,N_18642,N_16209);
or U21735 (N_21735,N_19819,N_19133);
xor U21736 (N_21736,N_18954,N_16161);
nand U21737 (N_21737,N_19494,N_19630);
xor U21738 (N_21738,N_16107,N_15424);
nand U21739 (N_21739,N_19997,N_17517);
and U21740 (N_21740,N_19856,N_17166);
and U21741 (N_21741,N_19115,N_15984);
xor U21742 (N_21742,N_19979,N_15770);
xnor U21743 (N_21743,N_18441,N_18216);
nand U21744 (N_21744,N_18843,N_18694);
xor U21745 (N_21745,N_19113,N_15316);
xnor U21746 (N_21746,N_15034,N_19184);
nor U21747 (N_21747,N_17458,N_16995);
nor U21748 (N_21748,N_16550,N_17142);
or U21749 (N_21749,N_16141,N_19669);
nor U21750 (N_21750,N_16556,N_17726);
xnor U21751 (N_21751,N_15864,N_18102);
and U21752 (N_21752,N_17949,N_17557);
and U21753 (N_21753,N_17466,N_19980);
nand U21754 (N_21754,N_16938,N_19879);
or U21755 (N_21755,N_17106,N_17079);
nand U21756 (N_21756,N_19973,N_16756);
or U21757 (N_21757,N_16746,N_16086);
and U21758 (N_21758,N_15389,N_17671);
and U21759 (N_21759,N_17834,N_18651);
xor U21760 (N_21760,N_18247,N_17614);
and U21761 (N_21761,N_19764,N_16522);
or U21762 (N_21762,N_19876,N_17202);
nand U21763 (N_21763,N_16134,N_18179);
xnor U21764 (N_21764,N_19081,N_18193);
nand U21765 (N_21765,N_19958,N_15448);
or U21766 (N_21766,N_16037,N_17268);
or U21767 (N_21767,N_16275,N_17632);
nand U21768 (N_21768,N_18368,N_19444);
or U21769 (N_21769,N_15244,N_19826);
nand U21770 (N_21770,N_17480,N_17589);
xnor U21771 (N_21771,N_17639,N_17292);
and U21772 (N_21772,N_17520,N_17148);
nor U21773 (N_21773,N_18256,N_19692);
nand U21774 (N_21774,N_19595,N_17605);
or U21775 (N_21775,N_19166,N_18403);
xor U21776 (N_21776,N_15809,N_17324);
nand U21777 (N_21777,N_15357,N_17238);
nand U21778 (N_21778,N_17978,N_18104);
nand U21779 (N_21779,N_18525,N_19211);
nor U21780 (N_21780,N_16569,N_15227);
xnor U21781 (N_21781,N_15511,N_19274);
or U21782 (N_21782,N_16615,N_18157);
and U21783 (N_21783,N_15112,N_16868);
and U21784 (N_21784,N_18405,N_18998);
nor U21785 (N_21785,N_18226,N_15695);
or U21786 (N_21786,N_19179,N_17584);
xor U21787 (N_21787,N_18699,N_15458);
nand U21788 (N_21788,N_15494,N_17549);
xor U21789 (N_21789,N_18771,N_15572);
nor U21790 (N_21790,N_18607,N_19735);
xor U21791 (N_21791,N_18829,N_15355);
xor U21792 (N_21792,N_15617,N_18548);
and U21793 (N_21793,N_18159,N_16532);
nand U21794 (N_21794,N_16739,N_19792);
xnor U21795 (N_21795,N_16108,N_19570);
xnor U21796 (N_21796,N_17685,N_15653);
or U21797 (N_21797,N_16590,N_17847);
xnor U21798 (N_21798,N_15804,N_19398);
and U21799 (N_21799,N_16515,N_16366);
xnor U21800 (N_21800,N_18618,N_16364);
or U21801 (N_21801,N_19332,N_17472);
or U21802 (N_21802,N_15493,N_16184);
or U21803 (N_21803,N_17001,N_18965);
xnor U21804 (N_21804,N_16004,N_19012);
and U21805 (N_21805,N_16949,N_18497);
or U21806 (N_21806,N_19930,N_18177);
nand U21807 (N_21807,N_15242,N_19271);
or U21808 (N_21808,N_16112,N_16750);
or U21809 (N_21809,N_17683,N_16710);
nand U21810 (N_21810,N_15147,N_19102);
xnor U21811 (N_21811,N_18002,N_15774);
xnor U21812 (N_21812,N_18777,N_16234);
and U21813 (N_21813,N_19956,N_19042);
and U21814 (N_21814,N_15633,N_17555);
and U21815 (N_21815,N_17641,N_17297);
xor U21816 (N_21816,N_17009,N_16745);
nand U21817 (N_21817,N_17889,N_18447);
nand U21818 (N_21818,N_19690,N_17241);
or U21819 (N_21819,N_19563,N_17678);
xnor U21820 (N_21820,N_19568,N_19203);
xnor U21821 (N_21821,N_16540,N_18436);
or U21822 (N_21822,N_17310,N_18986);
nor U21823 (N_21823,N_17528,N_18836);
or U21824 (N_21824,N_15941,N_17476);
or U21825 (N_21825,N_15797,N_16742);
or U21826 (N_21826,N_17846,N_16955);
xor U21827 (N_21827,N_18347,N_18238);
xor U21828 (N_21828,N_15965,N_18149);
and U21829 (N_21829,N_17820,N_15875);
and U21830 (N_21830,N_16242,N_19586);
nand U21831 (N_21831,N_17184,N_15487);
nand U21832 (N_21832,N_16564,N_19237);
nand U21833 (N_21833,N_15568,N_16513);
xor U21834 (N_21834,N_16389,N_15961);
and U21835 (N_21835,N_17216,N_16094);
nand U21836 (N_21836,N_17695,N_19748);
or U21837 (N_21837,N_18391,N_17468);
xnor U21838 (N_21838,N_18567,N_17344);
nand U21839 (N_21839,N_19960,N_15469);
or U21840 (N_21840,N_19342,N_16338);
xor U21841 (N_21841,N_19259,N_18415);
nand U21842 (N_21842,N_18438,N_17833);
nand U21843 (N_21843,N_19044,N_19901);
xor U21844 (N_21844,N_19577,N_17426);
or U21845 (N_21845,N_15500,N_17307);
nand U21846 (N_21846,N_17746,N_16680);
nand U21847 (N_21847,N_19918,N_18940);
nand U21848 (N_21848,N_17380,N_17935);
or U21849 (N_21849,N_19475,N_18074);
and U21850 (N_21850,N_15482,N_19418);
and U21851 (N_21851,N_18913,N_19230);
nand U21852 (N_21852,N_15922,N_19324);
nor U21853 (N_21853,N_15036,N_17459);
and U21854 (N_21854,N_16879,N_19827);
and U21855 (N_21855,N_15699,N_15185);
nor U21856 (N_21856,N_18328,N_19223);
xnor U21857 (N_21857,N_15939,N_15497);
xnor U21858 (N_21858,N_16359,N_17593);
or U21859 (N_21859,N_16178,N_16208);
xnor U21860 (N_21860,N_15987,N_15359);
and U21861 (N_21861,N_17263,N_19620);
nor U21862 (N_21862,N_18544,N_17819);
or U21863 (N_21863,N_15729,N_17888);
or U21864 (N_21864,N_19108,N_18164);
and U21865 (N_21865,N_19463,N_15327);
or U21866 (N_21866,N_17306,N_19900);
and U21867 (N_21867,N_19357,N_15696);
and U21868 (N_21868,N_16336,N_19047);
or U21869 (N_21869,N_17408,N_16304);
nand U21870 (N_21870,N_17198,N_16831);
xnor U21871 (N_21871,N_18476,N_15136);
nand U21872 (N_21872,N_17107,N_19364);
or U21873 (N_21873,N_15089,N_19089);
or U21874 (N_21874,N_18751,N_18577);
xor U21875 (N_21875,N_18147,N_15769);
nand U21876 (N_21876,N_15831,N_16572);
nand U21877 (N_21877,N_16111,N_19677);
or U21878 (N_21878,N_19329,N_19656);
or U21879 (N_21879,N_17464,N_17808);
nor U21880 (N_21880,N_16006,N_17280);
xnor U21881 (N_21881,N_15414,N_19769);
xnor U21882 (N_21882,N_15339,N_15033);
nor U21883 (N_21883,N_16061,N_18409);
nor U21884 (N_21884,N_17629,N_18270);
xor U21885 (N_21885,N_15901,N_17863);
xor U21886 (N_21886,N_16477,N_18975);
or U21887 (N_21887,N_16596,N_17740);
nand U21888 (N_21888,N_18955,N_19989);
and U21889 (N_21889,N_15577,N_16171);
nor U21890 (N_21890,N_17580,N_19155);
nor U21891 (N_21891,N_18194,N_18204);
xnor U21892 (N_21892,N_15942,N_17922);
nand U21893 (N_21893,N_16340,N_19759);
and U21894 (N_21894,N_18976,N_17825);
and U21895 (N_21895,N_19091,N_15158);
xnor U21896 (N_21896,N_16110,N_19663);
nand U21897 (N_21897,N_17052,N_15427);
and U21898 (N_21898,N_15069,N_17152);
xnor U21899 (N_21899,N_19749,N_16948);
or U21900 (N_21900,N_16320,N_19159);
or U21901 (N_21901,N_16725,N_16928);
or U21902 (N_21902,N_16768,N_18449);
xor U21903 (N_21903,N_16783,N_19575);
xor U21904 (N_21904,N_18469,N_17325);
nand U21905 (N_21905,N_15418,N_17918);
nand U21906 (N_21906,N_15188,N_15910);
nand U21907 (N_21907,N_19215,N_16747);
or U21908 (N_21908,N_17604,N_18454);
nand U21909 (N_21909,N_17787,N_18569);
or U21910 (N_21910,N_16192,N_19374);
and U21911 (N_21911,N_15255,N_16903);
nor U21912 (N_21912,N_19110,N_17973);
or U21913 (N_21913,N_16321,N_17946);
xor U21914 (N_21914,N_16355,N_18948);
and U21915 (N_21915,N_17438,N_15580);
xnor U21916 (N_21916,N_18156,N_19269);
and U21917 (N_21917,N_17314,N_19909);
nor U21918 (N_21918,N_16339,N_16626);
or U21919 (N_21919,N_18168,N_17987);
nor U21920 (N_21920,N_16624,N_18888);
nand U21921 (N_21921,N_16480,N_15009);
xnor U21922 (N_21922,N_17667,N_16628);
nor U21923 (N_21923,N_16378,N_17708);
or U21924 (N_21924,N_19170,N_19711);
or U21925 (N_21925,N_16700,N_19167);
nor U21926 (N_21926,N_19369,N_19052);
xnor U21927 (N_21927,N_16636,N_19924);
nand U21928 (N_21928,N_15280,N_18331);
nor U21929 (N_21929,N_18261,N_16481);
and U21930 (N_21930,N_18703,N_19277);
and U21931 (N_21931,N_15223,N_19430);
nor U21932 (N_21932,N_16788,N_19417);
nor U21933 (N_21933,N_15878,N_19347);
nand U21934 (N_21934,N_15459,N_16988);
or U21935 (N_21935,N_18935,N_15086);
or U21936 (N_21936,N_18625,N_15050);
nor U21937 (N_21937,N_15121,N_18993);
nor U21938 (N_21938,N_19991,N_15583);
nand U21939 (N_21939,N_18689,N_18886);
nand U21940 (N_21940,N_18148,N_16243);
nand U21941 (N_21941,N_17792,N_15483);
nand U21942 (N_21942,N_19415,N_19022);
or U21943 (N_21943,N_16316,N_18920);
or U21944 (N_21944,N_15613,N_16772);
or U21945 (N_21945,N_16493,N_16809);
xor U21946 (N_21946,N_18251,N_18901);
xnor U21947 (N_21947,N_16877,N_17416);
nand U21948 (N_21948,N_18696,N_16720);
nor U21949 (N_21949,N_15743,N_18079);
xnor U21950 (N_21950,N_16833,N_18596);
or U21951 (N_21951,N_16665,N_16537);
and U21952 (N_21952,N_17026,N_17826);
xor U21953 (N_21953,N_18979,N_17698);
or U21954 (N_21954,N_16003,N_17134);
nand U21955 (N_21955,N_16183,N_19733);
and U21956 (N_21956,N_19458,N_19606);
nor U21957 (N_21957,N_19588,N_16308);
and U21958 (N_21958,N_19842,N_19245);
and U21959 (N_21959,N_15180,N_15811);
or U21960 (N_21960,N_19739,N_15298);
or U21961 (N_21961,N_19217,N_16185);
nor U21962 (N_21962,N_15632,N_19855);
xnor U21963 (N_21963,N_15611,N_15788);
xor U21964 (N_21964,N_16946,N_16285);
nor U21965 (N_21965,N_18174,N_18614);
nand U21966 (N_21966,N_16646,N_18708);
or U21967 (N_21967,N_15620,N_17577);
nor U21968 (N_21968,N_17663,N_15663);
nor U21969 (N_21969,N_19718,N_18464);
nand U21970 (N_21970,N_15495,N_19564);
nand U21971 (N_21971,N_17345,N_17744);
and U21972 (N_21972,N_18208,N_15839);
or U21973 (N_21973,N_15609,N_17976);
or U21974 (N_21974,N_19890,N_16136);
nand U21975 (N_21975,N_15955,N_15194);
nand U21976 (N_21976,N_19304,N_16427);
nor U21977 (N_21977,N_19969,N_17785);
or U21978 (N_21978,N_19939,N_16137);
nand U21979 (N_21979,N_19041,N_19297);
nand U21980 (N_21980,N_15201,N_16741);
nor U21981 (N_21981,N_16755,N_19546);
and U21982 (N_21982,N_16180,N_16417);
nand U21983 (N_21983,N_19020,N_15947);
and U21984 (N_21984,N_18361,N_16874);
and U21985 (N_21985,N_19015,N_18545);
nor U21986 (N_21986,N_19573,N_17004);
xor U21987 (N_21987,N_19279,N_17906);
nor U21988 (N_21988,N_15678,N_15868);
and U21989 (N_21989,N_19077,N_15589);
nor U21990 (N_21990,N_19594,N_17634);
and U21991 (N_21991,N_16264,N_19420);
xnor U21992 (N_21992,N_19309,N_17146);
and U21993 (N_21993,N_18231,N_16804);
and U21994 (N_21994,N_15940,N_16857);
or U21995 (N_21995,N_16997,N_19574);
nand U21996 (N_21996,N_18114,N_16036);
nand U21997 (N_21997,N_15534,N_15525);
nand U21998 (N_21998,N_17957,N_19256);
nor U21999 (N_21999,N_19406,N_17893);
nand U22000 (N_22000,N_16303,N_15546);
or U22001 (N_22001,N_18422,N_17104);
xnor U22002 (N_22002,N_16446,N_16055);
and U22003 (N_22003,N_16293,N_17479);
nand U22004 (N_22004,N_19308,N_16909);
or U22005 (N_22005,N_17008,N_17454);
nand U22006 (N_22006,N_18401,N_19766);
nand U22007 (N_22007,N_17127,N_17429);
xnor U22008 (N_22008,N_19611,N_19850);
or U22009 (N_22009,N_16683,N_17095);
and U22010 (N_22010,N_16989,N_18579);
or U22011 (N_22011,N_19908,N_15960);
xnor U22012 (N_22012,N_18552,N_16416);
or U22013 (N_22013,N_19509,N_17366);
xor U22014 (N_22014,N_16413,N_18538);
or U22015 (N_22015,N_16642,N_19149);
nand U22016 (N_22016,N_18457,N_17948);
nand U22017 (N_22017,N_18160,N_18882);
and U22018 (N_22018,N_19228,N_17659);
xor U22019 (N_22019,N_15090,N_19933);
nor U22020 (N_22020,N_19678,N_19051);
and U22021 (N_22021,N_15508,N_18597);
or U22022 (N_22022,N_17689,N_17566);
nor U22023 (N_22023,N_15657,N_17145);
or U22024 (N_22024,N_17773,N_17055);
nor U22025 (N_22025,N_17091,N_17339);
nand U22026 (N_22026,N_19145,N_16908);
nor U22027 (N_22027,N_17272,N_16451);
nor U22028 (N_22028,N_18609,N_17064);
nand U22029 (N_22029,N_18333,N_15924);
xnor U22030 (N_22030,N_17664,N_19190);
nand U22031 (N_22031,N_17151,N_17990);
xor U22032 (N_22032,N_19528,N_19440);
or U22033 (N_22033,N_18819,N_17230);
nor U22034 (N_22034,N_18253,N_17986);
nor U22035 (N_22035,N_15226,N_17764);
nor U22036 (N_22036,N_19557,N_15501);
and U22037 (N_22037,N_19498,N_18863);
xor U22038 (N_22038,N_19036,N_17234);
nand U22039 (N_22039,N_18917,N_15284);
or U22040 (N_22040,N_19445,N_18799);
nand U22041 (N_22041,N_16722,N_18529);
nand U22042 (N_22042,N_18461,N_19104);
nand U22043 (N_22043,N_15800,N_19366);
nor U22044 (N_22044,N_17865,N_15642);
or U22045 (N_22045,N_18283,N_17487);
nor U22046 (N_22046,N_18623,N_16551);
xor U22047 (N_22047,N_19500,N_15312);
nor U22048 (N_22048,N_18914,N_19428);
nand U22049 (N_22049,N_17912,N_16844);
or U22050 (N_22050,N_18243,N_16839);
nor U22051 (N_22051,N_18151,N_19014);
nand U22052 (N_22052,N_16939,N_19393);
nor U22053 (N_22053,N_17611,N_16239);
and U22054 (N_22054,N_17982,N_15887);
nand U22055 (N_22055,N_15874,N_17722);
nand U22056 (N_22056,N_19968,N_19743);
and U22057 (N_22057,N_15499,N_17183);
nor U22058 (N_22058,N_18029,N_16667);
xnor U22059 (N_22059,N_16791,N_15668);
and U22060 (N_22060,N_16019,N_16148);
nand U22061 (N_22061,N_17335,N_18589);
and U22062 (N_22062,N_19898,N_16172);
nor U22063 (N_22063,N_19676,N_19355);
or U22064 (N_22064,N_17917,N_17937);
nor U22065 (N_22065,N_18479,N_18465);
xor U22066 (N_22066,N_18081,N_18754);
nand U22067 (N_22067,N_18816,N_15442);
and U22068 (N_22068,N_17778,N_16473);
nand U22069 (N_22069,N_17158,N_16734);
nand U22070 (N_22070,N_16911,N_19823);
xnor U22071 (N_22071,N_16044,N_19888);
nand U22072 (N_22072,N_18918,N_16457);
nor U22073 (N_22073,N_17727,N_15815);
nor U22074 (N_22074,N_18508,N_15697);
and U22075 (N_22075,N_18142,N_15461);
xor U22076 (N_22076,N_18023,N_18752);
nor U22077 (N_22077,N_17936,N_19543);
xnor U22078 (N_22078,N_17749,N_19943);
nor U22079 (N_22079,N_15373,N_15173);
nand U22080 (N_22080,N_17640,N_19263);
nand U22081 (N_22081,N_18184,N_18763);
and U22082 (N_22082,N_15431,N_16158);
xor U22083 (N_22083,N_19040,N_18030);
nand U22084 (N_22084,N_15621,N_19987);
and U22085 (N_22085,N_15439,N_16579);
nor U22086 (N_22086,N_19353,N_16001);
or U22087 (N_22087,N_16179,N_17809);
or U22088 (N_22088,N_15254,N_15923);
nor U22089 (N_22089,N_18706,N_18725);
xnor U22090 (N_22090,N_15744,N_15098);
nor U22091 (N_22091,N_16386,N_16051);
and U22092 (N_22092,N_16925,N_16224);
and U22093 (N_22093,N_15400,N_16715);
xor U22094 (N_22094,N_19226,N_15607);
or U22095 (N_22095,N_17908,N_19715);
and U22096 (N_22096,N_15808,N_15986);
nor U22097 (N_22097,N_15634,N_16156);
xnor U22098 (N_22098,N_15317,N_18341);
and U22099 (N_22099,N_16686,N_18937);
xor U22100 (N_22100,N_18343,N_15756);
or U22101 (N_22101,N_19752,N_15799);
nor U22102 (N_22102,N_16062,N_18684);
xor U22103 (N_22103,N_15739,N_17512);
and U22104 (N_22104,N_19600,N_16072);
xor U22105 (N_22105,N_17524,N_16599);
and U22106 (N_22106,N_18141,N_19201);
nor U22107 (N_22107,N_19750,N_19596);
xnor U22108 (N_22108,N_18306,N_16913);
and U22109 (N_22109,N_18424,N_19183);
xor U22110 (N_22110,N_17455,N_18304);
nor U22111 (N_22111,N_15681,N_18779);
nor U22112 (N_22112,N_15059,N_15777);
or U22113 (N_22113,N_16245,N_19818);
and U22114 (N_22114,N_15430,N_19556);
nor U22115 (N_22115,N_17254,N_17968);
nand U22116 (N_22116,N_16135,N_16186);
or U22117 (N_22117,N_17381,N_16229);
and U22118 (N_22118,N_17734,N_15844);
nor U22119 (N_22119,N_15394,N_15758);
xnor U22120 (N_22120,N_15709,N_15264);
nor U22121 (N_22121,N_19198,N_16176);
or U22122 (N_22122,N_15907,N_15446);
and U22123 (N_22123,N_16631,N_17171);
and U22124 (N_22124,N_19236,N_15361);
and U22125 (N_22125,N_16221,N_15047);
or U22126 (N_22126,N_16317,N_16917);
nand U22127 (N_22127,N_17837,N_16166);
or U22128 (N_22128,N_16187,N_16612);
xor U22129 (N_22129,N_16800,N_17209);
or U22130 (N_22130,N_18830,N_16452);
xnor U22131 (N_22131,N_19679,N_17943);
xnor U22132 (N_22132,N_16211,N_17546);
nand U22133 (N_22133,N_15594,N_18714);
nand U22134 (N_22134,N_16256,N_15820);
nor U22135 (N_22135,N_15591,N_15340);
nand U22136 (N_22136,N_17061,N_16329);
nor U22137 (N_22137,N_18655,N_15174);
and U22138 (N_22138,N_16900,N_19598);
and U22139 (N_22139,N_16132,N_16767);
xnor U22140 (N_22140,N_19291,N_19456);
and U22141 (N_22141,N_16781,N_18513);
or U22142 (N_22142,N_19985,N_18720);
or U22143 (N_22143,N_18897,N_19703);
xor U22144 (N_22144,N_15115,N_15993);
or U22145 (N_22145,N_18749,N_15854);
and U22146 (N_22146,N_17030,N_15843);
xnor U22147 (N_22147,N_15167,N_18351);
nor U22148 (N_22148,N_15540,N_15292);
nor U22149 (N_22149,N_17804,N_18480);
or U22150 (N_22150,N_18535,N_15784);
nand U22151 (N_22151,N_17765,N_19617);
and U22152 (N_22152,N_16432,N_19686);
xor U22153 (N_22153,N_15053,N_19948);
nor U22154 (N_22154,N_17620,N_18431);
nor U22155 (N_22155,N_19683,N_18987);
nor U22156 (N_22156,N_15706,N_16622);
and U22157 (N_22157,N_17673,N_17235);
xor U22158 (N_22158,N_16827,N_15429);
or U22159 (N_22159,N_19551,N_18573);
or U22160 (N_22160,N_19554,N_16543);
xnor U22161 (N_22161,N_15978,N_17160);
and U22162 (N_22162,N_16424,N_18419);
or U22163 (N_22163,N_18712,N_18653);
nor U22164 (N_22164,N_16647,N_19024);
nand U22165 (N_22165,N_19578,N_19860);
nor U22166 (N_22166,N_16878,N_16780);
xor U22167 (N_22167,N_17041,N_17072);
nor U22168 (N_22168,N_17981,N_16707);
xnor U22169 (N_22169,N_18408,N_16491);
and U22170 (N_22170,N_18299,N_18672);
and U22171 (N_22171,N_18482,N_19409);
nor U22172 (N_22172,N_17606,N_18884);
nor U22173 (N_22173,N_18158,N_16397);
xnor U22174 (N_22174,N_19962,N_15170);
nor U22175 (N_22175,N_15520,N_17278);
xor U22176 (N_22176,N_17121,N_17797);
nor U22177 (N_22177,N_17556,N_19204);
xor U22178 (N_22178,N_15897,N_17042);
and U22179 (N_22179,N_17930,N_16511);
xor U22180 (N_22180,N_16959,N_17283);
xor U22181 (N_22181,N_19043,N_17553);
nor U22182 (N_22182,N_15274,N_19654);
nand U22183 (N_22183,N_18659,N_15160);
nor U22184 (N_22184,N_18376,N_18635);
or U22185 (N_22185,N_18563,N_18740);
and U22186 (N_22186,N_19865,N_17775);
xnor U22187 (N_22187,N_19371,N_16968);
and U22188 (N_22188,N_19999,N_19652);
or U22189 (N_22189,N_15003,N_19727);
nor U22190 (N_22190,N_19067,N_17178);
and U22191 (N_22191,N_17767,N_19094);
or U22192 (N_22192,N_16460,N_17424);
xor U22193 (N_22193,N_17586,N_15447);
nor U22194 (N_22194,N_18459,N_16978);
nor U22195 (N_22195,N_18180,N_15995);
and U22196 (N_22196,N_19378,N_16627);
and U22197 (N_22197,N_15647,N_19317);
nand U22198 (N_22198,N_16119,N_17522);
xor U22199 (N_22199,N_17588,N_17331);
and U22200 (N_22200,N_19193,N_15701);
and U22201 (N_22201,N_15507,N_18125);
or U22202 (N_22202,N_15562,N_16270);
and U22203 (N_22203,N_17222,N_16032);
or U22204 (N_22204,N_15976,N_19066);
and U22205 (N_22205,N_18617,N_17139);
and U22206 (N_22206,N_15813,N_19432);
nand U22207 (N_22207,N_18206,N_17592);
or U22208 (N_22208,N_19561,N_18560);
nand U22209 (N_22209,N_17481,N_16740);
or U22210 (N_22210,N_19106,N_18012);
nand U22211 (N_22211,N_17320,N_16204);
and U22212 (N_22212,N_19736,N_18639);
and U22213 (N_22213,N_19899,N_16020);
xnor U22214 (N_22214,N_16640,N_18599);
and U22215 (N_22215,N_15111,N_16146);
or U22216 (N_22216,N_18237,N_16047);
and U22217 (N_22217,N_15011,N_17110);
or U22218 (N_22218,N_16125,N_18748);
and U22219 (N_22219,N_18203,N_19693);
xor U22220 (N_22220,N_15644,N_19608);
nor U22221 (N_22221,N_19518,N_17259);
nand U22222 (N_22222,N_15608,N_19519);
or U22223 (N_22223,N_17044,N_16915);
and U22224 (N_22224,N_17193,N_15467);
xnor U22225 (N_22225,N_17181,N_17410);
xor U22226 (N_22226,N_16345,N_16845);
and U22227 (N_22227,N_16547,N_19854);
xnor U22228 (N_22228,N_17118,N_19535);
or U22229 (N_22229,N_17413,N_15860);
or U22230 (N_22230,N_18014,N_18550);
or U22231 (N_22231,N_18467,N_19981);
and U22232 (N_22232,N_15691,N_17939);
nand U22233 (N_22233,N_19295,N_17185);
nor U22234 (N_22234,N_16677,N_17406);
and U22235 (N_22235,N_19068,N_18288);
xor U22236 (N_22236,N_18489,N_17475);
nand U22237 (N_22237,N_16614,N_16223);
xor U22238 (N_22238,N_19729,N_15856);
nor U22239 (N_22239,N_15029,N_15827);
nand U22240 (N_22240,N_15333,N_19859);
xnor U22241 (N_22241,N_19931,N_18494);
xnor U22242 (N_22242,N_17823,N_16495);
xnor U22243 (N_22243,N_16394,N_19802);
or U22244 (N_22244,N_16970,N_18988);
nor U22245 (N_22245,N_17316,N_17488);
nand U22246 (N_22246,N_16068,N_15376);
nor U22247 (N_22247,N_15543,N_19264);
nand U22248 (N_22248,N_18189,N_15504);
nor U22249 (N_22249,N_16817,N_15042);
xor U22250 (N_22250,N_18418,N_17430);
and U22251 (N_22251,N_15132,N_16942);
and U22252 (N_22252,N_18637,N_15559);
nand U22253 (N_22253,N_18622,N_17624);
xnor U22254 (N_22254,N_18272,N_16358);
xnor U22255 (N_22255,N_17920,N_19135);
nor U22256 (N_22256,N_16005,N_19481);
nand U22257 (N_22257,N_16174,N_19244);
nor U22258 (N_22258,N_19302,N_19974);
and U22259 (N_22259,N_18894,N_16422);
xor U22260 (N_22260,N_19804,N_19002);
or U22261 (N_22261,N_18020,N_17208);
xnor U22262 (N_22262,N_17919,N_16940);
nor U22263 (N_22263,N_15542,N_15204);
and U22264 (N_22264,N_16714,N_17456);
and U22265 (N_22265,N_15931,N_18739);
nand U22266 (N_22266,N_15291,N_17236);
or U22267 (N_22267,N_18334,N_19219);
nor U22268 (N_22268,N_18183,N_19336);
xor U22269 (N_22269,N_16875,N_15779);
nor U22270 (N_22270,N_17527,N_18503);
or U22271 (N_22271,N_17530,N_17264);
xor U22272 (N_22272,N_16637,N_15465);
or U22273 (N_22273,N_16056,N_19419);
xor U22274 (N_22274,N_15679,N_17269);
xnor U22275 (N_22275,N_16391,N_17583);
xor U22276 (N_22276,N_16202,N_19257);
nor U22277 (N_22277,N_16729,N_19920);
or U22278 (N_22278,N_19662,N_18244);
nand U22279 (N_22279,N_16436,N_16553);
or U22280 (N_22280,N_16595,N_15006);
xnor U22281 (N_22281,N_19581,N_17207);
nor U22282 (N_22282,N_19623,N_16947);
nor U22283 (N_22283,N_16349,N_15385);
or U22284 (N_22284,N_16523,N_19208);
or U22285 (N_22285,N_18143,N_17449);
or U22286 (N_22286,N_17262,N_15554);
or U22287 (N_22287,N_17832,N_16214);
or U22288 (N_22288,N_16288,N_15721);
xnor U22289 (N_22289,N_17402,N_18601);
and U22290 (N_22290,N_18543,N_19436);
and U22291 (N_22291,N_19095,N_18647);
nor U22292 (N_22292,N_16026,N_16830);
nor U22293 (N_22293,N_17688,N_15693);
nor U22294 (N_22294,N_18844,N_15349);
or U22295 (N_22295,N_15457,N_19222);
xor U22296 (N_22296,N_17653,N_16429);
and U22297 (N_22297,N_19601,N_18536);
nand U22298 (N_22298,N_17242,N_18096);
and U22299 (N_22299,N_16760,N_18313);
nor U22300 (N_22300,N_16118,N_18153);
and U22301 (N_22301,N_19742,N_18019);
nor U22302 (N_22302,N_17313,N_17887);
xor U22303 (N_22303,N_18717,N_15719);
nand U22304 (N_22304,N_17916,N_16069);
and U22305 (N_22305,N_16567,N_19421);
xnor U22306 (N_22306,N_18088,N_17065);
or U22307 (N_22307,N_15175,N_17701);
or U22308 (N_22308,N_18384,N_17666);
and U22309 (N_22309,N_15014,N_17394);
xnor U22310 (N_22310,N_16786,N_16000);
xnor U22311 (N_22311,N_18006,N_18129);
and U22312 (N_22312,N_19798,N_19359);
xor U22313 (N_22313,N_19116,N_15012);
and U22314 (N_22314,N_16501,N_15092);
nor U22315 (N_22315,N_19327,N_16717);
or U22316 (N_22316,N_18305,N_17233);
or U22317 (N_22317,N_15893,N_15766);
and U22318 (N_22318,N_15018,N_19346);
xor U22319 (N_22319,N_18276,N_18680);
nand U22320 (N_22320,N_16259,N_19808);
nand U22321 (N_22321,N_18207,N_18585);
nand U22322 (N_22322,N_16328,N_15563);
or U22323 (N_22323,N_18154,N_15819);
or U22324 (N_22324,N_15454,N_17120);
xor U22325 (N_22325,N_15762,N_15222);
and U22326 (N_22326,N_18960,N_17774);
and U22327 (N_22327,N_18323,N_17941);
and U22328 (N_22328,N_18574,N_17250);
nand U22329 (N_22329,N_18374,N_16691);
xor U22330 (N_22330,N_15645,N_17323);
and U22331 (N_22331,N_18033,N_15422);
nor U22332 (N_22332,N_19602,N_18404);
nand U22333 (N_22333,N_17921,N_19112);
or U22334 (N_22334,N_17433,N_16694);
nand U22335 (N_22335,N_18318,N_15001);
xnor U22336 (N_22336,N_16675,N_18112);
nand U22337 (N_22337,N_17453,N_19401);
nor U22338 (N_22338,N_15348,N_18731);
xnor U22339 (N_22339,N_16581,N_18868);
or U22340 (N_22340,N_19646,N_17094);
nor U22341 (N_22341,N_18460,N_16273);
xor U22342 (N_22342,N_18878,N_18516);
or U22343 (N_22343,N_17508,N_16261);
nand U22344 (N_22344,N_18769,N_19701);
and U22345 (N_22345,N_19192,N_17218);
and U22346 (N_22346,N_15303,N_16023);
xor U22347 (N_22347,N_16904,N_15345);
and U22348 (N_22348,N_16670,N_17391);
xnor U22349 (N_22349,N_18392,N_18510);
or U22350 (N_22350,N_18269,N_19448);
nor U22351 (N_22351,N_18046,N_17117);
xnor U22352 (N_22352,N_18797,N_17180);
nand U22353 (N_22353,N_15830,N_19433);
or U22354 (N_22354,N_16271,N_19169);
xnor U22355 (N_22355,N_16563,N_15913);
nand U22356 (N_22356,N_19666,N_18363);
or U22357 (N_22357,N_15824,N_17514);
xnor U22358 (N_22358,N_15787,N_16504);
xor U22359 (N_22359,N_17189,N_18939);
and U22360 (N_22360,N_18768,N_17760);
or U22361 (N_22361,N_15927,N_15502);
nand U22362 (N_22362,N_15048,N_17868);
nor U22363 (N_22363,N_18803,N_15636);
or U22364 (N_22364,N_19362,N_19168);
or U22365 (N_22365,N_16220,N_17597);
xnor U22366 (N_22366,N_15865,N_15982);
and U22367 (N_22367,N_15070,N_18865);
or U22368 (N_22368,N_16407,N_17062);
nand U22369 (N_22369,N_18250,N_15234);
xnor U22370 (N_22370,N_17687,N_18643);
and U22371 (N_22371,N_19427,N_15294);
xnor U22372 (N_22372,N_18101,N_17768);
or U22373 (N_22373,N_16484,N_18407);
and U22374 (N_22374,N_17231,N_19000);
xor U22375 (N_22375,N_19753,N_16360);
and U22376 (N_22376,N_15460,N_19914);
or U22377 (N_22377,N_17247,N_16488);
nand U22378 (N_22378,N_18638,N_19072);
nor U22379 (N_22379,N_16194,N_16296);
nand U22380 (N_22380,N_16621,N_18903);
and U22381 (N_22381,N_17682,N_18527);
or U22382 (N_22382,N_16400,N_19772);
or U22383 (N_22383,N_17213,N_16034);
nand U22384 (N_22384,N_15176,N_19873);
and U22385 (N_22385,N_18139,N_15315);
or U22386 (N_22386,N_15894,N_19220);
nor U22387 (N_22387,N_18395,N_19947);
and U22388 (N_22388,N_19088,N_16043);
and U22389 (N_22389,N_15935,N_19555);
or U22390 (N_22390,N_16042,N_17510);
and U22391 (N_22391,N_16816,N_16262);
nand U22392 (N_22392,N_18009,N_15310);
or U22393 (N_22393,N_16149,N_15243);
or U22394 (N_22394,N_19442,N_18952);
nand U22395 (N_22395,N_19816,N_15022);
nor U22396 (N_22396,N_15561,N_15388);
nor U22397 (N_22397,N_17419,N_19634);
or U22398 (N_22398,N_16785,N_16840);
nand U22399 (N_22399,N_16866,N_18707);
and U22400 (N_22400,N_17590,N_17363);
or U22401 (N_22401,N_15612,N_19231);
nor U22402 (N_22402,N_18111,N_19048);
nor U22403 (N_22403,N_17448,N_16983);
nand U22404 (N_22404,N_15934,N_18650);
nand U22405 (N_22405,N_16696,N_18426);
nand U22406 (N_22406,N_18235,N_16963);
xnor U22407 (N_22407,N_18297,N_15057);
and U22408 (N_22408,N_15876,N_16040);
and U22409 (N_22409,N_16611,N_17679);
nand U22410 (N_22410,N_15356,N_15855);
or U22411 (N_22411,N_18286,N_15471);
or U22412 (N_22412,N_18691,N_16442);
nor U22413 (N_22413,N_19467,N_18899);
and U22414 (N_22414,N_16067,N_17856);
and U22415 (N_22415,N_15260,N_18770);
nand U22416 (N_22416,N_19673,N_16748);
nor U22417 (N_22417,N_19367,N_15957);
nor U22418 (N_22418,N_15179,N_18198);
or U22419 (N_22419,N_18534,N_17496);
nand U22420 (N_22420,N_19074,N_19316);
xnor U22421 (N_22421,N_19158,N_15823);
xnor U22422 (N_22422,N_19026,N_16658);
or U22423 (N_22423,N_19975,N_15165);
and U22424 (N_22424,N_19762,N_17729);
or U22425 (N_22425,N_18788,N_16806);
nor U22426 (N_22426,N_16893,N_15522);
xnor U22427 (N_22427,N_16159,N_18367);
or U22428 (N_22428,N_16403,N_17478);
nor U22429 (N_22429,N_18953,N_16492);
nand U22430 (N_22430,N_19786,N_15675);
xnor U22431 (N_22431,N_18945,N_19310);
nand U22432 (N_22432,N_18008,N_19713);
nor U22433 (N_22433,N_18172,N_17412);
xor U22434 (N_22434,N_19033,N_18794);
nand U22435 (N_22435,N_19400,N_15015);
or U22436 (N_22436,N_17871,N_18451);
xnor U22437 (N_22437,N_19005,N_16021);
and U22438 (N_22438,N_16950,N_19775);
nand U22439 (N_22439,N_17998,N_18549);
xnor U22440 (N_22440,N_16971,N_19270);
xnor U22441 (N_22441,N_18781,N_17854);
xor U22442 (N_22442,N_15472,N_15441);
xnor U22443 (N_22443,N_19459,N_19084);
and U22444 (N_22444,N_18013,N_17891);
nor U22445 (N_22445,N_18277,N_19717);
and U22446 (N_22446,N_17169,N_17045);
xnor U22447 (N_22447,N_18200,N_17375);
or U22448 (N_22448,N_15017,N_19707);
xor U22449 (N_22449,N_18486,N_19682);
nor U22450 (N_22450,N_16130,N_16163);
or U22451 (N_22451,N_19846,N_17631);
and U22452 (N_22452,N_16793,N_18245);
and U22453 (N_22453,N_19659,N_18933);
xor U22454 (N_22454,N_16571,N_18814);
nand U22455 (N_22455,N_17068,N_19153);
and U22456 (N_22456,N_17963,N_15013);
nor U22457 (N_22457,N_17608,N_19253);
nor U22458 (N_22458,N_16219,N_19737);
nand U22459 (N_22459,N_17190,N_19385);
xor U22460 (N_22460,N_16373,N_18321);
nor U22461 (N_22461,N_18485,N_17838);
xnor U22462 (N_22462,N_17308,N_19885);
or U22463 (N_22463,N_18848,N_16201);
and U22464 (N_22464,N_15853,N_15738);
xor U22465 (N_22465,N_15909,N_19548);
nand U22466 (N_22466,N_19527,N_19566);
nor U22467 (N_22467,N_18795,N_16295);
and U22468 (N_22468,N_17102,N_18852);
nand U22469 (N_22469,N_17515,N_16960);
nand U22470 (N_22470,N_17902,N_16867);
xor U22471 (N_22471,N_19249,N_17155);
nand U22472 (N_22472,N_18220,N_17537);
nor U22473 (N_22473,N_15479,N_18726);
nor U22474 (N_22474,N_17194,N_18862);
or U22475 (N_22475,N_18820,N_16660);
nand U22476 (N_22476,N_18282,N_17507);
or U22477 (N_22477,N_19660,N_16415);
or U22478 (N_22478,N_18167,N_17829);
or U22479 (N_22479,N_18861,N_18271);
xnor U22480 (N_22480,N_17697,N_15852);
and U22481 (N_22481,N_16542,N_18239);
nand U22482 (N_22482,N_19389,N_19512);
nand U22483 (N_22483,N_19060,N_19871);
nand U22484 (N_22484,N_19605,N_19313);
nor U22485 (N_22485,N_15570,N_19614);
nor U22486 (N_22486,N_16485,N_18860);
xor U22487 (N_22487,N_17626,N_18514);
nand U22488 (N_22488,N_19784,N_18423);
and U22489 (N_22489,N_15382,N_18857);
xor U22490 (N_22490,N_18840,N_15428);
xor U22491 (N_22491,N_15231,N_19907);
xor U22492 (N_22492,N_16648,N_19425);
and U22493 (N_22493,N_17359,N_16090);
or U22494 (N_22494,N_16087,N_15318);
nand U22495 (N_22495,N_15708,N_16476);
or U22496 (N_22496,N_17389,N_16490);
xor U22497 (N_22497,N_18824,N_18980);
nand U22498 (N_22498,N_16776,N_17677);
nand U22499 (N_22499,N_17257,N_15205);
nand U22500 (N_22500,N_16159,N_15744);
nand U22501 (N_22501,N_18473,N_17347);
or U22502 (N_22502,N_16439,N_16827);
or U22503 (N_22503,N_15448,N_15786);
xnor U22504 (N_22504,N_19589,N_18460);
nand U22505 (N_22505,N_17078,N_16886);
xnor U22506 (N_22506,N_18381,N_15441);
nor U22507 (N_22507,N_18440,N_17416);
or U22508 (N_22508,N_18316,N_15040);
xor U22509 (N_22509,N_16222,N_15258);
and U22510 (N_22510,N_18901,N_15115);
or U22511 (N_22511,N_18030,N_17076);
and U22512 (N_22512,N_15809,N_18265);
nand U22513 (N_22513,N_16369,N_19910);
or U22514 (N_22514,N_17013,N_17420);
xor U22515 (N_22515,N_16370,N_16927);
and U22516 (N_22516,N_19554,N_16435);
and U22517 (N_22517,N_19599,N_18211);
and U22518 (N_22518,N_18185,N_18582);
nor U22519 (N_22519,N_19970,N_15206);
nand U22520 (N_22520,N_19619,N_18926);
or U22521 (N_22521,N_19089,N_17613);
or U22522 (N_22522,N_17960,N_15905);
or U22523 (N_22523,N_16143,N_16513);
xnor U22524 (N_22524,N_18588,N_18858);
and U22525 (N_22525,N_17115,N_17072);
xnor U22526 (N_22526,N_15201,N_15330);
or U22527 (N_22527,N_15002,N_18637);
nor U22528 (N_22528,N_17167,N_18280);
nand U22529 (N_22529,N_15838,N_16596);
or U22530 (N_22530,N_18441,N_15070);
and U22531 (N_22531,N_15312,N_17603);
or U22532 (N_22532,N_19380,N_15976);
xor U22533 (N_22533,N_17239,N_16242);
and U22534 (N_22534,N_19044,N_18738);
and U22535 (N_22535,N_18758,N_19217);
nor U22536 (N_22536,N_17113,N_17727);
or U22537 (N_22537,N_18826,N_15027);
nor U22538 (N_22538,N_18379,N_17058);
nor U22539 (N_22539,N_19178,N_15645);
xnor U22540 (N_22540,N_17881,N_15929);
or U22541 (N_22541,N_16034,N_19254);
nor U22542 (N_22542,N_19867,N_18315);
nor U22543 (N_22543,N_15071,N_15275);
nor U22544 (N_22544,N_15067,N_15117);
and U22545 (N_22545,N_17186,N_18788);
and U22546 (N_22546,N_18790,N_19104);
nor U22547 (N_22547,N_19647,N_16533);
nor U22548 (N_22548,N_19176,N_18760);
nor U22549 (N_22549,N_17381,N_15663);
or U22550 (N_22550,N_18882,N_19365);
and U22551 (N_22551,N_17717,N_17169);
nor U22552 (N_22552,N_18747,N_15094);
nand U22553 (N_22553,N_17537,N_16131);
xor U22554 (N_22554,N_17490,N_19204);
or U22555 (N_22555,N_19349,N_18468);
xor U22556 (N_22556,N_18348,N_16849);
xor U22557 (N_22557,N_15011,N_18947);
xor U22558 (N_22558,N_18149,N_16780);
nor U22559 (N_22559,N_16957,N_16224);
nand U22560 (N_22560,N_19459,N_18657);
or U22561 (N_22561,N_19171,N_15322);
or U22562 (N_22562,N_18062,N_19866);
xnor U22563 (N_22563,N_19404,N_18108);
or U22564 (N_22564,N_19078,N_19959);
xor U22565 (N_22565,N_17851,N_16336);
xor U22566 (N_22566,N_19255,N_17200);
and U22567 (N_22567,N_17346,N_17643);
nand U22568 (N_22568,N_17066,N_18473);
nor U22569 (N_22569,N_16794,N_17282);
or U22570 (N_22570,N_18312,N_18523);
and U22571 (N_22571,N_17772,N_17353);
nor U22572 (N_22572,N_15905,N_19404);
nand U22573 (N_22573,N_19857,N_19480);
nand U22574 (N_22574,N_19709,N_19625);
or U22575 (N_22575,N_17591,N_19452);
xor U22576 (N_22576,N_17320,N_17210);
nor U22577 (N_22577,N_17946,N_16466);
or U22578 (N_22578,N_15664,N_15346);
or U22579 (N_22579,N_17272,N_18865);
xor U22580 (N_22580,N_17372,N_18636);
xnor U22581 (N_22581,N_16891,N_19643);
or U22582 (N_22582,N_17645,N_16075);
nor U22583 (N_22583,N_17613,N_18949);
nor U22584 (N_22584,N_16598,N_16178);
or U22585 (N_22585,N_17311,N_18700);
nor U22586 (N_22586,N_18236,N_17344);
or U22587 (N_22587,N_16333,N_16025);
nor U22588 (N_22588,N_19520,N_17877);
or U22589 (N_22589,N_15690,N_18306);
or U22590 (N_22590,N_16908,N_19828);
nor U22591 (N_22591,N_19075,N_17286);
xor U22592 (N_22592,N_15526,N_18681);
and U22593 (N_22593,N_16233,N_17244);
or U22594 (N_22594,N_19437,N_17238);
or U22595 (N_22595,N_16525,N_15923);
or U22596 (N_22596,N_15066,N_16168);
or U22597 (N_22597,N_17631,N_17513);
and U22598 (N_22598,N_17422,N_15196);
nand U22599 (N_22599,N_17148,N_18753);
nor U22600 (N_22600,N_19348,N_15739);
or U22601 (N_22601,N_17739,N_18184);
nor U22602 (N_22602,N_18720,N_16011);
nor U22603 (N_22603,N_15719,N_17886);
nor U22604 (N_22604,N_19262,N_18704);
nand U22605 (N_22605,N_16394,N_17773);
and U22606 (N_22606,N_19807,N_19465);
or U22607 (N_22607,N_18001,N_15912);
nand U22608 (N_22608,N_19123,N_16804);
and U22609 (N_22609,N_17779,N_19584);
nand U22610 (N_22610,N_18024,N_15195);
or U22611 (N_22611,N_18385,N_18894);
xor U22612 (N_22612,N_15776,N_17416);
and U22613 (N_22613,N_16392,N_18409);
nand U22614 (N_22614,N_17241,N_19845);
or U22615 (N_22615,N_16968,N_15313);
nand U22616 (N_22616,N_19178,N_19208);
or U22617 (N_22617,N_16694,N_17423);
xnor U22618 (N_22618,N_15828,N_16934);
xor U22619 (N_22619,N_15910,N_19511);
or U22620 (N_22620,N_16433,N_17656);
xnor U22621 (N_22621,N_17747,N_18362);
and U22622 (N_22622,N_15462,N_15719);
and U22623 (N_22623,N_17721,N_15400);
nor U22624 (N_22624,N_15377,N_17975);
nor U22625 (N_22625,N_18401,N_18069);
and U22626 (N_22626,N_16778,N_18663);
or U22627 (N_22627,N_17340,N_16589);
and U22628 (N_22628,N_15733,N_16498);
and U22629 (N_22629,N_15008,N_15888);
xnor U22630 (N_22630,N_18627,N_17123);
nor U22631 (N_22631,N_19221,N_15701);
nand U22632 (N_22632,N_19726,N_16614);
xnor U22633 (N_22633,N_17304,N_15352);
and U22634 (N_22634,N_19411,N_16963);
and U22635 (N_22635,N_15977,N_18988);
and U22636 (N_22636,N_18935,N_18545);
nand U22637 (N_22637,N_17014,N_15119);
xnor U22638 (N_22638,N_18854,N_18428);
and U22639 (N_22639,N_19707,N_16386);
and U22640 (N_22640,N_19356,N_15918);
nor U22641 (N_22641,N_15547,N_17606);
and U22642 (N_22642,N_15443,N_18440);
nand U22643 (N_22643,N_19853,N_17221);
nor U22644 (N_22644,N_16918,N_19570);
xor U22645 (N_22645,N_17589,N_18455);
xor U22646 (N_22646,N_17128,N_18024);
nand U22647 (N_22647,N_17434,N_17315);
nand U22648 (N_22648,N_19475,N_19639);
nand U22649 (N_22649,N_15502,N_15713);
and U22650 (N_22650,N_18690,N_19059);
and U22651 (N_22651,N_18681,N_17596);
nor U22652 (N_22652,N_18101,N_19691);
xor U22653 (N_22653,N_19823,N_17622);
nand U22654 (N_22654,N_16673,N_19964);
nand U22655 (N_22655,N_19807,N_17305);
nor U22656 (N_22656,N_18435,N_17132);
nor U22657 (N_22657,N_17694,N_17677);
and U22658 (N_22658,N_19068,N_16073);
nor U22659 (N_22659,N_15287,N_18406);
or U22660 (N_22660,N_16202,N_17342);
xnor U22661 (N_22661,N_19403,N_19992);
nor U22662 (N_22662,N_19164,N_19230);
and U22663 (N_22663,N_16712,N_18240);
or U22664 (N_22664,N_16753,N_15071);
or U22665 (N_22665,N_15552,N_16166);
and U22666 (N_22666,N_16447,N_19909);
or U22667 (N_22667,N_18904,N_18847);
or U22668 (N_22668,N_18586,N_15209);
nand U22669 (N_22669,N_15003,N_19606);
or U22670 (N_22670,N_16792,N_16384);
or U22671 (N_22671,N_18270,N_17293);
xor U22672 (N_22672,N_15830,N_16525);
nor U22673 (N_22673,N_16031,N_18569);
nor U22674 (N_22674,N_16042,N_16169);
or U22675 (N_22675,N_17230,N_17150);
xnor U22676 (N_22676,N_16749,N_19054);
and U22677 (N_22677,N_16423,N_16706);
nor U22678 (N_22678,N_19787,N_19419);
or U22679 (N_22679,N_15419,N_15534);
nor U22680 (N_22680,N_19726,N_18345);
xnor U22681 (N_22681,N_19642,N_18420);
nor U22682 (N_22682,N_19868,N_15355);
or U22683 (N_22683,N_15017,N_17291);
and U22684 (N_22684,N_16034,N_16806);
nand U22685 (N_22685,N_19745,N_17056);
nand U22686 (N_22686,N_18605,N_19219);
nand U22687 (N_22687,N_17044,N_15525);
nand U22688 (N_22688,N_16487,N_19176);
or U22689 (N_22689,N_17421,N_16283);
and U22690 (N_22690,N_16218,N_15246);
or U22691 (N_22691,N_17719,N_16001);
xor U22692 (N_22692,N_18323,N_18955);
or U22693 (N_22693,N_19073,N_16550);
and U22694 (N_22694,N_17511,N_15973);
xnor U22695 (N_22695,N_17575,N_18638);
nand U22696 (N_22696,N_18525,N_18432);
and U22697 (N_22697,N_18206,N_19964);
or U22698 (N_22698,N_16346,N_15180);
and U22699 (N_22699,N_17795,N_17816);
nand U22700 (N_22700,N_18153,N_16110);
xor U22701 (N_22701,N_17343,N_15934);
nand U22702 (N_22702,N_19554,N_19588);
nor U22703 (N_22703,N_16313,N_15635);
or U22704 (N_22704,N_15394,N_16529);
and U22705 (N_22705,N_17831,N_18487);
nand U22706 (N_22706,N_19712,N_19367);
nand U22707 (N_22707,N_17488,N_17538);
and U22708 (N_22708,N_18257,N_18859);
and U22709 (N_22709,N_16478,N_19201);
nor U22710 (N_22710,N_15082,N_17922);
nand U22711 (N_22711,N_15029,N_18400);
or U22712 (N_22712,N_18308,N_17265);
nor U22713 (N_22713,N_16802,N_15225);
nor U22714 (N_22714,N_15512,N_17516);
nand U22715 (N_22715,N_15714,N_19489);
and U22716 (N_22716,N_15420,N_16975);
nand U22717 (N_22717,N_16255,N_19038);
nor U22718 (N_22718,N_15884,N_18120);
xnor U22719 (N_22719,N_18866,N_15569);
nand U22720 (N_22720,N_19614,N_19297);
nand U22721 (N_22721,N_16715,N_15664);
nor U22722 (N_22722,N_15321,N_17248);
and U22723 (N_22723,N_15515,N_19037);
xor U22724 (N_22724,N_18018,N_18339);
nor U22725 (N_22725,N_19735,N_16643);
nor U22726 (N_22726,N_18622,N_16655);
nor U22727 (N_22727,N_16225,N_16843);
nand U22728 (N_22728,N_17130,N_15767);
or U22729 (N_22729,N_18950,N_17798);
nand U22730 (N_22730,N_16669,N_16318);
nand U22731 (N_22731,N_18665,N_19061);
or U22732 (N_22732,N_19010,N_17625);
nor U22733 (N_22733,N_18629,N_19815);
xnor U22734 (N_22734,N_15917,N_18651);
or U22735 (N_22735,N_15188,N_16459);
or U22736 (N_22736,N_15740,N_17357);
nand U22737 (N_22737,N_19218,N_17296);
xor U22738 (N_22738,N_18442,N_15215);
nor U22739 (N_22739,N_17774,N_17385);
or U22740 (N_22740,N_17963,N_15496);
xnor U22741 (N_22741,N_15511,N_17198);
xnor U22742 (N_22742,N_19620,N_16277);
nor U22743 (N_22743,N_15738,N_19874);
xor U22744 (N_22744,N_19275,N_19246);
nor U22745 (N_22745,N_16095,N_18993);
and U22746 (N_22746,N_19452,N_17500);
or U22747 (N_22747,N_15278,N_17659);
xor U22748 (N_22748,N_15819,N_17118);
or U22749 (N_22749,N_19204,N_17795);
and U22750 (N_22750,N_16449,N_19193);
and U22751 (N_22751,N_17895,N_18685);
and U22752 (N_22752,N_18903,N_19928);
or U22753 (N_22753,N_18531,N_15083);
and U22754 (N_22754,N_17249,N_15615);
or U22755 (N_22755,N_19830,N_18192);
or U22756 (N_22756,N_18354,N_19315);
or U22757 (N_22757,N_17219,N_16789);
nand U22758 (N_22758,N_19931,N_17986);
nor U22759 (N_22759,N_15319,N_18069);
and U22760 (N_22760,N_18788,N_16570);
nand U22761 (N_22761,N_15860,N_15213);
and U22762 (N_22762,N_18952,N_16853);
nand U22763 (N_22763,N_17309,N_17996);
or U22764 (N_22764,N_19309,N_16339);
and U22765 (N_22765,N_19165,N_18776);
nor U22766 (N_22766,N_18763,N_15569);
and U22767 (N_22767,N_15938,N_16409);
nand U22768 (N_22768,N_15173,N_15641);
and U22769 (N_22769,N_17624,N_18403);
nand U22770 (N_22770,N_18231,N_17737);
nor U22771 (N_22771,N_17508,N_16013);
and U22772 (N_22772,N_19847,N_17519);
xor U22773 (N_22773,N_18388,N_18465);
and U22774 (N_22774,N_18415,N_15730);
nand U22775 (N_22775,N_16975,N_15685);
and U22776 (N_22776,N_18157,N_15278);
nand U22777 (N_22777,N_15478,N_18635);
or U22778 (N_22778,N_17794,N_19654);
and U22779 (N_22779,N_18140,N_18463);
or U22780 (N_22780,N_19004,N_17329);
or U22781 (N_22781,N_15356,N_19647);
nand U22782 (N_22782,N_16442,N_15151);
or U22783 (N_22783,N_16843,N_17562);
and U22784 (N_22784,N_18926,N_18542);
xor U22785 (N_22785,N_16151,N_17673);
nand U22786 (N_22786,N_18433,N_16121);
nor U22787 (N_22787,N_16769,N_19552);
nor U22788 (N_22788,N_16958,N_15584);
or U22789 (N_22789,N_19528,N_17021);
or U22790 (N_22790,N_15365,N_17646);
or U22791 (N_22791,N_18965,N_15264);
or U22792 (N_22792,N_18658,N_16720);
and U22793 (N_22793,N_19986,N_17950);
nor U22794 (N_22794,N_18824,N_18376);
xor U22795 (N_22795,N_15596,N_19463);
and U22796 (N_22796,N_17666,N_17754);
xor U22797 (N_22797,N_18351,N_18899);
or U22798 (N_22798,N_16159,N_17254);
nor U22799 (N_22799,N_19924,N_17756);
nand U22800 (N_22800,N_19675,N_15932);
and U22801 (N_22801,N_16905,N_16285);
xnor U22802 (N_22802,N_17534,N_18142);
nor U22803 (N_22803,N_17254,N_19991);
and U22804 (N_22804,N_16515,N_19630);
and U22805 (N_22805,N_19160,N_18561);
xnor U22806 (N_22806,N_15853,N_16561);
xnor U22807 (N_22807,N_19286,N_16276);
nand U22808 (N_22808,N_15892,N_15466);
and U22809 (N_22809,N_18885,N_17365);
nor U22810 (N_22810,N_15998,N_19845);
nor U22811 (N_22811,N_16075,N_19777);
nor U22812 (N_22812,N_15968,N_15253);
xnor U22813 (N_22813,N_17332,N_15337);
or U22814 (N_22814,N_19355,N_15806);
nand U22815 (N_22815,N_19971,N_15747);
nand U22816 (N_22816,N_18463,N_18065);
nor U22817 (N_22817,N_15985,N_18615);
and U22818 (N_22818,N_19931,N_15942);
nor U22819 (N_22819,N_15487,N_16271);
or U22820 (N_22820,N_19324,N_19477);
or U22821 (N_22821,N_15690,N_16761);
or U22822 (N_22822,N_16896,N_16312);
or U22823 (N_22823,N_17635,N_16121);
and U22824 (N_22824,N_18081,N_16156);
and U22825 (N_22825,N_16145,N_15415);
nor U22826 (N_22826,N_15964,N_15124);
or U22827 (N_22827,N_15856,N_15129);
nand U22828 (N_22828,N_16802,N_16350);
and U22829 (N_22829,N_18327,N_16726);
nor U22830 (N_22830,N_18530,N_17075);
xnor U22831 (N_22831,N_19701,N_19035);
or U22832 (N_22832,N_16738,N_18517);
nor U22833 (N_22833,N_19539,N_18398);
and U22834 (N_22834,N_15142,N_16453);
nor U22835 (N_22835,N_18774,N_15871);
nand U22836 (N_22836,N_15656,N_18561);
xor U22837 (N_22837,N_18773,N_18047);
or U22838 (N_22838,N_18062,N_16927);
nand U22839 (N_22839,N_16093,N_16817);
nand U22840 (N_22840,N_17543,N_15736);
nor U22841 (N_22841,N_16480,N_18367);
or U22842 (N_22842,N_17419,N_15298);
or U22843 (N_22843,N_18638,N_19509);
xor U22844 (N_22844,N_16921,N_18523);
nand U22845 (N_22845,N_16378,N_15076);
xor U22846 (N_22846,N_16536,N_17086);
and U22847 (N_22847,N_15932,N_19297);
nor U22848 (N_22848,N_16401,N_16550);
nor U22849 (N_22849,N_19584,N_17331);
nor U22850 (N_22850,N_16457,N_15946);
nor U22851 (N_22851,N_19786,N_17165);
nand U22852 (N_22852,N_18419,N_16267);
nor U22853 (N_22853,N_17135,N_15654);
and U22854 (N_22854,N_16179,N_18090);
nand U22855 (N_22855,N_18360,N_19832);
xor U22856 (N_22856,N_16415,N_15496);
nand U22857 (N_22857,N_17478,N_15436);
nor U22858 (N_22858,N_15219,N_17095);
nand U22859 (N_22859,N_19437,N_15995);
nand U22860 (N_22860,N_19383,N_15988);
xor U22861 (N_22861,N_15218,N_17796);
xnor U22862 (N_22862,N_15279,N_17874);
nor U22863 (N_22863,N_16023,N_17537);
or U22864 (N_22864,N_17041,N_19186);
nor U22865 (N_22865,N_19367,N_16875);
or U22866 (N_22866,N_19214,N_15242);
nor U22867 (N_22867,N_15857,N_18241);
nand U22868 (N_22868,N_15704,N_15019);
or U22869 (N_22869,N_17137,N_16145);
nor U22870 (N_22870,N_18438,N_17868);
xor U22871 (N_22871,N_19932,N_18288);
or U22872 (N_22872,N_19834,N_19452);
nor U22873 (N_22873,N_18030,N_15112);
or U22874 (N_22874,N_17163,N_15928);
and U22875 (N_22875,N_15672,N_18140);
and U22876 (N_22876,N_15327,N_18808);
or U22877 (N_22877,N_15104,N_15246);
and U22878 (N_22878,N_18279,N_18836);
and U22879 (N_22879,N_19305,N_16594);
nor U22880 (N_22880,N_16932,N_19458);
nand U22881 (N_22881,N_16789,N_19655);
nand U22882 (N_22882,N_15788,N_18351);
nor U22883 (N_22883,N_16193,N_18277);
or U22884 (N_22884,N_18855,N_15489);
and U22885 (N_22885,N_15558,N_18330);
and U22886 (N_22886,N_17500,N_17355);
xor U22887 (N_22887,N_15298,N_19636);
xor U22888 (N_22888,N_17344,N_19674);
nand U22889 (N_22889,N_17858,N_17211);
or U22890 (N_22890,N_19941,N_16839);
xor U22891 (N_22891,N_17280,N_17895);
xor U22892 (N_22892,N_19401,N_15758);
nand U22893 (N_22893,N_19655,N_18650);
nor U22894 (N_22894,N_18460,N_19812);
and U22895 (N_22895,N_17990,N_17260);
and U22896 (N_22896,N_19287,N_17496);
nand U22897 (N_22897,N_15344,N_17726);
and U22898 (N_22898,N_19723,N_19249);
nor U22899 (N_22899,N_19423,N_15104);
and U22900 (N_22900,N_18463,N_15195);
xnor U22901 (N_22901,N_17087,N_15378);
and U22902 (N_22902,N_16745,N_15633);
and U22903 (N_22903,N_17520,N_18042);
nor U22904 (N_22904,N_18350,N_17667);
nand U22905 (N_22905,N_18387,N_19823);
and U22906 (N_22906,N_17361,N_16250);
nor U22907 (N_22907,N_15487,N_18298);
xnor U22908 (N_22908,N_18773,N_15800);
nor U22909 (N_22909,N_16222,N_16902);
nand U22910 (N_22910,N_15958,N_17728);
or U22911 (N_22911,N_15907,N_17026);
xnor U22912 (N_22912,N_16051,N_16283);
or U22913 (N_22913,N_16513,N_18715);
nand U22914 (N_22914,N_18552,N_15601);
nand U22915 (N_22915,N_15234,N_18554);
xnor U22916 (N_22916,N_17436,N_19129);
or U22917 (N_22917,N_18245,N_15278);
or U22918 (N_22918,N_17452,N_17106);
xnor U22919 (N_22919,N_17646,N_16256);
or U22920 (N_22920,N_19170,N_15107);
nor U22921 (N_22921,N_18553,N_15469);
and U22922 (N_22922,N_19999,N_16602);
or U22923 (N_22923,N_18326,N_16555);
and U22924 (N_22924,N_19141,N_15877);
nand U22925 (N_22925,N_17748,N_19974);
xor U22926 (N_22926,N_15618,N_17072);
nand U22927 (N_22927,N_17494,N_16875);
nor U22928 (N_22928,N_15753,N_15835);
or U22929 (N_22929,N_19836,N_17132);
and U22930 (N_22930,N_15738,N_17603);
xnor U22931 (N_22931,N_18836,N_16686);
nand U22932 (N_22932,N_19549,N_15490);
nor U22933 (N_22933,N_15527,N_19656);
nor U22934 (N_22934,N_19530,N_15712);
nor U22935 (N_22935,N_19761,N_18539);
or U22936 (N_22936,N_16798,N_18888);
or U22937 (N_22937,N_15892,N_16831);
or U22938 (N_22938,N_19676,N_18476);
nand U22939 (N_22939,N_15502,N_15963);
and U22940 (N_22940,N_18529,N_16055);
nor U22941 (N_22941,N_19485,N_17699);
nor U22942 (N_22942,N_16443,N_15158);
xor U22943 (N_22943,N_19301,N_16125);
or U22944 (N_22944,N_16288,N_18424);
nor U22945 (N_22945,N_16392,N_16129);
nor U22946 (N_22946,N_16239,N_18245);
xnor U22947 (N_22947,N_16497,N_18779);
and U22948 (N_22948,N_15980,N_17003);
nor U22949 (N_22949,N_19909,N_16248);
nand U22950 (N_22950,N_17725,N_18489);
nand U22951 (N_22951,N_16666,N_17776);
nand U22952 (N_22952,N_19933,N_18175);
xnor U22953 (N_22953,N_16005,N_15268);
or U22954 (N_22954,N_19795,N_18717);
xor U22955 (N_22955,N_18448,N_19218);
nand U22956 (N_22956,N_16695,N_19815);
xor U22957 (N_22957,N_17541,N_18981);
nor U22958 (N_22958,N_18400,N_19188);
or U22959 (N_22959,N_19051,N_18641);
or U22960 (N_22960,N_16177,N_19659);
nor U22961 (N_22961,N_18536,N_16967);
and U22962 (N_22962,N_18151,N_15047);
nand U22963 (N_22963,N_18605,N_18009);
or U22964 (N_22964,N_18279,N_19451);
xor U22965 (N_22965,N_19426,N_17386);
xnor U22966 (N_22966,N_18596,N_16972);
nand U22967 (N_22967,N_19878,N_19533);
nand U22968 (N_22968,N_17553,N_17400);
nand U22969 (N_22969,N_18721,N_16250);
or U22970 (N_22970,N_17841,N_17148);
nand U22971 (N_22971,N_16105,N_16014);
nand U22972 (N_22972,N_15257,N_15845);
nor U22973 (N_22973,N_18879,N_16375);
or U22974 (N_22974,N_17378,N_19458);
nand U22975 (N_22975,N_16913,N_19817);
nand U22976 (N_22976,N_18262,N_18543);
or U22977 (N_22977,N_19829,N_16868);
xnor U22978 (N_22978,N_17440,N_17251);
nand U22979 (N_22979,N_15882,N_16834);
nand U22980 (N_22980,N_16450,N_19450);
or U22981 (N_22981,N_19058,N_18032);
nand U22982 (N_22982,N_15072,N_19042);
and U22983 (N_22983,N_19239,N_17168);
nor U22984 (N_22984,N_15096,N_18501);
and U22985 (N_22985,N_17708,N_16800);
and U22986 (N_22986,N_15262,N_17942);
nand U22987 (N_22987,N_15538,N_17422);
xor U22988 (N_22988,N_18815,N_18951);
or U22989 (N_22989,N_18887,N_16093);
xnor U22990 (N_22990,N_18518,N_15135);
nor U22991 (N_22991,N_18753,N_19706);
and U22992 (N_22992,N_16084,N_16445);
nor U22993 (N_22993,N_16848,N_19321);
nand U22994 (N_22994,N_15078,N_15179);
xnor U22995 (N_22995,N_15720,N_15259);
and U22996 (N_22996,N_16813,N_18642);
or U22997 (N_22997,N_18757,N_18606);
or U22998 (N_22998,N_19102,N_18171);
or U22999 (N_22999,N_19306,N_17167);
xor U23000 (N_23000,N_18314,N_16309);
and U23001 (N_23001,N_18301,N_18861);
nand U23002 (N_23002,N_19123,N_19336);
nand U23003 (N_23003,N_18946,N_19460);
or U23004 (N_23004,N_19833,N_17214);
nand U23005 (N_23005,N_16665,N_17543);
or U23006 (N_23006,N_16987,N_16587);
and U23007 (N_23007,N_16781,N_17817);
xor U23008 (N_23008,N_16891,N_16829);
nand U23009 (N_23009,N_16046,N_15926);
xor U23010 (N_23010,N_15003,N_15994);
nand U23011 (N_23011,N_15922,N_18285);
xor U23012 (N_23012,N_15433,N_17895);
nand U23013 (N_23013,N_16803,N_18023);
xor U23014 (N_23014,N_16255,N_16821);
and U23015 (N_23015,N_18816,N_18274);
nor U23016 (N_23016,N_16194,N_17567);
xor U23017 (N_23017,N_19359,N_15802);
nand U23018 (N_23018,N_18112,N_15939);
or U23019 (N_23019,N_17388,N_16117);
nor U23020 (N_23020,N_18915,N_19128);
nand U23021 (N_23021,N_15734,N_17686);
nand U23022 (N_23022,N_17622,N_16565);
nor U23023 (N_23023,N_15271,N_17709);
xor U23024 (N_23024,N_17547,N_17113);
and U23025 (N_23025,N_17160,N_15404);
xnor U23026 (N_23026,N_16140,N_18236);
and U23027 (N_23027,N_15468,N_19869);
and U23028 (N_23028,N_15931,N_16432);
nor U23029 (N_23029,N_18845,N_15241);
and U23030 (N_23030,N_17379,N_18181);
nand U23031 (N_23031,N_18430,N_19576);
nor U23032 (N_23032,N_17719,N_18506);
nand U23033 (N_23033,N_15044,N_16040);
or U23034 (N_23034,N_17656,N_16939);
and U23035 (N_23035,N_18131,N_17891);
xor U23036 (N_23036,N_19263,N_18013);
and U23037 (N_23037,N_16492,N_19690);
nand U23038 (N_23038,N_19307,N_19620);
nand U23039 (N_23039,N_16556,N_16367);
xor U23040 (N_23040,N_17084,N_16399);
or U23041 (N_23041,N_19059,N_16007);
or U23042 (N_23042,N_15837,N_15144);
and U23043 (N_23043,N_19670,N_16495);
xor U23044 (N_23044,N_19632,N_16346);
nor U23045 (N_23045,N_18692,N_17764);
nand U23046 (N_23046,N_16903,N_18395);
or U23047 (N_23047,N_18251,N_18371);
nor U23048 (N_23048,N_17881,N_16436);
and U23049 (N_23049,N_19758,N_16064);
or U23050 (N_23050,N_19006,N_15292);
and U23051 (N_23051,N_17128,N_17904);
nor U23052 (N_23052,N_17475,N_15134);
or U23053 (N_23053,N_19731,N_17886);
nand U23054 (N_23054,N_18947,N_17890);
xnor U23055 (N_23055,N_18177,N_15266);
and U23056 (N_23056,N_17886,N_19907);
or U23057 (N_23057,N_19508,N_19615);
or U23058 (N_23058,N_19936,N_18554);
nand U23059 (N_23059,N_17881,N_15147);
xor U23060 (N_23060,N_19563,N_17710);
nor U23061 (N_23061,N_16821,N_16487);
nand U23062 (N_23062,N_17351,N_18958);
or U23063 (N_23063,N_15003,N_19785);
or U23064 (N_23064,N_18394,N_18038);
and U23065 (N_23065,N_18628,N_18128);
xor U23066 (N_23066,N_17686,N_16363);
nand U23067 (N_23067,N_19982,N_17671);
or U23068 (N_23068,N_17014,N_15923);
or U23069 (N_23069,N_15564,N_16642);
or U23070 (N_23070,N_16332,N_15328);
nor U23071 (N_23071,N_19478,N_17777);
or U23072 (N_23072,N_19911,N_15403);
xnor U23073 (N_23073,N_18279,N_15493);
nand U23074 (N_23074,N_16188,N_16964);
nand U23075 (N_23075,N_16716,N_18785);
nand U23076 (N_23076,N_19583,N_17030);
and U23077 (N_23077,N_17854,N_15372);
nand U23078 (N_23078,N_18934,N_15274);
nor U23079 (N_23079,N_16794,N_18103);
and U23080 (N_23080,N_19179,N_18304);
nor U23081 (N_23081,N_15380,N_17507);
nand U23082 (N_23082,N_19012,N_15284);
nor U23083 (N_23083,N_17049,N_18165);
and U23084 (N_23084,N_18331,N_19651);
nand U23085 (N_23085,N_16483,N_18906);
nor U23086 (N_23086,N_15112,N_17988);
or U23087 (N_23087,N_19243,N_18986);
and U23088 (N_23088,N_16572,N_16266);
nand U23089 (N_23089,N_19011,N_17891);
nor U23090 (N_23090,N_15331,N_19758);
and U23091 (N_23091,N_19015,N_16067);
and U23092 (N_23092,N_17941,N_19294);
or U23093 (N_23093,N_19349,N_19786);
and U23094 (N_23094,N_15078,N_16092);
or U23095 (N_23095,N_18858,N_17626);
or U23096 (N_23096,N_18831,N_15303);
or U23097 (N_23097,N_19543,N_15663);
and U23098 (N_23098,N_19728,N_16184);
nand U23099 (N_23099,N_16028,N_15860);
nor U23100 (N_23100,N_19507,N_15082);
and U23101 (N_23101,N_15696,N_15871);
or U23102 (N_23102,N_19161,N_16363);
nor U23103 (N_23103,N_15833,N_15060);
nand U23104 (N_23104,N_19440,N_19748);
nand U23105 (N_23105,N_17189,N_17050);
or U23106 (N_23106,N_16715,N_15857);
or U23107 (N_23107,N_17348,N_18555);
and U23108 (N_23108,N_18304,N_17830);
xnor U23109 (N_23109,N_17432,N_16012);
and U23110 (N_23110,N_17122,N_16038);
nand U23111 (N_23111,N_16969,N_17141);
nor U23112 (N_23112,N_18105,N_16524);
nor U23113 (N_23113,N_16125,N_15970);
nor U23114 (N_23114,N_15584,N_16678);
and U23115 (N_23115,N_16446,N_18840);
xor U23116 (N_23116,N_17027,N_15317);
xor U23117 (N_23117,N_19446,N_17797);
xnor U23118 (N_23118,N_17011,N_17511);
nor U23119 (N_23119,N_18239,N_15118);
and U23120 (N_23120,N_17491,N_15928);
and U23121 (N_23121,N_17200,N_19754);
xnor U23122 (N_23122,N_15975,N_15575);
xor U23123 (N_23123,N_15808,N_15738);
nand U23124 (N_23124,N_18322,N_19238);
xor U23125 (N_23125,N_17971,N_15506);
and U23126 (N_23126,N_16317,N_19090);
xnor U23127 (N_23127,N_19321,N_17274);
xor U23128 (N_23128,N_19306,N_16553);
nand U23129 (N_23129,N_17643,N_18130);
xor U23130 (N_23130,N_19769,N_17745);
nor U23131 (N_23131,N_17974,N_15440);
nand U23132 (N_23132,N_17370,N_19557);
nor U23133 (N_23133,N_18181,N_18202);
nor U23134 (N_23134,N_15061,N_15532);
nand U23135 (N_23135,N_15797,N_17311);
nand U23136 (N_23136,N_18121,N_16355);
nor U23137 (N_23137,N_15221,N_17659);
nor U23138 (N_23138,N_19382,N_16429);
nor U23139 (N_23139,N_19484,N_15581);
xor U23140 (N_23140,N_17199,N_15105);
nor U23141 (N_23141,N_18482,N_15493);
and U23142 (N_23142,N_15057,N_19658);
and U23143 (N_23143,N_16404,N_19720);
or U23144 (N_23144,N_18977,N_15725);
nor U23145 (N_23145,N_15290,N_15068);
xnor U23146 (N_23146,N_19429,N_16965);
or U23147 (N_23147,N_16894,N_17455);
nor U23148 (N_23148,N_15611,N_18544);
xnor U23149 (N_23149,N_19328,N_17953);
or U23150 (N_23150,N_16265,N_17719);
nor U23151 (N_23151,N_15306,N_18306);
or U23152 (N_23152,N_18337,N_17212);
or U23153 (N_23153,N_17498,N_19331);
nand U23154 (N_23154,N_19642,N_19760);
nor U23155 (N_23155,N_19301,N_19054);
or U23156 (N_23156,N_15399,N_16556);
or U23157 (N_23157,N_16014,N_19490);
xor U23158 (N_23158,N_15163,N_18244);
nor U23159 (N_23159,N_17280,N_18628);
xnor U23160 (N_23160,N_19845,N_17243);
nand U23161 (N_23161,N_18962,N_17244);
and U23162 (N_23162,N_16472,N_19539);
and U23163 (N_23163,N_15691,N_16033);
xnor U23164 (N_23164,N_18043,N_17353);
nand U23165 (N_23165,N_19704,N_16862);
or U23166 (N_23166,N_17672,N_18776);
and U23167 (N_23167,N_15741,N_16308);
and U23168 (N_23168,N_15821,N_19213);
xnor U23169 (N_23169,N_17012,N_18078);
and U23170 (N_23170,N_15988,N_18624);
and U23171 (N_23171,N_16423,N_17440);
or U23172 (N_23172,N_16071,N_19105);
or U23173 (N_23173,N_19843,N_17524);
nand U23174 (N_23174,N_17533,N_19168);
and U23175 (N_23175,N_15984,N_15356);
nor U23176 (N_23176,N_15629,N_18849);
xnor U23177 (N_23177,N_15607,N_18302);
nand U23178 (N_23178,N_19220,N_16699);
or U23179 (N_23179,N_17406,N_16118);
xor U23180 (N_23180,N_18240,N_19944);
and U23181 (N_23181,N_19818,N_18809);
and U23182 (N_23182,N_16437,N_16415);
and U23183 (N_23183,N_16661,N_17600);
or U23184 (N_23184,N_19222,N_17851);
nand U23185 (N_23185,N_15928,N_15229);
nor U23186 (N_23186,N_15329,N_17627);
nand U23187 (N_23187,N_16111,N_18081);
nor U23188 (N_23188,N_15786,N_19825);
nor U23189 (N_23189,N_17506,N_19481);
nand U23190 (N_23190,N_17313,N_17232);
nand U23191 (N_23191,N_19359,N_19170);
and U23192 (N_23192,N_17942,N_19646);
xnor U23193 (N_23193,N_17057,N_19875);
or U23194 (N_23194,N_17681,N_17400);
or U23195 (N_23195,N_17417,N_16763);
nand U23196 (N_23196,N_16828,N_17547);
nand U23197 (N_23197,N_19359,N_15420);
xor U23198 (N_23198,N_16302,N_17648);
nor U23199 (N_23199,N_17224,N_18822);
xor U23200 (N_23200,N_16073,N_15050);
or U23201 (N_23201,N_16241,N_19443);
nor U23202 (N_23202,N_16485,N_16835);
xor U23203 (N_23203,N_18760,N_15008);
nor U23204 (N_23204,N_17725,N_16442);
nand U23205 (N_23205,N_19731,N_19124);
and U23206 (N_23206,N_18109,N_18261);
nor U23207 (N_23207,N_16147,N_17294);
or U23208 (N_23208,N_16063,N_16587);
nand U23209 (N_23209,N_15806,N_18343);
nand U23210 (N_23210,N_19575,N_16316);
nor U23211 (N_23211,N_18854,N_16708);
xnor U23212 (N_23212,N_18912,N_18442);
xor U23213 (N_23213,N_15294,N_15843);
xor U23214 (N_23214,N_16308,N_15552);
and U23215 (N_23215,N_16457,N_17258);
or U23216 (N_23216,N_17482,N_15017);
nor U23217 (N_23217,N_17254,N_16855);
and U23218 (N_23218,N_17977,N_16521);
nor U23219 (N_23219,N_17925,N_19154);
nor U23220 (N_23220,N_15973,N_15310);
nor U23221 (N_23221,N_18843,N_16606);
nand U23222 (N_23222,N_17652,N_15431);
nor U23223 (N_23223,N_19477,N_15675);
nor U23224 (N_23224,N_19598,N_19430);
and U23225 (N_23225,N_16055,N_17072);
xor U23226 (N_23226,N_18197,N_17721);
and U23227 (N_23227,N_19899,N_15025);
nand U23228 (N_23228,N_15378,N_19196);
and U23229 (N_23229,N_17882,N_16968);
or U23230 (N_23230,N_18993,N_16696);
or U23231 (N_23231,N_15318,N_16960);
and U23232 (N_23232,N_17732,N_19154);
nor U23233 (N_23233,N_19247,N_17223);
xnor U23234 (N_23234,N_17315,N_18001);
xnor U23235 (N_23235,N_18427,N_15202);
and U23236 (N_23236,N_17113,N_18159);
or U23237 (N_23237,N_17583,N_19246);
xnor U23238 (N_23238,N_15265,N_19850);
or U23239 (N_23239,N_19220,N_15863);
and U23240 (N_23240,N_15650,N_16232);
xor U23241 (N_23241,N_18963,N_15571);
and U23242 (N_23242,N_15972,N_19900);
or U23243 (N_23243,N_18540,N_19708);
xnor U23244 (N_23244,N_19915,N_19617);
or U23245 (N_23245,N_15906,N_19501);
and U23246 (N_23246,N_17915,N_18548);
nand U23247 (N_23247,N_19229,N_17870);
nand U23248 (N_23248,N_16290,N_15080);
nand U23249 (N_23249,N_16015,N_17537);
and U23250 (N_23250,N_17668,N_18251);
and U23251 (N_23251,N_15965,N_17652);
nand U23252 (N_23252,N_16504,N_17188);
nand U23253 (N_23253,N_19539,N_16860);
xor U23254 (N_23254,N_17630,N_19629);
nor U23255 (N_23255,N_19478,N_19390);
nor U23256 (N_23256,N_15527,N_17852);
nor U23257 (N_23257,N_15051,N_16057);
or U23258 (N_23258,N_18184,N_18468);
nor U23259 (N_23259,N_18646,N_19161);
and U23260 (N_23260,N_17149,N_18815);
nor U23261 (N_23261,N_17946,N_17195);
and U23262 (N_23262,N_16896,N_17885);
nor U23263 (N_23263,N_19057,N_18815);
nor U23264 (N_23264,N_15845,N_17946);
and U23265 (N_23265,N_16913,N_17314);
nor U23266 (N_23266,N_19585,N_17047);
xnor U23267 (N_23267,N_19502,N_17980);
nor U23268 (N_23268,N_16505,N_16348);
xnor U23269 (N_23269,N_16616,N_16375);
nand U23270 (N_23270,N_19528,N_18007);
or U23271 (N_23271,N_19780,N_17772);
or U23272 (N_23272,N_19938,N_16248);
nor U23273 (N_23273,N_18789,N_15445);
nor U23274 (N_23274,N_17192,N_16244);
nand U23275 (N_23275,N_17288,N_19588);
nand U23276 (N_23276,N_15002,N_18822);
or U23277 (N_23277,N_18299,N_18709);
nand U23278 (N_23278,N_15812,N_18755);
or U23279 (N_23279,N_19594,N_18656);
xnor U23280 (N_23280,N_17033,N_18891);
and U23281 (N_23281,N_19803,N_16682);
nand U23282 (N_23282,N_17240,N_19860);
xnor U23283 (N_23283,N_16000,N_18094);
or U23284 (N_23284,N_16634,N_15488);
nor U23285 (N_23285,N_17786,N_16181);
xnor U23286 (N_23286,N_17510,N_19679);
nand U23287 (N_23287,N_15361,N_15504);
xnor U23288 (N_23288,N_18023,N_16295);
or U23289 (N_23289,N_16514,N_15172);
nor U23290 (N_23290,N_17863,N_16892);
xnor U23291 (N_23291,N_17250,N_19555);
nand U23292 (N_23292,N_16922,N_18574);
nor U23293 (N_23293,N_17831,N_18300);
and U23294 (N_23294,N_15740,N_15412);
and U23295 (N_23295,N_18362,N_15001);
nor U23296 (N_23296,N_18775,N_16348);
or U23297 (N_23297,N_18877,N_16887);
or U23298 (N_23298,N_17239,N_16386);
nor U23299 (N_23299,N_19356,N_15834);
xor U23300 (N_23300,N_18372,N_16747);
and U23301 (N_23301,N_17681,N_18725);
xor U23302 (N_23302,N_18561,N_16832);
nand U23303 (N_23303,N_16914,N_16379);
nor U23304 (N_23304,N_19563,N_17682);
nor U23305 (N_23305,N_15779,N_16719);
xnor U23306 (N_23306,N_19285,N_17024);
nand U23307 (N_23307,N_17663,N_18495);
nand U23308 (N_23308,N_15764,N_15446);
xor U23309 (N_23309,N_18405,N_19756);
nand U23310 (N_23310,N_19825,N_17609);
nand U23311 (N_23311,N_15394,N_19959);
nor U23312 (N_23312,N_16763,N_18470);
nand U23313 (N_23313,N_15988,N_18266);
nand U23314 (N_23314,N_16050,N_17428);
and U23315 (N_23315,N_16235,N_18767);
nand U23316 (N_23316,N_16545,N_16688);
or U23317 (N_23317,N_17816,N_15620);
and U23318 (N_23318,N_19441,N_17345);
xor U23319 (N_23319,N_19092,N_18158);
or U23320 (N_23320,N_15405,N_15879);
nand U23321 (N_23321,N_18501,N_16059);
nor U23322 (N_23322,N_17158,N_18328);
or U23323 (N_23323,N_17581,N_19772);
nand U23324 (N_23324,N_15514,N_15157);
and U23325 (N_23325,N_19909,N_19363);
and U23326 (N_23326,N_18931,N_19383);
nand U23327 (N_23327,N_15042,N_16642);
and U23328 (N_23328,N_16806,N_15184);
or U23329 (N_23329,N_17013,N_19290);
and U23330 (N_23330,N_15064,N_17263);
and U23331 (N_23331,N_16187,N_17413);
nand U23332 (N_23332,N_17548,N_15907);
nor U23333 (N_23333,N_18404,N_19145);
or U23334 (N_23334,N_18054,N_15471);
nand U23335 (N_23335,N_17858,N_15966);
xor U23336 (N_23336,N_15340,N_18800);
and U23337 (N_23337,N_18952,N_17029);
nor U23338 (N_23338,N_16714,N_18401);
xor U23339 (N_23339,N_16750,N_16773);
nor U23340 (N_23340,N_16186,N_18536);
nor U23341 (N_23341,N_16295,N_19539);
xnor U23342 (N_23342,N_17232,N_15284);
xor U23343 (N_23343,N_19208,N_19691);
xnor U23344 (N_23344,N_15455,N_18997);
xnor U23345 (N_23345,N_18606,N_16420);
or U23346 (N_23346,N_19797,N_18879);
nor U23347 (N_23347,N_15395,N_18580);
or U23348 (N_23348,N_19768,N_18011);
nor U23349 (N_23349,N_19289,N_18922);
nor U23350 (N_23350,N_16497,N_18393);
and U23351 (N_23351,N_19919,N_17740);
xor U23352 (N_23352,N_17001,N_17204);
or U23353 (N_23353,N_18307,N_18444);
xor U23354 (N_23354,N_18872,N_19606);
or U23355 (N_23355,N_18909,N_15050);
nor U23356 (N_23356,N_19728,N_17687);
nand U23357 (N_23357,N_16162,N_15093);
xor U23358 (N_23358,N_16311,N_15997);
and U23359 (N_23359,N_16184,N_16393);
nand U23360 (N_23360,N_18925,N_19442);
and U23361 (N_23361,N_16691,N_19715);
nor U23362 (N_23362,N_15442,N_16173);
and U23363 (N_23363,N_15067,N_15712);
nand U23364 (N_23364,N_15104,N_16661);
nand U23365 (N_23365,N_19882,N_15876);
or U23366 (N_23366,N_16605,N_18417);
nand U23367 (N_23367,N_19924,N_17330);
nor U23368 (N_23368,N_17414,N_19648);
and U23369 (N_23369,N_19849,N_17378);
or U23370 (N_23370,N_17377,N_17391);
xnor U23371 (N_23371,N_15368,N_19899);
nor U23372 (N_23372,N_17287,N_18479);
nor U23373 (N_23373,N_17172,N_17678);
xor U23374 (N_23374,N_18391,N_17144);
or U23375 (N_23375,N_16773,N_18491);
or U23376 (N_23376,N_18247,N_19587);
and U23377 (N_23377,N_18736,N_15568);
nand U23378 (N_23378,N_15058,N_18729);
and U23379 (N_23379,N_19417,N_16487);
nor U23380 (N_23380,N_19357,N_15873);
nand U23381 (N_23381,N_19565,N_16768);
and U23382 (N_23382,N_18322,N_17165);
nor U23383 (N_23383,N_16989,N_18968);
nand U23384 (N_23384,N_19480,N_16281);
xnor U23385 (N_23385,N_16421,N_16176);
xor U23386 (N_23386,N_15927,N_16790);
nand U23387 (N_23387,N_18602,N_16444);
and U23388 (N_23388,N_19382,N_15914);
or U23389 (N_23389,N_16802,N_19998);
and U23390 (N_23390,N_16873,N_19387);
nor U23391 (N_23391,N_18014,N_16137);
xnor U23392 (N_23392,N_16737,N_15511);
and U23393 (N_23393,N_19957,N_17696);
xor U23394 (N_23394,N_19366,N_19839);
nand U23395 (N_23395,N_15808,N_17516);
xnor U23396 (N_23396,N_19817,N_16376);
xnor U23397 (N_23397,N_15004,N_19295);
and U23398 (N_23398,N_15311,N_16463);
nor U23399 (N_23399,N_16390,N_19613);
nand U23400 (N_23400,N_15169,N_19320);
nor U23401 (N_23401,N_18807,N_15645);
xnor U23402 (N_23402,N_16096,N_17879);
nor U23403 (N_23403,N_15512,N_19701);
nor U23404 (N_23404,N_16676,N_15397);
and U23405 (N_23405,N_17529,N_16291);
xor U23406 (N_23406,N_15943,N_17058);
and U23407 (N_23407,N_18177,N_18333);
or U23408 (N_23408,N_17052,N_17730);
xnor U23409 (N_23409,N_19486,N_18864);
nand U23410 (N_23410,N_15232,N_16557);
or U23411 (N_23411,N_17685,N_17533);
nand U23412 (N_23412,N_17052,N_15953);
xnor U23413 (N_23413,N_17448,N_18747);
nor U23414 (N_23414,N_15792,N_18388);
nor U23415 (N_23415,N_17563,N_15590);
or U23416 (N_23416,N_16512,N_18749);
or U23417 (N_23417,N_17286,N_15341);
nand U23418 (N_23418,N_18682,N_17586);
xnor U23419 (N_23419,N_17483,N_19578);
nand U23420 (N_23420,N_17742,N_19446);
nor U23421 (N_23421,N_18199,N_18936);
or U23422 (N_23422,N_15418,N_19831);
xor U23423 (N_23423,N_17629,N_16136);
or U23424 (N_23424,N_15821,N_17187);
or U23425 (N_23425,N_15675,N_15412);
or U23426 (N_23426,N_17866,N_17404);
and U23427 (N_23427,N_17835,N_17612);
nor U23428 (N_23428,N_16622,N_17660);
and U23429 (N_23429,N_18865,N_17526);
xor U23430 (N_23430,N_16140,N_19684);
or U23431 (N_23431,N_17983,N_16482);
nor U23432 (N_23432,N_15729,N_19780);
and U23433 (N_23433,N_16921,N_18979);
nand U23434 (N_23434,N_18850,N_19880);
nand U23435 (N_23435,N_15999,N_15249);
nand U23436 (N_23436,N_15424,N_16333);
nor U23437 (N_23437,N_19232,N_19109);
or U23438 (N_23438,N_18492,N_17038);
xor U23439 (N_23439,N_17727,N_19031);
nor U23440 (N_23440,N_19623,N_16526);
nand U23441 (N_23441,N_15803,N_19601);
nand U23442 (N_23442,N_16621,N_16223);
nand U23443 (N_23443,N_16212,N_16716);
nand U23444 (N_23444,N_18224,N_15891);
nand U23445 (N_23445,N_19627,N_17149);
nand U23446 (N_23446,N_19394,N_19449);
and U23447 (N_23447,N_17296,N_19499);
nand U23448 (N_23448,N_16463,N_18479);
nor U23449 (N_23449,N_19200,N_15240);
nand U23450 (N_23450,N_15634,N_15452);
xnor U23451 (N_23451,N_17246,N_18318);
and U23452 (N_23452,N_15254,N_16135);
xnor U23453 (N_23453,N_16353,N_19084);
or U23454 (N_23454,N_15103,N_19068);
nand U23455 (N_23455,N_17510,N_17546);
or U23456 (N_23456,N_16534,N_16404);
or U23457 (N_23457,N_19270,N_19579);
xor U23458 (N_23458,N_15650,N_16843);
or U23459 (N_23459,N_19137,N_15646);
nand U23460 (N_23460,N_17520,N_19649);
nand U23461 (N_23461,N_16169,N_15364);
or U23462 (N_23462,N_15492,N_19131);
or U23463 (N_23463,N_15631,N_18532);
nor U23464 (N_23464,N_15082,N_18217);
xor U23465 (N_23465,N_15717,N_19930);
nor U23466 (N_23466,N_16184,N_15325);
xor U23467 (N_23467,N_17993,N_18938);
or U23468 (N_23468,N_19425,N_19526);
nand U23469 (N_23469,N_16365,N_16096);
xnor U23470 (N_23470,N_15846,N_18548);
nand U23471 (N_23471,N_16775,N_17753);
xnor U23472 (N_23472,N_17371,N_18482);
xor U23473 (N_23473,N_15892,N_18877);
nand U23474 (N_23474,N_19819,N_15384);
nor U23475 (N_23475,N_18616,N_19849);
and U23476 (N_23476,N_15909,N_16628);
nand U23477 (N_23477,N_18268,N_19611);
xnor U23478 (N_23478,N_19025,N_17085);
nor U23479 (N_23479,N_16008,N_15167);
xor U23480 (N_23480,N_16728,N_18877);
nand U23481 (N_23481,N_15712,N_16106);
or U23482 (N_23482,N_17497,N_15784);
nor U23483 (N_23483,N_16129,N_19195);
xnor U23484 (N_23484,N_18909,N_19167);
and U23485 (N_23485,N_15691,N_19696);
nor U23486 (N_23486,N_16040,N_19090);
nand U23487 (N_23487,N_15394,N_15360);
and U23488 (N_23488,N_16622,N_18080);
nor U23489 (N_23489,N_15431,N_16670);
xnor U23490 (N_23490,N_16867,N_18959);
nand U23491 (N_23491,N_19163,N_16350);
or U23492 (N_23492,N_15446,N_15550);
and U23493 (N_23493,N_17557,N_15502);
nor U23494 (N_23494,N_18674,N_15445);
and U23495 (N_23495,N_16051,N_19364);
and U23496 (N_23496,N_17143,N_18675);
or U23497 (N_23497,N_17701,N_19059);
or U23498 (N_23498,N_16736,N_16963);
xnor U23499 (N_23499,N_18172,N_19820);
or U23500 (N_23500,N_17362,N_19372);
nor U23501 (N_23501,N_18716,N_17204);
xor U23502 (N_23502,N_16462,N_18430);
or U23503 (N_23503,N_16641,N_16438);
xnor U23504 (N_23504,N_19849,N_19658);
or U23505 (N_23505,N_16822,N_16692);
nor U23506 (N_23506,N_16528,N_19408);
or U23507 (N_23507,N_18074,N_19262);
xnor U23508 (N_23508,N_15132,N_16027);
and U23509 (N_23509,N_19961,N_16234);
nor U23510 (N_23510,N_15072,N_15496);
xor U23511 (N_23511,N_18583,N_17652);
nand U23512 (N_23512,N_17267,N_15997);
and U23513 (N_23513,N_18040,N_16461);
nor U23514 (N_23514,N_17426,N_16548);
nor U23515 (N_23515,N_19863,N_18297);
nand U23516 (N_23516,N_19004,N_16999);
nor U23517 (N_23517,N_18841,N_16088);
xnor U23518 (N_23518,N_15248,N_15435);
or U23519 (N_23519,N_15550,N_15751);
and U23520 (N_23520,N_19959,N_15778);
nor U23521 (N_23521,N_15551,N_18581);
nor U23522 (N_23522,N_18974,N_17514);
xnor U23523 (N_23523,N_18962,N_17589);
nand U23524 (N_23524,N_15490,N_18159);
nor U23525 (N_23525,N_19395,N_18429);
xnor U23526 (N_23526,N_16419,N_19182);
or U23527 (N_23527,N_16682,N_18469);
nor U23528 (N_23528,N_15477,N_18248);
xor U23529 (N_23529,N_16424,N_16007);
nand U23530 (N_23530,N_16808,N_16726);
and U23531 (N_23531,N_17159,N_16909);
nand U23532 (N_23532,N_15141,N_17648);
nor U23533 (N_23533,N_19143,N_16688);
nor U23534 (N_23534,N_19623,N_16419);
or U23535 (N_23535,N_15817,N_16588);
xor U23536 (N_23536,N_19287,N_16204);
nand U23537 (N_23537,N_19827,N_18544);
xnor U23538 (N_23538,N_15642,N_16112);
nand U23539 (N_23539,N_18909,N_15633);
or U23540 (N_23540,N_16304,N_15394);
xor U23541 (N_23541,N_15979,N_19502);
nor U23542 (N_23542,N_15826,N_18310);
xnor U23543 (N_23543,N_18469,N_18675);
nor U23544 (N_23544,N_15114,N_16662);
xor U23545 (N_23545,N_17130,N_15743);
or U23546 (N_23546,N_16385,N_18058);
nor U23547 (N_23547,N_15709,N_15894);
nor U23548 (N_23548,N_16390,N_15947);
nand U23549 (N_23549,N_19799,N_19401);
nor U23550 (N_23550,N_18817,N_18389);
and U23551 (N_23551,N_18629,N_17538);
and U23552 (N_23552,N_17876,N_17051);
or U23553 (N_23553,N_18781,N_17720);
nand U23554 (N_23554,N_15871,N_15187);
nor U23555 (N_23555,N_18394,N_16876);
nand U23556 (N_23556,N_15234,N_16223);
nand U23557 (N_23557,N_18742,N_16051);
and U23558 (N_23558,N_19599,N_15861);
nand U23559 (N_23559,N_16834,N_17831);
nand U23560 (N_23560,N_17700,N_18608);
or U23561 (N_23561,N_15581,N_15917);
nor U23562 (N_23562,N_17690,N_19174);
and U23563 (N_23563,N_17434,N_15106);
nand U23564 (N_23564,N_19089,N_18306);
xor U23565 (N_23565,N_15544,N_17176);
nand U23566 (N_23566,N_18854,N_15465);
nor U23567 (N_23567,N_17548,N_18457);
xor U23568 (N_23568,N_16726,N_16701);
and U23569 (N_23569,N_15968,N_15810);
nor U23570 (N_23570,N_17951,N_17273);
and U23571 (N_23571,N_16523,N_16378);
and U23572 (N_23572,N_17720,N_18512);
and U23573 (N_23573,N_18398,N_18071);
and U23574 (N_23574,N_16364,N_18740);
nand U23575 (N_23575,N_17418,N_18972);
nand U23576 (N_23576,N_19116,N_18895);
and U23577 (N_23577,N_18587,N_15554);
or U23578 (N_23578,N_19859,N_15027);
nand U23579 (N_23579,N_18779,N_18193);
and U23580 (N_23580,N_16368,N_18668);
and U23581 (N_23581,N_18052,N_18262);
xor U23582 (N_23582,N_19983,N_19658);
nand U23583 (N_23583,N_19407,N_16433);
or U23584 (N_23584,N_18180,N_16152);
and U23585 (N_23585,N_16208,N_18619);
and U23586 (N_23586,N_18075,N_18022);
and U23587 (N_23587,N_16932,N_17138);
nor U23588 (N_23588,N_17652,N_17339);
nand U23589 (N_23589,N_16217,N_18818);
or U23590 (N_23590,N_18532,N_16018);
nand U23591 (N_23591,N_19140,N_18314);
xnor U23592 (N_23592,N_17557,N_18810);
or U23593 (N_23593,N_15524,N_19343);
or U23594 (N_23594,N_16773,N_19057);
nand U23595 (N_23595,N_18733,N_16092);
nand U23596 (N_23596,N_18933,N_19948);
nand U23597 (N_23597,N_18712,N_17536);
or U23598 (N_23598,N_16679,N_17064);
and U23599 (N_23599,N_17388,N_17035);
nand U23600 (N_23600,N_17483,N_19016);
or U23601 (N_23601,N_17933,N_18807);
nor U23602 (N_23602,N_18238,N_15795);
and U23603 (N_23603,N_19314,N_16435);
or U23604 (N_23604,N_16854,N_15533);
or U23605 (N_23605,N_19125,N_15236);
nor U23606 (N_23606,N_17780,N_18678);
and U23607 (N_23607,N_18609,N_16834);
or U23608 (N_23608,N_19606,N_19205);
and U23609 (N_23609,N_18680,N_15389);
and U23610 (N_23610,N_17232,N_19463);
nor U23611 (N_23611,N_18896,N_18097);
nand U23612 (N_23612,N_19109,N_16869);
nand U23613 (N_23613,N_17972,N_17979);
or U23614 (N_23614,N_17722,N_19254);
xnor U23615 (N_23615,N_15164,N_15526);
xnor U23616 (N_23616,N_16049,N_15287);
xor U23617 (N_23617,N_18374,N_16307);
nor U23618 (N_23618,N_15819,N_19653);
xor U23619 (N_23619,N_18995,N_15306);
xor U23620 (N_23620,N_18151,N_17111);
xnor U23621 (N_23621,N_15911,N_15596);
or U23622 (N_23622,N_18005,N_16245);
nor U23623 (N_23623,N_15763,N_19981);
xnor U23624 (N_23624,N_15343,N_18794);
and U23625 (N_23625,N_16547,N_17045);
nand U23626 (N_23626,N_18233,N_15386);
xor U23627 (N_23627,N_16026,N_18630);
nand U23628 (N_23628,N_17844,N_17305);
nor U23629 (N_23629,N_17169,N_19604);
and U23630 (N_23630,N_18937,N_16460);
xor U23631 (N_23631,N_15727,N_16161);
or U23632 (N_23632,N_18320,N_16657);
nand U23633 (N_23633,N_18562,N_18354);
and U23634 (N_23634,N_19271,N_15865);
or U23635 (N_23635,N_16352,N_17010);
and U23636 (N_23636,N_18042,N_16905);
and U23637 (N_23637,N_17493,N_18514);
nor U23638 (N_23638,N_18845,N_18434);
nand U23639 (N_23639,N_16515,N_15414);
nand U23640 (N_23640,N_19574,N_19716);
xnor U23641 (N_23641,N_19039,N_18659);
or U23642 (N_23642,N_15541,N_18692);
nor U23643 (N_23643,N_17440,N_17832);
xnor U23644 (N_23644,N_19574,N_15629);
xnor U23645 (N_23645,N_18092,N_19762);
nand U23646 (N_23646,N_17333,N_19424);
or U23647 (N_23647,N_18083,N_18715);
nand U23648 (N_23648,N_15106,N_15304);
or U23649 (N_23649,N_16318,N_19236);
or U23650 (N_23650,N_19015,N_18529);
and U23651 (N_23651,N_15203,N_16325);
nor U23652 (N_23652,N_16938,N_16928);
nor U23653 (N_23653,N_17364,N_18633);
nand U23654 (N_23654,N_17340,N_16922);
and U23655 (N_23655,N_15319,N_18186);
or U23656 (N_23656,N_16811,N_15638);
nor U23657 (N_23657,N_19980,N_16884);
or U23658 (N_23658,N_19161,N_18927);
and U23659 (N_23659,N_17604,N_16257);
and U23660 (N_23660,N_19268,N_15389);
nand U23661 (N_23661,N_19363,N_16072);
nand U23662 (N_23662,N_15382,N_16527);
nand U23663 (N_23663,N_19506,N_15018);
nor U23664 (N_23664,N_16961,N_19778);
xor U23665 (N_23665,N_16042,N_18897);
and U23666 (N_23666,N_17497,N_18984);
nand U23667 (N_23667,N_15869,N_17813);
and U23668 (N_23668,N_18322,N_18157);
nand U23669 (N_23669,N_18665,N_16571);
nor U23670 (N_23670,N_17239,N_19320);
nor U23671 (N_23671,N_18328,N_17950);
or U23672 (N_23672,N_17575,N_15940);
or U23673 (N_23673,N_17654,N_19182);
nor U23674 (N_23674,N_18355,N_16068);
nand U23675 (N_23675,N_17441,N_17254);
or U23676 (N_23676,N_17898,N_19471);
and U23677 (N_23677,N_17622,N_15165);
nand U23678 (N_23678,N_18346,N_15100);
and U23679 (N_23679,N_16298,N_15572);
xnor U23680 (N_23680,N_16897,N_16922);
and U23681 (N_23681,N_16421,N_17248);
and U23682 (N_23682,N_19965,N_18919);
xnor U23683 (N_23683,N_16463,N_19662);
nand U23684 (N_23684,N_17183,N_16094);
or U23685 (N_23685,N_15151,N_19265);
nand U23686 (N_23686,N_18189,N_16425);
or U23687 (N_23687,N_18080,N_17649);
and U23688 (N_23688,N_17766,N_17049);
nand U23689 (N_23689,N_15460,N_17253);
nand U23690 (N_23690,N_18330,N_18638);
and U23691 (N_23691,N_15368,N_15903);
xnor U23692 (N_23692,N_16104,N_18024);
and U23693 (N_23693,N_18266,N_17653);
or U23694 (N_23694,N_19045,N_18172);
and U23695 (N_23695,N_15000,N_18041);
nand U23696 (N_23696,N_16896,N_15437);
nor U23697 (N_23697,N_15482,N_16417);
and U23698 (N_23698,N_19811,N_17080);
and U23699 (N_23699,N_17702,N_16812);
nor U23700 (N_23700,N_15730,N_19287);
nand U23701 (N_23701,N_15871,N_16477);
xnor U23702 (N_23702,N_17041,N_15509);
xnor U23703 (N_23703,N_15877,N_15039);
nor U23704 (N_23704,N_15838,N_19715);
xor U23705 (N_23705,N_18561,N_15157);
nor U23706 (N_23706,N_17718,N_17969);
nand U23707 (N_23707,N_16628,N_17799);
or U23708 (N_23708,N_18937,N_19050);
nor U23709 (N_23709,N_17539,N_19689);
nor U23710 (N_23710,N_18230,N_19165);
and U23711 (N_23711,N_17402,N_18623);
nand U23712 (N_23712,N_18371,N_19275);
nor U23713 (N_23713,N_15848,N_18971);
or U23714 (N_23714,N_15422,N_15528);
nand U23715 (N_23715,N_18530,N_16773);
nor U23716 (N_23716,N_18004,N_16339);
xnor U23717 (N_23717,N_18848,N_16114);
nor U23718 (N_23718,N_15634,N_15253);
xnor U23719 (N_23719,N_18534,N_18578);
xor U23720 (N_23720,N_15480,N_18933);
nor U23721 (N_23721,N_15475,N_18845);
or U23722 (N_23722,N_17228,N_18072);
xnor U23723 (N_23723,N_18784,N_19022);
nand U23724 (N_23724,N_19445,N_18405);
xnor U23725 (N_23725,N_15422,N_16309);
nand U23726 (N_23726,N_16160,N_15799);
or U23727 (N_23727,N_17720,N_16276);
nor U23728 (N_23728,N_19907,N_16920);
xnor U23729 (N_23729,N_16241,N_16992);
or U23730 (N_23730,N_19943,N_18923);
or U23731 (N_23731,N_15644,N_18088);
xor U23732 (N_23732,N_19574,N_19785);
and U23733 (N_23733,N_15883,N_15665);
and U23734 (N_23734,N_19021,N_17419);
nand U23735 (N_23735,N_18887,N_17835);
xnor U23736 (N_23736,N_18388,N_15000);
xor U23737 (N_23737,N_18521,N_17095);
nand U23738 (N_23738,N_18401,N_17763);
nor U23739 (N_23739,N_17847,N_15769);
nand U23740 (N_23740,N_19997,N_17469);
or U23741 (N_23741,N_15381,N_19068);
nand U23742 (N_23742,N_16597,N_17743);
nand U23743 (N_23743,N_16916,N_19693);
nand U23744 (N_23744,N_15691,N_19219);
and U23745 (N_23745,N_16018,N_18738);
nand U23746 (N_23746,N_18139,N_15712);
xor U23747 (N_23747,N_19763,N_17851);
nand U23748 (N_23748,N_17557,N_16607);
nor U23749 (N_23749,N_15452,N_16272);
nor U23750 (N_23750,N_15029,N_17803);
nor U23751 (N_23751,N_16634,N_18896);
or U23752 (N_23752,N_16701,N_19053);
and U23753 (N_23753,N_17569,N_18976);
nor U23754 (N_23754,N_19917,N_19915);
nand U23755 (N_23755,N_17057,N_17516);
nand U23756 (N_23756,N_15671,N_15340);
and U23757 (N_23757,N_17176,N_19838);
or U23758 (N_23758,N_18696,N_19236);
nor U23759 (N_23759,N_18147,N_16467);
xor U23760 (N_23760,N_19002,N_17884);
nor U23761 (N_23761,N_18932,N_15496);
xnor U23762 (N_23762,N_16264,N_17818);
xor U23763 (N_23763,N_19111,N_18749);
xor U23764 (N_23764,N_15384,N_17916);
nand U23765 (N_23765,N_16177,N_16181);
nand U23766 (N_23766,N_16501,N_17526);
and U23767 (N_23767,N_15067,N_18809);
and U23768 (N_23768,N_18632,N_17224);
nor U23769 (N_23769,N_16765,N_16472);
nor U23770 (N_23770,N_16804,N_19076);
nand U23771 (N_23771,N_15957,N_17681);
and U23772 (N_23772,N_16521,N_18355);
nor U23773 (N_23773,N_15742,N_15514);
nor U23774 (N_23774,N_15975,N_19436);
and U23775 (N_23775,N_19413,N_17506);
and U23776 (N_23776,N_17931,N_19785);
nand U23777 (N_23777,N_15341,N_19590);
nor U23778 (N_23778,N_19645,N_16795);
and U23779 (N_23779,N_19736,N_18101);
xor U23780 (N_23780,N_16752,N_19592);
nor U23781 (N_23781,N_19964,N_16799);
nor U23782 (N_23782,N_18554,N_18742);
nor U23783 (N_23783,N_19961,N_19299);
or U23784 (N_23784,N_19755,N_16558);
nor U23785 (N_23785,N_19227,N_16631);
xor U23786 (N_23786,N_16424,N_16455);
nand U23787 (N_23787,N_18739,N_19148);
or U23788 (N_23788,N_16430,N_17145);
and U23789 (N_23789,N_17037,N_16813);
xor U23790 (N_23790,N_19291,N_15646);
nand U23791 (N_23791,N_19555,N_15317);
and U23792 (N_23792,N_19955,N_16470);
and U23793 (N_23793,N_18294,N_18388);
and U23794 (N_23794,N_18631,N_19996);
xnor U23795 (N_23795,N_19424,N_18241);
and U23796 (N_23796,N_15903,N_16825);
nor U23797 (N_23797,N_16511,N_17394);
nor U23798 (N_23798,N_19147,N_17800);
nand U23799 (N_23799,N_19872,N_18017);
nand U23800 (N_23800,N_18971,N_18777);
or U23801 (N_23801,N_17743,N_16140);
xor U23802 (N_23802,N_18697,N_18561);
nor U23803 (N_23803,N_18085,N_16447);
nand U23804 (N_23804,N_16291,N_18525);
nor U23805 (N_23805,N_19130,N_16067);
or U23806 (N_23806,N_16459,N_18809);
or U23807 (N_23807,N_16588,N_15823);
xnor U23808 (N_23808,N_19648,N_17487);
and U23809 (N_23809,N_19770,N_17046);
and U23810 (N_23810,N_18011,N_16150);
or U23811 (N_23811,N_16659,N_19220);
nor U23812 (N_23812,N_18103,N_19304);
or U23813 (N_23813,N_16394,N_15798);
xor U23814 (N_23814,N_18267,N_19489);
or U23815 (N_23815,N_19503,N_15007);
nor U23816 (N_23816,N_16164,N_19544);
xnor U23817 (N_23817,N_17716,N_16696);
nand U23818 (N_23818,N_16363,N_19830);
and U23819 (N_23819,N_16319,N_19911);
nand U23820 (N_23820,N_16356,N_18419);
xor U23821 (N_23821,N_16746,N_19700);
nand U23822 (N_23822,N_17402,N_19282);
or U23823 (N_23823,N_19580,N_16187);
and U23824 (N_23824,N_15909,N_17720);
nor U23825 (N_23825,N_19787,N_17364);
nor U23826 (N_23826,N_18886,N_18732);
nand U23827 (N_23827,N_16669,N_16566);
and U23828 (N_23828,N_15294,N_17992);
and U23829 (N_23829,N_17157,N_16306);
xor U23830 (N_23830,N_19900,N_15558);
and U23831 (N_23831,N_16959,N_19853);
and U23832 (N_23832,N_17673,N_19718);
xor U23833 (N_23833,N_17469,N_19325);
or U23834 (N_23834,N_18344,N_15110);
or U23835 (N_23835,N_18852,N_17836);
nand U23836 (N_23836,N_15783,N_18716);
and U23837 (N_23837,N_16907,N_16291);
xnor U23838 (N_23838,N_18160,N_16838);
nor U23839 (N_23839,N_16267,N_17771);
nand U23840 (N_23840,N_19908,N_17456);
nor U23841 (N_23841,N_18659,N_18436);
nor U23842 (N_23842,N_16855,N_15092);
xnor U23843 (N_23843,N_17702,N_19230);
and U23844 (N_23844,N_18399,N_19948);
or U23845 (N_23845,N_19436,N_19285);
or U23846 (N_23846,N_18806,N_18914);
xnor U23847 (N_23847,N_16110,N_16711);
and U23848 (N_23848,N_17748,N_16477);
nor U23849 (N_23849,N_17045,N_16243);
nand U23850 (N_23850,N_15919,N_18527);
xor U23851 (N_23851,N_16609,N_16856);
and U23852 (N_23852,N_19867,N_15593);
or U23853 (N_23853,N_18802,N_18808);
nand U23854 (N_23854,N_16872,N_15598);
or U23855 (N_23855,N_16860,N_17749);
nor U23856 (N_23856,N_19165,N_18005);
and U23857 (N_23857,N_17811,N_19187);
nand U23858 (N_23858,N_18691,N_15806);
xor U23859 (N_23859,N_18051,N_19656);
xnor U23860 (N_23860,N_19056,N_18454);
xor U23861 (N_23861,N_17165,N_15617);
nor U23862 (N_23862,N_16519,N_18745);
xor U23863 (N_23863,N_17769,N_16375);
xor U23864 (N_23864,N_17694,N_19300);
nand U23865 (N_23865,N_18944,N_15806);
xor U23866 (N_23866,N_19531,N_18192);
nor U23867 (N_23867,N_18209,N_17909);
nor U23868 (N_23868,N_18170,N_15821);
xnor U23869 (N_23869,N_19235,N_19251);
nand U23870 (N_23870,N_19107,N_18266);
or U23871 (N_23871,N_16037,N_17165);
or U23872 (N_23872,N_16365,N_16422);
and U23873 (N_23873,N_18560,N_15913);
nand U23874 (N_23874,N_15831,N_16281);
nor U23875 (N_23875,N_16444,N_17657);
xnor U23876 (N_23876,N_19807,N_18006);
or U23877 (N_23877,N_19515,N_16381);
or U23878 (N_23878,N_16283,N_17585);
or U23879 (N_23879,N_15679,N_17877);
or U23880 (N_23880,N_16411,N_16350);
nor U23881 (N_23881,N_19355,N_17212);
nand U23882 (N_23882,N_16077,N_17695);
xnor U23883 (N_23883,N_15784,N_15867);
and U23884 (N_23884,N_17258,N_17434);
or U23885 (N_23885,N_15258,N_19120);
nand U23886 (N_23886,N_16782,N_17368);
nor U23887 (N_23887,N_17503,N_16083);
or U23888 (N_23888,N_16781,N_19384);
and U23889 (N_23889,N_17698,N_17579);
or U23890 (N_23890,N_15039,N_19294);
and U23891 (N_23891,N_15845,N_18774);
nor U23892 (N_23892,N_16574,N_15799);
nand U23893 (N_23893,N_19177,N_17902);
nand U23894 (N_23894,N_16716,N_16150);
xor U23895 (N_23895,N_19532,N_18448);
nor U23896 (N_23896,N_16422,N_18685);
nor U23897 (N_23897,N_17061,N_16433);
nand U23898 (N_23898,N_18816,N_17706);
nor U23899 (N_23899,N_16620,N_16384);
nor U23900 (N_23900,N_17152,N_18965);
or U23901 (N_23901,N_16200,N_17718);
nor U23902 (N_23902,N_17156,N_18026);
nand U23903 (N_23903,N_16933,N_17293);
xor U23904 (N_23904,N_15985,N_17418);
or U23905 (N_23905,N_18874,N_17355);
and U23906 (N_23906,N_18728,N_18196);
xnor U23907 (N_23907,N_16120,N_17979);
or U23908 (N_23908,N_15736,N_15479);
xnor U23909 (N_23909,N_17265,N_19504);
nor U23910 (N_23910,N_17036,N_17589);
xor U23911 (N_23911,N_18659,N_16427);
and U23912 (N_23912,N_19944,N_16085);
xor U23913 (N_23913,N_16417,N_18906);
xnor U23914 (N_23914,N_19975,N_19307);
nand U23915 (N_23915,N_17759,N_19689);
or U23916 (N_23916,N_17831,N_19867);
nor U23917 (N_23917,N_15628,N_16911);
nor U23918 (N_23918,N_16261,N_19795);
nor U23919 (N_23919,N_17283,N_18144);
and U23920 (N_23920,N_15800,N_19235);
or U23921 (N_23921,N_18020,N_15979);
nand U23922 (N_23922,N_17315,N_16712);
and U23923 (N_23923,N_17545,N_19680);
and U23924 (N_23924,N_18006,N_19331);
or U23925 (N_23925,N_19133,N_19818);
and U23926 (N_23926,N_15560,N_17152);
nand U23927 (N_23927,N_17331,N_19733);
or U23928 (N_23928,N_16986,N_17016);
nand U23929 (N_23929,N_19910,N_19853);
nand U23930 (N_23930,N_19789,N_17711);
or U23931 (N_23931,N_17229,N_16673);
xor U23932 (N_23932,N_15924,N_16166);
or U23933 (N_23933,N_16067,N_17219);
and U23934 (N_23934,N_17182,N_18838);
and U23935 (N_23935,N_19090,N_17608);
nand U23936 (N_23936,N_19340,N_18316);
nor U23937 (N_23937,N_19070,N_19960);
and U23938 (N_23938,N_18201,N_17386);
nor U23939 (N_23939,N_19438,N_18532);
and U23940 (N_23940,N_15045,N_17035);
or U23941 (N_23941,N_19196,N_17087);
xnor U23942 (N_23942,N_15165,N_15486);
nor U23943 (N_23943,N_18215,N_19237);
nand U23944 (N_23944,N_19819,N_19687);
and U23945 (N_23945,N_18850,N_15889);
or U23946 (N_23946,N_15349,N_15993);
xnor U23947 (N_23947,N_15628,N_19285);
xor U23948 (N_23948,N_18847,N_18857);
and U23949 (N_23949,N_19881,N_17665);
nor U23950 (N_23950,N_16394,N_16374);
xor U23951 (N_23951,N_15356,N_17722);
and U23952 (N_23952,N_18337,N_17990);
or U23953 (N_23953,N_17802,N_16423);
xor U23954 (N_23954,N_19438,N_16930);
nor U23955 (N_23955,N_18476,N_19869);
xnor U23956 (N_23956,N_15899,N_15608);
xnor U23957 (N_23957,N_19132,N_17076);
xor U23958 (N_23958,N_18382,N_19340);
or U23959 (N_23959,N_18676,N_19507);
nor U23960 (N_23960,N_16066,N_15631);
nor U23961 (N_23961,N_17220,N_15471);
nand U23962 (N_23962,N_15585,N_17193);
and U23963 (N_23963,N_18946,N_15824);
and U23964 (N_23964,N_18625,N_17897);
xnor U23965 (N_23965,N_17421,N_16883);
nand U23966 (N_23966,N_15484,N_18404);
nand U23967 (N_23967,N_16995,N_15138);
and U23968 (N_23968,N_19312,N_17731);
nor U23969 (N_23969,N_16604,N_18744);
and U23970 (N_23970,N_16634,N_17246);
nand U23971 (N_23971,N_15982,N_18532);
and U23972 (N_23972,N_15397,N_16095);
nor U23973 (N_23973,N_19056,N_15457);
or U23974 (N_23974,N_16223,N_18720);
nor U23975 (N_23975,N_16001,N_17794);
or U23976 (N_23976,N_18376,N_17434);
nand U23977 (N_23977,N_19703,N_18632);
and U23978 (N_23978,N_15075,N_17791);
or U23979 (N_23979,N_16428,N_16523);
xnor U23980 (N_23980,N_16396,N_18600);
and U23981 (N_23981,N_15589,N_16055);
and U23982 (N_23982,N_16480,N_15215);
and U23983 (N_23983,N_19133,N_15076);
nor U23984 (N_23984,N_15051,N_18153);
xnor U23985 (N_23985,N_19586,N_17852);
or U23986 (N_23986,N_18091,N_17953);
and U23987 (N_23987,N_16549,N_15069);
xnor U23988 (N_23988,N_15523,N_16968);
xor U23989 (N_23989,N_19586,N_15091);
nand U23990 (N_23990,N_15568,N_19803);
nand U23991 (N_23991,N_19624,N_16774);
nor U23992 (N_23992,N_17492,N_15420);
nor U23993 (N_23993,N_18212,N_18065);
nand U23994 (N_23994,N_15054,N_18673);
or U23995 (N_23995,N_19617,N_19459);
and U23996 (N_23996,N_15904,N_18675);
xnor U23997 (N_23997,N_17233,N_17779);
xor U23998 (N_23998,N_17301,N_19931);
nor U23999 (N_23999,N_15065,N_17999);
nand U24000 (N_24000,N_15440,N_19072);
nand U24001 (N_24001,N_16769,N_16088);
or U24002 (N_24002,N_18903,N_19125);
nand U24003 (N_24003,N_18771,N_19447);
or U24004 (N_24004,N_15617,N_19682);
and U24005 (N_24005,N_19559,N_18454);
nand U24006 (N_24006,N_18535,N_19550);
nor U24007 (N_24007,N_18711,N_16994);
or U24008 (N_24008,N_15520,N_17852);
or U24009 (N_24009,N_17952,N_16930);
and U24010 (N_24010,N_17361,N_18680);
xnor U24011 (N_24011,N_18822,N_16605);
nor U24012 (N_24012,N_19008,N_15776);
nor U24013 (N_24013,N_15333,N_19432);
nand U24014 (N_24014,N_17410,N_16151);
nand U24015 (N_24015,N_15962,N_16678);
nor U24016 (N_24016,N_19033,N_17993);
and U24017 (N_24017,N_15866,N_16305);
nor U24018 (N_24018,N_17484,N_19845);
and U24019 (N_24019,N_15943,N_15042);
xor U24020 (N_24020,N_16451,N_19559);
nand U24021 (N_24021,N_16299,N_17171);
nor U24022 (N_24022,N_17255,N_16373);
nand U24023 (N_24023,N_17632,N_15332);
xor U24024 (N_24024,N_16927,N_19931);
nand U24025 (N_24025,N_18036,N_17257);
or U24026 (N_24026,N_16761,N_17060);
and U24027 (N_24027,N_15103,N_16271);
nand U24028 (N_24028,N_17155,N_15916);
xor U24029 (N_24029,N_15250,N_17745);
xnor U24030 (N_24030,N_19357,N_15614);
nor U24031 (N_24031,N_17377,N_18609);
xor U24032 (N_24032,N_17372,N_19731);
and U24033 (N_24033,N_15953,N_16896);
nand U24034 (N_24034,N_17307,N_18594);
nor U24035 (N_24035,N_15051,N_15650);
or U24036 (N_24036,N_18803,N_19973);
nor U24037 (N_24037,N_19171,N_17060);
or U24038 (N_24038,N_19877,N_17649);
nor U24039 (N_24039,N_18987,N_17072);
and U24040 (N_24040,N_16724,N_16977);
nand U24041 (N_24041,N_19445,N_16139);
and U24042 (N_24042,N_15395,N_17496);
nand U24043 (N_24043,N_19697,N_19112);
nor U24044 (N_24044,N_17880,N_17781);
or U24045 (N_24045,N_19125,N_18656);
or U24046 (N_24046,N_17016,N_15339);
nor U24047 (N_24047,N_19667,N_17160);
nand U24048 (N_24048,N_15423,N_19102);
or U24049 (N_24049,N_15124,N_17852);
xnor U24050 (N_24050,N_15951,N_16845);
and U24051 (N_24051,N_15857,N_15196);
and U24052 (N_24052,N_19447,N_15526);
nand U24053 (N_24053,N_17265,N_15474);
nor U24054 (N_24054,N_18400,N_16411);
and U24055 (N_24055,N_16051,N_19174);
and U24056 (N_24056,N_17095,N_16533);
nor U24057 (N_24057,N_16088,N_15781);
nand U24058 (N_24058,N_16354,N_19563);
or U24059 (N_24059,N_16773,N_17728);
nor U24060 (N_24060,N_19710,N_18594);
nand U24061 (N_24061,N_17681,N_15106);
nand U24062 (N_24062,N_17535,N_19836);
nor U24063 (N_24063,N_16020,N_18395);
or U24064 (N_24064,N_16112,N_15836);
xor U24065 (N_24065,N_16473,N_19430);
nand U24066 (N_24066,N_16514,N_19582);
nand U24067 (N_24067,N_15378,N_17718);
or U24068 (N_24068,N_18398,N_15897);
nand U24069 (N_24069,N_17242,N_17027);
or U24070 (N_24070,N_17134,N_17586);
xor U24071 (N_24071,N_19818,N_19191);
nand U24072 (N_24072,N_17322,N_19073);
xnor U24073 (N_24073,N_17358,N_18421);
xor U24074 (N_24074,N_18873,N_16600);
or U24075 (N_24075,N_18606,N_19726);
xnor U24076 (N_24076,N_16103,N_15352);
nor U24077 (N_24077,N_15716,N_15805);
xnor U24078 (N_24078,N_18086,N_17736);
and U24079 (N_24079,N_19578,N_17580);
nand U24080 (N_24080,N_16682,N_19059);
nand U24081 (N_24081,N_19533,N_15922);
or U24082 (N_24082,N_17038,N_16446);
or U24083 (N_24083,N_16607,N_15842);
nor U24084 (N_24084,N_19553,N_18711);
nand U24085 (N_24085,N_15983,N_16795);
nand U24086 (N_24086,N_16349,N_15613);
nor U24087 (N_24087,N_17945,N_17044);
xor U24088 (N_24088,N_17257,N_16714);
nand U24089 (N_24089,N_17587,N_17105);
nand U24090 (N_24090,N_19774,N_16621);
and U24091 (N_24091,N_17698,N_18545);
nor U24092 (N_24092,N_18484,N_18661);
nand U24093 (N_24093,N_15814,N_17831);
and U24094 (N_24094,N_19720,N_16769);
and U24095 (N_24095,N_16779,N_17635);
and U24096 (N_24096,N_18866,N_16366);
nor U24097 (N_24097,N_15434,N_18641);
or U24098 (N_24098,N_18254,N_15113);
xor U24099 (N_24099,N_17078,N_17275);
xnor U24100 (N_24100,N_15565,N_16662);
nor U24101 (N_24101,N_16035,N_15295);
or U24102 (N_24102,N_15076,N_15784);
xnor U24103 (N_24103,N_18096,N_17346);
nand U24104 (N_24104,N_19718,N_19662);
or U24105 (N_24105,N_19844,N_18718);
and U24106 (N_24106,N_15773,N_18482);
xnor U24107 (N_24107,N_19415,N_15153);
nor U24108 (N_24108,N_18032,N_17587);
nand U24109 (N_24109,N_17367,N_15105);
and U24110 (N_24110,N_15528,N_19707);
or U24111 (N_24111,N_19399,N_16794);
nand U24112 (N_24112,N_19412,N_18446);
nor U24113 (N_24113,N_18193,N_19705);
nand U24114 (N_24114,N_16755,N_19465);
nor U24115 (N_24115,N_17971,N_17473);
xnor U24116 (N_24116,N_15839,N_17245);
or U24117 (N_24117,N_19719,N_18961);
or U24118 (N_24118,N_18011,N_17421);
or U24119 (N_24119,N_19688,N_18019);
or U24120 (N_24120,N_17638,N_17554);
nor U24121 (N_24121,N_16015,N_18783);
or U24122 (N_24122,N_16575,N_18237);
nor U24123 (N_24123,N_18418,N_16736);
or U24124 (N_24124,N_17851,N_19910);
and U24125 (N_24125,N_19411,N_16730);
or U24126 (N_24126,N_15087,N_18563);
nand U24127 (N_24127,N_18878,N_15948);
or U24128 (N_24128,N_16737,N_15910);
or U24129 (N_24129,N_18400,N_18495);
nor U24130 (N_24130,N_16130,N_18228);
nor U24131 (N_24131,N_15829,N_17209);
nand U24132 (N_24132,N_15385,N_16016);
and U24133 (N_24133,N_17302,N_18185);
and U24134 (N_24134,N_18614,N_19713);
and U24135 (N_24135,N_16581,N_15154);
or U24136 (N_24136,N_15752,N_19668);
and U24137 (N_24137,N_15091,N_17955);
nand U24138 (N_24138,N_19937,N_18552);
nor U24139 (N_24139,N_19382,N_16827);
xor U24140 (N_24140,N_19284,N_16897);
nor U24141 (N_24141,N_17965,N_17404);
and U24142 (N_24142,N_19356,N_18212);
nand U24143 (N_24143,N_15561,N_16616);
nand U24144 (N_24144,N_18588,N_19382);
or U24145 (N_24145,N_19885,N_19744);
or U24146 (N_24146,N_19982,N_16094);
nand U24147 (N_24147,N_15535,N_16664);
nand U24148 (N_24148,N_18375,N_17037);
and U24149 (N_24149,N_17500,N_18407);
and U24150 (N_24150,N_19018,N_15280);
and U24151 (N_24151,N_17988,N_19398);
and U24152 (N_24152,N_19932,N_18114);
nor U24153 (N_24153,N_15674,N_16094);
or U24154 (N_24154,N_15690,N_15967);
nor U24155 (N_24155,N_15214,N_15845);
or U24156 (N_24156,N_15332,N_15424);
nand U24157 (N_24157,N_17622,N_19156);
or U24158 (N_24158,N_15395,N_17578);
xor U24159 (N_24159,N_18360,N_17122);
or U24160 (N_24160,N_17317,N_17600);
or U24161 (N_24161,N_17561,N_15725);
and U24162 (N_24162,N_16809,N_15214);
xor U24163 (N_24163,N_19758,N_16887);
or U24164 (N_24164,N_19315,N_18414);
or U24165 (N_24165,N_18240,N_16610);
nor U24166 (N_24166,N_17760,N_16989);
xnor U24167 (N_24167,N_18251,N_18818);
nand U24168 (N_24168,N_17631,N_15075);
nor U24169 (N_24169,N_19456,N_18171);
xnor U24170 (N_24170,N_16745,N_15651);
or U24171 (N_24171,N_18009,N_15874);
nand U24172 (N_24172,N_19987,N_19364);
or U24173 (N_24173,N_16289,N_18820);
xor U24174 (N_24174,N_19389,N_19353);
and U24175 (N_24175,N_18369,N_16661);
nand U24176 (N_24176,N_17784,N_16222);
and U24177 (N_24177,N_16686,N_15026);
xnor U24178 (N_24178,N_15936,N_17857);
nand U24179 (N_24179,N_17949,N_19416);
xnor U24180 (N_24180,N_19845,N_19807);
xnor U24181 (N_24181,N_15508,N_16868);
nor U24182 (N_24182,N_16019,N_19825);
nor U24183 (N_24183,N_16129,N_19683);
or U24184 (N_24184,N_18524,N_17812);
or U24185 (N_24185,N_19687,N_19050);
nor U24186 (N_24186,N_15209,N_17852);
xnor U24187 (N_24187,N_15842,N_16439);
nand U24188 (N_24188,N_19513,N_17787);
nor U24189 (N_24189,N_17847,N_16354);
xor U24190 (N_24190,N_15054,N_19192);
or U24191 (N_24191,N_19719,N_16428);
nand U24192 (N_24192,N_19955,N_15953);
or U24193 (N_24193,N_15366,N_19698);
or U24194 (N_24194,N_16683,N_17074);
xnor U24195 (N_24195,N_18309,N_17267);
nor U24196 (N_24196,N_19357,N_15216);
xnor U24197 (N_24197,N_16288,N_17950);
xor U24198 (N_24198,N_19300,N_17647);
nand U24199 (N_24199,N_17488,N_16247);
xnor U24200 (N_24200,N_15917,N_17842);
or U24201 (N_24201,N_19949,N_15586);
nand U24202 (N_24202,N_18070,N_16995);
nand U24203 (N_24203,N_19565,N_15231);
or U24204 (N_24204,N_15358,N_15549);
or U24205 (N_24205,N_15071,N_19388);
xnor U24206 (N_24206,N_17119,N_17960);
and U24207 (N_24207,N_19153,N_15975);
or U24208 (N_24208,N_18280,N_15828);
nand U24209 (N_24209,N_17499,N_16676);
or U24210 (N_24210,N_18192,N_19158);
or U24211 (N_24211,N_17113,N_15158);
nor U24212 (N_24212,N_19467,N_16217);
nor U24213 (N_24213,N_15959,N_16256);
and U24214 (N_24214,N_19416,N_15380);
nand U24215 (N_24215,N_19885,N_17115);
nor U24216 (N_24216,N_17512,N_19370);
nand U24217 (N_24217,N_17225,N_16552);
nand U24218 (N_24218,N_15971,N_18129);
xor U24219 (N_24219,N_18020,N_17610);
xor U24220 (N_24220,N_19176,N_16871);
and U24221 (N_24221,N_16146,N_18349);
or U24222 (N_24222,N_19564,N_16560);
and U24223 (N_24223,N_16916,N_19360);
nand U24224 (N_24224,N_17974,N_15067);
nor U24225 (N_24225,N_17456,N_15668);
nor U24226 (N_24226,N_17657,N_15626);
and U24227 (N_24227,N_16869,N_18418);
and U24228 (N_24228,N_16922,N_15442);
and U24229 (N_24229,N_17990,N_18443);
and U24230 (N_24230,N_19997,N_16209);
nand U24231 (N_24231,N_19555,N_18135);
or U24232 (N_24232,N_17489,N_19611);
nor U24233 (N_24233,N_18965,N_18629);
nor U24234 (N_24234,N_17026,N_17435);
or U24235 (N_24235,N_19387,N_18572);
xnor U24236 (N_24236,N_15727,N_15793);
and U24237 (N_24237,N_17573,N_19635);
or U24238 (N_24238,N_16434,N_19503);
and U24239 (N_24239,N_17545,N_15192);
xor U24240 (N_24240,N_17136,N_18191);
nand U24241 (N_24241,N_16352,N_15615);
nand U24242 (N_24242,N_16472,N_18839);
xnor U24243 (N_24243,N_15537,N_19097);
xnor U24244 (N_24244,N_15530,N_17264);
and U24245 (N_24245,N_18771,N_18690);
or U24246 (N_24246,N_15438,N_17610);
nor U24247 (N_24247,N_18960,N_15403);
nand U24248 (N_24248,N_17263,N_16543);
xor U24249 (N_24249,N_18773,N_18136);
nand U24250 (N_24250,N_17396,N_18690);
nor U24251 (N_24251,N_16758,N_18675);
xor U24252 (N_24252,N_19564,N_19430);
or U24253 (N_24253,N_16996,N_15678);
nand U24254 (N_24254,N_18656,N_19466);
nor U24255 (N_24255,N_15311,N_15666);
nor U24256 (N_24256,N_18459,N_16661);
nand U24257 (N_24257,N_18471,N_17996);
xor U24258 (N_24258,N_17192,N_15711);
nand U24259 (N_24259,N_19849,N_15490);
nor U24260 (N_24260,N_15311,N_15115);
and U24261 (N_24261,N_19759,N_18112);
nand U24262 (N_24262,N_19159,N_18855);
or U24263 (N_24263,N_16885,N_17575);
and U24264 (N_24264,N_16705,N_18366);
and U24265 (N_24265,N_16465,N_17864);
nor U24266 (N_24266,N_19467,N_17509);
xor U24267 (N_24267,N_16052,N_16939);
and U24268 (N_24268,N_17118,N_16893);
or U24269 (N_24269,N_15347,N_18244);
xnor U24270 (N_24270,N_19902,N_17134);
xor U24271 (N_24271,N_18307,N_18083);
xor U24272 (N_24272,N_15138,N_15743);
nand U24273 (N_24273,N_19870,N_18169);
nor U24274 (N_24274,N_15936,N_17027);
and U24275 (N_24275,N_19494,N_16210);
or U24276 (N_24276,N_18729,N_18171);
xor U24277 (N_24277,N_19043,N_15000);
nor U24278 (N_24278,N_16503,N_16817);
or U24279 (N_24279,N_15085,N_18361);
xor U24280 (N_24280,N_17560,N_19229);
xnor U24281 (N_24281,N_17889,N_18244);
and U24282 (N_24282,N_19095,N_16985);
and U24283 (N_24283,N_18001,N_19418);
or U24284 (N_24284,N_18124,N_16365);
and U24285 (N_24285,N_19186,N_18353);
nor U24286 (N_24286,N_18311,N_19526);
xor U24287 (N_24287,N_18722,N_16955);
nor U24288 (N_24288,N_17176,N_19544);
xnor U24289 (N_24289,N_19790,N_17072);
and U24290 (N_24290,N_19515,N_18786);
or U24291 (N_24291,N_16809,N_17558);
xor U24292 (N_24292,N_15150,N_15301);
nand U24293 (N_24293,N_17420,N_17389);
xnor U24294 (N_24294,N_19938,N_19912);
xor U24295 (N_24295,N_17616,N_16669);
nor U24296 (N_24296,N_18809,N_17791);
nor U24297 (N_24297,N_18483,N_16370);
nor U24298 (N_24298,N_18899,N_19087);
or U24299 (N_24299,N_17148,N_19256);
or U24300 (N_24300,N_15026,N_16833);
and U24301 (N_24301,N_19146,N_19544);
nand U24302 (N_24302,N_17862,N_16969);
and U24303 (N_24303,N_17051,N_18827);
and U24304 (N_24304,N_15809,N_15527);
nor U24305 (N_24305,N_15045,N_19626);
nand U24306 (N_24306,N_16795,N_16613);
nand U24307 (N_24307,N_16953,N_18322);
nand U24308 (N_24308,N_19063,N_16616);
or U24309 (N_24309,N_15252,N_16881);
and U24310 (N_24310,N_19026,N_18355);
nand U24311 (N_24311,N_16303,N_16445);
xor U24312 (N_24312,N_18136,N_16873);
and U24313 (N_24313,N_19255,N_16951);
or U24314 (N_24314,N_17113,N_15556);
nand U24315 (N_24315,N_17050,N_18545);
nand U24316 (N_24316,N_18371,N_18820);
nand U24317 (N_24317,N_19325,N_16162);
xnor U24318 (N_24318,N_15323,N_17917);
or U24319 (N_24319,N_17368,N_15724);
and U24320 (N_24320,N_18713,N_15147);
nand U24321 (N_24321,N_17305,N_15185);
or U24322 (N_24322,N_18564,N_19087);
nor U24323 (N_24323,N_19428,N_17282);
xor U24324 (N_24324,N_19191,N_15372);
or U24325 (N_24325,N_19871,N_17600);
nor U24326 (N_24326,N_15859,N_19441);
nand U24327 (N_24327,N_19326,N_19942);
and U24328 (N_24328,N_17327,N_15792);
nor U24329 (N_24329,N_18799,N_19221);
or U24330 (N_24330,N_18932,N_17282);
and U24331 (N_24331,N_19464,N_18042);
xnor U24332 (N_24332,N_18648,N_15926);
and U24333 (N_24333,N_15909,N_16124);
xor U24334 (N_24334,N_17942,N_19153);
xnor U24335 (N_24335,N_17503,N_15812);
xor U24336 (N_24336,N_17999,N_19500);
and U24337 (N_24337,N_15883,N_15661);
xor U24338 (N_24338,N_17264,N_15503);
xnor U24339 (N_24339,N_17293,N_17331);
and U24340 (N_24340,N_19924,N_19326);
xor U24341 (N_24341,N_19600,N_16801);
nor U24342 (N_24342,N_17964,N_15928);
nor U24343 (N_24343,N_18820,N_17318);
and U24344 (N_24344,N_17679,N_15300);
nand U24345 (N_24345,N_17811,N_17478);
and U24346 (N_24346,N_19413,N_16027);
nand U24347 (N_24347,N_16087,N_18567);
nand U24348 (N_24348,N_16711,N_17822);
or U24349 (N_24349,N_17629,N_19587);
xnor U24350 (N_24350,N_18628,N_18865);
nor U24351 (N_24351,N_15123,N_18592);
and U24352 (N_24352,N_17583,N_15698);
xor U24353 (N_24353,N_18906,N_16953);
nor U24354 (N_24354,N_16393,N_17336);
or U24355 (N_24355,N_17895,N_16127);
and U24356 (N_24356,N_18423,N_19113);
nand U24357 (N_24357,N_16596,N_16122);
nand U24358 (N_24358,N_17387,N_15000);
or U24359 (N_24359,N_15023,N_16941);
and U24360 (N_24360,N_16060,N_18500);
or U24361 (N_24361,N_15061,N_15084);
nand U24362 (N_24362,N_18902,N_15304);
nor U24363 (N_24363,N_15378,N_16805);
nand U24364 (N_24364,N_15179,N_16082);
nand U24365 (N_24365,N_19351,N_15029);
or U24366 (N_24366,N_15489,N_16646);
and U24367 (N_24367,N_15308,N_19767);
and U24368 (N_24368,N_16321,N_16493);
xnor U24369 (N_24369,N_16088,N_15008);
nand U24370 (N_24370,N_17497,N_17082);
and U24371 (N_24371,N_19358,N_18923);
and U24372 (N_24372,N_17269,N_15407);
xor U24373 (N_24373,N_15049,N_15065);
nand U24374 (N_24374,N_18706,N_16811);
and U24375 (N_24375,N_18397,N_19834);
nor U24376 (N_24376,N_16848,N_19012);
and U24377 (N_24377,N_19774,N_19875);
nor U24378 (N_24378,N_15916,N_18844);
and U24379 (N_24379,N_17741,N_17353);
nand U24380 (N_24380,N_17864,N_18733);
or U24381 (N_24381,N_16986,N_18745);
xor U24382 (N_24382,N_17057,N_19503);
nor U24383 (N_24383,N_19571,N_19897);
xnor U24384 (N_24384,N_16738,N_18968);
nor U24385 (N_24385,N_15002,N_18946);
nand U24386 (N_24386,N_15906,N_15829);
or U24387 (N_24387,N_15692,N_18771);
nor U24388 (N_24388,N_19151,N_19479);
or U24389 (N_24389,N_19213,N_19596);
nor U24390 (N_24390,N_15183,N_19291);
xnor U24391 (N_24391,N_19354,N_18646);
xnor U24392 (N_24392,N_18551,N_15677);
nor U24393 (N_24393,N_18603,N_16125);
xor U24394 (N_24394,N_15264,N_18488);
xor U24395 (N_24395,N_15704,N_15479);
nand U24396 (N_24396,N_17725,N_16341);
nand U24397 (N_24397,N_19125,N_17814);
nor U24398 (N_24398,N_17757,N_16347);
nor U24399 (N_24399,N_15066,N_16205);
or U24400 (N_24400,N_15905,N_17164);
nor U24401 (N_24401,N_18998,N_18303);
nand U24402 (N_24402,N_18196,N_17549);
xor U24403 (N_24403,N_18049,N_17567);
xnor U24404 (N_24404,N_16656,N_17554);
nand U24405 (N_24405,N_16394,N_17878);
and U24406 (N_24406,N_19764,N_18217);
and U24407 (N_24407,N_16876,N_18819);
nor U24408 (N_24408,N_15554,N_17129);
and U24409 (N_24409,N_16385,N_19605);
xor U24410 (N_24410,N_16428,N_16494);
and U24411 (N_24411,N_15849,N_19676);
nand U24412 (N_24412,N_16416,N_17334);
and U24413 (N_24413,N_16515,N_16741);
nand U24414 (N_24414,N_19728,N_19775);
nor U24415 (N_24415,N_15177,N_15747);
nand U24416 (N_24416,N_18565,N_15005);
or U24417 (N_24417,N_18282,N_16878);
and U24418 (N_24418,N_19545,N_18563);
or U24419 (N_24419,N_16646,N_19255);
xnor U24420 (N_24420,N_19910,N_19321);
and U24421 (N_24421,N_15570,N_19530);
xor U24422 (N_24422,N_18435,N_16759);
xor U24423 (N_24423,N_19961,N_16326);
nand U24424 (N_24424,N_16387,N_18314);
nor U24425 (N_24425,N_18229,N_18079);
nand U24426 (N_24426,N_19994,N_16105);
or U24427 (N_24427,N_15949,N_19810);
or U24428 (N_24428,N_18584,N_18537);
and U24429 (N_24429,N_17980,N_18691);
nor U24430 (N_24430,N_15884,N_18968);
xor U24431 (N_24431,N_17662,N_19945);
nor U24432 (N_24432,N_16981,N_18833);
nor U24433 (N_24433,N_18926,N_15756);
nand U24434 (N_24434,N_16909,N_15704);
and U24435 (N_24435,N_16834,N_15652);
or U24436 (N_24436,N_15710,N_15168);
xor U24437 (N_24437,N_16576,N_18987);
nand U24438 (N_24438,N_16421,N_16336);
nor U24439 (N_24439,N_15228,N_19570);
and U24440 (N_24440,N_18633,N_17629);
nor U24441 (N_24441,N_15295,N_15851);
nor U24442 (N_24442,N_16753,N_16708);
nor U24443 (N_24443,N_16874,N_16326);
or U24444 (N_24444,N_16578,N_15232);
or U24445 (N_24445,N_15836,N_15595);
nor U24446 (N_24446,N_15897,N_15948);
or U24447 (N_24447,N_17399,N_15346);
nor U24448 (N_24448,N_18115,N_17452);
nor U24449 (N_24449,N_19657,N_17131);
nor U24450 (N_24450,N_15107,N_16818);
xnor U24451 (N_24451,N_15326,N_19212);
nand U24452 (N_24452,N_15399,N_15141);
xnor U24453 (N_24453,N_17712,N_17864);
or U24454 (N_24454,N_18746,N_15355);
or U24455 (N_24455,N_16974,N_19151);
nand U24456 (N_24456,N_16011,N_16757);
and U24457 (N_24457,N_15512,N_17725);
nand U24458 (N_24458,N_19736,N_16133);
xnor U24459 (N_24459,N_18669,N_15538);
xnor U24460 (N_24460,N_17310,N_17284);
xor U24461 (N_24461,N_17245,N_15189);
nand U24462 (N_24462,N_16212,N_17972);
nor U24463 (N_24463,N_18016,N_15132);
and U24464 (N_24464,N_17957,N_19962);
and U24465 (N_24465,N_15218,N_17131);
or U24466 (N_24466,N_15489,N_18752);
nand U24467 (N_24467,N_15946,N_17198);
and U24468 (N_24468,N_18922,N_19268);
nand U24469 (N_24469,N_16633,N_18790);
nand U24470 (N_24470,N_15591,N_16308);
nor U24471 (N_24471,N_15276,N_17011);
nor U24472 (N_24472,N_17918,N_19283);
xnor U24473 (N_24473,N_19115,N_15772);
xnor U24474 (N_24474,N_15615,N_17119);
or U24475 (N_24475,N_19717,N_19243);
or U24476 (N_24476,N_15862,N_17964);
or U24477 (N_24477,N_15995,N_17350);
xnor U24478 (N_24478,N_19830,N_19599);
nor U24479 (N_24479,N_18772,N_19525);
and U24480 (N_24480,N_16716,N_15506);
nand U24481 (N_24481,N_16198,N_18363);
and U24482 (N_24482,N_18425,N_17315);
xnor U24483 (N_24483,N_15258,N_18866);
xnor U24484 (N_24484,N_15632,N_16698);
or U24485 (N_24485,N_18955,N_16745);
and U24486 (N_24486,N_15438,N_16484);
or U24487 (N_24487,N_17643,N_15300);
and U24488 (N_24488,N_18052,N_15811);
and U24489 (N_24489,N_17706,N_15654);
and U24490 (N_24490,N_15910,N_17502);
nand U24491 (N_24491,N_18324,N_15826);
or U24492 (N_24492,N_18829,N_18802);
and U24493 (N_24493,N_18668,N_15698);
and U24494 (N_24494,N_15799,N_15154);
or U24495 (N_24495,N_18755,N_15330);
xor U24496 (N_24496,N_19789,N_19458);
nand U24497 (N_24497,N_18022,N_17853);
and U24498 (N_24498,N_17058,N_17637);
and U24499 (N_24499,N_15214,N_15410);
and U24500 (N_24500,N_16252,N_19117);
xor U24501 (N_24501,N_18873,N_19917);
and U24502 (N_24502,N_16772,N_19007);
nor U24503 (N_24503,N_16774,N_15484);
nand U24504 (N_24504,N_15414,N_15473);
nand U24505 (N_24505,N_19805,N_19478);
and U24506 (N_24506,N_18471,N_19134);
and U24507 (N_24507,N_16516,N_18697);
nand U24508 (N_24508,N_18829,N_16373);
nor U24509 (N_24509,N_15140,N_15671);
and U24510 (N_24510,N_15810,N_18860);
and U24511 (N_24511,N_16466,N_19617);
and U24512 (N_24512,N_18881,N_18224);
nand U24513 (N_24513,N_16911,N_16984);
xor U24514 (N_24514,N_16429,N_19702);
or U24515 (N_24515,N_15135,N_18565);
and U24516 (N_24516,N_17357,N_16224);
and U24517 (N_24517,N_15190,N_18694);
or U24518 (N_24518,N_19059,N_15981);
nand U24519 (N_24519,N_16000,N_18386);
or U24520 (N_24520,N_17042,N_16594);
xor U24521 (N_24521,N_17337,N_17431);
or U24522 (N_24522,N_18778,N_18593);
and U24523 (N_24523,N_15598,N_15367);
or U24524 (N_24524,N_16465,N_16631);
nand U24525 (N_24525,N_16653,N_16770);
and U24526 (N_24526,N_18358,N_15533);
nor U24527 (N_24527,N_18186,N_15143);
and U24528 (N_24528,N_18437,N_17788);
xnor U24529 (N_24529,N_17534,N_17464);
xor U24530 (N_24530,N_19745,N_19783);
xor U24531 (N_24531,N_17836,N_16872);
xnor U24532 (N_24532,N_17714,N_19703);
nor U24533 (N_24533,N_16152,N_15440);
and U24534 (N_24534,N_16994,N_17605);
nor U24535 (N_24535,N_16579,N_16639);
nand U24536 (N_24536,N_18660,N_15814);
nor U24537 (N_24537,N_17441,N_16441);
nand U24538 (N_24538,N_18435,N_19772);
nand U24539 (N_24539,N_19545,N_16228);
xnor U24540 (N_24540,N_15031,N_15532);
nor U24541 (N_24541,N_19025,N_16155);
or U24542 (N_24542,N_17677,N_17779);
xnor U24543 (N_24543,N_16565,N_16289);
nor U24544 (N_24544,N_17416,N_16914);
and U24545 (N_24545,N_17255,N_17975);
nand U24546 (N_24546,N_15748,N_18639);
nor U24547 (N_24547,N_18833,N_18775);
nand U24548 (N_24548,N_18717,N_15487);
and U24549 (N_24549,N_16374,N_18837);
nor U24550 (N_24550,N_15155,N_18197);
xor U24551 (N_24551,N_15269,N_16565);
nor U24552 (N_24552,N_15969,N_18558);
nand U24553 (N_24553,N_17421,N_18866);
and U24554 (N_24554,N_15080,N_17210);
or U24555 (N_24555,N_17733,N_15427);
nor U24556 (N_24556,N_17576,N_19714);
xnor U24557 (N_24557,N_15034,N_18708);
and U24558 (N_24558,N_15336,N_16549);
and U24559 (N_24559,N_19640,N_18783);
and U24560 (N_24560,N_15688,N_19800);
or U24561 (N_24561,N_15652,N_17164);
xor U24562 (N_24562,N_16817,N_16209);
nor U24563 (N_24563,N_15190,N_19746);
xnor U24564 (N_24564,N_17457,N_17094);
nand U24565 (N_24565,N_18366,N_15296);
nor U24566 (N_24566,N_17622,N_17459);
or U24567 (N_24567,N_19982,N_17753);
and U24568 (N_24568,N_18288,N_19090);
nor U24569 (N_24569,N_19236,N_15720);
and U24570 (N_24570,N_19715,N_19681);
or U24571 (N_24571,N_15809,N_19827);
nand U24572 (N_24572,N_15555,N_15805);
and U24573 (N_24573,N_15437,N_16542);
nor U24574 (N_24574,N_19159,N_15597);
nor U24575 (N_24575,N_15711,N_18637);
or U24576 (N_24576,N_17308,N_16314);
nor U24577 (N_24577,N_18647,N_19466);
and U24578 (N_24578,N_19500,N_18467);
or U24579 (N_24579,N_16079,N_16973);
nand U24580 (N_24580,N_15561,N_18210);
or U24581 (N_24581,N_17278,N_18900);
nand U24582 (N_24582,N_16823,N_16236);
xnor U24583 (N_24583,N_16113,N_18587);
xor U24584 (N_24584,N_17197,N_15371);
nand U24585 (N_24585,N_16245,N_16344);
or U24586 (N_24586,N_19635,N_16655);
and U24587 (N_24587,N_15314,N_16834);
nor U24588 (N_24588,N_18681,N_16680);
xor U24589 (N_24589,N_15692,N_16755);
or U24590 (N_24590,N_16272,N_19774);
or U24591 (N_24591,N_16124,N_17466);
nor U24592 (N_24592,N_17431,N_17600);
nor U24593 (N_24593,N_16905,N_19929);
nand U24594 (N_24594,N_15428,N_15621);
xor U24595 (N_24595,N_16398,N_18628);
and U24596 (N_24596,N_17112,N_16177);
or U24597 (N_24597,N_19955,N_15912);
nand U24598 (N_24598,N_19102,N_15352);
or U24599 (N_24599,N_15419,N_17298);
nor U24600 (N_24600,N_16943,N_17447);
nand U24601 (N_24601,N_16648,N_18412);
xnor U24602 (N_24602,N_17316,N_17098);
or U24603 (N_24603,N_18570,N_19759);
nor U24604 (N_24604,N_15345,N_19316);
nand U24605 (N_24605,N_16703,N_15884);
or U24606 (N_24606,N_16922,N_15612);
nor U24607 (N_24607,N_19888,N_18887);
nor U24608 (N_24608,N_15529,N_16334);
nor U24609 (N_24609,N_19277,N_16135);
or U24610 (N_24610,N_17782,N_16564);
and U24611 (N_24611,N_17368,N_17387);
and U24612 (N_24612,N_17583,N_19000);
nor U24613 (N_24613,N_18488,N_17462);
and U24614 (N_24614,N_16377,N_17601);
nor U24615 (N_24615,N_18536,N_18772);
xnor U24616 (N_24616,N_18183,N_16880);
or U24617 (N_24617,N_17112,N_18780);
nand U24618 (N_24618,N_16217,N_16801);
and U24619 (N_24619,N_17549,N_15549);
and U24620 (N_24620,N_16186,N_15353);
nor U24621 (N_24621,N_17019,N_19838);
nor U24622 (N_24622,N_17492,N_17888);
and U24623 (N_24623,N_16691,N_17131);
nand U24624 (N_24624,N_15455,N_16622);
nand U24625 (N_24625,N_16871,N_16343);
nor U24626 (N_24626,N_18250,N_15176);
xnor U24627 (N_24627,N_18080,N_19374);
nor U24628 (N_24628,N_18430,N_18148);
and U24629 (N_24629,N_19868,N_16595);
nor U24630 (N_24630,N_15881,N_15319);
and U24631 (N_24631,N_16692,N_16059);
nand U24632 (N_24632,N_19313,N_17259);
xor U24633 (N_24633,N_19754,N_17437);
nand U24634 (N_24634,N_17292,N_15148);
nor U24635 (N_24635,N_17361,N_19883);
or U24636 (N_24636,N_16194,N_16640);
nor U24637 (N_24637,N_17598,N_16889);
nor U24638 (N_24638,N_15660,N_16130);
nor U24639 (N_24639,N_15598,N_18091);
and U24640 (N_24640,N_18299,N_19402);
or U24641 (N_24641,N_17555,N_18235);
xor U24642 (N_24642,N_19716,N_15826);
nand U24643 (N_24643,N_19701,N_16910);
nor U24644 (N_24644,N_19038,N_15590);
and U24645 (N_24645,N_16642,N_15064);
and U24646 (N_24646,N_16310,N_16947);
or U24647 (N_24647,N_15494,N_15520);
nor U24648 (N_24648,N_18475,N_18785);
nor U24649 (N_24649,N_19385,N_15351);
nor U24650 (N_24650,N_16105,N_17972);
xor U24651 (N_24651,N_16831,N_15307);
or U24652 (N_24652,N_18433,N_17688);
nor U24653 (N_24653,N_16583,N_16082);
nor U24654 (N_24654,N_16351,N_19468);
nand U24655 (N_24655,N_16565,N_17000);
or U24656 (N_24656,N_17756,N_15036);
and U24657 (N_24657,N_16780,N_16716);
nand U24658 (N_24658,N_15392,N_18936);
xnor U24659 (N_24659,N_19679,N_16341);
nand U24660 (N_24660,N_19147,N_19612);
nand U24661 (N_24661,N_17652,N_15450);
xor U24662 (N_24662,N_17847,N_16635);
nor U24663 (N_24663,N_15461,N_19472);
xor U24664 (N_24664,N_15075,N_19810);
and U24665 (N_24665,N_17658,N_19644);
xnor U24666 (N_24666,N_17172,N_15606);
or U24667 (N_24667,N_17762,N_17423);
and U24668 (N_24668,N_18119,N_18335);
nand U24669 (N_24669,N_16141,N_17509);
or U24670 (N_24670,N_15367,N_17534);
xnor U24671 (N_24671,N_18156,N_19669);
and U24672 (N_24672,N_15229,N_19876);
nor U24673 (N_24673,N_15238,N_15740);
or U24674 (N_24674,N_16137,N_17076);
nor U24675 (N_24675,N_17432,N_17777);
and U24676 (N_24676,N_15604,N_19777);
or U24677 (N_24677,N_17961,N_16972);
nand U24678 (N_24678,N_17442,N_16621);
and U24679 (N_24679,N_16502,N_15772);
or U24680 (N_24680,N_17840,N_17562);
nor U24681 (N_24681,N_19639,N_16441);
xnor U24682 (N_24682,N_19355,N_18879);
and U24683 (N_24683,N_16829,N_18856);
and U24684 (N_24684,N_16864,N_15297);
xnor U24685 (N_24685,N_18194,N_15765);
nor U24686 (N_24686,N_18679,N_15326);
nor U24687 (N_24687,N_15103,N_17634);
nor U24688 (N_24688,N_15126,N_16462);
nand U24689 (N_24689,N_18075,N_19215);
nand U24690 (N_24690,N_16047,N_18062);
xor U24691 (N_24691,N_15842,N_15896);
nor U24692 (N_24692,N_19078,N_15736);
or U24693 (N_24693,N_16906,N_18091);
nand U24694 (N_24694,N_16417,N_16154);
or U24695 (N_24695,N_17740,N_18849);
nor U24696 (N_24696,N_15001,N_17806);
and U24697 (N_24697,N_15845,N_15805);
nor U24698 (N_24698,N_15290,N_17005);
or U24699 (N_24699,N_16359,N_17914);
nor U24700 (N_24700,N_19895,N_16542);
nor U24701 (N_24701,N_19044,N_16327);
xnor U24702 (N_24702,N_18533,N_15836);
and U24703 (N_24703,N_18383,N_17711);
and U24704 (N_24704,N_17093,N_19327);
nor U24705 (N_24705,N_17779,N_17156);
and U24706 (N_24706,N_16730,N_18173);
or U24707 (N_24707,N_17787,N_19188);
and U24708 (N_24708,N_15274,N_17180);
and U24709 (N_24709,N_17771,N_18060);
xnor U24710 (N_24710,N_17041,N_17885);
nand U24711 (N_24711,N_19033,N_15977);
nand U24712 (N_24712,N_18376,N_17113);
xor U24713 (N_24713,N_16788,N_17701);
nand U24714 (N_24714,N_19999,N_18249);
nor U24715 (N_24715,N_15066,N_16965);
and U24716 (N_24716,N_17072,N_17438);
nand U24717 (N_24717,N_17593,N_17472);
and U24718 (N_24718,N_17453,N_18173);
nand U24719 (N_24719,N_17497,N_16145);
and U24720 (N_24720,N_17696,N_19947);
nor U24721 (N_24721,N_18047,N_18445);
xnor U24722 (N_24722,N_15078,N_17886);
nand U24723 (N_24723,N_17097,N_19559);
nand U24724 (N_24724,N_17427,N_19223);
nand U24725 (N_24725,N_16353,N_19919);
nand U24726 (N_24726,N_17469,N_19386);
nand U24727 (N_24727,N_15243,N_15000);
xor U24728 (N_24728,N_17218,N_17967);
xor U24729 (N_24729,N_16940,N_17669);
nor U24730 (N_24730,N_19825,N_15156);
nor U24731 (N_24731,N_19695,N_17108);
nor U24732 (N_24732,N_18061,N_19946);
xor U24733 (N_24733,N_18697,N_17712);
xnor U24734 (N_24734,N_16926,N_16075);
xor U24735 (N_24735,N_18419,N_16196);
or U24736 (N_24736,N_16664,N_15727);
nand U24737 (N_24737,N_18651,N_18940);
xor U24738 (N_24738,N_17607,N_19453);
or U24739 (N_24739,N_16084,N_17869);
and U24740 (N_24740,N_19074,N_19527);
nand U24741 (N_24741,N_15977,N_15230);
or U24742 (N_24742,N_16640,N_16070);
or U24743 (N_24743,N_15813,N_16035);
xnor U24744 (N_24744,N_18855,N_17432);
or U24745 (N_24745,N_17839,N_15822);
and U24746 (N_24746,N_15940,N_19845);
nor U24747 (N_24747,N_19457,N_16879);
xnor U24748 (N_24748,N_17478,N_17692);
nor U24749 (N_24749,N_16072,N_17679);
or U24750 (N_24750,N_18374,N_17569);
xnor U24751 (N_24751,N_18038,N_19642);
xnor U24752 (N_24752,N_16449,N_19727);
nor U24753 (N_24753,N_19537,N_17790);
nor U24754 (N_24754,N_15437,N_16665);
nor U24755 (N_24755,N_16797,N_15297);
and U24756 (N_24756,N_17145,N_19131);
or U24757 (N_24757,N_17683,N_15582);
and U24758 (N_24758,N_18265,N_16107);
nor U24759 (N_24759,N_16653,N_17467);
xnor U24760 (N_24760,N_18176,N_18074);
nor U24761 (N_24761,N_17202,N_17581);
nor U24762 (N_24762,N_17744,N_17762);
xnor U24763 (N_24763,N_19029,N_19031);
xnor U24764 (N_24764,N_16575,N_18739);
and U24765 (N_24765,N_16681,N_18278);
and U24766 (N_24766,N_16897,N_16644);
and U24767 (N_24767,N_18324,N_17667);
and U24768 (N_24768,N_19395,N_15566);
nor U24769 (N_24769,N_15678,N_16447);
xnor U24770 (N_24770,N_19416,N_16711);
and U24771 (N_24771,N_15501,N_15660);
and U24772 (N_24772,N_15451,N_15331);
xnor U24773 (N_24773,N_16264,N_16465);
or U24774 (N_24774,N_19877,N_18460);
nor U24775 (N_24775,N_16401,N_16968);
and U24776 (N_24776,N_17581,N_15492);
nand U24777 (N_24777,N_16654,N_17190);
and U24778 (N_24778,N_17208,N_15461);
or U24779 (N_24779,N_17573,N_17404);
xor U24780 (N_24780,N_17613,N_18791);
or U24781 (N_24781,N_19562,N_19766);
and U24782 (N_24782,N_19475,N_15785);
and U24783 (N_24783,N_16225,N_18199);
nand U24784 (N_24784,N_16794,N_18394);
xnor U24785 (N_24785,N_19427,N_18068);
nor U24786 (N_24786,N_19900,N_18677);
and U24787 (N_24787,N_15408,N_19287);
xnor U24788 (N_24788,N_18696,N_17682);
or U24789 (N_24789,N_17555,N_15384);
or U24790 (N_24790,N_19298,N_18112);
nor U24791 (N_24791,N_19445,N_18539);
xor U24792 (N_24792,N_15377,N_16532);
or U24793 (N_24793,N_16682,N_16084);
or U24794 (N_24794,N_17649,N_16262);
nor U24795 (N_24795,N_18972,N_18095);
nor U24796 (N_24796,N_17748,N_19400);
nand U24797 (N_24797,N_19566,N_19557);
nor U24798 (N_24798,N_18274,N_18359);
and U24799 (N_24799,N_16823,N_19888);
nand U24800 (N_24800,N_16367,N_15916);
and U24801 (N_24801,N_17298,N_16225);
or U24802 (N_24802,N_15335,N_15014);
nand U24803 (N_24803,N_16670,N_18905);
nand U24804 (N_24804,N_16191,N_16933);
and U24805 (N_24805,N_17323,N_19181);
nand U24806 (N_24806,N_16867,N_19876);
nand U24807 (N_24807,N_19335,N_18145);
xor U24808 (N_24808,N_18735,N_18132);
nand U24809 (N_24809,N_18900,N_17611);
xnor U24810 (N_24810,N_16075,N_15174);
and U24811 (N_24811,N_17426,N_18485);
nor U24812 (N_24812,N_18490,N_17946);
xnor U24813 (N_24813,N_18812,N_19040);
or U24814 (N_24814,N_18214,N_15919);
or U24815 (N_24815,N_19048,N_16199);
xor U24816 (N_24816,N_19013,N_18964);
nand U24817 (N_24817,N_19547,N_17217);
xor U24818 (N_24818,N_15993,N_19918);
xnor U24819 (N_24819,N_18895,N_18872);
and U24820 (N_24820,N_16866,N_17703);
xnor U24821 (N_24821,N_19782,N_15792);
and U24822 (N_24822,N_18702,N_17132);
nor U24823 (N_24823,N_15766,N_18958);
nor U24824 (N_24824,N_17120,N_16536);
and U24825 (N_24825,N_16391,N_16778);
and U24826 (N_24826,N_17876,N_17895);
nand U24827 (N_24827,N_16014,N_19023);
or U24828 (N_24828,N_19795,N_18641);
and U24829 (N_24829,N_16540,N_19501);
and U24830 (N_24830,N_18832,N_15778);
and U24831 (N_24831,N_15927,N_18105);
and U24832 (N_24832,N_15762,N_19658);
xor U24833 (N_24833,N_16030,N_15240);
xnor U24834 (N_24834,N_19667,N_19811);
nor U24835 (N_24835,N_17574,N_17215);
and U24836 (N_24836,N_17182,N_15763);
nand U24837 (N_24837,N_19186,N_16392);
xor U24838 (N_24838,N_15121,N_15631);
and U24839 (N_24839,N_17523,N_18358);
or U24840 (N_24840,N_19761,N_16378);
nand U24841 (N_24841,N_19002,N_17501);
xor U24842 (N_24842,N_18891,N_19278);
and U24843 (N_24843,N_17728,N_18602);
and U24844 (N_24844,N_17673,N_18708);
or U24845 (N_24845,N_18307,N_18540);
nor U24846 (N_24846,N_16083,N_16314);
or U24847 (N_24847,N_15153,N_17825);
or U24848 (N_24848,N_17034,N_15857);
nor U24849 (N_24849,N_17941,N_19818);
and U24850 (N_24850,N_15819,N_15924);
or U24851 (N_24851,N_18064,N_17072);
nand U24852 (N_24852,N_16823,N_16658);
xor U24853 (N_24853,N_16805,N_15808);
and U24854 (N_24854,N_16461,N_16084);
nand U24855 (N_24855,N_19264,N_16483);
nor U24856 (N_24856,N_16294,N_19301);
xor U24857 (N_24857,N_15107,N_15614);
nor U24858 (N_24858,N_15906,N_17067);
xnor U24859 (N_24859,N_15132,N_15863);
xnor U24860 (N_24860,N_17334,N_15183);
nor U24861 (N_24861,N_16429,N_18490);
and U24862 (N_24862,N_19377,N_16337);
xnor U24863 (N_24863,N_18861,N_18582);
xnor U24864 (N_24864,N_18149,N_17947);
nor U24865 (N_24865,N_19452,N_18489);
nor U24866 (N_24866,N_16249,N_19378);
and U24867 (N_24867,N_16185,N_17188);
nand U24868 (N_24868,N_15608,N_18938);
nand U24869 (N_24869,N_17047,N_19137);
and U24870 (N_24870,N_19795,N_15890);
xnor U24871 (N_24871,N_19118,N_19327);
xnor U24872 (N_24872,N_17285,N_19433);
nor U24873 (N_24873,N_15914,N_15162);
and U24874 (N_24874,N_16608,N_15584);
and U24875 (N_24875,N_18190,N_18124);
nor U24876 (N_24876,N_16803,N_16323);
and U24877 (N_24877,N_19437,N_15473);
nand U24878 (N_24878,N_17162,N_15601);
nand U24879 (N_24879,N_15950,N_16345);
or U24880 (N_24880,N_18597,N_19801);
nand U24881 (N_24881,N_17149,N_18950);
and U24882 (N_24882,N_15009,N_18229);
or U24883 (N_24883,N_16684,N_15746);
xor U24884 (N_24884,N_19124,N_19779);
nor U24885 (N_24885,N_16272,N_16927);
nand U24886 (N_24886,N_16447,N_17895);
nor U24887 (N_24887,N_16126,N_19812);
nor U24888 (N_24888,N_18234,N_15424);
and U24889 (N_24889,N_17635,N_15767);
and U24890 (N_24890,N_17098,N_16385);
or U24891 (N_24891,N_18362,N_19980);
xor U24892 (N_24892,N_15226,N_17528);
nor U24893 (N_24893,N_18534,N_17620);
nor U24894 (N_24894,N_18234,N_18951);
or U24895 (N_24895,N_19402,N_19135);
nand U24896 (N_24896,N_18341,N_19289);
and U24897 (N_24897,N_19846,N_19902);
xor U24898 (N_24898,N_17139,N_19259);
nor U24899 (N_24899,N_17583,N_18985);
nor U24900 (N_24900,N_17427,N_17186);
or U24901 (N_24901,N_18990,N_19451);
xor U24902 (N_24902,N_18919,N_18562);
or U24903 (N_24903,N_17544,N_17336);
and U24904 (N_24904,N_16593,N_19134);
xnor U24905 (N_24905,N_16581,N_18819);
and U24906 (N_24906,N_17464,N_15087);
xor U24907 (N_24907,N_17985,N_15842);
xor U24908 (N_24908,N_18810,N_19081);
and U24909 (N_24909,N_19627,N_19436);
nor U24910 (N_24910,N_19107,N_19173);
nand U24911 (N_24911,N_18129,N_16379);
nor U24912 (N_24912,N_17592,N_16069);
and U24913 (N_24913,N_18112,N_17376);
xor U24914 (N_24914,N_15829,N_19150);
nor U24915 (N_24915,N_18717,N_17667);
or U24916 (N_24916,N_16126,N_15412);
and U24917 (N_24917,N_18448,N_16131);
or U24918 (N_24918,N_15967,N_18864);
nand U24919 (N_24919,N_16068,N_16591);
xnor U24920 (N_24920,N_18506,N_19684);
and U24921 (N_24921,N_17239,N_19152);
nor U24922 (N_24922,N_17629,N_17607);
xnor U24923 (N_24923,N_19934,N_17127);
and U24924 (N_24924,N_15278,N_17763);
or U24925 (N_24925,N_19287,N_19325);
xnor U24926 (N_24926,N_17946,N_15415);
nor U24927 (N_24927,N_17835,N_16431);
xnor U24928 (N_24928,N_15962,N_18828);
nand U24929 (N_24929,N_17356,N_17591);
xnor U24930 (N_24930,N_18633,N_17092);
nor U24931 (N_24931,N_18292,N_16995);
or U24932 (N_24932,N_17225,N_16680);
nand U24933 (N_24933,N_19419,N_17425);
and U24934 (N_24934,N_18449,N_17718);
nor U24935 (N_24935,N_19226,N_19642);
nand U24936 (N_24936,N_15697,N_15834);
and U24937 (N_24937,N_19035,N_15369);
xor U24938 (N_24938,N_18225,N_19011);
or U24939 (N_24939,N_17544,N_15760);
nor U24940 (N_24940,N_15690,N_19298);
nor U24941 (N_24941,N_18818,N_17450);
xnor U24942 (N_24942,N_16957,N_19866);
nor U24943 (N_24943,N_19649,N_17210);
and U24944 (N_24944,N_15573,N_19863);
nor U24945 (N_24945,N_16356,N_18883);
nor U24946 (N_24946,N_17709,N_15030);
nor U24947 (N_24947,N_18488,N_19348);
nand U24948 (N_24948,N_18437,N_15021);
xnor U24949 (N_24949,N_19961,N_17571);
or U24950 (N_24950,N_16647,N_18016);
or U24951 (N_24951,N_15960,N_15505);
or U24952 (N_24952,N_18155,N_16522);
or U24953 (N_24953,N_19562,N_18287);
nand U24954 (N_24954,N_16651,N_18086);
and U24955 (N_24955,N_19064,N_15685);
xor U24956 (N_24956,N_15821,N_15247);
or U24957 (N_24957,N_18558,N_19527);
xor U24958 (N_24958,N_16538,N_16646);
nand U24959 (N_24959,N_17561,N_19065);
xnor U24960 (N_24960,N_16634,N_17816);
nand U24961 (N_24961,N_18060,N_15321);
xor U24962 (N_24962,N_18718,N_16089);
and U24963 (N_24963,N_19645,N_18434);
xnor U24964 (N_24964,N_19447,N_18566);
xnor U24965 (N_24965,N_18154,N_17521);
nor U24966 (N_24966,N_16853,N_16673);
nor U24967 (N_24967,N_16962,N_18270);
nand U24968 (N_24968,N_17136,N_17549);
nor U24969 (N_24969,N_15686,N_15257);
xnor U24970 (N_24970,N_15519,N_18649);
nor U24971 (N_24971,N_15686,N_18316);
or U24972 (N_24972,N_19745,N_15567);
nor U24973 (N_24973,N_18452,N_19090);
nand U24974 (N_24974,N_18027,N_15572);
nor U24975 (N_24975,N_17486,N_19417);
nand U24976 (N_24976,N_15666,N_16147);
and U24977 (N_24977,N_15397,N_19605);
and U24978 (N_24978,N_17111,N_17611);
nor U24979 (N_24979,N_18325,N_19209);
and U24980 (N_24980,N_19144,N_17437);
xnor U24981 (N_24981,N_15270,N_15346);
xor U24982 (N_24982,N_18178,N_17417);
xnor U24983 (N_24983,N_19621,N_17352);
and U24984 (N_24984,N_15230,N_15429);
and U24985 (N_24985,N_19677,N_15601);
nand U24986 (N_24986,N_18884,N_15406);
nor U24987 (N_24987,N_15910,N_19999);
and U24988 (N_24988,N_18269,N_19326);
nor U24989 (N_24989,N_17250,N_19372);
xnor U24990 (N_24990,N_17891,N_16190);
xor U24991 (N_24991,N_15423,N_16003);
or U24992 (N_24992,N_15125,N_16945);
and U24993 (N_24993,N_15671,N_15617);
xor U24994 (N_24994,N_18779,N_15455);
nand U24995 (N_24995,N_19084,N_17425);
nor U24996 (N_24996,N_15363,N_15654);
and U24997 (N_24997,N_19392,N_19881);
or U24998 (N_24998,N_16911,N_19933);
nor U24999 (N_24999,N_15179,N_16551);
nor U25000 (N_25000,N_24745,N_21388);
xnor U25001 (N_25001,N_21282,N_23081);
and U25002 (N_25002,N_21198,N_23313);
xor U25003 (N_25003,N_20239,N_20511);
nand U25004 (N_25004,N_21721,N_21000);
nand U25005 (N_25005,N_21977,N_24103);
xor U25006 (N_25006,N_22301,N_20722);
or U25007 (N_25007,N_24787,N_23272);
nor U25008 (N_25008,N_22770,N_22961);
and U25009 (N_25009,N_21710,N_22827);
nand U25010 (N_25010,N_24935,N_20611);
xnor U25011 (N_25011,N_21438,N_23171);
and U25012 (N_25012,N_24484,N_21760);
xor U25013 (N_25013,N_20122,N_21118);
xor U25014 (N_25014,N_20015,N_21523);
xor U25015 (N_25015,N_24381,N_21991);
xor U25016 (N_25016,N_22552,N_22597);
and U25017 (N_25017,N_22415,N_23705);
and U25018 (N_25018,N_20284,N_22820);
nand U25019 (N_25019,N_20497,N_20642);
nor U25020 (N_25020,N_20594,N_24404);
or U25021 (N_25021,N_22111,N_24122);
xor U25022 (N_25022,N_23973,N_24391);
nand U25023 (N_25023,N_22487,N_20016);
and U25024 (N_25024,N_24359,N_23472);
nand U25025 (N_25025,N_24407,N_21974);
or U25026 (N_25026,N_22678,N_23065);
and U25027 (N_25027,N_22299,N_21079);
xnor U25028 (N_25028,N_22499,N_23382);
xor U25029 (N_25029,N_21683,N_24215);
xor U25030 (N_25030,N_23282,N_22469);
xor U25031 (N_25031,N_23441,N_23002);
nor U25032 (N_25032,N_22927,N_24624);
xor U25033 (N_25033,N_20992,N_20235);
nor U25034 (N_25034,N_23617,N_22033);
nor U25035 (N_25035,N_21166,N_22830);
nor U25036 (N_25036,N_24152,N_23115);
xor U25037 (N_25037,N_24666,N_22443);
nand U25038 (N_25038,N_24064,N_23541);
nor U25039 (N_25039,N_21067,N_20853);
xor U25040 (N_25040,N_21706,N_20931);
or U25041 (N_25041,N_20614,N_22970);
or U25042 (N_25042,N_21866,N_22369);
nand U25043 (N_25043,N_24777,N_24298);
nor U25044 (N_25044,N_20859,N_23068);
xnor U25045 (N_25045,N_23330,N_22782);
xnor U25046 (N_25046,N_21491,N_21782);
or U25047 (N_25047,N_21183,N_23145);
or U25048 (N_25048,N_20954,N_22704);
nand U25049 (N_25049,N_23222,N_24327);
nand U25050 (N_25050,N_24952,N_22730);
and U25051 (N_25051,N_22540,N_21457);
xor U25052 (N_25052,N_24191,N_21854);
and U25053 (N_25053,N_20149,N_23135);
and U25054 (N_25054,N_22878,N_24490);
xnor U25055 (N_25055,N_23049,N_23519);
nand U25056 (N_25056,N_21646,N_23212);
or U25057 (N_25057,N_22658,N_21911);
nand U25058 (N_25058,N_20703,N_20257);
xnor U25059 (N_25059,N_24769,N_24920);
and U25060 (N_25060,N_23527,N_22412);
or U25061 (N_25061,N_21916,N_23084);
and U25062 (N_25062,N_24368,N_20130);
nor U25063 (N_25063,N_24740,N_21841);
nor U25064 (N_25064,N_20393,N_22953);
nand U25065 (N_25065,N_21595,N_23682);
nand U25066 (N_25066,N_24538,N_21535);
xor U25067 (N_25067,N_20255,N_21824);
nor U25068 (N_25068,N_22100,N_20182);
nand U25069 (N_25069,N_21377,N_20532);
nor U25070 (N_25070,N_24078,N_23545);
nor U25071 (N_25071,N_21694,N_22008);
nor U25072 (N_25072,N_23626,N_21046);
nand U25073 (N_25073,N_21026,N_22309);
and U25074 (N_25074,N_20377,N_24350);
and U25075 (N_25075,N_24402,N_24377);
nand U25076 (N_25076,N_20081,N_24523);
and U25077 (N_25077,N_20647,N_20870);
or U25078 (N_25078,N_20401,N_21141);
xnor U25079 (N_25079,N_20738,N_24856);
nand U25080 (N_25080,N_22910,N_20638);
and U25081 (N_25081,N_23418,N_23210);
xor U25082 (N_25082,N_24307,N_23616);
xor U25083 (N_25083,N_23742,N_22074);
or U25084 (N_25084,N_21101,N_24545);
or U25085 (N_25085,N_20430,N_24099);
nor U25086 (N_25086,N_22608,N_20460);
or U25087 (N_25087,N_22222,N_22615);
and U25088 (N_25088,N_22439,N_20335);
or U25089 (N_25089,N_24921,N_20482);
nor U25090 (N_25090,N_22146,N_21555);
or U25091 (N_25091,N_24123,N_23880);
nor U25092 (N_25092,N_20431,N_24694);
and U25093 (N_25093,N_21328,N_22472);
nand U25094 (N_25094,N_21990,N_23121);
nor U25095 (N_25095,N_20047,N_23345);
nand U25096 (N_25096,N_20515,N_21493);
and U25097 (N_25097,N_24847,N_24287);
and U25098 (N_25098,N_20330,N_21013);
and U25099 (N_25099,N_21704,N_23844);
xnor U25100 (N_25100,N_24770,N_24221);
and U25101 (N_25101,N_21981,N_24664);
or U25102 (N_25102,N_20767,N_23646);
xnor U25103 (N_25103,N_23846,N_21675);
and U25104 (N_25104,N_24303,N_20312);
xnor U25105 (N_25105,N_20058,N_22176);
xor U25106 (N_25106,N_20351,N_24255);
and U25107 (N_25107,N_21269,N_20832);
xnor U25108 (N_25108,N_24727,N_21467);
and U25109 (N_25109,N_20710,N_20171);
nand U25110 (N_25110,N_24764,N_20390);
nand U25111 (N_25111,N_22977,N_23079);
xor U25112 (N_25112,N_22248,N_20984);
nor U25113 (N_25113,N_24562,N_20543);
xor U25114 (N_25114,N_20461,N_20817);
and U25115 (N_25115,N_22598,N_20368);
xnor U25116 (N_25116,N_20571,N_23581);
nor U25117 (N_25117,N_20143,N_20061);
nor U25118 (N_25118,N_21811,N_20849);
nand U25119 (N_25119,N_24522,N_23580);
and U25120 (N_25120,N_22793,N_24521);
or U25121 (N_25121,N_21796,N_24370);
and U25122 (N_25122,N_21436,N_23673);
or U25123 (N_25123,N_21756,N_21909);
and U25124 (N_25124,N_24650,N_21835);
or U25125 (N_25125,N_23807,N_21879);
nor U25126 (N_25126,N_21507,N_22320);
nand U25127 (N_25127,N_23477,N_23924);
and U25128 (N_25128,N_23738,N_24412);
nand U25129 (N_25129,N_23398,N_20799);
xnor U25130 (N_25130,N_23565,N_23854);
or U25131 (N_25131,N_23420,N_23215);
nor U25132 (N_25132,N_24248,N_24912);
or U25133 (N_25133,N_23336,N_23730);
xnor U25134 (N_25134,N_22105,N_20729);
nor U25135 (N_25135,N_22705,N_20822);
or U25136 (N_25136,N_22509,N_23283);
nor U25137 (N_25137,N_23310,N_23062);
nor U25138 (N_25138,N_24133,N_23518);
and U25139 (N_25139,N_22959,N_23586);
and U25140 (N_25140,N_21908,N_24970);
or U25141 (N_25141,N_24448,N_24837);
nor U25142 (N_25142,N_24918,N_24037);
xnor U25143 (N_25143,N_23359,N_20165);
xor U25144 (N_25144,N_24803,N_23030);
and U25145 (N_25145,N_23090,N_23100);
or U25146 (N_25146,N_24372,N_23976);
and U25147 (N_25147,N_21725,N_21248);
and U25148 (N_25148,N_22913,N_20888);
and U25149 (N_25149,N_23813,N_23861);
or U25150 (N_25150,N_22520,N_24286);
nand U25151 (N_25151,N_20457,N_24949);
or U25152 (N_25152,N_24826,N_22502);
or U25153 (N_25153,N_21759,N_21330);
nor U25154 (N_25154,N_20452,N_22297);
xor U25155 (N_25155,N_24212,N_23899);
xnor U25156 (N_25156,N_23944,N_24534);
xor U25157 (N_25157,N_24177,N_20684);
nor U25158 (N_25158,N_23845,N_20475);
nor U25159 (N_25159,N_20116,N_22281);
xor U25160 (N_25160,N_24528,N_20289);
or U25161 (N_25161,N_20727,N_24138);
nand U25162 (N_25162,N_22543,N_22776);
xor U25163 (N_25163,N_23915,N_22319);
and U25164 (N_25164,N_24023,N_21015);
nor U25165 (N_25165,N_22138,N_21111);
and U25166 (N_25166,N_20740,N_21427);
nor U25167 (N_25167,N_20092,N_24786);
and U25168 (N_25168,N_23631,N_20785);
and U25169 (N_25169,N_24604,N_21016);
nor U25170 (N_25170,N_24956,N_20693);
xnor U25171 (N_25171,N_22724,N_20796);
and U25172 (N_25172,N_21913,N_24638);
and U25173 (N_25173,N_20499,N_22219);
xor U25174 (N_25174,N_20744,N_21790);
xnor U25175 (N_25175,N_20108,N_23059);
nor U25176 (N_25176,N_23599,N_20695);
and U25177 (N_25177,N_21424,N_22330);
and U25178 (N_25178,N_20947,N_24225);
xor U25179 (N_25179,N_22651,N_22584);
nand U25180 (N_25180,N_23715,N_21439);
nand U25181 (N_25181,N_22432,N_20798);
or U25182 (N_25182,N_22039,N_22424);
or U25183 (N_25183,N_20220,N_22789);
nor U25184 (N_25184,N_21559,N_24507);
nor U25185 (N_25185,N_22103,N_24348);
or U25186 (N_25186,N_23625,N_21834);
or U25187 (N_25187,N_23560,N_21476);
xor U25188 (N_25188,N_23908,N_22852);
xor U25189 (N_25189,N_24750,N_20121);
or U25190 (N_25190,N_24986,N_22433);
xnor U25191 (N_25191,N_23707,N_24774);
and U25192 (N_25192,N_23654,N_20236);
and U25193 (N_25193,N_24932,N_22191);
xnor U25194 (N_25194,N_24821,N_22168);
or U25195 (N_25195,N_22477,N_23525);
nor U25196 (N_25196,N_21784,N_21283);
or U25197 (N_25197,N_24473,N_24260);
xnor U25198 (N_25198,N_21090,N_21805);
nor U25199 (N_25199,N_23549,N_21946);
nand U25200 (N_25200,N_20297,N_22195);
nor U25201 (N_25201,N_24880,N_24382);
and U25202 (N_25202,N_24502,N_22802);
nand U25203 (N_25203,N_21413,N_21040);
xor U25204 (N_25204,N_20483,N_21024);
xnor U25205 (N_25205,N_20787,N_24100);
nor U25206 (N_25206,N_23832,N_23526);
or U25207 (N_25207,N_24200,N_24462);
xnor U25208 (N_25208,N_20552,N_20506);
and U25209 (N_25209,N_24478,N_21979);
nand U25210 (N_25210,N_22693,N_21754);
nor U25211 (N_25211,N_24074,N_23674);
and U25212 (N_25212,N_24397,N_21406);
or U25213 (N_25213,N_21028,N_24414);
nand U25214 (N_25214,N_24576,N_24275);
xor U25215 (N_25215,N_22924,N_20714);
or U25216 (N_25216,N_20656,N_24347);
xnor U25217 (N_25217,N_22925,N_23149);
nor U25218 (N_25218,N_22946,N_22044);
xnor U25219 (N_25219,N_21043,N_22339);
nand U25220 (N_25220,N_20355,N_21259);
nand U25221 (N_25221,N_20476,N_24127);
nand U25222 (N_25222,N_20986,N_24976);
nor U25223 (N_25223,N_20871,N_23797);
and U25224 (N_25224,N_23873,N_23781);
nand U25225 (N_25225,N_22649,N_22336);
nand U25226 (N_25226,N_20155,N_21478);
nor U25227 (N_25227,N_21787,N_21048);
xnor U25228 (N_25228,N_24366,N_22786);
nor U25229 (N_25229,N_24360,N_22032);
or U25230 (N_25230,N_23630,N_21082);
or U25231 (N_25231,N_23988,N_21757);
nor U25232 (N_25232,N_23902,N_24866);
xor U25233 (N_25233,N_20109,N_21679);
and U25234 (N_25234,N_21623,N_24006);
xnor U25235 (N_25235,N_24991,N_21110);
or U25236 (N_25236,N_23614,N_20129);
or U25237 (N_25237,N_20111,N_24852);
nor U25238 (N_25238,N_20494,N_21386);
or U25239 (N_25239,N_24306,N_22277);
and U25240 (N_25240,N_20365,N_22161);
xnor U25241 (N_25241,N_21156,N_24336);
and U25242 (N_25242,N_23403,N_22162);
or U25243 (N_25243,N_20914,N_22148);
xor U25244 (N_25244,N_24855,N_20559);
xnor U25245 (N_25245,N_24083,N_24539);
nand U25246 (N_25246,N_23139,N_21140);
and U25247 (N_25247,N_24483,N_23935);
nor U25248 (N_25248,N_24959,N_21394);
nand U25249 (N_25249,N_23177,N_24238);
nand U25250 (N_25250,N_23865,N_21812);
and U25251 (N_25251,N_22566,N_21634);
or U25252 (N_25252,N_21963,N_22674);
or U25253 (N_25253,N_20887,N_21772);
nand U25254 (N_25254,N_23265,N_20731);
xnor U25255 (N_25255,N_24120,N_23971);
nor U25256 (N_25256,N_20901,N_24536);
nor U25257 (N_25257,N_24311,N_24595);
and U25258 (N_25258,N_21465,N_22455);
and U25259 (N_25259,N_23633,N_24820);
xnor U25260 (N_25260,N_23461,N_21393);
nor U25261 (N_25261,N_23685,N_23702);
and U25262 (N_25262,N_20464,N_20200);
or U25263 (N_25263,N_23878,N_24645);
or U25264 (N_25264,N_20031,N_21437);
nand U25265 (N_25265,N_24457,N_21309);
xor U25266 (N_25266,N_24631,N_22885);
xor U25267 (N_25267,N_22861,N_21045);
and U25268 (N_25268,N_20449,N_23594);
nor U25269 (N_25269,N_20950,N_24456);
nand U25270 (N_25270,N_22533,N_23105);
or U25271 (N_25271,N_23304,N_24566);
nand U25272 (N_25272,N_24106,N_22104);
or U25273 (N_25273,N_22694,N_24889);
and U25274 (N_25274,N_21144,N_21629);
nand U25275 (N_25275,N_20724,N_21551);
xnor U25276 (N_25276,N_20999,N_20895);
and U25277 (N_25277,N_20180,N_24395);
nor U25278 (N_25278,N_21602,N_22828);
nor U25279 (N_25279,N_22722,N_22690);
and U25280 (N_25280,N_22147,N_23077);
nand U25281 (N_25281,N_20758,N_21355);
or U25282 (N_25282,N_22967,N_23713);
and U25283 (N_25283,N_23319,N_24273);
or U25284 (N_25284,N_22115,N_23666);
and U25285 (N_25285,N_20934,N_22485);
nand U25286 (N_25286,N_21795,N_22645);
nand U25287 (N_25287,N_24280,N_22059);
xnor U25288 (N_25288,N_21366,N_23669);
xnor U25289 (N_25289,N_21297,N_20565);
or U25290 (N_25290,N_24620,N_20846);
or U25291 (N_25291,N_24182,N_24213);
nor U25292 (N_25292,N_20359,N_23452);
and U25293 (N_25293,N_23196,N_21264);
nand U25294 (N_25294,N_22949,N_20343);
nand U25295 (N_25295,N_21321,N_22846);
or U25296 (N_25296,N_23697,N_24198);
nor U25297 (N_25297,N_24877,N_20117);
or U25298 (N_25298,N_20523,N_20959);
and U25299 (N_25299,N_23737,N_21041);
nor U25300 (N_25300,N_21052,N_20521);
xnor U25301 (N_25301,N_22132,N_20649);
nor U25302 (N_25302,N_22327,N_22560);
nand U25303 (N_25303,N_24008,N_24088);
nand U25304 (N_25304,N_20572,N_22200);
and U25305 (N_25305,N_21428,N_23369);
nor U25306 (N_25306,N_24527,N_23447);
nor U25307 (N_25307,N_23677,N_20309);
or U25308 (N_25308,N_23939,N_20604);
nor U25309 (N_25309,N_21687,N_23311);
xnor U25310 (N_25310,N_23401,N_20056);
and U25311 (N_25311,N_21800,N_24540);
xnor U25312 (N_25312,N_24897,N_23486);
nor U25313 (N_25313,N_20858,N_24227);
nor U25314 (N_25314,N_23089,N_22568);
nand U25315 (N_25315,N_24430,N_24868);
and U25316 (N_25316,N_21976,N_22960);
or U25317 (N_25317,N_22869,N_21578);
nor U25318 (N_25318,N_21189,N_22398);
or U25319 (N_25319,N_24957,N_23082);
nor U25320 (N_25320,N_22080,N_22733);
or U25321 (N_25321,N_21238,N_21997);
xnor U25322 (N_25322,N_23411,N_23800);
nor U25323 (N_25323,N_22594,N_21713);
and U25324 (N_25324,N_22224,N_24843);
xnor U25325 (N_25325,N_20928,N_24767);
xnor U25326 (N_25326,N_20779,N_24885);
nand U25327 (N_25327,N_24597,N_20286);
or U25328 (N_25328,N_21237,N_20933);
nand U25329 (N_25329,N_21865,N_22187);
xnor U25330 (N_25330,N_21218,N_23920);
xor U25331 (N_25331,N_23621,N_23957);
nor U25332 (N_25332,N_22585,N_21888);
and U25333 (N_25333,N_23812,N_20921);
and U25334 (N_25334,N_20020,N_21654);
xnor U25335 (N_25335,N_21587,N_24184);
or U25336 (N_25336,N_20545,N_20935);
or U25337 (N_25337,N_20011,N_23695);
or U25338 (N_25338,N_22565,N_24905);
and U25339 (N_25339,N_22778,N_24158);
nand U25340 (N_25340,N_21272,N_23406);
or U25341 (N_25341,N_24310,N_22091);
or U25342 (N_25342,N_21063,N_22947);
xor U25343 (N_25343,N_22557,N_21918);
nand U25344 (N_25344,N_21767,N_21980);
nor U25345 (N_25345,N_23814,N_22832);
or U25346 (N_25346,N_21186,N_22288);
xnor U25347 (N_25347,N_22895,N_21996);
and U25348 (N_25348,N_21160,N_24489);
nand U25349 (N_25349,N_20002,N_23760);
xor U25350 (N_25350,N_23003,N_24505);
and U25351 (N_25351,N_20749,N_22631);
or U25352 (N_25352,N_23236,N_20453);
and U25353 (N_25353,N_24076,N_24228);
xnor U25354 (N_25354,N_21745,N_20175);
and U25355 (N_25355,N_22049,N_20154);
and U25356 (N_25356,N_23153,N_21512);
nand U25357 (N_25357,N_20989,N_24572);
and U25358 (N_25358,N_24333,N_21382);
and U25359 (N_25359,N_24095,N_22024);
nor U25360 (N_25360,N_21290,N_21858);
and U25361 (N_25361,N_20184,N_24726);
nand U25362 (N_25362,N_21064,N_20367);
nor U25363 (N_25363,N_23710,N_20114);
xnor U25364 (N_25364,N_22289,N_22210);
or U25365 (N_25365,N_23204,N_20403);
or U25366 (N_25366,N_21674,N_23480);
or U25367 (N_25367,N_24474,N_24809);
or U25368 (N_25368,N_21983,N_24715);
nor U25369 (N_25369,N_21182,N_23493);
nor U25370 (N_25370,N_21137,N_24563);
xnor U25371 (N_25371,N_21825,N_21481);
nand U25372 (N_25372,N_23914,N_22069);
or U25373 (N_25373,N_24493,N_23629);
or U25374 (N_25374,N_23086,N_24676);
and U25375 (N_25375,N_23261,N_24771);
xor U25376 (N_25376,N_21022,N_21444);
or U25377 (N_25377,N_23628,N_22872);
or U25378 (N_25378,N_21071,N_24613);
or U25379 (N_25379,N_20007,N_22152);
xnor U25380 (N_25380,N_20411,N_24048);
and U25381 (N_25381,N_23749,N_24185);
and U25382 (N_25382,N_23799,N_22928);
nand U25383 (N_25383,N_23190,N_21263);
or U25384 (N_25384,N_21148,N_22030);
nand U25385 (N_25385,N_23442,N_23021);
nand U25386 (N_25386,N_24605,N_23798);
and U25387 (N_25387,N_21840,N_20361);
nor U25388 (N_25388,N_24374,N_20616);
xnor U25389 (N_25389,N_20067,N_22882);
xnor U25390 (N_25390,N_23469,N_21904);
and U25391 (N_25391,N_24043,N_20179);
and U25392 (N_25392,N_21032,N_23847);
nand U25393 (N_25393,N_23627,N_22285);
nor U25394 (N_25394,N_21116,N_20414);
nand U25395 (N_25395,N_20232,N_23026);
and U25396 (N_25396,N_23934,N_22506);
or U25397 (N_25397,N_21543,N_24199);
or U25398 (N_25398,N_24135,N_22078);
and U25399 (N_25399,N_22448,N_24601);
or U25400 (N_25400,N_22604,N_22655);
nor U25401 (N_25401,N_22648,N_24719);
xnor U25402 (N_25402,N_22613,N_24762);
nand U25403 (N_25403,N_23507,N_23980);
nand U25404 (N_25404,N_24141,N_24069);
nor U25405 (N_25405,N_20689,N_21487);
and U25406 (N_25406,N_23911,N_22708);
nor U25407 (N_25407,N_24222,N_23804);
nor U25408 (N_25408,N_24585,N_21047);
xnor U25409 (N_25409,N_21104,N_21716);
nand U25410 (N_25410,N_24600,N_22083);
xor U25411 (N_25411,N_21536,N_20544);
and U25412 (N_25412,N_24071,N_20160);
or U25413 (N_25413,N_21668,N_22262);
or U25414 (N_25414,N_21228,N_24284);
xnor U25415 (N_25415,N_20434,N_20864);
nand U25416 (N_25416,N_24926,N_23053);
or U25417 (N_25417,N_24156,N_22159);
nor U25418 (N_25418,N_21294,N_23664);
nand U25419 (N_25419,N_24394,N_24161);
and U25420 (N_25420,N_22976,N_24201);
and U25421 (N_25421,N_22201,N_23985);
or U25422 (N_25422,N_22257,N_20396);
and U25423 (N_25423,N_22729,N_23517);
nand U25424 (N_25424,N_23254,N_22466);
nor U25425 (N_25425,N_20503,N_23512);
nor U25426 (N_25426,N_24798,N_22984);
and U25427 (N_25427,N_24568,N_23922);
or U25428 (N_25428,N_24429,N_21868);
or U25429 (N_25429,N_21243,N_24279);
and U25430 (N_25430,N_22788,N_23427);
or U25431 (N_25431,N_20211,N_24709);
nor U25432 (N_25432,N_21097,N_23037);
xnor U25433 (N_25433,N_20209,N_23096);
and U25434 (N_25434,N_21372,N_22605);
and U25435 (N_25435,N_22242,N_20444);
or U25436 (N_25436,N_20610,N_23925);
or U25437 (N_25437,N_21972,N_20395);
and U25438 (N_25438,N_24934,N_20549);
nor U25439 (N_25439,N_22973,N_23963);
and U25440 (N_25440,N_21289,N_22562);
and U25441 (N_25441,N_21055,N_24070);
nor U25442 (N_25442,N_24881,N_20823);
or U25443 (N_25443,N_20620,N_21875);
nor U25444 (N_25444,N_22268,N_21752);
or U25445 (N_25445,N_24706,N_20905);
or U25446 (N_25446,N_20978,N_20485);
or U25447 (N_25447,N_23396,N_20314);
xor U25448 (N_25448,N_24371,N_21851);
or U25449 (N_25449,N_21459,N_23488);
nor U25450 (N_25450,N_24910,N_23424);
xnor U25451 (N_25451,N_23597,N_24357);
nor U25452 (N_25452,N_21220,N_20484);
or U25453 (N_25453,N_23645,N_23822);
nor U25454 (N_25454,N_21226,N_24685);
and U25455 (N_25455,N_24157,N_20400);
nor U25456 (N_25456,N_20378,N_21590);
nand U25457 (N_25457,N_23000,N_20436);
and U25458 (N_25458,N_22392,N_22018);
or U25459 (N_25459,N_20546,N_23205);
nand U25460 (N_25460,N_20215,N_23009);
or U25461 (N_25461,N_20890,N_24872);
nor U25462 (N_25462,N_23603,N_24558);
nor U25463 (N_25463,N_21842,N_23775);
and U25464 (N_25464,N_20227,N_22873);
or U25465 (N_25465,N_20174,N_23368);
xor U25466 (N_25466,N_21769,N_23387);
nor U25467 (N_25467,N_21336,N_24955);
and U25468 (N_25468,N_23719,N_24324);
nor U25469 (N_25469,N_23332,N_21054);
xor U25470 (N_25470,N_22462,N_24176);
xnor U25471 (N_25471,N_24827,N_21454);
or U25472 (N_25472,N_23166,N_21254);
nor U25473 (N_25473,N_24968,N_22130);
nor U25474 (N_25474,N_24463,N_23200);
xor U25475 (N_25475,N_20306,N_22000);
nor U25476 (N_25476,N_22429,N_21300);
xor U25477 (N_25477,N_23838,N_22348);
nor U25478 (N_25478,N_22932,N_20707);
nand U25479 (N_25479,N_21419,N_23324);
and U25480 (N_25480,N_24684,N_22246);
xnor U25481 (N_25481,N_23502,N_24349);
nor U25482 (N_25482,N_22899,N_23448);
and U25483 (N_25483,N_23979,N_24170);
nand U25484 (N_25484,N_20135,N_21030);
nand U25485 (N_25485,N_20037,N_24178);
xnor U25486 (N_25486,N_24708,N_24258);
nor U25487 (N_25487,N_22986,N_22774);
nand U25488 (N_25488,N_21849,N_20981);
or U25489 (N_25489,N_23439,N_24633);
nand U25490 (N_25490,N_21065,N_23958);
or U25491 (N_25491,N_22373,N_24654);
or U25492 (N_25492,N_20558,N_21876);
and U25493 (N_25493,N_24626,N_24254);
nand U25494 (N_25494,N_22792,N_23917);
nor U25495 (N_25495,N_22186,N_21447);
nand U25496 (N_25496,N_23223,N_20646);
or U25497 (N_25497,N_21608,N_24186);
and U25498 (N_25498,N_23591,N_20221);
or U25499 (N_25499,N_23843,N_21105);
xnor U25500 (N_25500,N_23791,N_23444);
or U25501 (N_25501,N_20666,N_23735);
nand U25502 (N_25502,N_21267,N_21936);
nand U25503 (N_25503,N_22101,N_21853);
or U25504 (N_25504,N_24229,N_20086);
xnor U25505 (N_25505,N_21216,N_23046);
xnor U25506 (N_25506,N_21932,N_20648);
xor U25507 (N_25507,N_23972,N_24683);
or U25508 (N_25508,N_23294,N_23011);
nor U25509 (N_25509,N_20605,N_22530);
nand U25510 (N_25510,N_20996,N_22914);
nand U25511 (N_25511,N_23022,N_21008);
nor U25512 (N_25512,N_20074,N_20674);
or U25513 (N_25513,N_24496,N_22823);
nor U25514 (N_25514,N_20014,N_20191);
or U25515 (N_25515,N_21338,N_21954);
or U25516 (N_25516,N_20726,N_23375);
nand U25517 (N_25517,N_22212,N_24834);
and U25518 (N_25518,N_20023,N_20124);
and U25519 (N_25519,N_22393,N_21720);
nand U25520 (N_25520,N_24044,N_21268);
nand U25521 (N_25521,N_20913,N_21942);
or U25522 (N_25522,N_21152,N_22264);
nand U25523 (N_25523,N_24791,N_22276);
and U25524 (N_25524,N_21662,N_23101);
nand U25525 (N_25525,N_23643,N_22022);
nand U25526 (N_25526,N_24197,N_22384);
and U25527 (N_25527,N_20911,N_22994);
nand U25528 (N_25528,N_20373,N_23724);
xnor U25529 (N_25529,N_22476,N_20326);
and U25530 (N_25530,N_20358,N_21532);
nand U25531 (N_25531,N_22449,N_21093);
nor U25532 (N_25532,N_21092,N_21761);
nor U25533 (N_25533,N_22360,N_24781);
and U25534 (N_25534,N_20421,N_21059);
and U25535 (N_25535,N_21766,N_22640);
nand U25536 (N_25536,N_22511,N_22982);
or U25537 (N_25537,N_22785,N_22575);
nand U25538 (N_25538,N_21322,N_24256);
nor U25539 (N_25539,N_23093,N_20219);
nand U25540 (N_25540,N_24183,N_21563);
nor U25541 (N_25541,N_21733,N_20697);
and U25542 (N_25542,N_24737,N_22985);
or U25543 (N_25543,N_23831,N_21074);
nand U25544 (N_25544,N_24615,N_24865);
nor U25545 (N_25545,N_24046,N_23242);
xor U25546 (N_25546,N_24365,N_24444);
nor U25547 (N_25547,N_24805,N_22418);
and U25548 (N_25548,N_23655,N_23912);
nor U25549 (N_25549,N_21534,N_23563);
or U25550 (N_25550,N_22290,N_24984);
nand U25551 (N_25551,N_24579,N_20806);
xor U25552 (N_25552,N_23918,N_23363);
nor U25553 (N_25553,N_20345,N_20525);
nand U25554 (N_25554,N_23712,N_23647);
nand U25555 (N_25555,N_20064,N_22437);
xor U25556 (N_25556,N_22736,N_22845);
and U25557 (N_25557,N_23458,N_22937);
and U25558 (N_25558,N_21901,N_23353);
nor U25559 (N_25559,N_23821,N_21978);
xor U25560 (N_25560,N_20944,N_22160);
nor U25561 (N_25561,N_23394,N_24239);
nand U25562 (N_25562,N_21605,N_20148);
nor U25563 (N_25563,N_23989,N_24065);
or U25564 (N_25564,N_24831,N_22865);
and U25565 (N_25565,N_21353,N_20754);
nor U25566 (N_25566,N_23170,N_22596);
nor U25567 (N_25567,N_22536,N_21554);
nor U25568 (N_25568,N_21609,N_24492);
and U25569 (N_25569,N_24796,N_21688);
xor U25570 (N_25570,N_21398,N_23243);
or U25571 (N_25571,N_21917,N_22208);
and U25572 (N_25572,N_23041,N_21776);
nand U25573 (N_25573,N_22417,N_21124);
nand U25574 (N_25574,N_23701,N_20385);
nor U25575 (N_25575,N_23228,N_21396);
xor U25576 (N_25576,N_21537,N_23227);
or U25577 (N_25577,N_23709,N_24824);
or U25578 (N_25578,N_22535,N_22909);
xor U25579 (N_25579,N_24590,N_24166);
xor U25580 (N_25580,N_20146,N_20467);
nor U25581 (N_25581,N_22305,N_22659);
and U25582 (N_25582,N_22696,N_24220);
or U25583 (N_25583,N_23887,N_21698);
nand U25584 (N_25584,N_21399,N_24148);
nand U25585 (N_25585,N_21864,N_20465);
and U25586 (N_25586,N_23747,N_22809);
nor U25587 (N_25587,N_22980,N_23191);
nor U25588 (N_25588,N_21184,N_20454);
nor U25589 (N_25589,N_21397,N_21181);
xnor U25590 (N_25590,N_21892,N_20048);
nand U25591 (N_25591,N_23462,N_22175);
nand U25592 (N_25592,N_24907,N_22076);
nand U25593 (N_25593,N_22060,N_21277);
nand U25594 (N_25594,N_21743,N_22529);
or U25595 (N_25595,N_23995,N_22085);
and U25596 (N_25596,N_24388,N_20994);
and U25597 (N_25597,N_24680,N_22790);
and U25598 (N_25598,N_24063,N_22108);
nand U25599 (N_25599,N_23870,N_23913);
and U25600 (N_25600,N_20059,N_22545);
or U25601 (N_25601,N_24844,N_20520);
or U25602 (N_25602,N_20202,N_22886);
xnor U25603 (N_25603,N_22874,N_22554);
and U25604 (N_25604,N_24015,N_24776);
or U25605 (N_25605,N_23379,N_22550);
nand U25606 (N_25606,N_20469,N_20397);
xnor U25607 (N_25607,N_21612,N_24479);
nand U25608 (N_25608,N_23860,N_24396);
and U25609 (N_25609,N_22062,N_22754);
and U25610 (N_25610,N_20163,N_20075);
nand U25611 (N_25611,N_20293,N_22758);
xor U25612 (N_25612,N_20915,N_21468);
nand U25613 (N_25613,N_21469,N_21881);
nor U25614 (N_25614,N_23970,N_22075);
xor U25615 (N_25615,N_21882,N_22410);
nor U25616 (N_25616,N_21636,N_20185);
and U25617 (N_25617,N_23073,N_21391);
nand U25618 (N_25618,N_21247,N_23225);
and U25619 (N_25619,N_20903,N_23900);
nand U25620 (N_25620,N_21597,N_20415);
or U25621 (N_25621,N_23095,N_22357);
xnor U25622 (N_25622,N_21677,N_23684);
xor U25623 (N_25623,N_22817,N_21432);
nor U25624 (N_25624,N_20582,N_22478);
or U25625 (N_25625,N_20516,N_22978);
and U25626 (N_25626,N_23606,N_20873);
nand U25627 (N_25627,N_22016,N_20248);
nor U25628 (N_25628,N_21009,N_20634);
or U25629 (N_25629,N_20133,N_21540);
nand U25630 (N_25630,N_20087,N_21162);
xor U25631 (N_25631,N_20567,N_23604);
nor U25632 (N_25632,N_21711,N_24115);
nor U25633 (N_25633,N_20807,N_20340);
nor U25634 (N_25634,N_23499,N_22050);
nand U25635 (N_25635,N_21486,N_20881);
and U25636 (N_25636,N_24111,N_22094);
and U25637 (N_25637,N_24981,N_23314);
nand U25638 (N_25638,N_22703,N_23257);
xnor U25639 (N_25639,N_20338,N_21193);
nor U25640 (N_25640,N_22266,N_23558);
or U25641 (N_25641,N_23696,N_21618);
xor U25642 (N_25642,N_24892,N_23850);
nor U25643 (N_25643,N_20893,N_20910);
xnor U25644 (N_25644,N_22639,N_23317);
or U25645 (N_25645,N_24282,N_22096);
nor U25646 (N_25646,N_20623,N_22833);
nor U25647 (N_25647,N_20249,N_24710);
nand U25648 (N_25648,N_23144,N_20203);
or U25649 (N_25649,N_21291,N_23683);
or U25650 (N_25650,N_21211,N_23136);
nand U25651 (N_25651,N_21197,N_20028);
nand U25652 (N_25652,N_22492,N_21221);
nor U25653 (N_25653,N_20815,N_21617);
nor U25654 (N_25654,N_23316,N_20426);
nor U25655 (N_25655,N_24361,N_21621);
nor U25656 (N_25656,N_23557,N_22541);
xor U25657 (N_25657,N_20537,N_23758);
xor U25658 (N_25658,N_23465,N_24504);
or U25659 (N_25659,N_23698,N_23347);
nor U25660 (N_25660,N_21889,N_23025);
nor U25661 (N_25661,N_23895,N_24418);
or U25662 (N_25662,N_22811,N_22627);
nand U25663 (N_25663,N_21526,N_21262);
or U25664 (N_25664,N_23632,N_24761);
or U25665 (N_25665,N_20865,N_24603);
or U25666 (N_25666,N_21027,N_20573);
or U25667 (N_25667,N_22444,N_20732);
nand U25668 (N_25668,N_24724,N_22172);
nand U25669 (N_25669,N_24721,N_23055);
nor U25670 (N_25670,N_20534,N_22364);
nor U25671 (N_25671,N_23307,N_22252);
nand U25672 (N_25672,N_21544,N_22066);
nand U25673 (N_25673,N_24084,N_23365);
xnor U25674 (N_25674,N_24979,N_24486);
nor U25675 (N_25675,N_24136,N_20548);
or U25676 (N_25676,N_21742,N_24704);
or U25677 (N_25677,N_20741,N_20681);
nor U25678 (N_25678,N_22328,N_24553);
nand U25679 (N_25679,N_24379,N_20372);
nand U25680 (N_25680,N_24196,N_21342);
nor U25681 (N_25681,N_21561,N_23069);
nand U25682 (N_25682,N_21645,N_24358);
and U25683 (N_25683,N_24808,N_24313);
xor U25684 (N_25684,N_23542,N_24508);
and U25685 (N_25685,N_22962,N_24380);
nand U25686 (N_25686,N_24139,N_22921);
or U25687 (N_25687,N_21313,N_20350);
nor U25688 (N_25688,N_20678,N_22218);
nor U25689 (N_25689,N_24050,N_22904);
xnor U25690 (N_25690,N_21356,N_21695);
nand U25691 (N_25691,N_23308,N_22067);
nand U25692 (N_25692,N_22211,N_23492);
xnor U25693 (N_25693,N_22621,N_23826);
and U25694 (N_25694,N_24373,N_23964);
nand U25695 (N_25695,N_21357,N_20387);
xor U25696 (N_25696,N_20592,N_21738);
or U25697 (N_25697,N_21707,N_22363);
nor U25698 (N_25698,N_20409,N_23932);
xnor U25699 (N_25699,N_22042,N_22512);
xnor U25700 (N_25700,N_23548,N_20217);
xor U25701 (N_25701,N_20971,N_23923);
nand U25702 (N_25702,N_24850,N_24697);
nor U25703 (N_25703,N_21011,N_22902);
nand U25704 (N_25704,N_24131,N_20353);
nor U25705 (N_25705,N_22454,N_21944);
and U25706 (N_25706,N_22374,N_24125);
and U25707 (N_25707,N_22063,N_24587);
or U25708 (N_25708,N_23898,N_22863);
nor U25709 (N_25709,N_21014,N_20627);
and U25710 (N_25710,N_24729,N_22856);
xnor U25711 (N_25711,N_24695,N_20900);
or U25712 (N_25712,N_21075,N_21485);
nand U25713 (N_25713,N_22670,N_20410);
nor U25714 (N_25714,N_22123,N_23926);
and U25715 (N_25715,N_23043,N_20794);
nor U25716 (N_25716,N_22151,N_20704);
nor U25717 (N_25717,N_22593,N_23667);
nand U25718 (N_25718,N_24421,N_22688);
and U25719 (N_25719,N_20137,N_23726);
and U25720 (N_25720,N_22835,N_24331);
nor U25721 (N_25721,N_20809,N_23164);
xor U25722 (N_25722,N_23176,N_20487);
or U25723 (N_25723,N_24698,N_22313);
nor U25724 (N_25724,N_24274,N_23023);
and U25725 (N_25725,N_21630,N_21145);
or U25726 (N_25726,N_23015,N_20765);
and U25727 (N_25727,N_22231,N_24612);
xor U25728 (N_25728,N_24319,N_22898);
and U25729 (N_25729,N_24416,N_24062);
and U25730 (N_25730,N_22796,N_22558);
xnor U25731 (N_25731,N_20652,N_20712);
nand U25732 (N_25732,N_23929,N_21236);
and U25733 (N_25733,N_21363,N_23454);
nor U25734 (N_25734,N_24398,N_21434);
nand U25735 (N_25735,N_24739,N_21208);
xor U25736 (N_25736,N_23768,N_20923);
and U25737 (N_25737,N_20489,N_20898);
and U25738 (N_25738,N_24117,N_24596);
nand U25739 (N_25739,N_20357,N_20246);
or U25740 (N_25740,N_24896,N_23506);
or U25741 (N_25741,N_24660,N_20804);
nand U25742 (N_25742,N_21227,N_20344);
and U25743 (N_25743,N_22436,N_24312);
or U25744 (N_25744,N_22644,N_20244);
or U25745 (N_25745,N_23270,N_23195);
and U25746 (N_25746,N_20909,N_20281);
and U25747 (N_25747,N_21653,N_23977);
or U25748 (N_25748,N_23856,N_24058);
nor U25749 (N_25749,N_21373,N_21012);
or U25750 (N_25750,N_20339,N_21951);
nand U25751 (N_25751,N_24410,N_21614);
nand U25752 (N_25752,N_23692,N_24335);
nand U25753 (N_25753,N_24126,N_21087);
nor U25754 (N_25754,N_20706,N_21987);
nand U25755 (N_25755,N_20459,N_22465);
nor U25756 (N_25756,N_22127,N_21775);
nor U25757 (N_25757,N_24175,N_24328);
xor U25758 (N_25758,N_24281,N_23390);
nand U25759 (N_25759,N_21299,N_21455);
nor U25760 (N_25760,N_23350,N_22498);
or U25761 (N_25761,N_20760,N_21723);
nor U25762 (N_25762,N_20561,N_24295);
xnor U25763 (N_25763,N_22570,N_22698);
nor U25764 (N_25764,N_22625,N_20651);
and U25765 (N_25765,N_24641,N_21814);
nor U25766 (N_25766,N_20617,N_21441);
and U25767 (N_25767,N_24634,N_24967);
xnor U25768 (N_25768,N_24592,N_20939);
xor U25769 (N_25769,N_24400,N_23623);
and U25770 (N_25770,N_21528,N_24742);
nand U25771 (N_25771,N_20283,N_24902);
or U25772 (N_25772,N_22842,N_21514);
xnor U25773 (N_25773,N_24231,N_24532);
nand U25774 (N_25774,N_21830,N_23278);
and U25775 (N_25775,N_24271,N_20522);
nand U25776 (N_25776,N_20276,N_23836);
nor U25777 (N_25777,N_20328,N_21903);
and U25778 (N_25778,N_21376,N_23658);
xor U25779 (N_25779,N_21524,N_20471);
nand U25780 (N_25780,N_21973,N_22521);
or U25781 (N_25781,N_21797,N_23315);
and U25782 (N_25782,N_23675,N_21333);
xnor U25783 (N_25783,N_22684,N_24216);
or U25784 (N_25784,N_21592,N_23638);
and U25785 (N_25785,N_22421,N_24096);
and U25786 (N_25786,N_24965,N_23717);
xnor U25787 (N_25787,N_24208,N_21142);
or U25788 (N_25788,N_23998,N_20946);
nand U25789 (N_25789,N_22135,N_22420);
nor U25790 (N_25790,N_24081,N_21195);
nor U25791 (N_25791,N_23165,N_24867);
and U25792 (N_25792,N_24290,N_24922);
and U25793 (N_25793,N_24701,N_24433);
and U25794 (N_25794,N_23635,N_23948);
or U25795 (N_25795,N_24147,N_23892);
xnor U25796 (N_25796,N_24586,N_21943);
xor U25797 (N_25797,N_23300,N_20323);
and U25798 (N_25798,N_21209,N_23947);
xnor U25799 (N_25799,N_23374,N_22496);
xor U25800 (N_25800,N_20138,N_21374);
and U25801 (N_25801,N_24759,N_24632);
nand U25802 (N_25802,N_21187,N_22038);
nand U25803 (N_25803,N_23183,N_24134);
nand U25804 (N_25804,N_21962,N_23779);
and U25805 (N_25805,N_21506,N_21036);
or U25806 (N_25806,N_20863,N_21948);
and U25807 (N_25807,N_24582,N_20833);
nand U25808 (N_25808,N_22931,N_21050);
nand U25809 (N_25809,N_24716,N_21874);
xor U25810 (N_25810,N_21084,N_24614);
or U25811 (N_25811,N_23301,N_22251);
xor U25812 (N_25812,N_22461,N_23148);
nand U25813 (N_25813,N_22620,N_24977);
or U25814 (N_25814,N_22458,N_20407);
xor U25815 (N_25815,N_21125,N_23708);
xnor U25816 (N_25816,N_24040,N_21665);
nand U25817 (N_25817,N_22731,N_22037);
nor U25818 (N_25818,N_22287,N_22810);
nand U25819 (N_25819,N_21863,N_21080);
nand U25820 (N_25820,N_23555,N_21113);
nand U25821 (N_25821,N_22838,N_20491);
nand U25822 (N_25822,N_21381,N_21123);
and U25823 (N_25823,N_22507,N_20958);
and U25824 (N_25824,N_20920,N_24236);
nor U25825 (N_25825,N_24818,N_22404);
and U25826 (N_25826,N_22347,N_20517);
nor U25827 (N_25827,N_21301,N_23772);
nor U25828 (N_25828,N_23325,N_23490);
nor U25829 (N_25829,N_23582,N_22523);
xor U25830 (N_25830,N_23494,N_24784);
and U25831 (N_25831,N_20034,N_21448);
nor U25832 (N_25832,N_22834,N_24802);
xnor U25833 (N_25833,N_22945,N_23787);
nor U25834 (N_25834,N_22473,N_22851);
xnor U25835 (N_25835,N_20088,N_20771);
or U25836 (N_25836,N_22957,N_23634);
and U25837 (N_25837,N_20418,N_21173);
nand U25838 (N_25838,N_21650,N_21337);
or U25839 (N_25839,N_23182,N_20132);
xnor U25840 (N_25840,N_22055,N_24649);
or U25841 (N_25841,N_23051,N_23681);
xor U25842 (N_25842,N_24810,N_21902);
xor U25843 (N_25843,N_20657,N_21852);
and U25844 (N_25844,N_24163,N_22791);
or U25845 (N_25845,N_20780,N_24937);
xor U25846 (N_25846,N_20479,N_22467);
and U25847 (N_25847,N_23785,N_20321);
and U25848 (N_25848,N_22929,N_23284);
nand U25849 (N_25849,N_23968,N_24415);
or U25850 (N_25850,N_21806,N_24980);
or U25851 (N_25851,N_24958,N_23431);
xnor U25852 (N_25852,N_24411,N_23128);
and U25853 (N_25853,N_24996,N_20095);
or U25854 (N_25854,N_23293,N_23117);
nor U25855 (N_25855,N_20750,N_22045);
xnor U25856 (N_25856,N_21802,N_20455);
and U25857 (N_25857,N_21940,N_21128);
nor U25858 (N_25858,N_24189,N_22471);
or U25859 (N_25859,N_23514,N_24034);
and U25860 (N_25860,N_21819,N_22906);
nand U25861 (N_25861,N_20973,N_23777);
nor U25862 (N_25862,N_22145,N_23916);
nand U25863 (N_25863,N_22381,N_21422);
or U25864 (N_25864,N_23152,N_24329);
and U25865 (N_25865,N_21697,N_23366);
xor U25866 (N_25866,N_24346,N_23686);
and U25867 (N_25867,N_22628,N_23722);
or U25868 (N_25868,N_24363,N_21359);
xor U25869 (N_25869,N_21007,N_20718);
nand U25870 (N_25870,N_23837,N_24985);
nor U25871 (N_25871,N_21727,N_21316);
xnor U25872 (N_25872,N_23780,N_23554);
or U25873 (N_25873,N_22574,N_20866);
nor U25874 (N_25874,N_23370,N_22518);
and U25875 (N_25875,N_24203,N_20379);
and U25876 (N_25876,N_21370,N_22377);
and U25877 (N_25877,N_23528,N_24941);
xor U25878 (N_25878,N_21246,N_22745);
xor U25879 (N_25879,N_20127,N_22302);
nand U25880 (N_25880,N_23376,N_22267);
and U25881 (N_25881,N_24661,N_20580);
or U25882 (N_25882,N_21741,N_23952);
and U25883 (N_25883,N_24190,N_21384);
and U25884 (N_25884,N_23192,N_21656);
or U25885 (N_25885,N_22493,N_23857);
and U25886 (N_25886,N_22995,N_24688);
and U25887 (N_25887,N_20204,N_21547);
nor U25888 (N_25888,N_23946,N_22337);
or U25889 (N_25889,N_24439,N_23032);
nand U25890 (N_25890,N_23754,N_22144);
nor U25891 (N_25891,N_23113,N_24763);
or U25892 (N_25892,N_21794,N_22316);
xnor U25893 (N_25893,N_22556,N_20768);
nand U25894 (N_25894,N_21085,N_20730);
or U25895 (N_25895,N_22366,N_22756);
xnor U25896 (N_25896,N_24027,N_24207);
xnor U25897 (N_25897,N_23393,N_23757);
xor U25898 (N_25898,N_24121,N_23335);
or U25899 (N_25899,N_24345,N_21693);
and U25900 (N_25900,N_24904,N_21678);
nand U25901 (N_25901,N_20560,N_21307);
or U25902 (N_25902,N_20263,N_23320);
nand U25903 (N_25903,N_21708,N_22821);
xor U25904 (N_25904,N_22142,N_23383);
xnor U25905 (N_25905,N_21174,N_20197);
and U25906 (N_25906,N_21106,N_23202);
xnor U25907 (N_25907,N_21395,N_24210);
nor U25908 (N_25908,N_20102,N_24017);
and U25909 (N_25909,N_24118,N_24944);
and U25910 (N_25910,N_21149,N_21497);
xor U25911 (N_25911,N_20581,N_24878);
or U25912 (N_25912,N_20183,N_22274);
and U25913 (N_25913,N_24807,N_23572);
and U25914 (N_25914,N_23173,N_21788);
nor U25915 (N_25915,N_21700,N_20272);
and U25916 (N_25916,N_24000,N_20789);
xnor U25917 (N_25917,N_22307,N_22579);
nand U25918 (N_25918,N_24938,N_24975);
or U25919 (N_25919,N_21746,N_23653);
or U25920 (N_25920,N_23276,N_22992);
or U25921 (N_25921,N_22516,N_22009);
nor U25922 (N_25922,N_23986,N_22282);
nor U25923 (N_25923,N_23326,N_23906);
nand U25924 (N_25924,N_20840,N_23108);
nor U25925 (N_25925,N_23928,N_21120);
and U25926 (N_25926,N_23879,N_23098);
nand U25927 (N_25927,N_21154,N_24906);
nand U25928 (N_25928,N_22092,N_20618);
or U25929 (N_25929,N_22390,N_22637);
nand U25930 (N_25930,N_22005,N_23966);
xnor U25931 (N_25931,N_20812,N_21780);
xnor U25932 (N_25932,N_23718,N_21647);
or U25933 (N_25933,N_23533,N_22095);
xor U25934 (N_25934,N_20788,N_20186);
nor U25935 (N_25935,N_21360,N_22133);
and U25936 (N_25936,N_22624,N_24884);
nand U25937 (N_25937,N_21603,N_23866);
nand U25938 (N_25938,N_22515,N_24960);
and U25939 (N_25939,N_20676,N_23515);
nand U25940 (N_25940,N_23849,N_23510);
nand U25941 (N_25941,N_21188,N_20391);
xnor U25942 (N_25942,N_22150,N_20813);
or U25943 (N_25943,N_23672,N_23238);
xnor U25944 (N_25944,N_23652,N_24869);
or U25945 (N_25945,N_20665,N_24499);
xor U25946 (N_25946,N_22561,N_24936);
nor U25947 (N_25947,N_22169,N_22781);
nor U25948 (N_25948,N_20319,N_24476);
or U25949 (N_25949,N_22199,N_20967);
and U25950 (N_25950,N_21826,N_20119);
or U25951 (N_25951,N_21546,N_22948);
nor U25952 (N_25952,N_20363,N_20847);
nand U25953 (N_25953,N_20301,N_24722);
or U25954 (N_25954,N_24469,N_23410);
or U25955 (N_25955,N_23150,N_24265);
xnor U25956 (N_25956,N_21584,N_22635);
or U25957 (N_25957,N_23853,N_20700);
and U25958 (N_25958,N_22753,N_24577);
nor U25959 (N_25959,N_21542,N_20206);
nor U25960 (N_25960,N_24277,N_23120);
or U25961 (N_25961,N_21442,N_21371);
nand U25962 (N_25962,N_23530,N_22401);
and U25963 (N_25963,N_22431,N_23720);
and U25964 (N_25964,N_24068,N_22943);
and U25965 (N_25965,N_23290,N_24928);
nor U25966 (N_25966,N_20844,N_23909);
or U25967 (N_25967,N_24738,N_23771);
xnor U25968 (N_25968,N_24130,N_23097);
nand U25969 (N_25969,N_24250,N_22021);
nor U25970 (N_25970,N_23094,N_20153);
nor U25971 (N_25971,N_24629,N_24972);
xor U25972 (N_25972,N_20805,N_20041);
nand U25973 (N_25973,N_22173,N_24766);
xnor U25974 (N_25974,N_23501,N_21827);
xor U25975 (N_25975,N_22329,N_23810);
or U25976 (N_25976,N_24090,N_23901);
and U25977 (N_25977,N_22572,N_24378);
or U25978 (N_25978,N_21318,N_20990);
xnor U25979 (N_25979,N_21751,N_24898);
xor U25980 (N_25980,N_23611,N_24501);
nand U25981 (N_25981,N_20247,N_22090);
and U25982 (N_25982,N_23087,N_22193);
and U25983 (N_25983,N_24151,N_22901);
nand U25984 (N_25984,N_20265,N_24635);
or U25985 (N_25985,N_23650,N_22093);
and U25986 (N_25986,N_24864,N_21724);
and U25987 (N_25987,N_23132,N_23050);
and U25988 (N_25988,N_24322,N_24780);
xor U25989 (N_25989,N_22107,N_23888);
nand U25990 (N_25990,N_23876,N_20874);
nor U25991 (N_25991,N_22291,N_23491);
and U25992 (N_25992,N_23434,N_21035);
nor U25993 (N_25993,N_21257,N_24537);
xnor U25994 (N_25994,N_24992,N_22553);
or U25995 (N_25995,N_24104,N_22178);
nor U25996 (N_25996,N_22413,N_22110);
or U25997 (N_25997,N_21099,N_22779);
nor U25998 (N_25998,N_23260,N_23414);
nor U25999 (N_25999,N_21292,N_21508);
nor U26000 (N_26000,N_20624,N_22603);
xor U26001 (N_26001,N_20004,N_24169);
nor U26002 (N_26002,N_22692,N_23214);
xor U26003 (N_26003,N_24693,N_24035);
nor U26004 (N_26004,N_21633,N_21850);
xor U26005 (N_26005,N_20360,N_21324);
xor U26006 (N_26006,N_23965,N_22416);
or U26007 (N_26007,N_21170,N_22588);
nand U26008 (N_26008,N_21098,N_21280);
xnor U26009 (N_26009,N_21907,N_22375);
nand U26010 (N_26010,N_21585,N_22430);
nand U26011 (N_26011,N_22713,N_22121);
or U26012 (N_26012,N_21327,N_21380);
nand U26013 (N_26013,N_21964,N_21915);
nor U26014 (N_26014,N_20103,N_21415);
or U26015 (N_26015,N_24393,N_20187);
xor U26016 (N_26016,N_20879,N_24014);
nor U26017 (N_26017,N_23388,N_21031);
nor U26018 (N_26018,N_23872,N_20977);
and U26019 (N_26019,N_23425,N_21433);
nand U26020 (N_26020,N_24675,N_22321);
or U26021 (N_26021,N_21002,N_23578);
nand U26022 (N_26022,N_22942,N_24114);
and U26023 (N_26023,N_20292,N_21843);
and U26024 (N_26024,N_22654,N_22858);
nor U26025 (N_26025,N_24753,N_22482);
xnor U26026 (N_26026,N_21664,N_21261);
nand U26027 (N_26027,N_22738,N_24144);
nor U26028 (N_26028,N_24434,N_23005);
xnor U26029 (N_26029,N_24861,N_20919);
nor U26030 (N_26030,N_21287,N_20514);
xnor U26031 (N_26031,N_22428,N_24801);
and U26032 (N_26032,N_20448,N_24961);
or U26033 (N_26033,N_24647,N_20268);
nor U26034 (N_26034,N_21495,N_21666);
or U26035 (N_26035,N_23983,N_24041);
or U26036 (N_26036,N_22814,N_21531);
nor U26037 (N_26037,N_22119,N_23537);
and U26038 (N_26038,N_23207,N_21339);
nand U26039 (N_26039,N_20210,N_21966);
nand U26040 (N_26040,N_24950,N_24720);
nor U26041 (N_26041,N_22259,N_22673);
or U26042 (N_26042,N_22767,N_20084);
and U26043 (N_26043,N_20042,N_24246);
and U26044 (N_26044,N_20929,N_20199);
and U26045 (N_26045,N_20316,N_24816);
xor U26046 (N_26046,N_24098,N_23704);
nand U26047 (N_26047,N_21250,N_21103);
nor U26048 (N_26048,N_24195,N_22368);
nor U26049 (N_26049,N_21607,N_20772);
nand U26050 (N_26050,N_21302,N_20428);
nand U26051 (N_26051,N_23999,N_22386);
nor U26052 (N_26052,N_20746,N_21449);
and U26053 (N_26053,N_23309,N_23752);
nand U26054 (N_26054,N_21762,N_23956);
and U26055 (N_26055,N_21541,N_23967);
xnor U26056 (N_26056,N_24011,N_21929);
and U26057 (N_26057,N_24643,N_24458);
xnor U26058 (N_26058,N_23445,N_23656);
nor U26059 (N_26059,N_22179,N_24253);
nor U26060 (N_26060,N_20876,N_22099);
and U26061 (N_26061,N_20589,N_24053);
nor U26062 (N_26062,N_20036,N_23744);
and U26063 (N_26063,N_23727,N_23443);
xor U26064 (N_26064,N_21729,N_20383);
nand U26065 (N_26065,N_23671,N_23001);
xnor U26066 (N_26066,N_24978,N_22197);
xnor U26067 (N_26067,N_22559,N_22527);
xor U26068 (N_26068,N_20432,N_22768);
or U26069 (N_26069,N_20677,N_20857);
or U26070 (N_26070,N_24245,N_20566);
nand U26071 (N_26071,N_22695,N_20518);
or U26072 (N_26072,N_22207,N_20425);
xnor U26073 (N_26073,N_24800,N_23233);
or U26074 (N_26074,N_20076,N_24734);
xnor U26075 (N_26075,N_22124,N_23060);
nor U26076 (N_26076,N_21114,N_23042);
nand U26077 (N_26077,N_20608,N_20504);
nor U26078 (N_26078,N_23143,N_23954);
or U26079 (N_26079,N_23271,N_22270);
and U26080 (N_26080,N_22848,N_23413);
xnor U26081 (N_26081,N_22610,N_21522);
nor U26082 (N_26082,N_24153,N_21564);
xor U26083 (N_26083,N_21062,N_24642);
nand U26084 (N_26084,N_23855,N_23590);
nor U26085 (N_26085,N_22682,N_23245);
nand U26086 (N_26086,N_23759,N_21658);
nor U26087 (N_26087,N_22306,N_22643);
xnor U26088 (N_26088,N_24129,N_21989);
nand U26089 (N_26089,N_20362,N_20830);
xor U26090 (N_26090,N_24651,N_21714);
and U26091 (N_26091,N_21323,N_21293);
xnor U26092 (N_26092,N_22171,N_24637);
xnor U26093 (N_26093,N_22839,N_24927);
and U26094 (N_26094,N_20423,N_20224);
nand U26095 (N_26095,N_22129,N_22720);
and U26096 (N_26096,N_24009,N_23897);
and U26097 (N_26097,N_21233,N_23355);
nand U26098 (N_26098,N_24217,N_24325);
xnor U26099 (N_26099,N_20044,N_22174);
nor U26100 (N_26100,N_22300,N_21616);
nor U26101 (N_26101,N_20766,N_21212);
or U26102 (N_26102,N_23882,N_20671);
nor U26103 (N_26103,N_23535,N_20176);
or U26104 (N_26104,N_23286,N_24619);
nand U26105 (N_26105,N_23839,N_23341);
nand U26106 (N_26106,N_22583,N_23516);
nor U26107 (N_26107,N_21317,N_22359);
and U26108 (N_26108,N_23244,N_24269);
and U26109 (N_26109,N_22763,N_23755);
nand U26110 (N_26110,N_23820,N_22244);
or U26111 (N_26111,N_21660,N_22889);
and U26112 (N_26112,N_22951,N_20783);
or U26113 (N_26113,N_24425,N_21718);
and U26114 (N_26114,N_23910,N_21443);
nor U26115 (N_26115,N_21925,N_22249);
nand U26116 (N_26116,N_21860,N_20166);
or U26117 (N_26117,N_22385,N_22230);
and U26118 (N_26118,N_21383,N_22650);
nor U26119 (N_26119,N_20063,N_23036);
or U26120 (N_26120,N_21837,N_24543);
nand U26121 (N_26121,N_20038,N_20717);
and U26122 (N_26122,N_24223,N_22883);
nor U26123 (N_26123,N_23035,N_20090);
nand U26124 (N_26124,N_21138,N_24453);
and U26125 (N_26125,N_24417,N_24873);
and U26126 (N_26126,N_24465,N_24047);
xor U26127 (N_26127,N_22488,N_21696);
nand U26128 (N_26128,N_24450,N_22577);
xnor U26129 (N_26129,N_22056,N_23399);
or U26130 (N_26130,N_24730,N_23945);
xor U26131 (N_26131,N_20307,N_20196);
nand U26132 (N_26132,N_24452,N_21306);
nand U26133 (N_26133,N_20317,N_20683);
nand U26134 (N_26134,N_24733,N_23012);
or U26135 (N_26135,N_22743,N_23663);
nor U26136 (N_26136,N_21435,N_23201);
xnor U26137 (N_26137,N_24304,N_21862);
nand U26138 (N_26138,N_21217,N_21791);
or U26139 (N_26139,N_22452,N_24628);
nor U26140 (N_26140,N_22669,N_21975);
and U26141 (N_26141,N_24778,N_24165);
xnor U26142 (N_26142,N_22675,N_23721);
or U26143 (N_26143,N_23381,N_24154);
and U26144 (N_26144,N_20472,N_21502);
xor U26145 (N_26145,N_23007,N_24627);
or U26146 (N_26146,N_23203,N_24779);
and U26147 (N_26147,N_20763,N_20381);
nand U26148 (N_26148,N_20101,N_22933);
and U26149 (N_26149,N_24723,N_20136);
xor U26150 (N_26150,N_21859,N_24107);
and U26151 (N_26151,N_21740,N_22818);
nand U26152 (N_26152,N_24606,N_23482);
nor U26153 (N_26153,N_24032,N_23657);
nand U26154 (N_26154,N_20869,N_24982);
xor U26155 (N_26155,N_22794,N_23942);
nor U26156 (N_26156,N_23116,N_24609);
nand U26157 (N_26157,N_22344,N_20948);
nand U26158 (N_26158,N_23543,N_23864);
or U26159 (N_26159,N_20105,N_20201);
xnor U26160 (N_26160,N_21573,N_21115);
nand U26161 (N_26161,N_20311,N_22548);
or U26162 (N_26162,N_20800,N_24475);
xor U26163 (N_26163,N_24700,N_22394);
xnor U26164 (N_26164,N_20463,N_20834);
or U26165 (N_26165,N_20139,N_23753);
xor U26166 (N_26166,N_21159,N_20445);
xor U26167 (N_26167,N_21755,N_22010);
and U26168 (N_26168,N_22043,N_23723);
nor U26169 (N_26169,N_21968,N_21245);
xor U26170 (N_26170,N_20083,N_22036);
and U26171 (N_26171,N_20134,N_21135);
or U26172 (N_26172,N_21877,N_24036);
nand U26173 (N_26173,N_23756,N_23239);
nand U26174 (N_26174,N_20541,N_21828);
nand U26175 (N_26175,N_20962,N_20538);
xor U26176 (N_26176,N_22840,N_20241);
nand U26177 (N_26177,N_23240,N_22638);
and U26178 (N_26178,N_21959,N_22283);
nand U26179 (N_26179,N_24480,N_20897);
and U26180 (N_26180,N_21928,N_20053);
or U26181 (N_26181,N_22065,N_22508);
and U26182 (N_26182,N_22905,N_21057);
xnor U26183 (N_26183,N_24886,N_23848);
and U26184 (N_26184,N_20769,N_21358);
or U26185 (N_26185,N_23569,N_20030);
nand U26186 (N_26186,N_21163,N_23852);
nor U26187 (N_26187,N_24468,N_24297);
and U26188 (N_26188,N_24242,N_21126);
and U26189 (N_26189,N_20917,N_24124);
xor U26190 (N_26190,N_20670,N_23226);
or U26191 (N_26191,N_20628,N_24192);
xnor U26192 (N_26192,N_20918,N_21669);
nor U26193 (N_26193,N_22864,N_23521);
xor U26194 (N_26194,N_21753,N_21496);
xor U26195 (N_26195,N_23884,N_20408);
nor U26196 (N_26196,N_23262,N_24731);
and U26197 (N_26197,N_21229,N_23571);
and U26198 (N_26198,N_20157,N_23279);
nor U26199 (N_26199,N_24146,N_20762);
and U26200 (N_26200,N_21286,N_23640);
nand U26201 (N_26201,N_22573,N_24257);
and U26202 (N_26202,N_23291,N_21169);
nand U26203 (N_26203,N_20120,N_22323);
or U26204 (N_26204,N_22391,N_23801);
and U26205 (N_26205,N_22877,N_24924);
nand U26206 (N_26206,N_23168,N_24460);
or U26207 (N_26207,N_24262,N_23074);
xnor U26208 (N_26208,N_24895,N_23764);
xor U26209 (N_26209,N_20192,N_22407);
or U26210 (N_26210,N_24149,N_22131);
xor U26211 (N_26211,N_20854,N_24947);
and U26212 (N_26212,N_21234,N_21821);
nor U26213 (N_26213,N_24020,N_20852);
nor U26214 (N_26214,N_21451,N_21214);
xor U26215 (N_26215,N_20299,N_23344);
nand U26216 (N_26216,N_21069,N_23295);
and U26217 (N_26217,N_22549,N_21822);
or U26218 (N_26218,N_21970,N_21804);
and U26219 (N_26219,N_22355,N_21249);
and U26220 (N_26220,N_22489,N_20956);
or U26221 (N_26221,N_24352,N_20473);
nor U26222 (N_26222,N_24858,N_21994);
xnor U26223 (N_26223,N_24888,N_20446);
xor U26224 (N_26224,N_20279,N_24119);
and U26225 (N_26225,N_21426,N_21139);
nand U26226 (N_26226,N_21632,N_23232);
and U26227 (N_26227,N_23984,N_21792);
xnor U26228 (N_26228,N_23636,N_22126);
or U26229 (N_26229,N_21950,N_23364);
nand U26230 (N_26230,N_20417,N_23766);
nor U26231 (N_26231,N_22213,N_24690);
and U26232 (N_26232,N_21922,N_21685);
xnor U26233 (N_26233,N_23251,N_22408);
xnor U26234 (N_26234,N_23481,N_22125);
nor U26235 (N_26235,N_22163,N_22258);
or U26236 (N_26236,N_21044,N_21311);
or U26237 (N_26237,N_21288,N_21935);
and U26238 (N_26238,N_22070,N_24829);
nand U26239 (N_26239,N_20222,N_24908);
or U26240 (N_26240,N_23404,N_20784);
nor U26241 (N_26241,N_24087,N_21610);
nor U26242 (N_26242,N_22709,N_22525);
xor U26243 (N_26243,N_22706,N_24341);
or U26244 (N_26244,N_23788,N_23498);
xnor U26245 (N_26245,N_22685,N_24512);
xor U26246 (N_26246,N_23896,N_20113);
or U26247 (N_26247,N_23825,N_24234);
xor U26248 (N_26248,N_22216,N_20528);
nand U26249 (N_26249,N_21314,N_21817);
nand U26250 (N_26250,N_23941,N_22721);
xor U26251 (N_26251,N_21461,N_23736);
xor U26252 (N_26252,N_21676,N_20751);
xnor U26253 (N_26253,N_22086,N_20068);
nand U26254 (N_26254,N_23137,N_20662);
nand U26255 (N_26255,N_24067,N_24589);
nor U26256 (N_26256,N_20303,N_24288);
nand U26257 (N_26257,N_22866,N_22907);
or U26258 (N_26258,N_21628,N_24879);
nand U26259 (N_26259,N_22766,N_21640);
or U26260 (N_26260,N_20519,N_23085);
nor U26261 (N_26261,N_20622,N_24001);
nor U26262 (N_26262,N_20229,N_20711);
nor U26263 (N_26263,N_22897,N_20991);
xor U26264 (N_26264,N_22372,N_23937);
or U26265 (N_26265,N_20713,N_20868);
or U26266 (N_26266,N_23157,N_22343);
nand U26267 (N_26267,N_20862,N_22403);
nand U26268 (N_26268,N_24917,N_24477);
nand U26269 (N_26269,N_21515,N_24524);
nor U26270 (N_26270,N_24387,N_21831);
nand U26271 (N_26271,N_22831,N_24760);
or U26272 (N_26272,N_24193,N_21266);
xor U26273 (N_26273,N_24644,N_22331);
nor U26274 (N_26274,N_21883,N_21278);
and U26275 (N_26275,N_22930,N_20082);
xor U26276 (N_26276,N_24386,N_20960);
xnor U26277 (N_26277,N_24385,N_21949);
xor U26278 (N_26278,N_21076,N_24549);
and U26279 (N_26279,N_21615,N_20837);
nand U26280 (N_26280,N_21320,N_21326);
xor U26281 (N_26281,N_24426,N_23596);
or U26282 (N_26282,N_21690,N_22979);
or U26283 (N_26283,N_22203,N_24655);
nor U26284 (N_26284,N_20650,N_20843);
and U26285 (N_26285,N_20889,N_20690);
xnor U26286 (N_26286,N_22198,N_22012);
nor U26287 (N_26287,N_21191,N_23397);
and U26288 (N_26288,N_21703,N_20261);
nor U26289 (N_26289,N_21734,N_20535);
nor U26290 (N_26290,N_20022,N_22813);
or U26291 (N_26291,N_22728,N_20555);
nor U26292 (N_26292,N_23568,N_22164);
or U26293 (N_26293,N_24962,N_21494);
or U26294 (N_26294,N_24799,N_22118);
and U26295 (N_26295,N_24167,N_22750);
and U26296 (N_26296,N_21818,N_21567);
or U26297 (N_26297,N_21456,N_21136);
and U26298 (N_26298,N_21213,N_24010);
nor U26299 (N_26299,N_20451,N_22435);
and U26300 (N_26300,N_23699,N_24756);
or U26301 (N_26301,N_23174,N_23474);
xor U26302 (N_26302,N_20699,N_23739);
or U26303 (N_26303,N_22481,N_21655);
nor U26304 (N_26304,N_21763,N_21927);
or U26305 (N_26305,N_20995,N_20938);
and U26306 (N_26306,N_20653,N_21533);
and U26307 (N_26307,N_23524,N_22470);
nand U26308 (N_26308,N_20831,N_20327);
nand U26309 (N_26309,N_21171,N_24919);
xnor U26310 (N_26310,N_20228,N_23078);
and U26311 (N_26311,N_21719,N_21446);
xor U26312 (N_26312,N_22500,N_21958);
nor U26313 (N_26313,N_24610,N_23459);
nand U26314 (N_26314,N_23004,N_24728);
and U26315 (N_26315,N_24929,N_23266);
or U26316 (N_26316,N_23927,N_20965);
and U26317 (N_26317,N_21235,N_24445);
nand U26318 (N_26318,N_21715,N_24667);
and U26319 (N_26319,N_20755,N_23817);
and U26320 (N_26320,N_23975,N_22614);
xor U26321 (N_26321,N_24233,N_22714);
nand U26322 (N_26322,N_24594,N_22544);
or U26323 (N_26323,N_24092,N_22916);
xnor U26324 (N_26324,N_22862,N_23318);
nor U26325 (N_26325,N_24830,N_21993);
nor U26326 (N_26326,N_20128,N_20635);
nand U26327 (N_26327,N_23808,N_24718);
xnor U26328 (N_26328,N_20716,N_24668);
nor U26329 (N_26329,N_21051,N_21385);
nor U26330 (N_26330,N_21652,N_20688);
nand U26331 (N_26331,N_21453,N_23496);
and U26332 (N_26332,N_20633,N_21726);
nor U26333 (N_26333,N_24573,N_20374);
and U26334 (N_26334,N_23466,N_23637);
and U26335 (N_26335,N_22141,N_21517);
and U26336 (N_26336,N_23373,N_20524);
nor U26337 (N_26337,N_22727,N_21222);
nor U26338 (N_26338,N_23767,N_20250);
and U26339 (N_26339,N_22167,N_23248);
nor U26340 (N_26340,N_23904,N_24732);
nand U26341 (N_26341,N_20899,N_21529);
xor U26342 (N_26342,N_24308,N_23536);
or U26343 (N_26343,N_23778,N_20433);
and U26344 (N_26344,N_21203,N_24289);
nor U26345 (N_26345,N_22204,N_20151);
nand U26346 (N_26346,N_24966,N_21937);
xnor U26347 (N_26347,N_24389,N_23765);
and U26348 (N_26348,N_24055,N_21134);
and U26349 (N_26349,N_20588,N_24520);
xor U26350 (N_26350,N_23455,N_21177);
or U26351 (N_26351,N_21984,N_21315);
and U26352 (N_26352,N_21368,N_21423);
nand U26353 (N_26353,N_20801,N_21933);
nand U26354 (N_26354,N_24464,N_24580);
and U26355 (N_26355,N_20194,N_21350);
nor U26356 (N_26356,N_22656,N_23570);
or U26357 (N_26357,N_23931,N_20826);
xor U26358 (N_26358,N_24857,N_22671);
xnor U26359 (N_26359,N_21673,N_23796);
nor U26360 (N_26360,N_22592,N_23794);
and U26361 (N_26361,N_24401,N_23197);
nand U26362 (N_26362,N_20329,N_23588);
nand U26363 (N_26363,N_24038,N_20606);
and U26364 (N_26364,N_23054,N_24235);
nor U26365 (N_26365,N_21281,N_20957);
xnor U26366 (N_26366,N_23179,N_20375);
and U26367 (N_26367,N_20759,N_22376);
nor U26368 (N_26368,N_22691,N_21416);
xnor U26369 (N_26369,N_21239,N_23264);
nand U26370 (N_26370,N_24743,N_23761);
xnor U26371 (N_26371,N_24658,N_23953);
xnor U26372 (N_26372,N_22723,N_20300);
xor U26373 (N_26373,N_22737,N_22011);
nor U26374 (N_26374,N_23819,N_20270);
and U26375 (N_26375,N_23556,N_23784);
and U26376 (N_26376,N_24672,N_21127);
or U26377 (N_26377,N_21480,N_22450);
xnor U26378 (N_26378,N_24663,N_21764);
and U26379 (N_26379,N_22797,N_22824);
xnor U26380 (N_26380,N_21596,N_20696);
or U26381 (N_26381,N_22975,N_22490);
or U26382 (N_26382,N_20231,N_24132);
or U26383 (N_26383,N_23217,N_23118);
xnor U26384 (N_26384,N_24602,N_23598);
nor U26385 (N_26385,N_22425,N_23505);
or U26386 (N_26386,N_20045,N_23520);
or U26387 (N_26387,N_23218,N_21705);
nand U26388 (N_26388,N_22993,N_22880);
nor U26389 (N_26389,N_24925,N_21516);
and U26390 (N_26390,N_23440,N_22279);
and U26391 (N_26391,N_23044,N_22271);
or U26392 (N_26392,N_21021,N_23660);
or U26393 (N_26393,N_20927,N_22822);
nor U26394 (N_26394,N_21096,N_22361);
nand U26395 (N_26395,N_21056,N_23255);
or U26396 (N_26396,N_23748,N_21095);
xor U26397 (N_26397,N_21861,N_20584);
xnor U26398 (N_26398,N_23862,N_23417);
xnor U26399 (N_26399,N_23547,N_22383);
or U26400 (N_26400,N_21520,N_21325);
nor U26401 (N_26401,N_23605,N_20060);
or U26402 (N_26402,N_24155,N_24002);
nor U26403 (N_26403,N_20660,N_21109);
and U26404 (N_26404,N_23436,N_23802);
nand U26405 (N_26405,N_23385,N_20851);
xnor U26406 (N_26406,N_20725,N_21408);
and U26407 (N_26407,N_21329,N_23905);
or U26408 (N_26408,N_21192,N_23209);
and U26409 (N_26409,N_22808,N_22602);
or U26410 (N_26410,N_23029,N_20207);
nor U26411 (N_26411,N_22689,N_21201);
nand U26412 (N_26412,N_21576,N_21130);
and U26413 (N_26413,N_24116,N_20107);
and U26414 (N_26414,N_21896,N_23833);
or U26415 (N_26415,N_24073,N_22939);
nand U26416 (N_26416,N_22742,N_23017);
xor U26417 (N_26417,N_21276,N_22185);
nor U26418 (N_26418,N_21833,N_21589);
and U26419 (N_26419,N_23040,N_22214);
nor U26420 (N_26420,N_23296,N_22777);
and U26421 (N_26421,N_24226,N_21680);
and U26422 (N_26422,N_21816,N_21934);
nor U26423 (N_26423,N_21518,N_22647);
and U26424 (N_26424,N_21663,N_23615);
or U26425 (N_26425,N_23357,N_20632);
xnor U26426 (N_26426,N_21332,N_22538);
and U26427 (N_26427,N_21768,N_21078);
nand U26428 (N_26428,N_21878,N_21750);
xnor U26429 (N_26429,N_21681,N_21598);
or U26430 (N_26430,N_20150,N_24890);
and U26431 (N_26431,N_21648,N_20302);
nand U26432 (N_26432,N_24691,N_22228);
nand U26433 (N_26433,N_20687,N_23579);
nor U26434 (N_26434,N_22426,N_22981);
xor U26435 (N_26435,N_21020,N_22989);
xnor U26436 (N_26436,N_20348,N_23776);
nor U26437 (N_26437,N_24268,N_22158);
and U26438 (N_26438,N_23725,N_24019);
nor U26439 (N_26439,N_21018,N_21722);
or U26440 (N_26440,N_24983,N_24735);
and U26441 (N_26441,N_24748,N_21960);
nand U26442 (N_26442,N_22563,N_22519);
xnor U26443 (N_26443,N_20427,N_22963);
nor U26444 (N_26444,N_23423,N_20795);
nor U26445 (N_26445,N_22294,N_22748);
xnor U26446 (N_26446,N_23163,N_23391);
or U26447 (N_26447,N_23172,N_23331);
or U26448 (N_26448,N_23371,N_22783);
or U26449 (N_26449,N_23540,N_22504);
nand U26450 (N_26450,N_24140,N_22025);
nand U26451 (N_26451,N_21793,N_20998);
or U26452 (N_26452,N_23334,N_21604);
xnor U26453 (N_26453,N_21219,N_20488);
nand U26454 (N_26454,N_23559,N_20234);
xnor U26455 (N_26455,N_20570,N_21176);
and U26456 (N_26456,N_20886,N_22202);
and U26457 (N_26457,N_23740,N_23875);
or U26458 (N_26458,N_22524,N_21504);
or U26459 (N_26459,N_23741,N_23337);
xnor U26460 (N_26460,N_23028,N_23883);
nand U26461 (N_26461,N_21077,N_22245);
nand U26462 (N_26462,N_23299,N_23103);
or U26463 (N_26463,N_22089,N_24403);
nand U26464 (N_26464,N_22956,N_24168);
or U26465 (N_26465,N_20352,N_21839);
xor U26466 (N_26466,N_22353,N_21712);
nor U26467 (N_26467,N_21379,N_24420);
nor U26468 (N_26468,N_22395,N_23478);
and U26469 (N_26469,N_22149,N_23618);
nand U26470 (N_26470,N_24405,N_20495);
nor U26471 (N_26471,N_20739,N_24574);
nor U26472 (N_26472,N_22711,N_21730);
nand U26473 (N_26473,N_20456,N_20963);
or U26474 (N_26474,N_20251,N_22154);
nand U26475 (N_26475,N_21086,N_24503);
or U26476 (N_26476,N_24526,N_20757);
and U26477 (N_26477,N_22664,N_21066);
or U26478 (N_26478,N_21748,N_24836);
nor U26479 (N_26479,N_20243,N_21620);
and U26480 (N_26480,N_23280,N_21998);
or U26481 (N_26481,N_24459,N_24162);
nor U26482 (N_26482,N_24578,N_21682);
or U26483 (N_26483,N_24533,N_20590);
nor U26484 (N_26484,N_20032,N_22295);
or U26485 (N_26485,N_22001,N_20147);
xor U26486 (N_26486,N_22632,N_20839);
and U26487 (N_26487,N_21691,N_20274);
and U26488 (N_26488,N_20527,N_23071);
nor U26489 (N_26489,N_21392,N_20542);
or U26490 (N_26490,N_21521,N_24823);
and U26491 (N_26491,N_20643,N_23651);
nand U26492 (N_26492,N_22944,N_21429);
nand U26493 (N_26493,N_23189,N_23476);
xnor U26494 (N_26494,N_23274,N_22582);
or U26495 (N_26495,N_24859,N_24682);
nand U26496 (N_26496,N_22397,N_20644);
nand U26497 (N_26497,N_24202,N_22667);
or U26498 (N_26498,N_23745,N_20443);
nand U26499 (N_26499,N_21553,N_22715);
and U26500 (N_26500,N_24454,N_20493);
xnor U26501 (N_26501,N_22806,N_23470);
and U26502 (N_26502,N_22137,N_22189);
nand U26503 (N_26503,N_22071,N_24541);
nor U26504 (N_26504,N_20679,N_23608);
nor U26505 (N_26505,N_21626,N_20140);
nor U26506 (N_26506,N_24509,N_20836);
xor U26507 (N_26507,N_24593,N_24525);
nand U26508 (N_26508,N_23877,N_23751);
nor U26509 (N_26509,N_23162,N_24173);
nand U26510 (N_26510,N_22272,N_22406);
nand U26511 (N_26511,N_24364,N_21644);
and U26512 (N_26512,N_21857,N_21347);
or U26513 (N_26513,N_20245,N_22676);
or U26514 (N_26514,N_22881,N_23620);
nor U26515 (N_26515,N_23099,N_23943);
or U26516 (N_26516,N_21982,N_20159);
and U26517 (N_26517,N_24741,N_21472);
xor U26518 (N_26518,N_21836,N_20478);
and U26519 (N_26519,N_23249,N_23566);
xor U26520 (N_26520,N_20969,N_20786);
or U26521 (N_26521,N_24259,N_22616);
or U26522 (N_26522,N_23489,N_24648);
nand U26523 (N_26523,N_23662,N_22073);
or U26524 (N_26524,N_24703,N_24440);
xor U26525 (N_26525,N_21789,N_23241);
nand U26526 (N_26526,N_20282,N_21470);
xor U26527 (N_26527,N_20104,N_23064);
or U26528 (N_26528,N_22182,N_22860);
nor U26529 (N_26529,N_22484,N_20035);
and U26530 (N_26530,N_24292,N_24514);
and U26531 (N_26531,N_24554,N_21781);
and U26532 (N_26532,N_23987,N_21129);
xnor U26533 (N_26533,N_24953,N_23940);
or U26534 (N_26534,N_23585,N_22346);
or U26535 (N_26535,N_21072,N_23851);
and U26536 (N_26536,N_23138,N_21049);
nand U26537 (N_26537,N_22340,N_20974);
nand U26538 (N_26538,N_22177,N_20569);
or U26539 (N_26539,N_22799,N_22112);
nand U26540 (N_26540,N_20017,N_20019);
nand U26541 (N_26541,N_22918,N_24326);
or U26542 (N_26542,N_20123,N_20659);
xor U26543 (N_26543,N_24518,N_22047);
nor U26544 (N_26544,N_24443,N_22784);
or U26545 (N_26545,N_24783,N_21823);
nor U26546 (N_26546,N_23061,N_21886);
or U26547 (N_26547,N_23038,N_21600);
xnor U26548 (N_26548,N_24113,N_22876);
nand U26549 (N_26549,N_20536,N_23321);
nand U26550 (N_26550,N_21599,N_20667);
and U26551 (N_26551,N_21728,N_20733);
xnor U26552 (N_26552,N_23538,N_24494);
or U26553 (N_26553,N_20158,N_20742);
nor U26554 (N_26554,N_24555,N_23828);
and U26555 (N_26555,N_24598,N_21375);
nor U26556 (N_26556,N_21207,N_21562);
nor U26557 (N_26557,N_23816,N_24355);
and U26558 (N_26558,N_23342,N_20547);
xor U26559 (N_26559,N_20737,N_24447);
or U26560 (N_26560,N_20420,N_20371);
and U26561 (N_26561,N_20429,N_22687);
nor U26562 (N_26562,N_22215,N_24974);
or U26563 (N_26563,N_23253,N_22338);
or U26564 (N_26564,N_24707,N_22890);
and U26565 (N_26565,N_23386,N_23193);
xor U26566 (N_26566,N_20226,N_24408);
and U26567 (N_26567,N_22241,N_23229);
or U26568 (N_26568,N_22345,N_23575);
xor U26569 (N_26569,N_21270,N_24351);
nand U26570 (N_26570,N_21894,N_21401);
nand U26571 (N_26571,N_20001,N_22352);
and U26572 (N_26572,N_24240,N_23122);
nand U26573 (N_26573,N_22609,N_24542);
and U26574 (N_26574,N_23289,N_22019);
or U26575 (N_26575,N_21404,N_23034);
xor U26576 (N_26576,N_22260,N_21405);
or U26577 (N_26577,N_23130,N_23056);
xnor U26578 (N_26578,N_21798,N_22015);
nand U26579 (N_26579,N_24516,N_22751);
nand U26580 (N_26580,N_23919,N_24089);
or U26581 (N_26581,N_24681,N_24772);
nand U26582 (N_26582,N_20291,N_24725);
or U26583 (N_26583,N_24670,N_20264);
xnor U26584 (N_26584,N_22497,N_22459);
or U26585 (N_26585,N_23460,N_21969);
or U26586 (N_26586,N_20458,N_22136);
or U26587 (N_26587,N_24828,N_24272);
xor U26588 (N_26588,N_22555,N_23546);
or U26589 (N_26589,N_20748,N_20308);
xor U26590 (N_26590,N_21556,N_22495);
xnor U26591 (N_26591,N_24636,N_24344);
or U26592 (N_26592,N_24142,N_24315);
nand U26593 (N_26593,N_22460,N_22887);
nand U26594 (N_26594,N_24206,N_23198);
or U26595 (N_26595,N_20803,N_21774);
nor U26596 (N_26596,N_20993,N_21895);
or U26597 (N_26597,N_22156,N_21122);
nand U26598 (N_26598,N_20238,N_22725);
or U26599 (N_26599,N_24930,N_24451);
or U26600 (N_26600,N_21232,N_21848);
or U26601 (N_26601,N_23303,N_22700);
and U26602 (N_26602,N_20000,N_20599);
nor U26603 (N_26603,N_23070,N_20715);
nor U26604 (N_26604,N_21686,N_23936);
xnor U26605 (N_26605,N_22077,N_22322);
or U26606 (N_26606,N_22315,N_24232);
and U26607 (N_26607,N_20046,N_23052);
and U26608 (N_26608,N_23991,N_24267);
nor U26609 (N_26609,N_20266,N_22926);
xor U26610 (N_26610,N_20949,N_23858);
xnor U26611 (N_26611,N_21244,N_22046);
and U26612 (N_26612,N_20966,N_20985);
xor U26613 (N_26613,N_22875,N_24564);
nor U26614 (N_26614,N_21606,N_20310);
nand U26615 (N_26615,N_24323,N_22801);
nand U26616 (N_26616,N_23622,N_20777);
or U26617 (N_26617,N_21899,N_23415);
or U26618 (N_26618,N_24320,N_21642);
and U26619 (N_26619,N_22441,N_24692);
nand U26620 (N_26620,N_23180,N_21464);
xor U26621 (N_26621,N_22634,N_23593);
nor U26622 (N_26622,N_24102,N_22569);
and U26623 (N_26623,N_24491,N_21172);
and U26624 (N_26624,N_20441,N_21019);
and U26625 (N_26625,N_23453,N_23426);
and U26626 (N_26626,N_24712,N_24012);
xor U26627 (N_26627,N_20005,N_23412);
or U26628 (N_26628,N_20131,N_21215);
xor U26629 (N_26629,N_22629,N_20275);
nor U26630 (N_26630,N_22275,N_24500);
nand U26631 (N_26631,N_23367,N_20835);
nand U26632 (N_26632,N_23706,N_21023);
nor U26633 (N_26633,N_24640,N_23362);
and U26634 (N_26634,N_20356,N_24584);
nand U26635 (N_26635,N_24057,N_23057);
xnor U26636 (N_26636,N_20078,N_24531);
xor U26637 (N_26637,N_24160,N_20556);
nand U26638 (N_26638,N_22370,N_21569);
xor U26639 (N_26639,N_21112,N_24079);
or U26640 (N_26640,N_23246,N_20930);
and U26641 (N_26641,N_24497,N_20477);
and U26642 (N_26642,N_21411,N_24075);
nor U26643 (N_26643,N_24989,N_20296);
and U26644 (N_26644,N_20603,N_24302);
and U26645 (N_26645,N_23312,N_20057);
and U26646 (N_26646,N_22362,N_21671);
nor U26647 (N_26647,N_21956,N_21778);
nand U26648 (N_26648,N_24794,N_22072);
or U26649 (N_26649,N_21053,N_23323);
and U26650 (N_26650,N_20698,N_21910);
xor U26651 (N_26651,N_24093,N_22702);
nand U26652 (N_26652,N_23349,N_20334);
or U26653 (N_26653,N_22292,N_20975);
or U26654 (N_26654,N_22999,N_21196);
nand U26655 (N_26655,N_20530,N_24811);
nand U26656 (N_26656,N_23711,N_20501);
and U26657 (N_26657,N_23834,N_23500);
or U26658 (N_26658,N_21400,N_23562);
xor U26659 (N_26659,N_23358,N_23058);
nand U26660 (N_26660,N_23356,N_24599);
and U26661 (N_26661,N_21295,N_20512);
or U26662 (N_26662,N_21637,N_22567);
xor U26663 (N_26663,N_20439,N_20173);
nand U26664 (N_26664,N_24674,N_21549);
xnor U26665 (N_26665,N_20115,N_21068);
and U26666 (N_26666,N_21029,N_22003);
or U26667 (N_26667,N_21362,N_20118);
xnor U26668 (N_26668,N_21025,N_22423);
or U26669 (N_26669,N_24466,N_21511);
nand U26670 (N_26670,N_24028,N_24042);
nor U26671 (N_26671,N_22955,N_24519);
or U26672 (N_26672,N_24893,N_20860);
or U26673 (N_26673,N_24406,N_22805);
or U26674 (N_26674,N_22657,N_22269);
and U26675 (N_26675,N_20563,N_23449);
nor U26676 (N_26676,N_22965,N_24383);
xnor U26677 (N_26677,N_23140,N_22235);
nor U26678 (N_26678,N_24314,N_24942);
nor U26679 (N_26679,N_24495,N_22920);
nor U26680 (N_26680,N_20856,N_20842);
and U26681 (N_26681,N_23479,N_20322);
nor U26682 (N_26682,N_23016,N_22505);
nor U26683 (N_26683,N_22236,N_20277);
nand U26684 (N_26684,N_21407,N_22192);
nor U26685 (N_26685,N_23668,N_22672);
nor U26686 (N_26686,N_23529,N_23665);
nand U26687 (N_26687,N_22514,N_24112);
or U26688 (N_26688,N_22990,N_22041);
nand U26689 (N_26689,N_24435,N_20596);
xor U26690 (N_26690,N_23250,N_23823);
or U26691 (N_26691,N_23868,N_20576);
and U26692 (N_26692,N_22052,N_24137);
nor U26693 (N_26693,N_20305,N_24591);
nand U26694 (N_26694,N_22974,N_22058);
xor U26695 (N_26695,N_22952,N_21702);
xor U26696 (N_26696,N_24021,N_21403);
nor U26697 (N_26697,N_23990,N_20639);
and U26698 (N_26698,N_24789,N_22209);
xnor U26699 (N_26699,N_23471,N_20369);
or U26700 (N_26700,N_22040,N_20450);
or U26701 (N_26701,N_24024,N_20937);
and U26702 (N_26702,N_21117,N_20069);
nand U26703 (N_26703,N_24330,N_23031);
and U26704 (N_26704,N_23694,N_22849);
xor U26705 (N_26705,N_24390,N_23551);
and U26706 (N_26706,N_24427,N_20325);
xor U26707 (N_26707,N_21765,N_22023);
and U26708 (N_26708,N_22004,N_20925);
nand U26709 (N_26709,N_22551,N_23809);
nand U26710 (N_26710,N_22807,N_22334);
and U26711 (N_26711,N_21354,N_22314);
xnor U26712 (N_26712,N_22064,N_20753);
or U26713 (N_26713,N_21349,N_22896);
nor U26714 (N_26714,N_24244,N_20821);
nand U26715 (N_26715,N_20892,N_21735);
and U26716 (N_26716,N_22683,N_24209);
nor U26717 (N_26717,N_21369,N_21808);
xnor U26718 (N_26718,N_21952,N_24422);
nor U26719 (N_26719,N_22116,N_21253);
nand U26720 (N_26720,N_21240,N_22623);
or U26721 (N_26721,N_21625,N_21341);
and U26722 (N_26722,N_22936,N_21500);
or U26723 (N_26723,N_24546,N_20637);
or U26724 (N_26724,N_21346,N_20315);
or U26725 (N_26725,N_20071,N_23997);
nor U26726 (N_26726,N_24841,N_21352);
xor U26727 (N_26727,N_22850,N_22532);
or U26728 (N_26728,N_21479,N_20942);
xnor U26729 (N_26729,N_21905,N_20331);
and U26730 (N_26730,N_23732,N_23509);
nand U26731 (N_26731,N_22586,N_23354);
nor U26732 (N_26732,N_20941,N_23574);
or U26733 (N_26733,N_24171,N_20225);
and U26734 (N_26734,N_21820,N_22474);
and U26735 (N_26735,N_21387,N_24705);
and U26736 (N_26736,N_23473,N_22253);
nor U26737 (N_26737,N_21872,N_23146);
and U26738 (N_26738,N_22699,N_22396);
and U26739 (N_26739,N_22447,N_20708);
nand U26740 (N_26740,N_21939,N_24172);
xnor U26741 (N_26741,N_22223,N_24933);
and U26742 (N_26742,N_23790,N_20791);
and U26743 (N_26743,N_23795,N_20747);
nor U26744 (N_26744,N_22680,N_20386);
and U26745 (N_26745,N_20052,N_20673);
nand U26746 (N_26746,N_23583,N_23595);
xor U26747 (N_26747,N_22795,N_24894);
and U26748 (N_26748,N_20907,N_24973);
or U26749 (N_26749,N_22804,N_23328);
or U26750 (N_26750,N_21367,N_24848);
or U26751 (N_26751,N_23221,N_21747);
and U26752 (N_26752,N_23584,N_20043);
or U26753 (N_26753,N_22987,N_22718);
or U26754 (N_26754,N_23298,N_24804);
nand U26755 (N_26755,N_22475,N_22547);
and U26756 (N_26756,N_23830,N_21430);
nor U26757 (N_26757,N_23789,N_24338);
nor U26758 (N_26758,N_21884,N_23327);
nand U26759 (N_26759,N_24045,N_21091);
and U26760 (N_26760,N_22029,N_23678);
xnor U26761 (N_26761,N_22580,N_21744);
and U26762 (N_26762,N_23889,N_23433);
nand U26763 (N_26763,N_23277,N_22517);
and U26764 (N_26764,N_22463,N_23088);
xnor U26765 (N_26765,N_20208,N_20630);
nor U26766 (N_26766,N_22028,N_21058);
or U26767 (N_26767,N_24775,N_21550);
or U26768 (N_26768,N_20288,N_24110);
xnor U26769 (N_26769,N_24657,N_23329);
and U26770 (N_26770,N_21568,N_23451);
nand U26771 (N_26771,N_22578,N_20721);
nand U26772 (N_26772,N_21474,N_20442);
nor U26773 (N_26773,N_24423,N_22760);
and U26774 (N_26774,N_22681,N_20077);
nor U26775 (N_26775,N_23601,N_23690);
and U26776 (N_26776,N_21431,N_23343);
or U26777 (N_26777,N_20205,N_20964);
xor U26778 (N_26778,N_24054,N_24097);
nand U26779 (N_26779,N_23487,N_20626);
nor U26780 (N_26780,N_24814,N_21150);
xnor U26781 (N_26781,N_20585,N_20924);
nand U26782 (N_26782,N_21017,N_22350);
and U26783 (N_26783,N_21167,N_23993);
and U26784 (N_26784,N_21440,N_22571);
nand U26785 (N_26785,N_22879,N_20332);
or U26786 (N_26786,N_24128,N_20049);
nor U26787 (N_26787,N_21265,N_20838);
or U26788 (N_26788,N_22479,N_24871);
nand U26789 (N_26789,N_20198,N_22546);
xnor U26790 (N_26790,N_21223,N_23933);
nand U26791 (N_26791,N_24940,N_24061);
or U26792 (N_26792,N_24903,N_22237);
and U26793 (N_26793,N_24987,N_20216);
or U26794 (N_26794,N_22351,N_21175);
and U26795 (N_26795,N_22844,N_20734);
or U26796 (N_26796,N_24300,N_22969);
xnor U26797 (N_26797,N_20280,N_23114);
nor U26798 (N_26798,N_20591,N_21255);
and U26799 (N_26799,N_24224,N_21155);
nor U26800 (N_26800,N_23091,N_21414);
and U26801 (N_26801,N_22744,N_20125);
nand U26802 (N_26802,N_20894,N_22031);
nor U26803 (N_26803,N_23504,N_21558);
and U26804 (N_26804,N_20273,N_22780);
nand U26805 (N_26805,N_23885,N_23805);
or U26806 (N_26806,N_21829,N_23142);
xor U26807 (N_26807,N_21157,N_22589);
and U26808 (N_26808,N_23978,N_23340);
and U26809 (N_26809,N_24159,N_23211);
xor U26810 (N_26810,N_20782,N_24790);
or U26811 (N_26811,N_23063,N_22757);
nor U26812 (N_26812,N_24384,N_20252);
or U26813 (N_26813,N_20508,N_22442);
xnor U26814 (N_26814,N_24854,N_22006);
nor U26815 (N_26815,N_24653,N_24266);
nand U26816 (N_26816,N_21570,N_22746);
or U26817 (N_26817,N_22194,N_22826);
and U26818 (N_26818,N_24832,N_21953);
nor U26819 (N_26819,N_21445,N_21736);
and U26820 (N_26820,N_20764,N_20574);
xor U26821 (N_26821,N_22102,N_21945);
xor U26822 (N_26822,N_20988,N_24150);
or U26823 (N_26823,N_21179,N_20062);
xnor U26824 (N_26824,N_23679,N_21343);
or U26825 (N_26825,N_23949,N_21777);
or U26826 (N_26826,N_20855,N_20912);
and U26827 (N_26827,N_21418,N_20029);
xor U26828 (N_26828,N_20557,N_23156);
nand U26829 (N_26829,N_21938,N_22387);
nand U26830 (N_26830,N_20287,N_22155);
or U26831 (N_26831,N_20416,N_22710);
or U26832 (N_26832,N_22233,N_20861);
and U26833 (N_26833,N_23039,N_21119);
xor U26834 (N_26834,N_23281,N_20692);
nor U26835 (N_26835,N_21565,N_22438);
or U26836 (N_26836,N_23676,N_21786);
or U26837 (N_26837,N_21838,N_24332);
xor U26838 (N_26838,N_24581,N_21108);
or U26839 (N_26839,N_22380,N_24022);
nand U26840 (N_26840,N_20577,N_20829);
nand U26841 (N_26841,N_23483,N_24559);
nor U26842 (N_26842,N_20709,N_23642);
and U26843 (N_26843,N_23532,N_21225);
or U26844 (N_26844,N_21845,N_20655);
xor U26845 (N_26845,N_24051,N_21185);
or U26846 (N_26846,N_24342,N_22734);
and U26847 (N_26847,N_22317,N_22663);
and U26848 (N_26848,N_23416,N_24339);
or U26849 (N_26849,N_21527,N_22595);
nor U26850 (N_26850,N_22451,N_24608);
or U26851 (N_26851,N_24840,N_21809);
and U26852 (N_26852,N_20240,N_24291);
nor U26853 (N_26853,N_22633,N_21887);
xnor U26854 (N_26854,N_20979,N_20597);
nand U26855 (N_26855,N_23208,N_20237);
and U26856 (N_26856,N_21912,N_22612);
and U26857 (N_26857,N_24317,N_22542);
nor U26858 (N_26858,N_23610,N_20775);
nor U26859 (N_26859,N_23544,N_21463);
or U26860 (N_26860,N_23592,N_24301);
and U26861 (N_26861,N_23769,N_22400);
nor U26862 (N_26862,N_24883,N_23824);
nor U26863 (N_26863,N_23561,N_20502);
and U26864 (N_26864,N_24091,N_22166);
nand U26865 (N_26865,N_20096,N_23774);
and U26866 (N_26866,N_24669,N_23352);
or U26867 (N_26867,N_23104,N_21252);
xnor U26868 (N_26868,N_24749,N_23409);
or U26869 (N_26869,N_20480,N_24782);
and U26870 (N_26870,N_23996,N_24376);
or U26871 (N_26871,N_23048,N_22310);
nand U26872 (N_26872,N_23346,N_24815);
or U26873 (N_26873,N_24109,N_24617);
and U26874 (N_26874,N_23827,N_23639);
and U26875 (N_26875,N_22847,N_21452);
xor U26876 (N_26876,N_23930,N_21924);
nor U26877 (N_26877,N_22217,N_21914);
and U26878 (N_26878,N_22326,N_21971);
or U26879 (N_26879,N_20943,N_23134);
xor U26880 (N_26880,N_22234,N_22908);
and U26881 (N_26881,N_23648,N_21147);
xor U26882 (N_26882,N_21498,N_24838);
and U26883 (N_26883,N_22190,N_21941);
xnor U26884 (N_26884,N_20720,N_23992);
and U26885 (N_26885,N_20878,N_21624);
nor U26886 (N_26886,N_24999,N_24622);
nor U26887 (N_26887,N_20883,N_24813);
nand U26888 (N_26888,N_21409,N_24819);
or U26889 (N_26889,N_21813,N_24205);
or U26890 (N_26890,N_23194,N_22564);
xor U26891 (N_26891,N_24174,N_23075);
nand U26892 (N_26892,N_21489,N_24164);
nand U26893 (N_26893,N_23955,N_20723);
nand U26894 (N_26894,N_20003,N_22816);
nand U26895 (N_26895,N_20404,N_24471);
xor U26896 (N_26896,N_24557,N_20735);
xnor U26897 (N_26897,N_23619,N_21638);
xor U26898 (N_26898,N_24863,N_22537);
nor U26899 (N_26899,N_23360,N_21897);
xor U26900 (N_26900,N_20953,N_20906);
xnor U26901 (N_26901,N_22884,N_24757);
and U26902 (N_26902,N_21566,N_21034);
or U26903 (N_26903,N_24747,N_24513);
xnor U26904 (N_26904,N_22273,N_20976);
nor U26905 (N_26905,N_20773,N_22894);
nor U26906 (N_26906,N_24625,N_24575);
nor U26907 (N_26907,N_23107,N_24845);
and U26908 (N_26908,N_21701,N_23457);
and U26909 (N_26909,N_20218,N_24862);
and U26910 (N_26910,N_23018,N_23161);
xor U26911 (N_26911,N_20669,N_22771);
and U26912 (N_26912,N_24029,N_24204);
or U26913 (N_26913,N_24687,N_22409);
nor U26914 (N_26914,N_23446,N_24746);
or U26915 (N_26915,N_22196,N_20033);
or U26916 (N_26916,N_24951,N_21258);
or U26917 (N_26917,N_21659,N_24033);
nor U26918 (N_26918,N_23231,N_24833);
nand U26919 (N_26919,N_24031,N_22677);
nand U26920 (N_26920,N_20761,N_20774);
nor U26921 (N_26921,N_21503,N_24887);
nand U26922 (N_26922,N_21482,N_22765);
nand U26923 (N_26923,N_22113,N_22773);
xnor U26924 (N_26924,N_21641,N_20178);
or U26925 (N_26925,N_20885,N_24891);
xnor U26926 (N_26926,N_24713,N_21499);
nand U26927 (N_26927,N_20902,N_24673);
nand U26928 (N_26928,N_23450,N_24510);
nand U26929 (N_26929,N_22958,N_23006);
or U26930 (N_26930,N_20848,N_23818);
and U26931 (N_26931,N_20904,N_20790);
and U26932 (N_26932,N_24337,N_22427);
or U26933 (N_26933,N_23169,N_22332);
xnor U26934 (N_26934,N_23576,N_23292);
or U26935 (N_26935,N_24702,N_22576);
nand U26936 (N_26936,N_24321,N_23786);
and U26937 (N_26937,N_24437,N_24679);
and U26938 (N_26938,N_21200,N_22434);
or U26939 (N_26939,N_23464,N_23600);
or U26940 (N_26940,N_20389,N_22117);
nor U26941 (N_26941,N_22747,N_24946);
xor U26942 (N_26942,N_21151,N_20728);
nand U26943 (N_26943,N_21509,N_22048);
nand U26944 (N_26944,N_24299,N_22825);
and U26945 (N_26945,N_23111,N_21256);
nand U26946 (N_26946,N_23237,N_21773);
or U26947 (N_26947,N_23770,N_20333);
nor U26948 (N_26948,N_21770,N_23167);
or U26949 (N_26949,N_22798,N_20661);
or U26950 (N_26950,N_22717,N_22188);
nand U26951 (N_26951,N_22318,N_20142);
or U26952 (N_26952,N_20719,N_23033);
and U26953 (N_26953,N_23762,N_24915);
or U26954 (N_26954,N_24630,N_20819);
nand U26955 (N_26955,N_22354,N_22888);
xnor U26956 (N_26956,N_21885,N_20055);
xnor U26957 (N_26957,N_21230,N_20440);
nand U26958 (N_26958,N_20845,N_20602);
xor U26959 (N_26959,N_20615,N_23252);
and U26960 (N_26960,N_20181,N_22855);
and U26961 (N_26961,N_22054,N_20167);
xnor U26962 (N_26962,N_23219,N_21900);
and U26963 (N_26963,N_22997,N_20997);
nand U26964 (N_26964,N_20189,N_23511);
nor U26965 (N_26965,N_21131,N_23994);
nor U26966 (N_26966,N_23792,N_24882);
xor U26967 (N_26967,N_24689,N_20936);
and U26968 (N_26968,N_23188,N_23230);
nand U26969 (N_26969,N_22053,N_24909);
nand U26970 (N_26970,N_20258,N_24016);
xnor U26971 (N_26971,N_20951,N_23045);
xor U26972 (N_26972,N_20500,N_21867);
nand U26973 (N_26973,N_20877,N_21271);
xnor U26974 (N_26974,N_24470,N_20190);
nor U26975 (N_26975,N_21519,N_24293);
xnor U26976 (N_26976,N_20388,N_22859);
or U26977 (N_26977,N_23407,N_24964);
or U26978 (N_26978,N_24870,N_22084);
nand U26979 (N_26979,N_24467,N_23159);
and U26980 (N_26980,N_22513,N_24899);
nor U26981 (N_26981,N_21583,N_20162);
nand U26982 (N_26982,N_21484,N_21365);
nor U26983 (N_26983,N_20170,N_21501);
nand U26984 (N_26984,N_20177,N_20254);
xor U26985 (N_26985,N_20896,N_22311);
xnor U26986 (N_26986,N_20298,N_21005);
nand U26987 (N_26987,N_22759,N_21425);
or U26988 (N_26988,N_23731,N_24797);
xnor U26989 (N_26989,N_21006,N_24849);
xor U26990 (N_26990,N_23959,N_24052);
nor U26991 (N_26991,N_24997,N_24860);
nor U26992 (N_26992,N_21143,N_23067);
xnor U26993 (N_26993,N_20290,N_24270);
or U26994 (N_26994,N_20230,N_22919);
nand U26995 (N_26995,N_21298,N_22686);
or U26996 (N_26996,N_22388,N_22900);
xnor U26997 (N_26997,N_24018,N_23297);
nor U26998 (N_26998,N_22165,N_22378);
nand U26999 (N_26999,N_20490,N_20884);
xnor U27000 (N_27000,N_21038,N_23573);
xnor U27001 (N_27001,N_20242,N_22243);
and U27002 (N_27002,N_24241,N_24343);
or U27003 (N_27003,N_21378,N_24030);
or U27004 (N_27004,N_21206,N_20882);
nand U27005 (N_27005,N_23158,N_20496);
nand U27006 (N_27006,N_20507,N_21732);
and U27007 (N_27007,N_21699,N_22002);
and U27008 (N_27008,N_24105,N_20050);
or U27009 (N_27009,N_20554,N_24812);
or U27010 (N_27010,N_23522,N_22679);
or U27011 (N_27011,N_22411,N_21749);
and U27012 (N_27012,N_22128,N_21488);
and U27013 (N_27013,N_24711,N_21389);
nor U27014 (N_27014,N_22280,N_21132);
or U27015 (N_27015,N_23287,N_20256);
or U27016 (N_27016,N_23456,N_22646);
xor U27017 (N_27017,N_21601,N_20702);
xor U27018 (N_27018,N_22868,N_22256);
nor U27019 (N_27019,N_23680,N_23106);
xnor U27020 (N_27020,N_23377,N_20168);
xor U27021 (N_27021,N_22205,N_23361);
or U27022 (N_27022,N_22503,N_23871);
or U27023 (N_27023,N_20612,N_24309);
and U27024 (N_27024,N_21305,N_21947);
nand U27025 (N_27025,N_24583,N_21999);
nor U27026 (N_27026,N_21870,N_21992);
and U27027 (N_27027,N_23392,N_24744);
nand U27028 (N_27028,N_20550,N_23072);
and U27029 (N_27029,N_20089,N_21513);
xor U27030 (N_27030,N_24362,N_21094);
nor U27031 (N_27031,N_20509,N_20422);
nor U27032 (N_27032,N_22617,N_22853);
and U27033 (N_27033,N_22414,N_23587);
nand U27034 (N_27034,N_20026,N_21492);
nor U27035 (N_27035,N_20926,N_23750);
and U27036 (N_27036,N_22735,N_21242);
or U27037 (N_27037,N_22446,N_20778);
nor U27038 (N_27038,N_20600,N_20824);
or U27039 (N_27039,N_23027,N_23119);
and U27040 (N_27040,N_24656,N_21010);
nor U27041 (N_27041,N_22601,N_20705);
and U27042 (N_27042,N_24795,N_24714);
nor U27043 (N_27043,N_22255,N_21471);
and U27044 (N_27044,N_20223,N_23008);
xnor U27045 (N_27045,N_21308,N_20468);
xor U27046 (N_27046,N_20553,N_20025);
nor U27047 (N_27047,N_20027,N_22841);
nor U27048 (N_27048,N_24247,N_22238);
and U27049 (N_27049,N_20505,N_21168);
nor U27050 (N_27050,N_22829,N_22456);
nand U27051 (N_27051,N_20595,N_20066);
and U27052 (N_27052,N_21231,N_20039);
xor U27053 (N_27053,N_23432,N_20645);
or U27054 (N_27054,N_23938,N_23728);
and U27055 (N_27055,N_22239,N_24913);
nor U27056 (N_27056,N_24994,N_23468);
nor U27057 (N_27057,N_22867,N_21591);
nand U27058 (N_27058,N_21955,N_24846);
nor U27059 (N_27059,N_20980,N_20161);
and U27060 (N_27060,N_20336,N_20621);
nand U27061 (N_27061,N_22619,N_24188);
or U27062 (N_27062,N_24025,N_22480);
or U27063 (N_27063,N_21689,N_21202);
and U27064 (N_27064,N_20583,N_22941);
xnor U27065 (N_27065,N_24340,N_21158);
nor U27066 (N_27066,N_21661,N_24004);
and U27067 (N_27067,N_24751,N_23806);
and U27068 (N_27068,N_23811,N_22764);
nand U27069 (N_27069,N_21505,N_20126);
and U27070 (N_27070,N_20970,N_20770);
and U27071 (N_27071,N_22787,N_23384);
nand U27072 (N_27072,N_23199,N_20640);
nor U27073 (N_27073,N_22082,N_20094);
nand U27074 (N_27074,N_23907,N_24547);
and U27075 (N_27075,N_23773,N_24334);
nor U27076 (N_27076,N_24588,N_23013);
and U27077 (N_27077,N_22697,N_21635);
and U27078 (N_27078,N_24243,N_20156);
nor U27079 (N_27079,N_20402,N_22278);
and U27080 (N_27080,N_22335,N_22304);
or U27081 (N_27081,N_24901,N_20609);
or U27082 (N_27082,N_22153,N_21510);
or U27083 (N_27083,N_21102,N_23348);
nor U27084 (N_27084,N_23463,N_22749);
xnor U27085 (N_27085,N_23693,N_21580);
nand U27086 (N_27086,N_21846,N_24080);
nand U27087 (N_27087,N_23552,N_20294);
and U27088 (N_27088,N_20406,N_22254);
nand U27089 (N_27089,N_24639,N_21284);
nor U27090 (N_27090,N_23893,N_20271);
nor U27091 (N_27091,N_21579,N_20073);
and U27092 (N_27092,N_23112,N_21088);
and U27093 (N_27093,N_20024,N_21574);
xnor U27094 (N_27094,N_20613,N_21651);
or U27095 (N_27095,N_24677,N_22590);
xnor U27096 (N_27096,N_23131,N_20098);
xor U27097 (N_27097,N_24261,N_22923);
or U27098 (N_27098,N_21303,N_23129);
and U27099 (N_27099,N_21807,N_22622);
xnor U27100 (N_27100,N_21146,N_21593);
and U27101 (N_27101,N_24194,N_22815);
xnor U27102 (N_27102,N_23405,N_24529);
nor U27103 (N_27103,N_24618,N_20394);
nor U27104 (N_27104,N_21462,N_20399);
xor U27105 (N_27105,N_21275,N_24607);
and U27106 (N_27106,N_21364,N_24551);
nor U27107 (N_27107,N_21458,N_24251);
nand U27108 (N_27108,N_24945,N_24441);
nor U27109 (N_27109,N_23224,N_21649);
and U27110 (N_27110,N_22665,N_23429);
nor U27111 (N_27111,N_22098,N_20085);
xnor U27112 (N_27112,N_20342,N_21107);
or U27113 (N_27113,N_24556,N_23607);
nor U27114 (N_27114,N_23372,N_22938);
nand U27115 (N_27115,N_23109,N_23609);
nand U27116 (N_27116,N_20663,N_24498);
or U27117 (N_27117,N_20065,N_21060);
nand U27118 (N_27118,N_22719,N_20526);
nand U27119 (N_27119,N_24218,N_23497);
nand U27120 (N_27120,N_21033,N_23982);
and U27121 (N_27121,N_22296,N_22922);
or U27122 (N_27122,N_20285,N_23010);
or U27123 (N_27123,N_23216,N_20435);
and U27124 (N_27124,N_20968,N_22701);
and U27125 (N_27125,N_22079,N_24754);
or U27126 (N_27126,N_24916,N_23874);
nand U27127 (N_27127,N_20955,N_22903);
nand U27128 (N_27128,N_22752,N_24876);
nand U27129 (N_27129,N_24487,N_24108);
or U27130 (N_27130,N_20529,N_21957);
nand U27131 (N_27131,N_21988,N_23147);
nor U27132 (N_27132,N_22581,N_24446);
nor U27133 (N_27133,N_23467,N_20827);
nand U27134 (N_27134,N_23567,N_23886);
nand U27135 (N_27135,N_23305,N_24438);
nor U27136 (N_27136,N_20675,N_23716);
nor U27137 (N_27137,N_22221,N_24822);
nand U27138 (N_27138,N_24659,N_24143);
xor U27139 (N_27139,N_22180,N_23891);
nor U27140 (N_27140,N_21205,N_24431);
xnor U27141 (N_27141,N_24752,N_23273);
or U27142 (N_27142,N_22057,N_23421);
nand U27143 (N_27143,N_20169,N_22983);
or U27144 (N_27144,N_23867,N_21241);
xnor U27145 (N_27145,N_22707,N_24993);
or U27146 (N_27146,N_21335,N_21042);
or U27147 (N_27147,N_20945,N_23644);
nor U27148 (N_27148,N_20533,N_23339);
and U27149 (N_27149,N_22035,N_21274);
xnor U27150 (N_27150,N_24066,N_24356);
and U27151 (N_27151,N_20575,N_20233);
and U27152 (N_27152,N_20213,N_24485);
nor U27153 (N_27153,N_21803,N_24998);
xnor U27154 (N_27154,N_21920,N_20278);
nand U27155 (N_27155,N_21003,N_24995);
xor U27156 (N_27156,N_21961,N_24755);
or U27157 (N_27157,N_21581,N_20370);
xor U27158 (N_27158,N_24971,N_23475);
and U27159 (N_27159,N_24571,N_24665);
and U27160 (N_27160,N_22140,N_22772);
nor U27161 (N_27161,N_22618,N_22871);
xnor U27162 (N_27162,N_21631,N_24249);
nor U27163 (N_27163,N_23275,N_22220);
or U27164 (N_27164,N_22170,N_22367);
and U27165 (N_27165,N_21594,N_24413);
nand U27166 (N_27166,N_23258,N_23288);
nand U27167 (N_27167,N_20636,N_22007);
nand U27168 (N_27168,N_24219,N_20586);
or U27169 (N_27169,N_21081,N_23539);
xnor U27170 (N_27170,N_23380,N_21530);
xnor U27171 (N_27171,N_20054,N_22935);
and U27172 (N_27172,N_23688,N_22892);
or U27173 (N_27173,N_23125,N_24758);
or U27174 (N_27174,N_23960,N_23378);
xnor U27175 (N_27175,N_20320,N_22652);
nor U27176 (N_27176,N_22587,N_21178);
and U27177 (N_27177,N_22229,N_23513);
or U27178 (N_27178,N_21931,N_23127);
and U27179 (N_27179,N_23550,N_23659);
nand U27180 (N_27180,N_24392,N_22893);
xnor U27181 (N_27181,N_22739,N_20354);
or U27182 (N_27182,N_24544,N_22405);
or U27183 (N_27183,N_20564,N_20013);
or U27184 (N_27184,N_20040,N_24662);
or U27185 (N_27185,N_20193,N_21627);
nor U27186 (N_27186,N_22998,N_22020);
xor U27187 (N_27187,N_22184,N_21783);
or U27188 (N_27188,N_21560,N_21709);
and U27189 (N_27189,N_24049,N_24939);
or U27190 (N_27190,N_22836,N_23981);
nor U27191 (N_27191,N_23333,N_20916);
nand U27192 (N_27192,N_22641,N_24911);
nor U27193 (N_27193,N_24652,N_21967);
nand U27194 (N_27194,N_22934,N_22755);
nand U27195 (N_27195,N_21331,N_20010);
xor U27196 (N_27196,N_22087,N_23485);
or U27197 (N_27197,N_22286,N_22630);
or U27198 (N_27198,N_24276,N_22971);
xor U27199 (N_27199,N_23835,N_23020);
and U27200 (N_27200,N_23256,N_23206);
nand U27201 (N_27201,N_22483,N_21758);
nor U27202 (N_27202,N_21348,N_21089);
or U27203 (N_27203,N_24094,N_22732);
xor U27204 (N_27204,N_21466,N_23187);
or U27205 (N_27205,N_21815,N_22653);
or U27206 (N_27206,N_22298,N_22097);
and U27207 (N_27207,N_21622,N_21779);
nand U27208 (N_27208,N_20814,N_20808);
nand U27209 (N_27209,N_21310,N_24283);
nand U27210 (N_27210,N_24931,N_21577);
nand U27211 (N_27211,N_20172,N_20593);
nand U27212 (N_27212,N_20872,N_24806);
xnor U27213 (N_27213,N_20961,N_24560);
or U27214 (N_27214,N_24530,N_24085);
nor U27215 (N_27215,N_21304,N_24428);
nand U27216 (N_27216,N_24990,N_22761);
or U27217 (N_27217,N_20658,N_20079);
and U27218 (N_27218,N_24923,N_24072);
or U27219 (N_27219,N_20145,N_22666);
and U27220 (N_27220,N_24565,N_20051);
nor U27221 (N_27221,N_20462,N_21001);
and U27222 (N_27222,N_22457,N_22966);
or U27223 (N_27223,N_20539,N_21810);
nor U27224 (N_27224,N_23083,N_23047);
and U27225 (N_27225,N_22950,N_20686);
or U27226 (N_27226,N_24296,N_24181);
xor U27227 (N_27227,N_22308,N_20304);
and U27228 (N_27228,N_22712,N_24264);
and U27229 (N_27229,N_24436,N_22026);
nor U27230 (N_27230,N_23613,N_23763);
or U27231 (N_27231,N_21210,N_24550);
nand U27232 (N_27232,N_22636,N_22534);
or U27233 (N_27233,N_20641,N_20816);
xor U27234 (N_27234,N_23523,N_20006);
and U27235 (N_27235,N_24842,N_23577);
or U27236 (N_27236,N_20260,N_24180);
and U27237 (N_27237,N_23102,N_22134);
and U27238 (N_27238,N_22014,N_24696);
nand U27239 (N_27239,N_20269,N_21260);
xor U27240 (N_27240,N_23175,N_21037);
nor U27241 (N_27241,N_22716,N_23703);
or U27242 (N_27242,N_22726,N_24621);
or U27243 (N_27243,N_20253,N_20195);
or U27244 (N_27244,N_22491,N_21930);
xnor U27245 (N_27245,N_24611,N_23484);
or U27246 (N_27246,N_24318,N_23024);
and U27247 (N_27247,N_20080,N_20802);
and U27248 (N_27248,N_21199,N_21855);
xor U27249 (N_27249,N_21538,N_24375);
nor U27250 (N_27250,N_24851,N_21161);
and U27251 (N_27251,N_21869,N_21133);
nand U27252 (N_27252,N_24792,N_20152);
or U27253 (N_27253,N_20664,N_24765);
nor U27254 (N_27254,N_21667,N_23624);
and U27255 (N_27255,N_24569,N_24449);
and U27256 (N_27256,N_22379,N_21279);
or U27257 (N_27257,N_20685,N_22324);
nand U27258 (N_27258,N_21856,N_21572);
or U27259 (N_27259,N_20587,N_20568);
or U27260 (N_27260,N_21525,N_24552);
nand U27261 (N_27261,N_21684,N_22626);
nor U27262 (N_27262,N_20349,N_23564);
xnor U27263 (N_27263,N_22954,N_21586);
or U27264 (N_27264,N_20097,N_24788);
or U27265 (N_27265,N_20841,N_20346);
nand U27266 (N_27266,N_21844,N_20694);
nor U27267 (N_27267,N_23921,N_20474);
nor U27268 (N_27268,N_21351,N_20820);
or U27269 (N_27269,N_22371,N_22510);
and U27270 (N_27270,N_21340,N_22740);
or U27271 (N_27271,N_21891,N_20850);
or U27272 (N_27272,N_21061,N_20466);
nand U27273 (N_27273,N_21923,N_24294);
xnor U27274 (N_27274,N_20313,N_23141);
xnor U27275 (N_27275,N_23531,N_21004);
nand U27276 (N_27276,N_21575,N_22183);
nor U27277 (N_27277,N_20295,N_24354);
or U27278 (N_27278,N_24187,N_23400);
or U27279 (N_27279,N_23395,N_20793);
nand U27280 (N_27280,N_20952,N_21582);
and U27281 (N_27281,N_23247,N_21073);
nor U27282 (N_27282,N_22263,N_24432);
xor U27283 (N_27283,N_22342,N_22422);
nor U27284 (N_27284,N_22522,N_21672);
nand U27285 (N_27285,N_22661,N_24853);
xnor U27286 (N_27286,N_20983,N_23553);
nand U27287 (N_27287,N_24481,N_24013);
nand U27288 (N_27288,N_23700,N_23080);
and U27289 (N_27289,N_24948,N_20413);
xor U27290 (N_27290,N_21412,N_22399);
nor U27291 (N_27291,N_22854,N_23220);
and U27292 (N_27292,N_20743,N_20470);
or U27293 (N_27293,N_22912,N_21344);
and U27294 (N_27294,N_22265,N_24316);
or U27295 (N_27295,N_24056,N_21898);
or U27296 (N_27296,N_22468,N_22531);
xor U27297 (N_27297,N_21771,N_24686);
nand U27298 (N_27298,N_21692,N_20008);
xnor U27299 (N_27299,N_23803,N_22157);
or U27300 (N_27300,N_24409,N_23181);
xor U27301 (N_27301,N_21639,N_22599);
xor U27302 (N_27302,N_23602,N_22775);
nor U27303 (N_27303,N_22857,N_24567);
nand U27304 (N_27304,N_22911,N_23869);
nand U27305 (N_27305,N_20144,N_23076);
xor U27306 (N_27306,N_23859,N_23435);
nand U27307 (N_27307,N_23419,N_23503);
xor U27308 (N_27308,N_21906,N_21880);
nand U27309 (N_27309,N_23123,N_22303);
nand U27310 (N_27310,N_21737,N_20337);
nand U27311 (N_27311,N_24717,N_23155);
xnor U27312 (N_27312,N_22642,N_20691);
xnor U27313 (N_27313,N_20112,N_22225);
nand U27314 (N_27314,N_22034,N_23962);
nor U27315 (N_27315,N_24954,N_21273);
nand U27316 (N_27316,N_23783,N_23160);
nor U27317 (N_27317,N_20106,N_23151);
or U27318 (N_27318,N_23437,N_20932);
nand U27319 (N_27319,N_20110,N_20598);
and U27320 (N_27320,N_20908,N_24874);
xnor U27321 (N_27321,N_24101,N_22611);
and U27322 (N_27322,N_20513,N_24353);
nor U27323 (N_27323,N_24623,N_20625);
xnor U27324 (N_27324,N_22600,N_23285);
and U27325 (N_27325,N_24825,N_21070);
nor U27326 (N_27326,N_24900,N_22284);
nand U27327 (N_27327,N_20447,N_20498);
or U27328 (N_27328,N_22988,N_21312);
xnor U27329 (N_27329,N_20341,N_20629);
xnor U27330 (N_27330,N_22261,N_22741);
or U27331 (N_27331,N_22528,N_21871);
xnor U27332 (N_27332,N_24399,N_24646);
nand U27333 (N_27333,N_24515,N_23734);
and U27334 (N_27334,N_21417,N_23234);
xnor U27335 (N_27335,N_20752,N_21986);
or U27336 (N_27336,N_22312,N_24442);
nor U27337 (N_27337,N_24472,N_22837);
xnor U27338 (N_27338,N_22081,N_21475);
nand U27339 (N_27339,N_20579,N_23438);
xnor U27340 (N_27340,N_21100,N_21251);
nand U27341 (N_27341,N_22964,N_21801);
xnor U27342 (N_27342,N_23815,N_20324);
and U27343 (N_27343,N_21832,N_21153);
and U27344 (N_27344,N_23408,N_22382);
or U27345 (N_27345,N_22494,N_22349);
nor U27346 (N_27346,N_22250,N_21785);
nor U27347 (N_27347,N_23495,N_24875);
xnor U27348 (N_27348,N_24511,N_22333);
nand U27349 (N_27349,N_20810,N_21402);
and U27350 (N_27350,N_20318,N_20438);
nor U27351 (N_27351,N_23829,N_22526);
nor U27352 (N_27352,N_20259,N_24488);
or U27353 (N_27353,N_22453,N_21390);
nor U27354 (N_27354,N_20481,N_22660);
xor U27355 (N_27355,N_21224,N_22812);
nor U27356 (N_27356,N_20867,N_22106);
xnor U27357 (N_27357,N_20212,N_24237);
nor U27358 (N_27358,N_23881,N_24616);
or U27359 (N_27359,N_22769,N_22068);
nor U27360 (N_27360,N_23661,N_20141);
nand U27361 (N_27361,N_20540,N_23534);
nand U27362 (N_27362,N_21731,N_24263);
nor U27363 (N_27363,N_23840,N_23110);
nand U27364 (N_27364,N_23863,N_20510);
nor U27365 (N_27365,N_20940,N_20021);
nand U27366 (N_27366,N_21670,N_22870);
nor U27367 (N_27367,N_24077,N_20631);
and U27368 (N_27368,N_22226,N_20776);
nor U27369 (N_27369,N_21450,N_24785);
nand U27370 (N_27370,N_22227,N_23974);
nor U27371 (N_27371,N_23589,N_23649);
xnor U27372 (N_27372,N_20012,N_24060);
or U27373 (N_27373,N_20492,N_20091);
and U27374 (N_27374,N_23969,N_20797);
nand U27375 (N_27375,N_21657,N_22915);
nor U27376 (N_27376,N_22143,N_21539);
xnor U27377 (N_27377,N_24506,N_20680);
nor U27378 (N_27378,N_21890,N_20654);
or U27379 (N_27379,N_21285,N_23430);
nand U27380 (N_27380,N_21552,N_20562);
nor U27381 (N_27381,N_23691,N_22501);
nand U27382 (N_27382,N_20424,N_21965);
nand U27383 (N_27383,N_22891,N_21483);
xor U27384 (N_27384,N_20811,N_24230);
or U27385 (N_27385,N_23689,N_23402);
or U27386 (N_27386,N_22445,N_23422);
nand U27387 (N_27387,N_20347,N_22591);
nor U27388 (N_27388,N_24026,N_20398);
or U27389 (N_27389,N_23259,N_24736);
nor U27390 (N_27390,N_23302,N_23019);
xnor U27391 (N_27391,N_22607,N_24252);
nor U27392 (N_27392,N_22917,N_20366);
nand U27393 (N_27393,N_20486,N_20380);
and U27394 (N_27394,N_22356,N_23322);
or U27395 (N_27395,N_24419,N_21083);
nand U27396 (N_27396,N_22247,N_23894);
nor U27397 (N_27397,N_20531,N_22662);
nand U27398 (N_27398,N_20987,N_24773);
nor U27399 (N_27399,N_21361,N_21164);
nand U27400 (N_27400,N_20364,N_24570);
nand U27401 (N_27401,N_24367,N_22341);
nand U27402 (N_27402,N_22991,N_20818);
nor U27403 (N_27403,N_24086,N_21893);
xnor U27404 (N_27404,N_21571,N_20100);
or U27405 (N_27405,N_21926,N_20781);
nor U27406 (N_27406,N_23269,N_20601);
nor U27407 (N_27407,N_23133,N_20188);
xor U27408 (N_27408,N_21180,N_23428);
xnor U27409 (N_27409,N_21995,N_20384);
and U27410 (N_27410,N_20828,N_22293);
nand U27411 (N_27411,N_22440,N_20405);
nand U27412 (N_27412,N_21919,N_22968);
xnor U27413 (N_27413,N_20262,N_24305);
nand U27414 (N_27414,N_21619,N_24179);
xnor U27415 (N_27415,N_21460,N_24285);
and U27416 (N_27416,N_24039,N_20093);
nor U27417 (N_27417,N_20099,N_23687);
or U27418 (N_27418,N_24548,N_22419);
or U27419 (N_27419,N_21548,N_20551);
nand U27420 (N_27420,N_20072,N_21039);
or U27421 (N_27421,N_22122,N_21194);
nor U27422 (N_27422,N_23841,N_23950);
or U27423 (N_27423,N_21319,N_21643);
or U27424 (N_27424,N_20792,N_21421);
or U27425 (N_27425,N_24517,N_23126);
nor U27426 (N_27426,N_22668,N_24963);
nand U27427 (N_27427,N_21420,N_20736);
nand U27428 (N_27428,N_22762,N_24059);
nand U27429 (N_27429,N_23508,N_22389);
xnor U27430 (N_27430,N_22181,N_24943);
nand U27431 (N_27431,N_23267,N_21717);
nand U27432 (N_27432,N_24969,N_23124);
xnor U27433 (N_27433,N_22109,N_21410);
and U27434 (N_27434,N_20701,N_21557);
xor U27435 (N_27435,N_22819,N_21121);
or U27436 (N_27436,N_24211,N_24007);
xor U27437 (N_27437,N_22232,N_22464);
and U27438 (N_27438,N_20875,N_22606);
xor U27439 (N_27439,N_23714,N_20412);
or U27440 (N_27440,N_20164,N_23338);
nand U27441 (N_27441,N_23729,N_20578);
nor U27442 (N_27442,N_21165,N_22061);
nor U27443 (N_27443,N_22139,N_21477);
nor U27444 (N_27444,N_20982,N_22358);
xor U27445 (N_27445,N_23733,N_24005);
or U27446 (N_27446,N_20745,N_20672);
xor U27447 (N_27447,N_23092,N_24793);
nor U27448 (N_27448,N_24835,N_23154);
nand U27449 (N_27449,N_22017,N_21739);
nand U27450 (N_27450,N_22539,N_22088);
and U27451 (N_27451,N_20891,N_21490);
nor U27452 (N_27452,N_24278,N_20070);
or U27453 (N_27453,N_24082,N_21296);
nor U27454 (N_27454,N_23842,N_22240);
or U27455 (N_27455,N_21334,N_20880);
nand U27456 (N_27456,N_24461,N_20607);
nand U27457 (N_27457,N_22206,N_22996);
nand U27458 (N_27458,N_22027,N_23186);
nand U27459 (N_27459,N_21473,N_24003);
and U27460 (N_27460,N_20668,N_23746);
and U27461 (N_27461,N_21921,N_20009);
or U27462 (N_27462,N_20392,N_23670);
or U27463 (N_27463,N_23351,N_21873);
nor U27464 (N_27464,N_24455,N_23178);
nor U27465 (N_27465,N_22325,N_23961);
nand U27466 (N_27466,N_22114,N_23903);
nor U27467 (N_27467,N_21985,N_20018);
xnor U27468 (N_27468,N_22800,N_20437);
and U27469 (N_27469,N_22803,N_20419);
xnor U27470 (N_27470,N_24817,N_20825);
nor U27471 (N_27471,N_24678,N_23793);
xnor U27472 (N_27472,N_20619,N_21190);
nand U27473 (N_27473,N_23184,N_23213);
xor U27474 (N_27474,N_24369,N_23782);
and U27475 (N_27475,N_22013,N_20214);
nor U27476 (N_27476,N_24424,N_22402);
nand U27477 (N_27477,N_23263,N_21611);
nand U27478 (N_27478,N_24214,N_21204);
xnor U27479 (N_27479,N_23185,N_23268);
nor U27480 (N_27480,N_21847,N_21588);
nor U27481 (N_27481,N_20267,N_20756);
nor U27482 (N_27482,N_23306,N_23641);
xnor U27483 (N_27483,N_23612,N_22972);
and U27484 (N_27484,N_20682,N_22051);
xor U27485 (N_27485,N_24561,N_21545);
or U27486 (N_27486,N_23014,N_22120);
nor U27487 (N_27487,N_20382,N_24768);
nor U27488 (N_27488,N_22843,N_22486);
nand U27489 (N_27489,N_22940,N_23743);
nor U27490 (N_27490,N_23066,N_23389);
or U27491 (N_27491,N_24988,N_24914);
and U27492 (N_27492,N_21613,N_21345);
nor U27493 (N_27493,N_23951,N_24699);
nor U27494 (N_27494,N_22365,N_20376);
nand U27495 (N_27495,N_24839,N_24671);
xnor U27496 (N_27496,N_21799,N_24535);
nand U27497 (N_27497,N_20922,N_23890);
xnor U27498 (N_27498,N_23235,N_24482);
nor U27499 (N_27499,N_20972,N_24145);
and U27500 (N_27500,N_24597,N_21266);
nor U27501 (N_27501,N_20437,N_22413);
nand U27502 (N_27502,N_24012,N_23958);
or U27503 (N_27503,N_20242,N_22200);
xnor U27504 (N_27504,N_22228,N_22236);
xor U27505 (N_27505,N_21542,N_22529);
xor U27506 (N_27506,N_20601,N_21074);
nor U27507 (N_27507,N_20814,N_20555);
nor U27508 (N_27508,N_24022,N_23351);
and U27509 (N_27509,N_21288,N_22136);
nor U27510 (N_27510,N_20129,N_24227);
xor U27511 (N_27511,N_24847,N_22753);
nand U27512 (N_27512,N_22884,N_22057);
nand U27513 (N_27513,N_24237,N_21960);
and U27514 (N_27514,N_23368,N_22944);
nand U27515 (N_27515,N_21999,N_21028);
nand U27516 (N_27516,N_22443,N_20214);
and U27517 (N_27517,N_21623,N_20679);
nand U27518 (N_27518,N_20763,N_24704);
nand U27519 (N_27519,N_24641,N_20197);
xnor U27520 (N_27520,N_23393,N_21866);
xor U27521 (N_27521,N_21944,N_20055);
or U27522 (N_27522,N_20427,N_23327);
and U27523 (N_27523,N_23577,N_23008);
or U27524 (N_27524,N_22984,N_21431);
and U27525 (N_27525,N_22239,N_23736);
xnor U27526 (N_27526,N_23236,N_24405);
nand U27527 (N_27527,N_24650,N_24112);
nand U27528 (N_27528,N_20763,N_21089);
xor U27529 (N_27529,N_23741,N_21591);
nor U27530 (N_27530,N_24950,N_20678);
nand U27531 (N_27531,N_20074,N_20448);
or U27532 (N_27532,N_20219,N_22747);
or U27533 (N_27533,N_21520,N_20313);
and U27534 (N_27534,N_20683,N_22055);
xnor U27535 (N_27535,N_22839,N_24208);
or U27536 (N_27536,N_23976,N_20165);
xor U27537 (N_27537,N_21413,N_20336);
nand U27538 (N_27538,N_21958,N_23458);
xor U27539 (N_27539,N_22536,N_22906);
nor U27540 (N_27540,N_24320,N_21717);
xor U27541 (N_27541,N_24790,N_24173);
nand U27542 (N_27542,N_24551,N_24830);
nand U27543 (N_27543,N_22842,N_21765);
or U27544 (N_27544,N_20675,N_24567);
and U27545 (N_27545,N_20143,N_20898);
nor U27546 (N_27546,N_20390,N_23293);
and U27547 (N_27547,N_21242,N_22815);
or U27548 (N_27548,N_20779,N_24371);
xor U27549 (N_27549,N_21760,N_24229);
or U27550 (N_27550,N_20853,N_24310);
xor U27551 (N_27551,N_22173,N_20972);
nand U27552 (N_27552,N_20165,N_22459);
or U27553 (N_27553,N_20128,N_20364);
or U27554 (N_27554,N_20404,N_20284);
xnor U27555 (N_27555,N_22120,N_23262);
nor U27556 (N_27556,N_20744,N_22551);
nand U27557 (N_27557,N_23482,N_23251);
nor U27558 (N_27558,N_20850,N_22936);
xnor U27559 (N_27559,N_20196,N_20188);
nor U27560 (N_27560,N_21434,N_22372);
and U27561 (N_27561,N_24642,N_23313);
xor U27562 (N_27562,N_24486,N_22297);
nor U27563 (N_27563,N_20608,N_21515);
xnor U27564 (N_27564,N_23904,N_20990);
and U27565 (N_27565,N_20102,N_24337);
xnor U27566 (N_27566,N_20458,N_20023);
xnor U27567 (N_27567,N_20382,N_20553);
nor U27568 (N_27568,N_24936,N_20975);
xor U27569 (N_27569,N_22546,N_22498);
and U27570 (N_27570,N_22368,N_23177);
nor U27571 (N_27571,N_22187,N_23274);
and U27572 (N_27572,N_23439,N_23837);
or U27573 (N_27573,N_24303,N_23148);
xor U27574 (N_27574,N_24213,N_22497);
and U27575 (N_27575,N_22238,N_24488);
nor U27576 (N_27576,N_21970,N_20903);
xor U27577 (N_27577,N_23583,N_21313);
nor U27578 (N_27578,N_20712,N_20048);
and U27579 (N_27579,N_24011,N_20071);
xor U27580 (N_27580,N_20701,N_22726);
and U27581 (N_27581,N_23934,N_23352);
or U27582 (N_27582,N_22506,N_24379);
or U27583 (N_27583,N_23379,N_21489);
or U27584 (N_27584,N_20367,N_20379);
and U27585 (N_27585,N_23054,N_21915);
and U27586 (N_27586,N_23513,N_22192);
nor U27587 (N_27587,N_24653,N_20020);
xor U27588 (N_27588,N_20884,N_21531);
xor U27589 (N_27589,N_24026,N_24911);
nor U27590 (N_27590,N_22089,N_21749);
or U27591 (N_27591,N_23855,N_24705);
nor U27592 (N_27592,N_22499,N_21681);
nand U27593 (N_27593,N_24905,N_21234);
or U27594 (N_27594,N_24659,N_20450);
and U27595 (N_27595,N_23460,N_22867);
nand U27596 (N_27596,N_23657,N_24092);
xor U27597 (N_27597,N_23758,N_24387);
and U27598 (N_27598,N_24008,N_23205);
nor U27599 (N_27599,N_21211,N_21036);
nor U27600 (N_27600,N_24660,N_24823);
and U27601 (N_27601,N_20655,N_22808);
xnor U27602 (N_27602,N_23167,N_20584);
nor U27603 (N_27603,N_20533,N_21689);
or U27604 (N_27604,N_21538,N_20128);
or U27605 (N_27605,N_20550,N_20505);
nor U27606 (N_27606,N_20362,N_24095);
and U27607 (N_27607,N_22979,N_20732);
xor U27608 (N_27608,N_24956,N_21808);
or U27609 (N_27609,N_23392,N_23446);
nand U27610 (N_27610,N_23328,N_20630);
nand U27611 (N_27611,N_22916,N_23919);
nand U27612 (N_27612,N_20295,N_22759);
nor U27613 (N_27613,N_22170,N_20447);
xnor U27614 (N_27614,N_21256,N_23077);
xnor U27615 (N_27615,N_20102,N_23908);
xnor U27616 (N_27616,N_21122,N_21430);
or U27617 (N_27617,N_22414,N_20597);
and U27618 (N_27618,N_21249,N_21716);
nand U27619 (N_27619,N_20667,N_24412);
and U27620 (N_27620,N_20478,N_23201);
nor U27621 (N_27621,N_21413,N_21885);
xor U27622 (N_27622,N_24076,N_20065);
and U27623 (N_27623,N_23555,N_24525);
and U27624 (N_27624,N_24335,N_21502);
and U27625 (N_27625,N_20120,N_23962);
nand U27626 (N_27626,N_23160,N_22182);
nor U27627 (N_27627,N_23935,N_24805);
and U27628 (N_27628,N_24402,N_20310);
nor U27629 (N_27629,N_20932,N_24465);
nor U27630 (N_27630,N_21016,N_20014);
and U27631 (N_27631,N_20485,N_23005);
nand U27632 (N_27632,N_23304,N_21774);
and U27633 (N_27633,N_21270,N_24044);
nand U27634 (N_27634,N_23637,N_22259);
nand U27635 (N_27635,N_22571,N_21830);
nor U27636 (N_27636,N_20542,N_22711);
and U27637 (N_27637,N_22761,N_23595);
nand U27638 (N_27638,N_22818,N_23808);
and U27639 (N_27639,N_24321,N_22928);
and U27640 (N_27640,N_21971,N_21847);
nand U27641 (N_27641,N_23812,N_20243);
nand U27642 (N_27642,N_23686,N_21020);
nand U27643 (N_27643,N_21463,N_23493);
nor U27644 (N_27644,N_24652,N_21445);
and U27645 (N_27645,N_21894,N_21093);
and U27646 (N_27646,N_20996,N_22066);
xnor U27647 (N_27647,N_24116,N_22521);
nand U27648 (N_27648,N_22540,N_21253);
nor U27649 (N_27649,N_20943,N_23124);
and U27650 (N_27650,N_23020,N_21086);
xor U27651 (N_27651,N_22696,N_22615);
and U27652 (N_27652,N_21471,N_21076);
or U27653 (N_27653,N_21722,N_21638);
nor U27654 (N_27654,N_24666,N_21067);
and U27655 (N_27655,N_23337,N_21544);
xor U27656 (N_27656,N_20127,N_20254);
or U27657 (N_27657,N_21345,N_23019);
xor U27658 (N_27658,N_20374,N_24316);
nor U27659 (N_27659,N_24516,N_20576);
and U27660 (N_27660,N_24866,N_24069);
or U27661 (N_27661,N_23777,N_21908);
or U27662 (N_27662,N_20737,N_21413);
nor U27663 (N_27663,N_20679,N_23882);
xnor U27664 (N_27664,N_21878,N_20248);
nor U27665 (N_27665,N_24552,N_20307);
or U27666 (N_27666,N_22757,N_24892);
nand U27667 (N_27667,N_24966,N_20796);
or U27668 (N_27668,N_20046,N_20552);
nand U27669 (N_27669,N_21237,N_24270);
xnor U27670 (N_27670,N_24832,N_24249);
and U27671 (N_27671,N_24170,N_24189);
or U27672 (N_27672,N_22226,N_21134);
nand U27673 (N_27673,N_22561,N_24753);
nor U27674 (N_27674,N_22053,N_21017);
nor U27675 (N_27675,N_21817,N_22467);
nor U27676 (N_27676,N_23420,N_23709);
or U27677 (N_27677,N_20433,N_23631);
xor U27678 (N_27678,N_20185,N_23609);
xnor U27679 (N_27679,N_21103,N_20148);
xnor U27680 (N_27680,N_23669,N_20487);
nor U27681 (N_27681,N_22184,N_20289);
nor U27682 (N_27682,N_24235,N_22275);
nand U27683 (N_27683,N_20159,N_24087);
and U27684 (N_27684,N_23385,N_23263);
and U27685 (N_27685,N_23532,N_23859);
nand U27686 (N_27686,N_22393,N_22307);
xor U27687 (N_27687,N_24492,N_21655);
and U27688 (N_27688,N_24948,N_23256);
nor U27689 (N_27689,N_24051,N_22791);
xor U27690 (N_27690,N_23281,N_20111);
or U27691 (N_27691,N_22486,N_24637);
and U27692 (N_27692,N_24997,N_20137);
nand U27693 (N_27693,N_23957,N_24016);
and U27694 (N_27694,N_20679,N_23300);
xor U27695 (N_27695,N_24992,N_23495);
or U27696 (N_27696,N_20326,N_24483);
nand U27697 (N_27697,N_22148,N_22438);
nand U27698 (N_27698,N_23944,N_22538);
nand U27699 (N_27699,N_23752,N_24947);
or U27700 (N_27700,N_20187,N_22362);
nor U27701 (N_27701,N_20889,N_20322);
nor U27702 (N_27702,N_23849,N_21556);
xnor U27703 (N_27703,N_20730,N_24573);
xnor U27704 (N_27704,N_23007,N_21378);
nor U27705 (N_27705,N_20086,N_20625);
xnor U27706 (N_27706,N_21245,N_20249);
xnor U27707 (N_27707,N_20902,N_24222);
and U27708 (N_27708,N_24935,N_23627);
nand U27709 (N_27709,N_23099,N_22417);
nor U27710 (N_27710,N_23085,N_22760);
xnor U27711 (N_27711,N_22342,N_20289);
and U27712 (N_27712,N_20424,N_22655);
and U27713 (N_27713,N_20084,N_20729);
xnor U27714 (N_27714,N_23998,N_21358);
xor U27715 (N_27715,N_22604,N_20575);
and U27716 (N_27716,N_22898,N_24130);
and U27717 (N_27717,N_21569,N_24599);
nand U27718 (N_27718,N_20286,N_23261);
or U27719 (N_27719,N_20378,N_20909);
or U27720 (N_27720,N_24748,N_21730);
xnor U27721 (N_27721,N_23029,N_21055);
and U27722 (N_27722,N_23374,N_23681);
and U27723 (N_27723,N_24025,N_24722);
xor U27724 (N_27724,N_20045,N_20001);
nor U27725 (N_27725,N_20221,N_21304);
xnor U27726 (N_27726,N_22926,N_23030);
or U27727 (N_27727,N_22773,N_22890);
or U27728 (N_27728,N_23660,N_20616);
nand U27729 (N_27729,N_24722,N_24806);
and U27730 (N_27730,N_24846,N_23683);
xor U27731 (N_27731,N_20073,N_20265);
nor U27732 (N_27732,N_22180,N_24526);
nor U27733 (N_27733,N_20371,N_24759);
nor U27734 (N_27734,N_21211,N_24006);
xor U27735 (N_27735,N_22149,N_22423);
and U27736 (N_27736,N_24959,N_23802);
or U27737 (N_27737,N_21706,N_23437);
nor U27738 (N_27738,N_20893,N_20198);
nor U27739 (N_27739,N_20685,N_23599);
and U27740 (N_27740,N_24160,N_20792);
nor U27741 (N_27741,N_23616,N_22861);
xor U27742 (N_27742,N_22275,N_20659);
and U27743 (N_27743,N_24330,N_20617);
or U27744 (N_27744,N_22783,N_22769);
xnor U27745 (N_27745,N_20441,N_20284);
and U27746 (N_27746,N_24859,N_23775);
nand U27747 (N_27747,N_24103,N_23963);
nor U27748 (N_27748,N_24678,N_21874);
and U27749 (N_27749,N_22355,N_20585);
nand U27750 (N_27750,N_21014,N_24920);
xor U27751 (N_27751,N_22732,N_21535);
nand U27752 (N_27752,N_23936,N_23290);
or U27753 (N_27753,N_22350,N_23591);
and U27754 (N_27754,N_23627,N_24973);
nand U27755 (N_27755,N_21777,N_22138);
nor U27756 (N_27756,N_20553,N_21365);
nand U27757 (N_27757,N_21682,N_20551);
or U27758 (N_27758,N_22542,N_24196);
nand U27759 (N_27759,N_23078,N_23357);
xnor U27760 (N_27760,N_20153,N_21659);
nor U27761 (N_27761,N_22460,N_22325);
nor U27762 (N_27762,N_24501,N_22615);
nor U27763 (N_27763,N_24370,N_24840);
nor U27764 (N_27764,N_20687,N_24299);
and U27765 (N_27765,N_21644,N_24195);
and U27766 (N_27766,N_24068,N_20475);
nand U27767 (N_27767,N_22324,N_22577);
nand U27768 (N_27768,N_20858,N_21494);
or U27769 (N_27769,N_22257,N_22532);
nand U27770 (N_27770,N_22053,N_23923);
or U27771 (N_27771,N_23903,N_22740);
nand U27772 (N_27772,N_22592,N_23440);
or U27773 (N_27773,N_23054,N_24357);
nor U27774 (N_27774,N_23896,N_20810);
or U27775 (N_27775,N_21217,N_21798);
nor U27776 (N_27776,N_21938,N_22852);
or U27777 (N_27777,N_23210,N_24734);
and U27778 (N_27778,N_24649,N_23039);
or U27779 (N_27779,N_24562,N_23342);
xor U27780 (N_27780,N_22157,N_24072);
nand U27781 (N_27781,N_22258,N_24898);
xnor U27782 (N_27782,N_21225,N_21138);
nand U27783 (N_27783,N_24508,N_22853);
nor U27784 (N_27784,N_20400,N_24996);
and U27785 (N_27785,N_20666,N_20915);
nand U27786 (N_27786,N_23739,N_20271);
or U27787 (N_27787,N_22379,N_22568);
nor U27788 (N_27788,N_20357,N_24807);
or U27789 (N_27789,N_22012,N_20136);
or U27790 (N_27790,N_20290,N_21521);
or U27791 (N_27791,N_23584,N_23432);
and U27792 (N_27792,N_23754,N_20005);
nor U27793 (N_27793,N_20787,N_24549);
nor U27794 (N_27794,N_21000,N_22544);
nand U27795 (N_27795,N_23867,N_22031);
and U27796 (N_27796,N_22009,N_20552);
xnor U27797 (N_27797,N_22534,N_24655);
and U27798 (N_27798,N_23174,N_24372);
xnor U27799 (N_27799,N_24874,N_23251);
or U27800 (N_27800,N_23128,N_23562);
and U27801 (N_27801,N_21885,N_21978);
or U27802 (N_27802,N_20437,N_22952);
nor U27803 (N_27803,N_24435,N_23017);
nor U27804 (N_27804,N_23809,N_20912);
nor U27805 (N_27805,N_22861,N_24193);
nor U27806 (N_27806,N_24991,N_20202);
and U27807 (N_27807,N_20327,N_22071);
and U27808 (N_27808,N_23901,N_21261);
and U27809 (N_27809,N_20296,N_23968);
nand U27810 (N_27810,N_24879,N_21836);
or U27811 (N_27811,N_21081,N_24796);
xor U27812 (N_27812,N_21681,N_21799);
nor U27813 (N_27813,N_21822,N_20612);
nand U27814 (N_27814,N_20512,N_23177);
nor U27815 (N_27815,N_24470,N_20992);
xnor U27816 (N_27816,N_22263,N_20157);
xnor U27817 (N_27817,N_23928,N_23625);
or U27818 (N_27818,N_24744,N_22284);
nor U27819 (N_27819,N_22273,N_22761);
xnor U27820 (N_27820,N_23431,N_23205);
nand U27821 (N_27821,N_24160,N_24024);
nand U27822 (N_27822,N_22370,N_24438);
or U27823 (N_27823,N_22599,N_22176);
nand U27824 (N_27824,N_22413,N_22177);
or U27825 (N_27825,N_23192,N_22116);
nor U27826 (N_27826,N_22574,N_24822);
or U27827 (N_27827,N_22823,N_20429);
and U27828 (N_27828,N_20690,N_21836);
and U27829 (N_27829,N_22761,N_22703);
nand U27830 (N_27830,N_22812,N_23012);
and U27831 (N_27831,N_22450,N_23297);
nor U27832 (N_27832,N_21901,N_23794);
nand U27833 (N_27833,N_21740,N_23975);
nor U27834 (N_27834,N_22619,N_24190);
and U27835 (N_27835,N_23523,N_22100);
and U27836 (N_27836,N_23710,N_21189);
and U27837 (N_27837,N_23044,N_22315);
nor U27838 (N_27838,N_21792,N_21456);
or U27839 (N_27839,N_24581,N_23189);
xor U27840 (N_27840,N_23370,N_20711);
xor U27841 (N_27841,N_20367,N_20728);
nand U27842 (N_27842,N_20713,N_24695);
xnor U27843 (N_27843,N_24828,N_20496);
or U27844 (N_27844,N_24461,N_23708);
nor U27845 (N_27845,N_20032,N_24955);
or U27846 (N_27846,N_24997,N_23375);
and U27847 (N_27847,N_23037,N_20874);
nor U27848 (N_27848,N_24389,N_24966);
xnor U27849 (N_27849,N_21992,N_24414);
or U27850 (N_27850,N_22344,N_22215);
and U27851 (N_27851,N_21229,N_23944);
or U27852 (N_27852,N_20591,N_22920);
and U27853 (N_27853,N_20123,N_24233);
and U27854 (N_27854,N_24110,N_21888);
nor U27855 (N_27855,N_21434,N_23479);
nor U27856 (N_27856,N_22996,N_22135);
xor U27857 (N_27857,N_20321,N_24880);
and U27858 (N_27858,N_24758,N_23319);
xnor U27859 (N_27859,N_23268,N_23114);
and U27860 (N_27860,N_22590,N_22575);
or U27861 (N_27861,N_23564,N_24737);
and U27862 (N_27862,N_21119,N_23648);
nand U27863 (N_27863,N_22785,N_22899);
or U27864 (N_27864,N_24354,N_23275);
nor U27865 (N_27865,N_22714,N_20431);
and U27866 (N_27866,N_20534,N_24106);
and U27867 (N_27867,N_21938,N_23977);
or U27868 (N_27868,N_23847,N_20455);
and U27869 (N_27869,N_20872,N_24961);
nand U27870 (N_27870,N_22770,N_21217);
xor U27871 (N_27871,N_24688,N_22628);
nor U27872 (N_27872,N_23272,N_20174);
nand U27873 (N_27873,N_22074,N_21750);
nor U27874 (N_27874,N_24527,N_20885);
nor U27875 (N_27875,N_24460,N_22383);
xor U27876 (N_27876,N_23409,N_23331);
or U27877 (N_27877,N_24736,N_21088);
xnor U27878 (N_27878,N_24648,N_21642);
xor U27879 (N_27879,N_23238,N_20204);
and U27880 (N_27880,N_21574,N_22740);
nor U27881 (N_27881,N_21569,N_23682);
or U27882 (N_27882,N_21636,N_21257);
xor U27883 (N_27883,N_22542,N_23267);
xor U27884 (N_27884,N_21877,N_20074);
nor U27885 (N_27885,N_23393,N_22199);
nand U27886 (N_27886,N_23146,N_22785);
nor U27887 (N_27887,N_21386,N_22071);
and U27888 (N_27888,N_22973,N_23278);
nand U27889 (N_27889,N_21046,N_20855);
and U27890 (N_27890,N_23659,N_24947);
nor U27891 (N_27891,N_24249,N_22473);
xnor U27892 (N_27892,N_21221,N_21287);
or U27893 (N_27893,N_20880,N_23826);
nor U27894 (N_27894,N_22674,N_21043);
xnor U27895 (N_27895,N_24014,N_21012);
or U27896 (N_27896,N_20009,N_20436);
nor U27897 (N_27897,N_23210,N_23798);
nor U27898 (N_27898,N_22577,N_23997);
and U27899 (N_27899,N_22036,N_22684);
nand U27900 (N_27900,N_23751,N_22547);
and U27901 (N_27901,N_22899,N_20208);
xor U27902 (N_27902,N_24793,N_22535);
nand U27903 (N_27903,N_22738,N_20334);
or U27904 (N_27904,N_22870,N_21171);
nor U27905 (N_27905,N_22223,N_24864);
or U27906 (N_27906,N_24593,N_21337);
nor U27907 (N_27907,N_21244,N_24020);
and U27908 (N_27908,N_22347,N_23724);
or U27909 (N_27909,N_21185,N_20088);
or U27910 (N_27910,N_24948,N_20816);
xor U27911 (N_27911,N_22587,N_20702);
nand U27912 (N_27912,N_24108,N_21130);
and U27913 (N_27913,N_21133,N_21866);
nand U27914 (N_27914,N_22877,N_23678);
xnor U27915 (N_27915,N_24005,N_22148);
nor U27916 (N_27916,N_24544,N_24322);
or U27917 (N_27917,N_24657,N_24091);
nand U27918 (N_27918,N_21343,N_23828);
or U27919 (N_27919,N_22186,N_21123);
nand U27920 (N_27920,N_22387,N_22326);
nor U27921 (N_27921,N_24357,N_23600);
xor U27922 (N_27922,N_20809,N_23555);
and U27923 (N_27923,N_21998,N_20323);
and U27924 (N_27924,N_23420,N_22999);
xnor U27925 (N_27925,N_21438,N_22124);
and U27926 (N_27926,N_21694,N_23213);
nand U27927 (N_27927,N_23853,N_21509);
or U27928 (N_27928,N_24356,N_21419);
nor U27929 (N_27929,N_20902,N_20548);
or U27930 (N_27930,N_23535,N_23353);
nand U27931 (N_27931,N_23877,N_22372);
or U27932 (N_27932,N_24705,N_24282);
or U27933 (N_27933,N_20451,N_21498);
nand U27934 (N_27934,N_21834,N_21863);
nor U27935 (N_27935,N_23467,N_21690);
and U27936 (N_27936,N_20283,N_20295);
nand U27937 (N_27937,N_23513,N_24456);
nand U27938 (N_27938,N_20600,N_21979);
xor U27939 (N_27939,N_22403,N_22011);
nor U27940 (N_27940,N_22961,N_23679);
and U27941 (N_27941,N_20716,N_21317);
and U27942 (N_27942,N_23415,N_23226);
nand U27943 (N_27943,N_20941,N_22674);
or U27944 (N_27944,N_21267,N_22197);
or U27945 (N_27945,N_24824,N_24022);
or U27946 (N_27946,N_24218,N_23784);
nand U27947 (N_27947,N_21277,N_22914);
and U27948 (N_27948,N_22439,N_24146);
or U27949 (N_27949,N_21670,N_23632);
xor U27950 (N_27950,N_21552,N_24745);
and U27951 (N_27951,N_24735,N_23700);
nand U27952 (N_27952,N_24040,N_20787);
xnor U27953 (N_27953,N_22519,N_22071);
xor U27954 (N_27954,N_21309,N_20245);
and U27955 (N_27955,N_21671,N_24227);
and U27956 (N_27956,N_22723,N_22687);
xor U27957 (N_27957,N_20108,N_23047);
or U27958 (N_27958,N_21014,N_23678);
and U27959 (N_27959,N_21321,N_20048);
xor U27960 (N_27960,N_24490,N_22384);
or U27961 (N_27961,N_20786,N_23945);
xor U27962 (N_27962,N_24532,N_20221);
and U27963 (N_27963,N_22544,N_22568);
nand U27964 (N_27964,N_21145,N_20853);
xor U27965 (N_27965,N_24242,N_22785);
and U27966 (N_27966,N_21940,N_22445);
xor U27967 (N_27967,N_20249,N_20995);
or U27968 (N_27968,N_22033,N_23068);
and U27969 (N_27969,N_21614,N_22659);
nor U27970 (N_27970,N_22952,N_23772);
nor U27971 (N_27971,N_24361,N_24450);
or U27972 (N_27972,N_24362,N_20222);
nand U27973 (N_27973,N_23615,N_22998);
nor U27974 (N_27974,N_21248,N_22617);
nor U27975 (N_27975,N_20604,N_24026);
xor U27976 (N_27976,N_21163,N_21780);
nand U27977 (N_27977,N_22768,N_20848);
and U27978 (N_27978,N_23513,N_21093);
xor U27979 (N_27979,N_24057,N_21609);
xor U27980 (N_27980,N_21693,N_22359);
xnor U27981 (N_27981,N_23696,N_21513);
nor U27982 (N_27982,N_24706,N_21090);
nand U27983 (N_27983,N_20828,N_22572);
nand U27984 (N_27984,N_20227,N_23187);
or U27985 (N_27985,N_21766,N_24991);
nor U27986 (N_27986,N_23227,N_20721);
or U27987 (N_27987,N_21218,N_20440);
or U27988 (N_27988,N_23357,N_24968);
nor U27989 (N_27989,N_23918,N_20116);
or U27990 (N_27990,N_21577,N_23151);
xor U27991 (N_27991,N_20736,N_22253);
nor U27992 (N_27992,N_22480,N_20552);
or U27993 (N_27993,N_20307,N_20490);
nor U27994 (N_27994,N_21625,N_22263);
nor U27995 (N_27995,N_21806,N_23494);
xnor U27996 (N_27996,N_23481,N_22326);
nand U27997 (N_27997,N_20519,N_24548);
xnor U27998 (N_27998,N_20266,N_23451);
xor U27999 (N_27999,N_20202,N_21065);
xnor U28000 (N_28000,N_22853,N_20626);
and U28001 (N_28001,N_20893,N_23506);
and U28002 (N_28002,N_24660,N_21489);
nand U28003 (N_28003,N_20141,N_23863);
or U28004 (N_28004,N_20288,N_24402);
and U28005 (N_28005,N_22129,N_24677);
or U28006 (N_28006,N_24012,N_22003);
xnor U28007 (N_28007,N_20690,N_22380);
or U28008 (N_28008,N_22636,N_22165);
and U28009 (N_28009,N_20226,N_22080);
or U28010 (N_28010,N_23032,N_21805);
and U28011 (N_28011,N_21724,N_20680);
and U28012 (N_28012,N_24851,N_20911);
xnor U28013 (N_28013,N_24713,N_20820);
nor U28014 (N_28014,N_23533,N_23919);
or U28015 (N_28015,N_22221,N_20745);
nor U28016 (N_28016,N_23419,N_22716);
nand U28017 (N_28017,N_20044,N_20183);
nor U28018 (N_28018,N_21863,N_21535);
xnor U28019 (N_28019,N_22227,N_24797);
and U28020 (N_28020,N_23295,N_21626);
nand U28021 (N_28021,N_20114,N_21394);
and U28022 (N_28022,N_20767,N_24762);
or U28023 (N_28023,N_24028,N_24726);
nor U28024 (N_28024,N_21588,N_24429);
nor U28025 (N_28025,N_22660,N_24592);
nor U28026 (N_28026,N_20463,N_24176);
and U28027 (N_28027,N_21238,N_20372);
and U28028 (N_28028,N_21385,N_23178);
nand U28029 (N_28029,N_24484,N_21938);
or U28030 (N_28030,N_24136,N_23310);
nor U28031 (N_28031,N_21425,N_20310);
or U28032 (N_28032,N_20579,N_21685);
or U28033 (N_28033,N_21550,N_24249);
nor U28034 (N_28034,N_21360,N_22176);
and U28035 (N_28035,N_21848,N_22683);
and U28036 (N_28036,N_21131,N_24644);
nor U28037 (N_28037,N_20316,N_24081);
nand U28038 (N_28038,N_23053,N_24897);
and U28039 (N_28039,N_24787,N_21355);
and U28040 (N_28040,N_22536,N_22943);
and U28041 (N_28041,N_21166,N_21614);
and U28042 (N_28042,N_23541,N_21515);
xor U28043 (N_28043,N_24136,N_23558);
or U28044 (N_28044,N_24206,N_23102);
or U28045 (N_28045,N_24487,N_21395);
xnor U28046 (N_28046,N_23380,N_22810);
or U28047 (N_28047,N_22319,N_23664);
and U28048 (N_28048,N_20220,N_21689);
xnor U28049 (N_28049,N_21952,N_22016);
nand U28050 (N_28050,N_22296,N_22100);
nand U28051 (N_28051,N_23996,N_23901);
nor U28052 (N_28052,N_21580,N_22140);
nor U28053 (N_28053,N_21643,N_23746);
nand U28054 (N_28054,N_22830,N_20380);
nand U28055 (N_28055,N_20654,N_22862);
nand U28056 (N_28056,N_24738,N_21402);
xor U28057 (N_28057,N_23362,N_20163);
nand U28058 (N_28058,N_20883,N_21523);
and U28059 (N_28059,N_22190,N_24630);
xor U28060 (N_28060,N_24717,N_24523);
nand U28061 (N_28061,N_21158,N_20865);
or U28062 (N_28062,N_21569,N_24574);
nor U28063 (N_28063,N_24281,N_21741);
or U28064 (N_28064,N_20267,N_22843);
nand U28065 (N_28065,N_20040,N_21919);
or U28066 (N_28066,N_23020,N_20587);
or U28067 (N_28067,N_20614,N_23199);
nor U28068 (N_28068,N_23652,N_21245);
xor U28069 (N_28069,N_21495,N_20270);
nand U28070 (N_28070,N_22910,N_21003);
xor U28071 (N_28071,N_21978,N_22579);
nor U28072 (N_28072,N_24427,N_24023);
or U28073 (N_28073,N_22121,N_23236);
or U28074 (N_28074,N_24822,N_21945);
and U28075 (N_28075,N_22460,N_21871);
or U28076 (N_28076,N_20647,N_21987);
and U28077 (N_28077,N_20591,N_23606);
and U28078 (N_28078,N_21304,N_21310);
or U28079 (N_28079,N_22445,N_24199);
xor U28080 (N_28080,N_24783,N_24394);
nand U28081 (N_28081,N_23502,N_23142);
or U28082 (N_28082,N_24284,N_20131);
and U28083 (N_28083,N_21634,N_22825);
nand U28084 (N_28084,N_23193,N_24733);
nand U28085 (N_28085,N_22613,N_24444);
or U28086 (N_28086,N_20447,N_22200);
and U28087 (N_28087,N_20163,N_20390);
and U28088 (N_28088,N_22588,N_21708);
nand U28089 (N_28089,N_22111,N_20625);
or U28090 (N_28090,N_23738,N_24601);
and U28091 (N_28091,N_22521,N_23261);
nand U28092 (N_28092,N_24071,N_21152);
nand U28093 (N_28093,N_22191,N_21690);
xor U28094 (N_28094,N_24028,N_22077);
and U28095 (N_28095,N_22037,N_23918);
nand U28096 (N_28096,N_22939,N_20127);
nor U28097 (N_28097,N_24478,N_22091);
xnor U28098 (N_28098,N_23312,N_21035);
nor U28099 (N_28099,N_22005,N_22475);
nand U28100 (N_28100,N_24066,N_24091);
nor U28101 (N_28101,N_24217,N_22506);
nor U28102 (N_28102,N_23358,N_23898);
and U28103 (N_28103,N_22832,N_24985);
and U28104 (N_28104,N_23224,N_23899);
or U28105 (N_28105,N_22775,N_20231);
or U28106 (N_28106,N_22059,N_21223);
nand U28107 (N_28107,N_22889,N_22426);
xnor U28108 (N_28108,N_22419,N_22451);
and U28109 (N_28109,N_24302,N_23292);
xor U28110 (N_28110,N_23557,N_22487);
nor U28111 (N_28111,N_21821,N_23450);
nor U28112 (N_28112,N_21818,N_22010);
and U28113 (N_28113,N_22321,N_20008);
nor U28114 (N_28114,N_20448,N_20381);
or U28115 (N_28115,N_22829,N_23906);
and U28116 (N_28116,N_23132,N_23927);
or U28117 (N_28117,N_22072,N_20371);
or U28118 (N_28118,N_23737,N_21386);
xor U28119 (N_28119,N_20035,N_21169);
xnor U28120 (N_28120,N_22564,N_20643);
or U28121 (N_28121,N_22470,N_23840);
xor U28122 (N_28122,N_22038,N_24452);
xor U28123 (N_28123,N_21692,N_24780);
nor U28124 (N_28124,N_21987,N_24690);
xnor U28125 (N_28125,N_21358,N_20633);
and U28126 (N_28126,N_23225,N_21897);
nor U28127 (N_28127,N_24812,N_21108);
nand U28128 (N_28128,N_21267,N_23976);
and U28129 (N_28129,N_21677,N_22924);
and U28130 (N_28130,N_24922,N_21332);
xnor U28131 (N_28131,N_24172,N_20509);
nand U28132 (N_28132,N_24216,N_24059);
nor U28133 (N_28133,N_24506,N_22563);
and U28134 (N_28134,N_20133,N_22601);
nand U28135 (N_28135,N_24551,N_20122);
nand U28136 (N_28136,N_20056,N_20082);
and U28137 (N_28137,N_23973,N_24593);
nand U28138 (N_28138,N_23092,N_22303);
nor U28139 (N_28139,N_24155,N_23995);
or U28140 (N_28140,N_21325,N_20847);
xnor U28141 (N_28141,N_24369,N_22600);
or U28142 (N_28142,N_24453,N_23846);
nor U28143 (N_28143,N_21538,N_23938);
xor U28144 (N_28144,N_22389,N_21765);
and U28145 (N_28145,N_22951,N_24986);
xor U28146 (N_28146,N_20737,N_21320);
and U28147 (N_28147,N_20863,N_22825);
or U28148 (N_28148,N_20143,N_23451);
nor U28149 (N_28149,N_22263,N_24289);
and U28150 (N_28150,N_24127,N_23626);
and U28151 (N_28151,N_24151,N_22286);
or U28152 (N_28152,N_21159,N_21500);
or U28153 (N_28153,N_20412,N_20923);
or U28154 (N_28154,N_21312,N_21906);
nand U28155 (N_28155,N_21663,N_23946);
and U28156 (N_28156,N_21226,N_22370);
xor U28157 (N_28157,N_21449,N_22105);
nor U28158 (N_28158,N_21782,N_24958);
xnor U28159 (N_28159,N_23348,N_22664);
or U28160 (N_28160,N_23494,N_21004);
or U28161 (N_28161,N_21877,N_24903);
nand U28162 (N_28162,N_20861,N_22214);
nand U28163 (N_28163,N_22965,N_23012);
or U28164 (N_28164,N_20030,N_22337);
nand U28165 (N_28165,N_20878,N_22362);
or U28166 (N_28166,N_21231,N_21847);
and U28167 (N_28167,N_21865,N_20359);
nand U28168 (N_28168,N_23331,N_22812);
xnor U28169 (N_28169,N_22630,N_20970);
xor U28170 (N_28170,N_23491,N_20202);
and U28171 (N_28171,N_24294,N_21197);
nand U28172 (N_28172,N_24982,N_23633);
nand U28173 (N_28173,N_24663,N_20908);
xnor U28174 (N_28174,N_24165,N_20102);
and U28175 (N_28175,N_24156,N_23069);
xnor U28176 (N_28176,N_24245,N_20110);
nand U28177 (N_28177,N_21913,N_24734);
and U28178 (N_28178,N_22810,N_24559);
or U28179 (N_28179,N_21225,N_23682);
nand U28180 (N_28180,N_22605,N_20567);
nor U28181 (N_28181,N_23227,N_20811);
nand U28182 (N_28182,N_22539,N_24508);
xnor U28183 (N_28183,N_23283,N_24366);
nor U28184 (N_28184,N_21973,N_22364);
xnor U28185 (N_28185,N_24921,N_23246);
nor U28186 (N_28186,N_20771,N_21516);
nor U28187 (N_28187,N_22694,N_20682);
xor U28188 (N_28188,N_21951,N_21323);
nor U28189 (N_28189,N_22731,N_24853);
nor U28190 (N_28190,N_21910,N_21498);
and U28191 (N_28191,N_24516,N_20686);
or U28192 (N_28192,N_21024,N_24739);
or U28193 (N_28193,N_24191,N_22731);
and U28194 (N_28194,N_23673,N_21664);
xnor U28195 (N_28195,N_20959,N_24988);
or U28196 (N_28196,N_24484,N_20372);
xnor U28197 (N_28197,N_24031,N_21399);
xor U28198 (N_28198,N_24648,N_21688);
nor U28199 (N_28199,N_20319,N_21774);
nor U28200 (N_28200,N_23638,N_20979);
nor U28201 (N_28201,N_20242,N_22951);
nor U28202 (N_28202,N_20066,N_24588);
nor U28203 (N_28203,N_22688,N_24461);
or U28204 (N_28204,N_23668,N_23537);
nand U28205 (N_28205,N_21061,N_20246);
nand U28206 (N_28206,N_23760,N_20224);
xnor U28207 (N_28207,N_20267,N_23461);
and U28208 (N_28208,N_20020,N_24731);
xor U28209 (N_28209,N_22487,N_23944);
nand U28210 (N_28210,N_22849,N_23168);
nand U28211 (N_28211,N_22265,N_24417);
nor U28212 (N_28212,N_20381,N_21278);
or U28213 (N_28213,N_22309,N_24300);
or U28214 (N_28214,N_24261,N_20642);
and U28215 (N_28215,N_20958,N_24794);
xnor U28216 (N_28216,N_21452,N_22889);
xor U28217 (N_28217,N_20259,N_21321);
xnor U28218 (N_28218,N_22386,N_21616);
nand U28219 (N_28219,N_21720,N_21333);
and U28220 (N_28220,N_22301,N_22848);
and U28221 (N_28221,N_24073,N_22449);
nor U28222 (N_28222,N_24507,N_20880);
and U28223 (N_28223,N_21186,N_20241);
xor U28224 (N_28224,N_22834,N_24917);
or U28225 (N_28225,N_24134,N_20962);
and U28226 (N_28226,N_24632,N_23585);
nand U28227 (N_28227,N_22825,N_21272);
and U28228 (N_28228,N_21030,N_21526);
or U28229 (N_28229,N_20606,N_24819);
or U28230 (N_28230,N_21158,N_24510);
xor U28231 (N_28231,N_23338,N_22860);
and U28232 (N_28232,N_23036,N_22543);
xnor U28233 (N_28233,N_20977,N_20501);
nor U28234 (N_28234,N_21415,N_21703);
or U28235 (N_28235,N_24211,N_24759);
and U28236 (N_28236,N_21383,N_22888);
or U28237 (N_28237,N_23321,N_21396);
or U28238 (N_28238,N_23103,N_20853);
xnor U28239 (N_28239,N_21644,N_22386);
and U28240 (N_28240,N_24763,N_20884);
nand U28241 (N_28241,N_23952,N_24898);
or U28242 (N_28242,N_23742,N_20646);
or U28243 (N_28243,N_24755,N_20831);
nand U28244 (N_28244,N_22900,N_24249);
nand U28245 (N_28245,N_23154,N_20525);
nor U28246 (N_28246,N_20655,N_22011);
xnor U28247 (N_28247,N_22577,N_22771);
or U28248 (N_28248,N_23054,N_22210);
nor U28249 (N_28249,N_22573,N_20229);
and U28250 (N_28250,N_24884,N_24332);
and U28251 (N_28251,N_20949,N_24089);
nor U28252 (N_28252,N_20336,N_21885);
xor U28253 (N_28253,N_20423,N_20730);
nand U28254 (N_28254,N_23686,N_20040);
nor U28255 (N_28255,N_22261,N_24153);
xor U28256 (N_28256,N_22518,N_20352);
nand U28257 (N_28257,N_24340,N_23055);
nand U28258 (N_28258,N_22993,N_23439);
nor U28259 (N_28259,N_23449,N_22511);
or U28260 (N_28260,N_23620,N_23182);
or U28261 (N_28261,N_22007,N_21516);
xnor U28262 (N_28262,N_24552,N_21532);
and U28263 (N_28263,N_24893,N_22125);
or U28264 (N_28264,N_21551,N_21999);
and U28265 (N_28265,N_23949,N_21709);
or U28266 (N_28266,N_23790,N_21701);
xor U28267 (N_28267,N_22189,N_21188);
and U28268 (N_28268,N_24788,N_23651);
or U28269 (N_28269,N_20921,N_24500);
and U28270 (N_28270,N_21688,N_23267);
xor U28271 (N_28271,N_21619,N_23292);
or U28272 (N_28272,N_23668,N_23965);
nand U28273 (N_28273,N_23729,N_21948);
and U28274 (N_28274,N_22679,N_23024);
or U28275 (N_28275,N_20312,N_24451);
xnor U28276 (N_28276,N_23086,N_21898);
nor U28277 (N_28277,N_23032,N_20797);
or U28278 (N_28278,N_22565,N_24318);
xnor U28279 (N_28279,N_22795,N_22502);
or U28280 (N_28280,N_20831,N_22380);
xnor U28281 (N_28281,N_20369,N_20726);
xor U28282 (N_28282,N_24134,N_21122);
nor U28283 (N_28283,N_22906,N_24911);
and U28284 (N_28284,N_21733,N_24204);
xnor U28285 (N_28285,N_23809,N_23728);
or U28286 (N_28286,N_20823,N_21336);
or U28287 (N_28287,N_20067,N_21141);
nor U28288 (N_28288,N_21235,N_22949);
and U28289 (N_28289,N_22372,N_20861);
or U28290 (N_28290,N_23973,N_22282);
nand U28291 (N_28291,N_23417,N_22829);
nand U28292 (N_28292,N_20213,N_22318);
or U28293 (N_28293,N_22586,N_22349);
or U28294 (N_28294,N_21580,N_21824);
nor U28295 (N_28295,N_21504,N_22179);
and U28296 (N_28296,N_21371,N_23548);
xnor U28297 (N_28297,N_20790,N_24154);
or U28298 (N_28298,N_21810,N_23068);
or U28299 (N_28299,N_21323,N_21533);
nor U28300 (N_28300,N_24588,N_21198);
nand U28301 (N_28301,N_20965,N_22607);
nor U28302 (N_28302,N_23429,N_20806);
nor U28303 (N_28303,N_23240,N_22764);
and U28304 (N_28304,N_21100,N_20072);
nand U28305 (N_28305,N_21360,N_23898);
and U28306 (N_28306,N_20555,N_22894);
xor U28307 (N_28307,N_22270,N_21086);
nor U28308 (N_28308,N_20957,N_24334);
nand U28309 (N_28309,N_24557,N_22106);
nor U28310 (N_28310,N_23670,N_21059);
nor U28311 (N_28311,N_21051,N_21017);
or U28312 (N_28312,N_20550,N_21496);
nor U28313 (N_28313,N_20904,N_24599);
nand U28314 (N_28314,N_22753,N_20561);
nand U28315 (N_28315,N_23086,N_20190);
or U28316 (N_28316,N_22245,N_21151);
or U28317 (N_28317,N_24597,N_22595);
xnor U28318 (N_28318,N_20650,N_24572);
nor U28319 (N_28319,N_21183,N_24473);
nor U28320 (N_28320,N_21902,N_23680);
nand U28321 (N_28321,N_24681,N_20085);
or U28322 (N_28322,N_21039,N_22277);
or U28323 (N_28323,N_22671,N_22344);
xor U28324 (N_28324,N_20981,N_23756);
nand U28325 (N_28325,N_22107,N_21486);
or U28326 (N_28326,N_23711,N_24661);
xnor U28327 (N_28327,N_24396,N_23261);
xnor U28328 (N_28328,N_20099,N_20060);
nor U28329 (N_28329,N_21765,N_23770);
or U28330 (N_28330,N_21070,N_22433);
or U28331 (N_28331,N_20904,N_20028);
or U28332 (N_28332,N_21618,N_20752);
nor U28333 (N_28333,N_23705,N_20583);
nand U28334 (N_28334,N_21518,N_22148);
and U28335 (N_28335,N_22617,N_20385);
nor U28336 (N_28336,N_23689,N_22246);
nand U28337 (N_28337,N_21970,N_22113);
or U28338 (N_28338,N_22764,N_23468);
nand U28339 (N_28339,N_22135,N_21560);
xor U28340 (N_28340,N_23111,N_20355);
nand U28341 (N_28341,N_23568,N_22067);
nand U28342 (N_28342,N_23363,N_24373);
and U28343 (N_28343,N_23607,N_20940);
or U28344 (N_28344,N_20277,N_22706);
nand U28345 (N_28345,N_21411,N_21476);
or U28346 (N_28346,N_24380,N_20480);
xor U28347 (N_28347,N_20960,N_20397);
and U28348 (N_28348,N_22408,N_22893);
or U28349 (N_28349,N_24479,N_20387);
xnor U28350 (N_28350,N_24181,N_21673);
and U28351 (N_28351,N_24662,N_22733);
nand U28352 (N_28352,N_23148,N_23140);
xnor U28353 (N_28353,N_23520,N_22948);
and U28354 (N_28354,N_24297,N_21615);
or U28355 (N_28355,N_23404,N_20382);
nor U28356 (N_28356,N_21073,N_22606);
or U28357 (N_28357,N_24790,N_20144);
and U28358 (N_28358,N_23896,N_23886);
xnor U28359 (N_28359,N_21912,N_21600);
nand U28360 (N_28360,N_20590,N_24611);
and U28361 (N_28361,N_22559,N_24712);
and U28362 (N_28362,N_24740,N_23729);
nand U28363 (N_28363,N_24618,N_24931);
and U28364 (N_28364,N_21761,N_22222);
nand U28365 (N_28365,N_22030,N_22136);
nor U28366 (N_28366,N_21250,N_23369);
xor U28367 (N_28367,N_21850,N_22385);
and U28368 (N_28368,N_24835,N_23601);
nor U28369 (N_28369,N_21043,N_22029);
xor U28370 (N_28370,N_23617,N_20969);
or U28371 (N_28371,N_24870,N_24826);
and U28372 (N_28372,N_23993,N_23337);
xor U28373 (N_28373,N_21262,N_24670);
nand U28374 (N_28374,N_24478,N_21272);
or U28375 (N_28375,N_21359,N_23983);
nor U28376 (N_28376,N_21572,N_24077);
nand U28377 (N_28377,N_22800,N_24231);
nand U28378 (N_28378,N_22015,N_20984);
and U28379 (N_28379,N_23842,N_23855);
nor U28380 (N_28380,N_20429,N_20803);
xnor U28381 (N_28381,N_21316,N_20358);
and U28382 (N_28382,N_22592,N_21702);
and U28383 (N_28383,N_23116,N_22428);
and U28384 (N_28384,N_23902,N_20338);
and U28385 (N_28385,N_23381,N_23738);
xor U28386 (N_28386,N_21675,N_20662);
nor U28387 (N_28387,N_22023,N_21802);
and U28388 (N_28388,N_22668,N_20245);
nand U28389 (N_28389,N_22734,N_20559);
nor U28390 (N_28390,N_20571,N_21878);
nand U28391 (N_28391,N_22714,N_21328);
xnor U28392 (N_28392,N_22574,N_21551);
xor U28393 (N_28393,N_22476,N_23757);
or U28394 (N_28394,N_23673,N_24109);
or U28395 (N_28395,N_22267,N_20101);
or U28396 (N_28396,N_21469,N_24482);
nand U28397 (N_28397,N_24832,N_21001);
nor U28398 (N_28398,N_24194,N_21370);
nor U28399 (N_28399,N_20562,N_21807);
and U28400 (N_28400,N_22075,N_21547);
xnor U28401 (N_28401,N_24178,N_20887);
nand U28402 (N_28402,N_21325,N_21618);
nand U28403 (N_28403,N_23253,N_23936);
and U28404 (N_28404,N_23615,N_22565);
xnor U28405 (N_28405,N_20116,N_21618);
nor U28406 (N_28406,N_20140,N_21309);
and U28407 (N_28407,N_22768,N_23646);
xor U28408 (N_28408,N_24895,N_21787);
nand U28409 (N_28409,N_21584,N_22876);
or U28410 (N_28410,N_20465,N_22105);
or U28411 (N_28411,N_23067,N_20302);
nand U28412 (N_28412,N_23310,N_21508);
or U28413 (N_28413,N_24907,N_23738);
or U28414 (N_28414,N_24308,N_22656);
and U28415 (N_28415,N_22048,N_21354);
nand U28416 (N_28416,N_21153,N_22044);
or U28417 (N_28417,N_24597,N_21558);
or U28418 (N_28418,N_22256,N_20799);
and U28419 (N_28419,N_23688,N_23297);
xor U28420 (N_28420,N_22330,N_22366);
and U28421 (N_28421,N_21367,N_22526);
nand U28422 (N_28422,N_23434,N_22873);
nand U28423 (N_28423,N_24907,N_21061);
nand U28424 (N_28424,N_21479,N_21727);
and U28425 (N_28425,N_23301,N_20888);
nor U28426 (N_28426,N_22762,N_22325);
and U28427 (N_28427,N_22450,N_24711);
nand U28428 (N_28428,N_20678,N_23165);
nor U28429 (N_28429,N_20073,N_24562);
nand U28430 (N_28430,N_24199,N_20239);
and U28431 (N_28431,N_22652,N_23708);
nor U28432 (N_28432,N_21085,N_24273);
nand U28433 (N_28433,N_23801,N_21155);
or U28434 (N_28434,N_22136,N_21374);
or U28435 (N_28435,N_22783,N_20961);
xor U28436 (N_28436,N_24495,N_20421);
nor U28437 (N_28437,N_20335,N_20151);
nand U28438 (N_28438,N_23099,N_22778);
nand U28439 (N_28439,N_20110,N_21896);
or U28440 (N_28440,N_20419,N_22771);
and U28441 (N_28441,N_20055,N_24867);
or U28442 (N_28442,N_23789,N_20763);
or U28443 (N_28443,N_24308,N_20821);
nor U28444 (N_28444,N_20164,N_20851);
xnor U28445 (N_28445,N_22199,N_22783);
nand U28446 (N_28446,N_24534,N_23817);
and U28447 (N_28447,N_20949,N_21662);
nand U28448 (N_28448,N_20015,N_22140);
nor U28449 (N_28449,N_20205,N_21291);
xnor U28450 (N_28450,N_24695,N_20392);
xnor U28451 (N_28451,N_21844,N_23905);
or U28452 (N_28452,N_24972,N_24185);
xor U28453 (N_28453,N_22181,N_21467);
nor U28454 (N_28454,N_21231,N_20382);
xnor U28455 (N_28455,N_21275,N_22451);
or U28456 (N_28456,N_22790,N_23670);
nor U28457 (N_28457,N_24927,N_24422);
xnor U28458 (N_28458,N_20844,N_22174);
xor U28459 (N_28459,N_20868,N_20251);
and U28460 (N_28460,N_21069,N_21635);
nor U28461 (N_28461,N_21610,N_20405);
or U28462 (N_28462,N_22806,N_23957);
nor U28463 (N_28463,N_20157,N_22649);
and U28464 (N_28464,N_23064,N_24099);
or U28465 (N_28465,N_20771,N_23397);
and U28466 (N_28466,N_23202,N_21323);
or U28467 (N_28467,N_22161,N_21246);
nor U28468 (N_28468,N_21558,N_22203);
and U28469 (N_28469,N_22785,N_23726);
or U28470 (N_28470,N_20071,N_22015);
nor U28471 (N_28471,N_23523,N_21361);
and U28472 (N_28472,N_24545,N_21526);
xor U28473 (N_28473,N_24206,N_21000);
nand U28474 (N_28474,N_22838,N_24153);
or U28475 (N_28475,N_24439,N_24297);
and U28476 (N_28476,N_21555,N_21093);
and U28477 (N_28477,N_20714,N_24178);
nor U28478 (N_28478,N_20915,N_22006);
nand U28479 (N_28479,N_24741,N_20273);
or U28480 (N_28480,N_20367,N_21828);
nand U28481 (N_28481,N_21147,N_20512);
nor U28482 (N_28482,N_20506,N_24283);
or U28483 (N_28483,N_22678,N_24597);
or U28484 (N_28484,N_22211,N_22061);
xnor U28485 (N_28485,N_22344,N_22045);
xnor U28486 (N_28486,N_22550,N_20555);
nor U28487 (N_28487,N_22218,N_24551);
nand U28488 (N_28488,N_22651,N_20041);
xor U28489 (N_28489,N_23049,N_22254);
and U28490 (N_28490,N_20556,N_20808);
and U28491 (N_28491,N_24061,N_24897);
and U28492 (N_28492,N_21314,N_21742);
nand U28493 (N_28493,N_21961,N_20880);
and U28494 (N_28494,N_23879,N_23141);
nor U28495 (N_28495,N_23809,N_24477);
or U28496 (N_28496,N_22194,N_20451);
xor U28497 (N_28497,N_21128,N_20096);
and U28498 (N_28498,N_23526,N_23926);
or U28499 (N_28499,N_20199,N_24306);
or U28500 (N_28500,N_23824,N_22914);
nand U28501 (N_28501,N_21493,N_24156);
xnor U28502 (N_28502,N_20351,N_22406);
xor U28503 (N_28503,N_21623,N_21663);
nand U28504 (N_28504,N_23313,N_20350);
nand U28505 (N_28505,N_22290,N_21021);
xor U28506 (N_28506,N_21862,N_22605);
nor U28507 (N_28507,N_23745,N_22771);
nand U28508 (N_28508,N_20819,N_22285);
or U28509 (N_28509,N_24023,N_20147);
and U28510 (N_28510,N_24685,N_20680);
or U28511 (N_28511,N_22702,N_23550);
xnor U28512 (N_28512,N_20610,N_21353);
xor U28513 (N_28513,N_21044,N_22175);
or U28514 (N_28514,N_21465,N_22515);
xor U28515 (N_28515,N_23342,N_24350);
and U28516 (N_28516,N_22027,N_21795);
and U28517 (N_28517,N_23502,N_23208);
and U28518 (N_28518,N_22016,N_23881);
nand U28519 (N_28519,N_21570,N_20517);
nor U28520 (N_28520,N_23430,N_22596);
and U28521 (N_28521,N_20655,N_22252);
nor U28522 (N_28522,N_24585,N_20795);
or U28523 (N_28523,N_23731,N_24704);
and U28524 (N_28524,N_22984,N_23655);
or U28525 (N_28525,N_21198,N_24618);
nand U28526 (N_28526,N_23351,N_21656);
nor U28527 (N_28527,N_24335,N_22192);
and U28528 (N_28528,N_24326,N_22800);
xnor U28529 (N_28529,N_20545,N_21363);
xnor U28530 (N_28530,N_24662,N_22180);
and U28531 (N_28531,N_21113,N_23205);
or U28532 (N_28532,N_23570,N_24422);
nand U28533 (N_28533,N_20171,N_22936);
and U28534 (N_28534,N_21572,N_20028);
and U28535 (N_28535,N_20448,N_22962);
and U28536 (N_28536,N_23607,N_21538);
nand U28537 (N_28537,N_23092,N_23082);
and U28538 (N_28538,N_24612,N_24683);
xnor U28539 (N_28539,N_21212,N_20665);
or U28540 (N_28540,N_21262,N_24472);
nand U28541 (N_28541,N_24399,N_21658);
and U28542 (N_28542,N_21750,N_20414);
or U28543 (N_28543,N_23480,N_21862);
and U28544 (N_28544,N_23936,N_20243);
or U28545 (N_28545,N_23456,N_24425);
nand U28546 (N_28546,N_24091,N_22962);
nand U28547 (N_28547,N_24163,N_21586);
or U28548 (N_28548,N_24561,N_21108);
nand U28549 (N_28549,N_23509,N_20814);
xnor U28550 (N_28550,N_23589,N_20222);
xor U28551 (N_28551,N_22076,N_23539);
xnor U28552 (N_28552,N_22772,N_20037);
or U28553 (N_28553,N_20693,N_23218);
or U28554 (N_28554,N_20273,N_21390);
nor U28555 (N_28555,N_23977,N_21812);
nor U28556 (N_28556,N_23357,N_23251);
nor U28557 (N_28557,N_24902,N_23943);
xnor U28558 (N_28558,N_21416,N_20257);
nand U28559 (N_28559,N_23987,N_20777);
and U28560 (N_28560,N_21277,N_24570);
nand U28561 (N_28561,N_23442,N_20724);
nor U28562 (N_28562,N_20477,N_22200);
nor U28563 (N_28563,N_20571,N_20364);
or U28564 (N_28564,N_24594,N_21968);
and U28565 (N_28565,N_22082,N_23829);
and U28566 (N_28566,N_20337,N_22059);
or U28567 (N_28567,N_22153,N_20867);
nand U28568 (N_28568,N_23483,N_23841);
nor U28569 (N_28569,N_22090,N_20121);
and U28570 (N_28570,N_24278,N_20499);
nand U28571 (N_28571,N_24499,N_23051);
and U28572 (N_28572,N_22448,N_21728);
nor U28573 (N_28573,N_24894,N_22635);
nor U28574 (N_28574,N_20246,N_20977);
or U28575 (N_28575,N_23470,N_20508);
nand U28576 (N_28576,N_23208,N_20442);
xnor U28577 (N_28577,N_21412,N_24809);
or U28578 (N_28578,N_24439,N_23812);
or U28579 (N_28579,N_22542,N_23467);
or U28580 (N_28580,N_24319,N_22777);
or U28581 (N_28581,N_22885,N_22266);
nor U28582 (N_28582,N_24462,N_20802);
nand U28583 (N_28583,N_21359,N_24117);
xor U28584 (N_28584,N_22076,N_23953);
and U28585 (N_28585,N_23624,N_21939);
and U28586 (N_28586,N_23278,N_21180);
xor U28587 (N_28587,N_21515,N_22504);
nor U28588 (N_28588,N_23553,N_22443);
nand U28589 (N_28589,N_21476,N_23549);
nand U28590 (N_28590,N_23358,N_23978);
nor U28591 (N_28591,N_23314,N_23795);
nor U28592 (N_28592,N_21038,N_21465);
xnor U28593 (N_28593,N_21953,N_20252);
nand U28594 (N_28594,N_20198,N_21178);
and U28595 (N_28595,N_20236,N_20722);
and U28596 (N_28596,N_23877,N_23875);
nand U28597 (N_28597,N_21391,N_22409);
and U28598 (N_28598,N_24697,N_23387);
xnor U28599 (N_28599,N_20148,N_22472);
nand U28600 (N_28600,N_21579,N_22309);
nand U28601 (N_28601,N_20323,N_24192);
nor U28602 (N_28602,N_22235,N_22927);
xor U28603 (N_28603,N_20085,N_22007);
or U28604 (N_28604,N_20144,N_23431);
nand U28605 (N_28605,N_24546,N_20602);
nand U28606 (N_28606,N_24970,N_22216);
xnor U28607 (N_28607,N_20310,N_20488);
nor U28608 (N_28608,N_20743,N_24768);
nand U28609 (N_28609,N_20543,N_24532);
nor U28610 (N_28610,N_21991,N_20588);
and U28611 (N_28611,N_24648,N_24042);
xnor U28612 (N_28612,N_23044,N_20252);
and U28613 (N_28613,N_21731,N_22761);
and U28614 (N_28614,N_23440,N_20479);
nor U28615 (N_28615,N_22681,N_21093);
xor U28616 (N_28616,N_20854,N_20819);
or U28617 (N_28617,N_20160,N_24878);
nor U28618 (N_28618,N_24527,N_20946);
nand U28619 (N_28619,N_22957,N_24851);
or U28620 (N_28620,N_21808,N_21732);
nor U28621 (N_28621,N_21744,N_23027);
or U28622 (N_28622,N_21247,N_22187);
nand U28623 (N_28623,N_22983,N_20193);
nand U28624 (N_28624,N_20521,N_22456);
xnor U28625 (N_28625,N_24925,N_23515);
xor U28626 (N_28626,N_21576,N_24221);
xnor U28627 (N_28627,N_23587,N_20015);
nor U28628 (N_28628,N_20103,N_24550);
nor U28629 (N_28629,N_22409,N_20971);
and U28630 (N_28630,N_20525,N_20390);
nor U28631 (N_28631,N_23999,N_22816);
or U28632 (N_28632,N_20996,N_23801);
xor U28633 (N_28633,N_24264,N_20063);
nor U28634 (N_28634,N_20040,N_24921);
xnor U28635 (N_28635,N_23249,N_20810);
nand U28636 (N_28636,N_23216,N_23770);
xor U28637 (N_28637,N_24590,N_20752);
or U28638 (N_28638,N_23715,N_23989);
nand U28639 (N_28639,N_22474,N_20240);
nor U28640 (N_28640,N_20013,N_24817);
and U28641 (N_28641,N_24375,N_21902);
nand U28642 (N_28642,N_23479,N_22491);
nand U28643 (N_28643,N_20002,N_22956);
xnor U28644 (N_28644,N_21434,N_21091);
nor U28645 (N_28645,N_22490,N_21136);
or U28646 (N_28646,N_23345,N_24309);
nor U28647 (N_28647,N_22948,N_23441);
xnor U28648 (N_28648,N_23602,N_24884);
or U28649 (N_28649,N_21388,N_21478);
and U28650 (N_28650,N_20720,N_21576);
and U28651 (N_28651,N_23952,N_20564);
nand U28652 (N_28652,N_21851,N_24353);
nor U28653 (N_28653,N_22987,N_21958);
nand U28654 (N_28654,N_22339,N_23209);
or U28655 (N_28655,N_23089,N_20599);
nor U28656 (N_28656,N_21856,N_20809);
or U28657 (N_28657,N_20938,N_22588);
or U28658 (N_28658,N_20398,N_22718);
nand U28659 (N_28659,N_20741,N_21114);
xor U28660 (N_28660,N_21584,N_23752);
and U28661 (N_28661,N_21038,N_21130);
and U28662 (N_28662,N_23363,N_24508);
nand U28663 (N_28663,N_21675,N_20380);
and U28664 (N_28664,N_24855,N_22640);
nor U28665 (N_28665,N_20724,N_22396);
and U28666 (N_28666,N_20892,N_20350);
nand U28667 (N_28667,N_24989,N_23532);
nand U28668 (N_28668,N_24195,N_22484);
or U28669 (N_28669,N_24883,N_20369);
nand U28670 (N_28670,N_21191,N_23416);
xor U28671 (N_28671,N_22139,N_20316);
nor U28672 (N_28672,N_20689,N_21516);
or U28673 (N_28673,N_20704,N_24071);
nor U28674 (N_28674,N_22432,N_23754);
and U28675 (N_28675,N_24714,N_23811);
nand U28676 (N_28676,N_21189,N_22828);
nand U28677 (N_28677,N_22917,N_22740);
nand U28678 (N_28678,N_22476,N_20213);
nor U28679 (N_28679,N_21730,N_23613);
and U28680 (N_28680,N_21821,N_22145);
nor U28681 (N_28681,N_24040,N_23671);
xor U28682 (N_28682,N_23106,N_20514);
xnor U28683 (N_28683,N_24677,N_22543);
nand U28684 (N_28684,N_24696,N_24250);
and U28685 (N_28685,N_23842,N_23664);
xnor U28686 (N_28686,N_24201,N_20152);
and U28687 (N_28687,N_20919,N_20589);
nand U28688 (N_28688,N_20144,N_20224);
nor U28689 (N_28689,N_20310,N_24663);
nand U28690 (N_28690,N_23947,N_23489);
nand U28691 (N_28691,N_24590,N_24426);
and U28692 (N_28692,N_21115,N_23833);
nor U28693 (N_28693,N_21193,N_21889);
nand U28694 (N_28694,N_24296,N_24866);
xnor U28695 (N_28695,N_24203,N_23005);
and U28696 (N_28696,N_21368,N_22763);
xor U28697 (N_28697,N_20767,N_22798);
nand U28698 (N_28698,N_21227,N_20455);
or U28699 (N_28699,N_22009,N_20013);
and U28700 (N_28700,N_24738,N_20961);
or U28701 (N_28701,N_24589,N_21894);
xnor U28702 (N_28702,N_22926,N_22630);
xnor U28703 (N_28703,N_22018,N_23281);
or U28704 (N_28704,N_21162,N_24924);
or U28705 (N_28705,N_22638,N_24949);
and U28706 (N_28706,N_20889,N_21182);
or U28707 (N_28707,N_23934,N_22279);
nand U28708 (N_28708,N_24033,N_22954);
xor U28709 (N_28709,N_22858,N_23181);
nor U28710 (N_28710,N_22703,N_24829);
xor U28711 (N_28711,N_24044,N_20871);
and U28712 (N_28712,N_22662,N_21763);
or U28713 (N_28713,N_24809,N_24267);
or U28714 (N_28714,N_23107,N_21674);
nor U28715 (N_28715,N_23034,N_20883);
and U28716 (N_28716,N_24837,N_23962);
or U28717 (N_28717,N_21992,N_22246);
nor U28718 (N_28718,N_22087,N_20623);
or U28719 (N_28719,N_23994,N_24004);
nor U28720 (N_28720,N_22974,N_20869);
and U28721 (N_28721,N_23055,N_23695);
nor U28722 (N_28722,N_22381,N_20142);
nand U28723 (N_28723,N_20391,N_21323);
nor U28724 (N_28724,N_21305,N_21308);
nor U28725 (N_28725,N_20629,N_20735);
nor U28726 (N_28726,N_24735,N_21644);
nor U28727 (N_28727,N_21351,N_20319);
nor U28728 (N_28728,N_20822,N_22383);
and U28729 (N_28729,N_24907,N_22439);
nand U28730 (N_28730,N_22115,N_23002);
nand U28731 (N_28731,N_23555,N_23430);
xor U28732 (N_28732,N_20472,N_23834);
or U28733 (N_28733,N_20621,N_20980);
and U28734 (N_28734,N_23329,N_23828);
xor U28735 (N_28735,N_21296,N_22625);
and U28736 (N_28736,N_20708,N_23191);
and U28737 (N_28737,N_23814,N_23510);
xor U28738 (N_28738,N_24099,N_21047);
nand U28739 (N_28739,N_21828,N_21820);
xnor U28740 (N_28740,N_21568,N_20023);
xnor U28741 (N_28741,N_21431,N_24353);
and U28742 (N_28742,N_22426,N_21777);
nor U28743 (N_28743,N_23943,N_24800);
or U28744 (N_28744,N_20787,N_22621);
or U28745 (N_28745,N_22607,N_24260);
nand U28746 (N_28746,N_24544,N_23796);
xor U28747 (N_28747,N_22313,N_24724);
nand U28748 (N_28748,N_23700,N_21025);
nand U28749 (N_28749,N_23186,N_20257);
nor U28750 (N_28750,N_21246,N_20436);
or U28751 (N_28751,N_21573,N_20551);
nand U28752 (N_28752,N_20453,N_21090);
or U28753 (N_28753,N_22858,N_24547);
xor U28754 (N_28754,N_22555,N_23260);
nand U28755 (N_28755,N_20734,N_20799);
nand U28756 (N_28756,N_22540,N_24198);
nand U28757 (N_28757,N_20982,N_23652);
or U28758 (N_28758,N_20211,N_23584);
or U28759 (N_28759,N_24989,N_24469);
xor U28760 (N_28760,N_23267,N_21863);
or U28761 (N_28761,N_21814,N_24554);
xnor U28762 (N_28762,N_20480,N_24386);
xor U28763 (N_28763,N_24365,N_24639);
xor U28764 (N_28764,N_24810,N_23858);
or U28765 (N_28765,N_22591,N_22950);
nor U28766 (N_28766,N_23411,N_23516);
xor U28767 (N_28767,N_24508,N_22627);
nand U28768 (N_28768,N_20684,N_21480);
or U28769 (N_28769,N_21953,N_24522);
xnor U28770 (N_28770,N_22013,N_24910);
and U28771 (N_28771,N_21271,N_22249);
xnor U28772 (N_28772,N_22327,N_23446);
or U28773 (N_28773,N_22499,N_23739);
nor U28774 (N_28774,N_22343,N_22440);
xnor U28775 (N_28775,N_20711,N_23789);
nand U28776 (N_28776,N_20009,N_23776);
or U28777 (N_28777,N_21828,N_23510);
and U28778 (N_28778,N_20931,N_20420);
nor U28779 (N_28779,N_20824,N_23378);
nand U28780 (N_28780,N_20367,N_21970);
nor U28781 (N_28781,N_21473,N_21190);
or U28782 (N_28782,N_20498,N_22152);
nor U28783 (N_28783,N_24866,N_23356);
xnor U28784 (N_28784,N_24736,N_22560);
and U28785 (N_28785,N_22286,N_22092);
or U28786 (N_28786,N_23628,N_21584);
or U28787 (N_28787,N_24563,N_23943);
xnor U28788 (N_28788,N_20703,N_21711);
or U28789 (N_28789,N_22625,N_21890);
and U28790 (N_28790,N_20188,N_21756);
nand U28791 (N_28791,N_23290,N_22430);
or U28792 (N_28792,N_24495,N_20150);
and U28793 (N_28793,N_22408,N_20805);
and U28794 (N_28794,N_22741,N_23176);
or U28795 (N_28795,N_23138,N_23476);
xor U28796 (N_28796,N_23129,N_22819);
and U28797 (N_28797,N_21089,N_24318);
and U28798 (N_28798,N_20636,N_23400);
nor U28799 (N_28799,N_20101,N_20431);
xnor U28800 (N_28800,N_24141,N_22404);
or U28801 (N_28801,N_20052,N_20260);
or U28802 (N_28802,N_22852,N_23245);
nand U28803 (N_28803,N_21084,N_20874);
nand U28804 (N_28804,N_23511,N_23703);
and U28805 (N_28805,N_21876,N_24395);
nand U28806 (N_28806,N_20898,N_24252);
or U28807 (N_28807,N_24850,N_22410);
nand U28808 (N_28808,N_22623,N_20037);
nor U28809 (N_28809,N_21305,N_20842);
and U28810 (N_28810,N_21070,N_20568);
nor U28811 (N_28811,N_22150,N_20408);
xor U28812 (N_28812,N_24406,N_24079);
nor U28813 (N_28813,N_21937,N_21586);
nand U28814 (N_28814,N_23641,N_20038);
nand U28815 (N_28815,N_20862,N_20009);
nor U28816 (N_28816,N_24940,N_24727);
xor U28817 (N_28817,N_23980,N_24183);
nor U28818 (N_28818,N_22972,N_24684);
xnor U28819 (N_28819,N_23406,N_22983);
nor U28820 (N_28820,N_20007,N_21600);
nor U28821 (N_28821,N_22242,N_24025);
nor U28822 (N_28822,N_23963,N_23176);
and U28823 (N_28823,N_22495,N_20178);
or U28824 (N_28824,N_22692,N_20734);
or U28825 (N_28825,N_21975,N_23161);
nand U28826 (N_28826,N_23583,N_22978);
nor U28827 (N_28827,N_22794,N_23792);
or U28828 (N_28828,N_24390,N_24290);
nand U28829 (N_28829,N_23185,N_23141);
xnor U28830 (N_28830,N_21856,N_21601);
xnor U28831 (N_28831,N_24803,N_23005);
xor U28832 (N_28832,N_20826,N_22060);
nand U28833 (N_28833,N_22751,N_22775);
nand U28834 (N_28834,N_20042,N_21705);
nor U28835 (N_28835,N_24395,N_22638);
nand U28836 (N_28836,N_20392,N_20693);
or U28837 (N_28837,N_21763,N_22320);
nor U28838 (N_28838,N_21161,N_24329);
nor U28839 (N_28839,N_21307,N_21884);
nand U28840 (N_28840,N_20144,N_22734);
nor U28841 (N_28841,N_23305,N_21731);
xnor U28842 (N_28842,N_21982,N_22293);
nand U28843 (N_28843,N_22721,N_21163);
and U28844 (N_28844,N_20354,N_24623);
and U28845 (N_28845,N_21521,N_24485);
nand U28846 (N_28846,N_22230,N_23975);
nand U28847 (N_28847,N_22969,N_24912);
xor U28848 (N_28848,N_22129,N_20727);
and U28849 (N_28849,N_20187,N_22018);
xnor U28850 (N_28850,N_22887,N_21423);
and U28851 (N_28851,N_20524,N_24300);
nor U28852 (N_28852,N_21790,N_23493);
xor U28853 (N_28853,N_24224,N_20019);
nand U28854 (N_28854,N_20971,N_21389);
nand U28855 (N_28855,N_21989,N_24773);
nor U28856 (N_28856,N_22672,N_24867);
nor U28857 (N_28857,N_21797,N_22446);
xor U28858 (N_28858,N_23360,N_22343);
and U28859 (N_28859,N_20653,N_24291);
or U28860 (N_28860,N_22025,N_24412);
nand U28861 (N_28861,N_21433,N_23478);
nand U28862 (N_28862,N_24300,N_22628);
and U28863 (N_28863,N_22250,N_20339);
xor U28864 (N_28864,N_24873,N_20400);
and U28865 (N_28865,N_22628,N_20532);
nand U28866 (N_28866,N_20593,N_24629);
or U28867 (N_28867,N_20194,N_24480);
and U28868 (N_28868,N_20882,N_23337);
nor U28869 (N_28869,N_23307,N_23970);
xor U28870 (N_28870,N_22892,N_22367);
or U28871 (N_28871,N_22172,N_21353);
and U28872 (N_28872,N_24157,N_20062);
nor U28873 (N_28873,N_20204,N_23465);
nand U28874 (N_28874,N_22832,N_20036);
or U28875 (N_28875,N_20193,N_20416);
xor U28876 (N_28876,N_21707,N_20696);
or U28877 (N_28877,N_21407,N_20166);
or U28878 (N_28878,N_23621,N_20616);
or U28879 (N_28879,N_24825,N_21522);
xor U28880 (N_28880,N_20086,N_23179);
xnor U28881 (N_28881,N_20721,N_22237);
xnor U28882 (N_28882,N_23036,N_24110);
nor U28883 (N_28883,N_23749,N_23115);
nor U28884 (N_28884,N_21256,N_22204);
nor U28885 (N_28885,N_21928,N_20681);
xnor U28886 (N_28886,N_24865,N_22506);
and U28887 (N_28887,N_24662,N_23922);
nand U28888 (N_28888,N_24854,N_24171);
nand U28889 (N_28889,N_20356,N_24599);
nand U28890 (N_28890,N_22085,N_21907);
nand U28891 (N_28891,N_21922,N_20301);
or U28892 (N_28892,N_23420,N_23925);
or U28893 (N_28893,N_23743,N_22872);
nor U28894 (N_28894,N_24142,N_21392);
nor U28895 (N_28895,N_20531,N_22237);
xor U28896 (N_28896,N_24489,N_21832);
nand U28897 (N_28897,N_24174,N_20948);
xnor U28898 (N_28898,N_22726,N_23697);
and U28899 (N_28899,N_21638,N_22557);
and U28900 (N_28900,N_23832,N_24477);
nor U28901 (N_28901,N_21478,N_23706);
or U28902 (N_28902,N_23037,N_24108);
nand U28903 (N_28903,N_24117,N_22330);
xor U28904 (N_28904,N_24050,N_24797);
nor U28905 (N_28905,N_23181,N_22230);
and U28906 (N_28906,N_24781,N_22454);
or U28907 (N_28907,N_21732,N_22972);
and U28908 (N_28908,N_24630,N_21154);
nand U28909 (N_28909,N_21406,N_21817);
xnor U28910 (N_28910,N_23896,N_23149);
and U28911 (N_28911,N_22860,N_23628);
nor U28912 (N_28912,N_21974,N_21712);
and U28913 (N_28913,N_24161,N_20571);
nand U28914 (N_28914,N_21862,N_21493);
or U28915 (N_28915,N_21964,N_21992);
nor U28916 (N_28916,N_22646,N_21866);
xor U28917 (N_28917,N_23420,N_21253);
nand U28918 (N_28918,N_23917,N_20658);
nor U28919 (N_28919,N_21880,N_20483);
and U28920 (N_28920,N_22727,N_21237);
xor U28921 (N_28921,N_24574,N_20787);
or U28922 (N_28922,N_22268,N_20305);
or U28923 (N_28923,N_24823,N_20291);
nor U28924 (N_28924,N_24653,N_23428);
xor U28925 (N_28925,N_20272,N_22908);
nand U28926 (N_28926,N_24672,N_23217);
nor U28927 (N_28927,N_21636,N_21294);
or U28928 (N_28928,N_21065,N_20931);
nand U28929 (N_28929,N_24270,N_22139);
and U28930 (N_28930,N_20046,N_24994);
xor U28931 (N_28931,N_20644,N_24095);
or U28932 (N_28932,N_22581,N_20173);
xnor U28933 (N_28933,N_20830,N_20229);
or U28934 (N_28934,N_23746,N_23270);
nand U28935 (N_28935,N_21205,N_24589);
or U28936 (N_28936,N_24496,N_23006);
xnor U28937 (N_28937,N_20764,N_21033);
or U28938 (N_28938,N_22754,N_20973);
and U28939 (N_28939,N_24275,N_20239);
xnor U28940 (N_28940,N_21579,N_22700);
nand U28941 (N_28941,N_21793,N_20363);
nor U28942 (N_28942,N_20855,N_20043);
and U28943 (N_28943,N_21991,N_22868);
nor U28944 (N_28944,N_20091,N_20847);
or U28945 (N_28945,N_22446,N_23613);
or U28946 (N_28946,N_20540,N_23686);
and U28947 (N_28947,N_20786,N_21390);
nand U28948 (N_28948,N_20692,N_22101);
xnor U28949 (N_28949,N_20029,N_20546);
nand U28950 (N_28950,N_24677,N_24232);
or U28951 (N_28951,N_20285,N_20287);
xor U28952 (N_28952,N_21626,N_23799);
nand U28953 (N_28953,N_20224,N_20431);
xnor U28954 (N_28954,N_23213,N_21955);
or U28955 (N_28955,N_23160,N_24371);
xnor U28956 (N_28956,N_24526,N_20111);
or U28957 (N_28957,N_24693,N_23716);
or U28958 (N_28958,N_20914,N_20178);
or U28959 (N_28959,N_24310,N_20501);
or U28960 (N_28960,N_24904,N_22371);
nor U28961 (N_28961,N_22991,N_24877);
and U28962 (N_28962,N_20679,N_21121);
or U28963 (N_28963,N_20223,N_24043);
or U28964 (N_28964,N_21758,N_22037);
nor U28965 (N_28965,N_21029,N_24601);
nand U28966 (N_28966,N_21166,N_21420);
nor U28967 (N_28967,N_24187,N_22434);
xnor U28968 (N_28968,N_23260,N_21374);
and U28969 (N_28969,N_20656,N_23336);
or U28970 (N_28970,N_21902,N_20941);
nand U28971 (N_28971,N_21248,N_22575);
xnor U28972 (N_28972,N_23541,N_22911);
nand U28973 (N_28973,N_20944,N_22839);
nand U28974 (N_28974,N_24544,N_24448);
and U28975 (N_28975,N_24357,N_20214);
nand U28976 (N_28976,N_24736,N_22110);
nor U28977 (N_28977,N_23730,N_24495);
and U28978 (N_28978,N_24478,N_21572);
or U28979 (N_28979,N_21970,N_23733);
and U28980 (N_28980,N_22598,N_21509);
or U28981 (N_28981,N_21235,N_21207);
nand U28982 (N_28982,N_23896,N_24934);
and U28983 (N_28983,N_23384,N_24880);
and U28984 (N_28984,N_22053,N_20627);
and U28985 (N_28985,N_21353,N_20834);
xor U28986 (N_28986,N_23687,N_20689);
nor U28987 (N_28987,N_24550,N_24772);
or U28988 (N_28988,N_23498,N_21251);
and U28989 (N_28989,N_21603,N_21251);
nand U28990 (N_28990,N_21968,N_23116);
nor U28991 (N_28991,N_20722,N_20571);
nand U28992 (N_28992,N_20739,N_20249);
and U28993 (N_28993,N_21895,N_21805);
nand U28994 (N_28994,N_20175,N_21763);
and U28995 (N_28995,N_22782,N_24467);
xnor U28996 (N_28996,N_22519,N_24589);
and U28997 (N_28997,N_22589,N_21465);
xnor U28998 (N_28998,N_24031,N_22103);
nor U28999 (N_28999,N_21107,N_23727);
and U29000 (N_29000,N_24331,N_20769);
or U29001 (N_29001,N_20380,N_24783);
nor U29002 (N_29002,N_21932,N_24744);
nor U29003 (N_29003,N_21305,N_24436);
and U29004 (N_29004,N_20526,N_21882);
and U29005 (N_29005,N_23520,N_23644);
nor U29006 (N_29006,N_22102,N_20655);
nand U29007 (N_29007,N_21146,N_22292);
nand U29008 (N_29008,N_21520,N_20946);
nor U29009 (N_29009,N_22817,N_22823);
xnor U29010 (N_29010,N_21661,N_21525);
xnor U29011 (N_29011,N_24292,N_20482);
and U29012 (N_29012,N_21465,N_23136);
xnor U29013 (N_29013,N_21051,N_24295);
nor U29014 (N_29014,N_22444,N_23588);
nor U29015 (N_29015,N_22585,N_21311);
or U29016 (N_29016,N_22263,N_22179);
and U29017 (N_29017,N_23362,N_20506);
nor U29018 (N_29018,N_20865,N_21116);
xnor U29019 (N_29019,N_24002,N_20522);
or U29020 (N_29020,N_24890,N_24173);
nand U29021 (N_29021,N_21836,N_22768);
or U29022 (N_29022,N_21402,N_20697);
xor U29023 (N_29023,N_22567,N_23385);
or U29024 (N_29024,N_22413,N_22156);
nand U29025 (N_29025,N_24098,N_23294);
nor U29026 (N_29026,N_22552,N_22114);
or U29027 (N_29027,N_22799,N_23547);
xnor U29028 (N_29028,N_20344,N_22503);
xnor U29029 (N_29029,N_24760,N_23273);
xor U29030 (N_29030,N_21451,N_24166);
nor U29031 (N_29031,N_23059,N_22041);
or U29032 (N_29032,N_22620,N_21144);
and U29033 (N_29033,N_21872,N_20742);
nand U29034 (N_29034,N_21343,N_22964);
and U29035 (N_29035,N_24279,N_20533);
and U29036 (N_29036,N_21382,N_20085);
and U29037 (N_29037,N_22780,N_22289);
nand U29038 (N_29038,N_23537,N_22780);
xor U29039 (N_29039,N_23891,N_21093);
or U29040 (N_29040,N_20485,N_20438);
or U29041 (N_29041,N_20753,N_24885);
nor U29042 (N_29042,N_23851,N_23942);
xor U29043 (N_29043,N_24915,N_24355);
xor U29044 (N_29044,N_21894,N_20098);
nand U29045 (N_29045,N_21040,N_24164);
or U29046 (N_29046,N_20262,N_22815);
and U29047 (N_29047,N_24101,N_23886);
or U29048 (N_29048,N_20255,N_21054);
or U29049 (N_29049,N_21447,N_20062);
or U29050 (N_29050,N_22344,N_20075);
xnor U29051 (N_29051,N_22140,N_23933);
nor U29052 (N_29052,N_21972,N_23701);
or U29053 (N_29053,N_24399,N_23746);
xnor U29054 (N_29054,N_24947,N_21869);
and U29055 (N_29055,N_21749,N_23462);
or U29056 (N_29056,N_24797,N_21504);
nand U29057 (N_29057,N_21682,N_24356);
nor U29058 (N_29058,N_21011,N_24732);
xor U29059 (N_29059,N_21692,N_22915);
and U29060 (N_29060,N_20003,N_21190);
or U29061 (N_29061,N_21831,N_23610);
xnor U29062 (N_29062,N_23154,N_22905);
nand U29063 (N_29063,N_23438,N_20754);
xor U29064 (N_29064,N_24489,N_23151);
nor U29065 (N_29065,N_24646,N_21956);
and U29066 (N_29066,N_22737,N_20848);
or U29067 (N_29067,N_23450,N_22371);
nand U29068 (N_29068,N_22347,N_21447);
or U29069 (N_29069,N_22039,N_23568);
and U29070 (N_29070,N_24065,N_20093);
nand U29071 (N_29071,N_21265,N_22376);
nand U29072 (N_29072,N_20626,N_22742);
nor U29073 (N_29073,N_23261,N_24598);
and U29074 (N_29074,N_21725,N_24048);
xnor U29075 (N_29075,N_21851,N_20380);
or U29076 (N_29076,N_23964,N_20707);
or U29077 (N_29077,N_21512,N_24913);
or U29078 (N_29078,N_21388,N_22403);
nor U29079 (N_29079,N_20233,N_20318);
xnor U29080 (N_29080,N_24664,N_24636);
or U29081 (N_29081,N_24349,N_21885);
and U29082 (N_29082,N_21342,N_22406);
and U29083 (N_29083,N_20656,N_23256);
or U29084 (N_29084,N_23551,N_22623);
xnor U29085 (N_29085,N_24279,N_20034);
xor U29086 (N_29086,N_24680,N_21356);
nand U29087 (N_29087,N_23737,N_23500);
nor U29088 (N_29088,N_24366,N_21644);
and U29089 (N_29089,N_23780,N_21515);
xor U29090 (N_29090,N_21701,N_22214);
and U29091 (N_29091,N_23028,N_23063);
and U29092 (N_29092,N_21298,N_21533);
nand U29093 (N_29093,N_22639,N_22855);
and U29094 (N_29094,N_24281,N_23857);
or U29095 (N_29095,N_24946,N_22862);
and U29096 (N_29096,N_23728,N_22672);
or U29097 (N_29097,N_21197,N_23176);
and U29098 (N_29098,N_22220,N_23768);
nand U29099 (N_29099,N_20727,N_22637);
or U29100 (N_29100,N_20351,N_20897);
xnor U29101 (N_29101,N_22561,N_22320);
xor U29102 (N_29102,N_22397,N_22811);
xnor U29103 (N_29103,N_24051,N_21783);
xor U29104 (N_29104,N_23008,N_24705);
and U29105 (N_29105,N_23760,N_21851);
nor U29106 (N_29106,N_21052,N_23762);
xor U29107 (N_29107,N_20948,N_23187);
or U29108 (N_29108,N_24044,N_24840);
or U29109 (N_29109,N_21939,N_24824);
nand U29110 (N_29110,N_21228,N_23262);
or U29111 (N_29111,N_22388,N_23975);
nand U29112 (N_29112,N_21148,N_21842);
nand U29113 (N_29113,N_24909,N_23847);
nand U29114 (N_29114,N_20196,N_24426);
and U29115 (N_29115,N_24598,N_24010);
nor U29116 (N_29116,N_24452,N_21832);
or U29117 (N_29117,N_24638,N_24747);
nand U29118 (N_29118,N_20696,N_24368);
nor U29119 (N_29119,N_20886,N_24651);
nand U29120 (N_29120,N_24393,N_24086);
or U29121 (N_29121,N_24240,N_21757);
nor U29122 (N_29122,N_20031,N_20620);
xor U29123 (N_29123,N_23193,N_21234);
and U29124 (N_29124,N_21226,N_23843);
and U29125 (N_29125,N_23940,N_20812);
nand U29126 (N_29126,N_24309,N_24492);
and U29127 (N_29127,N_24389,N_22198);
nor U29128 (N_29128,N_21037,N_24284);
or U29129 (N_29129,N_21260,N_23189);
or U29130 (N_29130,N_23507,N_23615);
xor U29131 (N_29131,N_23590,N_22103);
nand U29132 (N_29132,N_22906,N_20337);
and U29133 (N_29133,N_22052,N_21448);
and U29134 (N_29134,N_23510,N_20524);
xor U29135 (N_29135,N_24291,N_23124);
xor U29136 (N_29136,N_21944,N_21165);
nand U29137 (N_29137,N_22340,N_24350);
xor U29138 (N_29138,N_22604,N_24405);
or U29139 (N_29139,N_20943,N_24286);
and U29140 (N_29140,N_23593,N_21853);
nand U29141 (N_29141,N_22906,N_22036);
nand U29142 (N_29142,N_20380,N_23823);
nor U29143 (N_29143,N_20615,N_24967);
xor U29144 (N_29144,N_24850,N_21126);
and U29145 (N_29145,N_20188,N_20930);
xnor U29146 (N_29146,N_24443,N_21782);
nand U29147 (N_29147,N_23364,N_21855);
xnor U29148 (N_29148,N_20006,N_22851);
or U29149 (N_29149,N_22986,N_23205);
or U29150 (N_29150,N_20519,N_21582);
or U29151 (N_29151,N_21336,N_20422);
or U29152 (N_29152,N_24375,N_22326);
xnor U29153 (N_29153,N_22095,N_23219);
xnor U29154 (N_29154,N_24532,N_23609);
nand U29155 (N_29155,N_22847,N_21071);
or U29156 (N_29156,N_22385,N_22992);
xnor U29157 (N_29157,N_21967,N_24268);
nand U29158 (N_29158,N_22304,N_21395);
and U29159 (N_29159,N_20157,N_22573);
nor U29160 (N_29160,N_24221,N_24664);
and U29161 (N_29161,N_20437,N_22159);
xnor U29162 (N_29162,N_24475,N_24237);
xnor U29163 (N_29163,N_22671,N_22631);
xnor U29164 (N_29164,N_21765,N_22022);
nor U29165 (N_29165,N_22448,N_22167);
or U29166 (N_29166,N_20879,N_24832);
nor U29167 (N_29167,N_24881,N_23953);
or U29168 (N_29168,N_21755,N_24793);
and U29169 (N_29169,N_23336,N_21877);
nor U29170 (N_29170,N_22967,N_22270);
or U29171 (N_29171,N_22395,N_20667);
nand U29172 (N_29172,N_20547,N_23605);
nand U29173 (N_29173,N_24844,N_23186);
nor U29174 (N_29174,N_20415,N_23557);
or U29175 (N_29175,N_20780,N_22638);
xnor U29176 (N_29176,N_20948,N_21183);
xnor U29177 (N_29177,N_20936,N_24078);
xor U29178 (N_29178,N_21141,N_20328);
and U29179 (N_29179,N_23342,N_23021);
or U29180 (N_29180,N_22716,N_23093);
nand U29181 (N_29181,N_20698,N_21160);
nor U29182 (N_29182,N_24879,N_21995);
or U29183 (N_29183,N_20726,N_20083);
and U29184 (N_29184,N_20511,N_23972);
nand U29185 (N_29185,N_20102,N_22018);
xor U29186 (N_29186,N_20200,N_22901);
xor U29187 (N_29187,N_22263,N_20255);
xnor U29188 (N_29188,N_23155,N_24360);
xor U29189 (N_29189,N_20193,N_20310);
nand U29190 (N_29190,N_20222,N_21793);
or U29191 (N_29191,N_24388,N_20491);
and U29192 (N_29192,N_22311,N_23795);
xnor U29193 (N_29193,N_22940,N_20693);
nor U29194 (N_29194,N_21751,N_21000);
and U29195 (N_29195,N_22413,N_21516);
xnor U29196 (N_29196,N_20567,N_20359);
nor U29197 (N_29197,N_23887,N_23307);
nor U29198 (N_29198,N_22211,N_21612);
nand U29199 (N_29199,N_23378,N_23065);
nor U29200 (N_29200,N_22531,N_24427);
and U29201 (N_29201,N_24478,N_23688);
nand U29202 (N_29202,N_21730,N_22919);
nand U29203 (N_29203,N_23908,N_20727);
nand U29204 (N_29204,N_21432,N_22911);
nor U29205 (N_29205,N_24315,N_20520);
xor U29206 (N_29206,N_20774,N_21823);
xnor U29207 (N_29207,N_22548,N_24159);
or U29208 (N_29208,N_24558,N_20266);
nand U29209 (N_29209,N_24139,N_22124);
nor U29210 (N_29210,N_20555,N_21555);
xor U29211 (N_29211,N_24420,N_22405);
or U29212 (N_29212,N_23790,N_20777);
nand U29213 (N_29213,N_23543,N_23605);
and U29214 (N_29214,N_24606,N_22227);
nor U29215 (N_29215,N_24555,N_23704);
nor U29216 (N_29216,N_23155,N_21470);
and U29217 (N_29217,N_22706,N_20432);
xor U29218 (N_29218,N_22184,N_22128);
nand U29219 (N_29219,N_20537,N_23423);
xnor U29220 (N_29220,N_20781,N_20006);
xor U29221 (N_29221,N_21588,N_20682);
and U29222 (N_29222,N_21678,N_21119);
xnor U29223 (N_29223,N_22862,N_23302);
nand U29224 (N_29224,N_22473,N_22193);
nor U29225 (N_29225,N_23536,N_20899);
xor U29226 (N_29226,N_24165,N_21619);
and U29227 (N_29227,N_22645,N_20621);
xnor U29228 (N_29228,N_20442,N_21789);
xor U29229 (N_29229,N_20853,N_22189);
or U29230 (N_29230,N_24334,N_24037);
nand U29231 (N_29231,N_20392,N_22769);
or U29232 (N_29232,N_22263,N_22162);
or U29233 (N_29233,N_24080,N_22234);
nor U29234 (N_29234,N_22507,N_23109);
and U29235 (N_29235,N_23495,N_22402);
nor U29236 (N_29236,N_20129,N_23911);
nand U29237 (N_29237,N_23740,N_24689);
xnor U29238 (N_29238,N_22592,N_20874);
and U29239 (N_29239,N_23472,N_24947);
and U29240 (N_29240,N_23396,N_20417);
and U29241 (N_29241,N_24755,N_23528);
nor U29242 (N_29242,N_24338,N_23475);
and U29243 (N_29243,N_24867,N_20600);
nand U29244 (N_29244,N_22849,N_20826);
and U29245 (N_29245,N_23908,N_24884);
nand U29246 (N_29246,N_21694,N_22651);
xnor U29247 (N_29247,N_22544,N_20989);
and U29248 (N_29248,N_24444,N_23771);
nor U29249 (N_29249,N_23018,N_24160);
nand U29250 (N_29250,N_22776,N_23598);
nand U29251 (N_29251,N_22296,N_23018);
nor U29252 (N_29252,N_22390,N_23943);
and U29253 (N_29253,N_20902,N_20467);
nand U29254 (N_29254,N_21787,N_21925);
and U29255 (N_29255,N_22635,N_24688);
nand U29256 (N_29256,N_22717,N_23156);
nand U29257 (N_29257,N_22003,N_24790);
and U29258 (N_29258,N_21362,N_21441);
or U29259 (N_29259,N_22232,N_24516);
nand U29260 (N_29260,N_22594,N_23385);
nand U29261 (N_29261,N_22089,N_23912);
and U29262 (N_29262,N_24729,N_21795);
nor U29263 (N_29263,N_23142,N_21134);
nand U29264 (N_29264,N_21153,N_21074);
xnor U29265 (N_29265,N_24007,N_20355);
xor U29266 (N_29266,N_21572,N_22094);
xnor U29267 (N_29267,N_24988,N_23669);
nand U29268 (N_29268,N_20759,N_20949);
nor U29269 (N_29269,N_22115,N_20562);
nor U29270 (N_29270,N_20804,N_21750);
and U29271 (N_29271,N_20772,N_20765);
nand U29272 (N_29272,N_21500,N_21555);
or U29273 (N_29273,N_23000,N_21212);
or U29274 (N_29274,N_22627,N_23055);
or U29275 (N_29275,N_22261,N_24267);
nor U29276 (N_29276,N_22412,N_24841);
or U29277 (N_29277,N_20710,N_24276);
or U29278 (N_29278,N_24731,N_21576);
nand U29279 (N_29279,N_24241,N_23604);
xnor U29280 (N_29280,N_24578,N_24503);
and U29281 (N_29281,N_23198,N_23358);
or U29282 (N_29282,N_20971,N_20679);
nor U29283 (N_29283,N_20669,N_23281);
or U29284 (N_29284,N_22022,N_21225);
or U29285 (N_29285,N_21986,N_23424);
nand U29286 (N_29286,N_23166,N_21283);
nor U29287 (N_29287,N_22242,N_23113);
and U29288 (N_29288,N_23101,N_22568);
nand U29289 (N_29289,N_22817,N_23093);
and U29290 (N_29290,N_24342,N_20453);
or U29291 (N_29291,N_21407,N_21817);
nand U29292 (N_29292,N_21815,N_20700);
or U29293 (N_29293,N_23334,N_22113);
nand U29294 (N_29294,N_20769,N_22993);
xnor U29295 (N_29295,N_20028,N_23339);
and U29296 (N_29296,N_20628,N_22981);
xnor U29297 (N_29297,N_23763,N_21652);
nand U29298 (N_29298,N_22110,N_20808);
nor U29299 (N_29299,N_22718,N_20499);
xor U29300 (N_29300,N_22267,N_21717);
nand U29301 (N_29301,N_21832,N_22863);
or U29302 (N_29302,N_23315,N_20583);
xnor U29303 (N_29303,N_20617,N_22651);
or U29304 (N_29304,N_22428,N_22009);
nor U29305 (N_29305,N_21378,N_24661);
or U29306 (N_29306,N_23263,N_21723);
xor U29307 (N_29307,N_20150,N_22018);
nor U29308 (N_29308,N_21961,N_20165);
xnor U29309 (N_29309,N_22023,N_23531);
xnor U29310 (N_29310,N_24750,N_23631);
nor U29311 (N_29311,N_24084,N_23861);
nand U29312 (N_29312,N_22099,N_21149);
xnor U29313 (N_29313,N_22793,N_21403);
or U29314 (N_29314,N_24454,N_24648);
xnor U29315 (N_29315,N_23593,N_24042);
nor U29316 (N_29316,N_20977,N_20645);
and U29317 (N_29317,N_20686,N_24706);
and U29318 (N_29318,N_20305,N_23975);
xnor U29319 (N_29319,N_20010,N_23465);
nand U29320 (N_29320,N_20190,N_23606);
xnor U29321 (N_29321,N_21406,N_23007);
and U29322 (N_29322,N_24091,N_24750);
or U29323 (N_29323,N_24002,N_20528);
and U29324 (N_29324,N_23485,N_23577);
or U29325 (N_29325,N_20651,N_23391);
xor U29326 (N_29326,N_23207,N_24156);
nor U29327 (N_29327,N_20436,N_23015);
or U29328 (N_29328,N_21092,N_21977);
or U29329 (N_29329,N_23133,N_24382);
xor U29330 (N_29330,N_22247,N_21258);
xor U29331 (N_29331,N_22494,N_22241);
or U29332 (N_29332,N_20873,N_22813);
xor U29333 (N_29333,N_22064,N_23158);
nor U29334 (N_29334,N_21370,N_20765);
or U29335 (N_29335,N_20950,N_23064);
nor U29336 (N_29336,N_23664,N_20623);
xnor U29337 (N_29337,N_23034,N_23136);
or U29338 (N_29338,N_20359,N_21806);
nand U29339 (N_29339,N_20255,N_22137);
nand U29340 (N_29340,N_20888,N_22994);
xor U29341 (N_29341,N_24887,N_24805);
or U29342 (N_29342,N_24744,N_20063);
nand U29343 (N_29343,N_21757,N_24016);
nand U29344 (N_29344,N_22698,N_24128);
or U29345 (N_29345,N_22415,N_20628);
and U29346 (N_29346,N_21365,N_24083);
or U29347 (N_29347,N_22789,N_24555);
or U29348 (N_29348,N_21920,N_24088);
or U29349 (N_29349,N_22396,N_23345);
and U29350 (N_29350,N_23096,N_21789);
nand U29351 (N_29351,N_20961,N_23101);
or U29352 (N_29352,N_24106,N_21797);
or U29353 (N_29353,N_24086,N_23139);
or U29354 (N_29354,N_20472,N_21297);
xor U29355 (N_29355,N_20377,N_24003);
and U29356 (N_29356,N_20712,N_24217);
or U29357 (N_29357,N_20741,N_24087);
xnor U29358 (N_29358,N_20793,N_20839);
or U29359 (N_29359,N_24834,N_24833);
nand U29360 (N_29360,N_20597,N_20912);
and U29361 (N_29361,N_20910,N_22752);
nand U29362 (N_29362,N_23947,N_24547);
nor U29363 (N_29363,N_24742,N_23502);
nor U29364 (N_29364,N_23988,N_21924);
nor U29365 (N_29365,N_23001,N_24143);
or U29366 (N_29366,N_24290,N_21088);
nand U29367 (N_29367,N_21676,N_22597);
nand U29368 (N_29368,N_23522,N_23307);
xor U29369 (N_29369,N_20798,N_24880);
nor U29370 (N_29370,N_24954,N_24619);
and U29371 (N_29371,N_24054,N_21002);
or U29372 (N_29372,N_20646,N_23220);
or U29373 (N_29373,N_21570,N_22654);
or U29374 (N_29374,N_22818,N_22555);
nor U29375 (N_29375,N_21865,N_20970);
or U29376 (N_29376,N_24399,N_20752);
xor U29377 (N_29377,N_23916,N_20108);
nand U29378 (N_29378,N_23419,N_22411);
or U29379 (N_29379,N_21766,N_24521);
nand U29380 (N_29380,N_24023,N_24708);
nor U29381 (N_29381,N_24857,N_20356);
xnor U29382 (N_29382,N_24004,N_24842);
nand U29383 (N_29383,N_24358,N_22621);
nand U29384 (N_29384,N_21362,N_20536);
nand U29385 (N_29385,N_22295,N_23565);
xnor U29386 (N_29386,N_24121,N_23139);
nor U29387 (N_29387,N_20267,N_23957);
nor U29388 (N_29388,N_23618,N_24636);
and U29389 (N_29389,N_22936,N_20883);
or U29390 (N_29390,N_23413,N_23874);
nor U29391 (N_29391,N_21304,N_23660);
nand U29392 (N_29392,N_24117,N_23165);
nor U29393 (N_29393,N_22454,N_20306);
and U29394 (N_29394,N_23895,N_22533);
and U29395 (N_29395,N_23743,N_24005);
nand U29396 (N_29396,N_20610,N_24524);
and U29397 (N_29397,N_21411,N_21054);
and U29398 (N_29398,N_23688,N_21607);
nor U29399 (N_29399,N_20106,N_23008);
xnor U29400 (N_29400,N_20482,N_23589);
nand U29401 (N_29401,N_21661,N_24095);
xnor U29402 (N_29402,N_22229,N_21230);
nand U29403 (N_29403,N_23556,N_20317);
or U29404 (N_29404,N_21581,N_24514);
and U29405 (N_29405,N_21111,N_20637);
nor U29406 (N_29406,N_22355,N_21195);
nand U29407 (N_29407,N_21963,N_23967);
nand U29408 (N_29408,N_22427,N_24134);
or U29409 (N_29409,N_23463,N_23269);
nor U29410 (N_29410,N_22330,N_22952);
nor U29411 (N_29411,N_21071,N_21099);
and U29412 (N_29412,N_23491,N_22325);
or U29413 (N_29413,N_22592,N_21830);
nand U29414 (N_29414,N_24436,N_22646);
or U29415 (N_29415,N_23017,N_20724);
xnor U29416 (N_29416,N_23566,N_20441);
nand U29417 (N_29417,N_24775,N_23948);
xor U29418 (N_29418,N_23477,N_21632);
nor U29419 (N_29419,N_24067,N_24518);
or U29420 (N_29420,N_20099,N_24674);
and U29421 (N_29421,N_21626,N_24510);
and U29422 (N_29422,N_22828,N_21682);
xor U29423 (N_29423,N_20667,N_22906);
xnor U29424 (N_29424,N_22473,N_22610);
nor U29425 (N_29425,N_21626,N_22668);
nand U29426 (N_29426,N_21689,N_24339);
nor U29427 (N_29427,N_20543,N_23772);
or U29428 (N_29428,N_22628,N_21225);
nor U29429 (N_29429,N_21010,N_20646);
and U29430 (N_29430,N_20334,N_20252);
or U29431 (N_29431,N_21399,N_23570);
nand U29432 (N_29432,N_20688,N_22327);
xor U29433 (N_29433,N_23316,N_22826);
nand U29434 (N_29434,N_24641,N_20359);
nand U29435 (N_29435,N_20577,N_22288);
or U29436 (N_29436,N_21696,N_21405);
or U29437 (N_29437,N_23598,N_24929);
xnor U29438 (N_29438,N_21337,N_24024);
nor U29439 (N_29439,N_22280,N_20757);
xnor U29440 (N_29440,N_24081,N_22178);
or U29441 (N_29441,N_23582,N_21160);
nor U29442 (N_29442,N_21739,N_23367);
or U29443 (N_29443,N_20654,N_21246);
xor U29444 (N_29444,N_24182,N_21240);
nor U29445 (N_29445,N_23854,N_20232);
and U29446 (N_29446,N_24765,N_21630);
nor U29447 (N_29447,N_21022,N_20040);
or U29448 (N_29448,N_21844,N_23120);
nor U29449 (N_29449,N_20573,N_22348);
and U29450 (N_29450,N_23542,N_21614);
and U29451 (N_29451,N_22984,N_21967);
and U29452 (N_29452,N_21043,N_22624);
nand U29453 (N_29453,N_24772,N_21666);
nor U29454 (N_29454,N_22650,N_20047);
nand U29455 (N_29455,N_22153,N_20163);
or U29456 (N_29456,N_23925,N_20100);
or U29457 (N_29457,N_20962,N_20019);
xor U29458 (N_29458,N_20678,N_22554);
nor U29459 (N_29459,N_22932,N_23808);
and U29460 (N_29460,N_24921,N_22103);
nor U29461 (N_29461,N_23121,N_22663);
nor U29462 (N_29462,N_24726,N_23839);
nor U29463 (N_29463,N_20220,N_23809);
or U29464 (N_29464,N_21308,N_22745);
xor U29465 (N_29465,N_24667,N_24369);
nor U29466 (N_29466,N_20199,N_24915);
xnor U29467 (N_29467,N_23092,N_22094);
nor U29468 (N_29468,N_23060,N_21616);
and U29469 (N_29469,N_21830,N_20876);
xor U29470 (N_29470,N_24224,N_21693);
xor U29471 (N_29471,N_23799,N_20873);
nor U29472 (N_29472,N_23333,N_23737);
nor U29473 (N_29473,N_20505,N_23820);
nand U29474 (N_29474,N_24002,N_21064);
xor U29475 (N_29475,N_22132,N_23128);
nand U29476 (N_29476,N_23161,N_21834);
and U29477 (N_29477,N_23138,N_23706);
xor U29478 (N_29478,N_20741,N_20479);
nand U29479 (N_29479,N_24201,N_22698);
nand U29480 (N_29480,N_21453,N_24507);
or U29481 (N_29481,N_21778,N_20167);
nand U29482 (N_29482,N_24563,N_21157);
nor U29483 (N_29483,N_23039,N_22223);
nor U29484 (N_29484,N_21559,N_20440);
nand U29485 (N_29485,N_23347,N_22315);
nor U29486 (N_29486,N_22718,N_21816);
or U29487 (N_29487,N_20979,N_20101);
nand U29488 (N_29488,N_21931,N_24845);
nand U29489 (N_29489,N_20564,N_20198);
and U29490 (N_29490,N_20410,N_24638);
xor U29491 (N_29491,N_22773,N_23473);
and U29492 (N_29492,N_21242,N_23064);
nor U29493 (N_29493,N_20071,N_23626);
or U29494 (N_29494,N_23835,N_24179);
and U29495 (N_29495,N_23371,N_21470);
and U29496 (N_29496,N_22042,N_21824);
or U29497 (N_29497,N_22187,N_21387);
nor U29498 (N_29498,N_21888,N_20075);
nor U29499 (N_29499,N_23510,N_24725);
and U29500 (N_29500,N_21713,N_24146);
xnor U29501 (N_29501,N_20062,N_20319);
nor U29502 (N_29502,N_24658,N_24006);
or U29503 (N_29503,N_22368,N_22612);
xor U29504 (N_29504,N_20315,N_23821);
and U29505 (N_29505,N_24855,N_23747);
nor U29506 (N_29506,N_22079,N_20041);
or U29507 (N_29507,N_23725,N_20460);
or U29508 (N_29508,N_20748,N_22936);
or U29509 (N_29509,N_23914,N_24597);
nor U29510 (N_29510,N_23489,N_22556);
or U29511 (N_29511,N_21392,N_23547);
and U29512 (N_29512,N_24823,N_20199);
xor U29513 (N_29513,N_22649,N_23694);
nor U29514 (N_29514,N_22956,N_21152);
nand U29515 (N_29515,N_23499,N_22818);
nand U29516 (N_29516,N_20374,N_22640);
nand U29517 (N_29517,N_21559,N_24306);
nor U29518 (N_29518,N_20273,N_22146);
xnor U29519 (N_29519,N_21367,N_24976);
or U29520 (N_29520,N_21940,N_22585);
nor U29521 (N_29521,N_23099,N_23674);
nand U29522 (N_29522,N_20874,N_22660);
nand U29523 (N_29523,N_23049,N_21177);
nand U29524 (N_29524,N_22405,N_22392);
or U29525 (N_29525,N_20881,N_23521);
and U29526 (N_29526,N_22449,N_22277);
and U29527 (N_29527,N_23941,N_23402);
xnor U29528 (N_29528,N_20315,N_24832);
nand U29529 (N_29529,N_22473,N_24897);
or U29530 (N_29530,N_22689,N_21129);
and U29531 (N_29531,N_22191,N_21016);
and U29532 (N_29532,N_22709,N_20536);
or U29533 (N_29533,N_24362,N_22563);
nand U29534 (N_29534,N_21162,N_20499);
nand U29535 (N_29535,N_20282,N_24847);
or U29536 (N_29536,N_22868,N_21302);
and U29537 (N_29537,N_24905,N_20268);
and U29538 (N_29538,N_23543,N_24234);
and U29539 (N_29539,N_20389,N_24909);
or U29540 (N_29540,N_23796,N_23442);
nor U29541 (N_29541,N_22122,N_20266);
nand U29542 (N_29542,N_21171,N_24248);
xnor U29543 (N_29543,N_21645,N_21265);
xnor U29544 (N_29544,N_24835,N_24709);
xnor U29545 (N_29545,N_24733,N_22393);
xnor U29546 (N_29546,N_21141,N_24671);
nor U29547 (N_29547,N_21949,N_22134);
nor U29548 (N_29548,N_23984,N_20011);
and U29549 (N_29549,N_24427,N_22180);
xnor U29550 (N_29550,N_24744,N_20739);
or U29551 (N_29551,N_23844,N_20875);
nand U29552 (N_29552,N_24498,N_20569);
nor U29553 (N_29553,N_20761,N_23578);
xnor U29554 (N_29554,N_24082,N_21945);
or U29555 (N_29555,N_20793,N_20927);
nor U29556 (N_29556,N_24316,N_23106);
nand U29557 (N_29557,N_24210,N_23407);
xor U29558 (N_29558,N_22526,N_22141);
nand U29559 (N_29559,N_21400,N_20957);
and U29560 (N_29560,N_20252,N_21789);
xor U29561 (N_29561,N_20654,N_20645);
xnor U29562 (N_29562,N_23981,N_20575);
nand U29563 (N_29563,N_22044,N_21140);
or U29564 (N_29564,N_21916,N_23227);
xor U29565 (N_29565,N_24815,N_22321);
nand U29566 (N_29566,N_24224,N_22608);
or U29567 (N_29567,N_22249,N_23052);
or U29568 (N_29568,N_20944,N_22283);
nand U29569 (N_29569,N_23403,N_23168);
or U29570 (N_29570,N_21808,N_21005);
nand U29571 (N_29571,N_23761,N_23184);
xnor U29572 (N_29572,N_21022,N_21564);
nor U29573 (N_29573,N_20940,N_24388);
and U29574 (N_29574,N_20041,N_23778);
xor U29575 (N_29575,N_23602,N_21725);
nor U29576 (N_29576,N_22837,N_20974);
nor U29577 (N_29577,N_24722,N_23727);
nor U29578 (N_29578,N_21982,N_21858);
or U29579 (N_29579,N_24749,N_20009);
or U29580 (N_29580,N_23780,N_22015);
nor U29581 (N_29581,N_24952,N_22742);
nor U29582 (N_29582,N_20060,N_23291);
nand U29583 (N_29583,N_24959,N_21004);
nor U29584 (N_29584,N_20719,N_24928);
and U29585 (N_29585,N_24973,N_20363);
nor U29586 (N_29586,N_20285,N_20431);
or U29587 (N_29587,N_20239,N_22511);
nor U29588 (N_29588,N_21667,N_22237);
or U29589 (N_29589,N_24678,N_20660);
xor U29590 (N_29590,N_24496,N_20436);
or U29591 (N_29591,N_23710,N_24700);
xor U29592 (N_29592,N_24497,N_20721);
or U29593 (N_29593,N_21188,N_20506);
nor U29594 (N_29594,N_23905,N_20867);
xor U29595 (N_29595,N_20505,N_20189);
nand U29596 (N_29596,N_20836,N_20015);
xor U29597 (N_29597,N_21857,N_21128);
and U29598 (N_29598,N_21676,N_21683);
nor U29599 (N_29599,N_23960,N_24151);
xor U29600 (N_29600,N_24334,N_22743);
and U29601 (N_29601,N_20576,N_21132);
nand U29602 (N_29602,N_20860,N_20171);
xnor U29603 (N_29603,N_23439,N_22324);
nand U29604 (N_29604,N_24307,N_24536);
and U29605 (N_29605,N_22719,N_20719);
xnor U29606 (N_29606,N_21136,N_20938);
nand U29607 (N_29607,N_22980,N_20590);
xor U29608 (N_29608,N_21765,N_21567);
nand U29609 (N_29609,N_22400,N_22856);
or U29610 (N_29610,N_22515,N_24645);
xor U29611 (N_29611,N_23294,N_21271);
and U29612 (N_29612,N_20292,N_23531);
and U29613 (N_29613,N_23539,N_20359);
or U29614 (N_29614,N_22339,N_21156);
xnor U29615 (N_29615,N_24404,N_20375);
and U29616 (N_29616,N_21053,N_22451);
nand U29617 (N_29617,N_20801,N_22719);
xor U29618 (N_29618,N_21437,N_23486);
nor U29619 (N_29619,N_24356,N_24386);
nand U29620 (N_29620,N_24770,N_21212);
nor U29621 (N_29621,N_20422,N_20952);
and U29622 (N_29622,N_22394,N_23076);
nand U29623 (N_29623,N_23042,N_23610);
nand U29624 (N_29624,N_20786,N_20869);
nand U29625 (N_29625,N_20834,N_20769);
xor U29626 (N_29626,N_21988,N_21322);
nand U29627 (N_29627,N_23846,N_22981);
xor U29628 (N_29628,N_21514,N_23504);
nand U29629 (N_29629,N_23849,N_23161);
nand U29630 (N_29630,N_23994,N_21082);
and U29631 (N_29631,N_24720,N_20189);
nand U29632 (N_29632,N_20457,N_21743);
xor U29633 (N_29633,N_23972,N_20660);
or U29634 (N_29634,N_21881,N_20214);
and U29635 (N_29635,N_22105,N_24758);
or U29636 (N_29636,N_23425,N_22624);
or U29637 (N_29637,N_21599,N_20541);
nor U29638 (N_29638,N_20553,N_24385);
and U29639 (N_29639,N_24425,N_21790);
nor U29640 (N_29640,N_24750,N_24463);
and U29641 (N_29641,N_20595,N_23628);
xor U29642 (N_29642,N_22728,N_20710);
nor U29643 (N_29643,N_22115,N_22533);
xnor U29644 (N_29644,N_23230,N_20579);
nand U29645 (N_29645,N_23369,N_21413);
or U29646 (N_29646,N_21829,N_23487);
nand U29647 (N_29647,N_22454,N_22159);
xnor U29648 (N_29648,N_22736,N_22752);
or U29649 (N_29649,N_24796,N_23466);
xnor U29650 (N_29650,N_21311,N_20463);
xor U29651 (N_29651,N_23124,N_23265);
or U29652 (N_29652,N_22017,N_20791);
and U29653 (N_29653,N_21005,N_21153);
or U29654 (N_29654,N_20632,N_20286);
nor U29655 (N_29655,N_24449,N_20267);
and U29656 (N_29656,N_22478,N_21551);
nor U29657 (N_29657,N_20053,N_24320);
or U29658 (N_29658,N_22906,N_24808);
and U29659 (N_29659,N_23927,N_23431);
or U29660 (N_29660,N_23716,N_24031);
nor U29661 (N_29661,N_23910,N_23142);
and U29662 (N_29662,N_22819,N_23526);
nand U29663 (N_29663,N_24491,N_20541);
or U29664 (N_29664,N_21637,N_24147);
xor U29665 (N_29665,N_21046,N_20590);
xor U29666 (N_29666,N_20131,N_24292);
and U29667 (N_29667,N_24878,N_21905);
nand U29668 (N_29668,N_24029,N_22235);
and U29669 (N_29669,N_22647,N_20047);
and U29670 (N_29670,N_20833,N_24126);
and U29671 (N_29671,N_24472,N_24358);
and U29672 (N_29672,N_21808,N_21603);
or U29673 (N_29673,N_23991,N_22364);
and U29674 (N_29674,N_23978,N_20144);
nor U29675 (N_29675,N_21485,N_24017);
or U29676 (N_29676,N_21499,N_23913);
or U29677 (N_29677,N_21177,N_24783);
or U29678 (N_29678,N_22208,N_24694);
nand U29679 (N_29679,N_23466,N_23342);
or U29680 (N_29680,N_20575,N_24315);
nor U29681 (N_29681,N_24184,N_24042);
xor U29682 (N_29682,N_20360,N_20306);
and U29683 (N_29683,N_20871,N_22855);
and U29684 (N_29684,N_20472,N_23694);
and U29685 (N_29685,N_24157,N_22703);
nor U29686 (N_29686,N_24002,N_22556);
or U29687 (N_29687,N_23521,N_20530);
or U29688 (N_29688,N_24504,N_20124);
nand U29689 (N_29689,N_21636,N_21065);
nand U29690 (N_29690,N_24089,N_23345);
xor U29691 (N_29691,N_20166,N_24338);
xnor U29692 (N_29692,N_23366,N_22694);
nand U29693 (N_29693,N_20176,N_20130);
xor U29694 (N_29694,N_21550,N_21251);
and U29695 (N_29695,N_22567,N_24947);
nand U29696 (N_29696,N_22013,N_20839);
and U29697 (N_29697,N_21195,N_22151);
xor U29698 (N_29698,N_21934,N_24144);
and U29699 (N_29699,N_22889,N_21160);
nor U29700 (N_29700,N_22962,N_20525);
and U29701 (N_29701,N_22944,N_23358);
nor U29702 (N_29702,N_22954,N_24019);
nand U29703 (N_29703,N_22121,N_22565);
nand U29704 (N_29704,N_23835,N_21780);
xor U29705 (N_29705,N_22733,N_23439);
or U29706 (N_29706,N_20293,N_20626);
or U29707 (N_29707,N_23334,N_22039);
and U29708 (N_29708,N_23547,N_20527);
nor U29709 (N_29709,N_24140,N_21750);
or U29710 (N_29710,N_21583,N_22418);
xor U29711 (N_29711,N_20852,N_22718);
or U29712 (N_29712,N_22877,N_20758);
or U29713 (N_29713,N_21078,N_20742);
nand U29714 (N_29714,N_21943,N_21450);
nand U29715 (N_29715,N_21569,N_23477);
or U29716 (N_29716,N_20284,N_24771);
xor U29717 (N_29717,N_21192,N_20710);
nand U29718 (N_29718,N_23703,N_22471);
or U29719 (N_29719,N_21853,N_23929);
xnor U29720 (N_29720,N_20934,N_21797);
xor U29721 (N_29721,N_23800,N_20239);
nor U29722 (N_29722,N_24733,N_22251);
nor U29723 (N_29723,N_21018,N_23507);
xnor U29724 (N_29724,N_23232,N_20866);
or U29725 (N_29725,N_20965,N_23562);
or U29726 (N_29726,N_20228,N_21428);
xnor U29727 (N_29727,N_22409,N_21097);
and U29728 (N_29728,N_23395,N_24960);
or U29729 (N_29729,N_22148,N_20957);
nand U29730 (N_29730,N_23800,N_22439);
or U29731 (N_29731,N_21874,N_21250);
nand U29732 (N_29732,N_21268,N_24833);
and U29733 (N_29733,N_24931,N_20306);
nor U29734 (N_29734,N_23453,N_23604);
or U29735 (N_29735,N_23502,N_24210);
xnor U29736 (N_29736,N_22180,N_20748);
nor U29737 (N_29737,N_20300,N_24093);
nor U29738 (N_29738,N_20780,N_23489);
xor U29739 (N_29739,N_24362,N_21143);
or U29740 (N_29740,N_24318,N_23957);
and U29741 (N_29741,N_22059,N_23935);
nor U29742 (N_29742,N_24840,N_24801);
and U29743 (N_29743,N_20665,N_22750);
nor U29744 (N_29744,N_23231,N_23140);
or U29745 (N_29745,N_23692,N_20484);
nand U29746 (N_29746,N_20737,N_24706);
xnor U29747 (N_29747,N_20070,N_22196);
nand U29748 (N_29748,N_23432,N_24652);
and U29749 (N_29749,N_23625,N_21451);
and U29750 (N_29750,N_21016,N_24091);
nor U29751 (N_29751,N_23442,N_24710);
nand U29752 (N_29752,N_23347,N_20592);
nand U29753 (N_29753,N_21177,N_24036);
nand U29754 (N_29754,N_20773,N_23655);
nand U29755 (N_29755,N_22835,N_21322);
nand U29756 (N_29756,N_23864,N_20232);
and U29757 (N_29757,N_23569,N_23461);
nor U29758 (N_29758,N_21214,N_21992);
xor U29759 (N_29759,N_21047,N_22885);
xor U29760 (N_29760,N_23473,N_23574);
nor U29761 (N_29761,N_24343,N_24919);
nand U29762 (N_29762,N_21027,N_21816);
and U29763 (N_29763,N_24921,N_23664);
xnor U29764 (N_29764,N_23001,N_22988);
or U29765 (N_29765,N_24871,N_22450);
and U29766 (N_29766,N_24600,N_21696);
xnor U29767 (N_29767,N_21979,N_24414);
and U29768 (N_29768,N_20300,N_24391);
and U29769 (N_29769,N_24778,N_22012);
nand U29770 (N_29770,N_24404,N_21334);
xnor U29771 (N_29771,N_20855,N_20212);
and U29772 (N_29772,N_22290,N_23087);
nor U29773 (N_29773,N_20429,N_22940);
and U29774 (N_29774,N_22424,N_23279);
nor U29775 (N_29775,N_24119,N_21785);
xnor U29776 (N_29776,N_23230,N_21231);
nand U29777 (N_29777,N_21680,N_23619);
nand U29778 (N_29778,N_23944,N_21793);
nor U29779 (N_29779,N_22092,N_24116);
and U29780 (N_29780,N_22841,N_22797);
and U29781 (N_29781,N_23528,N_24271);
or U29782 (N_29782,N_24683,N_23713);
nor U29783 (N_29783,N_20175,N_20159);
xor U29784 (N_29784,N_20689,N_22436);
or U29785 (N_29785,N_21306,N_21520);
xor U29786 (N_29786,N_22379,N_23615);
nor U29787 (N_29787,N_22036,N_23273);
or U29788 (N_29788,N_21350,N_24567);
and U29789 (N_29789,N_23342,N_21324);
nand U29790 (N_29790,N_22637,N_20879);
nor U29791 (N_29791,N_24394,N_22678);
or U29792 (N_29792,N_23053,N_24370);
nand U29793 (N_29793,N_20490,N_20210);
and U29794 (N_29794,N_22183,N_24173);
or U29795 (N_29795,N_20082,N_22921);
xnor U29796 (N_29796,N_22772,N_20869);
nand U29797 (N_29797,N_24742,N_20647);
xnor U29798 (N_29798,N_20351,N_24500);
nand U29799 (N_29799,N_21719,N_23981);
xor U29800 (N_29800,N_22168,N_21257);
and U29801 (N_29801,N_21136,N_24470);
or U29802 (N_29802,N_21977,N_20674);
nor U29803 (N_29803,N_20514,N_23779);
and U29804 (N_29804,N_20846,N_20820);
or U29805 (N_29805,N_23669,N_22492);
nand U29806 (N_29806,N_24537,N_20942);
nor U29807 (N_29807,N_23518,N_21817);
nor U29808 (N_29808,N_20162,N_24615);
and U29809 (N_29809,N_22965,N_24519);
nor U29810 (N_29810,N_24264,N_23859);
xnor U29811 (N_29811,N_24514,N_22769);
nor U29812 (N_29812,N_23955,N_24595);
xnor U29813 (N_29813,N_22248,N_24036);
and U29814 (N_29814,N_20197,N_21525);
nand U29815 (N_29815,N_22662,N_20940);
nand U29816 (N_29816,N_20121,N_24068);
nor U29817 (N_29817,N_23475,N_21881);
or U29818 (N_29818,N_22464,N_20914);
nand U29819 (N_29819,N_21550,N_21968);
nand U29820 (N_29820,N_22708,N_21973);
or U29821 (N_29821,N_21888,N_21914);
and U29822 (N_29822,N_22256,N_22311);
and U29823 (N_29823,N_24795,N_20830);
xnor U29824 (N_29824,N_24649,N_20613);
nand U29825 (N_29825,N_23589,N_21594);
nor U29826 (N_29826,N_23183,N_24006);
or U29827 (N_29827,N_23193,N_23871);
nor U29828 (N_29828,N_23360,N_20056);
and U29829 (N_29829,N_20859,N_21105);
and U29830 (N_29830,N_21945,N_24701);
nand U29831 (N_29831,N_23920,N_24123);
or U29832 (N_29832,N_22628,N_23807);
nand U29833 (N_29833,N_20067,N_22181);
nand U29834 (N_29834,N_20150,N_24838);
nand U29835 (N_29835,N_22233,N_20812);
nor U29836 (N_29836,N_24263,N_22927);
and U29837 (N_29837,N_22050,N_21038);
or U29838 (N_29838,N_20346,N_20070);
and U29839 (N_29839,N_24296,N_20488);
and U29840 (N_29840,N_22558,N_21716);
and U29841 (N_29841,N_21784,N_20382);
or U29842 (N_29842,N_24474,N_24436);
nor U29843 (N_29843,N_23199,N_20537);
and U29844 (N_29844,N_21097,N_22032);
or U29845 (N_29845,N_23808,N_23555);
nor U29846 (N_29846,N_21903,N_22114);
or U29847 (N_29847,N_24196,N_22897);
xor U29848 (N_29848,N_20004,N_23718);
nor U29849 (N_29849,N_22344,N_22409);
and U29850 (N_29850,N_23663,N_24356);
nor U29851 (N_29851,N_21331,N_24476);
nand U29852 (N_29852,N_22151,N_24508);
nand U29853 (N_29853,N_20643,N_22756);
or U29854 (N_29854,N_20718,N_21975);
xnor U29855 (N_29855,N_23371,N_24625);
nand U29856 (N_29856,N_23203,N_20464);
and U29857 (N_29857,N_21843,N_23467);
xnor U29858 (N_29858,N_20409,N_24905);
xnor U29859 (N_29859,N_23348,N_24071);
and U29860 (N_29860,N_24631,N_20967);
nand U29861 (N_29861,N_24436,N_21834);
and U29862 (N_29862,N_23243,N_24093);
nor U29863 (N_29863,N_20711,N_23347);
nand U29864 (N_29864,N_20232,N_24853);
or U29865 (N_29865,N_23911,N_24194);
nand U29866 (N_29866,N_21029,N_23601);
xnor U29867 (N_29867,N_23959,N_22458);
and U29868 (N_29868,N_22616,N_20361);
and U29869 (N_29869,N_23417,N_23581);
nor U29870 (N_29870,N_23899,N_24958);
nor U29871 (N_29871,N_22453,N_20033);
nor U29872 (N_29872,N_22815,N_20860);
xnor U29873 (N_29873,N_21877,N_24348);
nand U29874 (N_29874,N_20896,N_22334);
nor U29875 (N_29875,N_20265,N_21414);
and U29876 (N_29876,N_22874,N_23435);
nand U29877 (N_29877,N_23395,N_20373);
nor U29878 (N_29878,N_20461,N_21959);
or U29879 (N_29879,N_22184,N_22663);
and U29880 (N_29880,N_20593,N_20280);
or U29881 (N_29881,N_24632,N_24868);
or U29882 (N_29882,N_23865,N_23532);
nand U29883 (N_29883,N_23241,N_21147);
and U29884 (N_29884,N_23638,N_24732);
nand U29885 (N_29885,N_23285,N_22964);
nand U29886 (N_29886,N_20595,N_24557);
nand U29887 (N_29887,N_22198,N_20845);
nor U29888 (N_29888,N_22104,N_20058);
and U29889 (N_29889,N_22472,N_20153);
nand U29890 (N_29890,N_23584,N_24965);
or U29891 (N_29891,N_23202,N_22312);
xor U29892 (N_29892,N_24028,N_23563);
or U29893 (N_29893,N_23711,N_20249);
or U29894 (N_29894,N_20695,N_23394);
nand U29895 (N_29895,N_23499,N_20277);
nor U29896 (N_29896,N_20448,N_21382);
or U29897 (N_29897,N_24777,N_20710);
or U29898 (N_29898,N_22196,N_21347);
or U29899 (N_29899,N_20230,N_22704);
xnor U29900 (N_29900,N_24443,N_22883);
nand U29901 (N_29901,N_21046,N_20828);
nand U29902 (N_29902,N_24879,N_23068);
xnor U29903 (N_29903,N_23655,N_21998);
or U29904 (N_29904,N_21621,N_21746);
or U29905 (N_29905,N_22633,N_20752);
nand U29906 (N_29906,N_23608,N_22440);
nand U29907 (N_29907,N_20512,N_20239);
nand U29908 (N_29908,N_23171,N_23824);
and U29909 (N_29909,N_21777,N_24305);
xnor U29910 (N_29910,N_21297,N_23299);
nand U29911 (N_29911,N_22043,N_23728);
nor U29912 (N_29912,N_21562,N_21413);
xor U29913 (N_29913,N_22845,N_20177);
and U29914 (N_29914,N_20572,N_24323);
or U29915 (N_29915,N_21998,N_23756);
nor U29916 (N_29916,N_24801,N_21909);
nor U29917 (N_29917,N_22927,N_24656);
xor U29918 (N_29918,N_22494,N_20148);
xor U29919 (N_29919,N_24395,N_22922);
and U29920 (N_29920,N_20858,N_20549);
nor U29921 (N_29921,N_21836,N_22040);
nand U29922 (N_29922,N_21448,N_22455);
or U29923 (N_29923,N_23223,N_21217);
or U29924 (N_29924,N_23508,N_23803);
or U29925 (N_29925,N_23168,N_22155);
and U29926 (N_29926,N_23597,N_21949);
or U29927 (N_29927,N_21058,N_20132);
nor U29928 (N_29928,N_22040,N_20213);
and U29929 (N_29929,N_21505,N_21568);
nor U29930 (N_29930,N_21679,N_23165);
xnor U29931 (N_29931,N_21714,N_20524);
and U29932 (N_29932,N_20390,N_21289);
nor U29933 (N_29933,N_20840,N_22309);
nand U29934 (N_29934,N_22487,N_21907);
xor U29935 (N_29935,N_22463,N_24454);
nand U29936 (N_29936,N_22332,N_23470);
nor U29937 (N_29937,N_24618,N_21721);
nor U29938 (N_29938,N_21148,N_21641);
xnor U29939 (N_29939,N_21252,N_24977);
and U29940 (N_29940,N_20729,N_20092);
or U29941 (N_29941,N_23629,N_20546);
nor U29942 (N_29942,N_22309,N_24203);
nor U29943 (N_29943,N_23846,N_20953);
xor U29944 (N_29944,N_21581,N_20235);
or U29945 (N_29945,N_24836,N_20541);
nor U29946 (N_29946,N_22953,N_21938);
nand U29947 (N_29947,N_24340,N_23801);
and U29948 (N_29948,N_21159,N_24162);
or U29949 (N_29949,N_23412,N_20159);
nand U29950 (N_29950,N_22528,N_22303);
or U29951 (N_29951,N_24097,N_21815);
nand U29952 (N_29952,N_20067,N_21398);
xor U29953 (N_29953,N_23582,N_22007);
xnor U29954 (N_29954,N_22911,N_20491);
or U29955 (N_29955,N_22812,N_24332);
or U29956 (N_29956,N_21929,N_24967);
xor U29957 (N_29957,N_22962,N_20426);
or U29958 (N_29958,N_22067,N_21354);
or U29959 (N_29959,N_22021,N_21288);
nand U29960 (N_29960,N_24781,N_23295);
or U29961 (N_29961,N_22281,N_20147);
and U29962 (N_29962,N_20935,N_24910);
or U29963 (N_29963,N_21879,N_24104);
nand U29964 (N_29964,N_24862,N_21361);
nand U29965 (N_29965,N_23669,N_22098);
xnor U29966 (N_29966,N_22385,N_22801);
xor U29967 (N_29967,N_20875,N_23098);
nand U29968 (N_29968,N_24380,N_22913);
nand U29969 (N_29969,N_21180,N_22896);
or U29970 (N_29970,N_20400,N_24215);
nor U29971 (N_29971,N_23716,N_21193);
or U29972 (N_29972,N_23497,N_24455);
xor U29973 (N_29973,N_23279,N_21083);
and U29974 (N_29974,N_20825,N_21870);
or U29975 (N_29975,N_23183,N_23849);
xor U29976 (N_29976,N_22698,N_22136);
nand U29977 (N_29977,N_21416,N_22785);
nand U29978 (N_29978,N_22677,N_22620);
xor U29979 (N_29979,N_23514,N_24721);
nand U29980 (N_29980,N_20383,N_21675);
or U29981 (N_29981,N_21819,N_23511);
nand U29982 (N_29982,N_21599,N_24650);
nand U29983 (N_29983,N_23576,N_21437);
and U29984 (N_29984,N_22584,N_23373);
or U29985 (N_29985,N_22944,N_22625);
nand U29986 (N_29986,N_23938,N_24451);
xor U29987 (N_29987,N_22849,N_23578);
xor U29988 (N_29988,N_24356,N_23170);
nand U29989 (N_29989,N_22982,N_24589);
nand U29990 (N_29990,N_20335,N_23645);
xnor U29991 (N_29991,N_21483,N_22778);
and U29992 (N_29992,N_23828,N_21840);
or U29993 (N_29993,N_23627,N_23169);
nand U29994 (N_29994,N_22610,N_24641);
or U29995 (N_29995,N_23970,N_24061);
nand U29996 (N_29996,N_21976,N_20471);
and U29997 (N_29997,N_24554,N_21669);
or U29998 (N_29998,N_22213,N_24147);
nand U29999 (N_29999,N_23922,N_23258);
nand UO_0 (O_0,N_29004,N_27611);
xnor UO_1 (O_1,N_27949,N_27095);
nand UO_2 (O_2,N_29411,N_25955);
and UO_3 (O_3,N_25684,N_25435);
or UO_4 (O_4,N_28064,N_28161);
or UO_5 (O_5,N_29323,N_25085);
xnor UO_6 (O_6,N_29465,N_27636);
and UO_7 (O_7,N_28881,N_29246);
nand UO_8 (O_8,N_25102,N_25365);
or UO_9 (O_9,N_28891,N_28402);
nor UO_10 (O_10,N_25392,N_26159);
and UO_11 (O_11,N_29588,N_25787);
nand UO_12 (O_12,N_28810,N_26205);
and UO_13 (O_13,N_25798,N_27271);
nor UO_14 (O_14,N_25146,N_27999);
nand UO_15 (O_15,N_29338,N_27437);
nand UO_16 (O_16,N_29256,N_28256);
and UO_17 (O_17,N_25277,N_26847);
xnor UO_18 (O_18,N_26081,N_25581);
nand UO_19 (O_19,N_27819,N_25422);
nand UO_20 (O_20,N_26718,N_29079);
or UO_21 (O_21,N_29819,N_25883);
nand UO_22 (O_22,N_27871,N_29421);
nor UO_23 (O_23,N_29230,N_25157);
xnor UO_24 (O_24,N_29867,N_29591);
nor UO_25 (O_25,N_25998,N_28215);
nor UO_26 (O_26,N_29706,N_29606);
nor UO_27 (O_27,N_29959,N_28198);
nand UO_28 (O_28,N_29351,N_25379);
nor UO_29 (O_29,N_28766,N_29417);
and UO_30 (O_30,N_25282,N_27017);
or UO_31 (O_31,N_25710,N_25922);
and UO_32 (O_32,N_29412,N_29687);
xnor UO_33 (O_33,N_25994,N_26894);
nor UO_34 (O_34,N_25292,N_29294);
xor UO_35 (O_35,N_25527,N_26985);
or UO_36 (O_36,N_28708,N_28454);
and UO_37 (O_37,N_28597,N_26280);
or UO_38 (O_38,N_29488,N_27328);
and UO_39 (O_39,N_26442,N_25566);
or UO_40 (O_40,N_25417,N_26478);
and UO_41 (O_41,N_28712,N_26922);
nor UO_42 (O_42,N_26225,N_27002);
xnor UO_43 (O_43,N_26038,N_25805);
xor UO_44 (O_44,N_26012,N_29646);
nand UO_45 (O_45,N_27458,N_29542);
nand UO_46 (O_46,N_25224,N_27235);
or UO_47 (O_47,N_27743,N_26759);
nand UO_48 (O_48,N_28382,N_29193);
nand UO_49 (O_49,N_28264,N_27136);
nand UO_50 (O_50,N_26704,N_26360);
and UO_51 (O_51,N_29430,N_26519);
and UO_52 (O_52,N_27716,N_25553);
and UO_53 (O_53,N_26450,N_26145);
nor UO_54 (O_54,N_28574,N_25313);
nand UO_55 (O_55,N_27762,N_27050);
nand UO_56 (O_56,N_29868,N_25041);
or UO_57 (O_57,N_26813,N_29413);
and UO_58 (O_58,N_26185,N_25385);
and UO_59 (O_59,N_25381,N_28341);
nand UO_60 (O_60,N_25999,N_28463);
and UO_61 (O_61,N_26914,N_28831);
nand UO_62 (O_62,N_25055,N_25668);
nor UO_63 (O_63,N_28527,N_27178);
nor UO_64 (O_64,N_29858,N_25728);
nand UO_65 (O_65,N_29396,N_25757);
xor UO_66 (O_66,N_29124,N_26177);
or UO_67 (O_67,N_29291,N_28591);
nand UO_68 (O_68,N_27444,N_26976);
nand UO_69 (O_69,N_25968,N_29777);
and UO_70 (O_70,N_28553,N_29344);
or UO_71 (O_71,N_25620,N_25791);
nand UO_72 (O_72,N_26164,N_29697);
and UO_73 (O_73,N_26314,N_29084);
or UO_74 (O_74,N_25984,N_29804);
or UO_75 (O_75,N_28009,N_29494);
and UO_76 (O_76,N_27013,N_25934);
nand UO_77 (O_77,N_29933,N_26792);
or UO_78 (O_78,N_28495,N_25168);
nor UO_79 (O_79,N_25554,N_26586);
and UO_80 (O_80,N_28320,N_27335);
xor UO_81 (O_81,N_28767,N_28787);
and UO_82 (O_82,N_27098,N_25500);
nand UO_83 (O_83,N_29418,N_25842);
xnor UO_84 (O_84,N_29899,N_25558);
xor UO_85 (O_85,N_28261,N_27372);
and UO_86 (O_86,N_27710,N_25175);
or UO_87 (O_87,N_28177,N_26046);
xor UO_88 (O_88,N_29290,N_25119);
xnor UO_89 (O_89,N_29707,N_28423);
or UO_90 (O_90,N_27477,N_29714);
nor UO_91 (O_91,N_28583,N_29767);
and UO_92 (O_92,N_25497,N_28386);
xnor UO_93 (O_93,N_27185,N_29221);
or UO_94 (O_94,N_28410,N_27826);
and UO_95 (O_95,N_25359,N_26458);
or UO_96 (O_96,N_27784,N_29519);
or UO_97 (O_97,N_25104,N_27311);
nand UO_98 (O_98,N_26260,N_27209);
xnor UO_99 (O_99,N_25606,N_27918);
nand UO_100 (O_100,N_29579,N_26666);
nor UO_101 (O_101,N_27786,N_29699);
nor UO_102 (O_102,N_26346,N_25541);
nor UO_103 (O_103,N_28941,N_26231);
or UO_104 (O_104,N_29717,N_27968);
nand UO_105 (O_105,N_28197,N_25735);
or UO_106 (O_106,N_26900,N_25966);
nor UO_107 (O_107,N_27373,N_29340);
or UO_108 (O_108,N_25248,N_29050);
xnor UO_109 (O_109,N_27977,N_29968);
nand UO_110 (O_110,N_25557,N_28796);
xnor UO_111 (O_111,N_26270,N_27677);
nand UO_112 (O_112,N_27575,N_29378);
nand UO_113 (O_113,N_26155,N_27839);
and UO_114 (O_114,N_25380,N_25651);
nand UO_115 (O_115,N_26253,N_28458);
or UO_116 (O_116,N_29181,N_27141);
nand UO_117 (O_117,N_28594,N_29503);
nand UO_118 (O_118,N_28052,N_26910);
or UO_119 (O_119,N_29524,N_27899);
or UO_120 (O_120,N_28826,N_27508);
or UO_121 (O_121,N_26301,N_27020);
nand UO_122 (O_122,N_29327,N_27772);
nand UO_123 (O_123,N_27281,N_26141);
xnor UO_124 (O_124,N_26644,N_29754);
xor UO_125 (O_125,N_25077,N_25584);
or UO_126 (O_126,N_28652,N_27589);
nand UO_127 (O_127,N_28180,N_26026);
xor UO_128 (O_128,N_26182,N_26619);
nand UO_129 (O_129,N_25540,N_28360);
or UO_130 (O_130,N_25614,N_26028);
or UO_131 (O_131,N_27551,N_28647);
and UO_132 (O_132,N_27962,N_26543);
xor UO_133 (O_133,N_27646,N_25401);
and UO_134 (O_134,N_26534,N_27440);
nand UO_135 (O_135,N_26802,N_26748);
and UO_136 (O_136,N_27253,N_29280);
and UO_137 (O_137,N_27851,N_27985);
nand UO_138 (O_138,N_25216,N_27672);
nor UO_139 (O_139,N_29750,N_29628);
xor UO_140 (O_140,N_25771,N_29244);
xor UO_141 (O_141,N_27715,N_29955);
or UO_142 (O_142,N_26023,N_26661);
nand UO_143 (O_143,N_27807,N_29207);
xnor UO_144 (O_144,N_26703,N_26475);
nand UO_145 (O_145,N_28589,N_27724);
nor UO_146 (O_146,N_26248,N_27180);
or UO_147 (O_147,N_25159,N_27401);
or UO_148 (O_148,N_26629,N_27693);
xor UO_149 (O_149,N_25743,N_29405);
or UO_150 (O_150,N_29424,N_27536);
nor UO_151 (O_151,N_27549,N_27601);
or UO_152 (O_152,N_27728,N_28867);
and UO_153 (O_153,N_26467,N_25658);
xor UO_154 (O_154,N_29609,N_25486);
or UO_155 (O_155,N_29170,N_29179);
nor UO_156 (O_156,N_28640,N_26364);
or UO_157 (O_157,N_25238,N_25799);
nor UO_158 (O_158,N_25496,N_29775);
nand UO_159 (O_159,N_25349,N_26656);
xnor UO_160 (O_160,N_29574,N_28559);
nand UO_161 (O_161,N_25773,N_28300);
and UO_162 (O_162,N_28966,N_26549);
xor UO_163 (O_163,N_26263,N_26927);
nand UO_164 (O_164,N_29060,N_27937);
xnor UO_165 (O_165,N_26669,N_27391);
or UO_166 (O_166,N_26842,N_26909);
xor UO_167 (O_167,N_28332,N_27315);
or UO_168 (O_168,N_28890,N_29624);
nor UO_169 (O_169,N_29477,N_28937);
nand UO_170 (O_170,N_29448,N_27358);
nor UO_171 (O_171,N_27932,N_25149);
nand UO_172 (O_172,N_26795,N_28724);
or UO_173 (O_173,N_26550,N_25666);
or UO_174 (O_174,N_29157,N_27245);
nand UO_175 (O_175,N_27658,N_25580);
and UO_176 (O_176,N_29737,N_25910);
or UO_177 (O_177,N_25258,N_25266);
nand UO_178 (O_178,N_28073,N_27800);
nor UO_179 (O_179,N_25640,N_28173);
nand UO_180 (O_180,N_25779,N_27431);
and UO_181 (O_181,N_25253,N_26431);
or UO_182 (O_182,N_28631,N_26339);
and UO_183 (O_183,N_25649,N_26864);
and UO_184 (O_184,N_25090,N_28380);
nor UO_185 (O_185,N_26489,N_25836);
or UO_186 (O_186,N_26818,N_26501);
or UO_187 (O_187,N_29657,N_26297);
nor UO_188 (O_188,N_26265,N_26216);
or UO_189 (O_189,N_28610,N_26076);
nand UO_190 (O_190,N_25869,N_28242);
nand UO_191 (O_191,N_27044,N_28419);
nand UO_192 (O_192,N_29969,N_27043);
and UO_193 (O_193,N_26585,N_26060);
xor UO_194 (O_194,N_27473,N_25488);
nor UO_195 (O_195,N_29390,N_25888);
and UO_196 (O_196,N_28619,N_29645);
and UO_197 (O_197,N_28883,N_25308);
or UO_198 (O_198,N_28845,N_28836);
and UO_199 (O_199,N_25702,N_26875);
nand UO_200 (O_200,N_29942,N_29202);
nand UO_201 (O_201,N_25671,N_26469);
or UO_202 (O_202,N_29009,N_27320);
and UO_203 (O_203,N_29753,N_27324);
nor UO_204 (O_204,N_26686,N_25720);
and UO_205 (O_205,N_26101,N_29065);
xnor UO_206 (O_206,N_26744,N_27892);
nand UO_207 (O_207,N_26485,N_26123);
nor UO_208 (O_208,N_29811,N_26781);
or UO_209 (O_209,N_25827,N_29473);
xor UO_210 (O_210,N_28493,N_27353);
nor UO_211 (O_211,N_25698,N_28475);
nand UO_212 (O_212,N_25324,N_26241);
and UO_213 (O_213,N_26685,N_29677);
or UO_214 (O_214,N_28224,N_25840);
and UO_215 (O_215,N_25474,N_26139);
or UO_216 (O_216,N_27507,N_27631);
nor UO_217 (O_217,N_27986,N_26390);
or UO_218 (O_218,N_27299,N_25029);
nand UO_219 (O_219,N_28804,N_25074);
xnor UO_220 (O_220,N_26142,N_27448);
and UO_221 (O_221,N_25348,N_25767);
nand UO_222 (O_222,N_27304,N_28905);
nor UO_223 (O_223,N_29878,N_28351);
nand UO_224 (O_224,N_26430,N_27598);
nor UO_225 (O_225,N_25515,N_27843);
xnor UO_226 (O_226,N_28540,N_27836);
nand UO_227 (O_227,N_26518,N_26162);
nor UO_228 (O_228,N_28479,N_27896);
nand UO_229 (O_229,N_27751,N_27198);
or UO_230 (O_230,N_25036,N_28279);
xor UO_231 (O_231,N_27689,N_26775);
xnor UO_232 (O_232,N_28289,N_26327);
xor UO_233 (O_233,N_26844,N_27614);
and UO_234 (O_234,N_29526,N_28538);
nor UO_235 (O_235,N_29178,N_25949);
nor UO_236 (O_236,N_25412,N_28006);
nor UO_237 (O_237,N_25592,N_27120);
nand UO_238 (O_238,N_27476,N_25001);
or UO_239 (O_239,N_28771,N_25636);
nor UO_240 (O_240,N_27132,N_25302);
or UO_241 (O_241,N_25096,N_25645);
nor UO_242 (O_242,N_25697,N_26342);
nand UO_243 (O_243,N_26020,N_27835);
nand UO_244 (O_244,N_28576,N_28319);
or UO_245 (O_245,N_25147,N_29691);
nand UO_246 (O_246,N_26257,N_27798);
nand UO_247 (O_247,N_26414,N_27778);
xnor UO_248 (O_248,N_26063,N_25415);
nor UO_249 (O_249,N_29077,N_25075);
and UO_250 (O_250,N_26895,N_27640);
xnor UO_251 (O_251,N_25492,N_29563);
and UO_252 (O_252,N_28872,N_26868);
xor UO_253 (O_253,N_28682,N_28666);
and UO_254 (O_254,N_27267,N_27058);
or UO_255 (O_255,N_29188,N_26244);
nor UO_256 (O_256,N_26646,N_27456);
xor UO_257 (O_257,N_29040,N_26183);
or UO_258 (O_258,N_27422,N_28513);
or UO_259 (O_259,N_27138,N_29683);
nor UO_260 (O_260,N_28762,N_26168);
or UO_261 (O_261,N_26069,N_26382);
nand UO_262 (O_262,N_29892,N_29423);
and UO_263 (O_263,N_28176,N_29884);
nor UO_264 (O_264,N_29748,N_29229);
nand UO_265 (O_265,N_27961,N_27505);
and UO_266 (O_266,N_28118,N_25115);
and UO_267 (O_267,N_26279,N_25221);
xor UO_268 (O_268,N_25199,N_29293);
xor UO_269 (O_269,N_28770,N_26799);
nand UO_270 (O_270,N_25375,N_27201);
or UO_271 (O_271,N_27106,N_26486);
xnor UO_272 (O_272,N_28698,N_28587);
and UO_273 (O_273,N_28888,N_25859);
xor UO_274 (O_274,N_28040,N_27880);
or UO_275 (O_275,N_26240,N_25953);
nand UO_276 (O_276,N_28798,N_25173);
or UO_277 (O_277,N_27517,N_25816);
nand UO_278 (O_278,N_27639,N_26783);
xor UO_279 (O_279,N_25863,N_25594);
xnor UO_280 (O_280,N_25367,N_27021);
nor UO_281 (O_281,N_29001,N_26548);
xor UO_282 (O_282,N_29794,N_27935);
and UO_283 (O_283,N_27648,N_27889);
or UO_284 (O_284,N_28748,N_25093);
nor UO_285 (O_285,N_25895,N_29635);
nor UO_286 (O_286,N_25366,N_25449);
or UO_287 (O_287,N_28756,N_25942);
nor UO_288 (O_288,N_25692,N_25897);
xnor UO_289 (O_289,N_26660,N_27171);
nor UO_290 (O_290,N_26740,N_28433);
or UO_291 (O_291,N_29847,N_29303);
nor UO_292 (O_292,N_29788,N_25761);
or UO_293 (O_293,N_29316,N_25034);
xnor UO_294 (O_294,N_26055,N_29665);
nor UO_295 (O_295,N_29130,N_28022);
nand UO_296 (O_296,N_26187,N_26989);
xnor UO_297 (O_297,N_25681,N_26239);
and UO_298 (O_298,N_29891,N_25194);
and UO_299 (O_299,N_25995,N_26150);
or UO_300 (O_300,N_28927,N_29204);
xnor UO_301 (O_301,N_25711,N_29778);
or UO_302 (O_302,N_28135,N_25874);
xnor UO_303 (O_303,N_29556,N_28144);
nor UO_304 (O_304,N_26305,N_25819);
nor UO_305 (O_305,N_26956,N_28859);
xnor UO_306 (O_306,N_28938,N_29926);
or UO_307 (O_307,N_27722,N_28633);
or UO_308 (O_308,N_27101,N_29605);
and UO_309 (O_309,N_29408,N_28949);
and UO_310 (O_310,N_25355,N_28719);
nand UO_311 (O_311,N_25975,N_28835);
xor UO_312 (O_312,N_29976,N_26546);
or UO_313 (O_313,N_25521,N_25650);
or UO_314 (O_314,N_29116,N_29099);
or UO_315 (O_315,N_27321,N_26603);
and UO_316 (O_316,N_28657,N_28954);
xor UO_317 (O_317,N_26705,N_26533);
nand UO_318 (O_318,N_25178,N_29101);
nand UO_319 (O_319,N_26878,N_27610);
or UO_320 (O_320,N_26338,N_25101);
or UO_321 (O_321,N_28885,N_27590);
xor UO_322 (O_322,N_26521,N_28194);
xor UO_323 (O_323,N_25271,N_29436);
and UO_324 (O_324,N_25120,N_25334);
xnor UO_325 (O_325,N_29560,N_28365);
xnor UO_326 (O_326,N_26291,N_27071);
nor UO_327 (O_327,N_25335,N_25220);
xnor UO_328 (O_328,N_25160,N_25089);
and UO_329 (O_329,N_25861,N_29527);
or UO_330 (O_330,N_29032,N_27958);
and UO_331 (O_331,N_27433,N_25233);
xnor UO_332 (O_332,N_27741,N_28057);
xor UO_333 (O_333,N_27602,N_25007);
and UO_334 (O_334,N_27497,N_26313);
and UO_335 (O_335,N_26275,N_27801);
xor UO_336 (O_336,N_26545,N_28229);
xor UO_337 (O_337,N_27654,N_25475);
xor UO_338 (O_338,N_28939,N_29225);
or UO_339 (O_339,N_29023,N_28361);
nand UO_340 (O_340,N_27666,N_28325);
xor UO_341 (O_341,N_25161,N_29371);
and UO_342 (O_342,N_28039,N_26919);
and UO_343 (O_343,N_27176,N_29007);
xnor UO_344 (O_344,N_26793,N_27822);
nand UO_345 (O_345,N_27107,N_26075);
and UO_346 (O_346,N_26427,N_27459);
and UO_347 (O_347,N_25240,N_29738);
nand UO_348 (O_348,N_25441,N_25807);
nand UO_349 (O_349,N_29272,N_27649);
and UO_350 (O_350,N_27965,N_29956);
xor UO_351 (O_351,N_28016,N_29156);
and UO_352 (O_352,N_27396,N_28107);
or UO_353 (O_353,N_26846,N_29607);
nor UO_354 (O_354,N_26093,N_25462);
or UO_355 (O_355,N_29318,N_26970);
and UO_356 (O_356,N_29342,N_25894);
or UO_357 (O_357,N_26609,N_28068);
or UO_358 (O_358,N_29307,N_26428);
nor UO_359 (O_359,N_25543,N_27055);
and UO_360 (O_360,N_27665,N_29839);
and UO_361 (O_361,N_26065,N_25165);
xnor UO_362 (O_362,N_27695,N_26607);
xor UO_363 (O_363,N_27768,N_27070);
nand UO_364 (O_364,N_28664,N_25709);
and UO_365 (O_365,N_28500,N_26833);
or UO_366 (O_366,N_26008,N_26932);
nand UO_367 (O_367,N_27014,N_28374);
nor UO_368 (O_368,N_29982,N_27637);
or UO_369 (O_369,N_26356,N_26329);
nand UO_370 (O_370,N_27696,N_27414);
nor UO_371 (O_371,N_29871,N_28496);
nor UO_372 (O_372,N_29639,N_29020);
xor UO_373 (O_373,N_26250,N_25418);
xnor UO_374 (O_374,N_26689,N_29627);
nor UO_375 (O_375,N_27090,N_28321);
nand UO_376 (O_376,N_25331,N_26676);
nand UO_377 (O_377,N_29584,N_27523);
nor UO_378 (O_378,N_26432,N_29948);
nand UO_379 (O_379,N_27690,N_25846);
or UO_380 (O_380,N_28847,N_25522);
nor UO_381 (O_381,N_27870,N_27399);
nand UO_382 (O_382,N_28362,N_26048);
xnor UO_383 (O_383,N_27876,N_27703);
xnor UO_384 (O_384,N_28800,N_28451);
nor UO_385 (O_385,N_29015,N_26973);
nor UO_386 (O_386,N_27467,N_27330);
and UO_387 (O_387,N_25058,N_26217);
nand UO_388 (O_388,N_27723,N_28252);
xor UO_389 (O_389,N_26196,N_26163);
nand UO_390 (O_390,N_29733,N_26706);
nor UO_391 (O_391,N_28662,N_28575);
nor UO_392 (O_392,N_27712,N_29110);
nor UO_393 (O_393,N_25320,N_26344);
or UO_394 (O_394,N_29837,N_29118);
and UO_395 (O_395,N_25634,N_29144);
and UO_396 (O_396,N_25124,N_26944);
and UO_397 (O_397,N_29541,N_27184);
or UO_398 (O_398,N_26321,N_25733);
xnor UO_399 (O_399,N_26707,N_28219);
nor UO_400 (O_400,N_26400,N_28673);
and UO_401 (O_401,N_26936,N_25621);
or UO_402 (O_402,N_29428,N_26653);
nand UO_403 (O_403,N_25826,N_29770);
nor UO_404 (O_404,N_27969,N_28926);
nor UO_405 (O_405,N_28685,N_26491);
or UO_406 (O_406,N_29636,N_26127);
and UO_407 (O_407,N_26268,N_25598);
xor UO_408 (O_408,N_27763,N_28731);
xor UO_409 (O_409,N_28822,N_29914);
xor UO_410 (O_410,N_27256,N_26210);
and UO_411 (O_411,N_29385,N_29026);
xor UO_412 (O_412,N_27332,N_27114);
nor UO_413 (O_413,N_27750,N_25063);
nand UO_414 (O_414,N_25914,N_26719);
nor UO_415 (O_415,N_28813,N_25516);
nand UO_416 (O_416,N_27901,N_29194);
nand UO_417 (O_417,N_26194,N_27490);
or UO_418 (O_418,N_26134,N_26935);
nor UO_419 (O_419,N_25502,N_28745);
nor UO_420 (O_420,N_25033,N_25834);
or UO_421 (O_421,N_29135,N_25166);
xor UO_422 (O_422,N_25509,N_29036);
xor UO_423 (O_423,N_26912,N_28047);
nand UO_424 (O_424,N_28750,N_28776);
xnor UO_425 (O_425,N_26304,N_29059);
nand UO_426 (O_426,N_25377,N_25996);
xnor UO_427 (O_427,N_26535,N_25900);
xor UO_428 (O_428,N_27177,N_28923);
xor UO_429 (O_429,N_26100,N_26153);
or UO_430 (O_430,N_29096,N_28537);
nor UO_431 (O_431,N_26045,N_26453);
xor UO_432 (O_432,N_29068,N_29128);
or UO_433 (O_433,N_27862,N_28946);
or UO_434 (O_434,N_25469,N_27699);
nor UO_435 (O_435,N_29616,N_28175);
xnor UO_436 (O_436,N_26276,N_25106);
and UO_437 (O_437,N_26790,N_26105);
or UO_438 (O_438,N_25629,N_26295);
nor UO_439 (O_439,N_29550,N_29719);
or UO_440 (O_440,N_28568,N_26133);
nand UO_441 (O_441,N_28049,N_29592);
and UO_442 (O_442,N_29994,N_26353);
and UO_443 (O_443,N_26882,N_26907);
nor UO_444 (O_444,N_28508,N_28084);
xor UO_445 (O_445,N_29793,N_26117);
and UO_446 (O_446,N_27694,N_26119);
nor UO_447 (O_447,N_28424,N_25425);
nand UO_448 (O_448,N_26865,N_26886);
xnor UO_449 (O_449,N_29952,N_27280);
and UO_450 (O_450,N_25847,N_26680);
and UO_451 (O_451,N_25588,N_27063);
nand UO_452 (O_452,N_29896,N_28687);
and UO_453 (O_453,N_26975,N_26939);
nor UO_454 (O_454,N_27331,N_25408);
nand UO_455 (O_455,N_26480,N_25915);
nand UO_456 (O_456,N_29445,N_28518);
and UO_457 (O_457,N_27834,N_29763);
or UO_458 (O_458,N_27126,N_25571);
nand UO_459 (O_459,N_26817,N_29276);
nor UO_460 (O_460,N_26222,N_27539);
xnor UO_461 (O_461,N_28406,N_25843);
nand UO_462 (O_462,N_28914,N_29910);
nand UO_463 (O_463,N_25751,N_25245);
and UO_464 (O_464,N_27584,N_25409);
or UO_465 (O_465,N_28048,N_25616);
or UO_466 (O_466,N_28742,N_28226);
nor UO_467 (O_467,N_29393,N_29735);
or UO_468 (O_468,N_27153,N_27576);
xor UO_469 (O_469,N_25289,N_26166);
nor UO_470 (O_470,N_27167,N_29983);
xor UO_471 (O_471,N_25822,N_29213);
nand UO_472 (O_472,N_29078,N_28803);
and UO_473 (O_473,N_26351,N_28014);
xnor UO_474 (O_474,N_28653,N_29829);
nand UO_475 (O_475,N_27895,N_28674);
or UO_476 (O_476,N_26099,N_27488);
xor UO_477 (O_477,N_25991,N_26892);
or UO_478 (O_478,N_25719,N_25973);
and UO_479 (O_479,N_25899,N_25964);
nor UO_480 (O_480,N_28412,N_28171);
xnor UO_481 (O_481,N_29484,N_28490);
or UO_482 (O_482,N_25740,N_29565);
nand UO_483 (O_483,N_25346,N_27556);
and UO_484 (O_484,N_28447,N_29022);
nand UO_485 (O_485,N_25078,N_27150);
nor UO_486 (O_486,N_27621,N_28728);
nor UO_487 (O_487,N_27343,N_29780);
xnor UO_488 (O_488,N_27947,N_27754);
xor UO_489 (O_489,N_28765,N_28227);
nor UO_490 (O_490,N_28050,N_27482);
xor UO_491 (O_491,N_25979,N_27673);
xnor UO_492 (O_492,N_28830,N_27592);
and UO_493 (O_493,N_25397,N_26654);
nor UO_494 (O_494,N_25215,N_27118);
xor UO_495 (O_495,N_29637,N_25184);
and UO_496 (O_496,N_27510,N_29838);
nor UO_497 (O_497,N_29715,N_28579);
nand UO_498 (O_498,N_29168,N_26403);
nand UO_499 (O_499,N_28864,N_26696);
and UO_500 (O_500,N_27309,N_26897);
xor UO_501 (O_501,N_29854,N_27365);
xnor UO_502 (O_502,N_26204,N_27349);
nand UO_503 (O_503,N_27973,N_29602);
nand UO_504 (O_504,N_28270,N_25971);
xnor UO_505 (O_505,N_28753,N_25918);
nor UO_506 (O_506,N_29450,N_26371);
xnor UO_507 (O_507,N_27036,N_27755);
or UO_508 (O_508,N_27500,N_27222);
nand UO_509 (O_509,N_26841,N_29089);
nand UO_510 (O_510,N_25809,N_29017);
nor UO_511 (O_511,N_28366,N_25057);
nor UO_512 (O_512,N_26316,N_27618);
nand UO_513 (O_513,N_27561,N_27405);
nor UO_514 (O_514,N_26622,N_29133);
xnor UO_515 (O_515,N_27630,N_28970);
and UO_516 (O_516,N_27368,N_29456);
xnor UO_517 (O_517,N_25311,N_29198);
and UO_518 (O_518,N_27221,N_25848);
or UO_519 (O_519,N_27912,N_28201);
and UO_520 (O_520,N_27173,N_28820);
or UO_521 (O_521,N_26537,N_25976);
nand UO_522 (O_522,N_29594,N_29284);
and UO_523 (O_523,N_27922,N_26899);
nand UO_524 (O_524,N_25031,N_28959);
nand UO_525 (O_525,N_26186,N_29082);
xor UO_526 (O_526,N_26971,N_29500);
or UO_527 (O_527,N_29785,N_26626);
nor UO_528 (O_528,N_28222,N_27116);
nor UO_529 (O_529,N_27019,N_28192);
and UO_530 (O_530,N_25977,N_26213);
xor UO_531 (O_531,N_29000,N_28134);
and UO_532 (O_532,N_29568,N_29803);
nand UO_533 (O_533,N_29905,N_26074);
xnor UO_534 (O_534,N_28861,N_27538);
nand UO_535 (O_535,N_28302,N_28672);
or UO_536 (O_536,N_27345,N_28465);
nand UO_537 (O_537,N_28623,N_25353);
or UO_538 (O_538,N_26831,N_27115);
xnor UO_539 (O_539,N_29362,N_25860);
or UO_540 (O_540,N_29160,N_25630);
or UO_541 (O_541,N_25021,N_28977);
xnor UO_542 (O_542,N_26710,N_28506);
or UO_543 (O_543,N_26395,N_27387);
nor UO_544 (O_544,N_26980,N_25028);
nand UO_545 (O_545,N_29196,N_26852);
nor UO_546 (O_546,N_25832,N_27298);
nand UO_547 (O_547,N_26621,N_26218);
nor UO_548 (O_548,N_25749,N_27407);
or UO_549 (O_549,N_26031,N_25717);
xor UO_550 (O_550,N_26730,N_28387);
nor UO_551 (O_551,N_27327,N_28277);
xor UO_552 (O_552,N_27068,N_27030);
xor UO_553 (O_553,N_25069,N_29578);
or UO_554 (O_554,N_27082,N_29523);
and UO_555 (O_555,N_25276,N_28541);
and UO_556 (O_556,N_26264,N_28809);
nand UO_557 (O_557,N_28695,N_25884);
or UO_558 (O_558,N_26800,N_29998);
or UO_559 (O_559,N_26633,N_29561);
xor UO_560 (O_560,N_28240,N_29262);
nand UO_561 (O_561,N_27216,N_25455);
and UO_562 (O_562,N_28523,N_27364);
xor UO_563 (O_563,N_25003,N_25940);
and UO_564 (O_564,N_27890,N_27042);
xor UO_565 (O_565,N_29950,N_26820);
xnor UO_566 (O_566,N_26372,N_25011);
nor UO_567 (O_567,N_28313,N_29384);
xor UO_568 (O_568,N_27297,N_28703);
and UO_569 (O_569,N_25081,N_26328);
or UO_570 (O_570,N_25369,N_25695);
nand UO_571 (O_571,N_25990,N_25326);
xnor UO_572 (O_572,N_25162,N_25685);
nor UO_573 (O_573,N_26735,N_25505);
nor UO_574 (O_574,N_28310,N_27874);
and UO_575 (O_575,N_28205,N_26021);
nand UO_576 (O_576,N_29521,N_29751);
and UO_577 (O_577,N_26592,N_26124);
nor UO_578 (O_578,N_28799,N_28667);
and UO_579 (O_579,N_29504,N_28886);
or UO_580 (O_580,N_26681,N_29097);
and UO_581 (O_581,N_25019,N_26331);
and UO_582 (O_582,N_26605,N_27130);
or UO_583 (O_583,N_25189,N_26345);
or UO_584 (O_584,N_28900,N_28160);
nand UO_585 (O_585,N_29790,N_28834);
nand UO_586 (O_586,N_25641,N_27838);
xnor UO_587 (O_587,N_25009,N_25841);
nand UO_588 (O_588,N_29885,N_26815);
xor UO_589 (O_589,N_28550,N_27902);
nand UO_590 (O_590,N_29274,N_25654);
nor UO_591 (O_591,N_29177,N_25983);
or UO_592 (O_592,N_25696,N_29723);
and UO_593 (O_593,N_29608,N_26363);
nor UO_594 (O_594,N_27052,N_26033);
nand UO_595 (O_595,N_28346,N_25706);
or UO_596 (O_596,N_28033,N_28641);
and UO_597 (O_597,N_27886,N_26623);
or UO_598 (O_598,N_27810,N_27830);
nand UO_599 (O_599,N_28096,N_27380);
xor UO_600 (O_600,N_26261,N_29805);
and UO_601 (O_601,N_26374,N_26287);
and UO_602 (O_602,N_29343,N_27217);
nand UO_603 (O_603,N_25192,N_25116);
or UO_604 (O_604,N_26758,N_26255);
and UO_605 (O_605,N_28741,N_26447);
and UO_606 (O_606,N_28760,N_27652);
xnor UO_607 (O_607,N_27322,N_26315);
nand UO_608 (O_608,N_27229,N_27733);
xor UO_609 (O_609,N_25913,N_25845);
nor UO_610 (O_610,N_27037,N_25008);
nor UO_611 (O_611,N_25477,N_25788);
nand UO_612 (O_612,N_28385,N_25098);
and UO_613 (O_613,N_28854,N_28123);
and UO_614 (O_614,N_29853,N_26195);
nor UO_615 (O_615,N_29852,N_29286);
xnor UO_616 (O_616,N_28440,N_29985);
and UO_617 (O_617,N_27499,N_26175);
or UO_618 (O_618,N_28392,N_26503);
xnor UO_619 (O_619,N_29127,N_26358);
nand UO_620 (O_620,N_28413,N_26034);
nor UO_621 (O_621,N_29978,N_25878);
xnor UO_622 (O_622,N_25204,N_29814);
nor UO_623 (O_623,N_26002,N_26029);
nand UO_624 (O_624,N_29145,N_28437);
xnor UO_625 (O_625,N_28778,N_25434);
nor UO_626 (O_626,N_26078,N_27752);
xor UO_627 (O_627,N_28738,N_25622);
and UO_628 (O_628,N_25775,N_26446);
or UO_629 (O_629,N_26006,N_28036);
xnor UO_630 (O_630,N_28120,N_26207);
nand UO_631 (O_631,N_27894,N_25176);
nand UO_632 (O_632,N_27520,N_25354);
and UO_633 (O_633,N_28649,N_28987);
and UO_634 (O_634,N_29622,N_25185);
and UO_635 (O_635,N_27620,N_27608);
nor UO_636 (O_636,N_29587,N_29085);
nor UO_637 (O_637,N_26479,N_27140);
and UO_638 (O_638,N_28116,N_26594);
nand UO_639 (O_639,N_28853,N_29031);
and UO_640 (O_640,N_28172,N_25793);
nand UO_641 (O_641,N_25993,N_26566);
or UO_642 (O_642,N_29442,N_25802);
nand UO_643 (O_643,N_27295,N_25792);
nand UO_644 (O_644,N_27319,N_26544);
nand UO_645 (O_645,N_27197,N_27785);
nor UO_646 (O_646,N_25235,N_28729);
and UO_647 (O_647,N_27558,N_28127);
nor UO_648 (O_648,N_29555,N_27936);
nor UO_649 (O_649,N_27053,N_26460);
or UO_650 (O_650,N_28411,N_25817);
nand UO_651 (O_651,N_28978,N_27707);
xor UO_652 (O_652,N_29237,N_27687);
or UO_653 (O_653,N_25902,N_26872);
and UO_654 (O_654,N_25446,N_26816);
xnor UO_655 (O_655,N_27831,N_27435);
nor UO_656 (O_656,N_28314,N_26916);
xnor UO_657 (O_657,N_28915,N_26924);
xor UO_658 (O_658,N_28863,N_29946);
nand UO_659 (O_659,N_28395,N_29358);
xor UO_660 (O_660,N_29849,N_26942);
xor UO_661 (O_661,N_27208,N_27072);
nand UO_662 (O_662,N_28654,N_25551);
nand UO_663 (O_663,N_26172,N_26017);
and UO_664 (O_664,N_27156,N_28292);
xor UO_665 (O_665,N_25426,N_26131);
xor UO_666 (O_666,N_28935,N_26913);
nand UO_667 (O_667,N_28678,N_29115);
xor UO_668 (O_668,N_25784,N_26674);
or UO_669 (O_669,N_27721,N_26402);
or UO_670 (O_670,N_27276,N_26409);
nand UO_671 (O_671,N_28422,N_28721);
nor UO_672 (O_672,N_25693,N_28442);
xor UO_673 (O_673,N_29419,N_29247);
nand UO_674 (O_674,N_29787,N_29782);
nand UO_675 (O_675,N_25273,N_28702);
and UO_676 (O_676,N_27516,N_25479);
nand UO_677 (O_677,N_29368,N_26979);
xor UO_678 (O_678,N_29328,N_25583);
and UO_679 (O_679,N_26373,N_25602);
and UO_680 (O_680,N_28995,N_27152);
xor UO_681 (O_681,N_25656,N_28059);
nand UO_682 (O_682,N_27641,N_25507);
nor UO_683 (O_683,N_26112,N_29459);
xor UO_684 (O_684,N_27502,N_26873);
nor UO_685 (O_685,N_25909,N_27760);
nand UO_686 (O_686,N_27739,N_25803);
nand UO_687 (O_687,N_26902,N_29652);
nor UO_688 (O_688,N_25285,N_26529);
and UO_689 (O_689,N_25601,N_27738);
nand UO_690 (O_690,N_27147,N_29306);
xor UO_691 (O_691,N_25625,N_25830);
xnor UO_692 (O_692,N_27662,N_27594);
and UO_693 (O_693,N_28851,N_27159);
nor UO_694 (O_694,N_27410,N_28095);
and UO_695 (O_695,N_29154,N_27306);
and UO_696 (O_696,N_28464,N_29146);
xnor UO_697 (O_697,N_28549,N_29766);
xor UO_698 (O_698,N_26836,N_25811);
or UO_699 (O_699,N_29902,N_26378);
or UO_700 (O_700,N_25203,N_27362);
and UO_701 (O_701,N_25323,N_26893);
or UO_702 (O_702,N_29648,N_25609);
xor UO_703 (O_703,N_25135,N_25631);
nand UO_704 (O_704,N_25373,N_25665);
and UO_705 (O_705,N_28195,N_29961);
nand UO_706 (O_706,N_25384,N_25188);
nor UO_707 (O_707,N_29136,N_26407);
or UO_708 (O_708,N_27770,N_29075);
or UO_709 (O_709,N_29016,N_28477);
xnor UO_710 (O_710,N_26234,N_28913);
nor UO_711 (O_711,N_25260,N_25789);
xnor UO_712 (O_712,N_28852,N_26884);
xor UO_713 (O_713,N_27092,N_25088);
and UO_714 (O_714,N_29768,N_27469);
xor UO_715 (O_715,N_26129,N_28593);
and UO_716 (O_716,N_28301,N_29251);
xnor UO_717 (O_717,N_29831,N_26826);
xnor UO_718 (O_718,N_27031,N_25347);
nor UO_719 (O_719,N_26408,N_27916);
nor UO_720 (O_720,N_25072,N_28817);
nand UO_721 (O_721,N_28114,N_27214);
nand UO_722 (O_722,N_27578,N_29585);
nor UO_723 (O_723,N_29433,N_25560);
nand UO_724 (O_724,N_27457,N_28485);
nand UO_725 (O_725,N_28216,N_26988);
nor UO_726 (O_726,N_25187,N_29440);
and UO_727 (O_727,N_27511,N_25988);
nand UO_728 (O_728,N_28482,N_28492);
and UO_729 (O_729,N_27411,N_26934);
and UO_730 (O_730,N_26597,N_27815);
nor UO_731 (O_731,N_28206,N_29489);
nor UO_732 (O_732,N_26388,N_25317);
or UO_733 (O_733,N_25084,N_29562);
and UO_734 (O_734,N_27904,N_26057);
or UO_735 (O_735,N_27190,N_26589);
xnor UO_736 (O_736,N_25091,N_25778);
and UO_737 (O_737,N_27817,N_26224);
nand UO_738 (O_738,N_29206,N_28684);
and UO_739 (O_739,N_25724,N_29600);
and UO_740 (O_740,N_28187,N_28725);
nand UO_741 (O_741,N_25056,N_28501);
nand UO_742 (O_742,N_29458,N_26835);
nor UO_743 (O_743,N_25197,N_28605);
and UO_744 (O_744,N_29641,N_25961);
and UO_745 (O_745,N_27504,N_28957);
or UO_746 (O_746,N_25404,N_26284);
or UO_747 (O_747,N_28326,N_29088);
and UO_748 (O_748,N_27325,N_28711);
xor UO_749 (O_749,N_27606,N_27352);
xnor UO_750 (O_750,N_25746,N_29166);
nand UO_751 (O_751,N_25738,N_26986);
nand UO_752 (O_752,N_26192,N_29334);
and UO_753 (O_753,N_29245,N_25201);
xnor UO_754 (O_754,N_28701,N_28012);
and UO_755 (O_755,N_25514,N_26786);
and UO_756 (O_756,N_27604,N_28691);
xnor UO_757 (O_757,N_26005,N_27472);
nor UO_758 (O_758,N_27416,N_25158);
and UO_759 (O_759,N_29326,N_28783);
or UO_760 (O_760,N_28470,N_29604);
xnor UO_761 (O_761,N_26564,N_25825);
xor UO_762 (O_762,N_26832,N_28990);
nor UO_763 (O_763,N_26051,N_27392);
or UO_764 (O_764,N_28903,N_27318);
nor UO_765 (O_765,N_26044,N_28309);
nor UO_766 (O_766,N_28061,N_27644);
nand UO_767 (O_767,N_26951,N_29776);
nor UO_768 (O_768,N_28035,N_27291);
and UO_769 (O_769,N_29314,N_26915);
nand UO_770 (O_770,N_25340,N_29784);
or UO_771 (O_771,N_26784,N_27314);
or UO_772 (O_772,N_29924,N_29512);
and UO_773 (O_773,N_29298,N_28162);
nand UO_774 (O_774,N_28491,N_27193);
nor UO_775 (O_775,N_28102,N_28910);
or UO_776 (O_776,N_27264,N_26606);
nand UO_777 (O_777,N_28965,N_27162);
and UO_778 (O_778,N_27746,N_29045);
xor UO_779 (O_779,N_29236,N_29283);
and UO_780 (O_780,N_25957,N_25981);
xnor UO_781 (O_781,N_28637,N_27521);
xnor UO_782 (O_782,N_26049,N_29481);
or UO_783 (O_783,N_26570,N_25518);
nor UO_784 (O_784,N_26639,N_29673);
and UO_785 (O_785,N_29506,N_25428);
or UO_786 (O_786,N_29631,N_25542);
nor UO_787 (O_787,N_28584,N_26354);
nor UO_788 (O_788,N_27847,N_27104);
and UO_789 (O_789,N_25639,N_25850);
nand UO_790 (O_790,N_28081,N_29138);
nand UO_791 (O_791,N_29980,N_26084);
nand UO_792 (O_792,N_25569,N_29669);
or UO_793 (O_793,N_26383,N_25016);
nor UO_794 (O_794,N_25877,N_26115);
or UO_795 (O_795,N_25229,N_27914);
and UO_796 (O_796,N_26655,N_26966);
nor UO_797 (O_797,N_28899,N_29629);
and UO_798 (O_798,N_29876,N_28934);
and UO_799 (O_799,N_27420,N_28401);
nand UO_800 (O_800,N_25241,N_28155);
nand UO_801 (O_801,N_29508,N_27869);
xor UO_802 (O_802,N_26420,N_25643);
xnor UO_803 (O_803,N_25919,N_28388);
xnor UO_804 (O_804,N_26256,N_27974);
or UO_805 (O_805,N_26776,N_26757);
and UO_806 (O_806,N_25338,N_26319);
or UO_807 (O_807,N_29414,N_29114);
nand UO_808 (O_808,N_25391,N_27883);
xor UO_809 (O_809,N_28067,N_27139);
xnor UO_810 (O_810,N_27375,N_25974);
nor UO_811 (O_811,N_26869,N_26303);
nand UO_812 (O_812,N_25786,N_29183);
nand UO_813 (O_813,N_26470,N_27006);
xnor UO_814 (O_814,N_26242,N_25246);
and UO_815 (O_815,N_25678,N_26532);
nor UO_816 (O_816,N_29125,N_26000);
xor UO_817 (O_817,N_29965,N_29522);
and UO_818 (O_818,N_28105,N_26659);
nor UO_819 (O_819,N_29501,N_26948);
nand UO_820 (O_820,N_26197,N_26302);
and UO_821 (O_821,N_29879,N_27480);
nand UO_822 (O_822,N_27527,N_27400);
nand UO_823 (O_823,N_29155,N_26160);
and UO_824 (O_824,N_28858,N_29552);
nand UO_825 (O_825,N_28316,N_29028);
or UO_826 (O_826,N_27725,N_25597);
and UO_827 (O_827,N_27691,N_28746);
xnor UO_828 (O_828,N_26611,N_27850);
and UO_829 (O_829,N_28772,N_26077);
nor UO_830 (O_830,N_28722,N_27857);
xnor UO_831 (O_831,N_26380,N_26281);
nand UO_832 (O_832,N_29809,N_29510);
and UO_833 (O_833,N_29895,N_26463);
xnor UO_834 (O_834,N_28250,N_29173);
nor UO_835 (O_835,N_25691,N_27357);
or UO_836 (O_836,N_25087,N_29640);
or UO_837 (O_837,N_29725,N_25905);
xnor UO_838 (O_838,N_28376,N_28489);
or UO_839 (O_839,N_26996,N_27356);
and UO_840 (O_840,N_26514,N_27853);
xnor UO_841 (O_841,N_27603,N_25890);
xor UO_842 (O_842,N_29996,N_26307);
nand UO_843 (O_843,N_26381,N_27142);
and UO_844 (O_844,N_25127,N_26226);
xor UO_845 (O_845,N_27438,N_28275);
or UO_846 (O_846,N_25181,N_26412);
nand UO_847 (O_847,N_27704,N_29577);
nor UO_848 (O_848,N_26122,N_27670);
and UO_849 (O_849,N_27821,N_27048);
or UO_850 (O_850,N_29241,N_28807);
nand UO_851 (O_851,N_28249,N_25682);
and UO_852 (O_852,N_28150,N_26928);
nand UO_853 (O_853,N_25242,N_29263);
or UO_854 (O_854,N_26616,N_26994);
nor UO_855 (O_855,N_29261,N_29575);
and UO_856 (O_856,N_29312,N_25596);
nand UO_857 (O_857,N_25332,N_26392);
xnor UO_858 (O_858,N_26251,N_27891);
nand UO_859 (O_859,N_28827,N_25935);
and UO_860 (O_860,N_26523,N_29043);
nand UO_861 (O_861,N_29216,N_25150);
nor UO_862 (O_862,N_28129,N_28925);
or UO_863 (O_863,N_26755,N_29200);
or UO_864 (O_864,N_25345,N_25287);
nand UO_865 (O_865,N_28359,N_29208);
nor UO_866 (O_866,N_28236,N_28692);
or UO_867 (O_867,N_27051,N_28015);
nor UO_868 (O_868,N_28897,N_25406);
or UO_869 (O_869,N_28873,N_26289);
or UO_870 (O_870,N_29397,N_29964);
xor UO_871 (O_871,N_25228,N_29012);
nor UO_872 (O_872,N_25451,N_25010);
xor UO_873 (O_873,N_26874,N_28381);
nor UO_874 (O_874,N_29826,N_26451);
and UO_875 (O_875,N_26959,N_28775);
xor UO_876 (O_876,N_25259,N_27868);
nand UO_877 (O_877,N_27957,N_26238);
and UO_878 (O_878,N_25278,N_26227);
nand UO_879 (O_879,N_25179,N_29643);
and UO_880 (O_880,N_26398,N_27946);
xnor UO_881 (O_881,N_28573,N_29499);
or UO_882 (O_882,N_28159,N_27102);
xnor UO_883 (O_883,N_25796,N_27844);
nor UO_884 (O_884,N_27212,N_29802);
nor UO_885 (O_885,N_29027,N_27661);
or UO_886 (O_886,N_26727,N_29210);
and UO_887 (O_887,N_26797,N_29546);
or UO_888 (O_888,N_29507,N_28021);
or UO_889 (O_889,N_25690,N_26269);
nand UO_890 (O_890,N_27697,N_26278);
nand UO_891 (O_891,N_28607,N_29139);
and UO_892 (O_892,N_27808,N_27305);
and UO_893 (O_893,N_26433,N_27659);
nand UO_894 (O_894,N_26498,N_26219);
nor UO_895 (O_895,N_28231,N_26796);
xor UO_896 (O_896,N_25210,N_26713);
nor UO_897 (O_897,N_29870,N_26384);
and UO_898 (O_898,N_27837,N_26571);
nor UO_899 (O_899,N_26788,N_28769);
xnor UO_900 (O_900,N_29439,N_28306);
and UO_901 (O_901,N_25109,N_27626);
or UO_902 (O_902,N_25871,N_28119);
nor UO_903 (O_903,N_29570,N_28260);
and UO_904 (O_904,N_29386,N_27232);
and UO_905 (O_905,N_27065,N_27781);
or UO_906 (O_906,N_28543,N_28730);
and UO_907 (O_907,N_27073,N_26721);
and UO_908 (O_908,N_29772,N_29223);
xor UO_909 (O_909,N_25352,N_27569);
xnor UO_910 (O_910,N_27591,N_26288);
xnor UO_911 (O_911,N_29679,N_26066);
xor UO_912 (O_912,N_28940,N_26778);
and UO_913 (O_913,N_25587,N_27960);
and UO_914 (O_914,N_26949,N_28971);
nand UO_915 (O_915,N_29253,N_29295);
or UO_916 (O_916,N_29731,N_27442);
xnor UO_917 (O_917,N_28986,N_27123);
xor UO_918 (O_918,N_28426,N_28335);
nand UO_919 (O_919,N_26881,N_27586);
xnor UO_920 (O_920,N_26426,N_28005);
nor UO_921 (O_921,N_25499,N_26090);
nand UO_922 (O_922,N_28768,N_28737);
or UO_923 (O_923,N_27284,N_28315);
xor UO_924 (O_924,N_27230,N_28663);
nand UO_925 (O_925,N_29363,N_27215);
nand UO_926 (O_926,N_26581,N_25667);
xor UO_927 (O_927,N_29619,N_26860);
nor UO_928 (O_928,N_28011,N_27287);
or UO_929 (O_929,N_29618,N_29740);
and UO_930 (O_930,N_25398,N_28906);
nor UO_931 (O_931,N_29469,N_27669);
and UO_932 (O_932,N_25297,N_28718);
nand UO_933 (O_933,N_28562,N_28478);
xor UO_934 (O_934,N_28536,N_29400);
nand UO_935 (O_935,N_25941,N_28268);
nand UO_936 (O_936,N_25208,N_25038);
xnor UO_937 (O_937,N_25431,N_29713);
nand UO_938 (O_938,N_26130,N_28077);
nor UO_939 (O_939,N_26156,N_27100);
xnor UO_940 (O_940,N_28000,N_27820);
and UO_941 (O_941,N_28601,N_27301);
nor UO_942 (O_942,N_28403,N_27954);
nand UO_943 (O_943,N_27047,N_28356);
or UO_944 (O_944,N_27720,N_25647);
xor UO_945 (O_945,N_27701,N_25211);
nand UO_946 (O_946,N_26449,N_27108);
xor UO_947 (O_947,N_27252,N_26734);
or UO_948 (O_948,N_28816,N_28244);
xor UO_949 (O_949,N_26953,N_27263);
nor UO_950 (O_950,N_27645,N_29755);
or UO_951 (O_951,N_28616,N_28908);
or UO_952 (O_952,N_26751,N_28348);
or UO_953 (O_953,N_26527,N_29668);
or UO_954 (O_954,N_28344,N_29977);
nor UO_955 (O_955,N_29148,N_28473);
nand UO_956 (O_956,N_27418,N_28397);
and UO_957 (O_957,N_29250,N_25312);
nor UO_958 (O_958,N_25524,N_27593);
xor UO_959 (O_959,N_25448,N_28818);
or UO_960 (O_960,N_28866,N_25926);
and UO_961 (O_961,N_25931,N_29791);
xnor UO_962 (O_962,N_27537,N_26500);
nand UO_963 (O_963,N_27110,N_25163);
xor UO_964 (O_964,N_28613,N_29476);
or UO_965 (O_965,N_26368,N_26513);
xnor UO_966 (O_966,N_26397,N_25837);
nor UO_967 (O_967,N_29387,N_29844);
nand UO_968 (O_968,N_27719,N_26672);
nor UO_969 (O_969,N_28080,N_27125);
or UO_970 (O_970,N_29310,N_26618);
nand UO_971 (O_971,N_25680,N_27445);
and UO_972 (O_972,N_28777,N_27628);
xor UO_973 (O_973,N_27852,N_26838);
and UO_974 (O_974,N_26054,N_26750);
and UO_975 (O_975,N_27244,N_26311);
xor UO_976 (O_976,N_26526,N_27385);
nor UO_977 (O_977,N_27317,N_29199);
xnor UO_978 (O_978,N_26435,N_27124);
nand UO_979 (O_979,N_25873,N_26885);
nand UO_980 (O_980,N_27466,N_29812);
or UO_981 (O_981,N_25864,N_25933);
nor UO_982 (O_982,N_27560,N_25766);
xnor UO_983 (O_983,N_28468,N_29761);
or UO_984 (O_984,N_29765,N_29920);
or UO_985 (O_985,N_26937,N_29692);
and UO_986 (O_986,N_28874,N_28153);
xor UO_987 (O_987,N_25167,N_26697);
xnor UO_988 (O_988,N_27761,N_26461);
nand UO_989 (O_989,N_29757,N_25526);
xnor UO_990 (O_990,N_27224,N_29862);
and UO_991 (O_991,N_29302,N_26845);
and UO_992 (O_992,N_26330,N_29861);
nor UO_993 (O_993,N_25866,N_27863);
nand UO_994 (O_994,N_29287,N_29391);
nand UO_995 (O_995,N_26508,N_26663);
or UO_996 (O_996,N_29169,N_25903);
xor UO_997 (O_997,N_27394,N_27419);
nor UO_998 (O_998,N_28739,N_27028);
nand UO_999 (O_999,N_27825,N_29822);
nand UO_1000 (O_1000,N_27934,N_25896);
nand UO_1001 (O_1001,N_26632,N_27228);
nand UO_1002 (O_1002,N_27683,N_29708);
and UO_1003 (O_1003,N_28764,N_28082);
and UO_1004 (O_1004,N_29090,N_26551);
xor UO_1005 (O_1005,N_26361,N_26670);
xnor UO_1006 (O_1006,N_26857,N_25950);
or UO_1007 (O_1007,N_27086,N_25407);
nand UO_1008 (O_1008,N_27128,N_28305);
or UO_1009 (O_1009,N_27981,N_25655);
and UO_1010 (O_1010,N_26348,N_29859);
xor UO_1011 (O_1011,N_29935,N_27971);
nand UO_1012 (O_1012,N_29598,N_25214);
and UO_1013 (O_1013,N_25128,N_28293);
and UO_1014 (O_1014,N_28519,N_26138);
nand UO_1015 (O_1015,N_26930,N_28782);
xor UO_1016 (O_1016,N_27441,N_27338);
nand UO_1017 (O_1017,N_28131,N_25829);
and UO_1018 (O_1018,N_26179,N_29346);
nand UO_1019 (O_1019,N_26274,N_28199);
and UO_1020 (O_1020,N_27023,N_25790);
nor UO_1021 (O_1021,N_26052,N_26125);
and UO_1022 (O_1022,N_26764,N_26567);
or UO_1023 (O_1023,N_25471,N_29132);
xor UO_1024 (O_1024,N_26152,N_26917);
and UO_1025 (O_1025,N_28697,N_27991);
nor UO_1026 (O_1026,N_26309,N_27938);
or UO_1027 (O_1027,N_28714,N_27550);
xnor UO_1028 (O_1028,N_27740,N_29372);
nand UO_1029 (O_1029,N_25776,N_25018);
xor UO_1030 (O_1030,N_27204,N_29409);
xnor UO_1031 (O_1031,N_28304,N_27265);
or UO_1032 (O_1032,N_27682,N_29907);
nor UO_1033 (O_1033,N_28425,N_29672);
nand UO_1034 (O_1034,N_26602,N_26741);
xor UO_1035 (O_1035,N_25610,N_26114);
and UO_1036 (O_1036,N_29927,N_27117);
nand UO_1037 (O_1037,N_25328,N_29845);
nand UO_1038 (O_1038,N_26807,N_28331);
nand UO_1039 (O_1039,N_25318,N_26804);
and UO_1040 (O_1040,N_29257,N_26285);
nor UO_1041 (O_1041,N_29887,N_25257);
nand UO_1042 (O_1042,N_28951,N_27027);
nor UO_1043 (O_1043,N_26334,N_25562);
nand UO_1044 (O_1044,N_29185,N_29345);
or UO_1045 (O_1045,N_28283,N_26931);
xor UO_1046 (O_1046,N_27905,N_27463);
xnor UO_1047 (O_1047,N_27452,N_25833);
and UO_1048 (O_1048,N_26448,N_27885);
nor UO_1049 (O_1049,N_26386,N_26471);
and UO_1050 (O_1050,N_27103,N_29163);
or UO_1051 (O_1051,N_26839,N_29543);
or UO_1052 (O_1052,N_29218,N_25694);
nand UO_1053 (O_1053,N_29589,N_25454);
and UO_1054 (O_1054,N_25963,N_29538);
xor UO_1055 (O_1055,N_27155,N_26497);
or UO_1056 (O_1056,N_25113,N_28024);
or UO_1057 (O_1057,N_28202,N_26563);
or UO_1058 (O_1058,N_28483,N_29149);
nor UO_1059 (O_1059,N_26766,N_26267);
nand UO_1060 (O_1060,N_25067,N_29437);
or UO_1061 (O_1061,N_25563,N_28604);
nor UO_1062 (O_1062,N_27449,N_28715);
and UO_1063 (O_1063,N_29799,N_28571);
nand UO_1064 (O_1064,N_28955,N_26714);
and UO_1065 (O_1065,N_27660,N_26001);
nor UO_1066 (O_1066,N_29332,N_26198);
nor UO_1067 (O_1067,N_26135,N_29900);
nor UO_1068 (O_1068,N_29264,N_25605);
and UO_1069 (O_1069,N_25337,N_25892);
nor UO_1070 (O_1070,N_28138,N_29300);
or UO_1071 (O_1071,N_28043,N_28004);
nor UO_1072 (O_1072,N_29051,N_26439);
xnor UO_1073 (O_1073,N_27623,N_28111);
xor UO_1074 (O_1074,N_28019,N_28615);
nand UO_1075 (O_1075,N_25987,N_25708);
xnor UO_1076 (O_1076,N_29712,N_29171);
nor UO_1077 (O_1077,N_26165,N_26904);
and UO_1078 (O_1078,N_26843,N_28122);
nand UO_1079 (O_1079,N_25364,N_27430);
nand UO_1080 (O_1080,N_28570,N_26733);
xor UO_1081 (O_1081,N_29472,N_29100);
nand UO_1082 (O_1082,N_25648,N_25363);
nand UO_1083 (O_1083,N_29704,N_29944);
nand UO_1084 (O_1084,N_29671,N_26015);
and UO_1085 (O_1085,N_25117,N_26193);
nand UO_1086 (O_1086,N_29487,N_26393);
or UO_1087 (O_1087,N_26791,N_29581);
nand UO_1088 (O_1088,N_28149,N_29582);
xnor UO_1089 (O_1089,N_27129,N_29086);
nor UO_1090 (O_1090,N_28870,N_25304);
or UO_1091 (O_1091,N_29842,N_26823);
nor UO_1092 (O_1092,N_26025,N_26889);
nor UO_1093 (O_1093,N_29756,N_29856);
nand UO_1094 (O_1094,N_27567,N_25753);
nor UO_1095 (O_1095,N_29655,N_26798);
xor UO_1096 (O_1096,N_29873,N_27787);
xnor UO_1097 (O_1097,N_28643,N_29685);
nand UO_1098 (O_1098,N_29449,N_25700);
and UO_1099 (O_1099,N_28415,N_26466);
or UO_1100 (O_1100,N_28840,N_26083);
nand UO_1101 (O_1101,N_26905,N_27069);
or UO_1102 (O_1102,N_29106,N_27833);
nand UO_1103 (O_1103,N_25099,N_29422);
xor UO_1104 (O_1104,N_26507,N_27062);
and UO_1105 (O_1105,N_25207,N_25765);
xnor UO_1106 (O_1106,N_27258,N_28868);
nand UO_1107 (O_1107,N_27379,N_26336);
or UO_1108 (O_1108,N_26073,N_25948);
or UO_1109 (O_1109,N_25399,N_29795);
nor UO_1110 (O_1110,N_28363,N_27060);
xnor UO_1111 (O_1111,N_27160,N_25481);
nor UO_1112 (O_1112,N_26943,N_27486);
nor UO_1113 (O_1113,N_29509,N_25818);
nand UO_1114 (O_1114,N_25568,N_29573);
nand UO_1115 (O_1115,N_26717,N_29150);
xor UO_1116 (O_1116,N_25059,N_27564);
nand UO_1117 (O_1117,N_26712,N_25429);
nor UO_1118 (O_1118,N_28487,N_26983);
or UO_1119 (O_1119,N_25820,N_26082);
and UO_1120 (O_1120,N_29482,N_28833);
xnor UO_1121 (O_1121,N_28404,N_26118);
nand UO_1122 (O_1122,N_29848,N_28298);
and UO_1123 (O_1123,N_25145,N_29309);
or UO_1124 (O_1124,N_28548,N_27206);
xnor UO_1125 (O_1125,N_26777,N_25756);
xor UO_1126 (O_1126,N_29092,N_27832);
nor UO_1127 (O_1127,N_29771,N_29462);
nor UO_1128 (O_1128,N_27432,N_29827);
nand UO_1129 (O_1129,N_26462,N_25660);
nor UO_1130 (O_1130,N_27625,N_28158);
xor UO_1131 (O_1131,N_25432,N_26030);
nand UO_1132 (O_1132,N_28763,N_29676);
nand UO_1133 (O_1133,N_26298,N_25148);
and UO_1134 (O_1134,N_27088,N_28294);
nor UO_1135 (O_1135,N_28030,N_27668);
nand UO_1136 (O_1136,N_28694,N_27749);
xor UO_1137 (O_1137,N_25844,N_29744);
and UO_1138 (O_1138,N_29240,N_27806);
nand UO_1139 (O_1139,N_25076,N_25747);
xor UO_1140 (O_1140,N_26173,N_28734);
xor UO_1141 (O_1141,N_29586,N_29747);
xor UO_1142 (O_1142,N_26610,N_25590);
and UO_1143 (O_1143,N_28524,N_26059);
and UO_1144 (O_1144,N_28399,N_26490);
nand UO_1145 (O_1145,N_28045,N_25851);
nor UO_1146 (O_1146,N_25064,N_28706);
nand UO_1147 (O_1147,N_25624,N_28113);
and UO_1148 (O_1148,N_28556,N_29117);
or UO_1149 (O_1149,N_29894,N_25513);
xnor UO_1150 (O_1150,N_27788,N_29866);
and UO_1151 (O_1151,N_26455,N_25582);
and UO_1152 (O_1152,N_25674,N_26923);
or UO_1153 (O_1153,N_25881,N_25122);
nand UO_1154 (O_1154,N_27524,N_25286);
or UO_1155 (O_1155,N_25236,N_29603);
nand UO_1156 (O_1156,N_26699,N_26861);
nor UO_1157 (O_1157,N_26377,N_26419);
and UO_1158 (O_1158,N_25300,N_28846);
or UO_1159 (O_1159,N_29662,N_29467);
nand UO_1160 (O_1160,N_29339,N_26539);
or UO_1161 (O_1161,N_25015,N_28688);
and UO_1162 (O_1162,N_26515,N_27953);
nor UO_1163 (O_1163,N_28156,N_26413);
nand UO_1164 (O_1164,N_25239,N_25932);
nand UO_1165 (O_1165,N_27681,N_27656);
nand UO_1166 (O_1166,N_26128,N_26582);
nor UO_1167 (O_1167,N_27266,N_25741);
xor UO_1168 (O_1168,N_27849,N_27545);
nor UO_1169 (O_1169,N_26530,N_29042);
nand UO_1170 (O_1170,N_27341,N_25256);
or UO_1171 (O_1171,N_27491,N_26600);
and UO_1172 (O_1172,N_25839,N_29214);
nand UO_1173 (O_1173,N_27312,N_29490);
or UO_1174 (O_1174,N_28996,N_29700);
nor UO_1175 (O_1175,N_26391,N_25298);
or UO_1176 (O_1176,N_25858,N_29019);
nor UO_1177 (O_1177,N_29454,N_26459);
xnor UO_1178 (O_1178,N_29407,N_28450);
nand UO_1179 (O_1179,N_25388,N_27684);
and UO_1180 (O_1180,N_29690,N_28909);
nor UO_1181 (O_1181,N_28056,N_29705);
or UO_1182 (O_1182,N_29464,N_28806);
and UO_1183 (O_1183,N_26890,N_27211);
nand UO_1184 (O_1184,N_27323,N_27667);
nand UO_1185 (O_1185,N_26888,N_26032);
nor UO_1186 (O_1186,N_27270,N_29457);
or UO_1187 (O_1187,N_27346,N_26188);
nand UO_1188 (O_1188,N_25887,N_29554);
and UO_1189 (O_1189,N_28106,N_28671);
nor UO_1190 (O_1190,N_26058,N_29817);
nor UO_1191 (O_1191,N_25712,N_28407);
and UO_1192 (O_1192,N_29243,N_25764);
or UO_1193 (O_1193,N_28880,N_25321);
nand UO_1194 (O_1194,N_26110,N_26424);
nand UO_1195 (O_1195,N_25947,N_29505);
nand UO_1196 (O_1196,N_27303,N_29932);
xor UO_1197 (O_1197,N_29872,N_26091);
or UO_1198 (O_1198,N_25254,N_29874);
xnor UO_1199 (O_1199,N_27846,N_25022);
or UO_1200 (O_1200,N_29989,N_26673);
and UO_1201 (O_1201,N_26266,N_27540);
nor UO_1202 (O_1202,N_28713,N_25485);
or UO_1203 (O_1203,N_27926,N_26387);
or UO_1204 (O_1204,N_28555,N_25281);
nand UO_1205 (O_1205,N_27427,N_28071);
and UO_1206 (O_1206,N_29709,N_28580);
nand UO_1207 (O_1207,N_29427,N_25755);
nand UO_1208 (O_1208,N_27532,N_27363);
or UO_1209 (O_1209,N_26190,N_28375);
and UO_1210 (O_1210,N_29703,N_28752);
and UO_1211 (O_1211,N_28705,N_27526);
nor UO_1212 (O_1212,N_29365,N_26596);
xnor UO_1213 (O_1213,N_25112,N_28747);
or UO_1214 (O_1214,N_27395,N_28645);
xor UO_1215 (O_1215,N_26590,N_26562);
nor UO_1216 (O_1216,N_26911,N_25937);
xor UO_1217 (O_1217,N_27487,N_29595);
nor UO_1218 (O_1218,N_25723,N_26612);
or UO_1219 (O_1219,N_26340,N_26443);
nor UO_1220 (O_1220,N_29260,N_25467);
or UO_1221 (O_1221,N_27827,N_26591);
nand UO_1222 (O_1222,N_25136,N_29992);
xor UO_1223 (O_1223,N_29002,N_28347);
or UO_1224 (O_1224,N_26317,N_28639);
and UO_1225 (O_1225,N_25828,N_29335);
nor UO_1226 (O_1226,N_26576,N_27040);
xor UO_1227 (O_1227,N_29320,N_28754);
xor UO_1228 (O_1228,N_25652,N_28794);
xor UO_1229 (O_1229,N_29774,N_26047);
nand UO_1230 (O_1230,N_28961,N_26824);
nor UO_1231 (O_1231,N_28832,N_25307);
xnor UO_1232 (O_1232,N_27685,N_26925);
xor UO_1233 (O_1233,N_28010,N_25519);
xnor UO_1234 (O_1234,N_25810,N_27111);
nor UO_1235 (O_1235,N_25303,N_27074);
xor UO_1236 (O_1236,N_25879,N_28948);
and UO_1237 (O_1237,N_29288,N_27326);
nand UO_1238 (O_1238,N_29654,N_25000);
and UO_1239 (O_1239,N_29836,N_26945);
nor UO_1240 (O_1240,N_27941,N_26604);
and UO_1241 (O_1241,N_25628,N_27413);
or UO_1242 (O_1242,N_27742,N_29108);
xnor UO_1243 (O_1243,N_25263,N_29141);
or UO_1244 (O_1244,N_27091,N_29281);
or UO_1245 (O_1245,N_28710,N_29516);
xor UO_1246 (O_1246,N_25284,N_25689);
and UO_1247 (O_1247,N_25325,N_27635);
nor UO_1248 (O_1248,N_26109,N_25050);
nor UO_1249 (O_1249,N_25376,N_28531);
or UO_1250 (O_1250,N_28869,N_28709);
or UO_1251 (O_1251,N_28079,N_27927);
xnor UO_1252 (O_1252,N_29821,N_28488);
nor UO_1253 (O_1253,N_29925,N_27951);
or UO_1254 (O_1254,N_29493,N_27767);
xnor UO_1255 (O_1255,N_28428,N_25472);
nor UO_1256 (O_1256,N_25670,N_25414);
and UO_1257 (O_1257,N_27254,N_27081);
nor UO_1258 (O_1258,N_28644,N_25371);
or UO_1259 (O_1259,N_25856,N_26667);
and UO_1260 (O_1260,N_28324,N_26294);
or UO_1261 (O_1261,N_25528,N_29373);
nand UO_1262 (O_1262,N_27079,N_29818);
xor UO_1263 (O_1263,N_28193,N_29651);
and UO_1264 (O_1264,N_29333,N_26310);
or UO_1265 (O_1265,N_26552,N_28062);
or UO_1266 (O_1266,N_25559,N_28223);
nand UO_1267 (O_1267,N_28497,N_27686);
and UO_1268 (O_1268,N_26867,N_26955);
and UO_1269 (O_1269,N_25748,N_29698);
nor UO_1270 (O_1270,N_25105,N_28191);
nor UO_1271 (O_1271,N_26136,N_27005);
nor UO_1272 (O_1272,N_25688,N_27813);
xnor UO_1273 (O_1273,N_28507,N_28823);
nand UO_1274 (O_1274,N_29883,N_29693);
nand UO_1275 (O_1275,N_28190,N_29270);
and UO_1276 (O_1276,N_26982,N_27000);
nor UO_1277 (O_1277,N_27557,N_28291);
nor UO_1278 (O_1278,N_26999,N_29444);
nor UO_1279 (O_1279,N_28204,N_25760);
or UO_1280 (O_1280,N_27008,N_29292);
nor UO_1281 (O_1281,N_28857,N_29806);
nor UO_1282 (O_1282,N_29539,N_27942);
nand UO_1283 (O_1283,N_26389,N_25480);
xor UO_1284 (O_1284,N_25868,N_27175);
nor UO_1285 (O_1285,N_26350,N_26668);
nor UO_1286 (O_1286,N_28773,N_26312);
nor UO_1287 (O_1287,N_26296,N_25437);
xor UO_1288 (O_1288,N_28353,N_28720);
xor UO_1289 (O_1289,N_25035,N_29701);
nand UO_1290 (O_1290,N_26811,N_26584);
and UO_1291 (O_1291,N_29227,N_26926);
and UO_1292 (O_1292,N_29081,N_28620);
nor UO_1293 (O_1293,N_29633,N_25305);
nor UO_1294 (O_1294,N_28805,N_29410);
or UO_1295 (O_1295,N_27568,N_28774);
or UO_1296 (O_1296,N_28658,N_27300);
and UO_1297 (O_1297,N_27484,N_27617);
nor UO_1298 (O_1298,N_25923,N_29813);
and UO_1299 (O_1299,N_28287,N_29808);
nor UO_1300 (O_1300,N_26089,N_26771);
or UO_1301 (O_1301,N_27634,N_27478);
nand UO_1302 (O_1302,N_25506,N_27003);
xnor UO_1303 (O_1303,N_27533,N_25137);
or UO_1304 (O_1304,N_29353,N_29957);
and UO_1305 (O_1305,N_25886,N_29716);
or UO_1306 (O_1306,N_26472,N_27577);
and UO_1307 (O_1307,N_25885,N_26399);
nor UO_1308 (O_1308,N_25024,N_28848);
and UO_1309 (O_1309,N_26417,N_25193);
nor UO_1310 (O_1310,N_26858,N_28931);
and UO_1311 (O_1311,N_29625,N_29979);
or UO_1312 (O_1312,N_29005,N_25854);
nand UO_1313 (O_1313,N_26773,N_29938);
nand UO_1314 (O_1314,N_28928,N_26014);
and UO_1315 (O_1315,N_28608,N_25027);
xor UO_1316 (O_1316,N_26728,N_29840);
or UO_1317 (O_1317,N_26202,N_28018);
xnor UO_1318 (O_1318,N_28209,N_29987);
and UO_1319 (O_1319,N_27039,N_25536);
nand UO_1320 (O_1320,N_26137,N_27615);
nand UO_1321 (O_1321,N_29906,N_29728);
or UO_1322 (O_1322,N_28408,N_28904);
or UO_1323 (O_1323,N_26042,N_27250);
nor UO_1324 (O_1324,N_28632,N_29759);
nand UO_1325 (O_1325,N_27348,N_29446);
xor UO_1326 (O_1326,N_28251,N_26682);
nand UO_1327 (O_1327,N_25463,N_25108);
and UO_1328 (O_1328,N_29881,N_25600);
or UO_1329 (O_1329,N_28112,N_27638);
or UO_1330 (O_1330,N_28179,N_29530);
or UO_1331 (O_1331,N_27917,N_25100);
or UO_1332 (O_1332,N_28486,N_25344);
or UO_1333 (O_1333,N_28661,N_27112);
or UO_1334 (O_1334,N_27292,N_27735);
nand UO_1335 (O_1335,N_26774,N_27421);
and UO_1336 (O_1336,N_25267,N_25420);
nand UO_1337 (O_1337,N_28808,N_27093);
xnor UO_1338 (O_1338,N_29833,N_29815);
nor UO_1339 (O_1339,N_25444,N_28952);
xor UO_1340 (O_1340,N_27709,N_27940);
nor UO_1341 (O_1341,N_25613,N_26473);
xnor UO_1342 (O_1342,N_25387,N_25929);
xor UO_1343 (O_1343,N_27194,N_27279);
or UO_1344 (O_1344,N_25534,N_29786);
nor UO_1345 (O_1345,N_26898,N_26349);
xnor UO_1346 (O_1346,N_28245,N_27597);
nor UO_1347 (O_1347,N_29724,N_27083);
and UO_1348 (O_1348,N_26385,N_25823);
nand UO_1349 (O_1349,N_28093,N_25758);
and UO_1350 (O_1350,N_26577,N_28683);
and UO_1351 (O_1351,N_27234,N_29192);
nor UO_1352 (O_1352,N_26962,N_26558);
nand UO_1353 (O_1353,N_26879,N_29741);
and UO_1354 (O_1354,N_27797,N_25612);
nor UO_1355 (O_1355,N_25917,N_26536);
xor UO_1356 (O_1356,N_26246,N_27997);
and UO_1357 (O_1357,N_28185,N_29215);
nand UO_1358 (O_1358,N_25617,N_28630);
or UO_1359 (O_1359,N_29517,N_27818);
xor UO_1360 (O_1360,N_25247,N_28182);
xor UO_1361 (O_1361,N_26960,N_25572);
or UO_1362 (O_1362,N_28484,N_25511);
nand UO_1363 (O_1363,N_25153,N_26003);
nand UO_1364 (O_1364,N_29277,N_29610);
xor UO_1365 (O_1365,N_28342,N_25546);
xor UO_1366 (O_1366,N_28733,N_27313);
and UO_1367 (O_1367,N_27409,N_25794);
or UO_1368 (O_1368,N_27402,N_29475);
and UO_1369 (O_1369,N_29597,N_28228);
xor UO_1370 (O_1370,N_28862,N_25261);
xor UO_1371 (O_1371,N_28002,N_26595);
xnor UO_1372 (O_1372,N_29599,N_27708);
and UO_1373 (O_1373,N_29534,N_25544);
nor UO_1374 (O_1374,N_28844,N_28849);
or UO_1375 (O_1375,N_26154,N_26615);
nand UO_1376 (O_1376,N_26516,N_28958);
xnor UO_1377 (O_1377,N_27732,N_26322);
xnor UO_1378 (O_1378,N_26370,N_27875);
xor UO_1379 (O_1379,N_25133,N_25770);
nand UO_1380 (O_1380,N_25291,N_29860);
or UO_1381 (O_1381,N_28369,N_29970);
nor UO_1382 (O_1382,N_25378,N_28850);
nor UO_1383 (O_1383,N_26724,N_27792);
xnor UO_1384 (O_1384,N_25250,N_29694);
or UO_1385 (O_1385,N_25389,N_27434);
nand UO_1386 (O_1386,N_29880,N_25213);
or UO_1387 (O_1387,N_28525,N_25230);
xor UO_1388 (O_1388,N_29656,N_25533);
nor UO_1389 (O_1389,N_28749,N_25329);
nand UO_1390 (O_1390,N_28337,N_27188);
and UO_1391 (O_1391,N_26464,N_29055);
or UO_1392 (O_1392,N_28668,N_29094);
nor UO_1393 (O_1393,N_25539,N_29266);
nand UO_1394 (O_1394,N_27496,N_29638);
or UO_1395 (O_1395,N_25269,N_28237);
and UO_1396 (O_1396,N_26474,N_26891);
nand UO_1397 (O_1397,N_26199,N_27881);
or UO_1398 (O_1398,N_29566,N_27334);
and UO_1399 (O_1399,N_28203,N_26004);
nand UO_1400 (O_1400,N_25548,N_28919);
nand UO_1401 (O_1401,N_27860,N_28265);
or UO_1402 (O_1402,N_28795,N_28349);
and UO_1403 (O_1403,N_28856,N_28405);
and UO_1404 (O_1404,N_29299,N_25872);
or UO_1405 (O_1405,N_26064,N_28611);
and UO_1406 (O_1406,N_27247,N_28037);
and UO_1407 (O_1407,N_28577,N_29564);
and UO_1408 (O_1408,N_25677,N_28956);
nand UO_1409 (O_1409,N_28308,N_26071);
nor UO_1410 (O_1410,N_29930,N_28103);
or UO_1411 (O_1411,N_26754,N_28284);
xor UO_1412 (O_1412,N_27588,N_26510);
nor UO_1413 (O_1413,N_25980,N_28117);
xor UO_1414 (O_1414,N_25750,N_25633);
nor UO_1415 (O_1415,N_28163,N_25227);
nand UO_1416 (O_1416,N_25020,N_29152);
nor UO_1417 (O_1417,N_27737,N_29478);
xnor UO_1418 (O_1418,N_29540,N_27581);
nand UO_1419 (O_1419,N_27225,N_28920);
or UO_1420 (O_1420,N_28090,N_29796);
and UO_1421 (O_1421,N_29054,N_28578);
and UO_1422 (O_1422,N_25956,N_25806);
and UO_1423 (O_1423,N_27948,N_25125);
nand UO_1424 (O_1424,N_25386,N_26812);
nor UO_1425 (O_1425,N_29620,N_28628);
xnor UO_1426 (O_1426,N_25048,N_25316);
xor UO_1427 (O_1427,N_27359,N_29126);
or UO_1428 (O_1428,N_27647,N_25978);
nor UO_1429 (O_1429,N_25336,N_27572);
xnor UO_1430 (O_1430,N_29680,N_28438);
and UO_1431 (O_1431,N_25274,N_29864);
nor UO_1432 (O_1432,N_27377,N_28917);
xor UO_1433 (O_1433,N_28825,N_28930);
nand UO_1434 (O_1434,N_26770,N_27757);
nor UO_1435 (O_1435,N_29308,N_25045);
and UO_1436 (O_1436,N_27423,N_26013);
nor UO_1437 (O_1437,N_28588,N_29187);
nand UO_1438 (O_1438,N_29131,N_25121);
nand UO_1439 (O_1439,N_27503,N_27542);
or UO_1440 (O_1440,N_26643,N_28648);
nand UO_1441 (O_1441,N_25576,N_27780);
nor UO_1442 (O_1442,N_26341,N_27970);
nand UO_1443 (O_1443,N_29869,N_28761);
xor UO_1444 (O_1444,N_28780,N_26247);
or UO_1445 (O_1445,N_29675,N_27443);
nor UO_1446 (O_1446,N_26333,N_26658);
xor UO_1447 (O_1447,N_25687,N_29186);
nand UO_1448 (O_1448,N_27541,N_28370);
xor UO_1449 (O_1449,N_25272,N_25062);
or UO_1450 (O_1450,N_28690,N_26620);
xnor UO_1451 (O_1451,N_29252,N_27534);
and UO_1452 (O_1452,N_29779,N_25290);
nand UO_1453 (O_1453,N_27903,N_27812);
and UO_1454 (O_1454,N_25002,N_26767);
or UO_1455 (O_1455,N_28246,N_28942);
nor UO_1456 (O_1456,N_27624,N_26151);
and UO_1457 (O_1457,N_27181,N_26429);
nor UO_1458 (O_1458,N_25547,N_25309);
or UO_1459 (O_1459,N_25356,N_28618);
nand UO_1460 (O_1460,N_26908,N_28707);
nand UO_1461 (O_1461,N_26016,N_27795);
or UO_1462 (O_1462,N_25433,N_29057);
and UO_1463 (O_1463,N_26743,N_26326);
xnor UO_1464 (O_1464,N_29918,N_26695);
nor UO_1465 (O_1465,N_28089,N_29420);
and UO_1466 (O_1466,N_25237,N_29742);
or UO_1467 (O_1467,N_25218,N_26410);
xor UO_1468 (O_1468,N_26638,N_29710);
nand UO_1469 (O_1469,N_26067,N_28472);
nor UO_1470 (O_1470,N_27189,N_28984);
nor UO_1471 (O_1471,N_27277,N_27756);
or UO_1472 (O_1472,N_27404,N_26825);
or UO_1473 (O_1473,N_29164,N_29810);
nand UO_1474 (O_1474,N_26061,N_25186);
nand UO_1475 (O_1475,N_28094,N_26206);
xor UO_1476 (O_1476,N_26499,N_28121);
or UO_1477 (O_1477,N_29518,N_28932);
and UO_1478 (O_1478,N_28184,N_27186);
nor UO_1479 (O_1479,N_27653,N_29255);
nor UO_1480 (O_1480,N_29855,N_27546);
nand UO_1481 (O_1481,N_29485,N_26555);
and UO_1482 (O_1482,N_26785,N_28026);
or UO_1483 (O_1483,N_26149,N_27172);
or UO_1484 (O_1484,N_28892,N_25555);
or UO_1485 (O_1485,N_27509,N_29195);
or UO_1486 (O_1486,N_26876,N_27711);
and UO_1487 (O_1487,N_25686,N_29916);
xor UO_1488 (O_1488,N_27494,N_28055);
nor UO_1489 (O_1489,N_28400,N_27544);
xor UO_1490 (O_1490,N_26806,N_26987);
and UO_1491 (O_1491,N_27811,N_25742);
nor UO_1492 (O_1492,N_25151,N_28295);
nor UO_1493 (O_1493,N_28614,N_27596);
nor UO_1494 (O_1494,N_25529,N_25043);
xnor UO_1495 (O_1495,N_25972,N_29549);
or UO_1496 (O_1496,N_29406,N_25642);
nand UO_1497 (O_1497,N_26072,N_25781);
xor UO_1498 (O_1498,N_25882,N_28126);
or UO_1499 (O_1499,N_25180,N_25936);
or UO_1500 (O_1500,N_26736,N_26108);
nand UO_1501 (O_1501,N_27243,N_29359);
or UO_1502 (O_1502,N_28526,N_25114);
and UO_1503 (O_1503,N_28140,N_27024);
nor UO_1504 (O_1504,N_29882,N_26147);
and UO_1505 (O_1505,N_25466,N_25333);
and UO_1506 (O_1506,N_26352,N_29745);
or UO_1507 (O_1507,N_27923,N_28345);
or UO_1508 (O_1508,N_28792,N_25659);
and UO_1509 (O_1509,N_25525,N_26557);
and UO_1510 (O_1510,N_28233,N_26896);
nand UO_1511 (O_1511,N_25339,N_28512);
and UO_1512 (O_1512,N_25483,N_26441);
nand UO_1513 (O_1513,N_27146,N_28323);
xnor UO_1514 (O_1514,N_26271,N_28452);
nor UO_1515 (O_1515,N_28178,N_29426);
and UO_1516 (O_1516,N_25545,N_25295);
xnor UO_1517 (O_1517,N_28098,N_27571);
and UO_1518 (O_1518,N_28759,N_29380);
xnor UO_1519 (O_1519,N_26665,N_26220);
xnor UO_1520 (O_1520,N_26853,N_25452);
nor UO_1521 (O_1521,N_26262,N_25646);
xor UO_1522 (O_1522,N_26308,N_28972);
nor UO_1523 (O_1523,N_25891,N_26229);
or UO_1524 (O_1524,N_26080,N_26484);
and UO_1525 (O_1525,N_26180,N_29954);
or UO_1526 (O_1526,N_29305,N_26762);
xor UO_1527 (O_1527,N_28200,N_26691);
nor UO_1528 (O_1528,N_27612,N_27978);
xnor UO_1529 (O_1529,N_28650,N_29590);
or UO_1530 (O_1530,N_27994,N_28716);
or UO_1531 (O_1531,N_29773,N_26201);
nand UO_1532 (O_1532,N_28896,N_26394);
nor UO_1533 (O_1533,N_28186,N_27213);
nand UO_1534 (O_1534,N_28839,N_27200);
and UO_1535 (O_1535,N_25725,N_28542);
nor UO_1536 (O_1536,N_29058,N_27702);
nor UO_1537 (O_1537,N_27878,N_29923);
or UO_1538 (O_1538,N_28969,N_29674);
nor UO_1539 (O_1539,N_29653,N_29121);
xnor UO_1540 (O_1540,N_28100,N_26143);
xnor UO_1541 (O_1541,N_27470,N_27627);
or UO_1542 (O_1542,N_25853,N_27865);
nor UO_1543 (O_1543,N_29931,N_28974);
nor UO_1544 (O_1544,N_28318,N_29492);
or UO_1545 (O_1545,N_25438,N_28007);
nand UO_1546 (O_1546,N_29617,N_28814);
and UO_1547 (O_1547,N_25374,N_29038);
nand UO_1548 (O_1548,N_27025,N_25638);
nand UO_1549 (O_1549,N_27383,N_28389);
nor UO_1550 (O_1550,N_27054,N_26855);
xor UO_1551 (O_1551,N_27984,N_29232);
xnor UO_1552 (O_1552,N_29781,N_25442);
xnor UO_1553 (O_1553,N_28558,N_28522);
or UO_1554 (O_1554,N_28373,N_29271);
nand UO_1555 (O_1555,N_27913,N_25795);
or UO_1556 (O_1556,N_29374,N_26272);
xor UO_1557 (O_1557,N_29525,N_29991);
nor UO_1558 (O_1558,N_29129,N_27269);
nor UO_1559 (O_1559,N_29463,N_29151);
nand UO_1560 (O_1560,N_28466,N_27972);
xor UO_1561 (O_1561,N_29468,N_25223);
nand UO_1562 (O_1562,N_27275,N_28439);
nand UO_1563 (O_1563,N_25727,N_29224);
xor UO_1564 (O_1564,N_27980,N_28569);
and UO_1565 (O_1565,N_27429,N_25152);
xor UO_1566 (O_1566,N_27774,N_25044);
xor UO_1567 (O_1567,N_25945,N_28517);
xor UO_1568 (O_1568,N_28076,N_27791);
nor UO_1569 (O_1569,N_27976,N_27759);
nor UO_1570 (O_1570,N_29403,N_28225);
nor UO_1571 (O_1571,N_25595,N_27531);
nor UO_1572 (O_1572,N_25556,N_29011);
nor UO_1573 (O_1573,N_26950,N_29008);
xor UO_1574 (O_1574,N_28181,N_28793);
or UO_1575 (O_1575,N_25464,N_28736);
or UO_1576 (O_1576,N_27022,N_26010);
nor UO_1577 (O_1577,N_27163,N_26678);
xor UO_1578 (O_1578,N_26282,N_26599);
and UO_1579 (O_1579,N_28330,N_26416);
nor UO_1580 (O_1580,N_29063,N_25183);
nand UO_1581 (O_1581,N_28686,N_27555);
xnor UO_1582 (O_1582,N_28430,N_27789);
nor UO_1583 (O_1583,N_28396,N_25169);
nor UO_1584 (O_1584,N_25959,N_26050);
nand UO_1585 (O_1585,N_27736,N_28446);
or UO_1586 (O_1586,N_28879,N_26221);
nand UO_1587 (O_1587,N_25177,N_28445);
or UO_1588 (O_1588,N_27246,N_26968);
xnor UO_1589 (O_1589,N_27038,N_25004);
nand UO_1590 (O_1590,N_26171,N_28003);
nor UO_1591 (O_1591,N_25604,N_27424);
nand UO_1592 (O_1592,N_25715,N_26249);
or UO_1593 (O_1593,N_28460,N_26146);
or UO_1594 (O_1594,N_25053,N_25907);
xnor UO_1595 (O_1595,N_26092,N_29943);
or UO_1596 (O_1596,N_25319,N_26870);
nor UO_1597 (O_1597,N_28924,N_29024);
xnor UO_1598 (O_1598,N_27249,N_25251);
and UO_1599 (O_1599,N_27664,N_29666);
nor UO_1600 (O_1600,N_27642,N_27134);
or UO_1601 (O_1601,N_29265,N_28976);
xor UO_1602 (O_1602,N_28384,N_29613);
nor UO_1603 (O_1603,N_28432,N_29820);
xor UO_1604 (O_1604,N_28355,N_25468);
or UO_1605 (O_1605,N_29035,N_28902);
nor UO_1606 (O_1606,N_27064,N_26992);
xor UO_1607 (O_1607,N_26722,N_25154);
xnor UO_1608 (O_1608,N_28973,N_27016);
and UO_1609 (O_1609,N_28280,N_27842);
nand UO_1610 (O_1610,N_26920,N_28638);
nor UO_1611 (O_1611,N_28665,N_26167);
or UO_1612 (O_1612,N_26043,N_28394);
nand UO_1613 (O_1613,N_27777,N_27944);
or UO_1614 (O_1614,N_25876,N_29112);
nand UO_1615 (O_1615,N_28042,N_28743);
nor UO_1616 (O_1616,N_26481,N_28060);
xor UO_1617 (O_1617,N_27979,N_25080);
nor UO_1618 (O_1618,N_25402,N_27915);
nor UO_1619 (O_1619,N_28983,N_26598);
nor UO_1620 (O_1620,N_25862,N_29681);
nor UO_1621 (O_1621,N_25134,N_25171);
or UO_1622 (O_1622,N_26468,N_27559);
nand UO_1623 (O_1623,N_29072,N_29175);
or UO_1624 (O_1624,N_26436,N_28207);
and UO_1625 (O_1625,N_27570,N_29120);
nor UO_1626 (O_1626,N_27489,N_28238);
nand UO_1627 (O_1627,N_28947,N_28821);
or UO_1628 (O_1628,N_27931,N_29474);
xor UO_1629 (O_1629,N_27133,N_26421);
nand UO_1630 (O_1630,N_27347,N_25111);
and UO_1631 (O_1631,N_26553,N_25928);
nand UO_1632 (O_1632,N_25405,N_26716);
nand UO_1633 (O_1633,N_27783,N_27543);
xor UO_1634 (O_1634,N_26365,N_29047);
xnor UO_1635 (O_1635,N_26174,N_27855);
and UO_1636 (O_1636,N_29003,N_25288);
or UO_1637 (O_1637,N_25675,N_28546);
xor UO_1638 (O_1638,N_28109,N_25453);
xnor UO_1639 (O_1639,N_28338,N_27945);
and UO_1640 (O_1640,N_29137,N_29835);
xor UO_1641 (O_1641,N_27471,N_28467);
xor UO_1642 (O_1642,N_29922,N_26997);
xor UO_1643 (O_1643,N_28174,N_27632);
nand UO_1644 (O_1644,N_26024,N_29285);
xnor UO_1645 (O_1645,N_29395,N_29030);
xor UO_1646 (O_1646,N_28142,N_27501);
nor UO_1647 (O_1647,N_29807,N_26779);
or UO_1648 (O_1648,N_29375,N_25664);
and UO_1649 (O_1649,N_26245,N_28565);
and UO_1650 (O_1650,N_29967,N_29739);
nor UO_1651 (O_1651,N_28895,N_28751);
nand UO_1652 (O_1652,N_29033,N_27692);
or UO_1653 (O_1653,N_27148,N_25005);
and UO_1654 (O_1654,N_29091,N_28327);
or UO_1655 (O_1655,N_28393,N_26323);
nand UO_1656 (O_1656,N_25531,N_29201);
nand UO_1657 (O_1657,N_29611,N_27461);
or UO_1658 (O_1658,N_29222,N_27210);
nand UO_1659 (O_1659,N_29851,N_29366);
xor UO_1660 (O_1660,N_25065,N_28829);
xnor UO_1661 (O_1661,N_26097,N_26677);
xor UO_1662 (O_1662,N_26933,N_28101);
xor UO_1663 (O_1663,N_27192,N_26849);
xor UO_1664 (O_1664,N_28070,N_27465);
nor UO_1665 (O_1665,N_27989,N_25927);
or UO_1666 (O_1666,N_27908,N_25206);
or UO_1667 (O_1667,N_25049,N_26120);
nor UO_1668 (O_1668,N_29953,N_29572);
and UO_1669 (O_1669,N_27775,N_28025);
or UO_1670 (O_1670,N_27548,N_28532);
or UO_1671 (O_1671,N_28732,N_27033);
nor UO_1672 (O_1672,N_28590,N_28421);
nand UO_1673 (O_1673,N_29401,N_28334);
nor UO_1674 (O_1674,N_26963,N_25904);
and UO_1675 (O_1675,N_29337,N_29797);
or UO_1676 (O_1676,N_26753,N_29736);
nor UO_1677 (O_1677,N_27170,N_28281);
nand UO_1678 (O_1678,N_28811,N_26228);
nand UO_1679 (O_1679,N_27262,N_28417);
xnor UO_1680 (O_1680,N_28901,N_26542);
nand UO_1681 (O_1681,N_29988,N_29732);
xor UO_1682 (O_1682,N_27061,N_28781);
and UO_1683 (O_1683,N_25110,N_25578);
or UO_1684 (O_1684,N_25637,N_28933);
or UO_1685 (O_1685,N_27329,N_27203);
xor UO_1686 (O_1686,N_27633,N_27099);
nor UO_1687 (O_1687,N_27943,N_26580);
nand UO_1688 (O_1688,N_26921,N_29069);
nand UO_1689 (O_1689,N_25857,N_29960);
xnor UO_1690 (O_1690,N_26492,N_26871);
nand UO_1691 (O_1691,N_28303,N_25608);
nor UO_1692 (O_1692,N_27378,N_26965);
nand UO_1693 (O_1693,N_25530,N_29105);
xor UO_1694 (O_1694,N_28480,N_26803);
or UO_1695 (O_1695,N_28435,N_26396);
nand UO_1696 (O_1696,N_25732,N_26019);
nor UO_1697 (O_1697,N_26972,N_29087);
and UO_1698 (O_1698,N_25212,N_26687);
nand UO_1699 (O_1699,N_25447,N_25992);
nand UO_1700 (O_1700,N_29986,N_28108);
or UO_1701 (O_1701,N_26834,N_26106);
nor UO_1702 (O_1702,N_27417,N_25704);
nand UO_1703 (O_1703,N_29336,N_29480);
nor UO_1704 (O_1704,N_26520,N_28696);
nand UO_1705 (O_1705,N_28087,N_26938);
xor UO_1706 (O_1706,N_28595,N_25306);
nor UO_1707 (O_1707,N_28262,N_25510);
nor UO_1708 (O_1708,N_29720,N_27450);
nand UO_1709 (O_1709,N_29502,N_27828);
xnor UO_1710 (O_1710,N_28276,N_25450);
or UO_1711 (O_1711,N_28572,N_29721);
and UO_1712 (O_1712,N_29496,N_28211);
xnor UO_1713 (O_1713,N_27492,N_26107);
nor UO_1714 (O_1714,N_26901,N_27460);
xnor UO_1715 (O_1715,N_28271,N_28214);
xnor UO_1716 (O_1716,N_27803,N_28894);
nor UO_1717 (O_1717,N_27447,N_28635);
xnor UO_1718 (O_1718,N_27731,N_27272);
or UO_1719 (O_1719,N_25275,N_29189);
nand UO_1720 (O_1720,N_28378,N_25759);
xnor UO_1721 (O_1721,N_28819,N_29109);
nor UO_1722 (O_1722,N_26320,N_25523);
nor UO_1723 (O_1723,N_26292,N_29219);
and UO_1724 (O_1724,N_25495,N_27293);
and UO_1725 (O_1725,N_25164,N_29498);
nor UO_1726 (O_1726,N_27933,N_26729);
and UO_1727 (O_1727,N_26742,N_27182);
nand UO_1728 (O_1728,N_26690,N_28032);
xnor UO_1729 (O_1729,N_26039,N_25821);
and UO_1730 (O_1730,N_29434,N_28092);
nor UO_1731 (O_1731,N_27077,N_25962);
and UO_1732 (O_1732,N_25564,N_27700);
and UO_1733 (O_1733,N_26862,N_25139);
or UO_1734 (O_1734,N_26233,N_25026);
xor UO_1735 (O_1735,N_27425,N_26079);
nor UO_1736 (O_1736,N_27078,N_27804);
and UO_1737 (O_1737,N_26243,N_25657);
and UO_1738 (O_1738,N_27714,N_25703);
and UO_1739 (O_1739,N_25265,N_29268);
nand UO_1740 (O_1740,N_26148,N_28234);
and UO_1741 (O_1741,N_25410,N_28533);
nor UO_1742 (O_1742,N_29911,N_29557);
nand UO_1743 (O_1743,N_27231,N_26828);
nand UO_1744 (O_1744,N_25294,N_28680);
or UO_1745 (O_1745,N_26588,N_26306);
nor UO_1746 (O_1746,N_26749,N_29074);
and UO_1747 (O_1747,N_28679,N_27196);
nand UO_1748 (O_1748,N_25255,N_27049);
nand UO_1749 (O_1749,N_25013,N_29995);
xor UO_1750 (O_1750,N_25737,N_27663);
nor UO_1751 (O_1751,N_29104,N_29451);
or UO_1752 (O_1752,N_25537,N_25457);
and UO_1753 (O_1753,N_27169,N_27563);
nor UO_1754 (O_1754,N_29684,N_29816);
xor UO_1755 (O_1755,N_28529,N_26406);
nand UO_1756 (O_1756,N_28677,N_25824);
nand UO_1757 (O_1757,N_26763,N_27310);
xnor UO_1758 (O_1758,N_29162,N_25390);
and UO_1759 (O_1759,N_28998,N_28441);
or UO_1760 (O_1760,N_25867,N_28547);
and UO_1761 (O_1761,N_27906,N_27464);
nand UO_1762 (O_1762,N_26230,N_27075);
or UO_1763 (O_1763,N_25615,N_26126);
and UO_1764 (O_1764,N_27493,N_29890);
xor UO_1765 (O_1765,N_25752,N_29888);
xor UO_1766 (O_1766,N_25092,N_25663);
or UO_1767 (O_1767,N_25797,N_28130);
nand UO_1768 (O_1768,N_27790,N_28379);
xnor UO_1769 (O_1769,N_29119,N_26415);
and UO_1770 (O_1770,N_29800,N_27029);
nand UO_1771 (O_1771,N_26505,N_28354);
nand UO_1772 (O_1772,N_29070,N_29416);
xor UO_1773 (O_1773,N_26693,N_28453);
nand UO_1774 (O_1774,N_25372,N_29041);
xnor UO_1775 (O_1775,N_25025,N_25370);
or UO_1776 (O_1776,N_25143,N_28797);
or UO_1777 (O_1777,N_29470,N_26961);
xnor UO_1778 (O_1778,N_28609,N_29172);
nand UO_1779 (O_1779,N_27481,N_28124);
nand UO_1780 (O_1780,N_27727,N_25722);
nand UO_1781 (O_1781,N_27239,N_28104);
xor UO_1782 (O_1782,N_29067,N_25517);
xnor UO_1783 (O_1783,N_27237,N_27959);
or UO_1784 (O_1784,N_27776,N_28991);
and UO_1785 (O_1785,N_28964,N_27982);
nand UO_1786 (O_1786,N_28812,N_26578);
xor UO_1787 (O_1787,N_28286,N_27168);
and UO_1788 (O_1788,N_27426,N_25244);
or UO_1789 (O_1789,N_27151,N_25925);
nand UO_1790 (O_1790,N_25938,N_27498);
xor UO_1791 (O_1791,N_25575,N_25661);
nor UO_1792 (O_1792,N_28596,N_28504);
xor UO_1793 (O_1793,N_26411,N_28560);
xnor UO_1794 (O_1794,N_25131,N_28317);
nor UO_1795 (O_1795,N_26357,N_27248);
or UO_1796 (O_1796,N_28336,N_28065);
or UO_1797 (O_1797,N_26094,N_26903);
nand UO_1798 (O_1798,N_27766,N_28051);
or UO_1799 (O_1799,N_28603,N_25489);
nand UO_1800 (O_1800,N_28535,N_28455);
and UO_1801 (O_1801,N_29431,N_26854);
or UO_1802 (O_1802,N_29897,N_25954);
and UO_1803 (O_1803,N_27135,N_28520);
xor UO_1804 (O_1804,N_25889,N_29623);
or UO_1805 (O_1805,N_27675,N_29254);
and UO_1806 (O_1806,N_28842,N_25754);
or UO_1807 (O_1807,N_25322,N_28503);
or UO_1808 (O_1808,N_27887,N_27829);
and UO_1809 (O_1809,N_28887,N_26086);
and UO_1810 (O_1810,N_29220,N_29553);
nand UO_1811 (O_1811,N_29383,N_28699);
nand UO_1812 (O_1812,N_27397,N_26579);
xnor UO_1813 (O_1813,N_27583,N_29140);
or UO_1814 (O_1814,N_25800,N_25943);
or UO_1815 (O_1815,N_25017,N_28078);
nor UO_1816 (O_1816,N_28072,N_28953);
nand UO_1817 (O_1817,N_25714,N_29319);
nand UO_1818 (O_1818,N_29404,N_28311);
xnor UO_1819 (O_1819,N_29898,N_29278);
xnor UO_1820 (O_1820,N_27514,N_25921);
and UO_1821 (O_1821,N_27910,N_27554);
nand UO_1822 (O_1822,N_26880,N_28296);
and UO_1823 (O_1823,N_29301,N_26789);
xnor UO_1824 (O_1824,N_28785,N_27342);
nand UO_1825 (O_1825,N_29080,N_28148);
xor UO_1826 (O_1826,N_28053,N_29921);
nand UO_1827 (O_1827,N_28462,N_28269);
or UO_1828 (O_1828,N_26929,N_28975);
or UO_1829 (O_1829,N_26851,N_26178);
nand UO_1830 (O_1830,N_29197,N_27799);
nor UO_1831 (O_1831,N_26140,N_27882);
nand UO_1832 (O_1832,N_27384,N_29912);
nor UO_1833 (O_1833,N_28023,N_25411);
xnor UO_1834 (O_1834,N_26157,N_26569);
or UO_1835 (O_1835,N_27240,N_28871);
xnor UO_1836 (O_1836,N_26634,N_25095);
xnor UO_1837 (O_1837,N_27187,N_29438);
and UO_1838 (O_1838,N_27975,N_27057);
or UO_1839 (O_1839,N_29217,N_26035);
or UO_1840 (O_1840,N_29659,N_28554);
or UO_1841 (O_1841,N_27925,N_25362);
xor UO_1842 (O_1842,N_28307,N_29486);
nor UO_1843 (O_1843,N_29642,N_28476);
xnor UO_1844 (O_1844,N_29825,N_27238);
nor UO_1845 (O_1845,N_27361,N_29231);
and UO_1846 (O_1846,N_26809,N_25052);
and UO_1847 (O_1847,N_29904,N_25482);
and UO_1848 (O_1848,N_28168,N_28878);
nand UO_1849 (O_1849,N_29682,N_26522);
xor UO_1850 (O_1850,N_26235,N_25051);
or UO_1851 (O_1851,N_29634,N_27143);
and UO_1852 (O_1852,N_25838,N_28257);
nor UO_1853 (O_1853,N_27145,N_28013);
or UO_1854 (O_1854,N_28625,N_25172);
nor UO_1855 (O_1855,N_27174,N_28263);
xnor UO_1856 (O_1856,N_29324,N_27113);
and UO_1857 (O_1857,N_25484,N_26494);
xor UO_1858 (O_1858,N_28099,N_29841);
or UO_1859 (O_1859,N_25683,N_27992);
and UO_1860 (O_1860,N_25421,N_25023);
and UO_1861 (O_1861,N_26688,N_28266);
nor UO_1862 (O_1862,N_28592,N_28717);
and UO_1863 (O_1863,N_28247,N_29275);
nand UO_1864 (O_1864,N_26850,N_26560);
or UO_1865 (O_1865,N_29893,N_28944);
nand UO_1866 (O_1866,N_28038,N_27308);
xnor UO_1867 (O_1867,N_27059,N_29928);
nand UO_1868 (O_1868,N_28801,N_29329);
and UO_1869 (O_1869,N_28889,N_26635);
and UO_1870 (O_1870,N_29537,N_27366);
nor UO_1871 (O_1871,N_28636,N_25721);
and UO_1872 (O_1872,N_27056,N_27371);
nand UO_1873 (O_1873,N_26191,N_29934);
nor UO_1874 (O_1874,N_26957,N_29580);
xnor UO_1875 (O_1875,N_25785,N_27283);
and UO_1876 (O_1876,N_27525,N_27164);
nand UO_1877 (O_1877,N_28254,N_28170);
xor UO_1878 (O_1878,N_29889,N_28802);
xnor UO_1879 (O_1879,N_29289,N_27251);
nor UO_1880 (O_1880,N_25039,N_26273);
or UO_1881 (O_1881,N_29966,N_27066);
xor UO_1882 (O_1882,N_29331,N_25593);
nor UO_1883 (O_1883,N_28755,N_28054);
xor UO_1884 (O_1884,N_29850,N_25126);
nand UO_1885 (O_1885,N_29095,N_28629);
or UO_1886 (O_1886,N_26808,N_27226);
xnor UO_1887 (O_1887,N_29630,N_28457);
xor UO_1888 (O_1888,N_25969,N_26132);
and UO_1889 (O_1889,N_28141,N_26502);
xor UO_1890 (O_1890,N_25357,N_27579);
and UO_1891 (O_1891,N_28448,N_25653);
and UO_1892 (O_1892,N_28985,N_27939);
nand UO_1893 (O_1893,N_28670,N_26946);
nand UO_1894 (O_1894,N_29267,N_27929);
nand UO_1895 (O_1895,N_26379,N_28981);
xor UO_1896 (O_1896,N_26102,N_29990);
or UO_1897 (O_1897,N_26095,N_27119);
or UO_1898 (O_1898,N_29364,N_27950);
or UO_1899 (O_1899,N_29249,N_26715);
or UO_1900 (O_1900,N_29165,N_27388);
xor UO_1901 (O_1901,N_28791,N_29399);
xnor UO_1902 (O_1902,N_25669,N_27011);
nor UO_1903 (O_1903,N_27930,N_29452);
and UO_1904 (O_1904,N_25094,N_29049);
nand UO_1905 (O_1905,N_25535,N_26636);
and UO_1906 (O_1906,N_25501,N_27771);
nand UO_1907 (O_1907,N_26541,N_27734);
and UO_1908 (O_1908,N_26877,N_25989);
or UO_1909 (O_1909,N_28582,N_29143);
xor UO_1910 (O_1910,N_29349,N_27032);
nand UO_1911 (O_1911,N_27302,N_27769);
and UO_1912 (O_1912,N_28471,N_29497);
and UO_1913 (O_1913,N_27007,N_29972);
nand UO_1914 (O_1914,N_26036,N_29322);
nor UO_1915 (O_1915,N_27085,N_25341);
nor UO_1916 (O_1916,N_27137,N_29239);
nand UO_1917 (O_1917,N_27599,N_26810);
or UO_1918 (O_1918,N_27340,N_29649);
and UO_1919 (O_1919,N_27513,N_28274);
xnor UO_1920 (O_1920,N_25142,N_27967);
xor UO_1921 (O_1921,N_26631,N_29226);
nand UO_1922 (O_1922,N_27001,N_28726);
and UO_1923 (O_1923,N_29536,N_27127);
and UO_1924 (O_1924,N_28145,N_27105);
xor UO_1925 (O_1925,N_25783,N_27515);
or UO_1926 (O_1926,N_29161,N_26840);
nand UO_1927 (O_1927,N_28329,N_27983);
nor UO_1928 (O_1928,N_25198,N_27084);
nand UO_1929 (O_1929,N_27191,N_27900);
and UO_1930 (O_1930,N_27046,N_25490);
nand UO_1931 (O_1931,N_27607,N_27273);
xnor UO_1932 (O_1932,N_26760,N_28147);
nand UO_1933 (O_1933,N_28427,N_29483);
nand UO_1934 (O_1934,N_26121,N_29471);
nor UO_1935 (O_1935,N_27990,N_29963);
xor UO_1936 (O_1936,N_26070,N_25460);
and UO_1937 (O_1937,N_28563,N_26575);
nand UO_1938 (O_1938,N_25231,N_25763);
nand UO_1939 (O_1939,N_27339,N_27406);
and UO_1940 (O_1940,N_27080,N_27382);
and UO_1941 (O_1941,N_28097,N_26725);
and UO_1942 (O_1942,N_27398,N_28943);
nor UO_1943 (O_1943,N_27360,N_26367);
nand UO_1944 (O_1944,N_26652,N_26827);
and UO_1945 (O_1945,N_26787,N_27547);
xor UO_1946 (O_1946,N_26116,N_27745);
or UO_1947 (O_1947,N_25217,N_28586);
nor UO_1948 (O_1948,N_27026,N_28248);
nor UO_1949 (O_1949,N_25870,N_29764);
and UO_1950 (O_1950,N_25729,N_28723);
and UO_1951 (O_1951,N_27706,N_28552);
or UO_1952 (O_1952,N_26780,N_28157);
xnor UO_1953 (O_1953,N_28086,N_29949);
nand UO_1954 (O_1954,N_27753,N_26700);
or UO_1955 (O_1955,N_25504,N_29962);
nor UO_1956 (O_1956,N_27207,N_28992);
xnor UO_1957 (O_1957,N_25436,N_26601);
xnor UO_1958 (O_1958,N_26401,N_26731);
and UO_1959 (O_1959,N_27963,N_29801);
and UO_1960 (O_1960,N_26746,N_29330);
and UO_1961 (O_1961,N_29123,N_25423);
and UO_1962 (O_1962,N_26176,N_26648);
xor UO_1963 (O_1963,N_28299,N_25066);
xnor UO_1964 (O_1964,N_25395,N_25443);
and UO_1965 (O_1965,N_25611,N_25579);
or UO_1966 (O_1966,N_28409,N_26022);
nand UO_1967 (O_1967,N_26087,N_29533);
nand UO_1968 (O_1968,N_27183,N_25952);
or UO_1969 (O_1969,N_26772,N_25130);
nand UO_1970 (O_1970,N_25299,N_28443);
or UO_1971 (O_1971,N_27657,N_27045);
or UO_1972 (O_1972,N_27879,N_29282);
nor UO_1973 (O_1973,N_28660,N_27909);
xnor UO_1974 (O_1974,N_26625,N_29361);
and UO_1975 (O_1975,N_26540,N_29945);
nor UO_1976 (O_1976,N_28267,N_26456);
or UO_1977 (O_1977,N_25644,N_27773);
nor UO_1978 (O_1978,N_25393,N_26637);
xor UO_1979 (O_1979,N_25268,N_29711);
nor UO_1980 (O_1980,N_26337,N_25769);
xnor UO_1981 (O_1981,N_29834,N_26283);
and UO_1982 (O_1982,N_26941,N_26184);
or UO_1983 (O_1983,N_25191,N_29686);
nor UO_1984 (O_1984,N_28481,N_25190);
nand UO_1985 (O_1985,N_29792,N_29915);
nor UO_1986 (O_1986,N_25768,N_29321);
xor UO_1987 (O_1987,N_27333,N_27242);
nor UO_1988 (O_1988,N_29044,N_28622);
nand UO_1989 (O_1989,N_25705,N_27713);
and UO_1990 (O_1990,N_28132,N_26444);
nor UO_1991 (O_1991,N_28058,N_27157);
xnor UO_1992 (O_1992,N_27650,N_27255);
nor UO_1993 (O_1993,N_29388,N_29903);
or UO_1994 (O_1994,N_28528,N_29688);
or UO_1995 (O_1995,N_26366,N_29209);
or UO_1996 (O_1996,N_29593,N_28979);
nand UO_1997 (O_1997,N_29702,N_26347);
or UO_1998 (O_1998,N_25713,N_27793);
nor UO_1999 (O_1999,N_29511,N_27009);
and UO_2000 (O_2000,N_27688,N_29435);
nor UO_2001 (O_2001,N_26011,N_26209);
nor UO_2002 (O_2002,N_28221,N_27864);
nor UO_2003 (O_2003,N_26487,N_28494);
xnor UO_2004 (O_2004,N_26801,N_28727);
or UO_2005 (O_2005,N_27552,N_27809);
nor UO_2006 (O_2006,N_28357,N_28530);
nor UO_2007 (O_2007,N_25814,N_28960);
nor UO_2008 (O_2008,N_27479,N_28350);
xnor UO_2009 (O_2009,N_28352,N_26830);
and UO_2010 (O_2010,N_28675,N_26053);
nor UO_2011 (O_2011,N_25097,N_28371);
nand UO_2012 (O_2012,N_29824,N_26649);
xor UO_2013 (O_2013,N_27412,N_29937);
xnor UO_2014 (O_2014,N_28333,N_26624);
nand UO_2015 (O_2015,N_25350,N_29071);
nor UO_2016 (O_2016,N_26085,N_29018);
nand UO_2017 (O_2017,N_25079,N_26765);
xor UO_2018 (O_2018,N_26212,N_29513);
or UO_2019 (O_2019,N_29762,N_26745);
nand UO_2020 (O_2020,N_29370,N_25849);
and UO_2021 (O_2021,N_25494,N_28218);
nand UO_2022 (O_2022,N_27260,N_26574);
nor UO_2023 (O_2023,N_29823,N_27316);
and UO_2024 (O_2024,N_27796,N_28511);
nor UO_2025 (O_2025,N_27840,N_28137);
nand UO_2026 (O_2026,N_27764,N_27454);
nor UO_2027 (O_2027,N_29997,N_29382);
and UO_2028 (O_2028,N_28420,N_27286);
or UO_2029 (O_2029,N_25073,N_28581);
nor UO_2030 (O_2030,N_29614,N_25586);
and UO_2031 (O_2031,N_26977,N_29929);
xnor UO_2032 (O_2032,N_28273,N_27121);
xor UO_2033 (O_2033,N_27651,N_27674);
nor UO_2034 (O_2034,N_28877,N_27698);
nor UO_2035 (O_2035,N_27453,N_25123);
xor UO_2036 (O_2036,N_29615,N_25054);
nand UO_2037 (O_2037,N_28232,N_29102);
nor UO_2038 (O_2038,N_29479,N_27920);
and UO_2039 (O_2039,N_26512,N_27220);
nor UO_2040 (O_2040,N_27528,N_25924);
xor UO_2041 (O_2041,N_28945,N_28634);
nor UO_2042 (O_2042,N_26531,N_26993);
nand UO_2043 (O_2043,N_26675,N_25461);
and UO_2044 (O_2044,N_25607,N_27518);
nand UO_2045 (O_2045,N_25916,N_28046);
xnor UO_2046 (O_2046,N_25315,N_28066);
and UO_2047 (O_2047,N_25478,N_28167);
nand UO_2048 (O_2048,N_28893,N_25264);
or UO_2049 (O_2049,N_26335,N_27907);
nor UO_2050 (O_2050,N_28514,N_28020);
or UO_2051 (O_2051,N_26252,N_25343);
nor UO_2052 (O_2052,N_26495,N_28340);
nand UO_2053 (O_2053,N_29153,N_26887);
xor UO_2054 (O_2054,N_29064,N_29548);
or UO_2055 (O_2055,N_29315,N_25912);
or UO_2056 (O_2056,N_29984,N_25138);
nor UO_2057 (O_2057,N_26454,N_29632);
nor UO_2058 (O_2058,N_28612,N_29297);
nor UO_2059 (O_2059,N_26761,N_29514);
xor UO_2060 (O_2060,N_29279,N_29381);
nand UO_2061 (O_2061,N_27294,N_29034);
or UO_2062 (O_2062,N_29529,N_29122);
xor UO_2063 (O_2063,N_28539,N_29846);
nand UO_2064 (O_2064,N_25416,N_29176);
and UO_2065 (O_2065,N_27655,N_28288);
or UO_2066 (O_2066,N_27109,N_27566);
or UO_2067 (O_2067,N_28444,N_25182);
xnor UO_2068 (O_2068,N_29743,N_27858);
or UO_2069 (O_2069,N_26496,N_28259);
nor UO_2070 (O_2070,N_28911,N_25006);
and UO_2071 (O_2071,N_28860,N_29341);
or UO_2072 (O_2072,N_27530,N_28217);
or UO_2073 (O_2073,N_29325,N_29103);
or UO_2074 (O_2074,N_29696,N_28285);
or UO_2075 (O_2075,N_25107,N_26984);
and UO_2076 (O_2076,N_26103,N_29913);
and UO_2077 (O_2077,N_28188,N_27219);
nand UO_2078 (O_2078,N_27573,N_29061);
and UO_2079 (O_2079,N_29304,N_25701);
nand UO_2080 (O_2080,N_26506,N_25400);
nor UO_2081 (O_2081,N_25944,N_29545);
xnor UO_2082 (O_2082,N_26701,N_28165);
or UO_2083 (O_2083,N_27403,N_29379);
nor UO_2084 (O_2084,N_26208,N_26040);
xnor UO_2085 (O_2085,N_25060,N_29644);
nand UO_2086 (O_2086,N_25745,N_26863);
and UO_2087 (O_2087,N_27595,N_28963);
nand UO_2088 (O_2088,N_27535,N_27336);
nand UO_2089 (O_2089,N_27227,N_27381);
nor UO_2090 (O_2090,N_27393,N_29443);
nor UO_2091 (O_2091,N_27483,N_28474);
nor UO_2092 (O_2092,N_25202,N_26293);
nor UO_2093 (O_2093,N_25086,N_25831);
xor UO_2094 (O_2094,N_25476,N_29394);
xnor UO_2095 (O_2095,N_27089,N_26739);
nor UO_2096 (O_2096,N_28980,N_27389);
nand UO_2097 (O_2097,N_25132,N_29752);
and UO_2098 (O_2098,N_29798,N_25908);
nand UO_2099 (O_2099,N_28551,N_28843);
and UO_2100 (O_2100,N_26457,N_26027);
nor UO_2101 (O_2101,N_28339,N_28431);
nand UO_2102 (O_2102,N_26538,N_27888);
and UO_2103 (O_2103,N_26990,N_28735);
nor UO_2104 (O_2104,N_25965,N_29830);
nor UO_2105 (O_2105,N_27485,N_25280);
xnor UO_2106 (O_2106,N_26068,N_28929);
xor UO_2107 (O_2107,N_25627,N_26088);
and UO_2108 (O_2108,N_29242,N_25744);
or UO_2109 (O_2109,N_28936,N_25061);
and UO_2110 (O_2110,N_28516,N_28183);
and UO_2111 (O_2111,N_27582,N_28757);
xor UO_2112 (O_2112,N_27679,N_29014);
nor UO_2113 (O_2113,N_26859,N_25368);
or UO_2114 (O_2114,N_29313,N_29212);
and UO_2115 (O_2115,N_29311,N_27955);
nand UO_2116 (O_2116,N_26488,N_29048);
or UO_2117 (O_2117,N_29886,N_27861);
nor UO_2118 (O_2118,N_27765,N_25835);
xnor UO_2119 (O_2119,N_26657,N_25736);
xnor UO_2120 (O_2120,N_27824,N_26524);
nand UO_2121 (O_2121,N_27616,N_25225);
nor UO_2122 (O_2122,N_25585,N_25699);
or UO_2123 (O_2123,N_27848,N_29520);
nand UO_2124 (O_2124,N_27386,N_25068);
or UO_2125 (O_2125,N_26723,N_28855);
nor UO_2126 (O_2126,N_29973,N_28390);
or UO_2127 (O_2127,N_25174,N_25730);
xnor UO_2128 (O_2128,N_25351,N_26504);
or UO_2129 (O_2129,N_29184,N_28567);
and UO_2130 (O_2130,N_28449,N_25394);
and UO_2131 (O_2131,N_26640,N_26111);
nand UO_2132 (O_2132,N_27619,N_29142);
or UO_2133 (O_2133,N_28358,N_26452);
and UO_2134 (O_2134,N_28681,N_27087);
or UO_2135 (O_2135,N_27823,N_29010);
and UO_2136 (O_2136,N_26158,N_28744);
nor UO_2137 (O_2137,N_28041,N_25982);
and UO_2138 (O_2138,N_27718,N_29727);
xor UO_2139 (O_2139,N_28617,N_26756);
xnor UO_2140 (O_2140,N_25439,N_26236);
nor UO_2141 (O_2141,N_25396,N_25503);
and UO_2142 (O_2142,N_27041,N_27859);
nand UO_2143 (O_2143,N_29269,N_25679);
xor UO_2144 (O_2144,N_27866,N_27307);
or UO_2145 (O_2145,N_29455,N_27609);
and UO_2146 (O_2146,N_26958,N_28461);
nand UO_2147 (O_2147,N_25550,N_26679);
xnor UO_2148 (O_2148,N_29098,N_27355);
xor UO_2149 (O_2149,N_27446,N_29093);
nor UO_2150 (O_2150,N_27553,N_28704);
xor UO_2151 (O_2151,N_28152,N_28416);
nand UO_2152 (O_2152,N_25812,N_25222);
nand UO_2153 (O_2153,N_27205,N_26726);
and UO_2154 (O_2154,N_26098,N_29013);
and UO_2155 (O_2155,N_28074,N_29901);
xor UO_2156 (O_2156,N_29909,N_26258);
and UO_2157 (O_2157,N_29491,N_26299);
xor UO_2158 (O_2158,N_26866,N_28091);
nand UO_2159 (O_2159,N_28391,N_25762);
or UO_2160 (O_2160,N_25565,N_27010);
and UO_2161 (O_2161,N_26254,N_25200);
nor UO_2162 (O_2162,N_27202,N_27035);
or UO_2163 (O_2163,N_28377,N_26702);
or UO_2164 (O_2164,N_29544,N_25985);
nand UO_2165 (O_2165,N_27816,N_28343);
nand UO_2166 (O_2166,N_27257,N_29233);
xnor UO_2167 (O_2167,N_28740,N_29670);
nand UO_2168 (O_2168,N_29663,N_27729);
nand UO_2169 (O_2169,N_28651,N_29056);
xor UO_2170 (O_2170,N_28364,N_25419);
nand UO_2171 (O_2171,N_29461,N_26422);
xor UO_2172 (O_2172,N_26007,N_28027);
and UO_2173 (O_2173,N_26170,N_28841);
or UO_2174 (O_2174,N_29495,N_29377);
nor UO_2175 (O_2175,N_27671,N_28031);
nor UO_2176 (O_2176,N_29936,N_26752);
or UO_2177 (O_2177,N_28962,N_29531);
nor UO_2178 (O_2178,N_28918,N_28521);
and UO_2179 (O_2179,N_27952,N_28436);
nor UO_2180 (O_2180,N_25603,N_25012);
nor UO_2181 (O_2181,N_25561,N_25739);
or UO_2182 (O_2182,N_28561,N_29947);
nor UO_2183 (O_2183,N_25591,N_27676);
or UO_2184 (O_2184,N_25718,N_26325);
and UO_2185 (O_2185,N_26694,N_29999);
and UO_2186 (O_2186,N_26511,N_26056);
nor UO_2187 (O_2187,N_25327,N_26782);
nor UO_2188 (O_2188,N_28212,N_28189);
nor UO_2189 (O_2189,N_27574,N_26104);
nand UO_2190 (O_2190,N_26232,N_25232);
nor UO_2191 (O_2191,N_29355,N_27841);
nand UO_2192 (O_2192,N_26711,N_26630);
nand UO_2193 (O_2193,N_29466,N_29398);
xor UO_2194 (O_2194,N_27367,N_26974);
nand UO_2195 (O_2195,N_27034,N_29689);
nand UO_2196 (O_2196,N_29664,N_29857);
or UO_2197 (O_2197,N_28598,N_28128);
nand UO_2198 (O_2198,N_27236,N_28434);
and UO_2199 (O_2199,N_25424,N_27274);
or UO_2200 (O_2200,N_28272,N_26805);
xnor UO_2201 (O_2201,N_28169,N_26628);
xnor UO_2202 (O_2202,N_25898,N_28258);
nand UO_2203 (O_2203,N_27451,N_29228);
and UO_2204 (O_2204,N_25618,N_29234);
nor UO_2205 (O_2205,N_29190,N_27354);
nand UO_2206 (O_2206,N_26200,N_26062);
or UO_2207 (O_2207,N_25234,N_27911);
nor UO_2208 (O_2208,N_28626,N_25382);
nor UO_2209 (O_2209,N_25815,N_28837);
or UO_2210 (O_2210,N_27278,N_26113);
nor UO_2211 (O_2211,N_28001,N_26918);
nor UO_2212 (O_2212,N_27259,N_26573);
xor UO_2213 (O_2213,N_29758,N_27012);
nor UO_2214 (O_2214,N_27261,N_25599);
xor UO_2215 (O_2215,N_29174,N_26343);
or UO_2216 (O_2216,N_25997,N_28824);
nand UO_2217 (O_2217,N_29441,N_25413);
xnor UO_2218 (O_2218,N_26662,N_26978);
nor UO_2219 (O_2219,N_26651,N_25383);
nor UO_2220 (O_2220,N_28689,N_29211);
and UO_2221 (O_2221,N_29939,N_27928);
and UO_2222 (O_2222,N_29021,N_28875);
or UO_2223 (O_2223,N_26332,N_29661);
and UO_2224 (O_2224,N_29083,N_27562);
and UO_2225 (O_2225,N_27094,N_26211);
and UO_2226 (O_2226,N_25804,N_26277);
or UO_2227 (O_2227,N_29660,N_26223);
nor UO_2228 (O_2228,N_28968,N_26376);
nor UO_2229 (O_2229,N_29974,N_25470);
nor UO_2230 (O_2230,N_29369,N_26814);
or UO_2231 (O_2231,N_25270,N_25283);
nor UO_2232 (O_2232,N_26369,N_26556);
xor UO_2233 (O_2233,N_28510,N_28566);
xor UO_2234 (O_2234,N_29053,N_29425);
xnor UO_2235 (O_2235,N_28239,N_26355);
nand UO_2236 (O_2236,N_27199,N_25901);
or UO_2237 (O_2237,N_26509,N_26698);
nand UO_2238 (O_2238,N_26375,N_28210);
nor UO_2239 (O_2239,N_25734,N_27678);
and UO_2240 (O_2240,N_27730,N_29730);
nand UO_2241 (O_2241,N_29532,N_25716);
or UO_2242 (O_2242,N_26737,N_29515);
xnor UO_2243 (O_2243,N_26732,N_27867);
nor UO_2244 (O_2244,N_27996,N_27877);
nor UO_2245 (O_2245,N_29006,N_27964);
nand UO_2246 (O_2246,N_25538,N_25459);
nand UO_2247 (O_2247,N_25243,N_28235);
or UO_2248 (O_2248,N_25782,N_29347);
nor UO_2249 (O_2249,N_25070,N_25226);
nor UO_2250 (O_2250,N_26318,N_26203);
or UO_2251 (O_2251,N_29971,N_25296);
or UO_2252 (O_2252,N_28624,N_27779);
nand UO_2253 (O_2253,N_26647,N_27726);
nor UO_2254 (O_2254,N_26613,N_28429);
nand UO_2255 (O_2255,N_28028,N_27758);
nor UO_2256 (O_2256,N_25570,N_28758);
nor UO_2257 (O_2257,N_26583,N_29569);
nor UO_2258 (O_2258,N_26967,N_29113);
xnor UO_2259 (O_2259,N_28110,N_25083);
and UO_2260 (O_2260,N_25552,N_25082);
or UO_2261 (O_2261,N_29843,N_26708);
nor UO_2262 (O_2262,N_28815,N_28125);
xnor UO_2263 (O_2263,N_25801,N_29182);
or UO_2264 (O_2264,N_25030,N_27218);
or UO_2265 (O_2265,N_28164,N_25358);
or UO_2266 (O_2266,N_27995,N_25573);
nor UO_2267 (O_2267,N_28290,N_26952);
nor UO_2268 (O_2268,N_29571,N_28368);
nor UO_2269 (O_2269,N_26300,N_29453);
nor UO_2270 (O_2270,N_26794,N_27161);
nor UO_2271 (O_2271,N_27289,N_25458);
xor UO_2272 (O_2272,N_25042,N_26214);
or UO_2273 (O_2273,N_28213,N_29650);
or UO_2274 (O_2274,N_25440,N_26684);
or UO_2275 (O_2275,N_25071,N_27415);
xnor UO_2276 (O_2276,N_29238,N_26641);
xnor UO_2277 (O_2277,N_28659,N_29389);
nor UO_2278 (O_2278,N_26995,N_29612);
nor UO_2279 (O_2279,N_26671,N_27344);
or UO_2280 (O_2280,N_26359,N_28328);
nand UO_2281 (O_2281,N_28655,N_27004);
and UO_2282 (O_2282,N_29357,N_25430);
or UO_2283 (O_2283,N_29235,N_26405);
nand UO_2284 (O_2284,N_25808,N_29076);
and UO_2285 (O_2285,N_26517,N_29066);
xnor UO_2286 (O_2286,N_26821,N_27369);
nor UO_2287 (O_2287,N_26650,N_25037);
nand UO_2288 (O_2288,N_27223,N_27428);
nand UO_2289 (O_2289,N_28034,N_28838);
xnor UO_2290 (O_2290,N_25014,N_25813);
or UO_2291 (O_2291,N_27455,N_27337);
nor UO_2292 (O_2292,N_29258,N_28166);
nand UO_2293 (O_2293,N_27987,N_27408);
nor UO_2294 (O_2294,N_27390,N_25487);
xnor UO_2295 (O_2295,N_28322,N_26144);
or UO_2296 (O_2296,N_25512,N_27233);
or UO_2297 (O_2297,N_29596,N_26954);
nor UO_2298 (O_2298,N_27680,N_28876);
nand UO_2299 (O_2299,N_29037,N_27921);
nand UO_2300 (O_2300,N_29828,N_25574);
nor UO_2301 (O_2301,N_26525,N_29350);
xor UO_2302 (O_2302,N_27613,N_26041);
nand UO_2303 (O_2303,N_26561,N_27587);
xor UO_2304 (O_2304,N_26568,N_28208);
and UO_2305 (O_2305,N_26883,N_28788);
and UO_2306 (O_2306,N_28255,N_25141);
or UO_2307 (O_2307,N_27956,N_28642);
or UO_2308 (O_2308,N_27268,N_28627);
xor UO_2309 (O_2309,N_26440,N_28459);
nor UO_2310 (O_2310,N_25252,N_26593);
and UO_2311 (O_2311,N_29317,N_29029);
or UO_2312 (O_2312,N_25140,N_25676);
or UO_2313 (O_2313,N_25262,N_25209);
or UO_2314 (O_2314,N_26404,N_27744);
and UO_2315 (O_2315,N_27374,N_25967);
and UO_2316 (O_2316,N_29746,N_28029);
xnor UO_2317 (O_2317,N_29975,N_29567);
nand UO_2318 (O_2318,N_29601,N_29356);
nor UO_2319 (O_2319,N_28997,N_26720);
xnor UO_2320 (O_2320,N_27076,N_25465);
and UO_2321 (O_2321,N_29415,N_27565);
nand UO_2322 (O_2322,N_29547,N_26425);
nor UO_2323 (O_2323,N_29528,N_29678);
or UO_2324 (O_2324,N_26709,N_25589);
nand UO_2325 (O_2325,N_27522,N_29941);
and UO_2326 (O_2326,N_28599,N_28278);
xnor UO_2327 (O_2327,N_28063,N_27158);
nor UO_2328 (O_2328,N_25731,N_29367);
and UO_2329 (O_2329,N_29447,N_29718);
xor UO_2330 (O_2330,N_26438,N_25549);
and UO_2331 (O_2331,N_27993,N_28008);
nand UO_2332 (O_2332,N_27018,N_26181);
or UO_2333 (O_2333,N_25852,N_28700);
or UO_2334 (O_2334,N_27705,N_26037);
and UO_2335 (O_2335,N_26096,N_26482);
nor UO_2336 (O_2336,N_26009,N_29205);
and UO_2337 (O_2337,N_29107,N_26940);
and UO_2338 (O_2338,N_27873,N_26169);
nor UO_2339 (O_2339,N_27814,N_27195);
or UO_2340 (O_2340,N_25567,N_29940);
or UO_2341 (O_2341,N_25508,N_26476);
nor UO_2342 (O_2342,N_25774,N_25491);
nor UO_2343 (O_2343,N_28017,N_29981);
and UO_2344 (O_2344,N_26991,N_28498);
xor UO_2345 (O_2345,N_27585,N_25577);
nor UO_2346 (O_2346,N_26614,N_25865);
nor UO_2347 (O_2347,N_27854,N_27097);
nand UO_2348 (O_2348,N_26493,N_29460);
nand UO_2349 (O_2349,N_26572,N_25893);
nor UO_2350 (O_2350,N_25046,N_29062);
nor UO_2351 (O_2351,N_25673,N_28676);
nand UO_2352 (O_2352,N_27495,N_29734);
nor UO_2353 (O_2353,N_25103,N_28967);
nand UO_2354 (O_2354,N_29348,N_26286);
nor UO_2355 (O_2355,N_26738,N_29832);
xnor UO_2356 (O_2356,N_25279,N_25040);
and UO_2357 (O_2357,N_25619,N_27350);
and UO_2358 (O_2358,N_27872,N_27067);
and UO_2359 (O_2359,N_27512,N_26189);
xnor UO_2360 (O_2360,N_27600,N_26418);
nand UO_2361 (O_2361,N_27782,N_28602);
nand UO_2362 (O_2362,N_28693,N_28669);
or UO_2363 (O_2363,N_27296,N_28784);
or UO_2364 (O_2364,N_28912,N_27529);
nand UO_2365 (O_2365,N_28898,N_25330);
xnor UO_2366 (O_2366,N_28133,N_28865);
or UO_2367 (O_2367,N_25930,N_28196);
or UO_2368 (O_2368,N_28243,N_26998);
xor UO_2369 (O_2369,N_29865,N_27475);
nand UO_2370 (O_2370,N_25249,N_26769);
xor UO_2371 (O_2371,N_28083,N_29875);
or UO_2372 (O_2372,N_25672,N_26822);
and UO_2373 (O_2373,N_29695,N_26565);
nor UO_2374 (O_2374,N_26664,N_29402);
or UO_2375 (O_2375,N_29354,N_25314);
xnor UO_2376 (O_2376,N_26829,N_25205);
or UO_2377 (O_2377,N_29667,N_26465);
and UO_2378 (O_2378,N_28383,N_25032);
nand UO_2379 (O_2379,N_25662,N_29248);
xnor UO_2380 (O_2380,N_28115,N_28916);
nand UO_2381 (O_2381,N_28088,N_25195);
xor UO_2382 (O_2382,N_26559,N_28790);
or UO_2383 (O_2383,N_27605,N_28253);
nor UO_2384 (O_2384,N_27805,N_27165);
xor UO_2385 (O_2385,N_27122,N_27506);
or UO_2386 (O_2386,N_27802,N_28075);
nor UO_2387 (O_2387,N_25342,N_27462);
nand UO_2388 (O_2388,N_25635,N_27622);
or UO_2389 (O_2389,N_25196,N_26445);
nor UO_2390 (O_2390,N_25946,N_25456);
nand UO_2391 (O_2391,N_29134,N_25986);
xor UO_2392 (O_2392,N_27998,N_25532);
xor UO_2393 (O_2393,N_28398,N_28621);
nand UO_2394 (O_2394,N_29769,N_27717);
or UO_2395 (O_2395,N_25047,N_29432);
nand UO_2396 (O_2396,N_27290,N_25906);
or UO_2397 (O_2397,N_26964,N_28069);
or UO_2398 (O_2398,N_25219,N_28786);
or UO_2399 (O_2399,N_26477,N_28534);
xor UO_2400 (O_2400,N_27519,N_27580);
or UO_2401 (O_2401,N_28545,N_25170);
or UO_2402 (O_2402,N_29863,N_29111);
xnor UO_2403 (O_2403,N_26947,N_25293);
nor UO_2404 (O_2404,N_25970,N_29583);
and UO_2405 (O_2405,N_25310,N_28469);
and UO_2406 (O_2406,N_29621,N_26617);
nand UO_2407 (O_2407,N_28146,N_26437);
and UO_2408 (O_2408,N_27154,N_26608);
nor UO_2409 (O_2409,N_26969,N_29259);
or UO_2410 (O_2410,N_27924,N_25626);
nor UO_2411 (O_2411,N_25726,N_25144);
nand UO_2412 (O_2412,N_27439,N_29626);
nand UO_2413 (O_2413,N_29191,N_28544);
and UO_2414 (O_2414,N_29919,N_28220);
and UO_2415 (O_2415,N_27015,N_28884);
nor UO_2416 (O_2416,N_29429,N_28297);
nor UO_2417 (O_2417,N_29147,N_28994);
and UO_2418 (O_2418,N_27370,N_26434);
or UO_2419 (O_2419,N_29376,N_29658);
nor UO_2420 (O_2420,N_27282,N_25361);
nand UO_2421 (O_2421,N_27629,N_28646);
and UO_2422 (O_2422,N_28557,N_25772);
xnor UO_2423 (O_2423,N_26362,N_26747);
nand UO_2424 (O_2424,N_27241,N_27897);
or UO_2425 (O_2425,N_26645,N_25520);
or UO_2426 (O_2426,N_28241,N_28828);
nand UO_2427 (O_2427,N_29159,N_28789);
xnor UO_2428 (O_2428,N_29576,N_27898);
xor UO_2429 (O_2429,N_28151,N_27794);
or UO_2430 (O_2430,N_28502,N_29273);
and UO_2431 (O_2431,N_28414,N_29025);
or UO_2432 (O_2432,N_27288,N_27884);
or UO_2433 (O_2433,N_28600,N_25155);
or UO_2434 (O_2434,N_28509,N_25403);
xnor UO_2435 (O_2435,N_25473,N_27988);
nand UO_2436 (O_2436,N_29360,N_28230);
nor UO_2437 (O_2437,N_29951,N_26237);
and UO_2438 (O_2438,N_29877,N_26215);
or UO_2439 (O_2439,N_27149,N_26161);
or UO_2440 (O_2440,N_28367,N_29783);
xor UO_2441 (O_2441,N_25129,N_27166);
nor UO_2442 (O_2442,N_26856,N_25855);
nor UO_2443 (O_2443,N_29722,N_29551);
xnor UO_2444 (O_2444,N_29180,N_25960);
or UO_2445 (O_2445,N_26848,N_26423);
and UO_2446 (O_2446,N_28136,N_29296);
or UO_2447 (O_2447,N_29073,N_28139);
and UO_2448 (O_2448,N_29729,N_27966);
or UO_2449 (O_2449,N_28606,N_29917);
nor UO_2450 (O_2450,N_28143,N_27131);
nor UO_2451 (O_2451,N_29203,N_28982);
or UO_2452 (O_2452,N_25445,N_28989);
nand UO_2453 (O_2453,N_25951,N_29558);
or UO_2454 (O_2454,N_26259,N_27096);
nand UO_2455 (O_2455,N_29726,N_28999);
nor UO_2456 (O_2456,N_29039,N_28907);
xnor UO_2457 (O_2457,N_26290,N_27285);
nand UO_2458 (O_2458,N_29993,N_25427);
and UO_2459 (O_2459,N_28456,N_25958);
nor UO_2460 (O_2460,N_29908,N_26528);
and UO_2461 (O_2461,N_29392,N_27919);
xnor UO_2462 (O_2462,N_29158,N_26819);
nand UO_2463 (O_2463,N_25156,N_26692);
or UO_2464 (O_2464,N_29167,N_25493);
and UO_2465 (O_2465,N_29749,N_28499);
nand UO_2466 (O_2466,N_26554,N_28418);
and UO_2467 (O_2467,N_27845,N_26683);
or UO_2468 (O_2468,N_29352,N_29052);
xnor UO_2469 (O_2469,N_27474,N_28312);
nand UO_2470 (O_2470,N_26981,N_29789);
nor UO_2471 (O_2471,N_27436,N_29046);
nand UO_2472 (O_2472,N_27856,N_26547);
xor UO_2473 (O_2473,N_29647,N_26324);
or UO_2474 (O_2474,N_28085,N_28154);
nand UO_2475 (O_2475,N_26483,N_25707);
nor UO_2476 (O_2476,N_26587,N_25920);
nor UO_2477 (O_2477,N_27144,N_26642);
or UO_2478 (O_2478,N_29535,N_26837);
nor UO_2479 (O_2479,N_29760,N_26018);
nor UO_2480 (O_2480,N_27893,N_28922);
xor UO_2481 (O_2481,N_25777,N_29958);
and UO_2482 (O_2482,N_27748,N_28656);
nor UO_2483 (O_2483,N_28505,N_25780);
nor UO_2484 (O_2484,N_25875,N_25118);
nand UO_2485 (O_2485,N_28779,N_25880);
nand UO_2486 (O_2486,N_28044,N_25498);
and UO_2487 (O_2487,N_26906,N_28564);
nand UO_2488 (O_2488,N_26768,N_25911);
and UO_2489 (O_2489,N_26627,N_29559);
and UO_2490 (O_2490,N_27351,N_27376);
nand UO_2491 (O_2491,N_28921,N_27643);
xor UO_2492 (O_2492,N_28282,N_25939);
nor UO_2493 (O_2493,N_28882,N_28372);
xnor UO_2494 (O_2494,N_28988,N_27468);
or UO_2495 (O_2495,N_25632,N_28993);
xnor UO_2496 (O_2496,N_27179,N_25360);
and UO_2497 (O_2497,N_28950,N_25623);
or UO_2498 (O_2498,N_27747,N_28585);
and UO_2499 (O_2499,N_25301,N_28515);
xnor UO_2500 (O_2500,N_29300,N_27085);
nand UO_2501 (O_2501,N_26788,N_28555);
nand UO_2502 (O_2502,N_26228,N_27972);
or UO_2503 (O_2503,N_26038,N_25645);
xnor UO_2504 (O_2504,N_26136,N_26468);
or UO_2505 (O_2505,N_29874,N_29328);
or UO_2506 (O_2506,N_28695,N_26570);
xnor UO_2507 (O_2507,N_28367,N_26062);
xor UO_2508 (O_2508,N_29777,N_28260);
or UO_2509 (O_2509,N_29213,N_28013);
nor UO_2510 (O_2510,N_29632,N_29013);
or UO_2511 (O_2511,N_25313,N_25567);
xnor UO_2512 (O_2512,N_25428,N_25743);
and UO_2513 (O_2513,N_27421,N_29916);
nand UO_2514 (O_2514,N_29356,N_29310);
nand UO_2515 (O_2515,N_29659,N_25580);
and UO_2516 (O_2516,N_29720,N_26741);
nand UO_2517 (O_2517,N_28292,N_29920);
nand UO_2518 (O_2518,N_26894,N_28172);
nand UO_2519 (O_2519,N_27774,N_27777);
nand UO_2520 (O_2520,N_25626,N_27904);
nor UO_2521 (O_2521,N_29008,N_26214);
or UO_2522 (O_2522,N_25340,N_29711);
or UO_2523 (O_2523,N_27594,N_29110);
and UO_2524 (O_2524,N_26520,N_27463);
nor UO_2525 (O_2525,N_28090,N_25787);
xnor UO_2526 (O_2526,N_28993,N_29333);
xor UO_2527 (O_2527,N_25548,N_27474);
nor UO_2528 (O_2528,N_29013,N_28508);
nor UO_2529 (O_2529,N_25051,N_26838);
and UO_2530 (O_2530,N_29106,N_25759);
and UO_2531 (O_2531,N_25682,N_25275);
or UO_2532 (O_2532,N_28564,N_29674);
or UO_2533 (O_2533,N_28355,N_25282);
or UO_2534 (O_2534,N_29201,N_28389);
or UO_2535 (O_2535,N_28238,N_27505);
xnor UO_2536 (O_2536,N_28551,N_28835);
nand UO_2537 (O_2537,N_26769,N_25602);
or UO_2538 (O_2538,N_29977,N_27900);
and UO_2539 (O_2539,N_25891,N_28929);
xor UO_2540 (O_2540,N_27222,N_27621);
and UO_2541 (O_2541,N_28750,N_26552);
and UO_2542 (O_2542,N_26274,N_29310);
and UO_2543 (O_2543,N_25824,N_27774);
nand UO_2544 (O_2544,N_28928,N_26175);
xnor UO_2545 (O_2545,N_26101,N_26195);
or UO_2546 (O_2546,N_26096,N_27726);
or UO_2547 (O_2547,N_28447,N_28845);
nand UO_2548 (O_2548,N_25063,N_26812);
nor UO_2549 (O_2549,N_29933,N_25492);
or UO_2550 (O_2550,N_25953,N_25777);
and UO_2551 (O_2551,N_29193,N_28566);
and UO_2552 (O_2552,N_25756,N_28702);
or UO_2553 (O_2553,N_25797,N_28523);
nor UO_2554 (O_2554,N_25881,N_27617);
nand UO_2555 (O_2555,N_25188,N_26616);
and UO_2556 (O_2556,N_26352,N_26971);
or UO_2557 (O_2557,N_25742,N_28879);
nand UO_2558 (O_2558,N_25931,N_29194);
and UO_2559 (O_2559,N_26137,N_27435);
nor UO_2560 (O_2560,N_27851,N_29726);
nand UO_2561 (O_2561,N_25674,N_26031);
nand UO_2562 (O_2562,N_28244,N_28287);
nor UO_2563 (O_2563,N_27620,N_27243);
nor UO_2564 (O_2564,N_29627,N_25806);
and UO_2565 (O_2565,N_29353,N_25451);
or UO_2566 (O_2566,N_29596,N_29138);
nand UO_2567 (O_2567,N_25322,N_28686);
and UO_2568 (O_2568,N_25915,N_27260);
or UO_2569 (O_2569,N_29138,N_28516);
xnor UO_2570 (O_2570,N_29714,N_25161);
and UO_2571 (O_2571,N_27291,N_28330);
nand UO_2572 (O_2572,N_26809,N_29516);
xor UO_2573 (O_2573,N_28489,N_26464);
nor UO_2574 (O_2574,N_28876,N_25345);
or UO_2575 (O_2575,N_29731,N_25969);
xnor UO_2576 (O_2576,N_27739,N_28675);
or UO_2577 (O_2577,N_27570,N_26445);
xnor UO_2578 (O_2578,N_27220,N_29916);
or UO_2579 (O_2579,N_26330,N_28322);
nor UO_2580 (O_2580,N_29230,N_29039);
or UO_2581 (O_2581,N_28516,N_26801);
nor UO_2582 (O_2582,N_29340,N_25699);
and UO_2583 (O_2583,N_27623,N_26544);
nor UO_2584 (O_2584,N_25505,N_29718);
nand UO_2585 (O_2585,N_29477,N_27683);
and UO_2586 (O_2586,N_27637,N_28204);
nand UO_2587 (O_2587,N_27378,N_27407);
or UO_2588 (O_2588,N_28560,N_27436);
xnor UO_2589 (O_2589,N_28194,N_27151);
xor UO_2590 (O_2590,N_28639,N_27250);
or UO_2591 (O_2591,N_27100,N_28677);
nor UO_2592 (O_2592,N_27605,N_28806);
nor UO_2593 (O_2593,N_28676,N_25945);
xnor UO_2594 (O_2594,N_26390,N_25326);
or UO_2595 (O_2595,N_28988,N_25800);
or UO_2596 (O_2596,N_29441,N_25512);
nand UO_2597 (O_2597,N_25856,N_25986);
xor UO_2598 (O_2598,N_25323,N_28194);
nor UO_2599 (O_2599,N_28149,N_27118);
and UO_2600 (O_2600,N_26763,N_26867);
nor UO_2601 (O_2601,N_26202,N_29526);
xor UO_2602 (O_2602,N_29827,N_26999);
or UO_2603 (O_2603,N_25290,N_28783);
and UO_2604 (O_2604,N_28424,N_28338);
or UO_2605 (O_2605,N_26221,N_29373);
or UO_2606 (O_2606,N_29147,N_29535);
nor UO_2607 (O_2607,N_26152,N_25831);
and UO_2608 (O_2608,N_26394,N_25036);
or UO_2609 (O_2609,N_26177,N_29412);
xor UO_2610 (O_2610,N_25049,N_26753);
xnor UO_2611 (O_2611,N_26555,N_28763);
nor UO_2612 (O_2612,N_28055,N_28436);
nor UO_2613 (O_2613,N_29906,N_25678);
and UO_2614 (O_2614,N_29614,N_27560);
nor UO_2615 (O_2615,N_25363,N_26739);
or UO_2616 (O_2616,N_27438,N_25526);
xnor UO_2617 (O_2617,N_29487,N_28602);
nor UO_2618 (O_2618,N_26135,N_28929);
nor UO_2619 (O_2619,N_25089,N_26785);
nand UO_2620 (O_2620,N_25039,N_25537);
xor UO_2621 (O_2621,N_26807,N_28772);
or UO_2622 (O_2622,N_28005,N_29939);
and UO_2623 (O_2623,N_29383,N_28073);
or UO_2624 (O_2624,N_26619,N_28919);
nor UO_2625 (O_2625,N_27437,N_28019);
or UO_2626 (O_2626,N_27789,N_26496);
or UO_2627 (O_2627,N_29625,N_26656);
and UO_2628 (O_2628,N_26818,N_27458);
xnor UO_2629 (O_2629,N_26133,N_27413);
nand UO_2630 (O_2630,N_25864,N_28425);
nor UO_2631 (O_2631,N_28334,N_25481);
nand UO_2632 (O_2632,N_27318,N_26994);
xor UO_2633 (O_2633,N_28993,N_29058);
xor UO_2634 (O_2634,N_27332,N_27383);
and UO_2635 (O_2635,N_28281,N_25916);
nand UO_2636 (O_2636,N_29451,N_28130);
nor UO_2637 (O_2637,N_28880,N_25507);
or UO_2638 (O_2638,N_25523,N_26485);
xor UO_2639 (O_2639,N_29607,N_28742);
nand UO_2640 (O_2640,N_25483,N_29326);
and UO_2641 (O_2641,N_27788,N_28733);
nand UO_2642 (O_2642,N_27839,N_25662);
and UO_2643 (O_2643,N_26797,N_29559);
nand UO_2644 (O_2644,N_27596,N_25331);
nand UO_2645 (O_2645,N_27637,N_25935);
and UO_2646 (O_2646,N_25847,N_26225);
nand UO_2647 (O_2647,N_28669,N_28890);
and UO_2648 (O_2648,N_28550,N_26439);
or UO_2649 (O_2649,N_27583,N_29743);
and UO_2650 (O_2650,N_28219,N_25019);
or UO_2651 (O_2651,N_29528,N_28439);
xor UO_2652 (O_2652,N_25015,N_29840);
nand UO_2653 (O_2653,N_26369,N_28781);
or UO_2654 (O_2654,N_29276,N_27589);
and UO_2655 (O_2655,N_28542,N_25492);
or UO_2656 (O_2656,N_29323,N_29795);
and UO_2657 (O_2657,N_25207,N_27851);
nor UO_2658 (O_2658,N_27700,N_27681);
nand UO_2659 (O_2659,N_25933,N_28727);
or UO_2660 (O_2660,N_28083,N_29120);
xor UO_2661 (O_2661,N_27646,N_25291);
or UO_2662 (O_2662,N_25195,N_25102);
nor UO_2663 (O_2663,N_29170,N_28574);
and UO_2664 (O_2664,N_29627,N_28367);
or UO_2665 (O_2665,N_25526,N_27122);
xnor UO_2666 (O_2666,N_27553,N_25916);
and UO_2667 (O_2667,N_29175,N_27981);
and UO_2668 (O_2668,N_26657,N_26251);
xor UO_2669 (O_2669,N_29952,N_26630);
nand UO_2670 (O_2670,N_25280,N_25970);
or UO_2671 (O_2671,N_27550,N_26314);
nand UO_2672 (O_2672,N_26400,N_29444);
nand UO_2673 (O_2673,N_27136,N_25018);
or UO_2674 (O_2674,N_29595,N_25871);
nor UO_2675 (O_2675,N_26675,N_26472);
nor UO_2676 (O_2676,N_28841,N_27781);
xnor UO_2677 (O_2677,N_28180,N_27808);
xnor UO_2678 (O_2678,N_29249,N_29488);
nand UO_2679 (O_2679,N_29025,N_25811);
nor UO_2680 (O_2680,N_28143,N_26810);
nor UO_2681 (O_2681,N_28927,N_26021);
and UO_2682 (O_2682,N_26760,N_29023);
nand UO_2683 (O_2683,N_29406,N_26714);
xor UO_2684 (O_2684,N_25588,N_27333);
xor UO_2685 (O_2685,N_26863,N_29934);
or UO_2686 (O_2686,N_25287,N_25024);
and UO_2687 (O_2687,N_29076,N_28159);
nand UO_2688 (O_2688,N_27250,N_26049);
nand UO_2689 (O_2689,N_26109,N_25743);
nand UO_2690 (O_2690,N_28887,N_25803);
or UO_2691 (O_2691,N_27301,N_28682);
nand UO_2692 (O_2692,N_27984,N_26510);
nor UO_2693 (O_2693,N_27065,N_29647);
nand UO_2694 (O_2694,N_27040,N_26259);
nand UO_2695 (O_2695,N_26876,N_27347);
nand UO_2696 (O_2696,N_26978,N_26119);
or UO_2697 (O_2697,N_29046,N_26439);
or UO_2698 (O_2698,N_27769,N_25857);
nor UO_2699 (O_2699,N_26418,N_26765);
nor UO_2700 (O_2700,N_27864,N_25947);
nor UO_2701 (O_2701,N_26639,N_26677);
nor UO_2702 (O_2702,N_27461,N_25744);
or UO_2703 (O_2703,N_27690,N_27588);
xor UO_2704 (O_2704,N_26083,N_27381);
or UO_2705 (O_2705,N_28383,N_27846);
and UO_2706 (O_2706,N_28476,N_26566);
nor UO_2707 (O_2707,N_28276,N_26171);
nor UO_2708 (O_2708,N_26153,N_26329);
nor UO_2709 (O_2709,N_27436,N_29075);
or UO_2710 (O_2710,N_25364,N_25210);
nand UO_2711 (O_2711,N_25358,N_25475);
nand UO_2712 (O_2712,N_26920,N_25415);
xor UO_2713 (O_2713,N_26664,N_26585);
nand UO_2714 (O_2714,N_29928,N_27004);
or UO_2715 (O_2715,N_27390,N_26238);
or UO_2716 (O_2716,N_27562,N_28269);
xor UO_2717 (O_2717,N_25865,N_26997);
nor UO_2718 (O_2718,N_25598,N_29126);
nor UO_2719 (O_2719,N_25665,N_26055);
and UO_2720 (O_2720,N_25171,N_28163);
nand UO_2721 (O_2721,N_25840,N_29971);
nor UO_2722 (O_2722,N_26600,N_26398);
and UO_2723 (O_2723,N_28447,N_26096);
xnor UO_2724 (O_2724,N_28925,N_26571);
nor UO_2725 (O_2725,N_26356,N_27316);
nand UO_2726 (O_2726,N_26122,N_27635);
xor UO_2727 (O_2727,N_25879,N_25553);
xnor UO_2728 (O_2728,N_26782,N_25952);
nand UO_2729 (O_2729,N_29957,N_27072);
and UO_2730 (O_2730,N_29444,N_29265);
and UO_2731 (O_2731,N_29744,N_29365);
nor UO_2732 (O_2732,N_29169,N_25938);
nand UO_2733 (O_2733,N_28808,N_26072);
nand UO_2734 (O_2734,N_26830,N_25008);
nor UO_2735 (O_2735,N_27806,N_29093);
xnor UO_2736 (O_2736,N_26842,N_27107);
nand UO_2737 (O_2737,N_28016,N_29041);
xnor UO_2738 (O_2738,N_27110,N_29886);
and UO_2739 (O_2739,N_27331,N_28074);
nand UO_2740 (O_2740,N_28623,N_27175);
and UO_2741 (O_2741,N_25429,N_28138);
nand UO_2742 (O_2742,N_29319,N_26353);
and UO_2743 (O_2743,N_25361,N_25265);
or UO_2744 (O_2744,N_27354,N_29985);
xnor UO_2745 (O_2745,N_29429,N_27895);
and UO_2746 (O_2746,N_29850,N_25556);
or UO_2747 (O_2747,N_26732,N_26275);
nand UO_2748 (O_2748,N_29661,N_28558);
and UO_2749 (O_2749,N_25865,N_26746);
or UO_2750 (O_2750,N_29137,N_29523);
xor UO_2751 (O_2751,N_26283,N_28656);
or UO_2752 (O_2752,N_29500,N_28071);
nor UO_2753 (O_2753,N_28684,N_27193);
or UO_2754 (O_2754,N_25100,N_27944);
or UO_2755 (O_2755,N_26846,N_29505);
and UO_2756 (O_2756,N_26671,N_27557);
nor UO_2757 (O_2757,N_29337,N_29468);
and UO_2758 (O_2758,N_28565,N_28023);
xnor UO_2759 (O_2759,N_26113,N_25955);
or UO_2760 (O_2760,N_28469,N_29134);
nor UO_2761 (O_2761,N_29719,N_25679);
and UO_2762 (O_2762,N_25658,N_29384);
and UO_2763 (O_2763,N_25769,N_25521);
xnor UO_2764 (O_2764,N_28814,N_27579);
nor UO_2765 (O_2765,N_28778,N_29667);
xor UO_2766 (O_2766,N_27703,N_27345);
and UO_2767 (O_2767,N_28310,N_27530);
nor UO_2768 (O_2768,N_28503,N_26688);
and UO_2769 (O_2769,N_28515,N_27041);
nand UO_2770 (O_2770,N_26976,N_26774);
xnor UO_2771 (O_2771,N_25248,N_29618);
and UO_2772 (O_2772,N_25984,N_29433);
and UO_2773 (O_2773,N_29220,N_27663);
nor UO_2774 (O_2774,N_28609,N_25333);
and UO_2775 (O_2775,N_26672,N_27331);
or UO_2776 (O_2776,N_27590,N_25396);
or UO_2777 (O_2777,N_26929,N_28327);
xnor UO_2778 (O_2778,N_25323,N_25714);
nand UO_2779 (O_2779,N_28642,N_27800);
or UO_2780 (O_2780,N_28378,N_28258);
xnor UO_2781 (O_2781,N_26818,N_27222);
xor UO_2782 (O_2782,N_28393,N_25734);
xnor UO_2783 (O_2783,N_27134,N_27714);
or UO_2784 (O_2784,N_28366,N_29297);
nor UO_2785 (O_2785,N_29676,N_26540);
xor UO_2786 (O_2786,N_28157,N_28780);
nand UO_2787 (O_2787,N_26398,N_27197);
xor UO_2788 (O_2788,N_26404,N_27094);
xnor UO_2789 (O_2789,N_29250,N_25730);
or UO_2790 (O_2790,N_29413,N_25085);
nand UO_2791 (O_2791,N_28988,N_29546);
or UO_2792 (O_2792,N_28494,N_27327);
or UO_2793 (O_2793,N_28325,N_27920);
xnor UO_2794 (O_2794,N_27706,N_29940);
nand UO_2795 (O_2795,N_25982,N_28333);
or UO_2796 (O_2796,N_27670,N_25900);
or UO_2797 (O_2797,N_26382,N_26205);
nand UO_2798 (O_2798,N_27110,N_29011);
xnor UO_2799 (O_2799,N_25975,N_26603);
or UO_2800 (O_2800,N_27612,N_26540);
or UO_2801 (O_2801,N_29043,N_26782);
xor UO_2802 (O_2802,N_26322,N_25143);
or UO_2803 (O_2803,N_28006,N_25033);
or UO_2804 (O_2804,N_27736,N_27455);
nand UO_2805 (O_2805,N_26031,N_25978);
or UO_2806 (O_2806,N_26480,N_27104);
or UO_2807 (O_2807,N_29334,N_27596);
nand UO_2808 (O_2808,N_27915,N_29308);
and UO_2809 (O_2809,N_29468,N_28710);
nand UO_2810 (O_2810,N_26315,N_26023);
or UO_2811 (O_2811,N_26820,N_25281);
and UO_2812 (O_2812,N_25969,N_26854);
or UO_2813 (O_2813,N_27762,N_26896);
and UO_2814 (O_2814,N_25748,N_25942);
nand UO_2815 (O_2815,N_29495,N_26066);
xnor UO_2816 (O_2816,N_25987,N_25501);
nor UO_2817 (O_2817,N_27241,N_25059);
nand UO_2818 (O_2818,N_27867,N_25188);
or UO_2819 (O_2819,N_29409,N_25063);
and UO_2820 (O_2820,N_28022,N_29878);
nor UO_2821 (O_2821,N_25684,N_25916);
xor UO_2822 (O_2822,N_28342,N_26831);
nand UO_2823 (O_2823,N_27765,N_27820);
xnor UO_2824 (O_2824,N_26520,N_28039);
xnor UO_2825 (O_2825,N_28864,N_27955);
nor UO_2826 (O_2826,N_29571,N_27231);
nor UO_2827 (O_2827,N_27568,N_29310);
xor UO_2828 (O_2828,N_27048,N_27935);
and UO_2829 (O_2829,N_26656,N_27471);
or UO_2830 (O_2830,N_25195,N_29897);
or UO_2831 (O_2831,N_26663,N_29714);
xor UO_2832 (O_2832,N_27708,N_29647);
nor UO_2833 (O_2833,N_28399,N_28822);
nand UO_2834 (O_2834,N_29235,N_27419);
xnor UO_2835 (O_2835,N_28433,N_29529);
xnor UO_2836 (O_2836,N_26592,N_29840);
nand UO_2837 (O_2837,N_26428,N_28937);
nand UO_2838 (O_2838,N_27639,N_27538);
nor UO_2839 (O_2839,N_25684,N_27205);
xor UO_2840 (O_2840,N_27000,N_28852);
xor UO_2841 (O_2841,N_29404,N_25500);
nor UO_2842 (O_2842,N_27588,N_26463);
and UO_2843 (O_2843,N_26609,N_27178);
or UO_2844 (O_2844,N_28617,N_26102);
and UO_2845 (O_2845,N_27472,N_25055);
xnor UO_2846 (O_2846,N_29775,N_29138);
or UO_2847 (O_2847,N_29916,N_25670);
nor UO_2848 (O_2848,N_25652,N_27086);
xnor UO_2849 (O_2849,N_25690,N_29195);
and UO_2850 (O_2850,N_28914,N_27292);
nor UO_2851 (O_2851,N_25945,N_29094);
and UO_2852 (O_2852,N_26262,N_28154);
nor UO_2853 (O_2853,N_29975,N_25547);
nand UO_2854 (O_2854,N_28595,N_27209);
nand UO_2855 (O_2855,N_28273,N_29733);
and UO_2856 (O_2856,N_27285,N_25758);
xnor UO_2857 (O_2857,N_26878,N_26882);
xor UO_2858 (O_2858,N_28269,N_29556);
and UO_2859 (O_2859,N_25790,N_29340);
and UO_2860 (O_2860,N_28356,N_26865);
nor UO_2861 (O_2861,N_25407,N_29092);
xor UO_2862 (O_2862,N_26537,N_25582);
or UO_2863 (O_2863,N_28245,N_29855);
and UO_2864 (O_2864,N_25976,N_26714);
xor UO_2865 (O_2865,N_26061,N_29513);
xor UO_2866 (O_2866,N_28103,N_27510);
nand UO_2867 (O_2867,N_28239,N_29616);
nor UO_2868 (O_2868,N_27960,N_29855);
nand UO_2869 (O_2869,N_26707,N_28283);
nand UO_2870 (O_2870,N_26298,N_29723);
nand UO_2871 (O_2871,N_28418,N_27750);
nor UO_2872 (O_2872,N_26789,N_26921);
and UO_2873 (O_2873,N_29454,N_28005);
nor UO_2874 (O_2874,N_28630,N_28307);
nor UO_2875 (O_2875,N_29314,N_26115);
nand UO_2876 (O_2876,N_28017,N_29136);
xnor UO_2877 (O_2877,N_25630,N_25418);
nor UO_2878 (O_2878,N_26363,N_25689);
or UO_2879 (O_2879,N_27287,N_27708);
nand UO_2880 (O_2880,N_29501,N_27600);
xnor UO_2881 (O_2881,N_27009,N_26919);
xor UO_2882 (O_2882,N_29398,N_28624);
nand UO_2883 (O_2883,N_28567,N_26516);
xor UO_2884 (O_2884,N_25099,N_25419);
nand UO_2885 (O_2885,N_27165,N_26932);
xor UO_2886 (O_2886,N_25175,N_26037);
xor UO_2887 (O_2887,N_28391,N_25907);
nand UO_2888 (O_2888,N_25878,N_26542);
nor UO_2889 (O_2889,N_25689,N_27840);
and UO_2890 (O_2890,N_28629,N_27302);
nor UO_2891 (O_2891,N_26053,N_27237);
and UO_2892 (O_2892,N_27326,N_25864);
xnor UO_2893 (O_2893,N_25739,N_28113);
and UO_2894 (O_2894,N_26580,N_28109);
xnor UO_2895 (O_2895,N_26512,N_28318);
xnor UO_2896 (O_2896,N_26190,N_26338);
or UO_2897 (O_2897,N_25756,N_27064);
and UO_2898 (O_2898,N_26418,N_25630);
and UO_2899 (O_2899,N_28827,N_25987);
nor UO_2900 (O_2900,N_27075,N_29332);
or UO_2901 (O_2901,N_28052,N_28405);
xor UO_2902 (O_2902,N_26218,N_27749);
nand UO_2903 (O_2903,N_27376,N_28616);
nand UO_2904 (O_2904,N_26661,N_28625);
or UO_2905 (O_2905,N_29867,N_28422);
nor UO_2906 (O_2906,N_29520,N_25716);
nand UO_2907 (O_2907,N_26896,N_28731);
and UO_2908 (O_2908,N_27389,N_28482);
and UO_2909 (O_2909,N_27405,N_27539);
nand UO_2910 (O_2910,N_29157,N_26849);
nor UO_2911 (O_2911,N_29878,N_25076);
nor UO_2912 (O_2912,N_25626,N_29199);
or UO_2913 (O_2913,N_27280,N_26915);
or UO_2914 (O_2914,N_27566,N_28812);
and UO_2915 (O_2915,N_28993,N_27684);
xnor UO_2916 (O_2916,N_25147,N_25208);
and UO_2917 (O_2917,N_29825,N_26874);
and UO_2918 (O_2918,N_26106,N_25240);
xnor UO_2919 (O_2919,N_29274,N_28724);
and UO_2920 (O_2920,N_27798,N_25953);
and UO_2921 (O_2921,N_29592,N_29204);
nand UO_2922 (O_2922,N_26984,N_29637);
nand UO_2923 (O_2923,N_26562,N_26662);
nand UO_2924 (O_2924,N_27897,N_28824);
nand UO_2925 (O_2925,N_25630,N_29643);
and UO_2926 (O_2926,N_29586,N_25711);
nand UO_2927 (O_2927,N_26152,N_28045);
xnor UO_2928 (O_2928,N_26185,N_27063);
xor UO_2929 (O_2929,N_28018,N_25272);
xnor UO_2930 (O_2930,N_25392,N_25010);
xnor UO_2931 (O_2931,N_28838,N_26299);
and UO_2932 (O_2932,N_25947,N_25461);
nor UO_2933 (O_2933,N_26034,N_28906);
and UO_2934 (O_2934,N_29071,N_26925);
or UO_2935 (O_2935,N_28458,N_25341);
or UO_2936 (O_2936,N_27183,N_29208);
or UO_2937 (O_2937,N_27989,N_29012);
nor UO_2938 (O_2938,N_25454,N_29320);
or UO_2939 (O_2939,N_26581,N_26303);
or UO_2940 (O_2940,N_26455,N_28764);
nand UO_2941 (O_2941,N_25287,N_26620);
xnor UO_2942 (O_2942,N_27780,N_25758);
nor UO_2943 (O_2943,N_27580,N_28724);
nand UO_2944 (O_2944,N_27341,N_28622);
xnor UO_2945 (O_2945,N_25630,N_26179);
nor UO_2946 (O_2946,N_28761,N_28520);
nand UO_2947 (O_2947,N_29168,N_28819);
and UO_2948 (O_2948,N_29490,N_25770);
nor UO_2949 (O_2949,N_28019,N_25929);
or UO_2950 (O_2950,N_27559,N_26073);
or UO_2951 (O_2951,N_27575,N_27112);
or UO_2952 (O_2952,N_25305,N_29162);
and UO_2953 (O_2953,N_26666,N_29105);
or UO_2954 (O_2954,N_27484,N_25090);
xnor UO_2955 (O_2955,N_29380,N_29392);
nor UO_2956 (O_2956,N_28411,N_27780);
nand UO_2957 (O_2957,N_25684,N_26616);
nor UO_2958 (O_2958,N_29496,N_26752);
or UO_2959 (O_2959,N_25555,N_27359);
xnor UO_2960 (O_2960,N_25757,N_25795);
and UO_2961 (O_2961,N_27222,N_27490);
or UO_2962 (O_2962,N_25754,N_25292);
and UO_2963 (O_2963,N_25841,N_26814);
xor UO_2964 (O_2964,N_26334,N_29770);
and UO_2965 (O_2965,N_28020,N_28502);
and UO_2966 (O_2966,N_26591,N_27116);
xor UO_2967 (O_2967,N_29471,N_29562);
or UO_2968 (O_2968,N_25843,N_25689);
nor UO_2969 (O_2969,N_27306,N_25689);
nor UO_2970 (O_2970,N_26012,N_26944);
nand UO_2971 (O_2971,N_26584,N_26222);
or UO_2972 (O_2972,N_28202,N_29257);
or UO_2973 (O_2973,N_26825,N_26544);
xnor UO_2974 (O_2974,N_26233,N_25415);
or UO_2975 (O_2975,N_25542,N_26005);
nor UO_2976 (O_2976,N_27815,N_25047);
or UO_2977 (O_2977,N_25259,N_27785);
or UO_2978 (O_2978,N_25196,N_25183);
nor UO_2979 (O_2979,N_28664,N_26320);
or UO_2980 (O_2980,N_25034,N_29135);
xor UO_2981 (O_2981,N_29180,N_26287);
xor UO_2982 (O_2982,N_27668,N_29601);
nand UO_2983 (O_2983,N_26062,N_25526);
nor UO_2984 (O_2984,N_25287,N_28594);
nand UO_2985 (O_2985,N_29522,N_29396);
nand UO_2986 (O_2986,N_27499,N_27771);
nand UO_2987 (O_2987,N_25274,N_25457);
nand UO_2988 (O_2988,N_26550,N_25867);
xor UO_2989 (O_2989,N_27350,N_27207);
nand UO_2990 (O_2990,N_25012,N_29918);
and UO_2991 (O_2991,N_26935,N_26790);
nand UO_2992 (O_2992,N_25601,N_25402);
or UO_2993 (O_2993,N_28437,N_26450);
and UO_2994 (O_2994,N_26170,N_29127);
and UO_2995 (O_2995,N_29547,N_25143);
nand UO_2996 (O_2996,N_28711,N_25296);
nand UO_2997 (O_2997,N_26453,N_28068);
nor UO_2998 (O_2998,N_25050,N_27261);
nand UO_2999 (O_2999,N_29372,N_26783);
nand UO_3000 (O_3000,N_27467,N_25379);
and UO_3001 (O_3001,N_29622,N_29686);
or UO_3002 (O_3002,N_26879,N_25900);
xnor UO_3003 (O_3003,N_27569,N_27911);
nor UO_3004 (O_3004,N_28230,N_26636);
and UO_3005 (O_3005,N_27188,N_28145);
nor UO_3006 (O_3006,N_28721,N_29223);
or UO_3007 (O_3007,N_25416,N_28099);
nor UO_3008 (O_3008,N_29919,N_28727);
or UO_3009 (O_3009,N_26977,N_26532);
and UO_3010 (O_3010,N_29548,N_27968);
and UO_3011 (O_3011,N_29183,N_29601);
or UO_3012 (O_3012,N_29706,N_25820);
xor UO_3013 (O_3013,N_29772,N_25743);
nand UO_3014 (O_3014,N_27861,N_29120);
xor UO_3015 (O_3015,N_25894,N_27414);
xnor UO_3016 (O_3016,N_25412,N_25592);
xnor UO_3017 (O_3017,N_27629,N_28159);
and UO_3018 (O_3018,N_27928,N_29081);
and UO_3019 (O_3019,N_25157,N_25227);
xnor UO_3020 (O_3020,N_26868,N_25723);
or UO_3021 (O_3021,N_25935,N_27109);
nor UO_3022 (O_3022,N_28841,N_28015);
and UO_3023 (O_3023,N_25652,N_29441);
and UO_3024 (O_3024,N_29705,N_26507);
or UO_3025 (O_3025,N_25017,N_29056);
nand UO_3026 (O_3026,N_27232,N_25670);
xor UO_3027 (O_3027,N_25156,N_29320);
nor UO_3028 (O_3028,N_26294,N_29665);
nand UO_3029 (O_3029,N_28648,N_26274);
or UO_3030 (O_3030,N_26267,N_25029);
xnor UO_3031 (O_3031,N_29149,N_28268);
nor UO_3032 (O_3032,N_27105,N_25685);
nand UO_3033 (O_3033,N_29023,N_28502);
nor UO_3034 (O_3034,N_27249,N_27411);
xor UO_3035 (O_3035,N_26155,N_25960);
and UO_3036 (O_3036,N_27481,N_26690);
nor UO_3037 (O_3037,N_26931,N_28674);
xor UO_3038 (O_3038,N_25306,N_25146);
or UO_3039 (O_3039,N_29481,N_28533);
nor UO_3040 (O_3040,N_29058,N_29054);
xnor UO_3041 (O_3041,N_27429,N_25818);
xor UO_3042 (O_3042,N_28357,N_26643);
or UO_3043 (O_3043,N_28860,N_28185);
and UO_3044 (O_3044,N_26206,N_29562);
and UO_3045 (O_3045,N_28488,N_25879);
nand UO_3046 (O_3046,N_29130,N_25817);
or UO_3047 (O_3047,N_29265,N_27193);
and UO_3048 (O_3048,N_27527,N_27025);
nand UO_3049 (O_3049,N_28706,N_28440);
or UO_3050 (O_3050,N_26328,N_26621);
and UO_3051 (O_3051,N_27977,N_28138);
or UO_3052 (O_3052,N_29765,N_28929);
nand UO_3053 (O_3053,N_25933,N_27838);
nor UO_3054 (O_3054,N_28001,N_25590);
nand UO_3055 (O_3055,N_29583,N_28865);
and UO_3056 (O_3056,N_25516,N_25011);
and UO_3057 (O_3057,N_26272,N_27708);
or UO_3058 (O_3058,N_28317,N_29254);
or UO_3059 (O_3059,N_28909,N_26742);
or UO_3060 (O_3060,N_29603,N_25308);
nand UO_3061 (O_3061,N_27653,N_27263);
nor UO_3062 (O_3062,N_28927,N_27307);
or UO_3063 (O_3063,N_28099,N_25981);
nand UO_3064 (O_3064,N_29205,N_27668);
nor UO_3065 (O_3065,N_29168,N_26832);
or UO_3066 (O_3066,N_26070,N_28987);
nor UO_3067 (O_3067,N_27534,N_26510);
nand UO_3068 (O_3068,N_29470,N_29643);
nand UO_3069 (O_3069,N_28172,N_26007);
nand UO_3070 (O_3070,N_28535,N_27068);
nor UO_3071 (O_3071,N_27020,N_27367);
nor UO_3072 (O_3072,N_27308,N_26788);
and UO_3073 (O_3073,N_26172,N_28468);
or UO_3074 (O_3074,N_27993,N_26118);
or UO_3075 (O_3075,N_26527,N_25786);
nand UO_3076 (O_3076,N_29404,N_27219);
and UO_3077 (O_3077,N_28395,N_29167);
or UO_3078 (O_3078,N_26319,N_27898);
and UO_3079 (O_3079,N_28995,N_27499);
xor UO_3080 (O_3080,N_25056,N_27881);
or UO_3081 (O_3081,N_29864,N_26709);
or UO_3082 (O_3082,N_28476,N_27343);
nor UO_3083 (O_3083,N_26356,N_29515);
nand UO_3084 (O_3084,N_28495,N_25629);
xnor UO_3085 (O_3085,N_29766,N_29281);
nand UO_3086 (O_3086,N_27350,N_25774);
nand UO_3087 (O_3087,N_29138,N_28725);
nor UO_3088 (O_3088,N_27007,N_28035);
nand UO_3089 (O_3089,N_27802,N_28700);
nand UO_3090 (O_3090,N_25467,N_29150);
or UO_3091 (O_3091,N_29397,N_29242);
nand UO_3092 (O_3092,N_28825,N_26308);
nand UO_3093 (O_3093,N_28322,N_25422);
and UO_3094 (O_3094,N_25123,N_27166);
nand UO_3095 (O_3095,N_25052,N_25863);
and UO_3096 (O_3096,N_28746,N_28398);
nand UO_3097 (O_3097,N_29372,N_28280);
nor UO_3098 (O_3098,N_28085,N_29390);
and UO_3099 (O_3099,N_28346,N_28344);
and UO_3100 (O_3100,N_27610,N_27288);
nand UO_3101 (O_3101,N_27821,N_27488);
xnor UO_3102 (O_3102,N_26963,N_26210);
nor UO_3103 (O_3103,N_28160,N_27468);
xor UO_3104 (O_3104,N_25884,N_25010);
and UO_3105 (O_3105,N_25401,N_28259);
nor UO_3106 (O_3106,N_25560,N_25839);
and UO_3107 (O_3107,N_27509,N_26014);
nand UO_3108 (O_3108,N_29734,N_25149);
or UO_3109 (O_3109,N_27906,N_28065);
and UO_3110 (O_3110,N_25753,N_29654);
or UO_3111 (O_3111,N_28360,N_26664);
and UO_3112 (O_3112,N_25701,N_27569);
and UO_3113 (O_3113,N_27600,N_27608);
xor UO_3114 (O_3114,N_25871,N_25942);
or UO_3115 (O_3115,N_26830,N_29178);
and UO_3116 (O_3116,N_26600,N_27686);
nor UO_3117 (O_3117,N_27724,N_27212);
xnor UO_3118 (O_3118,N_28023,N_27527);
nand UO_3119 (O_3119,N_25325,N_29750);
nor UO_3120 (O_3120,N_28282,N_28911);
nand UO_3121 (O_3121,N_28698,N_28311);
nand UO_3122 (O_3122,N_25169,N_25825);
and UO_3123 (O_3123,N_26978,N_26648);
and UO_3124 (O_3124,N_25343,N_29005);
or UO_3125 (O_3125,N_28914,N_28457);
xor UO_3126 (O_3126,N_25706,N_29095);
xnor UO_3127 (O_3127,N_28468,N_27596);
nor UO_3128 (O_3128,N_29166,N_25245);
xor UO_3129 (O_3129,N_28750,N_28555);
nand UO_3130 (O_3130,N_25754,N_28819);
or UO_3131 (O_3131,N_29153,N_28059);
nand UO_3132 (O_3132,N_25635,N_27369);
or UO_3133 (O_3133,N_25182,N_26255);
nor UO_3134 (O_3134,N_29145,N_26214);
nand UO_3135 (O_3135,N_28897,N_26032);
and UO_3136 (O_3136,N_26391,N_29837);
xnor UO_3137 (O_3137,N_27708,N_28036);
and UO_3138 (O_3138,N_25464,N_27942);
and UO_3139 (O_3139,N_28620,N_27743);
nor UO_3140 (O_3140,N_28625,N_28970);
and UO_3141 (O_3141,N_29224,N_26372);
nor UO_3142 (O_3142,N_26227,N_28033);
xor UO_3143 (O_3143,N_27483,N_26696);
xnor UO_3144 (O_3144,N_26174,N_29499);
or UO_3145 (O_3145,N_26256,N_25159);
or UO_3146 (O_3146,N_28870,N_26615);
nor UO_3147 (O_3147,N_29037,N_26115);
xnor UO_3148 (O_3148,N_29696,N_28903);
and UO_3149 (O_3149,N_29165,N_26461);
nand UO_3150 (O_3150,N_29366,N_29403);
xor UO_3151 (O_3151,N_29634,N_29537);
and UO_3152 (O_3152,N_25706,N_28184);
nor UO_3153 (O_3153,N_27188,N_25274);
or UO_3154 (O_3154,N_29030,N_26633);
xor UO_3155 (O_3155,N_26869,N_27835);
xnor UO_3156 (O_3156,N_29258,N_28563);
and UO_3157 (O_3157,N_29440,N_26788);
nand UO_3158 (O_3158,N_29626,N_28695);
xor UO_3159 (O_3159,N_26011,N_29956);
xnor UO_3160 (O_3160,N_26033,N_28333);
nand UO_3161 (O_3161,N_28818,N_28935);
nor UO_3162 (O_3162,N_28815,N_28624);
nor UO_3163 (O_3163,N_26205,N_28627);
xor UO_3164 (O_3164,N_28208,N_29753);
and UO_3165 (O_3165,N_29440,N_28998);
nor UO_3166 (O_3166,N_25912,N_29540);
nor UO_3167 (O_3167,N_26168,N_26208);
nand UO_3168 (O_3168,N_25990,N_25081);
xor UO_3169 (O_3169,N_25225,N_27557);
nand UO_3170 (O_3170,N_26970,N_28236);
and UO_3171 (O_3171,N_28793,N_29425);
nor UO_3172 (O_3172,N_25440,N_27424);
nor UO_3173 (O_3173,N_29136,N_26119);
or UO_3174 (O_3174,N_26411,N_25027);
xor UO_3175 (O_3175,N_27464,N_25151);
nand UO_3176 (O_3176,N_26082,N_25649);
xor UO_3177 (O_3177,N_28994,N_26589);
xor UO_3178 (O_3178,N_28533,N_26458);
xor UO_3179 (O_3179,N_25929,N_26434);
xor UO_3180 (O_3180,N_26384,N_29704);
nor UO_3181 (O_3181,N_29319,N_27624);
nor UO_3182 (O_3182,N_26955,N_26510);
nand UO_3183 (O_3183,N_28804,N_25490);
nand UO_3184 (O_3184,N_29726,N_28662);
and UO_3185 (O_3185,N_26728,N_25105);
nor UO_3186 (O_3186,N_26610,N_26745);
nor UO_3187 (O_3187,N_27660,N_26610);
xor UO_3188 (O_3188,N_29425,N_29471);
or UO_3189 (O_3189,N_29477,N_28598);
and UO_3190 (O_3190,N_25828,N_25675);
xor UO_3191 (O_3191,N_25780,N_27069);
nor UO_3192 (O_3192,N_27386,N_29457);
xor UO_3193 (O_3193,N_28268,N_26090);
nand UO_3194 (O_3194,N_26111,N_28872);
or UO_3195 (O_3195,N_25747,N_26917);
or UO_3196 (O_3196,N_26876,N_29470);
or UO_3197 (O_3197,N_29970,N_25857);
nor UO_3198 (O_3198,N_25807,N_25540);
xnor UO_3199 (O_3199,N_26746,N_25171);
nand UO_3200 (O_3200,N_28381,N_29019);
and UO_3201 (O_3201,N_26135,N_26683);
and UO_3202 (O_3202,N_29253,N_25710);
xor UO_3203 (O_3203,N_28308,N_26307);
xnor UO_3204 (O_3204,N_28144,N_27008);
and UO_3205 (O_3205,N_29574,N_25664);
nor UO_3206 (O_3206,N_27810,N_27430);
nor UO_3207 (O_3207,N_28695,N_26957);
and UO_3208 (O_3208,N_26861,N_29208);
or UO_3209 (O_3209,N_29071,N_27072);
nand UO_3210 (O_3210,N_26389,N_29389);
nand UO_3211 (O_3211,N_28619,N_26686);
xor UO_3212 (O_3212,N_29250,N_26926);
nor UO_3213 (O_3213,N_29789,N_26536);
nor UO_3214 (O_3214,N_29102,N_28149);
and UO_3215 (O_3215,N_28203,N_29517);
or UO_3216 (O_3216,N_29271,N_28951);
or UO_3217 (O_3217,N_26691,N_26422);
or UO_3218 (O_3218,N_29186,N_25029);
or UO_3219 (O_3219,N_27861,N_26853);
xor UO_3220 (O_3220,N_28964,N_29617);
xnor UO_3221 (O_3221,N_29310,N_26326);
nor UO_3222 (O_3222,N_26623,N_29319);
xnor UO_3223 (O_3223,N_29834,N_27112);
or UO_3224 (O_3224,N_28955,N_26735);
and UO_3225 (O_3225,N_26655,N_26604);
xnor UO_3226 (O_3226,N_29437,N_26227);
nand UO_3227 (O_3227,N_25829,N_26444);
or UO_3228 (O_3228,N_29277,N_28775);
nor UO_3229 (O_3229,N_26933,N_26385);
xnor UO_3230 (O_3230,N_26824,N_26420);
or UO_3231 (O_3231,N_25155,N_29142);
xor UO_3232 (O_3232,N_28885,N_27511);
or UO_3233 (O_3233,N_27506,N_28435);
and UO_3234 (O_3234,N_28705,N_28708);
and UO_3235 (O_3235,N_27838,N_27383);
xor UO_3236 (O_3236,N_25183,N_27991);
and UO_3237 (O_3237,N_26679,N_26218);
or UO_3238 (O_3238,N_26231,N_27861);
or UO_3239 (O_3239,N_28758,N_27191);
or UO_3240 (O_3240,N_25822,N_28594);
and UO_3241 (O_3241,N_29143,N_25545);
nand UO_3242 (O_3242,N_25930,N_29136);
nor UO_3243 (O_3243,N_29726,N_28630);
and UO_3244 (O_3244,N_26224,N_29331);
nor UO_3245 (O_3245,N_27218,N_28089);
and UO_3246 (O_3246,N_27713,N_26403);
or UO_3247 (O_3247,N_27293,N_25794);
nand UO_3248 (O_3248,N_29050,N_28651);
or UO_3249 (O_3249,N_26552,N_28548);
nand UO_3250 (O_3250,N_29768,N_26330);
nand UO_3251 (O_3251,N_26614,N_27691);
xor UO_3252 (O_3252,N_29216,N_29108);
nand UO_3253 (O_3253,N_28377,N_29086);
nor UO_3254 (O_3254,N_25672,N_29973);
nor UO_3255 (O_3255,N_29310,N_25314);
nand UO_3256 (O_3256,N_26616,N_25197);
xor UO_3257 (O_3257,N_29275,N_25662);
and UO_3258 (O_3258,N_29154,N_25626);
nand UO_3259 (O_3259,N_27843,N_28027);
xor UO_3260 (O_3260,N_29274,N_29367);
xnor UO_3261 (O_3261,N_25562,N_29696);
nor UO_3262 (O_3262,N_29259,N_28747);
nand UO_3263 (O_3263,N_29226,N_26732);
nor UO_3264 (O_3264,N_25586,N_26445);
nand UO_3265 (O_3265,N_25878,N_29971);
nor UO_3266 (O_3266,N_25594,N_26160);
nor UO_3267 (O_3267,N_25527,N_25993);
nor UO_3268 (O_3268,N_27765,N_25670);
nand UO_3269 (O_3269,N_26485,N_28055);
nand UO_3270 (O_3270,N_27969,N_27979);
nor UO_3271 (O_3271,N_27839,N_26986);
or UO_3272 (O_3272,N_26273,N_25628);
xnor UO_3273 (O_3273,N_26370,N_26814);
xor UO_3274 (O_3274,N_28649,N_27950);
nand UO_3275 (O_3275,N_28964,N_26915);
xnor UO_3276 (O_3276,N_26312,N_26500);
nand UO_3277 (O_3277,N_28091,N_29849);
xnor UO_3278 (O_3278,N_25769,N_25935);
and UO_3279 (O_3279,N_28187,N_25617);
and UO_3280 (O_3280,N_26031,N_28815);
nand UO_3281 (O_3281,N_28147,N_28547);
and UO_3282 (O_3282,N_29004,N_26942);
xor UO_3283 (O_3283,N_25665,N_29328);
or UO_3284 (O_3284,N_26984,N_27269);
xor UO_3285 (O_3285,N_26827,N_28013);
nor UO_3286 (O_3286,N_27504,N_28550);
nand UO_3287 (O_3287,N_26982,N_26790);
and UO_3288 (O_3288,N_26100,N_28803);
and UO_3289 (O_3289,N_29956,N_25907);
xnor UO_3290 (O_3290,N_26314,N_27015);
or UO_3291 (O_3291,N_29520,N_27970);
xor UO_3292 (O_3292,N_29680,N_25144);
or UO_3293 (O_3293,N_25621,N_25787);
and UO_3294 (O_3294,N_29895,N_29935);
nor UO_3295 (O_3295,N_28569,N_29784);
nand UO_3296 (O_3296,N_29902,N_25429);
xnor UO_3297 (O_3297,N_28029,N_25641);
nand UO_3298 (O_3298,N_25300,N_27760);
and UO_3299 (O_3299,N_27419,N_27151);
nand UO_3300 (O_3300,N_29099,N_26603);
or UO_3301 (O_3301,N_29007,N_26450);
xor UO_3302 (O_3302,N_25477,N_28388);
nor UO_3303 (O_3303,N_26680,N_28024);
or UO_3304 (O_3304,N_27874,N_27224);
and UO_3305 (O_3305,N_26038,N_27788);
or UO_3306 (O_3306,N_25382,N_27096);
and UO_3307 (O_3307,N_27180,N_28920);
xor UO_3308 (O_3308,N_28579,N_28385);
xnor UO_3309 (O_3309,N_27138,N_28985);
xnor UO_3310 (O_3310,N_29953,N_25273);
and UO_3311 (O_3311,N_26403,N_25184);
or UO_3312 (O_3312,N_28239,N_27755);
and UO_3313 (O_3313,N_26003,N_28551);
nor UO_3314 (O_3314,N_29759,N_25884);
nand UO_3315 (O_3315,N_28629,N_29984);
nand UO_3316 (O_3316,N_26606,N_28597);
nor UO_3317 (O_3317,N_26246,N_26100);
and UO_3318 (O_3318,N_28696,N_29182);
xor UO_3319 (O_3319,N_29621,N_26503);
nand UO_3320 (O_3320,N_25793,N_28858);
or UO_3321 (O_3321,N_27999,N_27244);
nor UO_3322 (O_3322,N_26788,N_25291);
nand UO_3323 (O_3323,N_25916,N_26364);
nor UO_3324 (O_3324,N_25657,N_28090);
xor UO_3325 (O_3325,N_28222,N_27097);
or UO_3326 (O_3326,N_29310,N_25594);
or UO_3327 (O_3327,N_27677,N_28126);
or UO_3328 (O_3328,N_25840,N_29175);
and UO_3329 (O_3329,N_27701,N_29727);
or UO_3330 (O_3330,N_26449,N_28238);
nor UO_3331 (O_3331,N_27195,N_26203);
nor UO_3332 (O_3332,N_28992,N_26281);
nand UO_3333 (O_3333,N_27928,N_28102);
xnor UO_3334 (O_3334,N_29009,N_28692);
nor UO_3335 (O_3335,N_26491,N_27392);
nand UO_3336 (O_3336,N_26647,N_28110);
xor UO_3337 (O_3337,N_25653,N_25647);
nor UO_3338 (O_3338,N_27718,N_28419);
and UO_3339 (O_3339,N_28177,N_25014);
nor UO_3340 (O_3340,N_28718,N_26482);
or UO_3341 (O_3341,N_28051,N_27216);
nor UO_3342 (O_3342,N_28104,N_28559);
and UO_3343 (O_3343,N_26099,N_27187);
nor UO_3344 (O_3344,N_28594,N_26172);
or UO_3345 (O_3345,N_29703,N_25199);
nand UO_3346 (O_3346,N_26665,N_26757);
nor UO_3347 (O_3347,N_25248,N_25412);
or UO_3348 (O_3348,N_27695,N_25185);
nor UO_3349 (O_3349,N_26503,N_27572);
nor UO_3350 (O_3350,N_29530,N_28328);
xor UO_3351 (O_3351,N_27581,N_25572);
and UO_3352 (O_3352,N_28507,N_27046);
xor UO_3353 (O_3353,N_26505,N_25800);
xor UO_3354 (O_3354,N_29448,N_29852);
and UO_3355 (O_3355,N_29431,N_29590);
xor UO_3356 (O_3356,N_29275,N_28143);
or UO_3357 (O_3357,N_27923,N_27893);
xnor UO_3358 (O_3358,N_25032,N_25396);
nor UO_3359 (O_3359,N_26872,N_27761);
nor UO_3360 (O_3360,N_25861,N_29484);
or UO_3361 (O_3361,N_26436,N_28347);
nand UO_3362 (O_3362,N_28915,N_26957);
and UO_3363 (O_3363,N_25590,N_25946);
nand UO_3364 (O_3364,N_29577,N_25871);
xor UO_3365 (O_3365,N_26427,N_25783);
nor UO_3366 (O_3366,N_27782,N_29875);
nand UO_3367 (O_3367,N_26780,N_26166);
or UO_3368 (O_3368,N_25539,N_28498);
xnor UO_3369 (O_3369,N_27911,N_25346);
and UO_3370 (O_3370,N_28582,N_26453);
and UO_3371 (O_3371,N_26571,N_27627);
nor UO_3372 (O_3372,N_28093,N_29573);
xor UO_3373 (O_3373,N_28740,N_27044);
or UO_3374 (O_3374,N_29137,N_28287);
nor UO_3375 (O_3375,N_29813,N_26879);
or UO_3376 (O_3376,N_25662,N_27545);
nor UO_3377 (O_3377,N_28412,N_25972);
and UO_3378 (O_3378,N_26273,N_29791);
and UO_3379 (O_3379,N_25327,N_29179);
xnor UO_3380 (O_3380,N_27852,N_26132);
and UO_3381 (O_3381,N_26279,N_29278);
and UO_3382 (O_3382,N_27052,N_28509);
nor UO_3383 (O_3383,N_28117,N_28612);
nor UO_3384 (O_3384,N_25348,N_27251);
nor UO_3385 (O_3385,N_28319,N_26758);
nor UO_3386 (O_3386,N_28487,N_25624);
or UO_3387 (O_3387,N_28443,N_28278);
nor UO_3388 (O_3388,N_25648,N_29715);
nand UO_3389 (O_3389,N_25319,N_25051);
and UO_3390 (O_3390,N_29569,N_26715);
nor UO_3391 (O_3391,N_26618,N_29434);
xnor UO_3392 (O_3392,N_26200,N_27642);
xnor UO_3393 (O_3393,N_25547,N_25015);
nand UO_3394 (O_3394,N_27593,N_27784);
xnor UO_3395 (O_3395,N_27562,N_29875);
and UO_3396 (O_3396,N_28354,N_28118);
or UO_3397 (O_3397,N_29438,N_29874);
and UO_3398 (O_3398,N_29693,N_29513);
nand UO_3399 (O_3399,N_27433,N_26263);
nor UO_3400 (O_3400,N_27072,N_27804);
and UO_3401 (O_3401,N_25908,N_25609);
or UO_3402 (O_3402,N_25675,N_28083);
xor UO_3403 (O_3403,N_27408,N_29502);
or UO_3404 (O_3404,N_27050,N_29461);
or UO_3405 (O_3405,N_28434,N_27088);
nor UO_3406 (O_3406,N_25443,N_25602);
and UO_3407 (O_3407,N_26829,N_26253);
and UO_3408 (O_3408,N_26514,N_25563);
nand UO_3409 (O_3409,N_26847,N_28745);
nor UO_3410 (O_3410,N_29827,N_25767);
nand UO_3411 (O_3411,N_25765,N_26890);
xor UO_3412 (O_3412,N_26516,N_25172);
nor UO_3413 (O_3413,N_26436,N_25279);
xor UO_3414 (O_3414,N_29172,N_26405);
nand UO_3415 (O_3415,N_28417,N_27850);
or UO_3416 (O_3416,N_26966,N_28956);
nand UO_3417 (O_3417,N_27857,N_25155);
and UO_3418 (O_3418,N_28275,N_29143);
or UO_3419 (O_3419,N_29686,N_29901);
nand UO_3420 (O_3420,N_25546,N_25714);
xor UO_3421 (O_3421,N_29712,N_26976);
or UO_3422 (O_3422,N_25397,N_29724);
and UO_3423 (O_3423,N_25189,N_25760);
nand UO_3424 (O_3424,N_29373,N_29789);
nand UO_3425 (O_3425,N_28847,N_28135);
nand UO_3426 (O_3426,N_29895,N_26895);
nor UO_3427 (O_3427,N_29617,N_26553);
nor UO_3428 (O_3428,N_29993,N_26953);
nor UO_3429 (O_3429,N_29794,N_27523);
nand UO_3430 (O_3430,N_26183,N_27011);
and UO_3431 (O_3431,N_29021,N_26413);
xor UO_3432 (O_3432,N_27561,N_28759);
and UO_3433 (O_3433,N_28030,N_25030);
or UO_3434 (O_3434,N_25147,N_26306);
nand UO_3435 (O_3435,N_29933,N_27786);
xnor UO_3436 (O_3436,N_29651,N_27933);
and UO_3437 (O_3437,N_28746,N_26688);
and UO_3438 (O_3438,N_25776,N_25789);
or UO_3439 (O_3439,N_28402,N_26645);
and UO_3440 (O_3440,N_28033,N_26255);
and UO_3441 (O_3441,N_25607,N_29633);
xnor UO_3442 (O_3442,N_26674,N_28778);
xor UO_3443 (O_3443,N_28280,N_29398);
nand UO_3444 (O_3444,N_27593,N_29992);
and UO_3445 (O_3445,N_26817,N_26708);
nand UO_3446 (O_3446,N_26730,N_29683);
or UO_3447 (O_3447,N_29319,N_25210);
nand UO_3448 (O_3448,N_29544,N_28374);
or UO_3449 (O_3449,N_27675,N_26793);
or UO_3450 (O_3450,N_25626,N_25718);
xor UO_3451 (O_3451,N_26759,N_29148);
nor UO_3452 (O_3452,N_29011,N_27108);
and UO_3453 (O_3453,N_27343,N_29029);
or UO_3454 (O_3454,N_27410,N_28385);
or UO_3455 (O_3455,N_26594,N_25707);
xor UO_3456 (O_3456,N_25637,N_25819);
nand UO_3457 (O_3457,N_26780,N_25374);
nand UO_3458 (O_3458,N_29009,N_26414);
nand UO_3459 (O_3459,N_26714,N_26469);
xnor UO_3460 (O_3460,N_26816,N_26643);
nor UO_3461 (O_3461,N_29459,N_27392);
or UO_3462 (O_3462,N_28346,N_28964);
nand UO_3463 (O_3463,N_27528,N_29816);
nand UO_3464 (O_3464,N_29282,N_25469);
nand UO_3465 (O_3465,N_25493,N_25907);
xnor UO_3466 (O_3466,N_25718,N_25528);
and UO_3467 (O_3467,N_29747,N_26593);
and UO_3468 (O_3468,N_25782,N_26578);
nand UO_3469 (O_3469,N_29070,N_25498);
or UO_3470 (O_3470,N_28973,N_25925);
nor UO_3471 (O_3471,N_28426,N_28980);
xor UO_3472 (O_3472,N_28684,N_29291);
xor UO_3473 (O_3473,N_25064,N_25104);
nand UO_3474 (O_3474,N_25772,N_26533);
and UO_3475 (O_3475,N_26174,N_26731);
or UO_3476 (O_3476,N_27761,N_28972);
nor UO_3477 (O_3477,N_27261,N_27582);
nor UO_3478 (O_3478,N_29693,N_29381);
and UO_3479 (O_3479,N_29619,N_29351);
xnor UO_3480 (O_3480,N_26253,N_29758);
nor UO_3481 (O_3481,N_25733,N_28623);
nand UO_3482 (O_3482,N_26854,N_28438);
and UO_3483 (O_3483,N_29613,N_27969);
or UO_3484 (O_3484,N_27392,N_25453);
xnor UO_3485 (O_3485,N_26923,N_25082);
nor UO_3486 (O_3486,N_26127,N_26704);
nand UO_3487 (O_3487,N_28095,N_27566);
nand UO_3488 (O_3488,N_26922,N_27936);
and UO_3489 (O_3489,N_27480,N_26417);
nor UO_3490 (O_3490,N_28637,N_28423);
or UO_3491 (O_3491,N_25119,N_29832);
or UO_3492 (O_3492,N_26676,N_26266);
nor UO_3493 (O_3493,N_28207,N_25642);
and UO_3494 (O_3494,N_25033,N_26446);
xor UO_3495 (O_3495,N_28949,N_26649);
nand UO_3496 (O_3496,N_26570,N_25997);
xnor UO_3497 (O_3497,N_29533,N_28941);
or UO_3498 (O_3498,N_26962,N_28459);
xor UO_3499 (O_3499,N_26814,N_28115);
endmodule